module basic_5000_50000_5000_5_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_2550,In_3379);
xnor U1 (N_1,In_4844,In_2206);
or U2 (N_2,In_1343,In_3166);
nor U3 (N_3,In_1926,In_3943);
or U4 (N_4,In_2121,In_1607);
or U5 (N_5,In_836,In_47);
and U6 (N_6,In_2447,In_4040);
xnor U7 (N_7,In_813,In_3447);
xor U8 (N_8,In_2053,In_2980);
or U9 (N_9,In_760,In_1042);
nor U10 (N_10,In_1157,In_2988);
nor U11 (N_11,In_2955,In_2004);
or U12 (N_12,In_3543,In_2355);
or U13 (N_13,In_3616,In_3392);
or U14 (N_14,In_292,In_136);
nor U15 (N_15,In_3830,In_1046);
nor U16 (N_16,In_243,In_1663);
nor U17 (N_17,In_1862,In_1187);
or U18 (N_18,In_4824,In_2630);
nand U19 (N_19,In_307,In_3787);
xnor U20 (N_20,In_2556,In_1714);
nor U21 (N_21,In_1296,In_1743);
nor U22 (N_22,In_1078,In_95);
nand U23 (N_23,In_601,In_4278);
or U24 (N_24,In_4447,In_758);
or U25 (N_25,In_4105,In_2962);
or U26 (N_26,In_2256,In_1589);
nand U27 (N_27,In_1949,In_174);
nor U28 (N_28,In_3007,In_947);
xor U29 (N_29,In_1581,In_1065);
xor U30 (N_30,In_1456,In_2932);
nor U31 (N_31,In_271,In_2662);
nand U32 (N_32,In_1236,In_4308);
or U33 (N_33,In_157,In_3280);
nand U34 (N_34,In_4221,In_3278);
nor U35 (N_35,In_1737,In_837);
nand U36 (N_36,In_3844,In_3937);
or U37 (N_37,In_2161,In_2003);
and U38 (N_38,In_2888,In_1326);
or U39 (N_39,In_2189,In_516);
nor U40 (N_40,In_3018,In_1339);
and U41 (N_41,In_4244,In_3919);
nand U42 (N_42,In_4056,In_4904);
xnor U43 (N_43,In_4047,In_860);
or U44 (N_44,In_3396,In_218);
or U45 (N_45,In_835,In_187);
xnor U46 (N_46,In_2611,In_1040);
nand U47 (N_47,In_4929,In_2387);
or U48 (N_48,In_4906,In_3870);
nand U49 (N_49,In_2947,In_2158);
or U50 (N_50,In_1508,In_2261);
and U51 (N_51,In_3227,In_4629);
and U52 (N_52,In_4184,In_2034);
nor U53 (N_53,In_2529,In_4551);
and U54 (N_54,In_229,In_4006);
nand U55 (N_55,In_2324,In_507);
xor U56 (N_56,In_3221,In_1869);
nor U57 (N_57,In_2996,In_428);
nor U58 (N_58,In_2184,In_1132);
nor U59 (N_59,In_2166,In_4375);
and U60 (N_60,In_968,In_816);
nor U61 (N_61,In_4924,In_4104);
nand U62 (N_62,In_2558,In_723);
nand U63 (N_63,In_955,In_1230);
xor U64 (N_64,In_1190,In_3667);
nor U65 (N_65,In_3001,In_4572);
or U66 (N_66,In_1016,In_2636);
nor U67 (N_67,In_4555,In_2938);
or U68 (N_68,In_3188,In_4579);
nand U69 (N_69,In_3163,In_636);
nand U70 (N_70,In_3359,In_4661);
nor U71 (N_71,In_4251,In_421);
nor U72 (N_72,In_1556,In_4949);
nor U73 (N_73,In_2594,In_3970);
and U74 (N_74,In_1590,In_4614);
nand U75 (N_75,In_2879,In_1734);
nor U76 (N_76,In_2358,In_4591);
nor U77 (N_77,In_2942,In_3313);
nand U78 (N_78,In_683,In_4806);
nand U79 (N_79,In_3495,In_253);
and U80 (N_80,In_252,In_146);
nand U81 (N_81,In_2647,In_1308);
nor U82 (N_82,In_4475,In_3631);
or U83 (N_83,In_3269,In_2212);
nand U84 (N_84,In_2840,In_3211);
nor U85 (N_85,In_4205,In_4137);
nor U86 (N_86,In_2799,In_744);
and U87 (N_87,In_2518,In_3663);
and U88 (N_88,In_4322,In_4708);
or U89 (N_89,In_333,In_2804);
or U90 (N_90,In_665,In_4074);
and U91 (N_91,In_1200,In_1971);
nand U92 (N_92,In_4073,In_2240);
or U93 (N_93,In_4165,In_2849);
or U94 (N_94,In_807,In_1282);
nand U95 (N_95,In_2390,In_4937);
nand U96 (N_96,In_2716,In_4717);
and U97 (N_97,In_1359,In_499);
and U98 (N_98,In_2234,In_4881);
nor U99 (N_99,In_2595,In_535);
or U100 (N_100,In_2743,In_200);
and U101 (N_101,In_2510,In_1863);
nand U102 (N_102,In_315,In_2273);
xnor U103 (N_103,In_2483,In_4240);
and U104 (N_104,In_702,In_1629);
xor U105 (N_105,In_1483,In_3824);
and U106 (N_106,In_1910,In_2675);
and U107 (N_107,In_2728,In_4296);
and U108 (N_108,In_1824,In_4116);
or U109 (N_109,In_2367,In_1283);
or U110 (N_110,In_1801,In_3526);
and U111 (N_111,In_2857,In_4640);
nand U112 (N_112,In_2741,In_1732);
nand U113 (N_113,In_2134,In_2628);
and U114 (N_114,In_3856,In_1060);
nand U115 (N_115,In_4784,In_3467);
nor U116 (N_116,In_4156,In_2200);
nor U117 (N_117,In_2719,In_3761);
and U118 (N_118,In_2022,In_2290);
and U119 (N_119,In_4927,In_4697);
xnor U120 (N_120,In_1764,In_3033);
nand U121 (N_121,In_1095,In_1034);
and U122 (N_122,In_871,In_4347);
nand U123 (N_123,In_1636,In_4242);
and U124 (N_124,In_2446,In_3426);
nand U125 (N_125,In_4190,In_2896);
nand U126 (N_126,In_4891,In_2971);
nand U127 (N_127,In_2026,In_1337);
nor U128 (N_128,In_1678,In_749);
or U129 (N_129,In_2123,In_1893);
nand U130 (N_130,In_2009,In_2615);
and U131 (N_131,In_4842,In_719);
and U132 (N_132,In_4663,In_3840);
nor U133 (N_133,In_97,In_2569);
or U134 (N_134,In_2393,In_1761);
and U135 (N_135,In_2427,In_2192);
or U136 (N_136,In_3774,In_1333);
nor U137 (N_137,In_148,In_2001);
xor U138 (N_138,In_101,In_88);
and U139 (N_139,In_2922,In_3608);
nand U140 (N_140,In_1840,In_2899);
nand U141 (N_141,In_2703,In_3080);
nor U142 (N_142,In_3423,In_734);
nand U143 (N_143,In_3993,In_1193);
and U144 (N_144,In_2450,In_3931);
and U145 (N_145,In_3884,In_1024);
or U146 (N_146,In_4998,In_1202);
or U147 (N_147,In_193,In_1396);
nand U148 (N_148,In_1806,In_4009);
nand U149 (N_149,In_4377,In_3129);
nand U150 (N_150,In_13,In_2856);
nor U151 (N_151,In_691,In_386);
or U152 (N_152,In_4491,In_3578);
and U153 (N_153,In_3030,In_3304);
nand U154 (N_154,In_2241,In_1523);
or U155 (N_155,In_293,In_4326);
nand U156 (N_156,In_878,In_642);
and U157 (N_157,In_129,In_4984);
xor U158 (N_158,In_677,In_1088);
or U159 (N_159,In_911,In_4658);
and U160 (N_160,In_3224,In_4399);
nand U161 (N_161,In_3653,In_3142);
or U162 (N_162,In_4029,In_684);
nand U163 (N_163,In_1344,In_2601);
xor U164 (N_164,In_2414,In_576);
nand U165 (N_165,In_2705,In_1891);
or U166 (N_166,In_2448,In_587);
or U167 (N_167,In_2765,In_3977);
nand U168 (N_168,In_3917,In_3590);
and U169 (N_169,In_4162,In_3266);
nand U170 (N_170,In_2991,In_3167);
and U171 (N_171,In_2858,In_1885);
and U172 (N_172,In_868,In_1574);
nand U173 (N_173,In_1979,In_571);
xnor U174 (N_174,In_1160,In_3854);
nor U175 (N_175,In_4204,In_2204);
and U176 (N_176,In_3716,In_1728);
or U177 (N_177,In_128,In_3721);
or U178 (N_178,In_3539,In_757);
nand U179 (N_179,In_1453,In_2909);
xnor U180 (N_180,In_2832,In_931);
nand U181 (N_181,In_4461,In_2043);
nor U182 (N_182,In_221,In_2638);
and U183 (N_183,In_1799,In_116);
nand U184 (N_184,In_4249,In_1443);
and U185 (N_185,In_2066,In_4354);
and U186 (N_186,In_3976,In_851);
nand U187 (N_187,In_2646,In_2291);
nand U188 (N_188,In_1002,In_3490);
nand U189 (N_189,In_4702,In_4186);
nand U190 (N_190,In_4690,In_4810);
nand U191 (N_191,In_1097,In_4489);
or U192 (N_192,In_1628,In_3113);
nand U193 (N_193,In_4504,In_1284);
and U194 (N_194,In_326,In_957);
and U195 (N_195,In_3400,In_4849);
nand U196 (N_196,In_2490,In_1830);
and U197 (N_197,In_4191,In_3918);
nor U198 (N_198,In_1825,In_775);
xnor U199 (N_199,In_2215,In_2092);
and U200 (N_200,In_4651,In_4867);
and U201 (N_201,In_2774,In_2178);
nand U202 (N_202,In_1672,In_3834);
or U203 (N_203,In_2788,In_2579);
nor U204 (N_204,In_455,In_3437);
and U205 (N_205,In_4339,In_1850);
and U206 (N_206,In_4526,In_4786);
and U207 (N_207,In_486,In_63);
or U208 (N_208,In_4766,In_1956);
nor U209 (N_209,In_461,In_1457);
nor U210 (N_210,In_2162,In_1140);
xor U211 (N_211,In_235,In_3503);
or U212 (N_212,In_4800,In_2864);
and U213 (N_213,In_1085,In_890);
or U214 (N_214,In_4360,In_2350);
or U215 (N_215,In_3074,In_2848);
nor U216 (N_216,In_410,In_49);
nor U217 (N_217,In_3604,In_1503);
and U218 (N_218,In_429,In_1127);
and U219 (N_219,In_3819,In_671);
and U220 (N_220,In_81,In_4751);
xor U221 (N_221,In_741,In_4017);
or U222 (N_222,In_4041,In_4058);
and U223 (N_223,In_378,In_805);
and U224 (N_224,In_2927,In_4902);
or U225 (N_225,In_3926,In_2380);
or U226 (N_226,In_359,In_4219);
xnor U227 (N_227,In_951,In_440);
nand U228 (N_228,In_2293,In_4532);
and U229 (N_229,In_1576,In_4674);
nand U230 (N_230,In_678,In_2208);
nand U231 (N_231,In_4306,In_2114);
or U232 (N_232,In_4024,In_3619);
or U233 (N_233,In_4746,In_3678);
nand U234 (N_234,In_1798,In_3201);
nor U235 (N_235,In_4159,In_1345);
and U236 (N_236,In_772,In_4404);
xnor U237 (N_237,In_4944,In_3393);
nand U238 (N_238,In_862,In_2258);
nand U239 (N_239,In_3570,In_3588);
and U240 (N_240,In_4852,In_3731);
and U241 (N_241,In_2784,In_4392);
or U242 (N_242,In_3660,In_474);
nor U243 (N_243,In_3331,In_2247);
and U244 (N_244,In_1470,In_2228);
and U245 (N_245,In_1747,In_1439);
nor U246 (N_246,In_1408,In_952);
and U247 (N_247,In_3461,In_2926);
or U248 (N_248,In_645,In_4601);
or U249 (N_249,In_4856,In_2400);
nand U250 (N_250,In_4862,In_942);
or U251 (N_251,In_4252,In_3336);
nand U252 (N_252,In_2918,In_2712);
nor U253 (N_253,In_436,In_2936);
nor U254 (N_254,In_1901,In_3361);
and U255 (N_255,In_120,In_1736);
nor U256 (N_256,In_2621,In_4598);
nand U257 (N_257,In_4291,In_3889);
and U258 (N_258,In_3115,In_2507);
nand U259 (N_259,In_818,In_1419);
nand U260 (N_260,In_4531,In_3628);
nand U261 (N_261,In_1955,In_2613);
or U262 (N_262,In_961,In_452);
or U263 (N_263,In_2429,In_3777);
or U264 (N_264,In_3428,In_4146);
and U265 (N_265,In_171,In_572);
nand U266 (N_266,In_2044,In_325);
nor U267 (N_267,In_1278,In_2140);
and U268 (N_268,In_4524,In_4947);
and U269 (N_269,In_3486,In_4631);
nor U270 (N_270,In_4272,In_964);
xnor U271 (N_271,In_4668,In_1310);
nand U272 (N_272,In_3814,In_3425);
and U273 (N_273,In_621,In_2090);
nand U274 (N_274,In_4028,In_1811);
or U275 (N_275,In_194,In_2316);
and U276 (N_276,In_1828,In_2827);
nor U277 (N_277,In_1683,In_72);
and U278 (N_278,In_4961,In_1990);
and U279 (N_279,In_177,In_2640);
nor U280 (N_280,In_244,In_309);
and U281 (N_281,In_2097,In_2893);
xnor U282 (N_282,In_4896,In_1101);
nor U283 (N_283,In_966,In_4565);
nand U284 (N_284,In_2660,In_1662);
nand U285 (N_285,In_4331,In_4883);
xnor U286 (N_286,In_1165,In_4550);
nand U287 (N_287,In_2199,In_4248);
or U288 (N_288,In_4036,In_1787);
and U289 (N_289,In_3499,In_1154);
xnor U290 (N_290,In_4216,In_585);
xor U291 (N_291,In_4164,In_3673);
xor U292 (N_292,In_470,In_3226);
nand U293 (N_293,In_2379,In_3921);
nor U294 (N_294,In_4126,In_2262);
or U295 (N_295,In_1188,In_1875);
and U296 (N_296,In_4600,In_4228);
and U297 (N_297,In_2369,In_2592);
or U298 (N_298,In_4429,In_2366);
and U299 (N_299,In_4070,In_1758);
or U300 (N_300,In_281,In_2722);
and U301 (N_301,In_524,In_2757);
and U302 (N_302,In_275,In_2421);
nand U303 (N_303,In_2702,In_2187);
nand U304 (N_304,In_3208,In_1091);
or U305 (N_305,In_503,In_2878);
xnor U306 (N_306,In_2431,In_2833);
nor U307 (N_307,In_145,In_2023);
and U308 (N_308,In_2913,In_449);
xnor U309 (N_309,In_1917,In_4954);
and U310 (N_310,In_1075,In_467);
nand U311 (N_311,In_987,In_2768);
nand U312 (N_312,In_3649,In_1981);
nor U313 (N_313,In_1192,In_3502);
or U314 (N_314,In_3207,In_4081);
and U315 (N_315,In_4868,In_3191);
or U316 (N_316,In_4854,In_1442);
or U317 (N_317,In_4076,In_2604);
nand U318 (N_318,In_2377,In_4473);
and U319 (N_319,In_613,In_4239);
nor U320 (N_320,In_1933,In_2508);
or U321 (N_321,In_3411,In_337);
nand U322 (N_322,In_2575,In_2157);
or U323 (N_323,In_2321,In_2378);
xor U324 (N_324,In_1660,In_3067);
and U325 (N_325,In_1888,In_948);
nand U326 (N_326,In_2693,In_2072);
nor U327 (N_327,In_542,In_2706);
nor U328 (N_328,In_655,In_2002);
nor U329 (N_329,In_4394,In_3969);
and U330 (N_330,In_56,In_3565);
nor U331 (N_331,In_492,In_4418);
and U332 (N_332,In_80,In_652);
or U333 (N_333,In_156,In_3200);
and U334 (N_334,In_1520,In_1013);
or U335 (N_335,In_1019,In_651);
nand U336 (N_336,In_4705,In_3333);
nor U337 (N_337,In_2707,In_2006);
and U338 (N_338,In_140,In_453);
and U339 (N_339,In_1751,In_1550);
nor U340 (N_340,In_4417,In_2317);
nand U341 (N_341,In_3763,In_4055);
nand U342 (N_342,In_4778,In_2627);
xor U343 (N_343,In_3541,In_4498);
or U344 (N_344,In_3452,In_2133);
nor U345 (N_345,In_1258,In_1571);
nor U346 (N_346,In_4292,In_3029);
nand U347 (N_347,In_534,In_465);
and U348 (N_348,In_4793,In_1380);
or U349 (N_349,In_1776,In_2533);
nand U350 (N_350,In_870,In_1890);
or U351 (N_351,In_2335,In_1991);
xnor U352 (N_352,In_4643,In_3020);
and U353 (N_353,In_4129,In_811);
nor U354 (N_354,In_1052,In_2946);
nand U355 (N_355,In_1564,In_3729);
nor U356 (N_356,In_2201,In_3929);
and U357 (N_357,In_1871,In_2889);
nand U358 (N_358,In_4264,In_3005);
and U359 (N_359,In_4845,In_1521);
nand U360 (N_360,In_3286,In_706);
and U361 (N_361,In_497,In_1591);
nand U362 (N_362,In_342,In_3132);
and U363 (N_363,In_3387,In_3966);
or U364 (N_364,In_3650,In_4514);
nand U365 (N_365,In_3624,In_2433);
and U366 (N_366,In_4507,In_1692);
nor U367 (N_367,In_861,In_418);
or U368 (N_368,In_2547,In_4142);
nand U369 (N_369,In_1001,In_1405);
xor U370 (N_370,In_3004,In_3505);
nor U371 (N_371,In_3700,In_4560);
nor U372 (N_372,In_99,In_1906);
or U373 (N_373,In_880,In_1210);
nand U374 (N_374,In_1814,In_3740);
and U375 (N_375,In_1818,In_688);
nand U376 (N_376,In_3670,In_2663);
and U377 (N_377,In_4315,In_2673);
and U378 (N_378,In_2027,In_2637);
and U379 (N_379,In_1849,In_2181);
nor U380 (N_380,In_2502,In_3143);
or U381 (N_381,In_2819,In_1530);
or U382 (N_382,In_1432,In_127);
nor U383 (N_383,In_971,In_2126);
nand U384 (N_384,In_1832,In_1653);
and U385 (N_385,In_604,In_3292);
and U386 (N_386,In_380,In_799);
nand U387 (N_387,In_4014,In_50);
nand U388 (N_388,In_2917,In_4411);
or U389 (N_389,In_4474,In_2504);
or U390 (N_390,In_273,In_3790);
nand U391 (N_391,In_103,In_3742);
nand U392 (N_392,In_1426,In_1673);
nand U393 (N_393,In_1739,In_3328);
and U394 (N_394,In_1725,In_4462);
or U395 (N_395,In_2924,In_4385);
or U396 (N_396,In_714,In_986);
nand U397 (N_397,In_3031,In_599);
nand U398 (N_398,In_464,In_4529);
xnor U399 (N_399,In_4195,In_4148);
nor U400 (N_400,In_119,In_2845);
or U401 (N_401,In_1434,In_504);
xnor U402 (N_402,In_3306,In_4945);
xor U403 (N_403,In_2347,In_1561);
and U404 (N_404,In_689,In_494);
nor U405 (N_405,In_2559,In_958);
and U406 (N_406,In_4988,In_3659);
and U407 (N_407,In_3924,In_4470);
or U408 (N_408,In_1070,In_2381);
xor U409 (N_409,In_2464,In_2843);
or U410 (N_410,In_1833,In_1755);
xor U411 (N_411,In_3934,In_4899);
nor U412 (N_412,In_568,In_939);
xor U413 (N_413,In_3219,In_3364);
and U414 (N_414,In_4995,In_3375);
nand U415 (N_415,In_573,In_1584);
nand U416 (N_416,In_3961,In_2781);
and U417 (N_417,In_703,In_3900);
nand U418 (N_418,In_1122,In_1375);
or U419 (N_419,In_1224,In_4646);
nand U420 (N_420,In_2417,In_3564);
nand U421 (N_421,In_2850,In_2211);
or U422 (N_422,In_4641,In_525);
xnor U423 (N_423,In_802,In_1228);
or U424 (N_424,In_916,In_2348);
nand U425 (N_425,In_1986,In_2315);
or U426 (N_426,In_4109,In_1942);
nand U427 (N_427,In_2154,In_3985);
and U428 (N_428,In_1079,In_4152);
nand U429 (N_429,In_1113,In_4613);
and U430 (N_430,In_924,In_618);
nand U431 (N_431,In_4727,In_2609);
nor U432 (N_432,In_3277,In_2407);
or U433 (N_433,In_3691,In_3014);
or U434 (N_434,In_3250,In_1648);
or U435 (N_435,In_2153,In_2237);
xnor U436 (N_436,In_3023,In_118);
xnor U437 (N_437,In_431,In_3383);
nand U438 (N_438,In_1050,In_3003);
nor U439 (N_439,In_213,In_1974);
nor U440 (N_440,In_182,In_4480);
or U441 (N_441,In_4194,In_3340);
or U442 (N_442,In_3881,In_388);
nor U443 (N_443,In_4969,In_4367);
nand U444 (N_444,In_1609,In_4089);
or U445 (N_445,In_3607,In_3714);
xor U446 (N_446,In_1350,In_2883);
and U447 (N_447,In_1305,In_3026);
or U448 (N_448,In_1529,In_4300);
nor U449 (N_449,In_690,In_4336);
and U450 (N_450,In_4022,In_3749);
nor U451 (N_451,In_1753,In_4909);
nand U452 (N_452,In_1216,In_3275);
nand U453 (N_453,In_4684,In_2645);
nor U454 (N_454,In_653,In_210);
nor U455 (N_455,In_3591,In_763);
nor U456 (N_456,In_4494,In_661);
nor U457 (N_457,In_4311,In_2249);
nand U458 (N_458,In_1543,In_3928);
nand U459 (N_459,In_4678,In_162);
nor U460 (N_460,In_4030,In_114);
nor U461 (N_461,In_2736,In_1448);
nor U462 (N_462,In_2182,In_1579);
nand U463 (N_463,In_2280,In_3089);
nor U464 (N_464,In_256,In_3764);
or U465 (N_465,In_4280,In_2438);
xnor U466 (N_466,In_2270,In_842);
and U467 (N_467,In_371,In_1491);
nand U468 (N_468,In_1365,In_1712);
nor U469 (N_469,In_3964,In_345);
and U470 (N_470,In_2288,In_4762);
nand U471 (N_471,In_4042,In_1959);
or U472 (N_472,In_3479,In_771);
and U473 (N_473,In_2163,In_4267);
xor U474 (N_474,In_566,In_747);
xnor U475 (N_475,In_4167,In_854);
xnor U476 (N_476,In_3458,In_1383);
nor U477 (N_477,In_2062,In_1655);
xor U478 (N_478,In_2058,In_1598);
or U479 (N_479,In_1297,In_3248);
nor U480 (N_480,In_3686,In_662);
or U481 (N_481,In_3688,In_2482);
nand U482 (N_482,In_2183,In_3672);
nand U483 (N_483,In_85,In_1487);
xnor U484 (N_484,In_45,In_2296);
and U485 (N_485,In_3193,In_175);
nand U486 (N_486,In_3178,In_2939);
nor U487 (N_487,In_1635,In_211);
and U488 (N_488,In_2582,In_4659);
or U489 (N_489,In_1341,In_4266);
and U490 (N_490,In_4145,In_4359);
and U491 (N_491,In_2961,In_2825);
and U492 (N_492,In_4825,In_1450);
nand U493 (N_493,In_1077,In_3391);
nor U494 (N_494,In_2359,In_1738);
nor U495 (N_495,In_1519,In_1185);
or U496 (N_496,In_117,In_4415);
nor U497 (N_497,In_237,In_2131);
nor U498 (N_498,In_4033,In_3885);
or U499 (N_499,In_2033,In_3100);
nor U500 (N_500,In_3338,In_1119);
or U501 (N_501,In_3600,In_3614);
nand U502 (N_502,In_4921,In_602);
nand U503 (N_503,In_491,In_1769);
nand U504 (N_504,In_4701,In_4213);
or U505 (N_505,In_4982,In_489);
nor U506 (N_506,In_1494,In_1051);
and U507 (N_507,In_1693,In_1676);
nor U508 (N_508,In_598,In_3035);
nand U509 (N_509,In_4941,In_2750);
or U510 (N_510,In_4530,In_2515);
nand U511 (N_511,In_2747,In_4134);
and U512 (N_512,In_929,In_2232);
and U513 (N_513,In_1746,In_3507);
xnor U514 (N_514,In_1126,In_3194);
nand U515 (N_515,In_424,In_1257);
nor U516 (N_516,In_2954,In_4181);
nor U517 (N_517,In_3903,In_1479);
and U518 (N_518,In_3750,In_549);
or U519 (N_519,In_4675,In_1622);
nand U520 (N_520,In_3645,In_591);
and U521 (N_521,In_4692,In_1829);
and U522 (N_522,In_1038,In_3335);
or U523 (N_523,In_4136,In_4325);
and U524 (N_524,In_1689,In_1357);
nand U525 (N_525,In_4860,In_4976);
nand U526 (N_526,In_4452,In_1545);
or U527 (N_527,In_959,In_4955);
nor U528 (N_528,In_4940,In_578);
or U529 (N_529,In_206,In_419);
nor U530 (N_530,In_1709,In_551);
nand U531 (N_531,In_2477,In_265);
or U532 (N_532,In_283,In_740);
nor U533 (N_533,In_780,In_2735);
or U534 (N_534,In_3360,In_2432);
xnor U535 (N_535,In_1295,In_896);
nor U536 (N_536,In_1407,In_1141);
nor U537 (N_537,In_3920,In_3620);
and U538 (N_538,In_4233,In_935);
nor U539 (N_539,In_833,In_433);
nor U540 (N_540,In_3572,In_4062);
xor U541 (N_541,In_1794,In_1110);
nand U542 (N_542,In_1199,In_2149);
or U543 (N_543,In_781,In_3747);
nand U544 (N_544,In_1469,In_3675);
or U545 (N_545,In_2088,In_2803);
nor U546 (N_546,In_296,In_2456);
and U547 (N_547,In_4905,In_4063);
or U548 (N_548,In_809,In_3520);
and U549 (N_549,In_2882,In_2019);
and U550 (N_550,In_960,In_0);
nand U551 (N_551,In_2872,In_1665);
and U552 (N_552,In_3972,In_1842);
xor U553 (N_553,In_993,In_441);
nor U554 (N_554,In_1909,In_630);
and U555 (N_555,In_3799,In_4269);
and U556 (N_556,In_1652,In_3707);
and U557 (N_557,In_1018,In_1117);
and U558 (N_558,In_2248,In_1307);
nand U559 (N_559,In_390,In_1715);
or U560 (N_560,In_1688,In_1221);
xor U561 (N_561,In_2548,In_4464);
and U562 (N_562,In_4911,In_2494);
nor U563 (N_563,In_4287,In_4051);
nor U564 (N_564,In_2224,In_3077);
xor U565 (N_565,In_1104,In_3470);
nand U566 (N_566,In_4543,In_4379);
or U567 (N_567,In_2462,In_4936);
nand U568 (N_568,In_2074,In_1169);
nor U569 (N_569,In_4485,In_216);
or U570 (N_570,In_4123,In_100);
nor U571 (N_571,In_2257,In_4241);
xnor U572 (N_572,In_203,In_4923);
nor U573 (N_573,In_1999,In_376);
nand U574 (N_574,In_1615,In_1962);
or U575 (N_575,In_4405,In_825);
and U576 (N_576,In_1784,In_1667);
nand U577 (N_577,In_4038,In_3753);
nor U578 (N_578,In_2301,In_3982);
and U579 (N_579,In_3181,In_8);
nand U580 (N_580,In_2976,In_856);
nor U581 (N_581,In_938,In_3404);
nor U582 (N_582,In_1691,In_4539);
or U583 (N_583,In_3161,In_4811);
and U584 (N_584,In_1473,In_2902);
nand U585 (N_585,In_3967,In_2685);
nor U586 (N_586,In_3587,In_974);
nor U587 (N_587,In_2852,In_2465);
nor U588 (N_588,In_3133,In_3258);
xor U589 (N_589,In_434,In_443);
or U590 (N_590,In_2875,In_4586);
xor U591 (N_591,In_1924,In_1848);
and U592 (N_592,In_1029,In_1044);
nor U593 (N_593,In_3679,In_356);
xor U594 (N_594,In_3725,In_4093);
or U595 (N_595,In_130,In_4174);
xor U596 (N_596,In_4730,In_2440);
nand U597 (N_597,In_3041,In_476);
nand U598 (N_598,In_2128,In_3756);
and U599 (N_599,In_1208,In_1496);
nand U600 (N_600,In_750,In_1235);
nand U601 (N_601,In_2260,In_736);
xnor U602 (N_602,In_3952,In_3318);
nor U603 (N_603,In_4343,In_4138);
and U604 (N_604,In_788,In_2691);
nand U605 (N_605,In_1250,In_4797);
nor U606 (N_606,In_897,In_4623);
nor U607 (N_607,In_3957,In_3012);
xnor U608 (N_608,In_1657,In_1300);
nand U609 (N_609,In_1834,In_2439);
or U610 (N_610,In_422,In_155);
nand U611 (N_611,In_1428,In_3685);
nand U612 (N_612,In_2354,In_4808);
and U613 (N_613,In_4423,In_3480);
nor U614 (N_614,In_3136,In_682);
or U615 (N_615,In_2255,In_552);
nand U616 (N_616,In_414,In_3481);
nor U617 (N_617,In_1524,In_647);
nand U618 (N_618,In_3366,In_3737);
nand U619 (N_619,In_635,In_1264);
nand U620 (N_620,In_328,In_1775);
or U621 (N_621,In_2901,In_4803);
and U622 (N_622,In_985,In_2061);
nor U623 (N_623,In_3424,In_2545);
xnor U624 (N_624,In_3945,In_2363);
nand U625 (N_625,In_2244,In_2336);
or U626 (N_626,In_1844,In_2130);
nor U627 (N_627,In_3925,In_1843);
nand U628 (N_628,In_1135,In_1941);
and U629 (N_629,In_3949,In_2950);
or U630 (N_630,In_403,In_4438);
and U631 (N_631,In_2413,In_4588);
or U632 (N_632,In_908,In_4889);
and U633 (N_633,In_2233,In_3394);
and U634 (N_634,In_4368,In_3542);
xor U635 (N_635,In_3710,In_2171);
or U636 (N_636,In_1347,In_820);
and U637 (N_637,In_377,In_2480);
or U638 (N_638,In_1953,In_1939);
nand U639 (N_639,In_2098,In_17);
and U640 (N_640,In_3463,In_1403);
and U641 (N_641,In_937,In_2415);
nand U642 (N_642,In_1705,In_3664);
xnor U643 (N_643,In_3744,In_3739);
and U644 (N_644,In_4618,In_4603);
or U645 (N_645,In_4482,In_4558);
nor U646 (N_646,In_2332,In_3775);
and U647 (N_647,In_2454,In_3283);
or U648 (N_648,In_124,In_1781);
nand U649 (N_649,In_4048,In_3537);
nand U650 (N_650,In_3898,In_4731);
or U651 (N_651,In_398,In_3858);
or U652 (N_652,In_4084,In_2442);
and U653 (N_653,In_2672,In_1446);
nor U654 (N_654,In_3755,In_2216);
nor U655 (N_655,In_3210,In_3641);
or U656 (N_656,In_22,In_4501);
nor U657 (N_657,In_3684,In_2631);
nand U658 (N_658,In_1376,In_396);
or U659 (N_659,In_1292,In_2283);
nor U660 (N_660,In_4773,In_3013);
nor U661 (N_661,In_1804,In_2085);
and U662 (N_662,In_1229,In_2488);
and U663 (N_663,In_1509,In_1687);
nor U664 (N_664,In_698,In_3654);
nand U665 (N_665,In_3021,In_4948);
nor U666 (N_666,In_3491,In_991);
and U667 (N_667,In_841,In_2517);
nand U668 (N_668,In_2109,In_3255);
and U669 (N_669,In_3228,In_3767);
nor U670 (N_670,In_294,In_456);
or U671 (N_671,In_2070,In_2345);
nand U672 (N_672,In_4149,In_3027);
nor U673 (N_673,In_417,In_579);
nor U674 (N_674,In_3104,In_1920);
or U675 (N_675,In_1076,In_934);
nand U676 (N_676,In_2639,In_2177);
nor U677 (N_677,In_634,In_3909);
or U678 (N_678,In_2175,In_387);
nor U679 (N_679,In_1325,In_2770);
and U680 (N_680,In_2082,In_412);
or U681 (N_681,In_291,In_3378);
or U682 (N_682,In_2668,In_4422);
or U683 (N_683,In_1301,In_2392);
and U684 (N_684,In_784,In_1697);
nor U685 (N_685,In_1717,In_4054);
or U686 (N_686,In_3709,In_263);
nand U687 (N_687,In_2563,In_953);
or U688 (N_688,In_3802,In_4865);
or U689 (N_689,In_1816,In_4435);
or U690 (N_690,In_4312,In_54);
or U691 (N_691,In_3000,In_537);
nor U692 (N_692,In_4742,In_318);
and U693 (N_693,In_3202,In_1286);
and U694 (N_694,In_3912,In_4439);
and U695 (N_695,In_478,In_1222);
or U696 (N_696,In_391,In_1867);
and U697 (N_697,In_1413,In_4283);
and U698 (N_698,In_4665,In_3914);
nor U699 (N_699,In_687,In_1055);
or U700 (N_700,In_303,In_3862);
or U701 (N_701,In_1402,In_518);
and U702 (N_702,In_3818,In_3549);
nand U703 (N_703,In_4619,In_329);
nand U704 (N_704,In_2641,In_3144);
and U705 (N_705,In_3443,In_1048);
and U706 (N_706,In_1580,In_2797);
and U707 (N_707,In_1386,In_3519);
nor U708 (N_708,In_2791,In_4943);
or U709 (N_709,In_241,In_4341);
nand U710 (N_710,In_2721,In_2769);
nand U711 (N_711,In_4789,In_1105);
and U712 (N_712,In_2554,In_4401);
or U713 (N_713,In_186,In_1103);
xnor U714 (N_714,In_4295,In_1668);
xor U715 (N_715,In_3849,In_43);
nand U716 (N_716,In_1602,In_4913);
nand U717 (N_717,In_2391,In_2463);
and U718 (N_718,In_2578,In_4039);
nand U719 (N_719,In_147,In_1633);
nand U720 (N_720,In_3867,In_1394);
and U721 (N_721,In_2013,In_2767);
or U722 (N_722,In_1964,In_1935);
nand U723 (N_723,In_3319,In_554);
or U724 (N_724,In_3209,In_198);
xnor U725 (N_725,In_4303,In_4425);
nand U726 (N_726,In_2051,In_4875);
and U727 (N_727,In_4656,In_3643);
nor U728 (N_728,In_2643,In_3613);
nand U729 (N_729,In_2710,In_2173);
nor U730 (N_730,In_4624,In_3847);
xnor U731 (N_731,In_1293,In_1853);
nor U732 (N_732,In_1931,In_4077);
and U733 (N_733,In_4434,In_2276);
nand U734 (N_734,In_295,In_70);
and U735 (N_735,In_2524,In_1472);
and U736 (N_736,In_79,In_4393);
or U737 (N_737,In_254,In_2295);
nand U738 (N_738,In_1791,In_2862);
nor U739 (N_739,In_2561,In_3979);
nor U740 (N_740,In_3152,In_4968);
nor U741 (N_741,In_2353,In_405);
nor U742 (N_742,In_278,In_92);
or U743 (N_743,In_3369,In_4476);
or U744 (N_744,In_1121,In_2597);
nor U745 (N_745,In_726,In_1894);
nand U746 (N_746,In_783,In_4500);
nor U747 (N_747,In_1695,In_1138);
or U748 (N_748,In_1249,In_266);
or U749 (N_749,In_4873,In_3098);
and U750 (N_750,In_1947,In_4928);
xnor U751 (N_751,In_3629,In_3546);
nand U752 (N_752,In_2514,In_746);
and U753 (N_753,In_1454,In_4430);
nor U754 (N_754,In_1460,In_1946);
nand U755 (N_755,In_3689,In_4064);
nand U756 (N_756,In_2505,In_755);
and U757 (N_757,In_2473,In_710);
or U758 (N_758,In_1189,In_2386);
or U759 (N_759,In_679,In_2018);
nor U760 (N_760,In_4271,In_1852);
xnor U761 (N_761,In_4983,In_3723);
xnor U762 (N_762,In_4007,In_770);
or U763 (N_763,In_2423,In_2174);
or U764 (N_764,In_3356,In_1730);
and U765 (N_765,In_4741,In_288);
nor U766 (N_766,In_4872,In_4044);
nand U767 (N_767,In_236,In_3138);
or U768 (N_768,In_2340,In_4801);
nor U769 (N_769,In_4043,In_108);
or U770 (N_770,In_1062,In_752);
nand U771 (N_771,In_626,In_4389);
and U772 (N_772,In_1594,In_1251);
and U773 (N_773,In_1003,In_1534);
and U774 (N_774,In_1136,In_859);
nor U775 (N_775,In_907,In_59);
nor U776 (N_776,In_2724,In_4671);
or U777 (N_777,In_657,In_4516);
nor U778 (N_778,In_3765,In_2614);
xnor U779 (N_779,In_1954,In_1393);
nor U780 (N_780,In_1355,In_4175);
xor U781 (N_781,In_4915,In_1817);
or U782 (N_782,In_1377,In_3079);
xnor U783 (N_783,In_2238,In_4580);
and U784 (N_784,In_3060,In_4169);
nor U785 (N_785,In_4901,In_4154);
nor U786 (N_786,In_3518,In_4599);
or U787 (N_787,In_2418,In_1565);
and U788 (N_788,In_180,In_4796);
and U789 (N_789,In_3122,In_2428);
or U790 (N_790,In_212,In_3488);
and U791 (N_791,In_3299,In_4686);
nor U792 (N_792,In_2306,In_2759);
nor U793 (N_793,In_2365,In_2282);
nor U794 (N_794,In_2397,In_4749);
or U795 (N_795,In_1694,In_3016);
nor U796 (N_796,In_1275,In_3241);
and U797 (N_797,In_33,In_2451);
and U798 (N_798,In_2607,In_4025);
nor U799 (N_799,In_3243,In_2060);
nor U800 (N_800,In_1256,In_2873);
xor U801 (N_801,In_567,In_3597);
and U802 (N_802,In_659,In_1723);
xor U803 (N_803,In_1299,In_1957);
and U804 (N_804,In_348,In_1444);
nor U805 (N_805,In_586,In_3343);
nand U806 (N_806,In_768,In_1856);
nor U807 (N_807,In_4918,In_4739);
and U808 (N_808,In_3037,In_885);
nand U809 (N_809,In_1908,In_324);
or U810 (N_810,In_1976,In_4534);
nor U811 (N_811,In_2087,In_4121);
nand U812 (N_812,In_2185,In_2221);
nand U813 (N_813,In_2119,In_4101);
and U814 (N_814,In_3154,In_2814);
or U815 (N_815,In_2606,In_4681);
xor U816 (N_816,In_2501,In_1093);
and U817 (N_817,In_1826,In_4733);
or U818 (N_818,In_2566,In_2963);
nor U819 (N_819,In_1731,In_276);
or U820 (N_820,In_4959,In_1729);
or U821 (N_821,In_1037,In_1248);
nor U822 (N_822,In_2300,In_2209);
nand U823 (N_823,In_3786,In_2069);
and U824 (N_824,In_3989,In_215);
nor U825 (N_825,In_1025,In_4130);
nand U826 (N_826,In_3377,In_1409);
nand U827 (N_827,In_1064,In_4199);
nor U828 (N_828,In_2570,In_4892);
nand U829 (N_829,In_1164,In_1782);
nor U830 (N_830,In_1465,In_93);
and U831 (N_831,In_4380,In_2867);
and U832 (N_832,In_4003,In_4799);
xnor U833 (N_833,In_3821,In_2577);
and U834 (N_834,In_4819,In_3915);
nor U835 (N_835,In_2682,In_900);
and U836 (N_836,In_1134,In_3873);
nand U837 (N_837,In_77,In_2021);
or U838 (N_838,In_4369,In_1560);
xor U839 (N_839,In_4528,In_1645);
or U840 (N_840,In_3785,In_1277);
or U841 (N_841,In_4031,In_664);
nor U842 (N_842,In_3851,In_4782);
and U843 (N_843,In_4790,In_3017);
or U844 (N_844,In_2975,In_4951);
and U845 (N_845,In_2373,In_4655);
and U846 (N_846,In_32,In_3285);
and U847 (N_847,In_1066,In_4090);
nand U848 (N_848,In_1203,In_2225);
or U849 (N_849,In_4361,In_1429);
nand U850 (N_850,In_3198,In_1674);
and U851 (N_851,In_1348,In_4250);
or U852 (N_852,In_1006,In_1887);
nor U853 (N_853,In_2993,In_2434);
or U854 (N_854,In_113,In_3184);
nand U855 (N_855,In_692,In_1351);
nand U856 (N_856,In_1879,In_3439);
and U857 (N_857,In_3442,In_4703);
or U858 (N_858,In_4625,In_4666);
xnor U859 (N_859,In_4391,In_4606);
xor U860 (N_860,In_3140,In_3724);
nor U861 (N_861,In_2602,In_1506);
nor U862 (N_862,In_3746,In_4034);
xor U863 (N_863,In_2610,In_2826);
nand U864 (N_864,In_2476,In_1613);
nor U865 (N_865,In_3084,In_1510);
nor U866 (N_866,In_469,In_4748);
nor U867 (N_867,In_1255,In_1124);
or U868 (N_868,In_3621,In_4979);
xor U869 (N_869,In_3085,In_970);
and U870 (N_870,In_4553,In_992);
xnor U871 (N_871,In_2560,In_927);
nand U872 (N_872,In_4728,In_713);
nand U873 (N_873,In_4187,In_4270);
nand U874 (N_874,In_1312,In_2143);
nand U875 (N_875,In_849,In_1027);
nor U876 (N_876,In_3992,In_4382);
nor U877 (N_877,In_1466,In_3010);
nand U878 (N_878,In_3081,In_2384);
nor U879 (N_879,In_4736,In_1324);
or U880 (N_880,In_3268,In_695);
or U881 (N_881,In_3203,In_2731);
and U882 (N_882,In_505,In_1030);
xnor U883 (N_883,In_3459,In_4974);
nand U884 (N_884,In_2105,In_3878);
and U885 (N_885,In_4820,In_4907);
nor U886 (N_886,In_2756,In_3817);
or U887 (N_887,In_976,In_361);
and U888 (N_888,In_2522,In_2531);
nor U889 (N_889,In_4903,In_2125);
or U890 (N_890,In_4719,In_3456);
and U891 (N_891,In_3875,In_3626);
and U892 (N_892,In_1938,In_3585);
and U893 (N_893,In_1627,In_921);
and U894 (N_894,In_1274,In_3477);
or U895 (N_895,In_2818,In_839);
or U896 (N_896,In_1374,In_3676);
or U897 (N_897,In_3501,In_1992);
xnor U898 (N_898,In_720,In_2969);
and U899 (N_899,In_3496,In_2210);
nor U900 (N_900,In_3326,In_468);
or U901 (N_901,In_2478,In_1225);
and U902 (N_902,In_2132,In_3853);
and U903 (N_903,In_623,In_681);
and U904 (N_904,In_4920,In_3701);
nand U905 (N_905,In_824,In_1512);
or U906 (N_906,In_1595,In_3307);
and U907 (N_907,In_2370,In_3722);
xor U908 (N_908,In_3231,In_3406);
xor U909 (N_909,In_776,In_3554);
nor U910 (N_910,In_646,In_149);
nor U911 (N_911,In_286,In_2536);
nand U912 (N_912,In_1183,In_3032);
or U913 (N_913,In_4721,In_1273);
and U914 (N_914,In_3932,In_999);
xnor U915 (N_915,In_1518,In_233);
and U916 (N_916,In_2905,In_4085);
nor U917 (N_917,In_4541,In_3139);
nor U918 (N_918,In_831,In_2269);
nor U919 (N_919,In_3720,In_4804);
xor U920 (N_920,In_2538,In_1500);
and U921 (N_921,In_2394,In_4362);
xor U922 (N_922,In_2666,In_4224);
or U923 (N_923,In_2371,In_3532);
xnor U924 (N_924,In_1838,In_4350);
nand U925 (N_925,In_4155,In_4567);
nand U926 (N_926,In_2959,In_2222);
nand U927 (N_927,In_3327,In_3803);
or U928 (N_928,In_815,In_4724);
nor U929 (N_929,In_1656,In_2259);
nor U930 (N_930,In_4390,In_1726);
xor U931 (N_931,In_1661,In_51);
or U932 (N_932,In_3410,In_2802);
xor U933 (N_933,In_4760,In_3172);
and U934 (N_934,In_3196,In_4052);
or U935 (N_935,In_3046,In_3344);
or U936 (N_936,In_3274,In_3256);
and U937 (N_937,In_4925,In_1669);
nand U938 (N_938,In_4397,In_1320);
and U939 (N_939,In_1802,In_4433);
nor U940 (N_940,In_998,In_1142);
nor U941 (N_941,In_1290,In_226);
xor U942 (N_942,In_3476,In_4492);
and U943 (N_943,In_1406,In_1765);
nand U944 (N_944,In_2086,In_1144);
or U945 (N_945,In_1624,In_1998);
and U946 (N_946,In_2093,In_2828);
nor U947 (N_947,In_163,In_1698);
nor U948 (N_948,In_2471,In_302);
and U949 (N_949,In_4119,In_1184);
or U950 (N_950,In_1043,In_4200);
nand U951 (N_951,In_269,In_4235);
and U952 (N_952,In_3868,In_4997);
or U953 (N_953,In_66,In_4060);
and U954 (N_954,In_69,In_2923);
or U955 (N_955,In_1658,In_341);
and U956 (N_956,In_4210,In_4814);
nand U957 (N_957,In_2933,In_2337);
nand U958 (N_958,In_2725,In_138);
nand U959 (N_959,In_1481,In_650);
nand U960 (N_960,In_2870,In_1317);
and U961 (N_961,In_4509,In_2539);
and U962 (N_962,In_2910,In_4585);
nand U963 (N_963,In_1596,In_3759);
xnor U964 (N_964,In_1318,In_4253);
nor U965 (N_965,In_4771,In_1585);
nor U966 (N_966,In_460,In_962);
nand U967 (N_967,In_590,In_4967);
xnor U968 (N_968,In_485,In_4537);
and U969 (N_969,In_712,In_4607);
or U970 (N_970,In_176,In_980);
nor U971 (N_971,In_2580,In_4346);
nor U972 (N_972,In_3697,In_2985);
or U973 (N_973,In_1438,In_2179);
nand U974 (N_974,In_4100,In_1572);
or U975 (N_975,In_2659,In_2498);
and U976 (N_976,In_517,In_133);
and U977 (N_977,In_4223,In_1356);
nor U978 (N_978,In_3671,In_4319);
and U979 (N_979,In_877,In_4768);
and U980 (N_980,In_2943,In_1021);
xnor U981 (N_981,In_1232,In_4163);
nand U982 (N_982,In_1762,In_600);
and U983 (N_983,In_4356,In_3848);
nand U984 (N_984,In_3741,In_196);
nor U985 (N_985,In_4682,In_1773);
nand U986 (N_986,In_308,In_4559);
nor U987 (N_987,In_202,In_4720);
nor U988 (N_988,In_615,In_3008);
nand U989 (N_989,In_4193,In_3105);
nor U990 (N_990,In_514,In_3986);
and U991 (N_991,In_3998,In_4914);
or U992 (N_992,In_28,In_62);
xnor U993 (N_993,In_4676,In_2100);
nor U994 (N_994,In_385,In_1554);
and U995 (N_995,In_3263,In_4538);
and U996 (N_996,In_4139,In_2912);
nor U997 (N_997,In_144,In_2796);
nor U998 (N_998,In_501,In_696);
or U999 (N_999,In_3417,In_339);
nor U1000 (N_1000,In_2738,In_4432);
or U1001 (N_1001,In_4798,In_2894);
and U1002 (N_1002,In_3300,In_4113);
nand U1003 (N_1003,In_2281,In_4178);
nand U1004 (N_1004,In_2811,In_1195);
and U1005 (N_1005,In_3511,In_3048);
and U1006 (N_1006,In_4989,In_3114);
nor U1007 (N_1007,In_426,In_1583);
nor U1008 (N_1008,In_9,In_4850);
nand U1009 (N_1009,In_3305,In_884);
nand U1010 (N_1010,In_4481,In_3757);
xnor U1011 (N_1011,In_372,In_1768);
xor U1012 (N_1012,In_4463,In_1032);
or U1013 (N_1013,In_4688,In_3386);
nand U1014 (N_1014,In_2921,In_1215);
nand U1015 (N_1015,In_3309,In_64);
xnor U1016 (N_1016,In_1148,In_2103);
and U1017 (N_1017,In_2644,In_4099);
or U1018 (N_1018,In_4758,In_1993);
nand U1019 (N_1019,In_2104,In_2325);
or U1020 (N_1020,In_3950,In_3713);
nand U1021 (N_1021,In_3665,In_477);
xnor U1022 (N_1022,In_4114,In_2815);
xnor U1023 (N_1023,In_2677,In_3638);
nand U1024 (N_1024,In_4348,In_3699);
nand U1025 (N_1025,In_2059,In_4628);
nor U1026 (N_1026,In_2493,In_289);
and U1027 (N_1027,In_4232,In_4592);
xnor U1028 (N_1028,In_1514,In_4289);
nor U1029 (N_1029,In_2168,In_90);
nand U1030 (N_1030,In_2147,In_4297);
or U1031 (N_1031,In_2470,In_1868);
xor U1032 (N_1032,In_3843,In_4885);
nand U1033 (N_1033,In_1567,In_4277);
nand U1034 (N_1034,In_979,In_1701);
nor U1035 (N_1035,In_2435,In_3066);
nand U1036 (N_1036,In_223,In_1677);
and U1037 (N_1037,In_1877,In_2401);
and U1038 (N_1038,In_2242,In_360);
nor U1039 (N_1039,In_777,In_2156);
nor U1040 (N_1040,In_3974,In_1485);
or U1041 (N_1041,In_2937,In_1896);
and U1042 (N_1042,In_1575,In_2964);
or U1043 (N_1043,In_4274,In_1358);
or U1044 (N_1044,In_1482,In_565);
xor U1045 (N_1045,In_1915,In_2629);
or U1046 (N_1046,In_978,In_1090);
nor U1047 (N_1047,In_4910,In_4775);
and U1048 (N_1048,In_4958,In_1995);
nor U1049 (N_1049,In_4575,In_898);
nor U1050 (N_1050,In_2491,In_3719);
nor U1051 (N_1051,In_1425,In_3942);
or U1052 (N_1052,In_4521,In_1153);
or U1053 (N_1053,In_1049,In_207);
nand U1054 (N_1054,In_619,In_2808);
nand U1055 (N_1055,In_4827,In_3529);
and U1056 (N_1056,In_4238,In_1322);
xor U1057 (N_1057,In_1499,In_4716);
and U1058 (N_1058,In_3891,In_844);
and U1059 (N_1059,In_5,In_4888);
nor U1060 (N_1060,In_84,In_57);
xnor U1061 (N_1061,In_1551,In_3237);
nor U1062 (N_1062,In_3427,In_4561);
and U1063 (N_1063,In_3380,In_4897);
nor U1064 (N_1064,In_3093,In_4313);
nand U1065 (N_1065,In_2903,In_4144);
or U1066 (N_1066,In_1125,In_4069);
and U1067 (N_1067,In_1489,In_4019);
or U1068 (N_1068,In_4342,In_4893);
or U1069 (N_1069,In_306,In_2755);
or U1070 (N_1070,In_2982,In_3581);
or U1071 (N_1071,In_2310,In_1026);
nor U1072 (N_1072,In_73,In_1982);
and U1073 (N_1073,In_803,In_2286);
or U1074 (N_1074,In_810,In_3101);
nand U1075 (N_1075,In_3251,In_16);
and U1076 (N_1076,In_161,In_4638);
or U1077 (N_1077,In_249,In_3323);
nor U1078 (N_1078,In_2714,In_4409);
and U1079 (N_1079,In_865,In_3087);
nand U1080 (N_1080,In_1700,In_4453);
nor U1081 (N_1081,In_1370,In_19);
and U1082 (N_1082,In_4895,In_3403);
and U1083 (N_1083,In_3448,In_2213);
nor U1084 (N_1084,In_1820,In_4332);
xnor U1085 (N_1085,In_3402,In_1089);
nand U1086 (N_1086,In_2351,In_603);
and U1087 (N_1087,In_4001,In_4032);
nand U1088 (N_1088,In_349,In_4783);
nand U1089 (N_1089,In_227,In_4838);
nor U1090 (N_1090,In_3451,In_3212);
nor U1091 (N_1091,In_4934,In_4609);
nor U1092 (N_1092,In_4078,In_2800);
nand U1093 (N_1093,In_759,In_1612);
nand U1094 (N_1094,In_4441,In_305);
xnor U1095 (N_1095,In_1311,In_967);
or U1096 (N_1096,In_1943,In_1900);
and U1097 (N_1097,In_4709,In_4518);
or U1098 (N_1098,In_2304,In_4189);
nand U1099 (N_1099,In_3002,In_4788);
or U1100 (N_1100,In_4352,In_4302);
nor U1101 (N_1101,In_2633,In_2739);
nand U1102 (N_1102,In_846,In_4533);
xnor U1103 (N_1103,In_197,In_4956);
and U1104 (N_1104,In_1643,In_1650);
nor U1105 (N_1105,In_4478,In_1934);
and U1106 (N_1106,In_3863,In_3232);
xor U1107 (N_1107,In_195,In_2245);
and U1108 (N_1108,In_1570,In_1555);
nor U1109 (N_1109,In_1014,In_620);
and U1110 (N_1110,In_3264,In_3555);
nor U1111 (N_1111,In_4851,In_201);
or U1112 (N_1112,In_660,In_4245);
nor U1113 (N_1113,In_392,In_3594);
nand U1114 (N_1114,In_3395,In_4887);
nand U1115 (N_1115,In_1513,In_4700);
or U1116 (N_1116,In_1793,In_1699);
and U1117 (N_1117,In_3137,In_3246);
and U1118 (N_1118,In_4227,In_641);
and U1119 (N_1119,In_3606,In_4386);
nor U1120 (N_1120,In_2038,In_4839);
nand U1121 (N_1121,In_4420,In_2585);
xor U1122 (N_1122,In_65,In_430);
nand U1123 (N_1123,In_2661,In_3230);
and U1124 (N_1124,In_3852,In_1262);
xor U1125 (N_1125,In_1684,In_1531);
nand U1126 (N_1126,In_3247,In_1254);
and U1127 (N_1127,In_2422,In_1098);
and U1128 (N_1128,In_4203,In_3061);
nand U1129 (N_1129,In_4027,In_4573);
or U1130 (N_1130,In_4630,In_3563);
or U1131 (N_1131,In_2289,In_4111);
or U1132 (N_1132,In_2546,In_3634);
xnor U1133 (N_1133,In_4396,In_2973);
xnor U1134 (N_1134,In_1930,In_1074);
nor U1135 (N_1135,In_2544,In_44);
and U1136 (N_1136,In_4972,In_2632);
and U1137 (N_1137,In_3556,In_4637);
and U1138 (N_1138,In_2029,In_553);
xor U1139 (N_1139,In_3622,In_135);
or U1140 (N_1140,In_2699,In_2050);
and U1141 (N_1141,In_1620,In_2624);
or U1142 (N_1142,In_3353,In_1864);
and U1143 (N_1143,In_1786,In_1597);
nand U1144 (N_1144,In_1537,In_458);
and U1145 (N_1145,In_875,In_298);
or U1146 (N_1146,In_592,In_3687);
nor U1147 (N_1147,In_512,In_3109);
nor U1148 (N_1148,In_1058,In_2865);
nand U1149 (N_1149,In_767,In_1831);
nand U1150 (N_1150,In_1836,In_1217);
and U1151 (N_1151,In_3696,In_191);
nand U1152 (N_1152,In_743,In_3469);
nand U1153 (N_1153,In_969,In_3317);
and U1154 (N_1154,In_2977,In_3839);
nand U1155 (N_1155,In_2500,In_1876);
xnor U1156 (N_1156,In_172,In_1017);
and U1157 (N_1157,In_2605,In_2650);
nor U1158 (N_1158,In_297,In_1720);
or U1159 (N_1159,In_3567,In_2844);
nand U1160 (N_1160,In_3103,In_2861);
nor U1161 (N_1161,In_3940,In_4371);
nor U1162 (N_1162,In_262,In_321);
or U1163 (N_1163,In_1646,In_3261);
or U1164 (N_1164,In_1186,In_574);
nand U1165 (N_1165,In_4962,In_1812);
nor U1166 (N_1166,In_3905,In_4770);
nand U1167 (N_1167,In_2983,In_1809);
and U1168 (N_1168,In_4428,In_2357);
nor U1169 (N_1169,In_2881,In_2998);
and U1170 (N_1170,In_327,In_384);
nand U1171 (N_1171,In_3524,In_423);
nor U1172 (N_1172,In_115,In_15);
nand U1173 (N_1173,In_2468,In_570);
nand U1174 (N_1174,In_4548,In_4993);
and U1175 (N_1175,In_2931,In_3534);
or U1176 (N_1176,In_3312,In_864);
nor U1177 (N_1177,In_2830,In_3493);
nand U1178 (N_1178,In_4122,In_932);
and U1179 (N_1179,In_945,In_2489);
xor U1180 (N_1180,In_3440,In_1059);
xnor U1181 (N_1181,In_1384,In_3310);
xnor U1182 (N_1182,In_4583,In_4135);
nor U1183 (N_1183,In_4931,In_4202);
nand U1184 (N_1184,In_2535,In_729);
or U1185 (N_1185,In_2101,In_41);
and U1186 (N_1186,In_2466,In_4563);
xor U1187 (N_1187,In_2202,In_2008);
xnor U1188 (N_1188,In_2176,In_728);
nand U1189 (N_1189,In_334,In_4459);
xor U1190 (N_1190,In_484,In_2253);
or U1191 (N_1191,In_1640,In_1269);
nand U1192 (N_1192,In_3610,In_3384);
or U1193 (N_1193,In_2530,In_2730);
and U1194 (N_1194,In_1504,In_2041);
or U1195 (N_1195,In_2145,In_2676);
xor U1196 (N_1196,In_995,In_1451);
nor U1197 (N_1197,In_3726,In_4456);
nor U1198 (N_1198,In_3257,In_1922);
or U1199 (N_1199,In_260,In_4349);
nand U1200 (N_1200,In_3260,In_2312);
nor U1201 (N_1201,In_2083,In_1128);
nand U1202 (N_1202,In_1923,In_672);
nor U1203 (N_1203,In_1800,In_3388);
xnor U1204 (N_1204,In_4919,In_3024);
nor U1205 (N_1205,In_4745,In_3528);
nor U1206 (N_1206,In_3295,In_1015);
nor U1207 (N_1207,In_3825,In_3933);
or U1208 (N_1208,In_3170,In_3800);
or U1209 (N_1209,In_340,In_1527);
xnor U1210 (N_1210,In_3164,In_96);
and U1211 (N_1211,In_617,In_3435);
or U1212 (N_1212,In_3036,In_1522);
or U1213 (N_1213,In_855,In_3213);
nand U1214 (N_1214,In_4841,In_3879);
and U1215 (N_1215,In_2457,In_4776);
or U1216 (N_1216,In_2549,In_4946);
and U1217 (N_1217,In_373,In_520);
nor U1218 (N_1218,In_1711,In_3475);
or U1219 (N_1219,In_3605,In_1918);
or U1220 (N_1220,In_3514,In_3368);
nor U1221 (N_1221,In_4107,In_1477);
and U1222 (N_1222,In_1371,In_2654);
nor U1223 (N_1223,In_362,In_21);
nand U1224 (N_1224,In_1261,In_3199);
and U1225 (N_1225,In_2364,In_3813);
xor U1226 (N_1226,In_3009,In_1547);
xnor U1227 (N_1227,In_2389,In_3325);
xor U1228 (N_1228,In_25,In_4722);
or U1229 (N_1229,In_4317,In_876);
and U1230 (N_1230,In_2520,In_3923);
and U1231 (N_1231,In_4220,In_251);
nor U1232 (N_1232,In_1133,In_1754);
nor U1233 (N_1233,In_742,In_2319);
or U1234 (N_1234,In_3651,In_3485);
nor U1235 (N_1235,In_4544,In_4329);
and U1236 (N_1236,In_3586,In_2557);
nand U1237 (N_1237,In_4977,In_3096);
and U1238 (N_1238,In_2235,In_564);
xnor U1239 (N_1239,In_1474,In_4321);
nor U1240 (N_1240,In_4305,In_1270);
or U1241 (N_1241,In_26,In_1424);
xor U1242 (N_1242,In_536,In_1315);
and U1243 (N_1243,In_2341,In_475);
and U1244 (N_1244,In_1243,In_4683);
or U1245 (N_1245,In_2512,In_393);
and U1246 (N_1246,In_350,In_2568);
or U1247 (N_1247,In_4273,In_3180);
nand U1248 (N_1248,In_169,In_1155);
nor U1249 (N_1249,In_941,In_2794);
or U1250 (N_1250,In_4986,In_4015);
nor U1251 (N_1251,In_2231,In_4437);
or U1252 (N_1252,In_3690,In_4664);
xnor U1253 (N_1253,In_1600,In_2479);
xnor U1254 (N_1254,In_4211,In_2045);
nand U1255 (N_1255,In_1410,In_4540);
xnor U1256 (N_1256,In_3253,In_4050);
or U1257 (N_1257,In_3603,In_1332);
nand U1258 (N_1258,In_4794,In_1492);
or U1259 (N_1259,In_268,In_2837);
nand U1260 (N_1260,In_320,In_1306);
xor U1261 (N_1261,In_2812,In_1548);
or U1262 (N_1262,In_2683,In_2838);
nand U1263 (N_1263,In_181,In_928);
and U1264 (N_1264,In_105,In_3281);
or U1265 (N_1265,In_673,In_3242);
nand U1266 (N_1266,In_1996,In_2404);
and U1267 (N_1267,In_2608,In_3473);
nor U1268 (N_1268,In_3471,In_2748);
nand U1269 (N_1269,In_3083,In_4201);
nand U1270 (N_1270,In_1378,In_4012);
or U1271 (N_1271,In_3574,In_3677);
or U1272 (N_1272,In_984,In_14);
xor U1273 (N_1273,In_2958,In_2084);
xor U1274 (N_1274,In_4617,In_2485);
nor U1275 (N_1275,In_4395,In_1381);
nor U1276 (N_1276,In_2111,In_1929);
and U1277 (N_1277,In_1681,In_1744);
and U1278 (N_1278,In_4835,In_1766);
or U1279 (N_1279,In_2246,In_4141);
nor U1280 (N_1280,In_3781,In_2409);
nor U1281 (N_1281,In_3045,In_3811);
nand U1282 (N_1282,In_2892,In_4176);
or U1283 (N_1283,In_4330,In_107);
xnor U1284 (N_1284,In_4837,In_3571);
or U1285 (N_1285,In_4595,In_4855);
nand U1286 (N_1286,In_4212,In_1634);
and U1287 (N_1287,In_1763,In_4020);
or U1288 (N_1288,In_847,In_1392);
and U1289 (N_1289,In_946,In_1706);
nand U1290 (N_1290,In_4455,In_2015);
or U1291 (N_1291,In_285,In_323);
xor U1292 (N_1292,In_2016,In_733);
and U1293 (N_1293,In_3782,In_1642);
nor U1294 (N_1294,In_3842,In_874);
or U1295 (N_1295,In_4351,In_2868);
and U1296 (N_1296,In_1212,In_1397);
xnor U1297 (N_1297,In_4932,In_4698);
and U1298 (N_1298,In_834,In_731);
and U1299 (N_1299,In_407,In_4807);
nor U1300 (N_1300,In_4458,In_2445);
and U1301 (N_1301,In_4013,In_1724);
nor U1302 (N_1302,In_2305,In_4446);
or U1303 (N_1303,In_3544,In_3569);
and U1304 (N_1304,In_3860,In_4761);
nand U1305 (N_1305,In_2376,In_1139);
or U1306 (N_1306,In_2410,In_3517);
nand U1307 (N_1307,In_3342,In_519);
nand U1308 (N_1308,In_4612,In_3073);
nand U1309 (N_1309,In_2968,In_1010);
nand U1310 (N_1310,In_12,In_1372);
or U1311 (N_1311,In_1150,In_2252);
nor U1312 (N_1312,In_521,In_2127);
nand U1313 (N_1313,In_3625,In_3156);
nor U1314 (N_1314,In_205,In_1855);
nor U1315 (N_1315,In_102,In_4687);
nor U1316 (N_1316,In_4087,In_1774);
nand U1317 (N_1317,In_4005,In_1319);
nand U1318 (N_1318,In_4179,In_4890);
and U1319 (N_1319,In_2067,In_1960);
or U1320 (N_1320,In_1145,In_1129);
or U1321 (N_1321,In_4590,In_1796);
or U1322 (N_1322,In_4234,In_3892);
nand U1323 (N_1323,In_1759,In_2360);
nand U1324 (N_1324,In_4818,In_2603);
nor U1325 (N_1325,In_1220,In_3095);
nor U1326 (N_1326,In_1735,In_3717);
or U1327 (N_1327,In_4215,In_3705);
nor U1328 (N_1328,In_2403,In_3128);
and U1329 (N_1329,In_594,In_693);
or U1330 (N_1330,In_3,In_178);
nand U1331 (N_1331,In_3205,In_3420);
or U1332 (N_1332,In_1951,In_3130);
and U1333 (N_1333,In_1967,In_4908);
or U1334 (N_1334,In_2642,In_1770);
nand U1335 (N_1335,In_3832,In_3441);
or U1336 (N_1336,In_2077,In_1420);
nor U1337 (N_1337,In_638,In_4769);
and U1338 (N_1338,In_4088,In_420);
and U1339 (N_1339,In_3596,In_3681);
nand U1340 (N_1340,In_3107,In_3874);
and U1341 (N_1341,In_490,In_4472);
nand U1342 (N_1342,In_2537,In_3195);
or U1343 (N_1343,In_1526,In_4158);
nor U1344 (N_1344,In_2314,In_3108);
xnor U1345 (N_1345,In_2986,In_1536);
and U1346 (N_1346,In_3229,In_2528);
and U1347 (N_1347,In_300,In_1081);
and U1348 (N_1348,In_1997,In_4964);
nor U1349 (N_1349,In_523,In_4735);
nand U1350 (N_1350,In_4787,In_219);
xor U1351 (N_1351,In_4900,In_3838);
nor U1352 (N_1352,In_153,In_2851);
xor U1353 (N_1353,In_346,In_46);
or U1354 (N_1354,In_832,In_3155);
nand U1355 (N_1355,In_2914,In_973);
and U1356 (N_1356,In_4268,In_3748);
or U1357 (N_1357,In_1123,In_2116);
xor U1358 (N_1358,In_2198,In_2342);
or U1359 (N_1359,In_1973,In_1925);
nand U1360 (N_1360,In_238,In_4057);
or U1361 (N_1361,In_4059,In_2775);
nor U1362 (N_1362,In_2904,In_540);
nand U1363 (N_1363,In_3110,In_2250);
or U1364 (N_1364,In_2571,In_444);
nor U1365 (N_1365,In_795,In_3350);
nand U1366 (N_1366,In_4180,In_4236);
nor U1367 (N_1367,In_3611,In_3994);
or U1368 (N_1368,In_3401,In_1084);
xor U1369 (N_1369,In_1227,In_3051);
and U1370 (N_1370,In_1719,In_529);
or U1371 (N_1371,In_843,In_413);
nor U1372 (N_1372,In_1984,In_2227);
nand U1373 (N_1373,In_2678,In_3457);
nand U1374 (N_1374,In_4576,In_4133);
nor U1375 (N_1375,In_4172,In_2226);
or U1376 (N_1376,In_4916,In_3938);
nand U1377 (N_1377,In_2588,In_1329);
or U1378 (N_1378,In_3935,In_904);
xor U1379 (N_1379,In_4582,In_547);
or U1380 (N_1380,In_3254,In_2590);
or U1381 (N_1381,In_1327,In_2778);
and U1382 (N_1382,In_4357,In_4334);
xnor U1383 (N_1383,In_164,In_311);
xnor U1384 (N_1384,In_2094,In_404);
nand U1385 (N_1385,In_2779,In_1892);
nor U1386 (N_1386,In_4779,In_3789);
xor U1387 (N_1387,In_1179,In_3598);
and U1388 (N_1388,In_3158,In_495);
nor U1389 (N_1389,In_4000,In_6);
nor U1390 (N_1390,In_500,In_3897);
and U1391 (N_1391,In_4707,In_4307);
or U1392 (N_1392,In_605,In_3648);
nand U1393 (N_1393,In_1353,In_432);
xor U1394 (N_1394,In_3282,In_3801);
and U1395 (N_1395,In_717,In_3149);
xor U1396 (N_1396,In_766,In_1194);
nand U1397 (N_1397,In_2220,In_4182);
and U1398 (N_1398,In_2042,In_3805);
xor U1399 (N_1399,In_4483,In_756);
nand U1400 (N_1400,In_4131,In_2135);
and U1401 (N_1401,In_2886,In_965);
nand U1402 (N_1402,In_190,In_2713);
and U1403 (N_1403,In_3769,In_111);
or U1404 (N_1404,In_2138,In_3019);
and U1405 (N_1405,In_3911,In_1242);
nor U1406 (N_1406,In_1907,In_1539);
nand U1407 (N_1407,In_2869,In_3560);
xnor U1408 (N_1408,In_4695,In_4832);
or U1409 (N_1409,In_2871,In_3438);
or U1410 (N_1410,In_4556,In_3623);
nor U1411 (N_1411,In_3760,In_1528);
nor U1412 (N_1412,In_894,In_3238);
nor U1413 (N_1413,In_3535,In_3736);
nor U1414 (N_1414,In_3357,In_2151);
and U1415 (N_1415,In_4685,In_1478);
and U1416 (N_1416,In_3421,In_4448);
nor U1417 (N_1417,In_4256,In_2679);
nor U1418 (N_1418,In_2737,In_1945);
nor U1419 (N_1419,In_1120,In_1461);
and U1420 (N_1420,In_2897,In_3043);
xor U1421 (N_1421,In_1532,In_1447);
nand U1422 (N_1422,In_2762,In_1149);
and U1423 (N_1423,In_1788,In_1516);
nand U1424 (N_1424,In_2617,In_2329);
and U1425 (N_1425,In_2760,In_3589);
nor U1426 (N_1426,In_1265,In_415);
or U1427 (N_1427,In_2320,In_4767);
nand U1428 (N_1428,In_4680,In_4479);
or U1429 (N_1429,In_282,In_1886);
or U1430 (N_1430,In_4520,In_3695);
nand U1431 (N_1431,In_4812,In_3052);
and U1432 (N_1432,In_2860,In_2035);
and U1433 (N_1433,In_1488,In_2207);
nor U1434 (N_1434,In_4723,In_4874);
or U1435 (N_1435,In_3414,In_1927);
and U1436 (N_1436,In_582,In_3547);
nor U1437 (N_1437,In_1404,In_1963);
nor U1438 (N_1438,In_2655,In_29);
or U1439 (N_1439,In_1592,In_1338);
or U1440 (N_1440,In_4337,In_4597);
nor U1441 (N_1441,In_4505,In_290);
nand U1442 (N_1442,In_1839,In_794);
xnor U1443 (N_1443,In_1937,In_3039);
xnor U1444 (N_1444,In_3293,In_4833);
and U1445 (N_1445,In_4933,In_2583);
nor U1446 (N_1446,In_2709,In_3561);
or U1447 (N_1447,In_4869,In_240);
or U1448 (N_1448,In_4581,In_167);
xnor U1449 (N_1449,In_189,In_1617);
or U1450 (N_1450,In_368,In_4781);
and U1451 (N_1451,In_3730,In_3303);
and U1452 (N_1452,In_790,In_86);
xor U1453 (N_1453,In_3962,In_1364);
nor U1454 (N_1454,In_3065,In_3576);
or U1455 (N_1455,In_1395,In_2935);
nand U1456 (N_1456,In_4952,In_608);
nor U1457 (N_1457,In_1789,In_3086);
nor U1458 (N_1458,In_1233,In_4966);
nor U1459 (N_1459,In_4258,In_1073);
or U1460 (N_1460,In_1020,In_1919);
or U1461 (N_1461,In_3829,In_39);
nor U1462 (N_1462,In_209,In_3872);
or U1463 (N_1463,In_2876,In_382);
and U1464 (N_1464,In_1619,In_3348);
and U1465 (N_1465,In_4795,In_416);
or U1466 (N_1466,In_3189,In_722);
nand U1467 (N_1467,In_3134,In_3025);
nand U1468 (N_1468,In_2966,In_1361);
and U1469 (N_1469,In_2667,In_3382);
or U1470 (N_1470,In_1797,In_2236);
and U1471 (N_1471,In_3223,In_4185);
and U1472 (N_1472,In_3047,In_1304);
and U1473 (N_1473,In_4953,In_915);
nor U1474 (N_1474,In_1382,In_3809);
and U1475 (N_1475,In_2929,In_3489);
nand U1476 (N_1476,In_2412,In_2080);
nor U1477 (N_1477,In_1198,In_2014);
nand U1478 (N_1478,In_1415,In_1421);
nand U1479 (N_1479,In_374,In_801);
nor U1480 (N_1480,In_3472,In_1280);
or U1481 (N_1481,In_3913,In_4094);
nand U1482 (N_1482,In_1036,In_3771);
and U1483 (N_1483,In_2031,In_3409);
and U1484 (N_1484,In_4118,In_4706);
nand U1485 (N_1485,In_3337,In_3762);
nor U1486 (N_1486,In_4260,In_2652);
nor U1487 (N_1487,In_425,In_217);
nand U1488 (N_1488,In_3363,In_4689);
nor U1489 (N_1489,In_1373,In_4021);
nor U1490 (N_1490,In_1671,In_2694);
nor U1491 (N_1491,In_4545,In_2472);
and U1492 (N_1492,In_3768,In_4108);
nor U1493 (N_1493,In_925,In_3904);
nor U1494 (N_1494,In_3980,In_1288);
nor U1495 (N_1495,In_4286,In_905);
nor U1496 (N_1496,In_1287,In_347);
nor U1497 (N_1497,In_4353,In_3954);
nand U1498 (N_1498,In_829,In_3869);
nor U1499 (N_1499,In_3390,In_3820);
nor U1500 (N_1500,In_1819,In_3944);
nor U1501 (N_1501,In_277,In_550);
or U1502 (N_1502,In_2239,In_4830);
nand U1503 (N_1503,In_4161,In_545);
xor U1504 (N_1504,In_3883,In_2142);
or U1505 (N_1505,In_154,In_1638);
or U1506 (N_1506,In_71,In_4805);
and U1507 (N_1507,In_3076,In_1644);
or U1508 (N_1508,In_2992,In_1061);
or U1509 (N_1509,In_2139,In_1437);
nand U1510 (N_1510,In_4318,In_3500);
nor U1511 (N_1511,In_739,In_1412);
xnor U1512 (N_1512,In_1880,In_1501);
nand U1513 (N_1513,In_2159,In_1005);
or U1514 (N_1514,In_2056,In_715);
nor U1515 (N_1515,In_3429,In_3592);
nor U1516 (N_1516,In_4495,In_3550);
or U1517 (N_1517,In_3828,In_381);
nor U1518 (N_1518,In_977,In_3880);
nor U1519 (N_1519,In_451,In_1563);
nor U1520 (N_1520,In_2900,In_4552);
nand U1521 (N_1521,In_131,In_1360);
or U1522 (N_1522,In_4570,In_3464);
xor U1523 (N_1523,In_3908,In_649);
or U1524 (N_1524,In_3332,In_1823);
or U1525 (N_1525,In_4992,In_2809);
nand U1526 (N_1526,In_887,In_2543);
nand U1527 (N_1527,In_708,In_538);
or U1528 (N_1528,In_2467,In_3334);
nand U1529 (N_1529,In_4261,In_1197);
nor U1530 (N_1530,In_1151,In_1162);
xor U1531 (N_1531,In_1260,In_4568);
and U1532 (N_1532,In_1631,In_3183);
nor U1533 (N_1533,In_1777,In_3106);
and U1534 (N_1534,In_2785,In_1004);
or U1535 (N_1535,In_988,In_4079);
and U1536 (N_1536,In_3548,In_2284);
nand U1537 (N_1537,In_797,In_3011);
or U1538 (N_1538,In_2398,In_3376);
and U1539 (N_1539,In_2308,In_3405);
or U1540 (N_1540,In_4364,In_1211);
and U1541 (N_1541,In_4922,In_2167);
and U1542 (N_1542,In_3419,In_4328);
or U1543 (N_1543,In_2443,In_515);
nor U1544 (N_1544,In_888,In_4971);
or U1545 (N_1545,In_4299,In_3668);
or U1546 (N_1546,In_1928,In_1808);
and U1547 (N_1547,In_2275,In_827);
nand U1548 (N_1548,In_3460,In_2063);
or U1549 (N_1549,In_3374,In_3028);
and U1550 (N_1550,In_513,In_3185);
xnor U1551 (N_1551,In_3656,In_234);
and U1552 (N_1552,In_1368,In_4209);
or U1553 (N_1553,In_4037,In_4517);
nor U1554 (N_1554,In_1851,In_840);
or U1555 (N_1555,In_4594,In_3022);
nand U1556 (N_1556,In_611,In_3072);
nor U1557 (N_1557,In_3833,In_3506);
nor U1558 (N_1558,In_2726,In_3522);
nor U1559 (N_1559,In_1568,In_2527);
and U1560 (N_1560,In_2789,In_3078);
nand U1561 (N_1561,In_1881,In_2374);
nand U1562 (N_1562,In_4886,In_853);
nor U1563 (N_1563,In_2956,In_4828);
nor U1564 (N_1564,In_4442,In_3265);
nor U1565 (N_1565,In_3218,In_3091);
nor U1566 (N_1566,In_395,In_3895);
or U1567 (N_1567,In_2555,In_3320);
xor U1568 (N_1568,In_789,In_1884);
or U1569 (N_1569,In_53,In_4604);
nand U1570 (N_1570,In_4632,In_950);
nand U1571 (N_1571,In_3646,In_4994);
and U1572 (N_1572,In_4247,In_4257);
nand U1573 (N_1573,In_1182,In_1803);
nand U1574 (N_1574,In_184,In_1741);
nand U1575 (N_1575,In_4068,In_1011);
xnor U1576 (N_1576,In_2940,In_4642);
nand U1577 (N_1577,In_3124,In_3145);
nor U1578 (N_1578,In_3617,In_3971);
nor U1579 (N_1579,In_2519,In_994);
and U1580 (N_1580,In_4208,In_2516);
or U1581 (N_1581,In_1507,In_4679);
nor U1582 (N_1582,In_3711,In_2425);
or U1583 (N_1583,In_2334,In_2196);
or U1584 (N_1584,In_4183,In_3141);
nor U1585 (N_1585,In_1247,In_4861);
nor U1586 (N_1586,In_3316,In_1335);
nor U1587 (N_1587,In_1544,In_2920);
nand U1588 (N_1588,In_3466,In_3551);
nor U1589 (N_1589,In_1623,In_204);
xor U1590 (N_1590,In_4853,In_972);
nor U1591 (N_1591,In_1167,In_232);
nand U1592 (N_1592,In_4106,In_3370);
nor U1593 (N_1593,In_1137,In_38);
nand U1594 (N_1594,In_67,In_4259);
xor U1595 (N_1595,In_1240,In_4644);
nor U1596 (N_1596,In_3436,In_4587);
or U1597 (N_1597,In_3666,In_3287);
and U1598 (N_1598,In_4206,In_817);
or U1599 (N_1599,In_3674,In_4431);
nand U1600 (N_1600,In_4822,In_4654);
xnor U1601 (N_1601,In_852,In_2406);
nand U1602 (N_1602,In_1577,In_2622);
or U1603 (N_1603,In_3160,In_4011);
nand U1604 (N_1604,In_3006,In_487);
nand U1605 (N_1605,In_751,In_27);
nand U1606 (N_1606,In_4626,In_258);
and U1607 (N_1607,In_3901,In_2499);
and U1608 (N_1608,In_230,In_4536);
nand U1609 (N_1609,In_1130,In_893);
or U1610 (N_1610,In_7,In_3798);
or U1611 (N_1611,In_3349,In_2805);
and U1612 (N_1612,In_654,In_4744);
nand U1613 (N_1613,In_125,In_3034);
nor U1614 (N_1614,In_480,In_3214);
nand U1615 (N_1615,In_3070,In_1175);
or U1616 (N_1616,In_2649,In_1980);
xnor U1617 (N_1617,In_3454,In_909);
nor U1618 (N_1618,In_3510,In_949);
or U1619 (N_1619,In_304,In_1983);
nor U1620 (N_1620,In_1352,In_1246);
nand U1621 (N_1621,In_3553,In_1621);
or U1622 (N_1622,In_2824,In_245);
nand U1623 (N_1623,In_1533,In_2684);
nor U1624 (N_1624,In_1092,In_606);
and U1625 (N_1625,In_3968,In_1115);
and U1626 (N_1626,In_610,In_2338);
or U1627 (N_1627,In_367,In_3773);
nor U1628 (N_1628,In_3346,In_2395);
nand U1629 (N_1629,In_151,In_4802);
or U1630 (N_1630,In_4018,In_3347);
nor U1631 (N_1631,In_3341,In_4002);
and U1632 (N_1632,In_1965,In_1245);
nor U1633 (N_1633,In_2430,In_1854);
and U1634 (N_1634,In_3984,In_2294);
and U1635 (N_1635,In_3148,In_1511);
nand U1636 (N_1636,In_1857,In_3094);
nand U1637 (N_1637,In_3064,In_91);
nor U1638 (N_1638,In_1659,In_3187);
and U1639 (N_1639,In_4884,In_648);
nor U1640 (N_1640,In_1173,In_4091);
and U1641 (N_1641,In_1727,In_242);
nand U1642 (N_1642,In_3990,In_1131);
nor U1643 (N_1643,In_1889,In_2898);
nand U1644 (N_1644,In_1289,In_1872);
nand U1645 (N_1645,In_732,In_1932);
nor U1646 (N_1646,In_1436,In_1266);
and U1647 (N_1647,In_48,In_3599);
or U1648 (N_1648,In_2665,In_2733);
and U1649 (N_1649,In_3698,In_2511);
xor U1650 (N_1650,In_4743,In_3151);
or U1651 (N_1651,In_1515,In_2322);
and U1652 (N_1652,In_1495,In_4314);
or U1653 (N_1653,In_4593,In_4649);
xor U1654 (N_1654,In_4980,In_3365);
nor U1655 (N_1655,In_4960,In_4414);
nand U1656 (N_1656,In_1704,In_3792);
nor U1657 (N_1657,In_1166,In_4639);
or U1658 (N_1658,In_2503,In_1994);
or U1659 (N_1659,In_1966,In_1552);
nor U1660 (N_1660,In_4578,In_822);
nand U1661 (N_1661,In_4188,In_2598);
and U1662 (N_1662,In_2424,In_1303);
nand U1663 (N_1663,In_2670,In_528);
nand U1664 (N_1664,In_3118,In_3533);
and U1665 (N_1665,In_3770,In_4285);
nand U1666 (N_1666,In_2564,In_3367);
or U1667 (N_1667,In_370,In_609);
xor U1668 (N_1668,In_804,In_2581);
xor U1669 (N_1669,In_1690,In_4112);
nor U1670 (N_1670,In_4817,In_3734);
nor U1671 (N_1671,In_1921,In_1790);
nand U1672 (N_1672,In_3111,In_2764);
or U1673 (N_1673,In_1733,In_1582);
or U1674 (N_1674,In_3794,In_773);
and U1675 (N_1675,In_656,In_4333);
or U1676 (N_1676,In_4620,In_1112);
and U1677 (N_1677,In_394,In_1944);
and U1678 (N_1678,In_1022,In_819);
nor U1679 (N_1679,In_4763,In_1106);
nand U1680 (N_1680,In_3416,In_3579);
nor U1681 (N_1681,In_3296,In_1174);
nor U1682 (N_1682,In_3399,In_3049);
nor U1683 (N_1683,In_2229,In_1213);
nand U1684 (N_1684,In_1614,In_583);
or U1685 (N_1685,In_707,In_3788);
or U1686 (N_1686,In_2949,In_2186);
nand U1687 (N_1687,In_4510,In_4677);
and U1688 (N_1688,In_3434,In_332);
nor U1689 (N_1689,In_3433,In_4323);
or U1690 (N_1690,In_1626,In_1039);
xor U1691 (N_1691,In_4049,In_248);
nand U1692 (N_1692,In_1950,In_2057);
nor U1693 (N_1693,In_2704,In_963);
nand U1694 (N_1694,In_4496,In_408);
nor U1695 (N_1695,In_1218,In_1);
and U1696 (N_1696,In_3823,In_830);
or U1697 (N_1697,In_3896,In_639);
xnor U1698 (N_1698,In_2110,In_563);
nand U1699 (N_1699,In_2323,In_3252);
and U1700 (N_1700,In_1100,In_4237);
nor U1701 (N_1701,In_2382,In_4571);
or U1702 (N_1702,In_3865,In_4963);
nand U1703 (N_1703,In_2877,In_2593);
nor U1704 (N_1704,In_3876,In_2573);
or U1705 (N_1705,In_2048,In_3582);
and U1706 (N_1706,In_2011,In_1031);
nor U1707 (N_1707,In_3062,In_4465);
and U1708 (N_1708,In_2908,In_1686);
nor U1709 (N_1709,In_3946,In_319);
and U1710 (N_1710,In_1336,In_112);
xor U1711 (N_1711,In_2715,In_838);
xnor U1712 (N_1712,In_2333,In_680);
nor U1713 (N_1713,In_1710,In_1316);
nor U1714 (N_1714,In_4071,In_4547);
nand U1715 (N_1715,In_1703,In_1009);
nand U1716 (N_1716,In_4098,In_1302);
nand U1717 (N_1717,In_2193,In_4128);
nor U1718 (N_1718,In_3116,In_2146);
nand U1719 (N_1719,In_4173,In_1158);
or U1720 (N_1720,In_2957,In_580);
nor U1721 (N_1721,In_1309,In_685);
nor U1722 (N_1722,In_3040,In_2327);
or U1723 (N_1723,In_2795,In_1497);
or U1724 (N_1724,In_2753,In_1557);
and U1725 (N_1725,In_1815,In_2155);
nand U1726 (N_1726,In_4218,In_3177);
nor U1727 (N_1727,In_1147,In_956);
or U1728 (N_1728,In_4691,In_2911);
xnor U1729 (N_1729,In_4426,In_2251);
and U1730 (N_1730,In_3702,In_791);
nor U1731 (N_1731,In_4847,In_926);
nor U1732 (N_1732,In_3754,In_399);
nand U1733 (N_1733,In_1430,In_1972);
xnor U1734 (N_1734,In_4834,In_1114);
xnor U1735 (N_1735,In_1958,In_1253);
nor U1736 (N_1736,In_2732,In_3509);
nor U1737 (N_1737,In_4566,In_3121);
xor U1738 (N_1738,In_3099,In_40);
or U1739 (N_1739,In_4621,In_616);
nand U1740 (N_1740,In_4857,In_4823);
nor U1741 (N_1741,In_4596,In_3706);
nand U1742 (N_1742,In_2619,In_2890);
and U1743 (N_1743,In_556,In_1611);
nand U1744 (N_1744,In_3412,In_2999);
and U1745 (N_1745,In_873,In_1163);
and U1746 (N_1746,In_280,In_87);
nand U1747 (N_1747,In_4290,In_3267);
nor U1748 (N_1748,In_3354,In_3680);
nor U1749 (N_1749,In_1989,In_2965);
nor U1750 (N_1750,In_1757,In_122);
or U1751 (N_1751,In_4217,In_4457);
nand U1752 (N_1752,In_4584,In_224);
nand U1753 (N_1753,In_2194,In_1366);
nor U1754 (N_1754,In_2930,In_2032);
or U1755 (N_1755,In_3204,In_2806);
nand U1756 (N_1756,In_2129,In_4729);
nand U1757 (N_1757,In_3497,In_2974);
nor U1758 (N_1758,In_3516,In_3602);
nor U1759 (N_1759,In_1363,In_1641);
and U1760 (N_1760,In_1389,In_463);
nand U1761 (N_1761,In_4996,In_4605);
xor U1762 (N_1762,In_4327,In_2915);
nand U1763 (N_1763,In_3965,In_2839);
nor U1764 (N_1764,In_3536,In_821);
nor U1765 (N_1765,In_1468,In_2458);
nor U1766 (N_1766,In_1423,In_3783);
and U1767 (N_1767,In_1827,In_727);
or U1768 (N_1768,In_990,In_481);
or U1769 (N_1769,In_725,In_4615);
nand U1770 (N_1770,In_2272,In_526);
or U1771 (N_1771,In_4279,In_310);
and U1772 (N_1772,In_397,In_2574);
or U1773 (N_1773,In_2263,In_1259);
nor U1774 (N_1774,In_4589,In_4293);
nor U1775 (N_1775,In_2055,In_4092);
and U1776 (N_1776,In_4301,In_4061);
and U1777 (N_1777,In_3311,In_3431);
nand U1778 (N_1778,In_3609,In_3112);
xnor U1779 (N_1779,In_4990,In_4710);
or U1780 (N_1780,In_1940,In_3692);
xor U1781 (N_1781,In_1480,In_4815);
or U1782 (N_1782,In_2551,In_4486);
or U1783 (N_1783,In_4493,In_3890);
or U1784 (N_1784,In_3637,In_546);
or U1785 (N_1785,In_4843,In_3056);
or U1786 (N_1786,In_3418,In_2071);
and U1787 (N_1787,In_3704,In_3069);
xor U1788 (N_1788,In_4046,In_1779);
nor U1789 (N_1789,In_74,In_3812);
and U1790 (N_1790,In_754,In_1252);
or U1791 (N_1791,In_4424,In_4072);
nand U1792 (N_1792,In_4413,In_845);
xor U1793 (N_1793,In_1605,In_1502);
or U1794 (N_1794,In_2553,In_3973);
xnor U1795 (N_1795,In_312,In_511);
nor U1796 (N_1796,In_2681,In_1903);
nand U1797 (N_1797,In_4878,In_1813);
nor U1798 (N_1798,In_3531,In_3432);
and U1799 (N_1799,In_4978,In_4870);
nand U1800 (N_1800,In_3630,In_1498);
nor U1801 (N_1801,In_2786,In_575);
or U1802 (N_1802,In_2297,In_1916);
and U1803 (N_1803,In_2776,In_483);
nand U1804 (N_1804,In_1369,In_2303);
nor U1805 (N_1805,In_3301,In_4381);
and U1806 (N_1806,In_2307,In_2591);
xor U1807 (N_1807,In_738,In_4840);
or U1808 (N_1808,In_4338,In_3523);
and U1809 (N_1809,In_2079,In_462);
and U1810 (N_1810,In_314,In_694);
or U1811 (N_1811,In_2866,In_3791);
nor U1812 (N_1812,In_389,In_666);
or U1813 (N_1813,In_2122,In_4987);
or U1814 (N_1814,In_1756,In_823);
nand U1815 (N_1815,In_4471,In_1845);
nor U1816 (N_1816,In_1054,In_1455);
xor U1817 (N_1817,In_121,In_2697);
or U1818 (N_1818,In_779,In_4562);
or U1819 (N_1819,In_2124,In_559);
or U1820 (N_1820,In_891,In_3991);
nand U1821 (N_1821,In_4378,In_2405);
and U1822 (N_1822,In_2847,In_2853);
nand U1823 (N_1823,In_3732,In_4450);
and U1824 (N_1824,In_764,In_2981);
and U1825 (N_1825,In_2599,In_2970);
nand U1826 (N_1826,In_4384,In_3225);
xor U1827 (N_1827,In_2278,In_1427);
nand U1828 (N_1828,In_11,In_2000);
nand U1829 (N_1829,In_3855,In_1588);
and U1830 (N_1830,In_3053,In_353);
or U1831 (N_1831,In_4939,In_1449);
and U1832 (N_1832,In_4829,In_4523);
and U1833 (N_1833,In_4421,In_4170);
nand U1834 (N_1834,In_954,In_2150);
nor U1835 (N_1835,In_2047,In_2701);
and U1836 (N_1836,In_3492,In_1072);
and U1837 (N_1837,In_3174,In_4866);
or U1838 (N_1838,In_2509,In_532);
or U1839 (N_1839,In_555,In_3836);
and U1840 (N_1840,In_4602,In_614);
nand U1841 (N_1841,In_3249,In_1388);
or U1842 (N_1842,In_1586,In_4750);
nand U1843 (N_1843,In_3627,In_1859);
nor U1844 (N_1844,In_2408,In_910);
and U1845 (N_1845,In_159,In_446);
or U1846 (N_1846,In_4813,In_989);
nand U1847 (N_1847,In_143,In_2330);
or U1848 (N_1848,In_1546,In_4755);
nand U1849 (N_1849,In_4693,In_3240);
nand U1850 (N_1850,In_3162,In_724);
nand U1851 (N_1851,In_697,In_2449);
xor U1852 (N_1852,In_1177,In_1285);
nor U1853 (N_1853,In_1541,In_3176);
and U1854 (N_1854,In_1749,In_192);
nand U1855 (N_1855,In_4935,In_1231);
nor U1856 (N_1856,In_3975,In_1161);
nor U1857 (N_1857,In_2223,In_2287);
or U1858 (N_1858,In_3482,In_4023);
or U1859 (N_1859,In_2396,In_3449);
nor U1860 (N_1860,In_2771,In_2362);
nor U1861 (N_1861,In_58,In_4229);
xnor U1862 (N_1862,In_4075,In_4086);
nor U1863 (N_1863,In_699,In_1566);
nand U1864 (N_1864,In_936,In_1399);
or U1865 (N_1865,In_4502,In_3146);
xor U1866 (N_1866,In_274,In_406);
nor U1867 (N_1867,In_3345,In_3291);
xor U1868 (N_1868,In_4115,In_4363);
and U1869 (N_1869,In_1007,In_4263);
nor U1870 (N_1870,In_3513,In_3850);
nor U1871 (N_1871,In_1400,In_2766);
xor U1872 (N_1872,In_4622,In_3837);
nor U1873 (N_1873,In_4230,In_137);
nor U1874 (N_1874,In_4650,In_2541);
or U1875 (N_1875,In_2584,In_1785);
and U1876 (N_1876,In_3804,In_2461);
xnor U1877 (N_1877,In_508,In_2190);
xor U1878 (N_1878,In_1599,In_4366);
or U1879 (N_1879,In_2842,In_1083);
nor U1880 (N_1880,In_3899,In_2994);
nand U1881 (N_1881,In_3615,In_2416);
nand U1882 (N_1882,In_4387,In_3557);
or U1883 (N_1883,In_4316,In_3397);
or U1884 (N_1884,In_3882,In_2277);
nand U1885 (N_1885,In_427,In_4816);
or U1886 (N_1886,In_2230,In_3846);
and U1887 (N_1887,In_3580,In_2020);
xnor U1888 (N_1888,In_2711,In_1822);
nand U1889 (N_1889,In_3197,In_3092);
and U1890 (N_1890,In_3123,In_1172);
and U1891 (N_1891,In_2907,In_466);
nor U1892 (N_1892,In_2997,In_3504);
or U1893 (N_1893,In_4991,In_872);
nor U1894 (N_1894,In_299,In_402);
nor U1895 (N_1895,In_3922,In_1143);
xnor U1896 (N_1896,In_1414,In_439);
nand U1897 (N_1897,In_4725,In_2420);
and U1898 (N_1898,In_2782,In_1713);
xnor U1899 (N_1899,In_1505,In_569);
nor U1900 (N_1900,In_944,In_4522);
xor U1901 (N_1901,In_982,In_336);
and U1902 (N_1902,In_539,In_4310);
and U1903 (N_1903,In_674,In_2180);
and U1904 (N_1904,In_808,In_2513);
nand U1905 (N_1905,In_1975,In_1610);
nor U1906 (N_1906,In_279,In_2274);
or U1907 (N_1907,In_4,In_4080);
and U1908 (N_1908,In_4365,In_2734);
nor U1909 (N_1909,In_640,In_3956);
or U1910 (N_1910,In_3147,In_2855);
xor U1911 (N_1911,In_2005,In_4309);
xnor U1912 (N_1912,In_3235,In_2068);
nand U1913 (N_1913,In_3498,In_1630);
nor U1914 (N_1914,In_3270,In_2460);
nor U1915 (N_1915,In_343,In_4222);
and U1916 (N_1916,In_4792,In_3640);
or U1917 (N_1917,In_3793,In_3779);
or U1918 (N_1918,In_4826,In_4120);
or U1919 (N_1919,In_543,In_4298);
and U1920 (N_1920,In_2978,In_1209);
or U1921 (N_1921,In_3727,In_3054);
nand U1922 (N_1922,In_1008,In_1205);
xor U1923 (N_1923,In_1033,In_1219);
xnor U1924 (N_1924,In_721,In_3930);
or U1925 (N_1925,In_3125,In_1159);
and U1926 (N_1926,In_4635,In_4734);
xnor U1927 (N_1927,In_981,In_2292);
or U1928 (N_1928,In_625,In_2820);
nor U1929 (N_1929,In_1778,In_2944);
nor U1930 (N_1930,In_179,In_4577);
or U1931 (N_1931,In_3298,In_1559);
nand U1932 (N_1932,In_1569,In_1238);
nor U1933 (N_1933,In_3559,In_2113);
nand U1934 (N_1934,In_364,In_1223);
and U1935 (N_1935,In_3948,In_4831);
nand U1936 (N_1936,In_2979,In_2565);
nor U1937 (N_1937,In_1608,In_1587);
and U1938 (N_1938,In_1988,In_4276);
nand U1939 (N_1939,In_3635,In_637);
nor U1940 (N_1940,In_1094,In_3999);
xnor U1941 (N_1941,In_357,In_4747);
xnor U1942 (N_1942,In_879,In_2118);
or U1943 (N_1943,In_4255,In_930);
xor U1944 (N_1944,In_4957,In_2801);
and U1945 (N_1945,In_4611,In_1281);
nand U1946 (N_1946,In_3958,In_1639);
xor U1947 (N_1947,In_1464,In_1618);
nand U1948 (N_1948,In_358,In_4320);
nand U1949 (N_1949,In_4231,In_301);
nor U1950 (N_1950,In_2475,In_2218);
or U1951 (N_1951,In_335,In_3939);
or U1952 (N_1952,In_3262,In_3192);
and U1953 (N_1953,In_709,In_2729);
and U1954 (N_1954,In_4477,In_3315);
nand U1955 (N_1955,In_2388,In_2754);
and U1956 (N_1956,In_1904,In_2780);
nand U1957 (N_1957,In_3978,In_4103);
nor U1958 (N_1958,In_1263,In_607);
nor U1959 (N_1959,In_37,In_4999);
nand U1960 (N_1960,In_793,In_2214);
or U1961 (N_1961,In_239,In_4647);
xor U1962 (N_1962,In_730,In_2375);
nand U1963 (N_1963,In_1116,In_2017);
or U1964 (N_1964,In_1874,In_923);
nand U1965 (N_1965,In_247,In_2120);
or U1966 (N_1966,In_1387,In_3220);
nand U1967 (N_1967,In_3682,In_4512);
or U1968 (N_1968,In_1201,In_1367);
or U1969 (N_1969,In_2773,In_2616);
and U1970 (N_1970,In_2328,In_98);
nor U1971 (N_1971,In_2521,In_4511);
or U1972 (N_1972,In_2073,In_168);
and U1973 (N_1973,In_4757,In_4546);
nor U1974 (N_1974,In_3530,In_531);
nand U1975 (N_1975,In_1298,In_4740);
and U1976 (N_1976,In_2037,In_1807);
and U1977 (N_1977,In_3795,In_3465);
or U1978 (N_1978,In_4981,In_1241);
nor U1979 (N_1979,In_2534,In_2576);
and U1980 (N_1980,In_2854,In_4408);
nor U1981 (N_1981,In_1654,In_943);
nor U1982 (N_1982,In_1107,In_4403);
nand U1983 (N_1983,In_4871,In_435);
xnor U1984 (N_1984,In_669,In_1053);
or U1985 (N_1985,In_2751,In_4876);
and U1986 (N_1986,In_2089,In_471);
nand U1987 (N_1987,In_2542,In_3236);
nand U1988 (N_1988,In_2311,In_3044);
and U1989 (N_1989,In_4973,In_3259);
nand U1990 (N_1990,In_3521,In_4225);
or U1991 (N_1991,In_3735,In_1835);
nor U1992 (N_1992,In_883,In_1987);
nand U1993 (N_1993,In_3190,In_1603);
or U1994 (N_1994,In_4053,In_632);
nand U1995 (N_1995,In_4660,In_36);
xor U1996 (N_1996,In_1416,In_3758);
nand U1997 (N_1997,In_2686,In_3487);
nand U1998 (N_1998,In_806,In_2717);
and U1999 (N_1999,In_2793,In_826);
or U2000 (N_2000,In_1647,In_2279);
nand U2001 (N_2001,In_2763,In_4673);
or U2002 (N_2002,In_3159,In_2887);
and U2003 (N_2003,In_3117,In_3718);
and U2004 (N_2004,In_1152,In_3527);
nand U2005 (N_2005,In_2264,In_4569);
nand U2006 (N_2006,In_2254,In_2863);
nand U2007 (N_2007,In_2078,In_3483);
or U2008 (N_2008,In_4419,In_3562);
and U2009 (N_2009,In_3636,In_2368);
nor U2010 (N_2010,In_4196,In_1087);
nand U2011 (N_2011,In_4370,In_3330);
nand U2012 (N_2012,In_3866,In_142);
or U2013 (N_2013,In_2625,In_2436);
xnor U2014 (N_2014,In_4610,In_4427);
or U2015 (N_2015,In_2160,In_2007);
nor U2016 (N_2016,In_4243,In_3894);
and U2017 (N_2017,In_4124,In_3450);
nand U2018 (N_2018,In_866,In_1664);
or U2019 (N_2019,In_2411,In_1651);
nor U2020 (N_2020,In_3941,In_4877);
or U2021 (N_2021,In_3408,In_3953);
and U2022 (N_2022,In_4608,In_450);
nand U2023 (N_2023,In_2925,In_4412);
nor U2024 (N_2024,In_787,In_1334);
and U2025 (N_2025,In_60,In_4207);
or U2026 (N_2026,In_109,In_1331);
and U2027 (N_2027,In_322,In_4004);
nor U2028 (N_2028,In_2885,In_2783);
xor U2029 (N_2029,In_3983,In_704);
or U2030 (N_2030,In_4372,In_4132);
xnor U2031 (N_2031,In_745,In_2723);
nand U2032 (N_2032,In_869,In_1431);
xnor U2033 (N_2033,In_4484,In_1063);
xor U2034 (N_2034,In_4726,In_2426);
or U2035 (N_2035,In_4265,In_2945);
nor U2036 (N_2036,In_3776,In_2012);
and U2037 (N_2037,In_711,In_4737);
and U2038 (N_2038,In_1841,In_3082);
and U2039 (N_2039,In_4340,In_4460);
nand U2040 (N_2040,In_2698,In_595);
or U2041 (N_2041,In_3097,In_317);
nand U2042 (N_2042,In_1056,In_4445);
nand U2043 (N_2043,In_3135,In_316);
nor U2044 (N_2044,In_4634,In_2054);
or U2045 (N_2045,In_1666,In_3119);
or U2046 (N_2046,In_1898,In_3276);
nand U2047 (N_2047,In_4657,In_2402);
or U2048 (N_2048,In_1899,In_2497);
and U2049 (N_2049,In_4711,In_4010);
and U2050 (N_2050,In_899,In_3871);
nor U2051 (N_2051,In_3808,In_4777);
or U2052 (N_2052,In_4880,In_18);
and U2053 (N_2053,In_4542,In_363);
or U2054 (N_2054,In_3963,In_1970);
nand U2055 (N_2055,In_4275,In_4574);
or U2056 (N_2056,In_1458,In_4168);
nand U2057 (N_2057,In_541,In_2941);
xor U2058 (N_2058,In_3893,In_1082);
or U2059 (N_2059,In_2891,In_4468);
or U2060 (N_2060,In_1905,In_3355);
nor U2061 (N_2061,In_3314,In_2816);
nand U2062 (N_2062,In_3857,In_2586);
nor U2063 (N_2063,In_2618,In_800);
xor U2064 (N_2064,In_493,In_2572);
nor U2065 (N_2065,In_2049,In_3445);
or U2066 (N_2066,In_983,In_173);
nor U2067 (N_2067,In_2951,In_917);
nor U2068 (N_2068,In_3371,In_786);
xnor U2069 (N_2069,In_3766,In_400);
or U2070 (N_2070,In_2552,In_2635);
nand U2071 (N_2071,In_448,In_4549);
nand U2072 (N_2072,In_3217,In_544);
or U2073 (N_2073,In_2136,In_581);
nor U2074 (N_2074,In_1821,In_912);
nand U2075 (N_2075,In_3088,In_2880);
or U2076 (N_2076,In_3150,In_2385);
or U2077 (N_2077,In_1354,In_4035);
nor U2078 (N_2078,In_1748,In_2268);
nor U2079 (N_2079,In_3907,In_4858);
nor U2080 (N_2080,In_502,In_4917);
nor U2081 (N_2081,In_4950,In_351);
nor U2082 (N_2082,In_1244,In_4304);
nand U2083 (N_2083,In_2841,In_1418);
and U2084 (N_2084,In_737,In_3633);
nor U2085 (N_2085,In_1760,In_643);
and U2086 (N_2086,In_1340,In_331);
and U2087 (N_2087,In_2169,In_1771);
nor U2088 (N_2088,In_4627,In_1057);
and U2089 (N_2089,In_588,In_3322);
or U2090 (N_2090,In_903,In_4198);
nand U2091 (N_2091,In_3385,In_4759);
nand U2092 (N_2092,In_4785,In_2829);
or U2093 (N_2093,In_188,In_4140);
nor U2094 (N_2094,In_1271,In_1805);
xor U2095 (N_2095,In_3422,In_82);
nand U2096 (N_2096,In_2859,In_1632);
xor U2097 (N_2097,In_4067,In_3389);
nand U2098 (N_2098,In_3324,In_4965);
nand U2099 (N_2099,In_2484,In_1772);
nand U2100 (N_2100,In_2164,In_2372);
nor U2101 (N_2101,In_2813,In_1968);
xor U2102 (N_2102,In_628,In_123);
xnor U2103 (N_2103,In_3290,In_2952);
xnor U2104 (N_2104,In_457,In_4753);
and U2105 (N_2105,In_3446,In_4026);
xor U2106 (N_2106,In_748,In_2589);
nor U2107 (N_2107,In_4772,In_4752);
xnor U2108 (N_2108,In_2064,In_2835);
or U2109 (N_2109,In_2344,In_4699);
and U2110 (N_2110,In_1342,In_4846);
xor U2111 (N_2111,In_3308,In_593);
nor U2112 (N_2112,In_3947,In_3955);
nor U2113 (N_2113,In_3271,In_126);
xor U2114 (N_2114,In_1593,In_4110);
and U2115 (N_2115,In_1696,In_4281);
and U2116 (N_2116,In_132,In_848);
xnor U2117 (N_2117,In_3661,In_2028);
or U2118 (N_2118,In_3127,In_2807);
and U2119 (N_2119,In_199,In_2102);
and U2120 (N_2120,In_1679,In_1601);
nand U2121 (N_2121,In_3289,In_4652);
xor U2122 (N_2122,In_1553,In_3887);
and U2123 (N_2123,In_3708,In_906);
and U2124 (N_2124,In_562,In_4127);
or U2125 (N_2125,In_597,In_3835);
nor U2126 (N_2126,In_1616,In_3372);
nand U2127 (N_2127,In_4616,In_2188);
or U2128 (N_2128,In_4696,In_2455);
xor U2129 (N_2129,In_3352,In_3222);
nor U2130 (N_2130,In_1490,In_411);
nand U2131 (N_2131,In_365,In_1538);
and U2132 (N_2132,In_1452,In_2496);
xnor U2133 (N_2133,In_3662,In_2046);
and U2134 (N_2134,In_584,In_1675);
or U2135 (N_2135,In_2486,In_1936);
xnor U2136 (N_2136,In_796,In_2792);
nand U2137 (N_2137,In_3618,In_895);
nand U2138 (N_2138,In_2671,In_4388);
nand U2139 (N_2139,In_828,In_2567);
nor U2140 (N_2140,In_454,In_1178);
nand U2141 (N_2141,In_158,In_4454);
nor U2142 (N_2142,In_1314,In_4143);
nor U2143 (N_2143,In_2948,In_2532);
or U2144 (N_2144,In_1176,In_675);
nor U2145 (N_2145,In_488,In_3902);
nor U2146 (N_2146,In_2934,In_3279);
xnor U2147 (N_2147,In_996,In_4809);
or U2148 (N_2148,In_2326,In_139);
and U2149 (N_2149,In_2526,In_1740);
nor U2150 (N_2150,In_1279,In_2656);
xor U2151 (N_2151,In_3153,In_3715);
and U2152 (N_2152,In_1068,In_4150);
nand U2153 (N_2153,In_3102,In_700);
or U2154 (N_2154,In_997,In_183);
xor U2155 (N_2155,In_3407,In_3494);
nor U2156 (N_2156,In_4859,In_533);
nor U2157 (N_2157,In_68,In_3981);
and U2158 (N_2158,In_1268,In_379);
or U2159 (N_2159,In_1860,In_3215);
and U2160 (N_2160,In_1291,In_2106);
and U2161 (N_2161,In_3669,In_3484);
and U2162 (N_2162,In_1625,In_1435);
nand U2163 (N_2163,In_2525,In_3566);
nor U2164 (N_2164,In_4527,In_4374);
nor U2165 (N_2165,In_10,In_4406);
or U2166 (N_2166,In_2953,In_2352);
nand U2167 (N_2167,In_4669,In_1878);
or U2168 (N_2168,In_3415,In_1028);
nor U2169 (N_2169,In_2039,In_231);
and U2170 (N_2170,In_4487,In_1445);
xor U2171 (N_2171,In_1012,In_1750);
xnor U2172 (N_2172,In_3886,In_4171);
nor U2173 (N_2173,In_3165,In_686);
nor U2174 (N_2174,In_814,In_658);
and U2175 (N_2175,In_83,In_3996);
nand U2176 (N_2176,In_1742,In_344);
or U2177 (N_2177,In_3272,In_1391);
or U2178 (N_2178,In_284,In_2695);
xnor U2179 (N_2179,In_3584,In_2600);
nor U2180 (N_2180,In_3297,In_858);
or U2181 (N_2181,In_4398,In_2474);
or U2182 (N_2182,In_3288,In_627);
and U2183 (N_2183,In_3632,In_4926);
nand U2184 (N_2184,In_4016,In_4754);
nand U2185 (N_2185,In_1237,In_473);
and U2186 (N_2186,In_4864,In_30);
nand U2187 (N_2187,In_225,In_3058);
nand U2188 (N_2188,In_762,In_1649);
or U2189 (N_2189,In_1385,In_2099);
xnor U2190 (N_2190,In_1398,In_2205);
and U2191 (N_2191,In_4942,In_530);
nand U2192 (N_2192,In_2298,In_61);
nor U2193 (N_2193,In_3575,In_1214);
xor U2194 (N_2194,In_442,In_1067);
or U2195 (N_2195,In_4214,In_4672);
xnor U2196 (N_2196,In_1156,In_1433);
nand U2197 (N_2197,In_1422,In_1109);
xor U2198 (N_2198,In_2523,In_2674);
nor U2199 (N_2199,In_892,In_3815);
or U2200 (N_2200,In_913,In_4894);
nor U2201 (N_2201,In_3797,In_3784);
nor U2202 (N_2202,In_3877,In_2772);
nand U2203 (N_2203,In_383,In_922);
nand U2204 (N_2204,In_3478,In_313);
or U2205 (N_2205,In_4358,In_3329);
xor U2206 (N_2206,In_867,In_1902);
xnor U2207 (N_2207,In_633,In_4821);
or U2208 (N_2208,In_1111,In_3462);
or U2209 (N_2209,In_2821,In_152);
or U2210 (N_2210,In_3244,In_4756);
nor U2211 (N_2211,In_1685,In_1680);
or U2212 (N_2212,In_89,In_2383);
nor U2213 (N_2213,In_3075,In_4117);
and U2214 (N_2214,In_2752,In_2846);
and U2215 (N_2215,In_4670,In_1171);
and U2216 (N_2216,In_2990,In_1573);
and U2217 (N_2217,In_3175,In_522);
xnor U2218 (N_2218,In_1099,In_3512);
nor U2219 (N_2219,In_2091,In_3169);
nor U2220 (N_2220,In_2987,In_2658);
and U2221 (N_2221,In_2349,In_4636);
xnor U2222 (N_2222,In_1493,In_2075);
or U2223 (N_2223,In_3601,In_1441);
nor U2224 (N_2224,In_3540,In_2459);
nor U2225 (N_2225,In_355,In_2339);
nor U2226 (N_2226,In_2265,In_2076);
nand U2227 (N_2227,In_4102,In_920);
or U2228 (N_2228,In_886,In_3373);
nand U2229 (N_2229,In_1328,In_2758);
nand U2230 (N_2230,In_1517,In_3796);
or U2231 (N_2231,In_2995,In_1401);
or U2232 (N_2232,In_1525,In_4653);
or U2233 (N_2233,In_3807,In_3059);
and U2234 (N_2234,In_2989,In_940);
or U2235 (N_2235,In_2203,In_1978);
or U2236 (N_2236,In_106,In_1604);
and U2237 (N_2237,In_479,In_4045);
nand U2238 (N_2238,In_2469,In_3988);
and U2239 (N_2239,In_4262,In_2441);
nand U2240 (N_2240,In_670,In_3381);
or U2241 (N_2241,In_3995,In_1866);
nand U2242 (N_2242,In_3644,In_3595);
and U2243 (N_2243,In_3302,In_663);
and U2244 (N_2244,In_4499,In_3179);
nand U2245 (N_2245,In_774,In_2361);
nand U2246 (N_2246,In_20,In_445);
or U2247 (N_2247,In_1558,In_3398);
and U2248 (N_2248,In_352,In_1707);
nand U2249 (N_2249,In_3577,In_3430);
or U2250 (N_2250,In_104,In_94);
or U2251 (N_2251,In_3245,In_4738);
nand U2252 (N_2252,In_4715,In_3545);
or U2253 (N_2253,In_3362,In_4443);
and U2254 (N_2254,In_1023,In_4525);
and U2255 (N_2255,In_4147,In_222);
xor U2256 (N_2256,In_2916,In_2823);
or U2257 (N_2257,In_668,In_4513);
or U2258 (N_2258,In_3987,In_2313);
nand U2259 (N_2259,In_2267,In_3703);
or U2260 (N_2260,In_437,In_401);
nor U2261 (N_2261,In_769,In_1272);
xnor U2262 (N_2262,In_1475,In_3959);
or U2263 (N_2263,In_857,In_1847);
nor U2264 (N_2264,In_644,In_667);
nor U2265 (N_2265,In_3772,In_933);
nor U2266 (N_2266,In_3568,In_3778);
and U2267 (N_2267,In_2115,In_4226);
xor U2268 (N_2268,In_3068,In_701);
or U2269 (N_2269,In_753,In_2919);
nand U2270 (N_2270,In_4554,In_3652);
nand U2271 (N_2271,In_1702,In_1181);
and U2272 (N_2272,In_3960,In_3455);
nand U2273 (N_2273,In_622,In_1837);
and U2274 (N_2274,In_4282,In_4177);
nor U2275 (N_2275,In_2141,In_4667);
xor U2276 (N_2276,In_4467,In_2777);
nand U2277 (N_2277,In_2984,In_1226);
nor U2278 (N_2278,In_2787,In_2331);
and U2279 (N_2279,In_4066,In_624);
or U2280 (N_2280,In_3916,In_3239);
or U2281 (N_2281,In_4879,In_3642);
nor U2282 (N_2282,In_4008,In_589);
nand U2283 (N_2283,In_1168,In_2967);
and U2284 (N_2284,In_1883,In_2623);
and U2285 (N_2285,In_577,In_1961);
nor U2286 (N_2286,In_1562,In_2495);
nand U2287 (N_2287,In_2596,In_270);
or U2288 (N_2288,In_2688,In_4469);
nor U2289 (N_2289,In_34,In_2895);
or U2290 (N_2290,In_4791,In_246);
nor U2291 (N_2291,In_1041,In_1191);
nor U2292 (N_2292,In_1047,In_4535);
or U2293 (N_2293,In_2720,In_2810);
or U2294 (N_2294,In_42,In_2745);
and U2295 (N_2295,In_55,In_1096);
nor U2296 (N_2296,In_2587,In_4410);
nand U2297 (N_2297,In_4400,In_3173);
and U2298 (N_2298,In_366,In_165);
or U2299 (N_2299,In_1870,In_267);
and U2300 (N_2300,In_1882,In_812);
and U2301 (N_2301,In_3515,In_4780);
nor U2302 (N_2302,In_272,In_506);
nor U2303 (N_2303,In_1417,In_24);
xor U2304 (N_2304,In_1294,In_1080);
nor U2305 (N_2305,In_3810,In_4192);
xor U2306 (N_2306,In_919,In_3859);
or U2307 (N_2307,In_2108,In_2740);
and U2308 (N_2308,In_4402,In_4416);
nand U2309 (N_2309,In_1721,In_4197);
nor U2310 (N_2310,In_4151,In_3538);
or U2311 (N_2311,In_447,In_2680);
nand U2312 (N_2312,In_4082,In_1810);
or U2313 (N_2313,In_3647,In_3738);
nor U2314 (N_2314,In_2651,In_141);
or U2315 (N_2315,In_557,In_1578);
xnor U2316 (N_2316,In_3071,In_3583);
nand U2317 (N_2317,In_1463,In_2960);
nor U2318 (N_2318,In_4157,In_4096);
or U2319 (N_2319,In_1267,In_1035);
or U2320 (N_2320,In_596,In_3951);
nand U2321 (N_2321,In_1767,In_527);
or U2322 (N_2322,In_2285,In_718);
xor U2323 (N_2323,In_2040,In_1752);
nand U2324 (N_2324,In_2928,In_3806);
nor U2325 (N_2325,In_75,In_612);
nor U2326 (N_2326,In_2742,In_3186);
nor U2327 (N_2327,In_881,In_2346);
or U2328 (N_2328,In_2302,In_4898);
and U2329 (N_2329,In_1146,In_4975);
nor U2330 (N_2330,In_3015,In_2266);
nor U2331 (N_2331,In_2036,In_2081);
and U2332 (N_2332,In_1346,In_110);
nand U2333 (N_2333,In_3171,In_3906);
and U2334 (N_2334,In_1440,In_3822);
or U2335 (N_2335,In_498,In_918);
nand U2336 (N_2336,In_2700,In_369);
nand U2337 (N_2337,In_1086,In_2444);
nor U2338 (N_2338,In_510,In_3639);
nand U2339 (N_2339,In_287,In_330);
xnor U2340 (N_2340,In_1462,In_2689);
nand U2341 (N_2341,In_4836,In_1484);
nor U2342 (N_2342,In_2065,In_2096);
or U2343 (N_2343,In_1549,In_1718);
nand U2344 (N_2344,In_1206,In_3233);
and U2345 (N_2345,In_2834,In_2112);
nand U2346 (N_2346,In_3693,In_2626);
and U2347 (N_2347,In_4444,In_4436);
xor U2348 (N_2348,In_1977,In_3845);
nor U2349 (N_2349,In_782,In_261);
nor U2350 (N_2350,In_3552,In_35);
nand U2351 (N_2351,In_1239,In_4097);
and U2352 (N_2352,In_4938,In_1276);
nand U2353 (N_2353,In_4774,In_4714);
or U2354 (N_2354,In_3657,In_4863);
or U2355 (N_2355,In_3038,In_2452);
and U2356 (N_2356,In_3358,In_257);
or U2357 (N_2357,In_2219,In_761);
or U2358 (N_2358,In_1313,In_78);
or U2359 (N_2359,In_1000,In_1471);
xnor U2360 (N_2360,In_4324,In_31);
nor U2361 (N_2361,In_2481,In_2419);
and U2362 (N_2362,In_166,In_4764);
or U2363 (N_2363,In_2399,In_3573);
and U2364 (N_2364,In_778,In_850);
nand U2365 (N_2365,In_1459,In_3182);
nor U2366 (N_2366,In_2148,In_1722);
and U2367 (N_2367,In_2744,In_375);
xor U2368 (N_2368,In_1204,In_409);
nand U2369 (N_2369,In_4662,In_1952);
nor U2370 (N_2370,In_2718,In_4648);
or U2371 (N_2371,In_2453,In_3733);
and U2372 (N_2372,In_2664,In_1913);
and U2373 (N_2373,In_4519,In_3090);
and U2374 (N_2374,In_705,In_914);
nor U2375 (N_2375,In_3888,In_1846);
nor U2376 (N_2376,In_2822,In_4713);
nand U2377 (N_2377,In_1379,In_4712);
or U2378 (N_2378,In_3525,In_3474);
nand U2379 (N_2379,In_1637,In_1914);
or U2380 (N_2380,In_2727,In_4930);
nand U2381 (N_2381,In_2708,In_2343);
nor U2382 (N_2382,In_4848,In_3751);
or U2383 (N_2383,In_1467,In_2318);
nor U2384 (N_2384,In_1180,In_4373);
nand U2385 (N_2385,In_4376,In_2817);
and U2386 (N_2386,In_4557,In_3157);
nand U2387 (N_2387,In_3321,In_2107);
nand U2388 (N_2388,In_4335,In_798);
nand U2389 (N_2389,In_2024,In_3120);
or U2390 (N_2390,In_1486,In_2271);
nor U2391 (N_2391,In_3593,In_2);
nor U2392 (N_2392,In_3131,In_3743);
and U2393 (N_2393,In_4344,In_1606);
or U2394 (N_2394,In_255,In_3063);
nor U2395 (N_2395,In_3216,In_459);
and U2396 (N_2396,In_4083,In_228);
and U2397 (N_2397,In_2309,In_3413);
and U2398 (N_2398,In_208,In_4503);
nor U2399 (N_2399,In_3558,In_863);
nand U2400 (N_2400,In_2144,In_3816);
nor U2401 (N_2401,In_1948,In_1330);
nand U2402 (N_2402,In_3826,In_185);
and U2403 (N_2403,In_4508,In_3294);
and U2404 (N_2404,In_2506,In_4765);
nand U2405 (N_2405,In_1108,In_1985);
nand U2406 (N_2406,In_1795,In_3831);
xnor U2407 (N_2407,In_735,In_4912);
nor U2408 (N_2408,In_2195,In_2030);
or U2409 (N_2409,In_2790,In_2172);
xnor U2410 (N_2410,In_3936,In_3780);
or U2411 (N_2411,In_1542,In_76);
nor U2412 (N_2412,In_3728,In_3508);
nor U2413 (N_2413,In_2972,In_1780);
nand U2414 (N_2414,In_1858,In_4497);
nor U2415 (N_2415,In_1873,In_629);
or U2416 (N_2416,In_214,In_3841);
and U2417 (N_2417,In_1682,In_438);
and U2418 (N_2418,In_2692,In_3168);
or U2419 (N_2419,In_1321,In_2749);
nor U2420 (N_2420,In_2798,In_4515);
and U2421 (N_2421,In_4704,In_3055);
nand U2422 (N_2422,In_170,In_2299);
nor U2423 (N_2423,In_3444,In_3658);
and U2424 (N_2424,In_220,In_4970);
and U2425 (N_2425,In_785,In_3339);
nand U2426 (N_2426,In_4125,In_3468);
nor U2427 (N_2427,In_3351,In_1362);
or U2428 (N_2428,In_1102,In_2761);
or U2429 (N_2429,In_4065,In_4645);
and U2430 (N_2430,In_4383,In_3827);
nor U2431 (N_2431,In_2831,In_3042);
nor U2432 (N_2432,In_2648,In_2052);
nand U2433 (N_2433,In_134,In_3284);
or U2434 (N_2434,In_3234,In_1069);
or U2435 (N_2435,In_1234,In_2836);
nor U2436 (N_2436,In_3927,In_4288);
nand U2437 (N_2437,In_882,In_2884);
nand U2438 (N_2438,In_975,In_3864);
nor U2439 (N_2439,In_1865,In_1071);
nand U2440 (N_2440,In_2197,In_3655);
nor U2441 (N_2441,In_901,In_1861);
or U2442 (N_2442,In_2152,In_3453);
nor U2443 (N_2443,In_3694,In_716);
or U2444 (N_2444,In_4407,In_2165);
xnor U2445 (N_2445,In_354,In_3057);
or U2446 (N_2446,In_4440,In_2487);
xnor U2447 (N_2447,In_1323,In_3683);
nor U2448 (N_2448,In_1792,In_509);
nor U2449 (N_2449,In_2492,In_250);
and U2450 (N_2450,In_4284,In_2612);
and U2451 (N_2451,In_2191,In_4985);
and U2452 (N_2452,In_2137,In_2746);
or U2453 (N_2453,In_160,In_482);
or U2454 (N_2454,In_1745,In_558);
or U2455 (N_2455,In_3745,In_4254);
nand U2456 (N_2456,In_3861,In_2657);
nor U2457 (N_2457,In_1895,In_3612);
and U2458 (N_2458,In_259,In_2437);
nor U2459 (N_2459,In_1783,In_4882);
nand U2460 (N_2460,In_792,In_4633);
nor U2461 (N_2461,In_4345,In_472);
or U2462 (N_2462,In_2696,In_902);
nor U2463 (N_2463,In_2170,In_4694);
and U2464 (N_2464,In_4718,In_1912);
nor U2465 (N_2465,In_1897,In_548);
nor U2466 (N_2466,In_3273,In_1911);
nor U2467 (N_2467,In_1196,In_2540);
and U2468 (N_2468,In_4490,In_1045);
nand U2469 (N_2469,In_23,In_2634);
and U2470 (N_2470,In_1411,In_2117);
xnor U2471 (N_2471,In_2653,In_561);
and U2472 (N_2472,In_4466,In_2874);
or U2473 (N_2473,In_4451,In_338);
and U2474 (N_2474,In_889,In_4449);
nand U2475 (N_2475,In_631,In_2217);
and U2476 (N_2476,In_2010,In_3997);
nand U2477 (N_2477,In_1708,In_264);
or U2478 (N_2478,In_2095,In_1118);
and U2479 (N_2479,In_676,In_1476);
nor U2480 (N_2480,In_496,In_2562);
or U2481 (N_2481,In_150,In_1349);
and U2482 (N_2482,In_2243,In_1969);
nand U2483 (N_2483,In_3050,In_765);
nand U2484 (N_2484,In_4506,In_4294);
nor U2485 (N_2485,In_3206,In_1535);
and U2486 (N_2486,In_1170,In_2025);
nor U2487 (N_2487,In_2690,In_560);
xnor U2488 (N_2488,In_1670,In_3712);
nor U2489 (N_2489,In_4488,In_4246);
xor U2490 (N_2490,In_4160,In_4153);
nor U2491 (N_2491,In_3752,In_2356);
nand U2492 (N_2492,In_3910,In_2669);
nor U2493 (N_2493,In_1207,In_4355);
and U2494 (N_2494,In_1390,In_1540);
xor U2495 (N_2495,In_2687,In_4166);
nand U2496 (N_2496,In_4732,In_2620);
xnor U2497 (N_2497,In_4564,In_4095);
or U2498 (N_2498,In_1716,In_3126);
or U2499 (N_2499,In_52,In_2906);
nand U2500 (N_2500,In_1241,In_2648);
xnor U2501 (N_2501,In_1045,In_2384);
nand U2502 (N_2502,In_92,In_356);
nand U2503 (N_2503,In_1747,In_1115);
and U2504 (N_2504,In_2315,In_2015);
or U2505 (N_2505,In_479,In_3646);
or U2506 (N_2506,In_3028,In_4130);
and U2507 (N_2507,In_869,In_595);
and U2508 (N_2508,In_4296,In_3057);
and U2509 (N_2509,In_4221,In_1011);
or U2510 (N_2510,In_209,In_1855);
nor U2511 (N_2511,In_2374,In_2464);
nor U2512 (N_2512,In_235,In_176);
xnor U2513 (N_2513,In_2088,In_4661);
and U2514 (N_2514,In_2398,In_1057);
nor U2515 (N_2515,In_1425,In_2357);
nand U2516 (N_2516,In_1765,In_180);
or U2517 (N_2517,In_32,In_4272);
and U2518 (N_2518,In_751,In_3115);
nor U2519 (N_2519,In_1772,In_1727);
or U2520 (N_2520,In_2301,In_4421);
and U2521 (N_2521,In_4185,In_3842);
and U2522 (N_2522,In_4291,In_4379);
nand U2523 (N_2523,In_4553,In_74);
and U2524 (N_2524,In_4314,In_4567);
nand U2525 (N_2525,In_4264,In_4706);
or U2526 (N_2526,In_3622,In_4075);
nand U2527 (N_2527,In_2210,In_1882);
nor U2528 (N_2528,In_4816,In_3303);
or U2529 (N_2529,In_1020,In_2403);
or U2530 (N_2530,In_3011,In_3604);
nor U2531 (N_2531,In_4187,In_3579);
and U2532 (N_2532,In_1032,In_275);
xnor U2533 (N_2533,In_1615,In_3956);
nand U2534 (N_2534,In_2063,In_2016);
or U2535 (N_2535,In_2927,In_1370);
nor U2536 (N_2536,In_3905,In_1056);
nor U2537 (N_2537,In_3508,In_4338);
nand U2538 (N_2538,In_4609,In_1772);
or U2539 (N_2539,In_667,In_4504);
and U2540 (N_2540,In_1309,In_1946);
xnor U2541 (N_2541,In_1090,In_3984);
or U2542 (N_2542,In_4352,In_846);
nor U2543 (N_2543,In_3723,In_4438);
nand U2544 (N_2544,In_1162,In_4630);
and U2545 (N_2545,In_4921,In_2977);
xnor U2546 (N_2546,In_2863,In_4609);
and U2547 (N_2547,In_2588,In_1793);
or U2548 (N_2548,In_3337,In_762);
nand U2549 (N_2549,In_631,In_3762);
nand U2550 (N_2550,In_3317,In_1617);
nand U2551 (N_2551,In_996,In_4865);
nand U2552 (N_2552,In_4913,In_4439);
or U2553 (N_2553,In_2682,In_2927);
nor U2554 (N_2554,In_2049,In_1767);
or U2555 (N_2555,In_3386,In_3843);
nand U2556 (N_2556,In_783,In_1264);
and U2557 (N_2557,In_3496,In_878);
nand U2558 (N_2558,In_3277,In_868);
or U2559 (N_2559,In_1179,In_2071);
nor U2560 (N_2560,In_4148,In_4140);
or U2561 (N_2561,In_4638,In_1029);
and U2562 (N_2562,In_3574,In_2247);
or U2563 (N_2563,In_1069,In_2169);
and U2564 (N_2564,In_3756,In_489);
nor U2565 (N_2565,In_1568,In_178);
or U2566 (N_2566,In_1810,In_897);
nor U2567 (N_2567,In_104,In_513);
nor U2568 (N_2568,In_4452,In_2996);
and U2569 (N_2569,In_596,In_1834);
nor U2570 (N_2570,In_4262,In_2398);
nor U2571 (N_2571,In_1256,In_2874);
nor U2572 (N_2572,In_2448,In_73);
nand U2573 (N_2573,In_2954,In_4142);
or U2574 (N_2574,In_167,In_4879);
nor U2575 (N_2575,In_4673,In_3503);
nand U2576 (N_2576,In_4854,In_4024);
nor U2577 (N_2577,In_993,In_3340);
or U2578 (N_2578,In_4009,In_4569);
and U2579 (N_2579,In_2491,In_1784);
nand U2580 (N_2580,In_3091,In_119);
and U2581 (N_2581,In_3172,In_2900);
xnor U2582 (N_2582,In_2044,In_228);
nand U2583 (N_2583,In_3751,In_1844);
and U2584 (N_2584,In_740,In_3955);
nand U2585 (N_2585,In_4895,In_1737);
and U2586 (N_2586,In_2125,In_2649);
and U2587 (N_2587,In_410,In_842);
or U2588 (N_2588,In_2250,In_3599);
or U2589 (N_2589,In_4357,In_3172);
and U2590 (N_2590,In_3936,In_3442);
nor U2591 (N_2591,In_3805,In_2690);
nand U2592 (N_2592,In_1019,In_1918);
nand U2593 (N_2593,In_322,In_631);
or U2594 (N_2594,In_4406,In_3849);
or U2595 (N_2595,In_3701,In_3036);
and U2596 (N_2596,In_2048,In_665);
nand U2597 (N_2597,In_4192,In_757);
nand U2598 (N_2598,In_4084,In_4102);
xnor U2599 (N_2599,In_1819,In_1624);
nor U2600 (N_2600,In_2980,In_1025);
and U2601 (N_2601,In_1853,In_4123);
nor U2602 (N_2602,In_3719,In_928);
nor U2603 (N_2603,In_768,In_4117);
nor U2604 (N_2604,In_1361,In_3811);
or U2605 (N_2605,In_2081,In_900);
nor U2606 (N_2606,In_2514,In_4068);
or U2607 (N_2607,In_3379,In_1515);
or U2608 (N_2608,In_18,In_4673);
or U2609 (N_2609,In_918,In_1516);
nor U2610 (N_2610,In_2982,In_4649);
nor U2611 (N_2611,In_1844,In_1106);
xnor U2612 (N_2612,In_1432,In_3058);
and U2613 (N_2613,In_17,In_1952);
or U2614 (N_2614,In_2176,In_626);
xnor U2615 (N_2615,In_1056,In_779);
nand U2616 (N_2616,In_1537,In_1615);
and U2617 (N_2617,In_1812,In_350);
nand U2618 (N_2618,In_53,In_4010);
or U2619 (N_2619,In_1948,In_946);
and U2620 (N_2620,In_3486,In_1398);
nor U2621 (N_2621,In_208,In_1082);
or U2622 (N_2622,In_3175,In_1669);
and U2623 (N_2623,In_3896,In_1187);
xor U2624 (N_2624,In_4826,In_506);
nor U2625 (N_2625,In_550,In_4909);
or U2626 (N_2626,In_4077,In_1804);
and U2627 (N_2627,In_1069,In_4750);
or U2628 (N_2628,In_3141,In_3885);
nor U2629 (N_2629,In_3870,In_4743);
nand U2630 (N_2630,In_3848,In_2780);
nor U2631 (N_2631,In_2924,In_133);
nand U2632 (N_2632,In_1594,In_1180);
or U2633 (N_2633,In_1786,In_4370);
and U2634 (N_2634,In_26,In_170);
nand U2635 (N_2635,In_3795,In_2564);
nor U2636 (N_2636,In_4451,In_860);
xnor U2637 (N_2637,In_2820,In_2278);
and U2638 (N_2638,In_1226,In_1675);
or U2639 (N_2639,In_1770,In_1527);
or U2640 (N_2640,In_3526,In_717);
or U2641 (N_2641,In_999,In_4634);
xor U2642 (N_2642,In_1920,In_3008);
xor U2643 (N_2643,In_519,In_4356);
nand U2644 (N_2644,In_3321,In_2482);
nor U2645 (N_2645,In_3845,In_4129);
nand U2646 (N_2646,In_1067,In_4466);
nand U2647 (N_2647,In_643,In_4565);
and U2648 (N_2648,In_4677,In_256);
nor U2649 (N_2649,In_23,In_3654);
or U2650 (N_2650,In_1000,In_1659);
nor U2651 (N_2651,In_2938,In_460);
and U2652 (N_2652,In_486,In_1875);
nor U2653 (N_2653,In_650,In_4149);
nand U2654 (N_2654,In_3426,In_1041);
nor U2655 (N_2655,In_1890,In_4889);
nand U2656 (N_2656,In_1607,In_3689);
or U2657 (N_2657,In_3939,In_1840);
or U2658 (N_2658,In_927,In_2338);
xnor U2659 (N_2659,In_1755,In_3514);
and U2660 (N_2660,In_3966,In_4722);
xor U2661 (N_2661,In_593,In_3915);
and U2662 (N_2662,In_3533,In_4882);
nand U2663 (N_2663,In_971,In_1848);
nor U2664 (N_2664,In_2545,In_2946);
and U2665 (N_2665,In_658,In_2953);
nand U2666 (N_2666,In_19,In_4760);
or U2667 (N_2667,In_3092,In_4533);
nand U2668 (N_2668,In_4559,In_60);
nor U2669 (N_2669,In_2231,In_1383);
nand U2670 (N_2670,In_867,In_834);
or U2671 (N_2671,In_947,In_2967);
nor U2672 (N_2672,In_3106,In_2196);
and U2673 (N_2673,In_2834,In_582);
or U2674 (N_2674,In_866,In_4497);
and U2675 (N_2675,In_3496,In_1201);
nand U2676 (N_2676,In_622,In_4694);
or U2677 (N_2677,In_2522,In_741);
xnor U2678 (N_2678,In_3745,In_1920);
nor U2679 (N_2679,In_2685,In_126);
nand U2680 (N_2680,In_3811,In_4737);
nor U2681 (N_2681,In_4867,In_4139);
nor U2682 (N_2682,In_1913,In_3055);
nor U2683 (N_2683,In_1488,In_4022);
or U2684 (N_2684,In_757,In_1531);
nand U2685 (N_2685,In_390,In_3412);
and U2686 (N_2686,In_1617,In_4712);
nand U2687 (N_2687,In_282,In_4225);
or U2688 (N_2688,In_2262,In_1975);
and U2689 (N_2689,In_999,In_1544);
and U2690 (N_2690,In_3252,In_4547);
and U2691 (N_2691,In_1500,In_1009);
nor U2692 (N_2692,In_1740,In_4098);
and U2693 (N_2693,In_1979,In_1912);
nor U2694 (N_2694,In_4970,In_4579);
or U2695 (N_2695,In_362,In_1778);
and U2696 (N_2696,In_550,In_4522);
or U2697 (N_2697,In_1660,In_4538);
and U2698 (N_2698,In_3188,In_2967);
nand U2699 (N_2699,In_3711,In_588);
nand U2700 (N_2700,In_3209,In_4413);
nand U2701 (N_2701,In_2167,In_4731);
nand U2702 (N_2702,In_2100,In_1394);
or U2703 (N_2703,In_1938,In_4711);
nor U2704 (N_2704,In_4290,In_496);
nor U2705 (N_2705,In_4234,In_4053);
nor U2706 (N_2706,In_4253,In_3645);
or U2707 (N_2707,In_3420,In_2240);
nor U2708 (N_2708,In_4957,In_2427);
nor U2709 (N_2709,In_1027,In_3604);
and U2710 (N_2710,In_1,In_2696);
or U2711 (N_2711,In_4052,In_1333);
or U2712 (N_2712,In_1577,In_2149);
nand U2713 (N_2713,In_4892,In_2809);
or U2714 (N_2714,In_210,In_909);
and U2715 (N_2715,In_1314,In_2188);
nor U2716 (N_2716,In_354,In_2971);
nand U2717 (N_2717,In_387,In_1979);
and U2718 (N_2718,In_227,In_212);
nor U2719 (N_2719,In_3839,In_4038);
or U2720 (N_2720,In_2444,In_4353);
xor U2721 (N_2721,In_3168,In_142);
nand U2722 (N_2722,In_1854,In_3783);
and U2723 (N_2723,In_4433,In_3332);
or U2724 (N_2724,In_1993,In_93);
and U2725 (N_2725,In_3833,In_4758);
and U2726 (N_2726,In_892,In_1902);
nand U2727 (N_2727,In_2967,In_4683);
nand U2728 (N_2728,In_4801,In_3312);
nor U2729 (N_2729,In_401,In_3479);
and U2730 (N_2730,In_3994,In_2567);
nand U2731 (N_2731,In_4232,In_3310);
and U2732 (N_2732,In_922,In_2983);
and U2733 (N_2733,In_860,In_1212);
nand U2734 (N_2734,In_924,In_1892);
xnor U2735 (N_2735,In_3876,In_1091);
nor U2736 (N_2736,In_96,In_723);
nor U2737 (N_2737,In_2378,In_4037);
xor U2738 (N_2738,In_3640,In_3693);
nand U2739 (N_2739,In_880,In_2562);
or U2740 (N_2740,In_1606,In_2301);
xnor U2741 (N_2741,In_969,In_4402);
or U2742 (N_2742,In_1739,In_476);
nor U2743 (N_2743,In_4635,In_442);
and U2744 (N_2744,In_3431,In_3571);
nor U2745 (N_2745,In_1581,In_4122);
nand U2746 (N_2746,In_4100,In_4690);
and U2747 (N_2747,In_3342,In_2721);
xnor U2748 (N_2748,In_2878,In_3125);
nor U2749 (N_2749,In_3978,In_3611);
nand U2750 (N_2750,In_754,In_4619);
or U2751 (N_2751,In_788,In_3446);
nor U2752 (N_2752,In_3769,In_1174);
xor U2753 (N_2753,In_957,In_500);
nor U2754 (N_2754,In_909,In_2551);
nor U2755 (N_2755,In_3685,In_1475);
xor U2756 (N_2756,In_4060,In_1617);
and U2757 (N_2757,In_64,In_1491);
and U2758 (N_2758,In_4392,In_280);
xor U2759 (N_2759,In_1076,In_4106);
nand U2760 (N_2760,In_2971,In_2079);
and U2761 (N_2761,In_2762,In_2170);
xor U2762 (N_2762,In_1111,In_4535);
or U2763 (N_2763,In_652,In_3278);
nor U2764 (N_2764,In_3176,In_1228);
or U2765 (N_2765,In_1888,In_2624);
nor U2766 (N_2766,In_4072,In_1458);
and U2767 (N_2767,In_1952,In_2379);
and U2768 (N_2768,In_2134,In_4859);
nand U2769 (N_2769,In_3359,In_2104);
and U2770 (N_2770,In_831,In_637);
nand U2771 (N_2771,In_4363,In_4187);
xor U2772 (N_2772,In_2683,In_2691);
and U2773 (N_2773,In_3328,In_898);
or U2774 (N_2774,In_3794,In_2694);
nand U2775 (N_2775,In_1848,In_1215);
xor U2776 (N_2776,In_4554,In_3995);
nand U2777 (N_2777,In_1321,In_35);
nand U2778 (N_2778,In_3735,In_3398);
nor U2779 (N_2779,In_3092,In_1928);
nand U2780 (N_2780,In_2107,In_1458);
nor U2781 (N_2781,In_4957,In_2829);
nand U2782 (N_2782,In_156,In_556);
nand U2783 (N_2783,In_4902,In_2035);
nand U2784 (N_2784,In_1936,In_105);
and U2785 (N_2785,In_3458,In_1904);
nor U2786 (N_2786,In_4575,In_2674);
or U2787 (N_2787,In_64,In_3213);
nor U2788 (N_2788,In_4559,In_3765);
or U2789 (N_2789,In_3711,In_3282);
and U2790 (N_2790,In_1320,In_4244);
and U2791 (N_2791,In_2434,In_881);
nor U2792 (N_2792,In_4675,In_3627);
xnor U2793 (N_2793,In_1245,In_1328);
nand U2794 (N_2794,In_3132,In_780);
or U2795 (N_2795,In_1401,In_4461);
xnor U2796 (N_2796,In_4216,In_4246);
and U2797 (N_2797,In_1143,In_407);
or U2798 (N_2798,In_4251,In_3447);
or U2799 (N_2799,In_4693,In_2916);
xor U2800 (N_2800,In_2353,In_1044);
and U2801 (N_2801,In_1986,In_1458);
or U2802 (N_2802,In_2670,In_4675);
or U2803 (N_2803,In_3403,In_4499);
and U2804 (N_2804,In_2228,In_3442);
and U2805 (N_2805,In_1525,In_4730);
and U2806 (N_2806,In_2995,In_2833);
xor U2807 (N_2807,In_4567,In_4537);
nand U2808 (N_2808,In_3858,In_4179);
nand U2809 (N_2809,In_2004,In_793);
or U2810 (N_2810,In_3262,In_162);
nand U2811 (N_2811,In_362,In_3936);
nor U2812 (N_2812,In_12,In_2127);
nor U2813 (N_2813,In_345,In_430);
or U2814 (N_2814,In_687,In_204);
or U2815 (N_2815,In_4359,In_904);
or U2816 (N_2816,In_2960,In_661);
xor U2817 (N_2817,In_1347,In_2041);
or U2818 (N_2818,In_2100,In_834);
and U2819 (N_2819,In_4926,In_4363);
and U2820 (N_2820,In_484,In_4764);
or U2821 (N_2821,In_938,In_125);
or U2822 (N_2822,In_2552,In_2912);
nand U2823 (N_2823,In_3572,In_4182);
nand U2824 (N_2824,In_4103,In_59);
xnor U2825 (N_2825,In_3139,In_488);
nand U2826 (N_2826,In_2506,In_1219);
nand U2827 (N_2827,In_271,In_1361);
xor U2828 (N_2828,In_4404,In_4523);
and U2829 (N_2829,In_2845,In_685);
nand U2830 (N_2830,In_3493,In_2983);
nor U2831 (N_2831,In_4280,In_1774);
and U2832 (N_2832,In_1758,In_2065);
xor U2833 (N_2833,In_1711,In_709);
nand U2834 (N_2834,In_4586,In_2162);
xnor U2835 (N_2835,In_4271,In_1769);
or U2836 (N_2836,In_1340,In_1546);
nor U2837 (N_2837,In_964,In_3001);
nand U2838 (N_2838,In_4320,In_3818);
or U2839 (N_2839,In_4974,In_1175);
or U2840 (N_2840,In_3103,In_4149);
and U2841 (N_2841,In_2410,In_360);
nand U2842 (N_2842,In_4076,In_2155);
and U2843 (N_2843,In_4132,In_4468);
nor U2844 (N_2844,In_887,In_203);
nor U2845 (N_2845,In_1219,In_1266);
and U2846 (N_2846,In_1395,In_4860);
and U2847 (N_2847,In_4524,In_551);
nor U2848 (N_2848,In_4271,In_3085);
nor U2849 (N_2849,In_1239,In_1169);
nor U2850 (N_2850,In_4234,In_2426);
nand U2851 (N_2851,In_881,In_237);
xor U2852 (N_2852,In_1581,In_2231);
nand U2853 (N_2853,In_2146,In_2640);
or U2854 (N_2854,In_940,In_3997);
nand U2855 (N_2855,In_4691,In_396);
or U2856 (N_2856,In_3302,In_3491);
or U2857 (N_2857,In_3799,In_1355);
and U2858 (N_2858,In_2874,In_1047);
xor U2859 (N_2859,In_2808,In_1280);
nand U2860 (N_2860,In_773,In_4742);
and U2861 (N_2861,In_4675,In_3562);
or U2862 (N_2862,In_3971,In_1373);
or U2863 (N_2863,In_3582,In_4933);
and U2864 (N_2864,In_4332,In_1252);
nor U2865 (N_2865,In_2993,In_1070);
nor U2866 (N_2866,In_716,In_4270);
and U2867 (N_2867,In_4446,In_2864);
and U2868 (N_2868,In_1331,In_2276);
or U2869 (N_2869,In_4539,In_3984);
or U2870 (N_2870,In_4824,In_745);
nand U2871 (N_2871,In_1282,In_1129);
or U2872 (N_2872,In_3249,In_2254);
or U2873 (N_2873,In_497,In_2736);
or U2874 (N_2874,In_4846,In_1232);
nand U2875 (N_2875,In_2032,In_702);
nor U2876 (N_2876,In_140,In_4025);
nor U2877 (N_2877,In_3819,In_3937);
and U2878 (N_2878,In_616,In_1807);
nand U2879 (N_2879,In_1604,In_498);
and U2880 (N_2880,In_4294,In_2049);
nor U2881 (N_2881,In_4350,In_1849);
nand U2882 (N_2882,In_1636,In_3773);
nand U2883 (N_2883,In_1937,In_1433);
nor U2884 (N_2884,In_2823,In_1862);
nand U2885 (N_2885,In_3661,In_1492);
nand U2886 (N_2886,In_3223,In_3159);
or U2887 (N_2887,In_2716,In_3198);
xnor U2888 (N_2888,In_3831,In_3775);
nor U2889 (N_2889,In_1157,In_2307);
nor U2890 (N_2890,In_1947,In_2847);
nand U2891 (N_2891,In_3006,In_3339);
nor U2892 (N_2892,In_2114,In_4295);
or U2893 (N_2893,In_2661,In_3851);
nand U2894 (N_2894,In_2821,In_1034);
nand U2895 (N_2895,In_66,In_2561);
or U2896 (N_2896,In_1372,In_3693);
nand U2897 (N_2897,In_3887,In_1989);
nor U2898 (N_2898,In_1190,In_1099);
and U2899 (N_2899,In_4524,In_4158);
or U2900 (N_2900,In_4152,In_4050);
xnor U2901 (N_2901,In_1591,In_167);
xnor U2902 (N_2902,In_4755,In_2661);
xor U2903 (N_2903,In_2369,In_1307);
and U2904 (N_2904,In_1940,In_741);
and U2905 (N_2905,In_559,In_3502);
and U2906 (N_2906,In_1240,In_2665);
and U2907 (N_2907,In_1936,In_4663);
or U2908 (N_2908,In_2678,In_4379);
and U2909 (N_2909,In_3023,In_2599);
nand U2910 (N_2910,In_4098,In_603);
nand U2911 (N_2911,In_3687,In_3315);
nor U2912 (N_2912,In_950,In_1806);
nand U2913 (N_2913,In_2103,In_3735);
and U2914 (N_2914,In_1188,In_703);
nand U2915 (N_2915,In_1201,In_2401);
nand U2916 (N_2916,In_893,In_4458);
nand U2917 (N_2917,In_1925,In_3237);
and U2918 (N_2918,In_4046,In_4108);
nor U2919 (N_2919,In_4265,In_1198);
and U2920 (N_2920,In_1159,In_2863);
and U2921 (N_2921,In_636,In_158);
nor U2922 (N_2922,In_2462,In_1485);
nor U2923 (N_2923,In_1265,In_211);
nor U2924 (N_2924,In_800,In_542);
or U2925 (N_2925,In_710,In_1553);
or U2926 (N_2926,In_3748,In_925);
nor U2927 (N_2927,In_3928,In_2914);
nand U2928 (N_2928,In_3342,In_4114);
nand U2929 (N_2929,In_795,In_3505);
or U2930 (N_2930,In_930,In_436);
and U2931 (N_2931,In_1092,In_3632);
nand U2932 (N_2932,In_499,In_237);
nand U2933 (N_2933,In_4721,In_4586);
and U2934 (N_2934,In_2631,In_4419);
and U2935 (N_2935,In_4084,In_2251);
nand U2936 (N_2936,In_2506,In_367);
xnor U2937 (N_2937,In_2345,In_3781);
and U2938 (N_2938,In_592,In_3427);
nor U2939 (N_2939,In_1154,In_309);
nor U2940 (N_2940,In_1943,In_969);
and U2941 (N_2941,In_2086,In_4832);
and U2942 (N_2942,In_1104,In_1512);
nand U2943 (N_2943,In_3652,In_267);
or U2944 (N_2944,In_3708,In_1731);
nor U2945 (N_2945,In_445,In_1889);
nor U2946 (N_2946,In_1009,In_1578);
nor U2947 (N_2947,In_448,In_4671);
nor U2948 (N_2948,In_3689,In_4560);
nand U2949 (N_2949,In_438,In_1177);
and U2950 (N_2950,In_3750,In_587);
and U2951 (N_2951,In_3281,In_2173);
nand U2952 (N_2952,In_3692,In_494);
and U2953 (N_2953,In_799,In_3150);
and U2954 (N_2954,In_1423,In_4161);
nand U2955 (N_2955,In_2764,In_3489);
or U2956 (N_2956,In_102,In_3733);
nand U2957 (N_2957,In_1663,In_2273);
or U2958 (N_2958,In_4292,In_1664);
nand U2959 (N_2959,In_120,In_4138);
and U2960 (N_2960,In_354,In_2470);
nand U2961 (N_2961,In_3733,In_4764);
nand U2962 (N_2962,In_2825,In_3164);
or U2963 (N_2963,In_1264,In_934);
nand U2964 (N_2964,In_4728,In_3055);
nand U2965 (N_2965,In_857,In_2588);
nor U2966 (N_2966,In_1311,In_4950);
nand U2967 (N_2967,In_3690,In_4985);
nand U2968 (N_2968,In_2159,In_3581);
and U2969 (N_2969,In_1151,In_3680);
and U2970 (N_2970,In_2389,In_1704);
nor U2971 (N_2971,In_3575,In_3673);
nor U2972 (N_2972,In_4564,In_2153);
or U2973 (N_2973,In_989,In_682);
or U2974 (N_2974,In_565,In_4086);
xor U2975 (N_2975,In_2474,In_4989);
nor U2976 (N_2976,In_4340,In_1467);
and U2977 (N_2977,In_2133,In_2677);
or U2978 (N_2978,In_2135,In_2700);
nand U2979 (N_2979,In_2701,In_3479);
nand U2980 (N_2980,In_2117,In_2594);
and U2981 (N_2981,In_1382,In_2775);
nand U2982 (N_2982,In_46,In_1149);
nand U2983 (N_2983,In_115,In_4237);
and U2984 (N_2984,In_3241,In_2840);
xor U2985 (N_2985,In_4195,In_212);
or U2986 (N_2986,In_3040,In_4157);
nand U2987 (N_2987,In_866,In_2563);
nand U2988 (N_2988,In_2798,In_426);
xor U2989 (N_2989,In_621,In_2112);
nor U2990 (N_2990,In_805,In_2070);
nor U2991 (N_2991,In_3176,In_2951);
nand U2992 (N_2992,In_1631,In_2279);
xor U2993 (N_2993,In_1540,In_510);
nand U2994 (N_2994,In_1077,In_2544);
nor U2995 (N_2995,In_4754,In_1140);
nor U2996 (N_2996,In_1443,In_743);
nor U2997 (N_2997,In_2767,In_125);
or U2998 (N_2998,In_2242,In_2762);
nand U2999 (N_2999,In_316,In_862);
xor U3000 (N_3000,In_4927,In_849);
and U3001 (N_3001,In_4844,In_3319);
nand U3002 (N_3002,In_140,In_152);
and U3003 (N_3003,In_2226,In_4979);
or U3004 (N_3004,In_4006,In_4345);
xnor U3005 (N_3005,In_458,In_1541);
nand U3006 (N_3006,In_3448,In_4017);
nand U3007 (N_3007,In_2029,In_1439);
nand U3008 (N_3008,In_4298,In_610);
xnor U3009 (N_3009,In_2958,In_4511);
and U3010 (N_3010,In_195,In_3561);
and U3011 (N_3011,In_3477,In_1120);
nor U3012 (N_3012,In_175,In_4083);
or U3013 (N_3013,In_4088,In_3739);
nand U3014 (N_3014,In_1162,In_2529);
nor U3015 (N_3015,In_3662,In_3866);
nand U3016 (N_3016,In_975,In_2654);
and U3017 (N_3017,In_170,In_3609);
and U3018 (N_3018,In_4063,In_4255);
or U3019 (N_3019,In_1151,In_1268);
and U3020 (N_3020,In_484,In_3261);
or U3021 (N_3021,In_3875,In_2403);
and U3022 (N_3022,In_2520,In_4755);
nand U3023 (N_3023,In_4904,In_4319);
and U3024 (N_3024,In_4638,In_4108);
or U3025 (N_3025,In_3216,In_3233);
and U3026 (N_3026,In_3234,In_3039);
nand U3027 (N_3027,In_1331,In_3092);
nor U3028 (N_3028,In_2817,In_3178);
or U3029 (N_3029,In_673,In_3866);
or U3030 (N_3030,In_4936,In_193);
nand U3031 (N_3031,In_4561,In_1091);
and U3032 (N_3032,In_2097,In_3580);
and U3033 (N_3033,In_2411,In_34);
or U3034 (N_3034,In_2333,In_2505);
xnor U3035 (N_3035,In_2609,In_835);
nor U3036 (N_3036,In_863,In_1939);
nor U3037 (N_3037,In_3985,In_3479);
and U3038 (N_3038,In_2251,In_2317);
and U3039 (N_3039,In_3215,In_3947);
or U3040 (N_3040,In_54,In_845);
and U3041 (N_3041,In_187,In_3639);
xor U3042 (N_3042,In_4621,In_3620);
nor U3043 (N_3043,In_2345,In_2694);
or U3044 (N_3044,In_33,In_69);
nand U3045 (N_3045,In_3408,In_798);
and U3046 (N_3046,In_4072,In_1830);
and U3047 (N_3047,In_301,In_1366);
or U3048 (N_3048,In_3345,In_3249);
or U3049 (N_3049,In_4158,In_4773);
and U3050 (N_3050,In_4122,In_4624);
xnor U3051 (N_3051,In_3839,In_3569);
or U3052 (N_3052,In_3696,In_1669);
nor U3053 (N_3053,In_2227,In_3929);
and U3054 (N_3054,In_978,In_3861);
or U3055 (N_3055,In_4377,In_327);
xnor U3056 (N_3056,In_4398,In_4723);
and U3057 (N_3057,In_2788,In_1217);
nand U3058 (N_3058,In_4247,In_1710);
nand U3059 (N_3059,In_4095,In_4830);
nand U3060 (N_3060,In_2908,In_1669);
nor U3061 (N_3061,In_2873,In_3579);
and U3062 (N_3062,In_3800,In_3332);
nand U3063 (N_3063,In_3821,In_1030);
or U3064 (N_3064,In_365,In_3656);
nor U3065 (N_3065,In_2430,In_613);
or U3066 (N_3066,In_4072,In_923);
nor U3067 (N_3067,In_4206,In_4221);
nand U3068 (N_3068,In_4467,In_2440);
nand U3069 (N_3069,In_1518,In_2067);
nor U3070 (N_3070,In_3108,In_1804);
nand U3071 (N_3071,In_2172,In_714);
nand U3072 (N_3072,In_2782,In_4722);
nor U3073 (N_3073,In_4951,In_1288);
xnor U3074 (N_3074,In_3374,In_151);
nand U3075 (N_3075,In_2952,In_3672);
nor U3076 (N_3076,In_1499,In_424);
xor U3077 (N_3077,In_873,In_2998);
nand U3078 (N_3078,In_1486,In_1899);
nand U3079 (N_3079,In_4166,In_2060);
or U3080 (N_3080,In_3426,In_3853);
nand U3081 (N_3081,In_2340,In_612);
nor U3082 (N_3082,In_1862,In_2654);
nor U3083 (N_3083,In_4954,In_4136);
nand U3084 (N_3084,In_3276,In_2620);
and U3085 (N_3085,In_2173,In_821);
or U3086 (N_3086,In_1564,In_3317);
and U3087 (N_3087,In_4283,In_3379);
nand U3088 (N_3088,In_3366,In_241);
and U3089 (N_3089,In_418,In_4711);
and U3090 (N_3090,In_839,In_2738);
nand U3091 (N_3091,In_3047,In_414);
nand U3092 (N_3092,In_145,In_3442);
nand U3093 (N_3093,In_4955,In_4723);
nand U3094 (N_3094,In_1406,In_814);
nor U3095 (N_3095,In_4463,In_618);
or U3096 (N_3096,In_3932,In_4031);
or U3097 (N_3097,In_1165,In_4847);
and U3098 (N_3098,In_1394,In_979);
nand U3099 (N_3099,In_4077,In_2083);
xnor U3100 (N_3100,In_1610,In_3664);
nand U3101 (N_3101,In_566,In_4701);
nor U3102 (N_3102,In_3645,In_3593);
or U3103 (N_3103,In_3970,In_2043);
and U3104 (N_3104,In_3713,In_3265);
and U3105 (N_3105,In_1992,In_2463);
nand U3106 (N_3106,In_2350,In_3808);
and U3107 (N_3107,In_3414,In_3029);
and U3108 (N_3108,In_1554,In_1260);
xnor U3109 (N_3109,In_4583,In_600);
and U3110 (N_3110,In_3074,In_2484);
or U3111 (N_3111,In_4547,In_4425);
or U3112 (N_3112,In_947,In_4707);
nand U3113 (N_3113,In_252,In_4174);
or U3114 (N_3114,In_4665,In_713);
nand U3115 (N_3115,In_3138,In_4685);
or U3116 (N_3116,In_4832,In_77);
xnor U3117 (N_3117,In_2883,In_1578);
nand U3118 (N_3118,In_165,In_2561);
and U3119 (N_3119,In_11,In_3467);
xor U3120 (N_3120,In_1317,In_569);
nand U3121 (N_3121,In_602,In_2828);
or U3122 (N_3122,In_1902,In_1114);
nor U3123 (N_3123,In_618,In_1014);
nor U3124 (N_3124,In_682,In_520);
or U3125 (N_3125,In_2444,In_3708);
xnor U3126 (N_3126,In_1342,In_503);
and U3127 (N_3127,In_2193,In_4033);
and U3128 (N_3128,In_3072,In_732);
nor U3129 (N_3129,In_1716,In_3915);
and U3130 (N_3130,In_2189,In_4823);
or U3131 (N_3131,In_4464,In_2581);
nor U3132 (N_3132,In_1359,In_4285);
or U3133 (N_3133,In_3105,In_559);
or U3134 (N_3134,In_4107,In_4157);
or U3135 (N_3135,In_262,In_2324);
or U3136 (N_3136,In_3603,In_4886);
nor U3137 (N_3137,In_2011,In_1825);
and U3138 (N_3138,In_3088,In_1610);
nor U3139 (N_3139,In_1018,In_2103);
xor U3140 (N_3140,In_1254,In_4487);
nor U3141 (N_3141,In_4907,In_4639);
nor U3142 (N_3142,In_2275,In_317);
nand U3143 (N_3143,In_3604,In_585);
xor U3144 (N_3144,In_3135,In_4774);
nand U3145 (N_3145,In_598,In_2241);
or U3146 (N_3146,In_1302,In_3666);
nor U3147 (N_3147,In_442,In_2105);
xor U3148 (N_3148,In_302,In_236);
and U3149 (N_3149,In_395,In_2341);
nor U3150 (N_3150,In_4259,In_4141);
and U3151 (N_3151,In_2529,In_4374);
nor U3152 (N_3152,In_1042,In_3342);
nor U3153 (N_3153,In_1510,In_4488);
nand U3154 (N_3154,In_3958,In_4697);
nor U3155 (N_3155,In_2233,In_883);
nand U3156 (N_3156,In_954,In_2655);
xor U3157 (N_3157,In_3429,In_1590);
nand U3158 (N_3158,In_3997,In_1961);
or U3159 (N_3159,In_995,In_4254);
nor U3160 (N_3160,In_4665,In_1098);
and U3161 (N_3161,In_1839,In_3243);
nor U3162 (N_3162,In_1788,In_2723);
nor U3163 (N_3163,In_3152,In_2589);
or U3164 (N_3164,In_379,In_1028);
nor U3165 (N_3165,In_4797,In_4945);
nand U3166 (N_3166,In_1228,In_809);
and U3167 (N_3167,In_2530,In_3927);
nor U3168 (N_3168,In_1122,In_4914);
or U3169 (N_3169,In_4330,In_4590);
nor U3170 (N_3170,In_3792,In_1573);
and U3171 (N_3171,In_2559,In_3103);
or U3172 (N_3172,In_2176,In_4877);
nor U3173 (N_3173,In_4714,In_3698);
and U3174 (N_3174,In_4383,In_3585);
or U3175 (N_3175,In_4954,In_4531);
nand U3176 (N_3176,In_277,In_3681);
nor U3177 (N_3177,In_4506,In_2959);
nand U3178 (N_3178,In_2551,In_3279);
and U3179 (N_3179,In_1891,In_2894);
and U3180 (N_3180,In_3075,In_975);
and U3181 (N_3181,In_4537,In_814);
nand U3182 (N_3182,In_2881,In_3624);
nand U3183 (N_3183,In_146,In_1880);
and U3184 (N_3184,In_1203,In_4281);
or U3185 (N_3185,In_2131,In_2390);
nand U3186 (N_3186,In_1504,In_1232);
or U3187 (N_3187,In_1495,In_702);
nand U3188 (N_3188,In_3024,In_4712);
and U3189 (N_3189,In_3551,In_2965);
xor U3190 (N_3190,In_2811,In_3877);
nand U3191 (N_3191,In_1748,In_4502);
nand U3192 (N_3192,In_823,In_1649);
and U3193 (N_3193,In_2041,In_4377);
xnor U3194 (N_3194,In_2228,In_692);
and U3195 (N_3195,In_308,In_2912);
nor U3196 (N_3196,In_1783,In_2015);
nor U3197 (N_3197,In_3048,In_1758);
nor U3198 (N_3198,In_4487,In_582);
nand U3199 (N_3199,In_1555,In_1644);
or U3200 (N_3200,In_1730,In_3177);
nand U3201 (N_3201,In_2607,In_3940);
and U3202 (N_3202,In_959,In_4879);
nand U3203 (N_3203,In_105,In_2193);
xor U3204 (N_3204,In_1628,In_1513);
and U3205 (N_3205,In_4105,In_2909);
or U3206 (N_3206,In_4205,In_4468);
nor U3207 (N_3207,In_1159,In_3052);
or U3208 (N_3208,In_1892,In_2319);
and U3209 (N_3209,In_3429,In_1453);
and U3210 (N_3210,In_2064,In_4505);
nand U3211 (N_3211,In_967,In_3523);
nand U3212 (N_3212,In_1656,In_2195);
and U3213 (N_3213,In_3404,In_1444);
and U3214 (N_3214,In_4825,In_671);
nand U3215 (N_3215,In_741,In_3186);
nand U3216 (N_3216,In_974,In_3182);
nor U3217 (N_3217,In_3674,In_2118);
or U3218 (N_3218,In_1400,In_257);
and U3219 (N_3219,In_4172,In_1953);
or U3220 (N_3220,In_2966,In_575);
nand U3221 (N_3221,In_4836,In_3092);
or U3222 (N_3222,In_3818,In_709);
or U3223 (N_3223,In_4744,In_4775);
and U3224 (N_3224,In_3170,In_710);
nand U3225 (N_3225,In_1537,In_681);
xor U3226 (N_3226,In_220,In_277);
nor U3227 (N_3227,In_686,In_232);
and U3228 (N_3228,In_1710,In_2658);
nor U3229 (N_3229,In_207,In_4301);
nor U3230 (N_3230,In_3963,In_3295);
nor U3231 (N_3231,In_3261,In_574);
or U3232 (N_3232,In_39,In_2539);
nand U3233 (N_3233,In_1464,In_4222);
nor U3234 (N_3234,In_2865,In_650);
and U3235 (N_3235,In_2060,In_3556);
nor U3236 (N_3236,In_4672,In_4029);
and U3237 (N_3237,In_4359,In_4176);
or U3238 (N_3238,In_8,In_3473);
xor U3239 (N_3239,In_2781,In_4880);
and U3240 (N_3240,In_1977,In_1239);
nand U3241 (N_3241,In_4852,In_3112);
or U3242 (N_3242,In_4466,In_4949);
nand U3243 (N_3243,In_1008,In_4024);
and U3244 (N_3244,In_1046,In_4892);
or U3245 (N_3245,In_150,In_2425);
and U3246 (N_3246,In_698,In_2111);
nand U3247 (N_3247,In_2421,In_2291);
or U3248 (N_3248,In_3376,In_4256);
nand U3249 (N_3249,In_204,In_4883);
nor U3250 (N_3250,In_2633,In_3644);
or U3251 (N_3251,In_4316,In_2111);
nor U3252 (N_3252,In_1110,In_183);
nand U3253 (N_3253,In_1129,In_4839);
and U3254 (N_3254,In_2340,In_3445);
or U3255 (N_3255,In_3820,In_3981);
nor U3256 (N_3256,In_1625,In_2038);
nor U3257 (N_3257,In_1543,In_1829);
xor U3258 (N_3258,In_1056,In_3478);
nor U3259 (N_3259,In_4403,In_3035);
nand U3260 (N_3260,In_1426,In_807);
and U3261 (N_3261,In_2101,In_3557);
nand U3262 (N_3262,In_4286,In_2324);
nor U3263 (N_3263,In_4629,In_2756);
and U3264 (N_3264,In_3825,In_420);
and U3265 (N_3265,In_4583,In_3949);
and U3266 (N_3266,In_2552,In_4414);
nor U3267 (N_3267,In_3854,In_3954);
nor U3268 (N_3268,In_3943,In_2073);
or U3269 (N_3269,In_2964,In_850);
nand U3270 (N_3270,In_412,In_664);
xor U3271 (N_3271,In_1140,In_4252);
nor U3272 (N_3272,In_520,In_3722);
or U3273 (N_3273,In_4796,In_4528);
nor U3274 (N_3274,In_1572,In_1830);
nor U3275 (N_3275,In_2292,In_2133);
nand U3276 (N_3276,In_1654,In_3064);
nor U3277 (N_3277,In_4477,In_1203);
or U3278 (N_3278,In_1034,In_4518);
xnor U3279 (N_3279,In_4541,In_405);
nor U3280 (N_3280,In_53,In_1730);
nand U3281 (N_3281,In_3347,In_2666);
and U3282 (N_3282,In_1859,In_3427);
and U3283 (N_3283,In_4648,In_1071);
xnor U3284 (N_3284,In_738,In_3118);
nor U3285 (N_3285,In_4850,In_39);
nor U3286 (N_3286,In_1694,In_1373);
or U3287 (N_3287,In_1327,In_1792);
nor U3288 (N_3288,In_3451,In_3622);
and U3289 (N_3289,In_1153,In_1809);
nand U3290 (N_3290,In_319,In_1233);
and U3291 (N_3291,In_3559,In_1640);
nand U3292 (N_3292,In_3188,In_3557);
nor U3293 (N_3293,In_3606,In_1021);
nor U3294 (N_3294,In_2992,In_4135);
nor U3295 (N_3295,In_2692,In_2759);
and U3296 (N_3296,In_3117,In_601);
nor U3297 (N_3297,In_2325,In_1237);
and U3298 (N_3298,In_307,In_3445);
nand U3299 (N_3299,In_1799,In_2533);
xor U3300 (N_3300,In_4012,In_1616);
nor U3301 (N_3301,In_4598,In_1423);
nand U3302 (N_3302,In_3846,In_854);
and U3303 (N_3303,In_795,In_2300);
nor U3304 (N_3304,In_3861,In_4187);
nor U3305 (N_3305,In_543,In_4544);
nor U3306 (N_3306,In_603,In_1454);
nand U3307 (N_3307,In_999,In_2696);
or U3308 (N_3308,In_133,In_892);
or U3309 (N_3309,In_4047,In_472);
nand U3310 (N_3310,In_982,In_4722);
and U3311 (N_3311,In_3762,In_206);
nor U3312 (N_3312,In_2162,In_568);
xor U3313 (N_3313,In_322,In_1407);
or U3314 (N_3314,In_2307,In_205);
nor U3315 (N_3315,In_1877,In_1473);
nand U3316 (N_3316,In_4495,In_1060);
nor U3317 (N_3317,In_3313,In_3829);
xor U3318 (N_3318,In_4341,In_4173);
nand U3319 (N_3319,In_1391,In_2153);
nand U3320 (N_3320,In_4141,In_2612);
or U3321 (N_3321,In_2603,In_4495);
nor U3322 (N_3322,In_3590,In_694);
or U3323 (N_3323,In_4252,In_2918);
nand U3324 (N_3324,In_477,In_90);
nor U3325 (N_3325,In_4942,In_1303);
nand U3326 (N_3326,In_4717,In_473);
and U3327 (N_3327,In_4852,In_1109);
nor U3328 (N_3328,In_933,In_1536);
or U3329 (N_3329,In_3655,In_3605);
xor U3330 (N_3330,In_22,In_914);
and U3331 (N_3331,In_2612,In_1024);
nand U3332 (N_3332,In_3162,In_1375);
nor U3333 (N_3333,In_2435,In_774);
xnor U3334 (N_3334,In_2063,In_3651);
nand U3335 (N_3335,In_1329,In_2495);
nor U3336 (N_3336,In_919,In_3980);
and U3337 (N_3337,In_3166,In_3100);
xor U3338 (N_3338,In_4263,In_2758);
nand U3339 (N_3339,In_711,In_2749);
xor U3340 (N_3340,In_4449,In_77);
nor U3341 (N_3341,In_743,In_4245);
or U3342 (N_3342,In_2159,In_652);
nor U3343 (N_3343,In_4086,In_691);
nor U3344 (N_3344,In_3515,In_4093);
or U3345 (N_3345,In_877,In_793);
and U3346 (N_3346,In_777,In_354);
xnor U3347 (N_3347,In_484,In_3930);
nor U3348 (N_3348,In_416,In_1977);
and U3349 (N_3349,In_3553,In_3723);
and U3350 (N_3350,In_4873,In_4401);
nor U3351 (N_3351,In_2054,In_3422);
nand U3352 (N_3352,In_669,In_326);
and U3353 (N_3353,In_4721,In_3760);
or U3354 (N_3354,In_3980,In_4275);
nand U3355 (N_3355,In_4350,In_1180);
nor U3356 (N_3356,In_1257,In_1508);
xnor U3357 (N_3357,In_3622,In_2050);
and U3358 (N_3358,In_487,In_2247);
nor U3359 (N_3359,In_4208,In_3470);
and U3360 (N_3360,In_2770,In_3867);
nor U3361 (N_3361,In_95,In_2969);
nor U3362 (N_3362,In_3407,In_585);
nand U3363 (N_3363,In_4926,In_890);
nor U3364 (N_3364,In_390,In_3606);
xnor U3365 (N_3365,In_2605,In_2005);
xnor U3366 (N_3366,In_1238,In_147);
nor U3367 (N_3367,In_1265,In_898);
and U3368 (N_3368,In_1637,In_4780);
nand U3369 (N_3369,In_2816,In_700);
xnor U3370 (N_3370,In_2553,In_2374);
nor U3371 (N_3371,In_4670,In_3158);
nand U3372 (N_3372,In_4147,In_3906);
nor U3373 (N_3373,In_4433,In_1013);
or U3374 (N_3374,In_3466,In_934);
or U3375 (N_3375,In_685,In_2774);
nand U3376 (N_3376,In_2794,In_4412);
and U3377 (N_3377,In_3645,In_3139);
or U3378 (N_3378,In_4612,In_4353);
xnor U3379 (N_3379,In_1004,In_4097);
and U3380 (N_3380,In_3051,In_3428);
nor U3381 (N_3381,In_3995,In_3992);
nand U3382 (N_3382,In_2636,In_3303);
xor U3383 (N_3383,In_1807,In_1552);
nand U3384 (N_3384,In_2929,In_2862);
and U3385 (N_3385,In_1597,In_2760);
nand U3386 (N_3386,In_412,In_3396);
nand U3387 (N_3387,In_2833,In_2521);
nor U3388 (N_3388,In_1871,In_384);
nor U3389 (N_3389,In_4717,In_1363);
or U3390 (N_3390,In_1745,In_3640);
nor U3391 (N_3391,In_2715,In_3302);
and U3392 (N_3392,In_4646,In_926);
nand U3393 (N_3393,In_535,In_3249);
and U3394 (N_3394,In_4488,In_540);
xnor U3395 (N_3395,In_1268,In_2363);
or U3396 (N_3396,In_3775,In_2586);
nor U3397 (N_3397,In_3041,In_1760);
or U3398 (N_3398,In_1314,In_2883);
or U3399 (N_3399,In_4900,In_1623);
nor U3400 (N_3400,In_3635,In_1623);
or U3401 (N_3401,In_1254,In_3903);
nor U3402 (N_3402,In_2910,In_1379);
nand U3403 (N_3403,In_1804,In_4909);
nand U3404 (N_3404,In_611,In_2713);
xor U3405 (N_3405,In_2408,In_770);
or U3406 (N_3406,In_3011,In_2192);
xnor U3407 (N_3407,In_2796,In_4603);
nor U3408 (N_3408,In_4382,In_4205);
nor U3409 (N_3409,In_118,In_3798);
and U3410 (N_3410,In_2832,In_3813);
nor U3411 (N_3411,In_4244,In_4480);
or U3412 (N_3412,In_191,In_2993);
nor U3413 (N_3413,In_4380,In_303);
and U3414 (N_3414,In_2201,In_4083);
nand U3415 (N_3415,In_3981,In_706);
nand U3416 (N_3416,In_3304,In_3589);
or U3417 (N_3417,In_4876,In_265);
xor U3418 (N_3418,In_4088,In_6);
and U3419 (N_3419,In_4990,In_4440);
or U3420 (N_3420,In_1289,In_2148);
nand U3421 (N_3421,In_3606,In_891);
nor U3422 (N_3422,In_1824,In_3645);
nand U3423 (N_3423,In_1077,In_1259);
nor U3424 (N_3424,In_1848,In_1193);
and U3425 (N_3425,In_3005,In_4976);
nor U3426 (N_3426,In_516,In_1231);
and U3427 (N_3427,In_2390,In_4444);
and U3428 (N_3428,In_119,In_651);
nand U3429 (N_3429,In_765,In_3334);
or U3430 (N_3430,In_4121,In_4351);
nand U3431 (N_3431,In_1185,In_4103);
or U3432 (N_3432,In_1262,In_1524);
or U3433 (N_3433,In_610,In_3813);
nand U3434 (N_3434,In_534,In_2290);
xor U3435 (N_3435,In_2437,In_1582);
nand U3436 (N_3436,In_25,In_3485);
or U3437 (N_3437,In_1039,In_1028);
or U3438 (N_3438,In_3019,In_902);
or U3439 (N_3439,In_593,In_364);
nand U3440 (N_3440,In_4193,In_2682);
nand U3441 (N_3441,In_1406,In_3445);
xnor U3442 (N_3442,In_2408,In_3297);
or U3443 (N_3443,In_1466,In_2673);
nand U3444 (N_3444,In_2234,In_2303);
or U3445 (N_3445,In_1911,In_3930);
and U3446 (N_3446,In_856,In_1984);
nor U3447 (N_3447,In_4801,In_4642);
nand U3448 (N_3448,In_2386,In_3766);
nand U3449 (N_3449,In_3074,In_3712);
and U3450 (N_3450,In_4683,In_4251);
nand U3451 (N_3451,In_1611,In_2476);
and U3452 (N_3452,In_3581,In_4622);
nand U3453 (N_3453,In_3314,In_1840);
or U3454 (N_3454,In_2514,In_1764);
and U3455 (N_3455,In_4560,In_2114);
xnor U3456 (N_3456,In_751,In_3597);
xor U3457 (N_3457,In_2488,In_2877);
nor U3458 (N_3458,In_2635,In_428);
xor U3459 (N_3459,In_127,In_4822);
or U3460 (N_3460,In_25,In_2523);
nand U3461 (N_3461,In_2221,In_4382);
or U3462 (N_3462,In_1596,In_415);
or U3463 (N_3463,In_410,In_226);
nor U3464 (N_3464,In_3834,In_1421);
or U3465 (N_3465,In_1039,In_1244);
xor U3466 (N_3466,In_3257,In_1175);
and U3467 (N_3467,In_4602,In_1005);
and U3468 (N_3468,In_1235,In_3481);
xnor U3469 (N_3469,In_3286,In_1044);
nand U3470 (N_3470,In_712,In_702);
nand U3471 (N_3471,In_2780,In_2376);
nor U3472 (N_3472,In_2387,In_3738);
or U3473 (N_3473,In_4371,In_1641);
nor U3474 (N_3474,In_2467,In_2272);
nand U3475 (N_3475,In_2706,In_3341);
or U3476 (N_3476,In_4934,In_1810);
xnor U3477 (N_3477,In_4241,In_944);
nor U3478 (N_3478,In_413,In_1532);
nor U3479 (N_3479,In_3383,In_4239);
or U3480 (N_3480,In_4837,In_4138);
and U3481 (N_3481,In_2007,In_2493);
and U3482 (N_3482,In_1354,In_2208);
or U3483 (N_3483,In_3367,In_4495);
or U3484 (N_3484,In_3068,In_2681);
and U3485 (N_3485,In_4810,In_1621);
nand U3486 (N_3486,In_2605,In_2397);
nor U3487 (N_3487,In_1614,In_3728);
nand U3488 (N_3488,In_4728,In_1825);
and U3489 (N_3489,In_721,In_786);
nand U3490 (N_3490,In_1450,In_2667);
nand U3491 (N_3491,In_202,In_1566);
and U3492 (N_3492,In_3238,In_2858);
or U3493 (N_3493,In_3655,In_3881);
and U3494 (N_3494,In_3471,In_1253);
xor U3495 (N_3495,In_3395,In_4704);
and U3496 (N_3496,In_4255,In_1102);
nand U3497 (N_3497,In_3717,In_2297);
nand U3498 (N_3498,In_1717,In_1672);
nor U3499 (N_3499,In_1945,In_698);
or U3500 (N_3500,In_4052,In_2617);
nand U3501 (N_3501,In_3911,In_4918);
and U3502 (N_3502,In_3928,In_3908);
nand U3503 (N_3503,In_320,In_2338);
or U3504 (N_3504,In_4226,In_2933);
and U3505 (N_3505,In_1167,In_1602);
nand U3506 (N_3506,In_1851,In_369);
or U3507 (N_3507,In_4328,In_657);
or U3508 (N_3508,In_3502,In_1802);
nor U3509 (N_3509,In_966,In_4313);
or U3510 (N_3510,In_949,In_3013);
nor U3511 (N_3511,In_3529,In_4308);
and U3512 (N_3512,In_3964,In_3167);
nor U3513 (N_3513,In_1186,In_3699);
xor U3514 (N_3514,In_895,In_4025);
nor U3515 (N_3515,In_2003,In_2752);
and U3516 (N_3516,In_4777,In_1452);
or U3517 (N_3517,In_1825,In_984);
or U3518 (N_3518,In_2541,In_4917);
nor U3519 (N_3519,In_2307,In_4406);
nand U3520 (N_3520,In_2744,In_4639);
xnor U3521 (N_3521,In_2481,In_799);
and U3522 (N_3522,In_3873,In_855);
or U3523 (N_3523,In_8,In_4477);
or U3524 (N_3524,In_3441,In_4577);
nor U3525 (N_3525,In_2336,In_1241);
and U3526 (N_3526,In_2699,In_3839);
and U3527 (N_3527,In_1270,In_3700);
or U3528 (N_3528,In_340,In_271);
nor U3529 (N_3529,In_3363,In_3844);
and U3530 (N_3530,In_1596,In_3788);
nor U3531 (N_3531,In_1078,In_4018);
and U3532 (N_3532,In_126,In_2225);
nand U3533 (N_3533,In_4738,In_4402);
and U3534 (N_3534,In_4470,In_3054);
and U3535 (N_3535,In_3777,In_1597);
or U3536 (N_3536,In_522,In_47);
nor U3537 (N_3537,In_2529,In_3751);
and U3538 (N_3538,In_3370,In_1436);
nor U3539 (N_3539,In_2745,In_4127);
nand U3540 (N_3540,In_1615,In_4715);
nand U3541 (N_3541,In_2717,In_3926);
or U3542 (N_3542,In_2645,In_4474);
nor U3543 (N_3543,In_568,In_3116);
xnor U3544 (N_3544,In_1133,In_2625);
or U3545 (N_3545,In_82,In_4252);
nand U3546 (N_3546,In_3092,In_1939);
or U3547 (N_3547,In_1144,In_1412);
xor U3548 (N_3548,In_4550,In_1163);
or U3549 (N_3549,In_3206,In_252);
or U3550 (N_3550,In_4943,In_4811);
nand U3551 (N_3551,In_4285,In_693);
or U3552 (N_3552,In_4370,In_1277);
or U3553 (N_3553,In_4790,In_1215);
nor U3554 (N_3554,In_1240,In_292);
nand U3555 (N_3555,In_1672,In_1684);
nand U3556 (N_3556,In_1906,In_206);
and U3557 (N_3557,In_2263,In_2880);
or U3558 (N_3558,In_2914,In_3901);
nand U3559 (N_3559,In_964,In_422);
or U3560 (N_3560,In_1705,In_4173);
nor U3561 (N_3561,In_970,In_1455);
nor U3562 (N_3562,In_4069,In_2655);
nand U3563 (N_3563,In_377,In_1515);
or U3564 (N_3564,In_2950,In_694);
nand U3565 (N_3565,In_3877,In_3833);
or U3566 (N_3566,In_1125,In_1043);
nor U3567 (N_3567,In_785,In_3781);
and U3568 (N_3568,In_161,In_256);
or U3569 (N_3569,In_1669,In_315);
nor U3570 (N_3570,In_1554,In_2512);
or U3571 (N_3571,In_1744,In_2489);
xnor U3572 (N_3572,In_4443,In_4119);
nand U3573 (N_3573,In_896,In_4553);
nand U3574 (N_3574,In_4298,In_1097);
xor U3575 (N_3575,In_1558,In_1197);
and U3576 (N_3576,In_1825,In_4341);
nor U3577 (N_3577,In_464,In_4461);
and U3578 (N_3578,In_3769,In_3251);
nand U3579 (N_3579,In_2694,In_4025);
nand U3580 (N_3580,In_3246,In_3294);
and U3581 (N_3581,In_4064,In_4634);
and U3582 (N_3582,In_1611,In_1020);
or U3583 (N_3583,In_3403,In_1608);
and U3584 (N_3584,In_1374,In_667);
nand U3585 (N_3585,In_2807,In_1321);
nor U3586 (N_3586,In_2146,In_1669);
or U3587 (N_3587,In_4513,In_1634);
nand U3588 (N_3588,In_533,In_2937);
xor U3589 (N_3589,In_207,In_52);
nor U3590 (N_3590,In_2515,In_1387);
or U3591 (N_3591,In_2763,In_1880);
xor U3592 (N_3592,In_3983,In_3585);
nand U3593 (N_3593,In_614,In_1871);
or U3594 (N_3594,In_2525,In_230);
and U3595 (N_3595,In_4702,In_3325);
and U3596 (N_3596,In_4979,In_2825);
xnor U3597 (N_3597,In_3322,In_4671);
xor U3598 (N_3598,In_522,In_1845);
xor U3599 (N_3599,In_3828,In_1708);
or U3600 (N_3600,In_332,In_1056);
and U3601 (N_3601,In_1342,In_2838);
xor U3602 (N_3602,In_2611,In_1666);
or U3603 (N_3603,In_198,In_602);
nand U3604 (N_3604,In_2801,In_1866);
and U3605 (N_3605,In_464,In_1160);
or U3606 (N_3606,In_3081,In_2343);
or U3607 (N_3607,In_4088,In_2552);
and U3608 (N_3608,In_3822,In_4074);
or U3609 (N_3609,In_2558,In_4989);
nor U3610 (N_3610,In_2762,In_3378);
or U3611 (N_3611,In_3418,In_440);
nand U3612 (N_3612,In_799,In_4480);
and U3613 (N_3613,In_4244,In_3814);
and U3614 (N_3614,In_3613,In_1356);
or U3615 (N_3615,In_1674,In_549);
or U3616 (N_3616,In_1602,In_2440);
or U3617 (N_3617,In_3174,In_1167);
nand U3618 (N_3618,In_1904,In_1389);
nor U3619 (N_3619,In_3029,In_300);
nor U3620 (N_3620,In_2309,In_2363);
and U3621 (N_3621,In_413,In_4005);
xnor U3622 (N_3622,In_1127,In_4665);
xnor U3623 (N_3623,In_703,In_745);
nand U3624 (N_3624,In_192,In_4686);
and U3625 (N_3625,In_917,In_4257);
or U3626 (N_3626,In_1858,In_3230);
and U3627 (N_3627,In_1140,In_4053);
nor U3628 (N_3628,In_365,In_2322);
and U3629 (N_3629,In_1734,In_1111);
xnor U3630 (N_3630,In_257,In_2256);
or U3631 (N_3631,In_1916,In_3421);
or U3632 (N_3632,In_771,In_2455);
xnor U3633 (N_3633,In_3261,In_1552);
or U3634 (N_3634,In_3558,In_566);
nor U3635 (N_3635,In_1643,In_661);
nor U3636 (N_3636,In_3982,In_2854);
nand U3637 (N_3637,In_4476,In_3765);
and U3638 (N_3638,In_1962,In_1233);
nand U3639 (N_3639,In_932,In_1908);
nor U3640 (N_3640,In_2943,In_67);
xnor U3641 (N_3641,In_4035,In_2495);
or U3642 (N_3642,In_3117,In_3599);
nor U3643 (N_3643,In_4141,In_3495);
nand U3644 (N_3644,In_3775,In_1277);
nor U3645 (N_3645,In_3361,In_598);
nand U3646 (N_3646,In_4007,In_1436);
and U3647 (N_3647,In_3167,In_3509);
and U3648 (N_3648,In_868,In_2491);
or U3649 (N_3649,In_3540,In_952);
nand U3650 (N_3650,In_1978,In_786);
or U3651 (N_3651,In_2284,In_4582);
nand U3652 (N_3652,In_3173,In_3137);
and U3653 (N_3653,In_789,In_3215);
or U3654 (N_3654,In_3654,In_3590);
or U3655 (N_3655,In_2588,In_2041);
nand U3656 (N_3656,In_1681,In_527);
or U3657 (N_3657,In_3921,In_3533);
nand U3658 (N_3658,In_2885,In_501);
nand U3659 (N_3659,In_4717,In_2434);
or U3660 (N_3660,In_18,In_1106);
nor U3661 (N_3661,In_1304,In_4587);
nand U3662 (N_3662,In_4882,In_4317);
nand U3663 (N_3663,In_2372,In_3018);
xor U3664 (N_3664,In_3945,In_270);
nor U3665 (N_3665,In_1088,In_1721);
nor U3666 (N_3666,In_2237,In_3664);
and U3667 (N_3667,In_331,In_2754);
nand U3668 (N_3668,In_2007,In_3071);
nand U3669 (N_3669,In_2291,In_4472);
or U3670 (N_3670,In_3386,In_2178);
and U3671 (N_3671,In_253,In_3793);
or U3672 (N_3672,In_3421,In_1130);
nand U3673 (N_3673,In_19,In_3269);
or U3674 (N_3674,In_2998,In_2108);
nor U3675 (N_3675,In_398,In_2345);
or U3676 (N_3676,In_1643,In_2618);
nand U3677 (N_3677,In_4273,In_2798);
and U3678 (N_3678,In_3781,In_3443);
and U3679 (N_3679,In_1416,In_1139);
nand U3680 (N_3680,In_3625,In_356);
nor U3681 (N_3681,In_3670,In_494);
xor U3682 (N_3682,In_3281,In_4244);
or U3683 (N_3683,In_4728,In_2799);
or U3684 (N_3684,In_3002,In_788);
nand U3685 (N_3685,In_3200,In_2958);
xor U3686 (N_3686,In_4512,In_3348);
nor U3687 (N_3687,In_570,In_3674);
or U3688 (N_3688,In_3344,In_2970);
and U3689 (N_3689,In_3334,In_3180);
nand U3690 (N_3690,In_123,In_4044);
and U3691 (N_3691,In_396,In_2913);
nor U3692 (N_3692,In_3897,In_102);
and U3693 (N_3693,In_2748,In_2853);
or U3694 (N_3694,In_2694,In_3113);
nand U3695 (N_3695,In_1138,In_2864);
nand U3696 (N_3696,In_1592,In_1347);
nand U3697 (N_3697,In_4752,In_1255);
xnor U3698 (N_3698,In_4244,In_858);
xnor U3699 (N_3699,In_2726,In_663);
or U3700 (N_3700,In_1325,In_4857);
nand U3701 (N_3701,In_76,In_4632);
or U3702 (N_3702,In_1928,In_4119);
nand U3703 (N_3703,In_1785,In_643);
nand U3704 (N_3704,In_4057,In_2488);
and U3705 (N_3705,In_491,In_4389);
nor U3706 (N_3706,In_1011,In_4790);
nand U3707 (N_3707,In_4924,In_211);
nor U3708 (N_3708,In_3820,In_3152);
nor U3709 (N_3709,In_4637,In_828);
xor U3710 (N_3710,In_502,In_2835);
or U3711 (N_3711,In_4111,In_2699);
xor U3712 (N_3712,In_462,In_2596);
or U3713 (N_3713,In_756,In_845);
xnor U3714 (N_3714,In_1782,In_2191);
nor U3715 (N_3715,In_4080,In_2995);
xnor U3716 (N_3716,In_1815,In_2987);
nor U3717 (N_3717,In_549,In_653);
or U3718 (N_3718,In_117,In_4015);
xor U3719 (N_3719,In_2034,In_1298);
and U3720 (N_3720,In_3808,In_710);
and U3721 (N_3721,In_2198,In_458);
nor U3722 (N_3722,In_3524,In_1807);
or U3723 (N_3723,In_3400,In_168);
nor U3724 (N_3724,In_2573,In_1052);
or U3725 (N_3725,In_2645,In_3638);
and U3726 (N_3726,In_2113,In_3112);
or U3727 (N_3727,In_1856,In_4400);
nand U3728 (N_3728,In_4094,In_635);
xor U3729 (N_3729,In_3635,In_1209);
and U3730 (N_3730,In_207,In_2038);
nor U3731 (N_3731,In_607,In_4207);
xor U3732 (N_3732,In_1446,In_4469);
or U3733 (N_3733,In_4502,In_3768);
nand U3734 (N_3734,In_3230,In_568);
nand U3735 (N_3735,In_4482,In_3380);
nand U3736 (N_3736,In_2502,In_4514);
or U3737 (N_3737,In_2650,In_127);
or U3738 (N_3738,In_493,In_933);
xnor U3739 (N_3739,In_3372,In_1681);
and U3740 (N_3740,In_4578,In_3766);
nand U3741 (N_3741,In_3469,In_3601);
nor U3742 (N_3742,In_762,In_1959);
xor U3743 (N_3743,In_4472,In_854);
nor U3744 (N_3744,In_4702,In_2371);
or U3745 (N_3745,In_4723,In_1159);
and U3746 (N_3746,In_2142,In_4848);
and U3747 (N_3747,In_2646,In_2733);
nand U3748 (N_3748,In_3419,In_2836);
xor U3749 (N_3749,In_1460,In_1713);
nor U3750 (N_3750,In_4818,In_1503);
nor U3751 (N_3751,In_568,In_3831);
or U3752 (N_3752,In_562,In_416);
and U3753 (N_3753,In_526,In_2620);
nand U3754 (N_3754,In_3536,In_2248);
and U3755 (N_3755,In_530,In_78);
xnor U3756 (N_3756,In_4500,In_3419);
xnor U3757 (N_3757,In_2567,In_4407);
or U3758 (N_3758,In_1955,In_2048);
and U3759 (N_3759,In_3291,In_2191);
nor U3760 (N_3760,In_2136,In_4759);
nor U3761 (N_3761,In_2111,In_409);
nor U3762 (N_3762,In_3614,In_309);
nor U3763 (N_3763,In_3163,In_3730);
nand U3764 (N_3764,In_4509,In_1902);
nand U3765 (N_3765,In_2340,In_4194);
or U3766 (N_3766,In_2856,In_1478);
nand U3767 (N_3767,In_3081,In_1577);
or U3768 (N_3768,In_570,In_2754);
xnor U3769 (N_3769,In_2324,In_2661);
nand U3770 (N_3770,In_2746,In_1431);
nor U3771 (N_3771,In_3478,In_4973);
nand U3772 (N_3772,In_528,In_4876);
nor U3773 (N_3773,In_2789,In_1275);
and U3774 (N_3774,In_4823,In_4312);
nand U3775 (N_3775,In_3076,In_2782);
nand U3776 (N_3776,In_3057,In_2943);
xnor U3777 (N_3777,In_1818,In_800);
or U3778 (N_3778,In_4868,In_2406);
or U3779 (N_3779,In_4477,In_4117);
nand U3780 (N_3780,In_2953,In_1854);
nand U3781 (N_3781,In_2305,In_412);
xor U3782 (N_3782,In_3067,In_711);
and U3783 (N_3783,In_1563,In_4018);
nor U3784 (N_3784,In_3019,In_1001);
nor U3785 (N_3785,In_3659,In_4439);
xor U3786 (N_3786,In_1677,In_3556);
nand U3787 (N_3787,In_4585,In_1190);
nand U3788 (N_3788,In_2539,In_3600);
nand U3789 (N_3789,In_4210,In_1840);
or U3790 (N_3790,In_3781,In_175);
nand U3791 (N_3791,In_4614,In_2452);
or U3792 (N_3792,In_2751,In_4212);
nand U3793 (N_3793,In_1893,In_2110);
or U3794 (N_3794,In_3615,In_1959);
nor U3795 (N_3795,In_1006,In_2576);
nor U3796 (N_3796,In_144,In_1568);
nand U3797 (N_3797,In_570,In_4180);
or U3798 (N_3798,In_4445,In_3662);
nor U3799 (N_3799,In_250,In_273);
nor U3800 (N_3800,In_4915,In_4539);
nor U3801 (N_3801,In_310,In_617);
or U3802 (N_3802,In_3600,In_1645);
nor U3803 (N_3803,In_2364,In_1887);
nor U3804 (N_3804,In_4728,In_3638);
or U3805 (N_3805,In_2815,In_4051);
and U3806 (N_3806,In_3825,In_2528);
or U3807 (N_3807,In_2040,In_2576);
xnor U3808 (N_3808,In_3213,In_795);
nor U3809 (N_3809,In_2412,In_1132);
and U3810 (N_3810,In_2121,In_3617);
and U3811 (N_3811,In_3432,In_1414);
nand U3812 (N_3812,In_2559,In_3966);
nand U3813 (N_3813,In_263,In_4836);
xnor U3814 (N_3814,In_4126,In_2672);
xnor U3815 (N_3815,In_1495,In_1886);
or U3816 (N_3816,In_2750,In_445);
nor U3817 (N_3817,In_1450,In_4400);
nor U3818 (N_3818,In_3837,In_4646);
or U3819 (N_3819,In_141,In_2164);
nor U3820 (N_3820,In_4200,In_3118);
and U3821 (N_3821,In_1983,In_993);
or U3822 (N_3822,In_2499,In_201);
and U3823 (N_3823,In_4394,In_1343);
or U3824 (N_3824,In_3156,In_3918);
or U3825 (N_3825,In_4386,In_901);
nor U3826 (N_3826,In_1178,In_410);
xnor U3827 (N_3827,In_1844,In_1434);
xor U3828 (N_3828,In_3962,In_2200);
and U3829 (N_3829,In_4862,In_3411);
nor U3830 (N_3830,In_261,In_4540);
nand U3831 (N_3831,In_5,In_1464);
nand U3832 (N_3832,In_3475,In_3006);
nand U3833 (N_3833,In_3057,In_4509);
or U3834 (N_3834,In_866,In_3560);
and U3835 (N_3835,In_325,In_1738);
nand U3836 (N_3836,In_4872,In_1807);
and U3837 (N_3837,In_1429,In_1483);
or U3838 (N_3838,In_943,In_2206);
or U3839 (N_3839,In_4108,In_2334);
nand U3840 (N_3840,In_2509,In_383);
nand U3841 (N_3841,In_3101,In_4714);
xor U3842 (N_3842,In_3668,In_2713);
or U3843 (N_3843,In_226,In_3487);
xnor U3844 (N_3844,In_2561,In_80);
and U3845 (N_3845,In_3807,In_1251);
nor U3846 (N_3846,In_4361,In_4376);
and U3847 (N_3847,In_1213,In_2278);
or U3848 (N_3848,In_2786,In_2453);
nor U3849 (N_3849,In_614,In_3745);
or U3850 (N_3850,In_170,In_3653);
and U3851 (N_3851,In_612,In_87);
and U3852 (N_3852,In_735,In_41);
xnor U3853 (N_3853,In_4668,In_3950);
and U3854 (N_3854,In_3680,In_2849);
nor U3855 (N_3855,In_4711,In_3979);
nor U3856 (N_3856,In_3483,In_2952);
or U3857 (N_3857,In_266,In_1355);
nor U3858 (N_3858,In_3249,In_2804);
and U3859 (N_3859,In_291,In_3038);
or U3860 (N_3860,In_669,In_2826);
nand U3861 (N_3861,In_2322,In_1);
nand U3862 (N_3862,In_3097,In_2618);
and U3863 (N_3863,In_1038,In_4597);
and U3864 (N_3864,In_2147,In_2474);
xnor U3865 (N_3865,In_4696,In_1105);
nand U3866 (N_3866,In_2993,In_307);
nor U3867 (N_3867,In_1942,In_2618);
nor U3868 (N_3868,In_4221,In_937);
xor U3869 (N_3869,In_4098,In_701);
nand U3870 (N_3870,In_222,In_1781);
and U3871 (N_3871,In_2092,In_326);
or U3872 (N_3872,In_639,In_2291);
nand U3873 (N_3873,In_1809,In_1765);
or U3874 (N_3874,In_2260,In_3504);
and U3875 (N_3875,In_4665,In_4096);
nand U3876 (N_3876,In_1167,In_2160);
and U3877 (N_3877,In_2279,In_451);
and U3878 (N_3878,In_2257,In_479);
or U3879 (N_3879,In_3769,In_1343);
xor U3880 (N_3880,In_2212,In_2287);
xnor U3881 (N_3881,In_3404,In_2126);
nor U3882 (N_3882,In_4757,In_4255);
nand U3883 (N_3883,In_4848,In_2278);
nand U3884 (N_3884,In_1976,In_669);
or U3885 (N_3885,In_692,In_4371);
and U3886 (N_3886,In_2869,In_4132);
xnor U3887 (N_3887,In_1198,In_1479);
nor U3888 (N_3888,In_2598,In_636);
nor U3889 (N_3889,In_4340,In_4486);
and U3890 (N_3890,In_2401,In_684);
or U3891 (N_3891,In_1469,In_3774);
and U3892 (N_3892,In_2971,In_2913);
nand U3893 (N_3893,In_1762,In_1674);
or U3894 (N_3894,In_2548,In_4071);
nor U3895 (N_3895,In_1940,In_361);
xnor U3896 (N_3896,In_1049,In_1232);
nand U3897 (N_3897,In_2834,In_1320);
xnor U3898 (N_3898,In_4845,In_2348);
nand U3899 (N_3899,In_1846,In_4325);
nor U3900 (N_3900,In_4001,In_1162);
nor U3901 (N_3901,In_1095,In_1789);
nand U3902 (N_3902,In_931,In_3641);
nor U3903 (N_3903,In_2902,In_1748);
nor U3904 (N_3904,In_2939,In_463);
and U3905 (N_3905,In_869,In_1456);
and U3906 (N_3906,In_994,In_2087);
nand U3907 (N_3907,In_76,In_972);
nor U3908 (N_3908,In_4900,In_3556);
nand U3909 (N_3909,In_3070,In_2418);
nand U3910 (N_3910,In_1417,In_567);
or U3911 (N_3911,In_1613,In_547);
nand U3912 (N_3912,In_836,In_2891);
nor U3913 (N_3913,In_3650,In_1884);
and U3914 (N_3914,In_4211,In_2523);
or U3915 (N_3915,In_1530,In_1190);
or U3916 (N_3916,In_2195,In_953);
nor U3917 (N_3917,In_4110,In_3592);
or U3918 (N_3918,In_1183,In_2165);
nor U3919 (N_3919,In_4394,In_2584);
or U3920 (N_3920,In_1400,In_3408);
xnor U3921 (N_3921,In_3168,In_1180);
or U3922 (N_3922,In_4103,In_3046);
and U3923 (N_3923,In_4611,In_2131);
xnor U3924 (N_3924,In_4362,In_1543);
or U3925 (N_3925,In_4691,In_2810);
xor U3926 (N_3926,In_1069,In_2048);
xnor U3927 (N_3927,In_876,In_3149);
nand U3928 (N_3928,In_1458,In_2834);
or U3929 (N_3929,In_4182,In_3608);
and U3930 (N_3930,In_2539,In_2456);
or U3931 (N_3931,In_4966,In_3330);
nor U3932 (N_3932,In_1023,In_4099);
or U3933 (N_3933,In_1022,In_2220);
nor U3934 (N_3934,In_2153,In_2889);
or U3935 (N_3935,In_2030,In_3090);
xor U3936 (N_3936,In_1791,In_889);
nand U3937 (N_3937,In_902,In_3220);
or U3938 (N_3938,In_3804,In_4692);
and U3939 (N_3939,In_830,In_1079);
nor U3940 (N_3940,In_2917,In_4619);
nand U3941 (N_3941,In_810,In_4373);
and U3942 (N_3942,In_2966,In_3553);
and U3943 (N_3943,In_2195,In_4955);
or U3944 (N_3944,In_2638,In_2218);
nor U3945 (N_3945,In_4077,In_1117);
or U3946 (N_3946,In_4165,In_1431);
xnor U3947 (N_3947,In_245,In_1806);
nand U3948 (N_3948,In_30,In_2749);
nor U3949 (N_3949,In_2812,In_1475);
nand U3950 (N_3950,In_1549,In_815);
and U3951 (N_3951,In_2271,In_4414);
nor U3952 (N_3952,In_281,In_2475);
nor U3953 (N_3953,In_1967,In_4446);
nor U3954 (N_3954,In_1163,In_1476);
nor U3955 (N_3955,In_4976,In_1609);
and U3956 (N_3956,In_4424,In_319);
nor U3957 (N_3957,In_4458,In_3405);
nand U3958 (N_3958,In_4968,In_1023);
and U3959 (N_3959,In_1691,In_2622);
and U3960 (N_3960,In_4457,In_4817);
nor U3961 (N_3961,In_2994,In_1779);
nand U3962 (N_3962,In_836,In_925);
nor U3963 (N_3963,In_1815,In_360);
and U3964 (N_3964,In_2881,In_273);
and U3965 (N_3965,In_4020,In_4992);
nand U3966 (N_3966,In_4175,In_2667);
or U3967 (N_3967,In_3336,In_1103);
nor U3968 (N_3968,In_1619,In_2953);
and U3969 (N_3969,In_1103,In_2119);
nor U3970 (N_3970,In_4868,In_1390);
and U3971 (N_3971,In_3500,In_3826);
nand U3972 (N_3972,In_2387,In_1013);
nand U3973 (N_3973,In_1421,In_1971);
xor U3974 (N_3974,In_985,In_2299);
or U3975 (N_3975,In_1673,In_4247);
nand U3976 (N_3976,In_3576,In_2451);
nand U3977 (N_3977,In_3100,In_2436);
or U3978 (N_3978,In_4077,In_3318);
nand U3979 (N_3979,In_275,In_338);
nor U3980 (N_3980,In_3855,In_978);
nand U3981 (N_3981,In_3809,In_740);
or U3982 (N_3982,In_529,In_3517);
nor U3983 (N_3983,In_4945,In_4626);
nor U3984 (N_3984,In_1315,In_2873);
nand U3985 (N_3985,In_2542,In_4445);
and U3986 (N_3986,In_1015,In_920);
and U3987 (N_3987,In_3775,In_2720);
and U3988 (N_3988,In_2856,In_2595);
nand U3989 (N_3989,In_2259,In_3106);
or U3990 (N_3990,In_4545,In_2831);
nor U3991 (N_3991,In_65,In_1346);
nand U3992 (N_3992,In_3521,In_4063);
nand U3993 (N_3993,In_255,In_3482);
nor U3994 (N_3994,In_627,In_619);
nand U3995 (N_3995,In_2908,In_1405);
nor U3996 (N_3996,In_1464,In_4942);
xor U3997 (N_3997,In_2329,In_2975);
or U3998 (N_3998,In_2735,In_493);
nand U3999 (N_3999,In_2049,In_906);
nand U4000 (N_4000,In_4150,In_1251);
nand U4001 (N_4001,In_4783,In_3764);
xnor U4002 (N_4002,In_2248,In_1563);
nor U4003 (N_4003,In_562,In_1392);
and U4004 (N_4004,In_1445,In_4627);
and U4005 (N_4005,In_1340,In_2691);
xnor U4006 (N_4006,In_2942,In_53);
xor U4007 (N_4007,In_2441,In_4319);
and U4008 (N_4008,In_3785,In_662);
nor U4009 (N_4009,In_4827,In_4110);
and U4010 (N_4010,In_1666,In_666);
nand U4011 (N_4011,In_2692,In_3198);
and U4012 (N_4012,In_4428,In_3177);
or U4013 (N_4013,In_4819,In_2125);
or U4014 (N_4014,In_1695,In_4722);
nand U4015 (N_4015,In_4553,In_2913);
and U4016 (N_4016,In_2733,In_692);
nor U4017 (N_4017,In_3658,In_1878);
xor U4018 (N_4018,In_2770,In_3445);
and U4019 (N_4019,In_4623,In_2547);
nand U4020 (N_4020,In_3701,In_1848);
and U4021 (N_4021,In_1042,In_2056);
nor U4022 (N_4022,In_2664,In_1343);
xor U4023 (N_4023,In_769,In_3474);
or U4024 (N_4024,In_4222,In_770);
and U4025 (N_4025,In_938,In_907);
and U4026 (N_4026,In_4723,In_2577);
and U4027 (N_4027,In_3831,In_1765);
nand U4028 (N_4028,In_1954,In_761);
xnor U4029 (N_4029,In_4213,In_3858);
nor U4030 (N_4030,In_1906,In_1397);
and U4031 (N_4031,In_766,In_1270);
nand U4032 (N_4032,In_2462,In_2526);
and U4033 (N_4033,In_2472,In_2525);
nor U4034 (N_4034,In_4606,In_1075);
xor U4035 (N_4035,In_423,In_1615);
or U4036 (N_4036,In_375,In_1544);
and U4037 (N_4037,In_4934,In_376);
or U4038 (N_4038,In_925,In_3405);
nand U4039 (N_4039,In_497,In_1670);
xnor U4040 (N_4040,In_2785,In_3351);
or U4041 (N_4041,In_4658,In_579);
and U4042 (N_4042,In_1837,In_3848);
and U4043 (N_4043,In_405,In_4813);
and U4044 (N_4044,In_4112,In_1222);
nand U4045 (N_4045,In_1222,In_2005);
xnor U4046 (N_4046,In_4448,In_4378);
nor U4047 (N_4047,In_660,In_585);
nand U4048 (N_4048,In_2817,In_958);
xnor U4049 (N_4049,In_1547,In_2472);
or U4050 (N_4050,In_234,In_2626);
xor U4051 (N_4051,In_488,In_1908);
nor U4052 (N_4052,In_4424,In_3316);
xor U4053 (N_4053,In_1076,In_2401);
and U4054 (N_4054,In_1736,In_1544);
or U4055 (N_4055,In_90,In_2360);
nor U4056 (N_4056,In_337,In_4120);
nor U4057 (N_4057,In_3430,In_4633);
or U4058 (N_4058,In_1515,In_2905);
nor U4059 (N_4059,In_3438,In_1773);
nand U4060 (N_4060,In_3505,In_4025);
nor U4061 (N_4061,In_3465,In_2462);
xnor U4062 (N_4062,In_4460,In_1756);
nor U4063 (N_4063,In_4586,In_4862);
and U4064 (N_4064,In_3823,In_1538);
nand U4065 (N_4065,In_2762,In_2278);
nand U4066 (N_4066,In_3175,In_4937);
nand U4067 (N_4067,In_4841,In_812);
nor U4068 (N_4068,In_2294,In_558);
or U4069 (N_4069,In_2306,In_1879);
and U4070 (N_4070,In_3683,In_2946);
and U4071 (N_4071,In_2216,In_3920);
nand U4072 (N_4072,In_3413,In_1309);
nor U4073 (N_4073,In_2794,In_2165);
nor U4074 (N_4074,In_2825,In_4106);
or U4075 (N_4075,In_2432,In_1242);
nor U4076 (N_4076,In_4635,In_3637);
nor U4077 (N_4077,In_3176,In_41);
and U4078 (N_4078,In_217,In_2682);
or U4079 (N_4079,In_1923,In_2595);
or U4080 (N_4080,In_1124,In_3854);
nand U4081 (N_4081,In_2566,In_2075);
and U4082 (N_4082,In_3410,In_3411);
nand U4083 (N_4083,In_4232,In_491);
nor U4084 (N_4084,In_1290,In_409);
nor U4085 (N_4085,In_1396,In_4424);
or U4086 (N_4086,In_48,In_4546);
nand U4087 (N_4087,In_2958,In_2858);
and U4088 (N_4088,In_74,In_760);
and U4089 (N_4089,In_1734,In_4591);
nand U4090 (N_4090,In_1998,In_769);
nor U4091 (N_4091,In_2565,In_2287);
nor U4092 (N_4092,In_4304,In_4980);
xor U4093 (N_4093,In_147,In_117);
nand U4094 (N_4094,In_497,In_3218);
and U4095 (N_4095,In_1353,In_633);
and U4096 (N_4096,In_1065,In_3731);
nor U4097 (N_4097,In_1891,In_235);
and U4098 (N_4098,In_171,In_3551);
and U4099 (N_4099,In_245,In_4076);
and U4100 (N_4100,In_4945,In_1033);
and U4101 (N_4101,In_1106,In_667);
or U4102 (N_4102,In_68,In_2588);
nand U4103 (N_4103,In_160,In_3368);
nand U4104 (N_4104,In_4270,In_4348);
nor U4105 (N_4105,In_3396,In_1423);
xor U4106 (N_4106,In_2759,In_271);
nand U4107 (N_4107,In_4009,In_4735);
nand U4108 (N_4108,In_2735,In_3678);
nor U4109 (N_4109,In_4373,In_2631);
or U4110 (N_4110,In_4224,In_3582);
or U4111 (N_4111,In_4470,In_216);
nand U4112 (N_4112,In_2966,In_2911);
nor U4113 (N_4113,In_763,In_2213);
nand U4114 (N_4114,In_864,In_2722);
or U4115 (N_4115,In_1866,In_1799);
nor U4116 (N_4116,In_2474,In_4907);
and U4117 (N_4117,In_3550,In_4109);
nand U4118 (N_4118,In_1425,In_416);
nor U4119 (N_4119,In_1438,In_976);
xnor U4120 (N_4120,In_592,In_4074);
and U4121 (N_4121,In_1394,In_4894);
or U4122 (N_4122,In_2293,In_3083);
or U4123 (N_4123,In_1474,In_4887);
or U4124 (N_4124,In_287,In_3770);
or U4125 (N_4125,In_3093,In_4045);
nand U4126 (N_4126,In_426,In_402);
nor U4127 (N_4127,In_1974,In_3615);
xnor U4128 (N_4128,In_1432,In_4929);
nand U4129 (N_4129,In_709,In_522);
nor U4130 (N_4130,In_1626,In_942);
nor U4131 (N_4131,In_2833,In_2667);
or U4132 (N_4132,In_2561,In_4218);
or U4133 (N_4133,In_55,In_558);
nand U4134 (N_4134,In_4331,In_32);
and U4135 (N_4135,In_3406,In_1077);
and U4136 (N_4136,In_3090,In_4953);
and U4137 (N_4137,In_4787,In_4322);
or U4138 (N_4138,In_2201,In_4507);
or U4139 (N_4139,In_4785,In_2487);
nor U4140 (N_4140,In_2728,In_1431);
and U4141 (N_4141,In_4618,In_4854);
nor U4142 (N_4142,In_2091,In_1366);
nand U4143 (N_4143,In_747,In_819);
nand U4144 (N_4144,In_4623,In_2521);
nor U4145 (N_4145,In_476,In_587);
and U4146 (N_4146,In_1566,In_3014);
nor U4147 (N_4147,In_1880,In_658);
or U4148 (N_4148,In_686,In_945);
and U4149 (N_4149,In_1555,In_4313);
nor U4150 (N_4150,In_19,In_4445);
or U4151 (N_4151,In_1746,In_278);
nand U4152 (N_4152,In_2388,In_689);
nor U4153 (N_4153,In_1789,In_4773);
nor U4154 (N_4154,In_3787,In_1723);
nor U4155 (N_4155,In_3381,In_2967);
nor U4156 (N_4156,In_3470,In_3286);
nor U4157 (N_4157,In_3944,In_771);
nor U4158 (N_4158,In_2531,In_3839);
nand U4159 (N_4159,In_2394,In_568);
nand U4160 (N_4160,In_3416,In_420);
nor U4161 (N_4161,In_3483,In_36);
and U4162 (N_4162,In_1567,In_3016);
nor U4163 (N_4163,In_3917,In_4220);
and U4164 (N_4164,In_2160,In_4263);
and U4165 (N_4165,In_4677,In_3062);
or U4166 (N_4166,In_1060,In_2285);
or U4167 (N_4167,In_1165,In_998);
and U4168 (N_4168,In_302,In_3233);
or U4169 (N_4169,In_2816,In_1959);
xor U4170 (N_4170,In_500,In_1511);
or U4171 (N_4171,In_3393,In_4536);
or U4172 (N_4172,In_1425,In_2890);
or U4173 (N_4173,In_4738,In_838);
nor U4174 (N_4174,In_3998,In_2160);
nor U4175 (N_4175,In_2605,In_4879);
and U4176 (N_4176,In_894,In_3511);
nand U4177 (N_4177,In_1482,In_2688);
and U4178 (N_4178,In_2119,In_3453);
nor U4179 (N_4179,In_2709,In_4531);
nand U4180 (N_4180,In_3055,In_452);
nor U4181 (N_4181,In_2296,In_1966);
nor U4182 (N_4182,In_29,In_605);
or U4183 (N_4183,In_3588,In_3585);
or U4184 (N_4184,In_2468,In_4028);
or U4185 (N_4185,In_3067,In_1658);
or U4186 (N_4186,In_2354,In_1371);
or U4187 (N_4187,In_952,In_3881);
or U4188 (N_4188,In_1952,In_2761);
nand U4189 (N_4189,In_3104,In_274);
nand U4190 (N_4190,In_2921,In_733);
or U4191 (N_4191,In_645,In_4549);
or U4192 (N_4192,In_4391,In_2670);
nand U4193 (N_4193,In_966,In_243);
and U4194 (N_4194,In_413,In_2968);
and U4195 (N_4195,In_2036,In_3111);
or U4196 (N_4196,In_2401,In_2486);
and U4197 (N_4197,In_2790,In_1566);
xor U4198 (N_4198,In_2630,In_2788);
or U4199 (N_4199,In_1045,In_722);
and U4200 (N_4200,In_3937,In_3052);
or U4201 (N_4201,In_4659,In_2197);
nand U4202 (N_4202,In_175,In_2776);
or U4203 (N_4203,In_386,In_1038);
nand U4204 (N_4204,In_2886,In_1950);
xnor U4205 (N_4205,In_4643,In_2471);
or U4206 (N_4206,In_2611,In_1317);
nor U4207 (N_4207,In_2222,In_4193);
or U4208 (N_4208,In_1952,In_2972);
xor U4209 (N_4209,In_4095,In_3650);
nor U4210 (N_4210,In_2000,In_3728);
xnor U4211 (N_4211,In_3185,In_2891);
nand U4212 (N_4212,In_1557,In_220);
or U4213 (N_4213,In_871,In_3275);
xnor U4214 (N_4214,In_4426,In_1693);
or U4215 (N_4215,In_3344,In_866);
xnor U4216 (N_4216,In_1648,In_806);
xnor U4217 (N_4217,In_211,In_190);
nand U4218 (N_4218,In_2484,In_1180);
or U4219 (N_4219,In_4507,In_2537);
nand U4220 (N_4220,In_1925,In_4669);
nand U4221 (N_4221,In_592,In_2084);
nor U4222 (N_4222,In_2524,In_3268);
nor U4223 (N_4223,In_431,In_326);
and U4224 (N_4224,In_255,In_4213);
and U4225 (N_4225,In_372,In_459);
or U4226 (N_4226,In_4761,In_2368);
nor U4227 (N_4227,In_2321,In_4116);
and U4228 (N_4228,In_3087,In_1007);
nor U4229 (N_4229,In_4304,In_3074);
or U4230 (N_4230,In_2418,In_4965);
and U4231 (N_4231,In_2355,In_1874);
or U4232 (N_4232,In_4051,In_545);
and U4233 (N_4233,In_3915,In_1385);
nor U4234 (N_4234,In_1520,In_4358);
nor U4235 (N_4235,In_2538,In_3117);
xor U4236 (N_4236,In_1519,In_1297);
nor U4237 (N_4237,In_104,In_3590);
nor U4238 (N_4238,In_2191,In_4603);
and U4239 (N_4239,In_3980,In_1617);
and U4240 (N_4240,In_2700,In_2786);
nand U4241 (N_4241,In_1096,In_49);
and U4242 (N_4242,In_4311,In_4520);
and U4243 (N_4243,In_4536,In_11);
and U4244 (N_4244,In_3543,In_4814);
and U4245 (N_4245,In_2053,In_1153);
nor U4246 (N_4246,In_3456,In_1547);
nand U4247 (N_4247,In_2503,In_2333);
nor U4248 (N_4248,In_449,In_3351);
or U4249 (N_4249,In_884,In_386);
xor U4250 (N_4250,In_1224,In_1230);
nand U4251 (N_4251,In_2220,In_4462);
and U4252 (N_4252,In_2882,In_4539);
nor U4253 (N_4253,In_1891,In_4214);
or U4254 (N_4254,In_2888,In_2996);
nand U4255 (N_4255,In_2113,In_4237);
nand U4256 (N_4256,In_3641,In_661);
or U4257 (N_4257,In_2592,In_2220);
nor U4258 (N_4258,In_3969,In_501);
nand U4259 (N_4259,In_1585,In_4723);
nand U4260 (N_4260,In_369,In_4175);
nor U4261 (N_4261,In_1180,In_4804);
or U4262 (N_4262,In_3627,In_4185);
and U4263 (N_4263,In_1952,In_2658);
or U4264 (N_4264,In_4082,In_2098);
and U4265 (N_4265,In_2147,In_4667);
nand U4266 (N_4266,In_1589,In_4139);
nand U4267 (N_4267,In_4291,In_4255);
nand U4268 (N_4268,In_3841,In_3551);
nand U4269 (N_4269,In_1293,In_2969);
nand U4270 (N_4270,In_77,In_1019);
and U4271 (N_4271,In_184,In_1503);
nor U4272 (N_4272,In_3298,In_275);
nand U4273 (N_4273,In_440,In_619);
and U4274 (N_4274,In_2592,In_1251);
or U4275 (N_4275,In_4505,In_4526);
xnor U4276 (N_4276,In_1498,In_4284);
and U4277 (N_4277,In_765,In_189);
or U4278 (N_4278,In_77,In_1885);
or U4279 (N_4279,In_4904,In_1810);
nand U4280 (N_4280,In_147,In_1889);
or U4281 (N_4281,In_131,In_3237);
nand U4282 (N_4282,In_1890,In_3246);
nor U4283 (N_4283,In_4503,In_1887);
nor U4284 (N_4284,In_2694,In_3944);
and U4285 (N_4285,In_3283,In_768);
nor U4286 (N_4286,In_2413,In_3583);
xor U4287 (N_4287,In_4606,In_916);
or U4288 (N_4288,In_1630,In_2067);
nor U4289 (N_4289,In_1383,In_99);
nand U4290 (N_4290,In_784,In_4762);
nor U4291 (N_4291,In_3099,In_592);
and U4292 (N_4292,In_1885,In_3626);
and U4293 (N_4293,In_3082,In_834);
xnor U4294 (N_4294,In_1894,In_1975);
nor U4295 (N_4295,In_1005,In_1274);
or U4296 (N_4296,In_129,In_756);
and U4297 (N_4297,In_2608,In_2688);
and U4298 (N_4298,In_4141,In_4586);
or U4299 (N_4299,In_1100,In_2430);
and U4300 (N_4300,In_3076,In_2156);
nor U4301 (N_4301,In_2008,In_4955);
and U4302 (N_4302,In_4714,In_4082);
or U4303 (N_4303,In_2589,In_201);
nor U4304 (N_4304,In_2078,In_2093);
or U4305 (N_4305,In_2146,In_1074);
or U4306 (N_4306,In_316,In_421);
nand U4307 (N_4307,In_8,In_2912);
or U4308 (N_4308,In_795,In_3542);
nand U4309 (N_4309,In_720,In_1589);
nand U4310 (N_4310,In_2257,In_2825);
nor U4311 (N_4311,In_883,In_3410);
or U4312 (N_4312,In_3473,In_1042);
nand U4313 (N_4313,In_1580,In_1039);
or U4314 (N_4314,In_4602,In_3445);
or U4315 (N_4315,In_2358,In_760);
and U4316 (N_4316,In_3715,In_4138);
or U4317 (N_4317,In_3354,In_4301);
nand U4318 (N_4318,In_498,In_1809);
or U4319 (N_4319,In_1306,In_3270);
and U4320 (N_4320,In_1062,In_2264);
nand U4321 (N_4321,In_883,In_1241);
nand U4322 (N_4322,In_4430,In_881);
and U4323 (N_4323,In_3502,In_298);
xor U4324 (N_4324,In_2384,In_961);
nand U4325 (N_4325,In_2437,In_4614);
xor U4326 (N_4326,In_3592,In_3932);
nor U4327 (N_4327,In_2231,In_161);
nor U4328 (N_4328,In_3853,In_707);
or U4329 (N_4329,In_1602,In_2334);
or U4330 (N_4330,In_3300,In_1151);
nor U4331 (N_4331,In_2254,In_4612);
or U4332 (N_4332,In_4400,In_1092);
and U4333 (N_4333,In_4954,In_1040);
nor U4334 (N_4334,In_3382,In_1836);
nand U4335 (N_4335,In_3466,In_3772);
nand U4336 (N_4336,In_2181,In_3058);
or U4337 (N_4337,In_1951,In_4936);
xor U4338 (N_4338,In_2946,In_1016);
or U4339 (N_4339,In_4812,In_4675);
or U4340 (N_4340,In_4441,In_3175);
nand U4341 (N_4341,In_1374,In_338);
or U4342 (N_4342,In_298,In_1476);
and U4343 (N_4343,In_476,In_803);
or U4344 (N_4344,In_650,In_2880);
and U4345 (N_4345,In_2500,In_3859);
nand U4346 (N_4346,In_3231,In_2157);
and U4347 (N_4347,In_633,In_3605);
xor U4348 (N_4348,In_1550,In_2619);
nand U4349 (N_4349,In_3731,In_75);
and U4350 (N_4350,In_1248,In_1312);
nand U4351 (N_4351,In_749,In_1237);
and U4352 (N_4352,In_4527,In_3611);
nor U4353 (N_4353,In_122,In_1663);
nor U4354 (N_4354,In_1278,In_3434);
or U4355 (N_4355,In_734,In_851);
nand U4356 (N_4356,In_2841,In_1367);
nand U4357 (N_4357,In_3533,In_2547);
nor U4358 (N_4358,In_1093,In_2866);
and U4359 (N_4359,In_3148,In_3851);
or U4360 (N_4360,In_4456,In_1638);
or U4361 (N_4361,In_1882,In_2722);
or U4362 (N_4362,In_2007,In_3308);
or U4363 (N_4363,In_1928,In_3546);
nor U4364 (N_4364,In_4102,In_2089);
nor U4365 (N_4365,In_700,In_3411);
xnor U4366 (N_4366,In_3566,In_4076);
nand U4367 (N_4367,In_4498,In_4320);
nand U4368 (N_4368,In_148,In_4430);
or U4369 (N_4369,In_3637,In_4485);
or U4370 (N_4370,In_4300,In_1732);
xor U4371 (N_4371,In_1250,In_2852);
or U4372 (N_4372,In_3684,In_1337);
xor U4373 (N_4373,In_3954,In_2034);
nor U4374 (N_4374,In_4025,In_2796);
or U4375 (N_4375,In_2409,In_1937);
xnor U4376 (N_4376,In_909,In_636);
xor U4377 (N_4377,In_4526,In_722);
xor U4378 (N_4378,In_1777,In_1400);
nor U4379 (N_4379,In_4752,In_3635);
nor U4380 (N_4380,In_2273,In_1868);
or U4381 (N_4381,In_2647,In_1321);
and U4382 (N_4382,In_905,In_1575);
and U4383 (N_4383,In_668,In_4819);
nand U4384 (N_4384,In_4511,In_4449);
nor U4385 (N_4385,In_804,In_1107);
nand U4386 (N_4386,In_2431,In_4378);
xor U4387 (N_4387,In_2264,In_1905);
and U4388 (N_4388,In_253,In_570);
nand U4389 (N_4389,In_2537,In_762);
or U4390 (N_4390,In_3552,In_1136);
and U4391 (N_4391,In_4156,In_172);
or U4392 (N_4392,In_3882,In_673);
nor U4393 (N_4393,In_2916,In_1134);
and U4394 (N_4394,In_1954,In_486);
nor U4395 (N_4395,In_2533,In_597);
nand U4396 (N_4396,In_4033,In_4534);
nand U4397 (N_4397,In_1210,In_349);
or U4398 (N_4398,In_3719,In_3492);
and U4399 (N_4399,In_3886,In_1304);
nand U4400 (N_4400,In_4149,In_1591);
xnor U4401 (N_4401,In_1195,In_4145);
or U4402 (N_4402,In_4254,In_1647);
or U4403 (N_4403,In_3904,In_3117);
and U4404 (N_4404,In_2586,In_1216);
nor U4405 (N_4405,In_4103,In_3605);
or U4406 (N_4406,In_2829,In_3944);
and U4407 (N_4407,In_4983,In_277);
nand U4408 (N_4408,In_1882,In_4508);
nand U4409 (N_4409,In_3164,In_4467);
and U4410 (N_4410,In_993,In_1887);
or U4411 (N_4411,In_479,In_853);
or U4412 (N_4412,In_3563,In_1138);
or U4413 (N_4413,In_4119,In_3001);
xor U4414 (N_4414,In_2257,In_3672);
nand U4415 (N_4415,In_4563,In_3443);
or U4416 (N_4416,In_3211,In_1692);
or U4417 (N_4417,In_3506,In_4078);
or U4418 (N_4418,In_604,In_4343);
and U4419 (N_4419,In_314,In_3768);
xor U4420 (N_4420,In_335,In_790);
and U4421 (N_4421,In_4127,In_3860);
and U4422 (N_4422,In_157,In_1254);
nor U4423 (N_4423,In_2133,In_3559);
nor U4424 (N_4424,In_579,In_1500);
or U4425 (N_4425,In_732,In_3026);
xor U4426 (N_4426,In_1271,In_1576);
xor U4427 (N_4427,In_1325,In_1847);
or U4428 (N_4428,In_4476,In_916);
nand U4429 (N_4429,In_1652,In_3049);
xnor U4430 (N_4430,In_3256,In_2136);
nor U4431 (N_4431,In_3640,In_4599);
and U4432 (N_4432,In_3159,In_1145);
nor U4433 (N_4433,In_3497,In_1770);
nor U4434 (N_4434,In_2629,In_4200);
xnor U4435 (N_4435,In_2471,In_2443);
and U4436 (N_4436,In_3953,In_3535);
nand U4437 (N_4437,In_619,In_4203);
nand U4438 (N_4438,In_2701,In_4485);
and U4439 (N_4439,In_2016,In_2272);
and U4440 (N_4440,In_432,In_1614);
and U4441 (N_4441,In_3034,In_4075);
xor U4442 (N_4442,In_47,In_229);
and U4443 (N_4443,In_212,In_2687);
or U4444 (N_4444,In_3260,In_1846);
or U4445 (N_4445,In_1548,In_1924);
and U4446 (N_4446,In_201,In_1086);
and U4447 (N_4447,In_4751,In_4549);
or U4448 (N_4448,In_59,In_692);
nand U4449 (N_4449,In_3987,In_3788);
nand U4450 (N_4450,In_3082,In_348);
nor U4451 (N_4451,In_4100,In_1357);
nand U4452 (N_4452,In_1596,In_1280);
nor U4453 (N_4453,In_2774,In_990);
xnor U4454 (N_4454,In_4870,In_2734);
nor U4455 (N_4455,In_4456,In_3684);
nand U4456 (N_4456,In_4029,In_198);
nor U4457 (N_4457,In_3687,In_1669);
and U4458 (N_4458,In_1112,In_559);
nand U4459 (N_4459,In_1300,In_311);
or U4460 (N_4460,In_4962,In_1794);
and U4461 (N_4461,In_711,In_1480);
and U4462 (N_4462,In_4065,In_3351);
and U4463 (N_4463,In_1292,In_436);
or U4464 (N_4464,In_2460,In_1106);
or U4465 (N_4465,In_3566,In_4446);
or U4466 (N_4466,In_4796,In_4731);
nand U4467 (N_4467,In_2623,In_3909);
or U4468 (N_4468,In_1310,In_1763);
nand U4469 (N_4469,In_449,In_4425);
and U4470 (N_4470,In_3180,In_1663);
and U4471 (N_4471,In_1309,In_2460);
or U4472 (N_4472,In_1179,In_636);
xor U4473 (N_4473,In_1284,In_1530);
xnor U4474 (N_4474,In_220,In_3084);
nand U4475 (N_4475,In_4720,In_2629);
nor U4476 (N_4476,In_3103,In_4044);
and U4477 (N_4477,In_1532,In_1564);
nor U4478 (N_4478,In_1503,In_894);
nor U4479 (N_4479,In_834,In_1999);
or U4480 (N_4480,In_4508,In_1629);
and U4481 (N_4481,In_608,In_1781);
xnor U4482 (N_4482,In_2034,In_386);
nor U4483 (N_4483,In_1095,In_9);
xnor U4484 (N_4484,In_2393,In_4996);
and U4485 (N_4485,In_4066,In_2370);
xor U4486 (N_4486,In_447,In_4241);
and U4487 (N_4487,In_4831,In_3347);
nand U4488 (N_4488,In_3456,In_266);
or U4489 (N_4489,In_1071,In_378);
or U4490 (N_4490,In_1498,In_2415);
or U4491 (N_4491,In_3771,In_2239);
nand U4492 (N_4492,In_4054,In_1437);
or U4493 (N_4493,In_1879,In_4331);
nand U4494 (N_4494,In_350,In_4675);
or U4495 (N_4495,In_3287,In_4924);
and U4496 (N_4496,In_2133,In_1435);
and U4497 (N_4497,In_4512,In_3501);
and U4498 (N_4498,In_4387,In_4815);
nor U4499 (N_4499,In_872,In_2112);
nand U4500 (N_4500,In_1971,In_1888);
or U4501 (N_4501,In_1379,In_4376);
and U4502 (N_4502,In_1402,In_1455);
nor U4503 (N_4503,In_141,In_1279);
nand U4504 (N_4504,In_972,In_4064);
nand U4505 (N_4505,In_1759,In_997);
nor U4506 (N_4506,In_1201,In_3972);
xor U4507 (N_4507,In_3690,In_3825);
xor U4508 (N_4508,In_3848,In_4486);
nor U4509 (N_4509,In_765,In_4611);
and U4510 (N_4510,In_746,In_4076);
nor U4511 (N_4511,In_1498,In_297);
nand U4512 (N_4512,In_4280,In_2820);
or U4513 (N_4513,In_3345,In_2809);
and U4514 (N_4514,In_44,In_1625);
and U4515 (N_4515,In_213,In_2192);
or U4516 (N_4516,In_4599,In_2622);
xor U4517 (N_4517,In_1991,In_2578);
and U4518 (N_4518,In_4987,In_459);
and U4519 (N_4519,In_3880,In_2216);
or U4520 (N_4520,In_4422,In_3634);
xor U4521 (N_4521,In_1041,In_520);
and U4522 (N_4522,In_4864,In_2651);
nand U4523 (N_4523,In_3814,In_4459);
nor U4524 (N_4524,In_2871,In_3927);
xnor U4525 (N_4525,In_971,In_3784);
or U4526 (N_4526,In_3118,In_927);
and U4527 (N_4527,In_3966,In_4590);
nand U4528 (N_4528,In_3154,In_512);
or U4529 (N_4529,In_2923,In_3734);
and U4530 (N_4530,In_435,In_1911);
or U4531 (N_4531,In_3696,In_328);
and U4532 (N_4532,In_1426,In_2059);
nor U4533 (N_4533,In_4449,In_3118);
nor U4534 (N_4534,In_2556,In_4331);
or U4535 (N_4535,In_1121,In_1927);
nand U4536 (N_4536,In_4447,In_741);
nor U4537 (N_4537,In_4576,In_273);
and U4538 (N_4538,In_3731,In_4566);
nor U4539 (N_4539,In_4539,In_2255);
nor U4540 (N_4540,In_483,In_2884);
and U4541 (N_4541,In_3023,In_4131);
or U4542 (N_4542,In_4254,In_3513);
or U4543 (N_4543,In_2623,In_30);
or U4544 (N_4544,In_1553,In_1147);
and U4545 (N_4545,In_557,In_2677);
nand U4546 (N_4546,In_2132,In_16);
nor U4547 (N_4547,In_4548,In_4409);
and U4548 (N_4548,In_396,In_4680);
nand U4549 (N_4549,In_1223,In_3347);
nand U4550 (N_4550,In_817,In_4333);
nand U4551 (N_4551,In_985,In_3116);
nand U4552 (N_4552,In_4657,In_2009);
nand U4553 (N_4553,In_2509,In_2492);
xnor U4554 (N_4554,In_2932,In_4597);
nor U4555 (N_4555,In_557,In_1712);
or U4556 (N_4556,In_2865,In_1147);
nand U4557 (N_4557,In_4746,In_1546);
xor U4558 (N_4558,In_4251,In_2490);
nand U4559 (N_4559,In_2555,In_925);
nor U4560 (N_4560,In_201,In_1140);
or U4561 (N_4561,In_1705,In_835);
and U4562 (N_4562,In_2470,In_4213);
nand U4563 (N_4563,In_2529,In_1070);
nand U4564 (N_4564,In_348,In_4539);
or U4565 (N_4565,In_2971,In_3291);
nor U4566 (N_4566,In_2199,In_3586);
or U4567 (N_4567,In_430,In_2622);
or U4568 (N_4568,In_4006,In_2962);
nor U4569 (N_4569,In_2572,In_3432);
and U4570 (N_4570,In_859,In_781);
and U4571 (N_4571,In_4487,In_4900);
or U4572 (N_4572,In_3648,In_2714);
xnor U4573 (N_4573,In_4131,In_3244);
nor U4574 (N_4574,In_4198,In_1947);
xnor U4575 (N_4575,In_1425,In_2173);
nor U4576 (N_4576,In_3670,In_379);
or U4577 (N_4577,In_4630,In_2770);
nor U4578 (N_4578,In_4093,In_3037);
or U4579 (N_4579,In_4211,In_3497);
or U4580 (N_4580,In_4332,In_4046);
nor U4581 (N_4581,In_4582,In_1003);
nand U4582 (N_4582,In_2599,In_1261);
and U4583 (N_4583,In_1507,In_2081);
nor U4584 (N_4584,In_439,In_4907);
and U4585 (N_4585,In_2103,In_2961);
or U4586 (N_4586,In_2598,In_4699);
or U4587 (N_4587,In_1429,In_568);
xor U4588 (N_4588,In_2606,In_879);
nand U4589 (N_4589,In_1393,In_2404);
and U4590 (N_4590,In_3945,In_4409);
and U4591 (N_4591,In_4094,In_1616);
nor U4592 (N_4592,In_1176,In_1509);
xor U4593 (N_4593,In_1154,In_3722);
and U4594 (N_4594,In_2703,In_3371);
nand U4595 (N_4595,In_3862,In_2470);
nor U4596 (N_4596,In_4648,In_314);
nand U4597 (N_4597,In_1161,In_475);
nor U4598 (N_4598,In_3329,In_3442);
xnor U4599 (N_4599,In_4208,In_1828);
nand U4600 (N_4600,In_1911,In_873);
and U4601 (N_4601,In_340,In_4688);
and U4602 (N_4602,In_4526,In_2414);
nor U4603 (N_4603,In_3403,In_2966);
nor U4604 (N_4604,In_2392,In_3068);
nand U4605 (N_4605,In_1566,In_4677);
nand U4606 (N_4606,In_2988,In_1022);
or U4607 (N_4607,In_2202,In_2221);
nand U4608 (N_4608,In_3600,In_3631);
xor U4609 (N_4609,In_3356,In_3126);
nor U4610 (N_4610,In_3383,In_3145);
or U4611 (N_4611,In_4302,In_4103);
xor U4612 (N_4612,In_2654,In_1287);
nor U4613 (N_4613,In_1496,In_2512);
nor U4614 (N_4614,In_4089,In_3732);
xor U4615 (N_4615,In_3492,In_762);
nor U4616 (N_4616,In_3950,In_2265);
nor U4617 (N_4617,In_2554,In_616);
nor U4618 (N_4618,In_3919,In_4573);
nand U4619 (N_4619,In_4410,In_3144);
nor U4620 (N_4620,In_2068,In_1548);
or U4621 (N_4621,In_1688,In_3689);
and U4622 (N_4622,In_1956,In_4025);
nand U4623 (N_4623,In_4081,In_4704);
or U4624 (N_4624,In_4106,In_3364);
nor U4625 (N_4625,In_4366,In_4616);
or U4626 (N_4626,In_4720,In_1430);
or U4627 (N_4627,In_3184,In_4270);
nor U4628 (N_4628,In_659,In_826);
or U4629 (N_4629,In_4045,In_4989);
nor U4630 (N_4630,In_1893,In_2721);
or U4631 (N_4631,In_1682,In_1396);
nand U4632 (N_4632,In_815,In_4186);
and U4633 (N_4633,In_297,In_1811);
or U4634 (N_4634,In_1587,In_3991);
xor U4635 (N_4635,In_2970,In_2134);
nor U4636 (N_4636,In_4476,In_4792);
nand U4637 (N_4637,In_587,In_1351);
nor U4638 (N_4638,In_2317,In_638);
and U4639 (N_4639,In_2270,In_2684);
and U4640 (N_4640,In_1830,In_3509);
nor U4641 (N_4641,In_2045,In_3815);
nand U4642 (N_4642,In_1317,In_2874);
or U4643 (N_4643,In_3339,In_2576);
nand U4644 (N_4644,In_4143,In_4110);
or U4645 (N_4645,In_2243,In_1749);
nand U4646 (N_4646,In_504,In_3782);
or U4647 (N_4647,In_399,In_542);
or U4648 (N_4648,In_3813,In_4073);
nor U4649 (N_4649,In_2414,In_3436);
or U4650 (N_4650,In_4943,In_818);
or U4651 (N_4651,In_4517,In_341);
nor U4652 (N_4652,In_2653,In_299);
nand U4653 (N_4653,In_2679,In_757);
xnor U4654 (N_4654,In_3051,In_7);
or U4655 (N_4655,In_612,In_164);
nand U4656 (N_4656,In_832,In_444);
nand U4657 (N_4657,In_3821,In_3026);
xor U4658 (N_4658,In_3541,In_4302);
nor U4659 (N_4659,In_3845,In_4441);
nor U4660 (N_4660,In_537,In_3828);
and U4661 (N_4661,In_1890,In_1630);
nor U4662 (N_4662,In_4612,In_900);
xor U4663 (N_4663,In_2895,In_1528);
nand U4664 (N_4664,In_4741,In_3931);
nor U4665 (N_4665,In_357,In_789);
nor U4666 (N_4666,In_4183,In_365);
xor U4667 (N_4667,In_827,In_3044);
or U4668 (N_4668,In_1317,In_386);
and U4669 (N_4669,In_3313,In_484);
nor U4670 (N_4670,In_3359,In_2764);
nand U4671 (N_4671,In_440,In_4471);
or U4672 (N_4672,In_2175,In_2388);
and U4673 (N_4673,In_1243,In_369);
xor U4674 (N_4674,In_4659,In_687);
nor U4675 (N_4675,In_2103,In_1793);
nand U4676 (N_4676,In_635,In_2008);
or U4677 (N_4677,In_345,In_1524);
and U4678 (N_4678,In_3074,In_1136);
nor U4679 (N_4679,In_4896,In_1419);
nand U4680 (N_4680,In_1428,In_241);
nor U4681 (N_4681,In_1882,In_3655);
or U4682 (N_4682,In_4832,In_2852);
or U4683 (N_4683,In_4014,In_3058);
xor U4684 (N_4684,In_2632,In_4774);
nand U4685 (N_4685,In_3414,In_4223);
or U4686 (N_4686,In_2220,In_4871);
and U4687 (N_4687,In_2697,In_1274);
and U4688 (N_4688,In_221,In_4298);
nor U4689 (N_4689,In_946,In_4999);
and U4690 (N_4690,In_1550,In_1563);
and U4691 (N_4691,In_844,In_4181);
or U4692 (N_4692,In_4816,In_2731);
nor U4693 (N_4693,In_3764,In_286);
and U4694 (N_4694,In_3075,In_3527);
nand U4695 (N_4695,In_151,In_3974);
nand U4696 (N_4696,In_3474,In_4045);
and U4697 (N_4697,In_3295,In_345);
and U4698 (N_4698,In_215,In_3654);
or U4699 (N_4699,In_2612,In_4123);
and U4700 (N_4700,In_538,In_382);
nor U4701 (N_4701,In_1300,In_4239);
nor U4702 (N_4702,In_2678,In_4430);
nand U4703 (N_4703,In_2580,In_4763);
nor U4704 (N_4704,In_338,In_4171);
nand U4705 (N_4705,In_3464,In_1335);
nand U4706 (N_4706,In_1986,In_502);
and U4707 (N_4707,In_4740,In_1240);
and U4708 (N_4708,In_474,In_1231);
nand U4709 (N_4709,In_3808,In_3613);
nand U4710 (N_4710,In_4900,In_1639);
xnor U4711 (N_4711,In_4439,In_2218);
and U4712 (N_4712,In_108,In_1584);
nor U4713 (N_4713,In_4451,In_629);
nor U4714 (N_4714,In_4897,In_1084);
and U4715 (N_4715,In_3169,In_1460);
nor U4716 (N_4716,In_2573,In_4573);
nor U4717 (N_4717,In_637,In_4856);
or U4718 (N_4718,In_4360,In_1862);
nor U4719 (N_4719,In_4935,In_4031);
and U4720 (N_4720,In_4059,In_355);
and U4721 (N_4721,In_2970,In_1367);
xor U4722 (N_4722,In_411,In_2276);
nand U4723 (N_4723,In_1565,In_1888);
nand U4724 (N_4724,In_1491,In_1656);
nand U4725 (N_4725,In_1062,In_1024);
nand U4726 (N_4726,In_1131,In_3245);
nand U4727 (N_4727,In_1616,In_2663);
or U4728 (N_4728,In_3283,In_2158);
nor U4729 (N_4729,In_2348,In_3135);
nor U4730 (N_4730,In_3585,In_948);
xnor U4731 (N_4731,In_4774,In_2024);
or U4732 (N_4732,In_2599,In_2991);
or U4733 (N_4733,In_1286,In_457);
nor U4734 (N_4734,In_534,In_1317);
nor U4735 (N_4735,In_4388,In_1519);
nor U4736 (N_4736,In_3635,In_1109);
nor U4737 (N_4737,In_1448,In_1875);
and U4738 (N_4738,In_4489,In_2261);
or U4739 (N_4739,In_2094,In_4166);
nand U4740 (N_4740,In_909,In_2971);
nand U4741 (N_4741,In_244,In_1978);
and U4742 (N_4742,In_2808,In_241);
and U4743 (N_4743,In_3035,In_4951);
nand U4744 (N_4744,In_2880,In_914);
or U4745 (N_4745,In_97,In_3435);
or U4746 (N_4746,In_1945,In_4597);
and U4747 (N_4747,In_2781,In_1573);
and U4748 (N_4748,In_1704,In_927);
xor U4749 (N_4749,In_4053,In_503);
nor U4750 (N_4750,In_519,In_200);
nand U4751 (N_4751,In_275,In_1690);
and U4752 (N_4752,In_433,In_91);
nand U4753 (N_4753,In_1808,In_2407);
nand U4754 (N_4754,In_1920,In_1706);
nand U4755 (N_4755,In_2618,In_2708);
or U4756 (N_4756,In_3368,In_7);
nand U4757 (N_4757,In_4324,In_1551);
or U4758 (N_4758,In_332,In_2006);
and U4759 (N_4759,In_685,In_135);
and U4760 (N_4760,In_3430,In_658);
nand U4761 (N_4761,In_3935,In_4962);
or U4762 (N_4762,In_1713,In_1175);
and U4763 (N_4763,In_1730,In_1624);
nand U4764 (N_4764,In_126,In_4834);
nand U4765 (N_4765,In_1007,In_870);
nand U4766 (N_4766,In_3560,In_3620);
or U4767 (N_4767,In_835,In_1451);
or U4768 (N_4768,In_1608,In_42);
nand U4769 (N_4769,In_4390,In_1172);
nor U4770 (N_4770,In_970,In_3354);
and U4771 (N_4771,In_1326,In_4787);
nand U4772 (N_4772,In_2129,In_2444);
nand U4773 (N_4773,In_1364,In_2488);
or U4774 (N_4774,In_111,In_599);
nor U4775 (N_4775,In_114,In_3829);
and U4776 (N_4776,In_840,In_4317);
nand U4777 (N_4777,In_1661,In_3239);
and U4778 (N_4778,In_212,In_1753);
xnor U4779 (N_4779,In_3141,In_5);
and U4780 (N_4780,In_3309,In_1701);
nor U4781 (N_4781,In_1036,In_1992);
and U4782 (N_4782,In_1372,In_388);
nor U4783 (N_4783,In_4776,In_295);
nor U4784 (N_4784,In_1164,In_4236);
nand U4785 (N_4785,In_481,In_3205);
xnor U4786 (N_4786,In_4555,In_4761);
and U4787 (N_4787,In_829,In_378);
and U4788 (N_4788,In_2018,In_1729);
xor U4789 (N_4789,In_271,In_2280);
nand U4790 (N_4790,In_909,In_4522);
and U4791 (N_4791,In_114,In_683);
or U4792 (N_4792,In_1588,In_1820);
and U4793 (N_4793,In_3051,In_284);
nand U4794 (N_4794,In_1917,In_1292);
or U4795 (N_4795,In_813,In_3652);
and U4796 (N_4796,In_796,In_56);
or U4797 (N_4797,In_2811,In_819);
nand U4798 (N_4798,In_2995,In_883);
or U4799 (N_4799,In_3197,In_2479);
or U4800 (N_4800,In_3377,In_2016);
or U4801 (N_4801,In_4746,In_853);
nor U4802 (N_4802,In_719,In_3352);
and U4803 (N_4803,In_2434,In_1851);
nand U4804 (N_4804,In_182,In_4189);
nor U4805 (N_4805,In_340,In_3783);
and U4806 (N_4806,In_988,In_3222);
and U4807 (N_4807,In_430,In_4334);
xor U4808 (N_4808,In_3089,In_2767);
and U4809 (N_4809,In_4368,In_4164);
or U4810 (N_4810,In_4541,In_380);
nor U4811 (N_4811,In_2669,In_4453);
and U4812 (N_4812,In_23,In_870);
nor U4813 (N_4813,In_3564,In_3802);
and U4814 (N_4814,In_511,In_3626);
and U4815 (N_4815,In_3308,In_875);
nand U4816 (N_4816,In_4152,In_2330);
or U4817 (N_4817,In_2202,In_4741);
and U4818 (N_4818,In_1496,In_1861);
xor U4819 (N_4819,In_4751,In_1960);
and U4820 (N_4820,In_2196,In_1767);
and U4821 (N_4821,In_4146,In_1033);
or U4822 (N_4822,In_954,In_3497);
nor U4823 (N_4823,In_3168,In_4898);
nand U4824 (N_4824,In_718,In_404);
and U4825 (N_4825,In_1826,In_4818);
xnor U4826 (N_4826,In_3074,In_4852);
nor U4827 (N_4827,In_1334,In_2681);
and U4828 (N_4828,In_1946,In_2462);
nand U4829 (N_4829,In_2048,In_375);
and U4830 (N_4830,In_4525,In_1850);
nand U4831 (N_4831,In_1289,In_1822);
xor U4832 (N_4832,In_4210,In_2656);
nor U4833 (N_4833,In_57,In_2232);
and U4834 (N_4834,In_1051,In_519);
xor U4835 (N_4835,In_4680,In_1152);
nand U4836 (N_4836,In_3800,In_1923);
and U4837 (N_4837,In_2209,In_3034);
nand U4838 (N_4838,In_390,In_1408);
or U4839 (N_4839,In_3768,In_3634);
or U4840 (N_4840,In_2905,In_4337);
or U4841 (N_4841,In_1348,In_4582);
xnor U4842 (N_4842,In_4,In_4521);
nor U4843 (N_4843,In_206,In_3344);
nand U4844 (N_4844,In_3449,In_3710);
nand U4845 (N_4845,In_297,In_1349);
or U4846 (N_4846,In_2669,In_4826);
nand U4847 (N_4847,In_1755,In_2623);
nand U4848 (N_4848,In_2995,In_2074);
or U4849 (N_4849,In_3074,In_4536);
or U4850 (N_4850,In_3719,In_3469);
nor U4851 (N_4851,In_387,In_909);
nand U4852 (N_4852,In_1811,In_4694);
and U4853 (N_4853,In_4698,In_1585);
nor U4854 (N_4854,In_1805,In_3836);
or U4855 (N_4855,In_3900,In_1782);
nand U4856 (N_4856,In_2201,In_894);
nor U4857 (N_4857,In_371,In_4101);
nor U4858 (N_4858,In_3179,In_3310);
or U4859 (N_4859,In_2287,In_4789);
or U4860 (N_4860,In_4271,In_4149);
nand U4861 (N_4861,In_3539,In_4004);
xnor U4862 (N_4862,In_3700,In_4416);
nor U4863 (N_4863,In_4149,In_4721);
or U4864 (N_4864,In_128,In_2657);
nor U4865 (N_4865,In_3066,In_3517);
nor U4866 (N_4866,In_2219,In_3011);
or U4867 (N_4867,In_3831,In_3626);
or U4868 (N_4868,In_2176,In_3654);
nand U4869 (N_4869,In_2351,In_218);
and U4870 (N_4870,In_4163,In_3161);
or U4871 (N_4871,In_4736,In_1436);
or U4872 (N_4872,In_223,In_909);
and U4873 (N_4873,In_770,In_1816);
and U4874 (N_4874,In_1998,In_2769);
nor U4875 (N_4875,In_1179,In_3008);
nor U4876 (N_4876,In_2319,In_160);
and U4877 (N_4877,In_4617,In_3472);
or U4878 (N_4878,In_4426,In_4389);
nor U4879 (N_4879,In_1740,In_3683);
and U4880 (N_4880,In_4318,In_823);
and U4881 (N_4881,In_671,In_1117);
nor U4882 (N_4882,In_3101,In_598);
nand U4883 (N_4883,In_2499,In_190);
and U4884 (N_4884,In_2374,In_2901);
and U4885 (N_4885,In_1363,In_933);
or U4886 (N_4886,In_4829,In_265);
or U4887 (N_4887,In_853,In_3051);
and U4888 (N_4888,In_4097,In_1518);
and U4889 (N_4889,In_1384,In_3873);
and U4890 (N_4890,In_1096,In_4779);
or U4891 (N_4891,In_3,In_2409);
or U4892 (N_4892,In_333,In_416);
nand U4893 (N_4893,In_89,In_3856);
xnor U4894 (N_4894,In_2844,In_2406);
or U4895 (N_4895,In_3374,In_2425);
and U4896 (N_4896,In_4547,In_2197);
or U4897 (N_4897,In_4194,In_723);
nor U4898 (N_4898,In_1429,In_4432);
nand U4899 (N_4899,In_3679,In_2758);
or U4900 (N_4900,In_3442,In_2403);
or U4901 (N_4901,In_3231,In_3746);
nor U4902 (N_4902,In_4849,In_2924);
or U4903 (N_4903,In_1232,In_4293);
or U4904 (N_4904,In_740,In_2956);
nand U4905 (N_4905,In_3573,In_3616);
nand U4906 (N_4906,In_1777,In_2932);
and U4907 (N_4907,In_1739,In_569);
nand U4908 (N_4908,In_1952,In_2047);
or U4909 (N_4909,In_4415,In_2275);
nor U4910 (N_4910,In_2970,In_4946);
nand U4911 (N_4911,In_4477,In_282);
nand U4912 (N_4912,In_4365,In_2181);
nor U4913 (N_4913,In_138,In_3216);
and U4914 (N_4914,In_4979,In_4563);
or U4915 (N_4915,In_1230,In_3130);
nand U4916 (N_4916,In_1949,In_2778);
xor U4917 (N_4917,In_1786,In_2588);
nand U4918 (N_4918,In_83,In_4598);
nor U4919 (N_4919,In_1714,In_556);
nor U4920 (N_4920,In_3619,In_2680);
xnor U4921 (N_4921,In_4392,In_1107);
or U4922 (N_4922,In_2389,In_4455);
nand U4923 (N_4923,In_4258,In_421);
nor U4924 (N_4924,In_3061,In_3804);
nor U4925 (N_4925,In_393,In_4689);
and U4926 (N_4926,In_3074,In_1218);
nor U4927 (N_4927,In_4941,In_2584);
or U4928 (N_4928,In_1732,In_3815);
nand U4929 (N_4929,In_4896,In_1550);
or U4930 (N_4930,In_1678,In_1759);
and U4931 (N_4931,In_2158,In_2371);
nand U4932 (N_4932,In_2284,In_2399);
or U4933 (N_4933,In_2557,In_275);
nand U4934 (N_4934,In_4277,In_196);
nor U4935 (N_4935,In_772,In_2466);
nand U4936 (N_4936,In_4233,In_1804);
nand U4937 (N_4937,In_3077,In_2839);
nand U4938 (N_4938,In_266,In_4746);
nor U4939 (N_4939,In_1704,In_107);
nor U4940 (N_4940,In_3491,In_4165);
and U4941 (N_4941,In_2182,In_858);
or U4942 (N_4942,In_2776,In_694);
xor U4943 (N_4943,In_3286,In_4919);
and U4944 (N_4944,In_187,In_2954);
or U4945 (N_4945,In_3239,In_1998);
or U4946 (N_4946,In_4696,In_1739);
or U4947 (N_4947,In_64,In_3886);
nor U4948 (N_4948,In_1361,In_3425);
or U4949 (N_4949,In_3371,In_2166);
and U4950 (N_4950,In_1031,In_4875);
nand U4951 (N_4951,In_3216,In_2655);
nor U4952 (N_4952,In_3990,In_763);
nand U4953 (N_4953,In_2479,In_3750);
and U4954 (N_4954,In_1536,In_2403);
and U4955 (N_4955,In_4289,In_2497);
and U4956 (N_4956,In_1306,In_4986);
nor U4957 (N_4957,In_2005,In_4918);
and U4958 (N_4958,In_3816,In_4778);
nor U4959 (N_4959,In_3044,In_70);
and U4960 (N_4960,In_2473,In_3923);
nand U4961 (N_4961,In_4119,In_1667);
xor U4962 (N_4962,In_901,In_2861);
and U4963 (N_4963,In_4713,In_3475);
xor U4964 (N_4964,In_4010,In_2204);
nor U4965 (N_4965,In_592,In_4020);
nor U4966 (N_4966,In_4146,In_2349);
and U4967 (N_4967,In_4616,In_518);
and U4968 (N_4968,In_4387,In_3899);
nand U4969 (N_4969,In_859,In_2640);
and U4970 (N_4970,In_4900,In_1312);
and U4971 (N_4971,In_4071,In_464);
or U4972 (N_4972,In_4451,In_3480);
nand U4973 (N_4973,In_3134,In_1903);
or U4974 (N_4974,In_4978,In_1185);
nor U4975 (N_4975,In_4135,In_2673);
nand U4976 (N_4976,In_263,In_4149);
nand U4977 (N_4977,In_3541,In_2050);
xor U4978 (N_4978,In_1709,In_2605);
or U4979 (N_4979,In_973,In_581);
or U4980 (N_4980,In_4187,In_3730);
nor U4981 (N_4981,In_2407,In_602);
or U4982 (N_4982,In_3459,In_3138);
or U4983 (N_4983,In_2981,In_3026);
nand U4984 (N_4984,In_325,In_2911);
or U4985 (N_4985,In_4896,In_1159);
and U4986 (N_4986,In_994,In_866);
or U4987 (N_4987,In_716,In_1747);
nor U4988 (N_4988,In_4576,In_2199);
and U4989 (N_4989,In_4875,In_4284);
or U4990 (N_4990,In_711,In_1716);
nor U4991 (N_4991,In_1221,In_4585);
and U4992 (N_4992,In_756,In_3018);
or U4993 (N_4993,In_2860,In_2245);
nand U4994 (N_4994,In_2984,In_292);
nand U4995 (N_4995,In_332,In_2743);
or U4996 (N_4996,In_395,In_4368);
and U4997 (N_4997,In_3571,In_3859);
and U4998 (N_4998,In_3893,In_4105);
or U4999 (N_4999,In_998,In_1575);
and U5000 (N_5000,In_3,In_2969);
nand U5001 (N_5001,In_1984,In_3174);
nor U5002 (N_5002,In_127,In_3005);
nor U5003 (N_5003,In_1889,In_1789);
xnor U5004 (N_5004,In_1245,In_1614);
or U5005 (N_5005,In_1752,In_353);
and U5006 (N_5006,In_4405,In_3478);
xnor U5007 (N_5007,In_2538,In_4869);
nand U5008 (N_5008,In_3250,In_1709);
xnor U5009 (N_5009,In_1166,In_2568);
nand U5010 (N_5010,In_3735,In_1507);
or U5011 (N_5011,In_2739,In_2871);
and U5012 (N_5012,In_4058,In_4464);
or U5013 (N_5013,In_2290,In_234);
or U5014 (N_5014,In_4738,In_3711);
nor U5015 (N_5015,In_2869,In_796);
nor U5016 (N_5016,In_1499,In_4538);
and U5017 (N_5017,In_4553,In_1516);
nor U5018 (N_5018,In_2428,In_3445);
or U5019 (N_5019,In_3992,In_3310);
or U5020 (N_5020,In_3723,In_1844);
or U5021 (N_5021,In_4490,In_219);
and U5022 (N_5022,In_1946,In_381);
xor U5023 (N_5023,In_3716,In_1596);
nor U5024 (N_5024,In_3199,In_2608);
and U5025 (N_5025,In_370,In_767);
and U5026 (N_5026,In_3443,In_2741);
nand U5027 (N_5027,In_3966,In_3063);
or U5028 (N_5028,In_3380,In_1368);
and U5029 (N_5029,In_2311,In_583);
nand U5030 (N_5030,In_4534,In_4764);
and U5031 (N_5031,In_2748,In_1335);
and U5032 (N_5032,In_4020,In_66);
nand U5033 (N_5033,In_287,In_2766);
xnor U5034 (N_5034,In_4780,In_3058);
or U5035 (N_5035,In_3333,In_3877);
nor U5036 (N_5036,In_3301,In_75);
nand U5037 (N_5037,In_2202,In_2124);
or U5038 (N_5038,In_198,In_2310);
nand U5039 (N_5039,In_4239,In_2025);
nor U5040 (N_5040,In_923,In_3863);
nor U5041 (N_5041,In_1072,In_3239);
nor U5042 (N_5042,In_1965,In_1296);
nor U5043 (N_5043,In_4193,In_3957);
nand U5044 (N_5044,In_3450,In_2133);
xnor U5045 (N_5045,In_149,In_2892);
and U5046 (N_5046,In_4994,In_1487);
nor U5047 (N_5047,In_3910,In_111);
nor U5048 (N_5048,In_291,In_818);
and U5049 (N_5049,In_4044,In_2696);
nor U5050 (N_5050,In_1355,In_3866);
nor U5051 (N_5051,In_2158,In_4211);
or U5052 (N_5052,In_844,In_4441);
nor U5053 (N_5053,In_4117,In_3384);
or U5054 (N_5054,In_4746,In_2758);
nand U5055 (N_5055,In_3387,In_116);
nand U5056 (N_5056,In_2460,In_3432);
nand U5057 (N_5057,In_3547,In_4033);
nand U5058 (N_5058,In_1540,In_968);
nand U5059 (N_5059,In_2827,In_1108);
nand U5060 (N_5060,In_1734,In_5);
nand U5061 (N_5061,In_2010,In_3066);
nor U5062 (N_5062,In_4334,In_2274);
and U5063 (N_5063,In_4317,In_2878);
nand U5064 (N_5064,In_1400,In_2119);
xnor U5065 (N_5065,In_1165,In_3736);
nor U5066 (N_5066,In_2250,In_96);
nor U5067 (N_5067,In_1584,In_2643);
or U5068 (N_5068,In_1843,In_1778);
or U5069 (N_5069,In_916,In_2880);
and U5070 (N_5070,In_1141,In_1761);
and U5071 (N_5071,In_2584,In_4113);
nor U5072 (N_5072,In_3662,In_1602);
and U5073 (N_5073,In_4987,In_2417);
and U5074 (N_5074,In_4961,In_1444);
nor U5075 (N_5075,In_4794,In_1776);
and U5076 (N_5076,In_1121,In_422);
nand U5077 (N_5077,In_4282,In_1531);
xnor U5078 (N_5078,In_4903,In_1310);
nand U5079 (N_5079,In_4884,In_552);
nand U5080 (N_5080,In_3576,In_3061);
or U5081 (N_5081,In_1520,In_2387);
nand U5082 (N_5082,In_428,In_259);
xor U5083 (N_5083,In_4403,In_4576);
nor U5084 (N_5084,In_1531,In_3485);
and U5085 (N_5085,In_4769,In_4283);
nor U5086 (N_5086,In_3586,In_2216);
and U5087 (N_5087,In_191,In_3159);
nand U5088 (N_5088,In_1804,In_3007);
or U5089 (N_5089,In_4877,In_1414);
nand U5090 (N_5090,In_3649,In_997);
and U5091 (N_5091,In_4618,In_3153);
and U5092 (N_5092,In_3828,In_383);
nor U5093 (N_5093,In_3634,In_2200);
or U5094 (N_5094,In_3679,In_916);
and U5095 (N_5095,In_2174,In_3928);
or U5096 (N_5096,In_1605,In_4294);
nand U5097 (N_5097,In_288,In_2674);
and U5098 (N_5098,In_1879,In_1553);
nand U5099 (N_5099,In_536,In_3771);
or U5100 (N_5100,In_4957,In_4201);
xnor U5101 (N_5101,In_3493,In_2412);
nor U5102 (N_5102,In_2691,In_2464);
and U5103 (N_5103,In_1423,In_986);
nand U5104 (N_5104,In_1984,In_4611);
xnor U5105 (N_5105,In_4455,In_3789);
nand U5106 (N_5106,In_3923,In_2076);
nor U5107 (N_5107,In_2717,In_2891);
and U5108 (N_5108,In_1690,In_833);
xnor U5109 (N_5109,In_3490,In_80);
nor U5110 (N_5110,In_3211,In_2991);
nor U5111 (N_5111,In_2105,In_4795);
xor U5112 (N_5112,In_4495,In_2026);
and U5113 (N_5113,In_1662,In_3128);
and U5114 (N_5114,In_1730,In_4116);
xnor U5115 (N_5115,In_3929,In_4749);
and U5116 (N_5116,In_4728,In_1839);
or U5117 (N_5117,In_2542,In_1732);
or U5118 (N_5118,In_1462,In_1752);
nand U5119 (N_5119,In_3989,In_1998);
nand U5120 (N_5120,In_388,In_4890);
or U5121 (N_5121,In_4737,In_2996);
and U5122 (N_5122,In_3518,In_4662);
nand U5123 (N_5123,In_4915,In_1848);
nor U5124 (N_5124,In_4456,In_1809);
nand U5125 (N_5125,In_2984,In_3735);
or U5126 (N_5126,In_2123,In_3756);
nor U5127 (N_5127,In_1866,In_2274);
and U5128 (N_5128,In_400,In_4498);
and U5129 (N_5129,In_4180,In_4859);
and U5130 (N_5130,In_3783,In_959);
xor U5131 (N_5131,In_3853,In_1955);
nor U5132 (N_5132,In_4121,In_4502);
nand U5133 (N_5133,In_3993,In_3986);
nor U5134 (N_5134,In_3976,In_720);
nor U5135 (N_5135,In_3122,In_2031);
nor U5136 (N_5136,In_2692,In_2232);
or U5137 (N_5137,In_4026,In_1373);
or U5138 (N_5138,In_3862,In_1189);
nor U5139 (N_5139,In_2038,In_4373);
nand U5140 (N_5140,In_4064,In_2376);
or U5141 (N_5141,In_1747,In_3448);
or U5142 (N_5142,In_486,In_3566);
nor U5143 (N_5143,In_1664,In_760);
nor U5144 (N_5144,In_1736,In_3687);
and U5145 (N_5145,In_4762,In_3342);
or U5146 (N_5146,In_1287,In_2405);
xnor U5147 (N_5147,In_3692,In_4756);
nor U5148 (N_5148,In_4322,In_597);
and U5149 (N_5149,In_2288,In_4520);
or U5150 (N_5150,In_4321,In_531);
nand U5151 (N_5151,In_4654,In_2745);
and U5152 (N_5152,In_2118,In_183);
nand U5153 (N_5153,In_4740,In_2306);
and U5154 (N_5154,In_1520,In_3346);
and U5155 (N_5155,In_2689,In_4118);
nand U5156 (N_5156,In_3581,In_4827);
nor U5157 (N_5157,In_3014,In_442);
nor U5158 (N_5158,In_3928,In_2507);
nand U5159 (N_5159,In_16,In_2440);
and U5160 (N_5160,In_3607,In_1137);
or U5161 (N_5161,In_1237,In_3477);
nor U5162 (N_5162,In_3425,In_3137);
or U5163 (N_5163,In_4620,In_2358);
nand U5164 (N_5164,In_3257,In_706);
nand U5165 (N_5165,In_1120,In_408);
and U5166 (N_5166,In_556,In_326);
nand U5167 (N_5167,In_2480,In_2705);
nand U5168 (N_5168,In_249,In_1013);
or U5169 (N_5169,In_4034,In_4713);
nand U5170 (N_5170,In_2515,In_3486);
or U5171 (N_5171,In_1825,In_4683);
and U5172 (N_5172,In_4885,In_2298);
nor U5173 (N_5173,In_564,In_123);
and U5174 (N_5174,In_2495,In_4402);
nor U5175 (N_5175,In_67,In_483);
or U5176 (N_5176,In_458,In_684);
and U5177 (N_5177,In_2427,In_454);
nand U5178 (N_5178,In_3780,In_4399);
xnor U5179 (N_5179,In_3194,In_1981);
and U5180 (N_5180,In_4706,In_1068);
or U5181 (N_5181,In_2521,In_4849);
or U5182 (N_5182,In_1729,In_1129);
and U5183 (N_5183,In_1610,In_4787);
or U5184 (N_5184,In_905,In_3140);
nor U5185 (N_5185,In_4401,In_1192);
nand U5186 (N_5186,In_1174,In_707);
nor U5187 (N_5187,In_3337,In_160);
xor U5188 (N_5188,In_4170,In_408);
nor U5189 (N_5189,In_1272,In_3552);
or U5190 (N_5190,In_1645,In_3497);
nor U5191 (N_5191,In_357,In_2133);
and U5192 (N_5192,In_2187,In_1314);
or U5193 (N_5193,In_2142,In_3665);
nor U5194 (N_5194,In_2888,In_2989);
or U5195 (N_5195,In_3162,In_2235);
xnor U5196 (N_5196,In_3768,In_2701);
xor U5197 (N_5197,In_3345,In_2155);
and U5198 (N_5198,In_1513,In_3149);
or U5199 (N_5199,In_304,In_2366);
and U5200 (N_5200,In_4066,In_1928);
xor U5201 (N_5201,In_172,In_4505);
xor U5202 (N_5202,In_3530,In_962);
nand U5203 (N_5203,In_4851,In_2156);
or U5204 (N_5204,In_3333,In_3181);
and U5205 (N_5205,In_4551,In_226);
and U5206 (N_5206,In_1243,In_1823);
nand U5207 (N_5207,In_2933,In_4134);
nor U5208 (N_5208,In_3096,In_3068);
or U5209 (N_5209,In_1689,In_4992);
nand U5210 (N_5210,In_546,In_1833);
nand U5211 (N_5211,In_3011,In_890);
nor U5212 (N_5212,In_1682,In_1545);
or U5213 (N_5213,In_2482,In_817);
nand U5214 (N_5214,In_3872,In_2181);
nand U5215 (N_5215,In_1424,In_860);
or U5216 (N_5216,In_596,In_4453);
and U5217 (N_5217,In_1227,In_744);
nor U5218 (N_5218,In_4228,In_3606);
or U5219 (N_5219,In_4143,In_1573);
xor U5220 (N_5220,In_818,In_2524);
nand U5221 (N_5221,In_1068,In_1897);
nand U5222 (N_5222,In_4231,In_785);
and U5223 (N_5223,In_398,In_1966);
xnor U5224 (N_5224,In_3100,In_3954);
nand U5225 (N_5225,In_4981,In_85);
nor U5226 (N_5226,In_2635,In_1252);
nor U5227 (N_5227,In_385,In_1371);
nor U5228 (N_5228,In_4571,In_4831);
xor U5229 (N_5229,In_1028,In_3059);
nor U5230 (N_5230,In_864,In_3963);
nand U5231 (N_5231,In_3899,In_1203);
and U5232 (N_5232,In_2886,In_2537);
and U5233 (N_5233,In_2828,In_3884);
nor U5234 (N_5234,In_688,In_1226);
and U5235 (N_5235,In_1046,In_4466);
and U5236 (N_5236,In_347,In_837);
or U5237 (N_5237,In_2256,In_710);
nand U5238 (N_5238,In_208,In_4954);
nand U5239 (N_5239,In_2235,In_3884);
nor U5240 (N_5240,In_1492,In_523);
nor U5241 (N_5241,In_143,In_3974);
xnor U5242 (N_5242,In_4265,In_3733);
nand U5243 (N_5243,In_1325,In_897);
nand U5244 (N_5244,In_1506,In_854);
nor U5245 (N_5245,In_2418,In_1330);
nor U5246 (N_5246,In_4631,In_1068);
or U5247 (N_5247,In_3903,In_2588);
nand U5248 (N_5248,In_542,In_2063);
and U5249 (N_5249,In_103,In_4788);
and U5250 (N_5250,In_4556,In_3684);
and U5251 (N_5251,In_3144,In_3202);
xor U5252 (N_5252,In_3076,In_3837);
nand U5253 (N_5253,In_2389,In_707);
and U5254 (N_5254,In_1087,In_3561);
nor U5255 (N_5255,In_4296,In_2058);
xor U5256 (N_5256,In_310,In_2337);
and U5257 (N_5257,In_3339,In_4540);
nand U5258 (N_5258,In_1795,In_4918);
and U5259 (N_5259,In_4823,In_352);
nand U5260 (N_5260,In_144,In_2034);
and U5261 (N_5261,In_2130,In_2387);
nand U5262 (N_5262,In_2944,In_188);
nand U5263 (N_5263,In_2356,In_3744);
nor U5264 (N_5264,In_4241,In_1333);
xor U5265 (N_5265,In_4358,In_1591);
nor U5266 (N_5266,In_2152,In_4711);
xor U5267 (N_5267,In_4933,In_805);
nor U5268 (N_5268,In_3527,In_4305);
or U5269 (N_5269,In_3644,In_3654);
xnor U5270 (N_5270,In_3991,In_2065);
or U5271 (N_5271,In_2045,In_3603);
nor U5272 (N_5272,In_4727,In_1635);
nand U5273 (N_5273,In_173,In_4929);
nand U5274 (N_5274,In_1188,In_775);
nor U5275 (N_5275,In_4243,In_1424);
and U5276 (N_5276,In_1750,In_4453);
nor U5277 (N_5277,In_2003,In_3833);
nand U5278 (N_5278,In_3544,In_4393);
and U5279 (N_5279,In_4633,In_3900);
or U5280 (N_5280,In_4346,In_3868);
nor U5281 (N_5281,In_4464,In_4832);
nor U5282 (N_5282,In_2411,In_2814);
or U5283 (N_5283,In_1278,In_938);
nand U5284 (N_5284,In_2330,In_4016);
or U5285 (N_5285,In_524,In_708);
nand U5286 (N_5286,In_173,In_3110);
and U5287 (N_5287,In_1300,In_4410);
and U5288 (N_5288,In_2409,In_852);
or U5289 (N_5289,In_904,In_2616);
or U5290 (N_5290,In_4795,In_4160);
nand U5291 (N_5291,In_1088,In_4969);
nand U5292 (N_5292,In_973,In_1917);
nand U5293 (N_5293,In_4497,In_2888);
nand U5294 (N_5294,In_2401,In_1775);
nand U5295 (N_5295,In_2358,In_2646);
nand U5296 (N_5296,In_12,In_4406);
nor U5297 (N_5297,In_2921,In_237);
xor U5298 (N_5298,In_2076,In_1997);
nor U5299 (N_5299,In_2641,In_2665);
nand U5300 (N_5300,In_4697,In_2625);
nand U5301 (N_5301,In_1181,In_2843);
nor U5302 (N_5302,In_3646,In_4036);
nand U5303 (N_5303,In_2448,In_1001);
nand U5304 (N_5304,In_1741,In_4775);
or U5305 (N_5305,In_3483,In_3477);
nor U5306 (N_5306,In_2402,In_1471);
or U5307 (N_5307,In_2419,In_3111);
and U5308 (N_5308,In_2996,In_436);
and U5309 (N_5309,In_1483,In_1625);
nor U5310 (N_5310,In_4130,In_1638);
xnor U5311 (N_5311,In_2059,In_2042);
nand U5312 (N_5312,In_3894,In_1749);
and U5313 (N_5313,In_39,In_2905);
xor U5314 (N_5314,In_1256,In_2460);
nor U5315 (N_5315,In_223,In_4915);
nand U5316 (N_5316,In_4505,In_237);
nand U5317 (N_5317,In_3426,In_34);
nor U5318 (N_5318,In_1826,In_2836);
or U5319 (N_5319,In_3917,In_4051);
nand U5320 (N_5320,In_1101,In_3135);
nor U5321 (N_5321,In_926,In_4044);
or U5322 (N_5322,In_2893,In_3600);
nor U5323 (N_5323,In_2761,In_4425);
and U5324 (N_5324,In_3853,In_1023);
nand U5325 (N_5325,In_4931,In_1388);
nand U5326 (N_5326,In_1060,In_4758);
nand U5327 (N_5327,In_4311,In_2665);
and U5328 (N_5328,In_448,In_1375);
xor U5329 (N_5329,In_1325,In_1820);
or U5330 (N_5330,In_559,In_2229);
nand U5331 (N_5331,In_4095,In_987);
or U5332 (N_5332,In_3266,In_4614);
xnor U5333 (N_5333,In_40,In_4100);
nor U5334 (N_5334,In_1625,In_1778);
nand U5335 (N_5335,In_1001,In_1142);
nor U5336 (N_5336,In_2712,In_2513);
xnor U5337 (N_5337,In_891,In_1109);
xor U5338 (N_5338,In_4400,In_2398);
nor U5339 (N_5339,In_2790,In_122);
or U5340 (N_5340,In_4409,In_1022);
nor U5341 (N_5341,In_237,In_4048);
nand U5342 (N_5342,In_4959,In_1015);
or U5343 (N_5343,In_4599,In_1613);
nand U5344 (N_5344,In_2094,In_2866);
or U5345 (N_5345,In_318,In_2045);
nand U5346 (N_5346,In_4143,In_2112);
or U5347 (N_5347,In_4827,In_4892);
nand U5348 (N_5348,In_1957,In_2069);
xnor U5349 (N_5349,In_2545,In_4162);
nor U5350 (N_5350,In_4010,In_3130);
nand U5351 (N_5351,In_2621,In_4675);
and U5352 (N_5352,In_104,In_4913);
and U5353 (N_5353,In_2155,In_4765);
nand U5354 (N_5354,In_1745,In_672);
and U5355 (N_5355,In_3986,In_3094);
nor U5356 (N_5356,In_3457,In_4140);
or U5357 (N_5357,In_1844,In_1942);
or U5358 (N_5358,In_2618,In_2107);
nand U5359 (N_5359,In_1756,In_4705);
or U5360 (N_5360,In_238,In_778);
and U5361 (N_5361,In_2985,In_3);
nand U5362 (N_5362,In_4636,In_1670);
or U5363 (N_5363,In_110,In_3684);
or U5364 (N_5364,In_4426,In_4284);
nand U5365 (N_5365,In_2930,In_4601);
or U5366 (N_5366,In_1347,In_4340);
nand U5367 (N_5367,In_1777,In_4568);
or U5368 (N_5368,In_2738,In_3141);
and U5369 (N_5369,In_2063,In_1451);
nor U5370 (N_5370,In_2783,In_136);
or U5371 (N_5371,In_2924,In_1161);
xnor U5372 (N_5372,In_1785,In_635);
nand U5373 (N_5373,In_536,In_2334);
nor U5374 (N_5374,In_774,In_755);
nor U5375 (N_5375,In_563,In_1261);
or U5376 (N_5376,In_3957,In_3117);
and U5377 (N_5377,In_2203,In_1124);
and U5378 (N_5378,In_2227,In_1994);
nand U5379 (N_5379,In_3646,In_3070);
or U5380 (N_5380,In_1366,In_680);
and U5381 (N_5381,In_4800,In_4037);
and U5382 (N_5382,In_4742,In_2733);
or U5383 (N_5383,In_3644,In_2799);
nand U5384 (N_5384,In_2477,In_4546);
nand U5385 (N_5385,In_3835,In_1605);
or U5386 (N_5386,In_2918,In_2742);
and U5387 (N_5387,In_401,In_4760);
nor U5388 (N_5388,In_1189,In_4745);
xnor U5389 (N_5389,In_2884,In_3437);
xor U5390 (N_5390,In_4298,In_2926);
and U5391 (N_5391,In_243,In_3899);
and U5392 (N_5392,In_4651,In_2365);
nor U5393 (N_5393,In_905,In_2816);
or U5394 (N_5394,In_3072,In_3570);
nand U5395 (N_5395,In_1810,In_2704);
nand U5396 (N_5396,In_2271,In_3088);
nand U5397 (N_5397,In_3566,In_3440);
and U5398 (N_5398,In_388,In_1660);
or U5399 (N_5399,In_4648,In_1080);
and U5400 (N_5400,In_1583,In_4537);
nor U5401 (N_5401,In_1802,In_4166);
nor U5402 (N_5402,In_1132,In_933);
nand U5403 (N_5403,In_2137,In_1570);
and U5404 (N_5404,In_2813,In_2732);
nor U5405 (N_5405,In_2946,In_182);
nor U5406 (N_5406,In_1300,In_4948);
nand U5407 (N_5407,In_3595,In_2786);
and U5408 (N_5408,In_168,In_2103);
nor U5409 (N_5409,In_3670,In_1002);
xnor U5410 (N_5410,In_3530,In_2238);
or U5411 (N_5411,In_3348,In_1407);
nor U5412 (N_5412,In_4645,In_4435);
and U5413 (N_5413,In_3866,In_1389);
or U5414 (N_5414,In_3795,In_3934);
nand U5415 (N_5415,In_3371,In_2375);
xor U5416 (N_5416,In_1606,In_3880);
nor U5417 (N_5417,In_432,In_4747);
nand U5418 (N_5418,In_4060,In_3948);
and U5419 (N_5419,In_1466,In_1899);
nand U5420 (N_5420,In_3043,In_3031);
nand U5421 (N_5421,In_951,In_41);
or U5422 (N_5422,In_3091,In_1671);
nor U5423 (N_5423,In_2096,In_466);
or U5424 (N_5424,In_697,In_2630);
nor U5425 (N_5425,In_1639,In_4982);
xnor U5426 (N_5426,In_2417,In_144);
nand U5427 (N_5427,In_4282,In_2544);
nand U5428 (N_5428,In_67,In_2182);
and U5429 (N_5429,In_4186,In_1163);
xor U5430 (N_5430,In_1176,In_3669);
nand U5431 (N_5431,In_997,In_3702);
nor U5432 (N_5432,In_2086,In_2207);
nor U5433 (N_5433,In_1338,In_3021);
and U5434 (N_5434,In_308,In_659);
and U5435 (N_5435,In_2699,In_50);
and U5436 (N_5436,In_1442,In_503);
nand U5437 (N_5437,In_2953,In_3799);
nand U5438 (N_5438,In_1569,In_2169);
nand U5439 (N_5439,In_4999,In_2026);
and U5440 (N_5440,In_1376,In_4940);
nand U5441 (N_5441,In_1758,In_2776);
nor U5442 (N_5442,In_4132,In_2296);
and U5443 (N_5443,In_4565,In_3608);
nor U5444 (N_5444,In_1083,In_1851);
and U5445 (N_5445,In_4237,In_3202);
or U5446 (N_5446,In_4777,In_4027);
and U5447 (N_5447,In_4515,In_2338);
xor U5448 (N_5448,In_3340,In_466);
nor U5449 (N_5449,In_1677,In_3063);
or U5450 (N_5450,In_126,In_2809);
nor U5451 (N_5451,In_1366,In_4145);
xor U5452 (N_5452,In_1139,In_1656);
or U5453 (N_5453,In_4888,In_2980);
nor U5454 (N_5454,In_2704,In_1080);
and U5455 (N_5455,In_4930,In_4846);
nand U5456 (N_5456,In_1243,In_1179);
nor U5457 (N_5457,In_1935,In_1830);
or U5458 (N_5458,In_3401,In_1763);
xnor U5459 (N_5459,In_3130,In_1794);
nand U5460 (N_5460,In_4275,In_3214);
nand U5461 (N_5461,In_417,In_4147);
nor U5462 (N_5462,In_241,In_2307);
and U5463 (N_5463,In_720,In_3547);
nor U5464 (N_5464,In_544,In_3469);
nand U5465 (N_5465,In_63,In_961);
and U5466 (N_5466,In_72,In_2213);
or U5467 (N_5467,In_2699,In_2021);
or U5468 (N_5468,In_2177,In_4761);
nor U5469 (N_5469,In_1493,In_93);
nor U5470 (N_5470,In_1242,In_1375);
nand U5471 (N_5471,In_2000,In_904);
or U5472 (N_5472,In_2789,In_670);
nand U5473 (N_5473,In_1245,In_2493);
and U5474 (N_5474,In_4577,In_4538);
nand U5475 (N_5475,In_4870,In_2878);
xor U5476 (N_5476,In_3205,In_4499);
nor U5477 (N_5477,In_3259,In_4412);
or U5478 (N_5478,In_2667,In_1671);
or U5479 (N_5479,In_157,In_3371);
nand U5480 (N_5480,In_427,In_4466);
nand U5481 (N_5481,In_4099,In_2086);
xnor U5482 (N_5482,In_452,In_2264);
and U5483 (N_5483,In_4722,In_2629);
nand U5484 (N_5484,In_1031,In_1276);
nand U5485 (N_5485,In_1573,In_2179);
nor U5486 (N_5486,In_1361,In_3480);
or U5487 (N_5487,In_2563,In_2959);
and U5488 (N_5488,In_3940,In_2994);
or U5489 (N_5489,In_1959,In_42);
and U5490 (N_5490,In_2104,In_2891);
xnor U5491 (N_5491,In_164,In_3251);
and U5492 (N_5492,In_3727,In_3102);
and U5493 (N_5493,In_1533,In_1396);
nand U5494 (N_5494,In_2484,In_2162);
and U5495 (N_5495,In_3256,In_2033);
and U5496 (N_5496,In_2151,In_1762);
and U5497 (N_5497,In_1307,In_2968);
or U5498 (N_5498,In_814,In_4781);
or U5499 (N_5499,In_3597,In_3198);
xnor U5500 (N_5500,In_2917,In_2867);
and U5501 (N_5501,In_4424,In_193);
and U5502 (N_5502,In_4785,In_4359);
nor U5503 (N_5503,In_680,In_569);
nor U5504 (N_5504,In_1425,In_2049);
nor U5505 (N_5505,In_4107,In_1393);
or U5506 (N_5506,In_3494,In_1209);
nand U5507 (N_5507,In_4222,In_3671);
xor U5508 (N_5508,In_3360,In_2999);
and U5509 (N_5509,In_111,In_4679);
and U5510 (N_5510,In_4248,In_4210);
nand U5511 (N_5511,In_889,In_1711);
and U5512 (N_5512,In_4319,In_1344);
xnor U5513 (N_5513,In_3157,In_4751);
and U5514 (N_5514,In_564,In_3937);
nand U5515 (N_5515,In_3336,In_94);
nand U5516 (N_5516,In_4126,In_658);
and U5517 (N_5517,In_154,In_1662);
nor U5518 (N_5518,In_990,In_1153);
nor U5519 (N_5519,In_2423,In_3139);
xor U5520 (N_5520,In_3308,In_4599);
nand U5521 (N_5521,In_4333,In_1693);
nor U5522 (N_5522,In_4825,In_906);
nand U5523 (N_5523,In_3046,In_3001);
nand U5524 (N_5524,In_2457,In_4926);
xnor U5525 (N_5525,In_1988,In_3857);
nor U5526 (N_5526,In_2104,In_32);
and U5527 (N_5527,In_1750,In_488);
or U5528 (N_5528,In_1854,In_705);
or U5529 (N_5529,In_2467,In_2229);
or U5530 (N_5530,In_788,In_517);
nand U5531 (N_5531,In_4536,In_3063);
nor U5532 (N_5532,In_4027,In_3566);
and U5533 (N_5533,In_2017,In_3151);
or U5534 (N_5534,In_2961,In_3396);
and U5535 (N_5535,In_3488,In_4900);
or U5536 (N_5536,In_4958,In_3530);
nor U5537 (N_5537,In_4156,In_4740);
nor U5538 (N_5538,In_1791,In_1321);
nand U5539 (N_5539,In_46,In_2542);
or U5540 (N_5540,In_247,In_4031);
nor U5541 (N_5541,In_2007,In_3152);
or U5542 (N_5542,In_2942,In_1029);
nor U5543 (N_5543,In_3690,In_582);
or U5544 (N_5544,In_3771,In_1945);
and U5545 (N_5545,In_4595,In_4314);
xnor U5546 (N_5546,In_3810,In_3701);
and U5547 (N_5547,In_372,In_2781);
and U5548 (N_5548,In_3019,In_205);
and U5549 (N_5549,In_3288,In_2738);
or U5550 (N_5550,In_1690,In_1439);
xor U5551 (N_5551,In_1805,In_88);
nor U5552 (N_5552,In_2435,In_4529);
and U5553 (N_5553,In_1887,In_2153);
nand U5554 (N_5554,In_1482,In_2475);
nand U5555 (N_5555,In_3904,In_2313);
and U5556 (N_5556,In_2032,In_3066);
nor U5557 (N_5557,In_256,In_1542);
or U5558 (N_5558,In_2670,In_4656);
and U5559 (N_5559,In_1416,In_4763);
and U5560 (N_5560,In_928,In_1029);
nor U5561 (N_5561,In_1847,In_3879);
nand U5562 (N_5562,In_3657,In_247);
nor U5563 (N_5563,In_3466,In_2630);
nor U5564 (N_5564,In_1772,In_3142);
and U5565 (N_5565,In_4851,In_3628);
nand U5566 (N_5566,In_2051,In_4391);
xnor U5567 (N_5567,In_1441,In_2108);
nor U5568 (N_5568,In_4426,In_550);
nand U5569 (N_5569,In_1016,In_2028);
nand U5570 (N_5570,In_1581,In_4039);
and U5571 (N_5571,In_718,In_3239);
xor U5572 (N_5572,In_1347,In_2735);
nor U5573 (N_5573,In_1280,In_30);
or U5574 (N_5574,In_2929,In_643);
nand U5575 (N_5575,In_3639,In_1507);
nor U5576 (N_5576,In_4347,In_699);
nand U5577 (N_5577,In_413,In_3768);
nand U5578 (N_5578,In_128,In_2361);
and U5579 (N_5579,In_699,In_1512);
and U5580 (N_5580,In_2538,In_680);
nor U5581 (N_5581,In_2983,In_3956);
or U5582 (N_5582,In_544,In_4484);
or U5583 (N_5583,In_4328,In_3602);
and U5584 (N_5584,In_4383,In_1703);
nand U5585 (N_5585,In_4952,In_3126);
or U5586 (N_5586,In_1031,In_234);
nand U5587 (N_5587,In_4757,In_2467);
and U5588 (N_5588,In_2339,In_990);
and U5589 (N_5589,In_880,In_2290);
or U5590 (N_5590,In_2393,In_1722);
and U5591 (N_5591,In_1692,In_4118);
or U5592 (N_5592,In_4350,In_3313);
and U5593 (N_5593,In_4547,In_362);
and U5594 (N_5594,In_54,In_3279);
nand U5595 (N_5595,In_1390,In_4915);
nand U5596 (N_5596,In_1574,In_3887);
and U5597 (N_5597,In_3200,In_476);
nand U5598 (N_5598,In_2783,In_4092);
nand U5599 (N_5599,In_1467,In_2264);
and U5600 (N_5600,In_4275,In_2746);
or U5601 (N_5601,In_1392,In_267);
or U5602 (N_5602,In_4208,In_859);
nor U5603 (N_5603,In_629,In_1205);
nand U5604 (N_5604,In_1710,In_2683);
nand U5605 (N_5605,In_2237,In_1039);
or U5606 (N_5606,In_2913,In_1760);
nor U5607 (N_5607,In_4217,In_4131);
and U5608 (N_5608,In_2301,In_4730);
nor U5609 (N_5609,In_1776,In_3892);
nand U5610 (N_5610,In_2503,In_714);
and U5611 (N_5611,In_82,In_4074);
nor U5612 (N_5612,In_3692,In_1498);
xor U5613 (N_5613,In_2810,In_2200);
xnor U5614 (N_5614,In_123,In_1603);
nor U5615 (N_5615,In_3501,In_1845);
and U5616 (N_5616,In_3853,In_4257);
nor U5617 (N_5617,In_3300,In_4087);
or U5618 (N_5618,In_1708,In_2517);
nor U5619 (N_5619,In_2230,In_2081);
xor U5620 (N_5620,In_4984,In_3718);
nor U5621 (N_5621,In_3311,In_4662);
or U5622 (N_5622,In_1003,In_3572);
and U5623 (N_5623,In_13,In_4420);
or U5624 (N_5624,In_2360,In_2068);
nand U5625 (N_5625,In_1404,In_2065);
nor U5626 (N_5626,In_3758,In_4914);
and U5627 (N_5627,In_3704,In_2685);
nand U5628 (N_5628,In_3811,In_2502);
nand U5629 (N_5629,In_749,In_3708);
nor U5630 (N_5630,In_1991,In_2881);
nand U5631 (N_5631,In_3359,In_4690);
xor U5632 (N_5632,In_1876,In_471);
nand U5633 (N_5633,In_1974,In_237);
or U5634 (N_5634,In_4457,In_1261);
nand U5635 (N_5635,In_3533,In_3687);
nand U5636 (N_5636,In_4884,In_4592);
or U5637 (N_5637,In_2852,In_3159);
or U5638 (N_5638,In_4671,In_3803);
nand U5639 (N_5639,In_755,In_942);
nand U5640 (N_5640,In_3282,In_2274);
nor U5641 (N_5641,In_2766,In_2967);
nand U5642 (N_5642,In_4242,In_233);
nand U5643 (N_5643,In_2836,In_1255);
or U5644 (N_5644,In_3000,In_510);
or U5645 (N_5645,In_4566,In_3330);
and U5646 (N_5646,In_4804,In_751);
nor U5647 (N_5647,In_1097,In_2380);
and U5648 (N_5648,In_3761,In_4674);
and U5649 (N_5649,In_4473,In_3235);
nand U5650 (N_5650,In_3835,In_742);
and U5651 (N_5651,In_329,In_343);
or U5652 (N_5652,In_4103,In_3630);
xnor U5653 (N_5653,In_1498,In_4264);
or U5654 (N_5654,In_2692,In_2710);
nor U5655 (N_5655,In_1975,In_3559);
xor U5656 (N_5656,In_954,In_591);
nor U5657 (N_5657,In_4054,In_2798);
nor U5658 (N_5658,In_2104,In_2369);
xnor U5659 (N_5659,In_2544,In_1575);
and U5660 (N_5660,In_4677,In_3906);
or U5661 (N_5661,In_2153,In_1645);
or U5662 (N_5662,In_4873,In_2654);
or U5663 (N_5663,In_1894,In_1885);
and U5664 (N_5664,In_2948,In_4447);
nor U5665 (N_5665,In_4680,In_18);
nor U5666 (N_5666,In_1851,In_2000);
or U5667 (N_5667,In_706,In_800);
and U5668 (N_5668,In_2540,In_1237);
xnor U5669 (N_5669,In_1457,In_4967);
nand U5670 (N_5670,In_1942,In_1833);
nand U5671 (N_5671,In_3013,In_2157);
and U5672 (N_5672,In_3316,In_3679);
and U5673 (N_5673,In_2297,In_3855);
xnor U5674 (N_5674,In_4198,In_455);
xor U5675 (N_5675,In_1278,In_4333);
or U5676 (N_5676,In_3404,In_308);
nor U5677 (N_5677,In_450,In_2104);
and U5678 (N_5678,In_960,In_3082);
and U5679 (N_5679,In_4220,In_94);
and U5680 (N_5680,In_2271,In_4233);
nor U5681 (N_5681,In_2634,In_407);
and U5682 (N_5682,In_2068,In_386);
or U5683 (N_5683,In_4005,In_1976);
nor U5684 (N_5684,In_4883,In_1616);
and U5685 (N_5685,In_1255,In_2922);
nor U5686 (N_5686,In_1480,In_2524);
nand U5687 (N_5687,In_4678,In_3291);
or U5688 (N_5688,In_4166,In_4914);
nand U5689 (N_5689,In_2291,In_4703);
and U5690 (N_5690,In_582,In_212);
nand U5691 (N_5691,In_1987,In_639);
and U5692 (N_5692,In_3877,In_2498);
and U5693 (N_5693,In_4461,In_1567);
nand U5694 (N_5694,In_2520,In_4552);
and U5695 (N_5695,In_3431,In_4254);
nand U5696 (N_5696,In_3789,In_3596);
nor U5697 (N_5697,In_1693,In_955);
nor U5698 (N_5698,In_4334,In_4729);
nor U5699 (N_5699,In_2380,In_3965);
and U5700 (N_5700,In_2624,In_3535);
xnor U5701 (N_5701,In_1768,In_2649);
or U5702 (N_5702,In_52,In_3405);
and U5703 (N_5703,In_934,In_544);
and U5704 (N_5704,In_4327,In_3896);
nand U5705 (N_5705,In_736,In_3890);
nand U5706 (N_5706,In_1265,In_742);
nand U5707 (N_5707,In_687,In_2175);
nor U5708 (N_5708,In_771,In_4547);
nor U5709 (N_5709,In_2367,In_2038);
nor U5710 (N_5710,In_742,In_2020);
or U5711 (N_5711,In_744,In_496);
or U5712 (N_5712,In_1588,In_4154);
nand U5713 (N_5713,In_1609,In_4552);
nor U5714 (N_5714,In_4287,In_4212);
nor U5715 (N_5715,In_515,In_3844);
and U5716 (N_5716,In_3777,In_4666);
and U5717 (N_5717,In_1399,In_4371);
nor U5718 (N_5718,In_2447,In_1623);
xor U5719 (N_5719,In_990,In_1417);
or U5720 (N_5720,In_2282,In_3688);
xor U5721 (N_5721,In_3539,In_4954);
nand U5722 (N_5722,In_3002,In_3709);
nand U5723 (N_5723,In_4151,In_3256);
nand U5724 (N_5724,In_3225,In_1860);
nand U5725 (N_5725,In_758,In_830);
and U5726 (N_5726,In_2824,In_3547);
and U5727 (N_5727,In_4936,In_3992);
nand U5728 (N_5728,In_2618,In_132);
nor U5729 (N_5729,In_2277,In_328);
nand U5730 (N_5730,In_883,In_4889);
nor U5731 (N_5731,In_82,In_4251);
nor U5732 (N_5732,In_2773,In_3053);
and U5733 (N_5733,In_3368,In_1054);
and U5734 (N_5734,In_2096,In_1834);
nand U5735 (N_5735,In_692,In_3355);
and U5736 (N_5736,In_3179,In_2301);
xor U5737 (N_5737,In_257,In_4395);
nor U5738 (N_5738,In_1571,In_281);
and U5739 (N_5739,In_3999,In_1085);
or U5740 (N_5740,In_1865,In_4372);
nand U5741 (N_5741,In_1688,In_4222);
xnor U5742 (N_5742,In_2472,In_4942);
nand U5743 (N_5743,In_2581,In_4245);
and U5744 (N_5744,In_3764,In_4260);
xnor U5745 (N_5745,In_1249,In_1345);
nor U5746 (N_5746,In_3334,In_4508);
and U5747 (N_5747,In_1566,In_1731);
or U5748 (N_5748,In_623,In_4000);
nor U5749 (N_5749,In_256,In_885);
nand U5750 (N_5750,In_1294,In_1524);
nor U5751 (N_5751,In_4162,In_3384);
or U5752 (N_5752,In_1173,In_2455);
and U5753 (N_5753,In_871,In_374);
nand U5754 (N_5754,In_2241,In_3865);
nor U5755 (N_5755,In_2854,In_3241);
nand U5756 (N_5756,In_2428,In_4048);
nand U5757 (N_5757,In_2979,In_1299);
and U5758 (N_5758,In_1713,In_1627);
xnor U5759 (N_5759,In_24,In_1759);
xor U5760 (N_5760,In_1364,In_1854);
or U5761 (N_5761,In_2631,In_1386);
or U5762 (N_5762,In_597,In_1294);
nand U5763 (N_5763,In_809,In_4122);
xnor U5764 (N_5764,In_1720,In_1844);
and U5765 (N_5765,In_2044,In_3810);
nand U5766 (N_5766,In_3967,In_1870);
nand U5767 (N_5767,In_1061,In_3561);
and U5768 (N_5768,In_4488,In_1615);
and U5769 (N_5769,In_1758,In_2999);
xnor U5770 (N_5770,In_3556,In_2353);
nand U5771 (N_5771,In_4958,In_36);
nand U5772 (N_5772,In_4058,In_2154);
or U5773 (N_5773,In_4206,In_3054);
nor U5774 (N_5774,In_2990,In_3729);
nand U5775 (N_5775,In_4539,In_3398);
and U5776 (N_5776,In_4518,In_2265);
xor U5777 (N_5777,In_3716,In_143);
nor U5778 (N_5778,In_4729,In_2474);
nand U5779 (N_5779,In_811,In_1030);
nor U5780 (N_5780,In_3418,In_1031);
or U5781 (N_5781,In_4842,In_2256);
and U5782 (N_5782,In_3674,In_4479);
and U5783 (N_5783,In_4469,In_2365);
nand U5784 (N_5784,In_49,In_4126);
xnor U5785 (N_5785,In_293,In_4484);
nor U5786 (N_5786,In_1326,In_3917);
nand U5787 (N_5787,In_4478,In_413);
and U5788 (N_5788,In_421,In_1924);
nor U5789 (N_5789,In_2725,In_263);
nor U5790 (N_5790,In_3439,In_1874);
xnor U5791 (N_5791,In_3418,In_1299);
nor U5792 (N_5792,In_890,In_4790);
xor U5793 (N_5793,In_1026,In_4437);
nor U5794 (N_5794,In_1041,In_1884);
nand U5795 (N_5795,In_2844,In_2588);
nand U5796 (N_5796,In_2204,In_278);
nor U5797 (N_5797,In_2202,In_1844);
or U5798 (N_5798,In_2391,In_3338);
xnor U5799 (N_5799,In_3481,In_3087);
and U5800 (N_5800,In_4668,In_2268);
xnor U5801 (N_5801,In_3742,In_767);
or U5802 (N_5802,In_3657,In_2904);
nand U5803 (N_5803,In_3494,In_3332);
nor U5804 (N_5804,In_1961,In_2252);
nand U5805 (N_5805,In_164,In_4537);
and U5806 (N_5806,In_4209,In_3999);
and U5807 (N_5807,In_1308,In_1210);
and U5808 (N_5808,In_2396,In_3431);
nor U5809 (N_5809,In_4951,In_2006);
nand U5810 (N_5810,In_527,In_2470);
or U5811 (N_5811,In_1556,In_2774);
nand U5812 (N_5812,In_3857,In_4943);
and U5813 (N_5813,In_102,In_3711);
and U5814 (N_5814,In_4994,In_4788);
nor U5815 (N_5815,In_574,In_524);
or U5816 (N_5816,In_4900,In_3363);
or U5817 (N_5817,In_2662,In_2343);
and U5818 (N_5818,In_2302,In_2989);
or U5819 (N_5819,In_1249,In_3561);
nand U5820 (N_5820,In_4481,In_3112);
or U5821 (N_5821,In_3041,In_626);
nand U5822 (N_5822,In_4789,In_4953);
and U5823 (N_5823,In_3405,In_1414);
xor U5824 (N_5824,In_2795,In_1986);
nand U5825 (N_5825,In_582,In_363);
or U5826 (N_5826,In_2007,In_2012);
nand U5827 (N_5827,In_4648,In_648);
nand U5828 (N_5828,In_4201,In_3805);
nand U5829 (N_5829,In_2888,In_2587);
nor U5830 (N_5830,In_4928,In_2330);
and U5831 (N_5831,In_266,In_4511);
and U5832 (N_5832,In_829,In_403);
or U5833 (N_5833,In_3082,In_1138);
and U5834 (N_5834,In_4594,In_3813);
and U5835 (N_5835,In_3762,In_1861);
or U5836 (N_5836,In_1409,In_3768);
or U5837 (N_5837,In_3347,In_658);
or U5838 (N_5838,In_4803,In_4631);
nand U5839 (N_5839,In_2506,In_516);
nor U5840 (N_5840,In_3589,In_891);
nand U5841 (N_5841,In_2295,In_4918);
or U5842 (N_5842,In_244,In_4829);
and U5843 (N_5843,In_1408,In_2263);
or U5844 (N_5844,In_2733,In_4022);
or U5845 (N_5845,In_3655,In_1993);
or U5846 (N_5846,In_3855,In_2442);
or U5847 (N_5847,In_3625,In_379);
and U5848 (N_5848,In_3223,In_3371);
and U5849 (N_5849,In_249,In_2548);
nor U5850 (N_5850,In_4216,In_3890);
xnor U5851 (N_5851,In_3100,In_241);
and U5852 (N_5852,In_2907,In_4186);
xor U5853 (N_5853,In_4872,In_2394);
or U5854 (N_5854,In_4876,In_2701);
nor U5855 (N_5855,In_1715,In_1626);
xor U5856 (N_5856,In_1086,In_4942);
and U5857 (N_5857,In_3666,In_4545);
nor U5858 (N_5858,In_444,In_4904);
nor U5859 (N_5859,In_3319,In_319);
nand U5860 (N_5860,In_1833,In_3401);
and U5861 (N_5861,In_3327,In_2745);
or U5862 (N_5862,In_3499,In_3456);
or U5863 (N_5863,In_2695,In_4300);
or U5864 (N_5864,In_887,In_3467);
xor U5865 (N_5865,In_562,In_4526);
or U5866 (N_5866,In_2064,In_3773);
and U5867 (N_5867,In_221,In_3388);
or U5868 (N_5868,In_3011,In_1894);
nor U5869 (N_5869,In_3193,In_4626);
nor U5870 (N_5870,In_491,In_2110);
xor U5871 (N_5871,In_309,In_3693);
xor U5872 (N_5872,In_3920,In_447);
or U5873 (N_5873,In_4968,In_3971);
or U5874 (N_5874,In_4806,In_3734);
or U5875 (N_5875,In_2754,In_362);
nor U5876 (N_5876,In_3537,In_3284);
nand U5877 (N_5877,In_4848,In_2247);
nand U5878 (N_5878,In_3947,In_4524);
and U5879 (N_5879,In_3786,In_1375);
and U5880 (N_5880,In_2794,In_3533);
nor U5881 (N_5881,In_3006,In_3186);
nand U5882 (N_5882,In_1767,In_3997);
and U5883 (N_5883,In_3386,In_1620);
nor U5884 (N_5884,In_342,In_2221);
nand U5885 (N_5885,In_935,In_1329);
nor U5886 (N_5886,In_3262,In_265);
or U5887 (N_5887,In_1992,In_3751);
and U5888 (N_5888,In_3437,In_4974);
and U5889 (N_5889,In_4899,In_3117);
nand U5890 (N_5890,In_4016,In_2891);
or U5891 (N_5891,In_2738,In_950);
nand U5892 (N_5892,In_187,In_3050);
xnor U5893 (N_5893,In_2082,In_4354);
or U5894 (N_5894,In_2473,In_2803);
nand U5895 (N_5895,In_4391,In_4619);
nor U5896 (N_5896,In_1248,In_721);
nor U5897 (N_5897,In_2307,In_1811);
and U5898 (N_5898,In_56,In_1993);
or U5899 (N_5899,In_1912,In_4389);
nand U5900 (N_5900,In_3358,In_1542);
nor U5901 (N_5901,In_17,In_748);
nand U5902 (N_5902,In_4873,In_133);
or U5903 (N_5903,In_1405,In_945);
and U5904 (N_5904,In_3683,In_2767);
and U5905 (N_5905,In_373,In_981);
nor U5906 (N_5906,In_1298,In_2294);
and U5907 (N_5907,In_1128,In_921);
or U5908 (N_5908,In_1471,In_2672);
and U5909 (N_5909,In_2548,In_4554);
and U5910 (N_5910,In_526,In_4076);
and U5911 (N_5911,In_4631,In_2320);
nand U5912 (N_5912,In_185,In_557);
nand U5913 (N_5913,In_3714,In_1927);
nand U5914 (N_5914,In_3435,In_852);
nand U5915 (N_5915,In_2381,In_1056);
or U5916 (N_5916,In_2767,In_4132);
and U5917 (N_5917,In_2282,In_3428);
and U5918 (N_5918,In_3940,In_3994);
nand U5919 (N_5919,In_4759,In_2830);
and U5920 (N_5920,In_102,In_2017);
xnor U5921 (N_5921,In_2867,In_4760);
and U5922 (N_5922,In_2879,In_350);
nand U5923 (N_5923,In_4011,In_714);
nor U5924 (N_5924,In_3816,In_2043);
nor U5925 (N_5925,In_2425,In_4209);
and U5926 (N_5926,In_2265,In_3662);
or U5927 (N_5927,In_4163,In_4159);
nand U5928 (N_5928,In_4018,In_1746);
and U5929 (N_5929,In_134,In_2962);
and U5930 (N_5930,In_3585,In_1739);
nor U5931 (N_5931,In_1143,In_4930);
nor U5932 (N_5932,In_2460,In_3311);
nor U5933 (N_5933,In_3523,In_2955);
nor U5934 (N_5934,In_2270,In_4792);
nor U5935 (N_5935,In_2052,In_3374);
nor U5936 (N_5936,In_1693,In_633);
xnor U5937 (N_5937,In_1995,In_4472);
and U5938 (N_5938,In_2686,In_4968);
and U5939 (N_5939,In_2053,In_446);
or U5940 (N_5940,In_1844,In_3448);
and U5941 (N_5941,In_3664,In_4732);
nand U5942 (N_5942,In_2585,In_3299);
or U5943 (N_5943,In_1109,In_4311);
or U5944 (N_5944,In_2588,In_3971);
nor U5945 (N_5945,In_2691,In_3418);
or U5946 (N_5946,In_4101,In_2377);
nor U5947 (N_5947,In_1091,In_91);
nand U5948 (N_5948,In_1072,In_3559);
and U5949 (N_5949,In_780,In_4858);
and U5950 (N_5950,In_4119,In_2035);
nor U5951 (N_5951,In_1346,In_3284);
or U5952 (N_5952,In_2345,In_4534);
xnor U5953 (N_5953,In_2713,In_550);
nand U5954 (N_5954,In_1176,In_4670);
nand U5955 (N_5955,In_2789,In_4320);
and U5956 (N_5956,In_3985,In_4804);
nor U5957 (N_5957,In_4250,In_4706);
and U5958 (N_5958,In_830,In_3374);
xnor U5959 (N_5959,In_3947,In_1242);
and U5960 (N_5960,In_1636,In_3459);
or U5961 (N_5961,In_4251,In_708);
and U5962 (N_5962,In_592,In_382);
xor U5963 (N_5963,In_2530,In_253);
nor U5964 (N_5964,In_2877,In_1574);
nand U5965 (N_5965,In_51,In_2310);
nor U5966 (N_5966,In_1840,In_2681);
and U5967 (N_5967,In_1695,In_4144);
or U5968 (N_5968,In_4271,In_1399);
and U5969 (N_5969,In_4440,In_679);
or U5970 (N_5970,In_18,In_1400);
or U5971 (N_5971,In_4005,In_4353);
and U5972 (N_5972,In_395,In_1985);
nand U5973 (N_5973,In_771,In_3624);
nor U5974 (N_5974,In_2714,In_3157);
and U5975 (N_5975,In_2868,In_2882);
or U5976 (N_5976,In_4169,In_585);
or U5977 (N_5977,In_4317,In_4704);
and U5978 (N_5978,In_2267,In_3916);
nand U5979 (N_5979,In_3536,In_4777);
or U5980 (N_5980,In_2980,In_191);
nand U5981 (N_5981,In_4025,In_2604);
xor U5982 (N_5982,In_1679,In_4565);
and U5983 (N_5983,In_1077,In_701);
or U5984 (N_5984,In_354,In_1125);
nor U5985 (N_5985,In_2607,In_2724);
nand U5986 (N_5986,In_2258,In_426);
nand U5987 (N_5987,In_4933,In_3364);
xnor U5988 (N_5988,In_574,In_1262);
xor U5989 (N_5989,In_2521,In_2641);
xor U5990 (N_5990,In_2516,In_2617);
and U5991 (N_5991,In_1534,In_2264);
nor U5992 (N_5992,In_4443,In_3947);
and U5993 (N_5993,In_41,In_2987);
or U5994 (N_5994,In_1995,In_740);
nand U5995 (N_5995,In_3678,In_57);
or U5996 (N_5996,In_2262,In_1591);
xor U5997 (N_5997,In_2191,In_8);
nand U5998 (N_5998,In_4819,In_372);
xor U5999 (N_5999,In_4849,In_3542);
or U6000 (N_6000,In_3364,In_1905);
and U6001 (N_6001,In_2313,In_6);
or U6002 (N_6002,In_1260,In_3012);
nand U6003 (N_6003,In_4050,In_3438);
and U6004 (N_6004,In_1850,In_59);
nand U6005 (N_6005,In_605,In_468);
or U6006 (N_6006,In_1106,In_1415);
or U6007 (N_6007,In_4123,In_3714);
and U6008 (N_6008,In_2297,In_3156);
xnor U6009 (N_6009,In_2318,In_1101);
nand U6010 (N_6010,In_2795,In_2420);
or U6011 (N_6011,In_2967,In_4227);
and U6012 (N_6012,In_1014,In_4148);
or U6013 (N_6013,In_4955,In_531);
or U6014 (N_6014,In_3950,In_4121);
or U6015 (N_6015,In_4036,In_3719);
nand U6016 (N_6016,In_547,In_2323);
nor U6017 (N_6017,In_2986,In_4045);
nand U6018 (N_6018,In_1119,In_3986);
and U6019 (N_6019,In_3765,In_2500);
nand U6020 (N_6020,In_1616,In_4352);
and U6021 (N_6021,In_2607,In_3913);
and U6022 (N_6022,In_1060,In_1981);
nand U6023 (N_6023,In_212,In_1646);
xor U6024 (N_6024,In_874,In_3325);
or U6025 (N_6025,In_3084,In_265);
and U6026 (N_6026,In_4671,In_3849);
or U6027 (N_6027,In_2811,In_2616);
and U6028 (N_6028,In_3483,In_2696);
nor U6029 (N_6029,In_472,In_2157);
nand U6030 (N_6030,In_1370,In_2045);
nor U6031 (N_6031,In_1171,In_3445);
nand U6032 (N_6032,In_2678,In_127);
and U6033 (N_6033,In_4628,In_3438);
nand U6034 (N_6034,In_1664,In_1966);
xor U6035 (N_6035,In_2879,In_1122);
or U6036 (N_6036,In_3211,In_4312);
and U6037 (N_6037,In_4056,In_2933);
nor U6038 (N_6038,In_2906,In_368);
nor U6039 (N_6039,In_1317,In_1380);
nor U6040 (N_6040,In_4316,In_114);
or U6041 (N_6041,In_1843,In_3691);
nor U6042 (N_6042,In_3900,In_2450);
and U6043 (N_6043,In_3571,In_478);
nor U6044 (N_6044,In_248,In_2257);
or U6045 (N_6045,In_142,In_3069);
nor U6046 (N_6046,In_4293,In_3047);
nand U6047 (N_6047,In_3021,In_1029);
and U6048 (N_6048,In_3184,In_1296);
nand U6049 (N_6049,In_4154,In_2027);
and U6050 (N_6050,In_980,In_4839);
nand U6051 (N_6051,In_3377,In_3079);
nor U6052 (N_6052,In_1436,In_2200);
nor U6053 (N_6053,In_2413,In_3286);
nand U6054 (N_6054,In_2638,In_2071);
nand U6055 (N_6055,In_1208,In_1538);
nand U6056 (N_6056,In_4482,In_802);
and U6057 (N_6057,In_612,In_1868);
nor U6058 (N_6058,In_588,In_4016);
nand U6059 (N_6059,In_1145,In_4912);
nand U6060 (N_6060,In_525,In_2428);
and U6061 (N_6061,In_3858,In_1352);
and U6062 (N_6062,In_621,In_2212);
nand U6063 (N_6063,In_4801,In_3556);
and U6064 (N_6064,In_3944,In_4085);
nor U6065 (N_6065,In_4516,In_4839);
and U6066 (N_6066,In_288,In_3863);
nand U6067 (N_6067,In_804,In_1554);
or U6068 (N_6068,In_4279,In_2334);
nor U6069 (N_6069,In_1527,In_4430);
nand U6070 (N_6070,In_2295,In_1373);
or U6071 (N_6071,In_227,In_4445);
and U6072 (N_6072,In_1081,In_3629);
nor U6073 (N_6073,In_276,In_3616);
nor U6074 (N_6074,In_279,In_2575);
or U6075 (N_6075,In_4657,In_1581);
and U6076 (N_6076,In_3338,In_4879);
nor U6077 (N_6077,In_170,In_190);
and U6078 (N_6078,In_739,In_4253);
nand U6079 (N_6079,In_947,In_3471);
nand U6080 (N_6080,In_31,In_2943);
and U6081 (N_6081,In_124,In_3463);
nand U6082 (N_6082,In_4444,In_264);
nand U6083 (N_6083,In_3975,In_3628);
or U6084 (N_6084,In_559,In_4175);
nor U6085 (N_6085,In_4013,In_2730);
and U6086 (N_6086,In_135,In_3679);
or U6087 (N_6087,In_973,In_3222);
nor U6088 (N_6088,In_174,In_2858);
nand U6089 (N_6089,In_1119,In_2930);
nor U6090 (N_6090,In_4476,In_2565);
nor U6091 (N_6091,In_132,In_4955);
nor U6092 (N_6092,In_3713,In_4337);
nor U6093 (N_6093,In_4060,In_1421);
nor U6094 (N_6094,In_2202,In_2237);
or U6095 (N_6095,In_321,In_1517);
nor U6096 (N_6096,In_489,In_1242);
nand U6097 (N_6097,In_3959,In_1150);
nand U6098 (N_6098,In_1292,In_2208);
and U6099 (N_6099,In_549,In_4250);
or U6100 (N_6100,In_4210,In_534);
nor U6101 (N_6101,In_2163,In_500);
nor U6102 (N_6102,In_2423,In_4940);
xnor U6103 (N_6103,In_2594,In_4643);
or U6104 (N_6104,In_2274,In_4768);
and U6105 (N_6105,In_1838,In_3090);
nor U6106 (N_6106,In_825,In_1841);
or U6107 (N_6107,In_3838,In_2569);
and U6108 (N_6108,In_979,In_4558);
xnor U6109 (N_6109,In_2414,In_2886);
and U6110 (N_6110,In_3524,In_2227);
nor U6111 (N_6111,In_1348,In_262);
or U6112 (N_6112,In_2954,In_3977);
and U6113 (N_6113,In_74,In_4648);
nor U6114 (N_6114,In_2904,In_265);
or U6115 (N_6115,In_1622,In_3126);
and U6116 (N_6116,In_3023,In_2299);
nand U6117 (N_6117,In_3922,In_3875);
nor U6118 (N_6118,In_1480,In_3256);
nand U6119 (N_6119,In_1265,In_2045);
and U6120 (N_6120,In_594,In_1140);
or U6121 (N_6121,In_4051,In_1210);
or U6122 (N_6122,In_1086,In_1940);
nor U6123 (N_6123,In_1655,In_2045);
xnor U6124 (N_6124,In_4379,In_2328);
and U6125 (N_6125,In_4977,In_3307);
nand U6126 (N_6126,In_2409,In_511);
or U6127 (N_6127,In_2089,In_2141);
and U6128 (N_6128,In_1424,In_483);
nand U6129 (N_6129,In_1366,In_595);
nand U6130 (N_6130,In_1698,In_2515);
nand U6131 (N_6131,In_2696,In_3248);
nor U6132 (N_6132,In_2099,In_610);
nor U6133 (N_6133,In_2868,In_439);
nor U6134 (N_6134,In_1901,In_1669);
or U6135 (N_6135,In_988,In_2482);
nor U6136 (N_6136,In_2225,In_4049);
nand U6137 (N_6137,In_2286,In_4951);
nor U6138 (N_6138,In_2948,In_1737);
nor U6139 (N_6139,In_557,In_2031);
nor U6140 (N_6140,In_1853,In_1894);
nand U6141 (N_6141,In_3268,In_1335);
and U6142 (N_6142,In_421,In_3699);
nor U6143 (N_6143,In_1073,In_719);
xor U6144 (N_6144,In_4928,In_4370);
or U6145 (N_6145,In_4831,In_1892);
nand U6146 (N_6146,In_4398,In_1764);
and U6147 (N_6147,In_2549,In_235);
nor U6148 (N_6148,In_4938,In_3428);
nand U6149 (N_6149,In_2235,In_210);
xor U6150 (N_6150,In_254,In_1070);
or U6151 (N_6151,In_4164,In_346);
or U6152 (N_6152,In_4368,In_1259);
nand U6153 (N_6153,In_4210,In_387);
and U6154 (N_6154,In_779,In_4423);
nor U6155 (N_6155,In_1335,In_2117);
nor U6156 (N_6156,In_1631,In_4603);
and U6157 (N_6157,In_2468,In_168);
nor U6158 (N_6158,In_3231,In_3119);
xnor U6159 (N_6159,In_982,In_961);
nor U6160 (N_6160,In_3964,In_619);
nand U6161 (N_6161,In_4791,In_440);
nor U6162 (N_6162,In_4962,In_4363);
and U6163 (N_6163,In_56,In_4408);
xnor U6164 (N_6164,In_3700,In_2940);
xnor U6165 (N_6165,In_417,In_1316);
nand U6166 (N_6166,In_3349,In_842);
nor U6167 (N_6167,In_3167,In_2787);
or U6168 (N_6168,In_3762,In_2130);
nor U6169 (N_6169,In_1239,In_3430);
or U6170 (N_6170,In_1674,In_1172);
or U6171 (N_6171,In_1185,In_3049);
and U6172 (N_6172,In_2002,In_2210);
and U6173 (N_6173,In_1583,In_4542);
and U6174 (N_6174,In_2490,In_4974);
nand U6175 (N_6175,In_44,In_2392);
nor U6176 (N_6176,In_3521,In_34);
or U6177 (N_6177,In_819,In_1655);
nand U6178 (N_6178,In_4936,In_4321);
or U6179 (N_6179,In_4942,In_3160);
or U6180 (N_6180,In_4421,In_2257);
or U6181 (N_6181,In_1352,In_2723);
nor U6182 (N_6182,In_2001,In_1117);
nand U6183 (N_6183,In_811,In_1306);
nor U6184 (N_6184,In_326,In_3320);
nand U6185 (N_6185,In_3548,In_4254);
and U6186 (N_6186,In_1075,In_746);
nor U6187 (N_6187,In_4343,In_760);
and U6188 (N_6188,In_317,In_4295);
or U6189 (N_6189,In_3279,In_2524);
nor U6190 (N_6190,In_4986,In_2723);
nor U6191 (N_6191,In_4199,In_2473);
or U6192 (N_6192,In_3811,In_3830);
nor U6193 (N_6193,In_3035,In_4806);
or U6194 (N_6194,In_775,In_1627);
nor U6195 (N_6195,In_4395,In_1095);
xor U6196 (N_6196,In_1091,In_524);
nor U6197 (N_6197,In_2053,In_4908);
xor U6198 (N_6198,In_2421,In_4071);
and U6199 (N_6199,In_4808,In_1345);
and U6200 (N_6200,In_3674,In_4126);
xnor U6201 (N_6201,In_476,In_247);
or U6202 (N_6202,In_4745,In_4269);
nand U6203 (N_6203,In_4250,In_1088);
nand U6204 (N_6204,In_1565,In_3357);
or U6205 (N_6205,In_4716,In_806);
or U6206 (N_6206,In_1488,In_221);
and U6207 (N_6207,In_3274,In_1812);
xnor U6208 (N_6208,In_2359,In_4783);
nor U6209 (N_6209,In_1509,In_2952);
nand U6210 (N_6210,In_303,In_3256);
nor U6211 (N_6211,In_1454,In_4183);
nand U6212 (N_6212,In_3356,In_1602);
nand U6213 (N_6213,In_2707,In_960);
nand U6214 (N_6214,In_864,In_164);
and U6215 (N_6215,In_3456,In_3054);
or U6216 (N_6216,In_2187,In_1573);
or U6217 (N_6217,In_2742,In_3032);
and U6218 (N_6218,In_1645,In_4052);
or U6219 (N_6219,In_765,In_4994);
and U6220 (N_6220,In_3805,In_2980);
nand U6221 (N_6221,In_3796,In_3736);
nor U6222 (N_6222,In_4801,In_3028);
or U6223 (N_6223,In_3372,In_4011);
nor U6224 (N_6224,In_2832,In_2911);
and U6225 (N_6225,In_3142,In_3857);
xor U6226 (N_6226,In_25,In_240);
and U6227 (N_6227,In_906,In_824);
nor U6228 (N_6228,In_4106,In_3812);
and U6229 (N_6229,In_2512,In_571);
and U6230 (N_6230,In_2468,In_1450);
or U6231 (N_6231,In_3752,In_3546);
xor U6232 (N_6232,In_2332,In_848);
or U6233 (N_6233,In_3301,In_4231);
or U6234 (N_6234,In_631,In_3368);
or U6235 (N_6235,In_1979,In_699);
nor U6236 (N_6236,In_893,In_869);
nand U6237 (N_6237,In_2623,In_2092);
nand U6238 (N_6238,In_2145,In_163);
and U6239 (N_6239,In_1459,In_4637);
nand U6240 (N_6240,In_498,In_982);
and U6241 (N_6241,In_3938,In_4729);
nand U6242 (N_6242,In_2153,In_1885);
nand U6243 (N_6243,In_1075,In_3193);
and U6244 (N_6244,In_1408,In_1473);
and U6245 (N_6245,In_110,In_754);
nor U6246 (N_6246,In_3565,In_4574);
xor U6247 (N_6247,In_4820,In_4278);
and U6248 (N_6248,In_4032,In_3592);
nand U6249 (N_6249,In_2311,In_3570);
nand U6250 (N_6250,In_2034,In_2798);
and U6251 (N_6251,In_4295,In_2122);
nor U6252 (N_6252,In_2001,In_1135);
xor U6253 (N_6253,In_2130,In_3602);
nor U6254 (N_6254,In_1433,In_4020);
and U6255 (N_6255,In_4908,In_2655);
nor U6256 (N_6256,In_3891,In_4149);
nand U6257 (N_6257,In_3486,In_907);
nand U6258 (N_6258,In_416,In_287);
nor U6259 (N_6259,In_4686,In_4629);
xnor U6260 (N_6260,In_319,In_4917);
xnor U6261 (N_6261,In_2150,In_4394);
or U6262 (N_6262,In_1008,In_3873);
nand U6263 (N_6263,In_2774,In_2225);
and U6264 (N_6264,In_3355,In_1865);
nor U6265 (N_6265,In_1225,In_1954);
xnor U6266 (N_6266,In_3589,In_3362);
or U6267 (N_6267,In_4634,In_278);
xor U6268 (N_6268,In_4055,In_4109);
nand U6269 (N_6269,In_1835,In_2840);
and U6270 (N_6270,In_2947,In_3524);
or U6271 (N_6271,In_1896,In_160);
xor U6272 (N_6272,In_1348,In_2686);
nor U6273 (N_6273,In_350,In_1486);
nor U6274 (N_6274,In_1670,In_2826);
nor U6275 (N_6275,In_68,In_2657);
and U6276 (N_6276,In_3400,In_3933);
nand U6277 (N_6277,In_3085,In_2508);
and U6278 (N_6278,In_1636,In_1568);
or U6279 (N_6279,In_1064,In_3917);
nand U6280 (N_6280,In_4913,In_2627);
xnor U6281 (N_6281,In_2926,In_1340);
nand U6282 (N_6282,In_2766,In_112);
or U6283 (N_6283,In_4784,In_2469);
nor U6284 (N_6284,In_4281,In_655);
or U6285 (N_6285,In_3655,In_1660);
and U6286 (N_6286,In_188,In_663);
or U6287 (N_6287,In_1018,In_2481);
or U6288 (N_6288,In_19,In_683);
nand U6289 (N_6289,In_1535,In_2622);
nor U6290 (N_6290,In_3428,In_2226);
nor U6291 (N_6291,In_1709,In_4854);
or U6292 (N_6292,In_2826,In_862);
nand U6293 (N_6293,In_2355,In_688);
and U6294 (N_6294,In_3586,In_4698);
or U6295 (N_6295,In_316,In_3406);
or U6296 (N_6296,In_3907,In_454);
nor U6297 (N_6297,In_4867,In_1351);
or U6298 (N_6298,In_1643,In_1680);
nand U6299 (N_6299,In_3527,In_3517);
or U6300 (N_6300,In_4041,In_3893);
nand U6301 (N_6301,In_2266,In_2893);
nand U6302 (N_6302,In_2683,In_1065);
xor U6303 (N_6303,In_4877,In_3633);
and U6304 (N_6304,In_1215,In_4057);
nand U6305 (N_6305,In_4090,In_2313);
nand U6306 (N_6306,In_820,In_3341);
or U6307 (N_6307,In_1857,In_4591);
and U6308 (N_6308,In_1674,In_4298);
nand U6309 (N_6309,In_282,In_750);
and U6310 (N_6310,In_1134,In_2024);
or U6311 (N_6311,In_2586,In_2904);
nand U6312 (N_6312,In_4412,In_667);
and U6313 (N_6313,In_4080,In_4610);
nor U6314 (N_6314,In_4698,In_909);
nor U6315 (N_6315,In_4423,In_1465);
or U6316 (N_6316,In_1655,In_4641);
nand U6317 (N_6317,In_714,In_4737);
nor U6318 (N_6318,In_2368,In_474);
nor U6319 (N_6319,In_640,In_990);
or U6320 (N_6320,In_4125,In_729);
xor U6321 (N_6321,In_3122,In_1915);
nor U6322 (N_6322,In_1320,In_2778);
or U6323 (N_6323,In_71,In_3048);
and U6324 (N_6324,In_3778,In_1179);
nor U6325 (N_6325,In_2083,In_4322);
nand U6326 (N_6326,In_4256,In_1589);
or U6327 (N_6327,In_191,In_3752);
and U6328 (N_6328,In_2149,In_537);
xor U6329 (N_6329,In_3778,In_4342);
or U6330 (N_6330,In_1342,In_3200);
or U6331 (N_6331,In_963,In_911);
xnor U6332 (N_6332,In_1173,In_1843);
and U6333 (N_6333,In_1365,In_2302);
and U6334 (N_6334,In_1172,In_3190);
or U6335 (N_6335,In_4547,In_3976);
and U6336 (N_6336,In_1820,In_3864);
or U6337 (N_6337,In_2164,In_4314);
nand U6338 (N_6338,In_1561,In_2744);
or U6339 (N_6339,In_3621,In_4866);
nand U6340 (N_6340,In_4620,In_4096);
nor U6341 (N_6341,In_2008,In_1273);
and U6342 (N_6342,In_2961,In_777);
xnor U6343 (N_6343,In_8,In_2800);
nand U6344 (N_6344,In_1642,In_4791);
nor U6345 (N_6345,In_2595,In_1232);
nor U6346 (N_6346,In_4129,In_3743);
and U6347 (N_6347,In_122,In_3624);
xnor U6348 (N_6348,In_295,In_463);
or U6349 (N_6349,In_638,In_4605);
and U6350 (N_6350,In_1868,In_1918);
nand U6351 (N_6351,In_1075,In_4079);
and U6352 (N_6352,In_3587,In_3311);
nand U6353 (N_6353,In_1697,In_593);
nand U6354 (N_6354,In_4482,In_3675);
or U6355 (N_6355,In_1084,In_2366);
or U6356 (N_6356,In_4661,In_2592);
nand U6357 (N_6357,In_4109,In_360);
and U6358 (N_6358,In_3633,In_1033);
or U6359 (N_6359,In_1854,In_328);
or U6360 (N_6360,In_3080,In_1788);
nor U6361 (N_6361,In_733,In_1107);
and U6362 (N_6362,In_663,In_911);
or U6363 (N_6363,In_4474,In_4381);
and U6364 (N_6364,In_2111,In_1420);
nor U6365 (N_6365,In_4244,In_4634);
nor U6366 (N_6366,In_18,In_3796);
or U6367 (N_6367,In_159,In_648);
nor U6368 (N_6368,In_4064,In_607);
xnor U6369 (N_6369,In_3293,In_1435);
nor U6370 (N_6370,In_1991,In_4304);
nor U6371 (N_6371,In_1645,In_1053);
nor U6372 (N_6372,In_2080,In_3686);
and U6373 (N_6373,In_3921,In_2478);
and U6374 (N_6374,In_2903,In_2183);
and U6375 (N_6375,In_4998,In_1612);
or U6376 (N_6376,In_1630,In_1753);
nor U6377 (N_6377,In_672,In_4253);
and U6378 (N_6378,In_3430,In_1412);
xnor U6379 (N_6379,In_3301,In_1394);
nand U6380 (N_6380,In_1401,In_2805);
and U6381 (N_6381,In_4388,In_4695);
or U6382 (N_6382,In_4892,In_2227);
or U6383 (N_6383,In_101,In_1092);
or U6384 (N_6384,In_3127,In_2439);
xor U6385 (N_6385,In_1753,In_2497);
xor U6386 (N_6386,In_4464,In_4297);
nor U6387 (N_6387,In_4170,In_1851);
nand U6388 (N_6388,In_4547,In_201);
nor U6389 (N_6389,In_4822,In_2704);
nor U6390 (N_6390,In_3170,In_3953);
and U6391 (N_6391,In_1773,In_4054);
nor U6392 (N_6392,In_3089,In_3213);
nor U6393 (N_6393,In_2018,In_517);
nand U6394 (N_6394,In_4377,In_384);
nand U6395 (N_6395,In_2356,In_181);
or U6396 (N_6396,In_1223,In_1625);
nand U6397 (N_6397,In_4825,In_2791);
or U6398 (N_6398,In_4744,In_969);
nor U6399 (N_6399,In_4981,In_4040);
nor U6400 (N_6400,In_4971,In_599);
xnor U6401 (N_6401,In_889,In_4236);
and U6402 (N_6402,In_218,In_2794);
xor U6403 (N_6403,In_3752,In_681);
or U6404 (N_6404,In_3010,In_4405);
nand U6405 (N_6405,In_4585,In_4269);
or U6406 (N_6406,In_4165,In_3872);
nor U6407 (N_6407,In_864,In_914);
nand U6408 (N_6408,In_3456,In_4302);
nor U6409 (N_6409,In_2588,In_1738);
and U6410 (N_6410,In_3701,In_4819);
nand U6411 (N_6411,In_1990,In_607);
and U6412 (N_6412,In_4375,In_1752);
and U6413 (N_6413,In_4244,In_66);
and U6414 (N_6414,In_3708,In_3120);
or U6415 (N_6415,In_1908,In_3930);
nand U6416 (N_6416,In_9,In_3130);
or U6417 (N_6417,In_2514,In_3226);
nor U6418 (N_6418,In_3167,In_1819);
xnor U6419 (N_6419,In_4963,In_4613);
nor U6420 (N_6420,In_4300,In_4488);
or U6421 (N_6421,In_3225,In_2999);
and U6422 (N_6422,In_2292,In_2583);
nor U6423 (N_6423,In_1802,In_1557);
or U6424 (N_6424,In_2463,In_1490);
and U6425 (N_6425,In_4695,In_4325);
or U6426 (N_6426,In_3494,In_400);
nor U6427 (N_6427,In_1761,In_3373);
nand U6428 (N_6428,In_2164,In_2513);
nand U6429 (N_6429,In_4173,In_1144);
or U6430 (N_6430,In_2893,In_3406);
and U6431 (N_6431,In_2842,In_2692);
and U6432 (N_6432,In_2887,In_2640);
nand U6433 (N_6433,In_3372,In_3852);
nand U6434 (N_6434,In_976,In_1612);
and U6435 (N_6435,In_1835,In_2802);
nand U6436 (N_6436,In_3445,In_4434);
and U6437 (N_6437,In_2068,In_3436);
nand U6438 (N_6438,In_4549,In_1268);
and U6439 (N_6439,In_3664,In_1629);
or U6440 (N_6440,In_1886,In_1472);
or U6441 (N_6441,In_4294,In_4345);
and U6442 (N_6442,In_4678,In_3071);
or U6443 (N_6443,In_1856,In_3979);
and U6444 (N_6444,In_3081,In_3197);
nor U6445 (N_6445,In_2833,In_1497);
nand U6446 (N_6446,In_3398,In_307);
and U6447 (N_6447,In_1467,In_1058);
nor U6448 (N_6448,In_4784,In_3719);
or U6449 (N_6449,In_3194,In_98);
nor U6450 (N_6450,In_3118,In_3473);
xnor U6451 (N_6451,In_1611,In_3018);
nand U6452 (N_6452,In_733,In_1643);
and U6453 (N_6453,In_2329,In_4632);
nor U6454 (N_6454,In_2477,In_1282);
and U6455 (N_6455,In_700,In_4494);
or U6456 (N_6456,In_3341,In_2335);
nand U6457 (N_6457,In_1523,In_747);
or U6458 (N_6458,In_2706,In_3595);
or U6459 (N_6459,In_2532,In_4242);
nand U6460 (N_6460,In_4344,In_3718);
and U6461 (N_6461,In_218,In_3472);
nand U6462 (N_6462,In_3969,In_2594);
or U6463 (N_6463,In_851,In_882);
nand U6464 (N_6464,In_422,In_2152);
and U6465 (N_6465,In_4955,In_3391);
or U6466 (N_6466,In_4622,In_1922);
nand U6467 (N_6467,In_3016,In_3323);
nor U6468 (N_6468,In_643,In_2328);
nand U6469 (N_6469,In_2885,In_3775);
nor U6470 (N_6470,In_2757,In_2928);
nand U6471 (N_6471,In_2101,In_4558);
nand U6472 (N_6472,In_4294,In_4310);
xor U6473 (N_6473,In_395,In_2269);
nand U6474 (N_6474,In_3785,In_4903);
or U6475 (N_6475,In_4766,In_4974);
nand U6476 (N_6476,In_1917,In_3362);
nor U6477 (N_6477,In_2926,In_4750);
and U6478 (N_6478,In_3411,In_2732);
and U6479 (N_6479,In_3072,In_3778);
nor U6480 (N_6480,In_3033,In_3247);
nor U6481 (N_6481,In_1887,In_1738);
nor U6482 (N_6482,In_1196,In_2329);
or U6483 (N_6483,In_258,In_2251);
nor U6484 (N_6484,In_3794,In_1624);
or U6485 (N_6485,In_3488,In_3912);
nor U6486 (N_6486,In_1667,In_458);
nand U6487 (N_6487,In_2681,In_1354);
or U6488 (N_6488,In_4236,In_1424);
or U6489 (N_6489,In_3800,In_3572);
nor U6490 (N_6490,In_746,In_1382);
nand U6491 (N_6491,In_2022,In_2531);
and U6492 (N_6492,In_2323,In_3376);
and U6493 (N_6493,In_772,In_2163);
nor U6494 (N_6494,In_1735,In_2162);
nor U6495 (N_6495,In_127,In_3380);
or U6496 (N_6496,In_4319,In_3021);
xor U6497 (N_6497,In_183,In_2621);
and U6498 (N_6498,In_1899,In_2267);
or U6499 (N_6499,In_1222,In_1642);
and U6500 (N_6500,In_1221,In_3428);
nand U6501 (N_6501,In_1506,In_1024);
or U6502 (N_6502,In_2573,In_2608);
xor U6503 (N_6503,In_3314,In_894);
and U6504 (N_6504,In_2336,In_3100);
and U6505 (N_6505,In_3736,In_966);
nand U6506 (N_6506,In_8,In_1431);
or U6507 (N_6507,In_1125,In_3822);
nor U6508 (N_6508,In_1728,In_1987);
and U6509 (N_6509,In_3085,In_4465);
and U6510 (N_6510,In_3453,In_4695);
nand U6511 (N_6511,In_4526,In_2283);
nand U6512 (N_6512,In_4348,In_3873);
nor U6513 (N_6513,In_198,In_964);
nor U6514 (N_6514,In_1855,In_1620);
nor U6515 (N_6515,In_920,In_2103);
xnor U6516 (N_6516,In_228,In_3665);
or U6517 (N_6517,In_3985,In_3961);
and U6518 (N_6518,In_1714,In_4841);
xnor U6519 (N_6519,In_1262,In_3837);
nand U6520 (N_6520,In_1802,In_2241);
nor U6521 (N_6521,In_2598,In_4875);
and U6522 (N_6522,In_3882,In_516);
and U6523 (N_6523,In_2107,In_1990);
xnor U6524 (N_6524,In_3984,In_2380);
or U6525 (N_6525,In_4757,In_4068);
or U6526 (N_6526,In_2169,In_642);
nor U6527 (N_6527,In_1181,In_4554);
nor U6528 (N_6528,In_89,In_101);
or U6529 (N_6529,In_2147,In_3187);
and U6530 (N_6530,In_3351,In_1641);
nand U6531 (N_6531,In_12,In_4342);
nor U6532 (N_6532,In_4530,In_1085);
and U6533 (N_6533,In_4262,In_4748);
nand U6534 (N_6534,In_3073,In_3681);
nor U6535 (N_6535,In_2894,In_4183);
or U6536 (N_6536,In_1580,In_3750);
and U6537 (N_6537,In_2868,In_1546);
nand U6538 (N_6538,In_4324,In_1824);
and U6539 (N_6539,In_190,In_4660);
or U6540 (N_6540,In_1663,In_4806);
nor U6541 (N_6541,In_425,In_3994);
or U6542 (N_6542,In_4757,In_4602);
or U6543 (N_6543,In_2088,In_3994);
and U6544 (N_6544,In_3199,In_4413);
and U6545 (N_6545,In_4063,In_2334);
nor U6546 (N_6546,In_650,In_2529);
xnor U6547 (N_6547,In_540,In_1401);
nor U6548 (N_6548,In_2463,In_4855);
nor U6549 (N_6549,In_2110,In_4290);
or U6550 (N_6550,In_857,In_770);
nor U6551 (N_6551,In_4875,In_3497);
nor U6552 (N_6552,In_2707,In_121);
nand U6553 (N_6553,In_2985,In_2614);
xnor U6554 (N_6554,In_1779,In_4424);
nor U6555 (N_6555,In_3079,In_1925);
or U6556 (N_6556,In_2010,In_2403);
xnor U6557 (N_6557,In_2984,In_2496);
and U6558 (N_6558,In_2050,In_1301);
and U6559 (N_6559,In_1795,In_3743);
nand U6560 (N_6560,In_1452,In_2278);
xnor U6561 (N_6561,In_2346,In_4734);
or U6562 (N_6562,In_3209,In_2469);
or U6563 (N_6563,In_255,In_2433);
nand U6564 (N_6564,In_1171,In_2865);
xnor U6565 (N_6565,In_4533,In_2526);
xnor U6566 (N_6566,In_449,In_4416);
and U6567 (N_6567,In_529,In_4903);
nor U6568 (N_6568,In_1469,In_3840);
or U6569 (N_6569,In_2539,In_2721);
xor U6570 (N_6570,In_1358,In_1583);
nand U6571 (N_6571,In_2895,In_2023);
or U6572 (N_6572,In_4553,In_2023);
nor U6573 (N_6573,In_4327,In_2555);
nand U6574 (N_6574,In_505,In_4888);
nor U6575 (N_6575,In_3674,In_2163);
and U6576 (N_6576,In_4334,In_2211);
nand U6577 (N_6577,In_4748,In_2446);
nor U6578 (N_6578,In_3836,In_3025);
xor U6579 (N_6579,In_2125,In_1911);
nand U6580 (N_6580,In_647,In_3987);
xnor U6581 (N_6581,In_1627,In_3778);
nand U6582 (N_6582,In_920,In_1942);
nor U6583 (N_6583,In_50,In_18);
nor U6584 (N_6584,In_3141,In_1289);
nand U6585 (N_6585,In_4673,In_4657);
or U6586 (N_6586,In_4088,In_252);
nand U6587 (N_6587,In_4324,In_2260);
or U6588 (N_6588,In_3755,In_167);
nor U6589 (N_6589,In_1873,In_4070);
or U6590 (N_6590,In_2816,In_2420);
or U6591 (N_6591,In_2941,In_2494);
nor U6592 (N_6592,In_2420,In_4413);
and U6593 (N_6593,In_510,In_2128);
nor U6594 (N_6594,In_1899,In_2245);
and U6595 (N_6595,In_1759,In_1233);
or U6596 (N_6596,In_641,In_4463);
and U6597 (N_6597,In_4409,In_1486);
or U6598 (N_6598,In_511,In_4815);
or U6599 (N_6599,In_596,In_3264);
nand U6600 (N_6600,In_4202,In_686);
and U6601 (N_6601,In_3592,In_280);
nand U6602 (N_6602,In_3824,In_836);
xnor U6603 (N_6603,In_4174,In_1111);
and U6604 (N_6604,In_4016,In_2356);
or U6605 (N_6605,In_1034,In_2544);
nor U6606 (N_6606,In_1559,In_531);
and U6607 (N_6607,In_2507,In_386);
nor U6608 (N_6608,In_4857,In_1048);
and U6609 (N_6609,In_3144,In_2679);
xnor U6610 (N_6610,In_2935,In_526);
and U6611 (N_6611,In_3004,In_3232);
nand U6612 (N_6612,In_94,In_3464);
nor U6613 (N_6613,In_1955,In_2933);
nand U6614 (N_6614,In_3140,In_167);
nand U6615 (N_6615,In_88,In_2439);
and U6616 (N_6616,In_4653,In_638);
or U6617 (N_6617,In_2140,In_4171);
nor U6618 (N_6618,In_417,In_648);
and U6619 (N_6619,In_4557,In_3830);
and U6620 (N_6620,In_3402,In_2765);
xnor U6621 (N_6621,In_942,In_309);
and U6622 (N_6622,In_1463,In_2731);
or U6623 (N_6623,In_4403,In_272);
nor U6624 (N_6624,In_439,In_4400);
or U6625 (N_6625,In_4441,In_2739);
or U6626 (N_6626,In_4704,In_3198);
or U6627 (N_6627,In_1751,In_3074);
and U6628 (N_6628,In_2012,In_3115);
nor U6629 (N_6629,In_4796,In_4030);
or U6630 (N_6630,In_364,In_3104);
or U6631 (N_6631,In_984,In_4559);
or U6632 (N_6632,In_4534,In_3109);
nand U6633 (N_6633,In_2336,In_4432);
or U6634 (N_6634,In_3449,In_4601);
and U6635 (N_6635,In_4609,In_2269);
nand U6636 (N_6636,In_385,In_1982);
nand U6637 (N_6637,In_4517,In_2341);
and U6638 (N_6638,In_4558,In_3999);
or U6639 (N_6639,In_598,In_2513);
nor U6640 (N_6640,In_4640,In_3894);
or U6641 (N_6641,In_4275,In_1740);
and U6642 (N_6642,In_3322,In_1111);
and U6643 (N_6643,In_2394,In_2703);
or U6644 (N_6644,In_2934,In_1590);
xor U6645 (N_6645,In_4147,In_605);
and U6646 (N_6646,In_2820,In_4495);
and U6647 (N_6647,In_737,In_4914);
and U6648 (N_6648,In_431,In_3425);
nand U6649 (N_6649,In_2719,In_747);
or U6650 (N_6650,In_619,In_4615);
and U6651 (N_6651,In_3101,In_4249);
nor U6652 (N_6652,In_2386,In_2372);
xnor U6653 (N_6653,In_484,In_287);
xor U6654 (N_6654,In_1244,In_1395);
xor U6655 (N_6655,In_175,In_2870);
nand U6656 (N_6656,In_1178,In_743);
and U6657 (N_6657,In_3305,In_2701);
and U6658 (N_6658,In_1235,In_1841);
or U6659 (N_6659,In_2197,In_4251);
nand U6660 (N_6660,In_3330,In_49);
nand U6661 (N_6661,In_4296,In_1519);
nand U6662 (N_6662,In_4401,In_34);
nand U6663 (N_6663,In_3711,In_4802);
or U6664 (N_6664,In_4393,In_4851);
or U6665 (N_6665,In_3984,In_502);
or U6666 (N_6666,In_3703,In_2535);
nor U6667 (N_6667,In_133,In_2036);
nand U6668 (N_6668,In_2802,In_3827);
nor U6669 (N_6669,In_3677,In_1458);
xnor U6670 (N_6670,In_3597,In_4280);
or U6671 (N_6671,In_3804,In_230);
and U6672 (N_6672,In_342,In_4001);
nor U6673 (N_6673,In_1057,In_4934);
nand U6674 (N_6674,In_143,In_2820);
nor U6675 (N_6675,In_2967,In_313);
nor U6676 (N_6676,In_3209,In_4811);
or U6677 (N_6677,In_4575,In_4528);
and U6678 (N_6678,In_3766,In_2735);
nand U6679 (N_6679,In_3695,In_4355);
and U6680 (N_6680,In_3227,In_1000);
or U6681 (N_6681,In_4872,In_3396);
or U6682 (N_6682,In_3574,In_2933);
nand U6683 (N_6683,In_1807,In_4662);
nand U6684 (N_6684,In_3031,In_1102);
nor U6685 (N_6685,In_228,In_4196);
or U6686 (N_6686,In_2753,In_2291);
and U6687 (N_6687,In_3553,In_756);
nand U6688 (N_6688,In_976,In_1367);
or U6689 (N_6689,In_3885,In_3865);
and U6690 (N_6690,In_1574,In_609);
and U6691 (N_6691,In_3309,In_217);
xnor U6692 (N_6692,In_1068,In_1161);
and U6693 (N_6693,In_1577,In_600);
or U6694 (N_6694,In_3963,In_1635);
or U6695 (N_6695,In_549,In_2575);
nand U6696 (N_6696,In_3113,In_1818);
nor U6697 (N_6697,In_2413,In_3469);
nand U6698 (N_6698,In_2437,In_3047);
nand U6699 (N_6699,In_882,In_2114);
nor U6700 (N_6700,In_1903,In_4342);
and U6701 (N_6701,In_3653,In_2671);
nor U6702 (N_6702,In_2049,In_757);
nand U6703 (N_6703,In_4560,In_722);
and U6704 (N_6704,In_3871,In_959);
or U6705 (N_6705,In_4204,In_4664);
xor U6706 (N_6706,In_3786,In_619);
nand U6707 (N_6707,In_1803,In_1406);
xnor U6708 (N_6708,In_3309,In_4093);
xnor U6709 (N_6709,In_2675,In_926);
nor U6710 (N_6710,In_1085,In_2173);
nand U6711 (N_6711,In_83,In_4400);
and U6712 (N_6712,In_1996,In_4500);
and U6713 (N_6713,In_4697,In_2319);
and U6714 (N_6714,In_3147,In_4726);
nor U6715 (N_6715,In_126,In_446);
xnor U6716 (N_6716,In_870,In_149);
nor U6717 (N_6717,In_3254,In_4694);
nand U6718 (N_6718,In_4445,In_1975);
nor U6719 (N_6719,In_1861,In_3052);
and U6720 (N_6720,In_794,In_3068);
nor U6721 (N_6721,In_2512,In_4248);
xnor U6722 (N_6722,In_1805,In_87);
nor U6723 (N_6723,In_2717,In_3135);
or U6724 (N_6724,In_122,In_1437);
nand U6725 (N_6725,In_2157,In_506);
nand U6726 (N_6726,In_1696,In_4928);
nand U6727 (N_6727,In_1414,In_1208);
nand U6728 (N_6728,In_1259,In_1326);
and U6729 (N_6729,In_1110,In_2054);
or U6730 (N_6730,In_4405,In_2763);
and U6731 (N_6731,In_3630,In_4788);
and U6732 (N_6732,In_3564,In_4833);
nand U6733 (N_6733,In_3314,In_3011);
nor U6734 (N_6734,In_4770,In_3865);
nor U6735 (N_6735,In_236,In_311);
nand U6736 (N_6736,In_4933,In_2003);
xnor U6737 (N_6737,In_1594,In_4449);
nor U6738 (N_6738,In_1799,In_1358);
or U6739 (N_6739,In_3691,In_3069);
xnor U6740 (N_6740,In_1208,In_1044);
nor U6741 (N_6741,In_400,In_3443);
xor U6742 (N_6742,In_2728,In_3864);
and U6743 (N_6743,In_1163,In_1983);
or U6744 (N_6744,In_1246,In_4442);
or U6745 (N_6745,In_950,In_1358);
xor U6746 (N_6746,In_2933,In_3482);
nand U6747 (N_6747,In_3608,In_1947);
or U6748 (N_6748,In_3136,In_4714);
or U6749 (N_6749,In_4973,In_2103);
and U6750 (N_6750,In_828,In_2056);
nor U6751 (N_6751,In_3412,In_2914);
nand U6752 (N_6752,In_1804,In_1718);
nand U6753 (N_6753,In_4566,In_2614);
and U6754 (N_6754,In_3913,In_2841);
or U6755 (N_6755,In_2516,In_472);
and U6756 (N_6756,In_1372,In_797);
or U6757 (N_6757,In_2090,In_4922);
or U6758 (N_6758,In_2128,In_3418);
nor U6759 (N_6759,In_985,In_3214);
and U6760 (N_6760,In_3362,In_3209);
or U6761 (N_6761,In_139,In_2224);
and U6762 (N_6762,In_1095,In_188);
and U6763 (N_6763,In_4283,In_1433);
and U6764 (N_6764,In_2108,In_3755);
or U6765 (N_6765,In_4706,In_2038);
nand U6766 (N_6766,In_1079,In_2216);
nor U6767 (N_6767,In_1080,In_1763);
nand U6768 (N_6768,In_1052,In_1635);
nor U6769 (N_6769,In_4404,In_2388);
nor U6770 (N_6770,In_2440,In_1789);
or U6771 (N_6771,In_1087,In_1786);
and U6772 (N_6772,In_4455,In_4593);
nand U6773 (N_6773,In_3371,In_4779);
nand U6774 (N_6774,In_524,In_3624);
nor U6775 (N_6775,In_1759,In_3353);
nor U6776 (N_6776,In_1336,In_1704);
or U6777 (N_6777,In_2388,In_3716);
and U6778 (N_6778,In_979,In_4346);
or U6779 (N_6779,In_3278,In_146);
or U6780 (N_6780,In_221,In_3136);
nor U6781 (N_6781,In_3840,In_3114);
nor U6782 (N_6782,In_4182,In_79);
xnor U6783 (N_6783,In_4452,In_4811);
nand U6784 (N_6784,In_2071,In_1953);
or U6785 (N_6785,In_3761,In_2554);
nor U6786 (N_6786,In_2796,In_2246);
nor U6787 (N_6787,In_2942,In_3392);
or U6788 (N_6788,In_2447,In_3774);
and U6789 (N_6789,In_212,In_4904);
and U6790 (N_6790,In_452,In_591);
nand U6791 (N_6791,In_4991,In_3404);
or U6792 (N_6792,In_3714,In_4871);
and U6793 (N_6793,In_4946,In_4132);
nand U6794 (N_6794,In_2263,In_2273);
or U6795 (N_6795,In_1604,In_2295);
nand U6796 (N_6796,In_632,In_487);
or U6797 (N_6797,In_1717,In_4812);
and U6798 (N_6798,In_4504,In_1651);
and U6799 (N_6799,In_2843,In_3400);
or U6800 (N_6800,In_3964,In_2276);
or U6801 (N_6801,In_3740,In_542);
or U6802 (N_6802,In_2987,In_2455);
nand U6803 (N_6803,In_856,In_950);
nor U6804 (N_6804,In_3820,In_3231);
xnor U6805 (N_6805,In_4994,In_3211);
or U6806 (N_6806,In_685,In_2672);
nand U6807 (N_6807,In_4212,In_3171);
nand U6808 (N_6808,In_2407,In_3101);
and U6809 (N_6809,In_2381,In_4310);
or U6810 (N_6810,In_759,In_4474);
nand U6811 (N_6811,In_1205,In_1402);
nor U6812 (N_6812,In_3777,In_4967);
nor U6813 (N_6813,In_3728,In_3086);
nor U6814 (N_6814,In_71,In_2891);
nor U6815 (N_6815,In_2992,In_3709);
and U6816 (N_6816,In_657,In_305);
and U6817 (N_6817,In_119,In_3964);
nand U6818 (N_6818,In_1732,In_188);
and U6819 (N_6819,In_678,In_4263);
or U6820 (N_6820,In_2652,In_3409);
nor U6821 (N_6821,In_2452,In_3072);
nor U6822 (N_6822,In_3297,In_3901);
and U6823 (N_6823,In_2148,In_3418);
nand U6824 (N_6824,In_2967,In_4923);
xnor U6825 (N_6825,In_3398,In_119);
nor U6826 (N_6826,In_507,In_2281);
nand U6827 (N_6827,In_4961,In_2593);
or U6828 (N_6828,In_2566,In_3708);
nand U6829 (N_6829,In_4701,In_1332);
xnor U6830 (N_6830,In_70,In_673);
nand U6831 (N_6831,In_1266,In_3970);
and U6832 (N_6832,In_1261,In_3537);
or U6833 (N_6833,In_2775,In_2329);
and U6834 (N_6834,In_890,In_1317);
nand U6835 (N_6835,In_2450,In_713);
nor U6836 (N_6836,In_4119,In_3276);
and U6837 (N_6837,In_1774,In_1446);
nor U6838 (N_6838,In_1056,In_2715);
nand U6839 (N_6839,In_74,In_3723);
or U6840 (N_6840,In_4804,In_2025);
nor U6841 (N_6841,In_42,In_2421);
or U6842 (N_6842,In_4591,In_194);
or U6843 (N_6843,In_2371,In_86);
nand U6844 (N_6844,In_4514,In_2218);
or U6845 (N_6845,In_4056,In_4136);
or U6846 (N_6846,In_3355,In_4269);
or U6847 (N_6847,In_3637,In_1485);
nand U6848 (N_6848,In_4527,In_3862);
nor U6849 (N_6849,In_1204,In_2409);
nand U6850 (N_6850,In_3503,In_2190);
nor U6851 (N_6851,In_1076,In_358);
or U6852 (N_6852,In_4442,In_1425);
xor U6853 (N_6853,In_2671,In_2237);
nor U6854 (N_6854,In_1839,In_4251);
and U6855 (N_6855,In_1712,In_4425);
nand U6856 (N_6856,In_2157,In_466);
xor U6857 (N_6857,In_107,In_608);
and U6858 (N_6858,In_2967,In_478);
and U6859 (N_6859,In_4892,In_1883);
or U6860 (N_6860,In_1622,In_1629);
nand U6861 (N_6861,In_1959,In_4598);
nor U6862 (N_6862,In_428,In_4864);
nand U6863 (N_6863,In_1989,In_1522);
nor U6864 (N_6864,In_1888,In_870);
nand U6865 (N_6865,In_2858,In_4956);
and U6866 (N_6866,In_332,In_4081);
and U6867 (N_6867,In_4067,In_453);
or U6868 (N_6868,In_4146,In_2594);
or U6869 (N_6869,In_2681,In_3492);
nand U6870 (N_6870,In_679,In_2642);
nor U6871 (N_6871,In_4671,In_2987);
or U6872 (N_6872,In_1350,In_2820);
nor U6873 (N_6873,In_2123,In_1151);
xnor U6874 (N_6874,In_2908,In_2169);
nand U6875 (N_6875,In_1473,In_1533);
or U6876 (N_6876,In_854,In_1806);
or U6877 (N_6877,In_3914,In_2897);
nor U6878 (N_6878,In_2655,In_156);
xnor U6879 (N_6879,In_3711,In_4230);
nand U6880 (N_6880,In_2480,In_2604);
nand U6881 (N_6881,In_1266,In_1359);
and U6882 (N_6882,In_506,In_1502);
nor U6883 (N_6883,In_3541,In_1024);
nand U6884 (N_6884,In_3318,In_4611);
nand U6885 (N_6885,In_3300,In_309);
nor U6886 (N_6886,In_3923,In_2594);
nand U6887 (N_6887,In_1643,In_2770);
and U6888 (N_6888,In_3799,In_3476);
and U6889 (N_6889,In_790,In_2250);
nor U6890 (N_6890,In_3116,In_3588);
and U6891 (N_6891,In_575,In_2572);
nor U6892 (N_6892,In_3480,In_1080);
nand U6893 (N_6893,In_3921,In_1705);
and U6894 (N_6894,In_1311,In_1991);
or U6895 (N_6895,In_2008,In_563);
or U6896 (N_6896,In_4264,In_4753);
and U6897 (N_6897,In_2060,In_1290);
or U6898 (N_6898,In_1711,In_3096);
or U6899 (N_6899,In_318,In_1218);
nor U6900 (N_6900,In_2863,In_2);
nand U6901 (N_6901,In_3492,In_1632);
xor U6902 (N_6902,In_892,In_2023);
nor U6903 (N_6903,In_4028,In_3169);
xnor U6904 (N_6904,In_4126,In_3589);
and U6905 (N_6905,In_4495,In_2677);
xor U6906 (N_6906,In_4344,In_1294);
nor U6907 (N_6907,In_3497,In_3928);
nand U6908 (N_6908,In_2664,In_2028);
nand U6909 (N_6909,In_3140,In_2208);
and U6910 (N_6910,In_2293,In_4369);
nand U6911 (N_6911,In_3839,In_4683);
and U6912 (N_6912,In_542,In_2054);
nand U6913 (N_6913,In_1867,In_4724);
or U6914 (N_6914,In_1668,In_1961);
nand U6915 (N_6915,In_297,In_248);
nand U6916 (N_6916,In_2368,In_2221);
nor U6917 (N_6917,In_4340,In_3415);
or U6918 (N_6918,In_3502,In_2215);
and U6919 (N_6919,In_4990,In_435);
nand U6920 (N_6920,In_4646,In_3883);
nand U6921 (N_6921,In_4935,In_2696);
or U6922 (N_6922,In_785,In_303);
or U6923 (N_6923,In_1366,In_2885);
and U6924 (N_6924,In_1723,In_2442);
xor U6925 (N_6925,In_4962,In_1829);
or U6926 (N_6926,In_2116,In_508);
and U6927 (N_6927,In_1479,In_1254);
nor U6928 (N_6928,In_2853,In_126);
or U6929 (N_6929,In_2926,In_2309);
nor U6930 (N_6930,In_1801,In_3774);
xnor U6931 (N_6931,In_2582,In_2560);
and U6932 (N_6932,In_2097,In_1039);
and U6933 (N_6933,In_352,In_3418);
nand U6934 (N_6934,In_3019,In_2408);
and U6935 (N_6935,In_3961,In_4819);
or U6936 (N_6936,In_729,In_1411);
nand U6937 (N_6937,In_4733,In_2170);
or U6938 (N_6938,In_2879,In_4129);
and U6939 (N_6939,In_4492,In_1160);
nand U6940 (N_6940,In_4801,In_519);
nor U6941 (N_6941,In_976,In_4790);
and U6942 (N_6942,In_2998,In_1529);
nor U6943 (N_6943,In_2868,In_3540);
nand U6944 (N_6944,In_3123,In_490);
nand U6945 (N_6945,In_4647,In_1835);
and U6946 (N_6946,In_1641,In_416);
nand U6947 (N_6947,In_2840,In_2128);
nor U6948 (N_6948,In_872,In_3335);
or U6949 (N_6949,In_2469,In_220);
nand U6950 (N_6950,In_3724,In_4976);
or U6951 (N_6951,In_3701,In_1026);
xnor U6952 (N_6952,In_4496,In_1046);
and U6953 (N_6953,In_1169,In_2865);
nor U6954 (N_6954,In_687,In_2784);
or U6955 (N_6955,In_916,In_1987);
and U6956 (N_6956,In_1823,In_1251);
nand U6957 (N_6957,In_1479,In_2128);
nor U6958 (N_6958,In_1159,In_612);
nand U6959 (N_6959,In_3975,In_2610);
or U6960 (N_6960,In_2798,In_3425);
or U6961 (N_6961,In_3872,In_479);
nand U6962 (N_6962,In_734,In_662);
or U6963 (N_6963,In_3756,In_511);
nor U6964 (N_6964,In_412,In_1689);
and U6965 (N_6965,In_2780,In_4815);
nor U6966 (N_6966,In_3349,In_4401);
or U6967 (N_6967,In_4747,In_3440);
nor U6968 (N_6968,In_2420,In_4275);
nor U6969 (N_6969,In_272,In_4566);
and U6970 (N_6970,In_2113,In_3826);
nor U6971 (N_6971,In_249,In_647);
nor U6972 (N_6972,In_662,In_470);
nand U6973 (N_6973,In_1710,In_1761);
nand U6974 (N_6974,In_607,In_3663);
nor U6975 (N_6975,In_72,In_2195);
nor U6976 (N_6976,In_2586,In_3473);
and U6977 (N_6977,In_4077,In_241);
or U6978 (N_6978,In_355,In_4036);
and U6979 (N_6979,In_1522,In_2194);
nand U6980 (N_6980,In_3141,In_3115);
nor U6981 (N_6981,In_3963,In_2267);
nor U6982 (N_6982,In_4241,In_2276);
or U6983 (N_6983,In_1553,In_2249);
xor U6984 (N_6984,In_4149,In_3805);
nor U6985 (N_6985,In_709,In_2925);
or U6986 (N_6986,In_1156,In_538);
or U6987 (N_6987,In_792,In_1846);
or U6988 (N_6988,In_4430,In_4851);
nor U6989 (N_6989,In_2159,In_3509);
nor U6990 (N_6990,In_4866,In_1016);
or U6991 (N_6991,In_1438,In_2319);
and U6992 (N_6992,In_484,In_2159);
and U6993 (N_6993,In_2933,In_182);
and U6994 (N_6994,In_3851,In_4203);
or U6995 (N_6995,In_3966,In_549);
and U6996 (N_6996,In_1700,In_4802);
or U6997 (N_6997,In_2010,In_4503);
nand U6998 (N_6998,In_2386,In_4786);
and U6999 (N_6999,In_4513,In_1168);
nand U7000 (N_7000,In_2872,In_2133);
nand U7001 (N_7001,In_3344,In_3762);
nand U7002 (N_7002,In_109,In_1729);
xnor U7003 (N_7003,In_2103,In_4910);
or U7004 (N_7004,In_4348,In_2472);
nand U7005 (N_7005,In_1702,In_1300);
nand U7006 (N_7006,In_4553,In_4954);
nor U7007 (N_7007,In_4282,In_378);
nand U7008 (N_7008,In_2063,In_2676);
nor U7009 (N_7009,In_3728,In_2483);
or U7010 (N_7010,In_4540,In_4842);
or U7011 (N_7011,In_1171,In_2878);
or U7012 (N_7012,In_4139,In_1963);
or U7013 (N_7013,In_2260,In_945);
and U7014 (N_7014,In_2728,In_2471);
and U7015 (N_7015,In_1745,In_2246);
or U7016 (N_7016,In_1936,In_2124);
nor U7017 (N_7017,In_3118,In_2721);
or U7018 (N_7018,In_4926,In_1924);
nor U7019 (N_7019,In_4212,In_1298);
nand U7020 (N_7020,In_1784,In_1516);
nor U7021 (N_7021,In_3610,In_447);
nor U7022 (N_7022,In_2403,In_4228);
nand U7023 (N_7023,In_3059,In_4477);
nor U7024 (N_7024,In_300,In_1322);
nor U7025 (N_7025,In_2380,In_2000);
or U7026 (N_7026,In_1710,In_2977);
nor U7027 (N_7027,In_831,In_2587);
nand U7028 (N_7028,In_4002,In_4958);
or U7029 (N_7029,In_2587,In_1525);
or U7030 (N_7030,In_732,In_4263);
or U7031 (N_7031,In_1733,In_2906);
nor U7032 (N_7032,In_1572,In_3719);
and U7033 (N_7033,In_4538,In_4275);
nor U7034 (N_7034,In_2432,In_4217);
and U7035 (N_7035,In_4977,In_2148);
or U7036 (N_7036,In_368,In_2740);
nand U7037 (N_7037,In_3250,In_1035);
or U7038 (N_7038,In_2143,In_2395);
and U7039 (N_7039,In_3331,In_2763);
or U7040 (N_7040,In_3068,In_2395);
and U7041 (N_7041,In_809,In_3794);
or U7042 (N_7042,In_1118,In_4533);
and U7043 (N_7043,In_2962,In_2664);
nand U7044 (N_7044,In_262,In_2070);
nand U7045 (N_7045,In_308,In_1052);
nor U7046 (N_7046,In_97,In_2390);
and U7047 (N_7047,In_823,In_2506);
nor U7048 (N_7048,In_63,In_58);
and U7049 (N_7049,In_2497,In_766);
and U7050 (N_7050,In_2445,In_4325);
nand U7051 (N_7051,In_2113,In_3661);
nor U7052 (N_7052,In_3876,In_2043);
or U7053 (N_7053,In_2740,In_3108);
nor U7054 (N_7054,In_3135,In_114);
or U7055 (N_7055,In_138,In_3907);
nand U7056 (N_7056,In_2209,In_2983);
and U7057 (N_7057,In_3679,In_2742);
nor U7058 (N_7058,In_4474,In_1617);
xnor U7059 (N_7059,In_2557,In_2558);
and U7060 (N_7060,In_4124,In_2266);
nor U7061 (N_7061,In_1303,In_2264);
nor U7062 (N_7062,In_4101,In_1910);
xnor U7063 (N_7063,In_3107,In_2649);
and U7064 (N_7064,In_4946,In_2652);
and U7065 (N_7065,In_2752,In_2036);
nand U7066 (N_7066,In_3076,In_1202);
nand U7067 (N_7067,In_2614,In_3677);
nor U7068 (N_7068,In_31,In_2422);
and U7069 (N_7069,In_4105,In_4241);
xnor U7070 (N_7070,In_3482,In_3905);
nor U7071 (N_7071,In_2279,In_169);
xnor U7072 (N_7072,In_2361,In_188);
nor U7073 (N_7073,In_4272,In_2246);
nand U7074 (N_7074,In_3020,In_2223);
or U7075 (N_7075,In_1751,In_4301);
and U7076 (N_7076,In_4795,In_2599);
nor U7077 (N_7077,In_3445,In_2628);
nand U7078 (N_7078,In_3252,In_443);
nand U7079 (N_7079,In_4889,In_2459);
nand U7080 (N_7080,In_780,In_1859);
nand U7081 (N_7081,In_4302,In_1952);
and U7082 (N_7082,In_542,In_4171);
xor U7083 (N_7083,In_626,In_2865);
and U7084 (N_7084,In_3347,In_4965);
and U7085 (N_7085,In_2749,In_4724);
nand U7086 (N_7086,In_1543,In_181);
and U7087 (N_7087,In_2405,In_565);
nor U7088 (N_7088,In_836,In_1053);
nand U7089 (N_7089,In_4142,In_2202);
nor U7090 (N_7090,In_2776,In_4081);
nand U7091 (N_7091,In_79,In_2341);
or U7092 (N_7092,In_3344,In_4151);
xnor U7093 (N_7093,In_2221,In_508);
nor U7094 (N_7094,In_3888,In_2802);
or U7095 (N_7095,In_4362,In_2695);
nor U7096 (N_7096,In_1006,In_218);
or U7097 (N_7097,In_2460,In_1320);
nand U7098 (N_7098,In_561,In_3950);
or U7099 (N_7099,In_1310,In_3396);
or U7100 (N_7100,In_531,In_396);
or U7101 (N_7101,In_1129,In_3897);
and U7102 (N_7102,In_448,In_4356);
nor U7103 (N_7103,In_4849,In_268);
nor U7104 (N_7104,In_3542,In_3443);
nand U7105 (N_7105,In_1544,In_3035);
nand U7106 (N_7106,In_4811,In_441);
and U7107 (N_7107,In_4531,In_4050);
or U7108 (N_7108,In_2277,In_1606);
nand U7109 (N_7109,In_3582,In_2353);
and U7110 (N_7110,In_1402,In_1576);
nor U7111 (N_7111,In_1859,In_4172);
xor U7112 (N_7112,In_2805,In_619);
nor U7113 (N_7113,In_3895,In_351);
nand U7114 (N_7114,In_1833,In_4207);
nand U7115 (N_7115,In_2957,In_4846);
or U7116 (N_7116,In_4084,In_2205);
xnor U7117 (N_7117,In_3778,In_1855);
or U7118 (N_7118,In_4404,In_875);
nor U7119 (N_7119,In_3299,In_3710);
xnor U7120 (N_7120,In_1133,In_4798);
nand U7121 (N_7121,In_3504,In_61);
nor U7122 (N_7122,In_4827,In_1274);
nor U7123 (N_7123,In_3372,In_3208);
or U7124 (N_7124,In_2534,In_4280);
or U7125 (N_7125,In_3047,In_3534);
and U7126 (N_7126,In_2111,In_1073);
and U7127 (N_7127,In_3758,In_1091);
nor U7128 (N_7128,In_104,In_1430);
and U7129 (N_7129,In_705,In_3702);
xor U7130 (N_7130,In_615,In_790);
or U7131 (N_7131,In_3331,In_2197);
nor U7132 (N_7132,In_1433,In_1553);
and U7133 (N_7133,In_1020,In_4026);
nor U7134 (N_7134,In_2268,In_2683);
or U7135 (N_7135,In_1915,In_4441);
and U7136 (N_7136,In_1402,In_3533);
nand U7137 (N_7137,In_925,In_958);
nand U7138 (N_7138,In_2562,In_833);
nor U7139 (N_7139,In_204,In_4233);
or U7140 (N_7140,In_3054,In_48);
nand U7141 (N_7141,In_455,In_3424);
xnor U7142 (N_7142,In_4494,In_1694);
and U7143 (N_7143,In_2375,In_152);
nand U7144 (N_7144,In_121,In_4824);
xnor U7145 (N_7145,In_350,In_4714);
or U7146 (N_7146,In_1092,In_4673);
nand U7147 (N_7147,In_1532,In_1954);
and U7148 (N_7148,In_120,In_1835);
and U7149 (N_7149,In_2854,In_4495);
nor U7150 (N_7150,In_2476,In_3421);
and U7151 (N_7151,In_1884,In_4956);
and U7152 (N_7152,In_3834,In_1788);
nand U7153 (N_7153,In_201,In_3394);
xor U7154 (N_7154,In_2646,In_198);
or U7155 (N_7155,In_3191,In_160);
and U7156 (N_7156,In_2916,In_3796);
nor U7157 (N_7157,In_3153,In_4208);
nor U7158 (N_7158,In_3567,In_430);
xor U7159 (N_7159,In_1707,In_1874);
nor U7160 (N_7160,In_1426,In_270);
and U7161 (N_7161,In_3744,In_4301);
or U7162 (N_7162,In_781,In_1762);
and U7163 (N_7163,In_2552,In_988);
or U7164 (N_7164,In_3929,In_68);
nand U7165 (N_7165,In_1189,In_826);
and U7166 (N_7166,In_884,In_3147);
nand U7167 (N_7167,In_4732,In_578);
nor U7168 (N_7168,In_465,In_2754);
nor U7169 (N_7169,In_362,In_1337);
nand U7170 (N_7170,In_1044,In_801);
nand U7171 (N_7171,In_3322,In_2326);
nand U7172 (N_7172,In_1617,In_3454);
nand U7173 (N_7173,In_558,In_3862);
xnor U7174 (N_7174,In_3588,In_1803);
nor U7175 (N_7175,In_3060,In_1199);
and U7176 (N_7176,In_4772,In_2327);
and U7177 (N_7177,In_1373,In_1076);
nand U7178 (N_7178,In_2551,In_3790);
or U7179 (N_7179,In_3091,In_4983);
nor U7180 (N_7180,In_43,In_4761);
nand U7181 (N_7181,In_167,In_599);
nor U7182 (N_7182,In_2230,In_1161);
and U7183 (N_7183,In_930,In_655);
and U7184 (N_7184,In_4026,In_2924);
nand U7185 (N_7185,In_1610,In_734);
or U7186 (N_7186,In_3382,In_224);
nand U7187 (N_7187,In_3240,In_243);
and U7188 (N_7188,In_3057,In_2983);
or U7189 (N_7189,In_174,In_600);
nor U7190 (N_7190,In_4307,In_3965);
nor U7191 (N_7191,In_3094,In_2646);
and U7192 (N_7192,In_3628,In_4676);
nand U7193 (N_7193,In_3357,In_4541);
nand U7194 (N_7194,In_278,In_2578);
nand U7195 (N_7195,In_2411,In_3690);
or U7196 (N_7196,In_1080,In_749);
or U7197 (N_7197,In_3383,In_2030);
nand U7198 (N_7198,In_3661,In_685);
nand U7199 (N_7199,In_2026,In_4835);
nand U7200 (N_7200,In_4099,In_703);
and U7201 (N_7201,In_1353,In_192);
or U7202 (N_7202,In_2124,In_1540);
or U7203 (N_7203,In_2794,In_2365);
nor U7204 (N_7204,In_1126,In_3125);
and U7205 (N_7205,In_1368,In_2738);
nor U7206 (N_7206,In_4646,In_1674);
nor U7207 (N_7207,In_1937,In_1187);
or U7208 (N_7208,In_3831,In_1811);
nand U7209 (N_7209,In_812,In_376);
or U7210 (N_7210,In_1904,In_2322);
nor U7211 (N_7211,In_432,In_2972);
nand U7212 (N_7212,In_4408,In_335);
nand U7213 (N_7213,In_794,In_2971);
and U7214 (N_7214,In_3463,In_2972);
or U7215 (N_7215,In_4655,In_4120);
nor U7216 (N_7216,In_945,In_1266);
or U7217 (N_7217,In_2310,In_4685);
or U7218 (N_7218,In_2477,In_2878);
nor U7219 (N_7219,In_1723,In_1395);
nor U7220 (N_7220,In_1987,In_3786);
and U7221 (N_7221,In_1866,In_505);
and U7222 (N_7222,In_616,In_846);
and U7223 (N_7223,In_48,In_1101);
xor U7224 (N_7224,In_3836,In_1860);
nor U7225 (N_7225,In_769,In_2801);
nor U7226 (N_7226,In_1891,In_2083);
and U7227 (N_7227,In_1460,In_2014);
or U7228 (N_7228,In_4559,In_1175);
nor U7229 (N_7229,In_4367,In_1172);
or U7230 (N_7230,In_4113,In_3817);
and U7231 (N_7231,In_2770,In_736);
nor U7232 (N_7232,In_2016,In_194);
xnor U7233 (N_7233,In_2716,In_1958);
xnor U7234 (N_7234,In_3022,In_4037);
nand U7235 (N_7235,In_4803,In_2125);
xor U7236 (N_7236,In_3580,In_3493);
nor U7237 (N_7237,In_4747,In_2206);
nor U7238 (N_7238,In_2926,In_3638);
xor U7239 (N_7239,In_4013,In_3247);
and U7240 (N_7240,In_965,In_2001);
nand U7241 (N_7241,In_3359,In_1271);
xnor U7242 (N_7242,In_1188,In_4994);
or U7243 (N_7243,In_2617,In_4453);
nand U7244 (N_7244,In_2483,In_631);
nor U7245 (N_7245,In_188,In_2526);
and U7246 (N_7246,In_931,In_2991);
or U7247 (N_7247,In_2549,In_1243);
nand U7248 (N_7248,In_1741,In_2664);
nor U7249 (N_7249,In_3747,In_4898);
xnor U7250 (N_7250,In_3595,In_1264);
nand U7251 (N_7251,In_4636,In_4281);
nand U7252 (N_7252,In_3273,In_3397);
nor U7253 (N_7253,In_4178,In_4011);
nor U7254 (N_7254,In_734,In_576);
nand U7255 (N_7255,In_3275,In_2285);
or U7256 (N_7256,In_3948,In_2604);
or U7257 (N_7257,In_354,In_4154);
and U7258 (N_7258,In_3729,In_2604);
nand U7259 (N_7259,In_2394,In_2507);
xnor U7260 (N_7260,In_4343,In_3827);
or U7261 (N_7261,In_2512,In_3971);
or U7262 (N_7262,In_3222,In_249);
and U7263 (N_7263,In_2911,In_605);
or U7264 (N_7264,In_1339,In_4225);
or U7265 (N_7265,In_712,In_2412);
and U7266 (N_7266,In_4766,In_4756);
and U7267 (N_7267,In_1206,In_4844);
or U7268 (N_7268,In_2710,In_4079);
nor U7269 (N_7269,In_3785,In_2510);
and U7270 (N_7270,In_690,In_717);
nand U7271 (N_7271,In_252,In_873);
and U7272 (N_7272,In_726,In_4436);
nand U7273 (N_7273,In_3179,In_15);
nand U7274 (N_7274,In_4329,In_371);
nand U7275 (N_7275,In_3046,In_1336);
nand U7276 (N_7276,In_958,In_3706);
and U7277 (N_7277,In_3221,In_4875);
nand U7278 (N_7278,In_3810,In_2114);
nor U7279 (N_7279,In_4545,In_1796);
nand U7280 (N_7280,In_3137,In_1619);
nor U7281 (N_7281,In_3117,In_1773);
nand U7282 (N_7282,In_3960,In_4326);
nand U7283 (N_7283,In_515,In_2847);
nand U7284 (N_7284,In_384,In_2437);
or U7285 (N_7285,In_3126,In_1450);
and U7286 (N_7286,In_3960,In_4968);
nand U7287 (N_7287,In_1499,In_1073);
nor U7288 (N_7288,In_1777,In_1361);
nor U7289 (N_7289,In_448,In_458);
xnor U7290 (N_7290,In_1981,In_3541);
or U7291 (N_7291,In_4966,In_4770);
and U7292 (N_7292,In_4035,In_1463);
nand U7293 (N_7293,In_3996,In_4464);
and U7294 (N_7294,In_3705,In_2499);
or U7295 (N_7295,In_4549,In_3297);
and U7296 (N_7296,In_4145,In_3978);
nand U7297 (N_7297,In_2190,In_1255);
nor U7298 (N_7298,In_1796,In_4433);
xor U7299 (N_7299,In_2580,In_4339);
xnor U7300 (N_7300,In_2452,In_2730);
nand U7301 (N_7301,In_4365,In_1546);
nor U7302 (N_7302,In_3007,In_4244);
or U7303 (N_7303,In_1829,In_252);
nand U7304 (N_7304,In_3730,In_3262);
or U7305 (N_7305,In_2608,In_4825);
nor U7306 (N_7306,In_1377,In_4023);
nor U7307 (N_7307,In_2298,In_223);
nor U7308 (N_7308,In_4631,In_2766);
and U7309 (N_7309,In_2536,In_279);
or U7310 (N_7310,In_3762,In_1260);
xor U7311 (N_7311,In_1921,In_3117);
xor U7312 (N_7312,In_1399,In_2613);
or U7313 (N_7313,In_685,In_1262);
and U7314 (N_7314,In_1565,In_3145);
nor U7315 (N_7315,In_2519,In_3968);
and U7316 (N_7316,In_4749,In_3899);
nand U7317 (N_7317,In_4392,In_2659);
nor U7318 (N_7318,In_1158,In_4082);
nor U7319 (N_7319,In_667,In_2204);
nor U7320 (N_7320,In_99,In_4006);
and U7321 (N_7321,In_1951,In_187);
nor U7322 (N_7322,In_2964,In_1049);
and U7323 (N_7323,In_682,In_3621);
or U7324 (N_7324,In_2994,In_463);
or U7325 (N_7325,In_973,In_1368);
nand U7326 (N_7326,In_2151,In_2894);
and U7327 (N_7327,In_2854,In_1282);
or U7328 (N_7328,In_1273,In_3845);
nand U7329 (N_7329,In_396,In_1576);
nand U7330 (N_7330,In_2898,In_4443);
nor U7331 (N_7331,In_4876,In_83);
or U7332 (N_7332,In_4595,In_1329);
and U7333 (N_7333,In_4088,In_2582);
or U7334 (N_7334,In_15,In_274);
xor U7335 (N_7335,In_1257,In_1105);
or U7336 (N_7336,In_2059,In_3751);
and U7337 (N_7337,In_209,In_391);
xnor U7338 (N_7338,In_2227,In_3510);
nor U7339 (N_7339,In_4114,In_2364);
nand U7340 (N_7340,In_1215,In_3291);
nor U7341 (N_7341,In_4586,In_1744);
or U7342 (N_7342,In_4806,In_2221);
nand U7343 (N_7343,In_1888,In_591);
xor U7344 (N_7344,In_1684,In_63);
or U7345 (N_7345,In_4777,In_2019);
and U7346 (N_7346,In_2294,In_1133);
or U7347 (N_7347,In_4733,In_3963);
or U7348 (N_7348,In_1737,In_2189);
nand U7349 (N_7349,In_2602,In_2278);
and U7350 (N_7350,In_3568,In_3928);
and U7351 (N_7351,In_643,In_3592);
or U7352 (N_7352,In_4510,In_2026);
nand U7353 (N_7353,In_1087,In_892);
or U7354 (N_7354,In_185,In_4127);
nor U7355 (N_7355,In_3376,In_187);
nor U7356 (N_7356,In_2293,In_2563);
or U7357 (N_7357,In_4715,In_1834);
and U7358 (N_7358,In_54,In_1949);
nor U7359 (N_7359,In_440,In_3624);
nand U7360 (N_7360,In_1123,In_375);
or U7361 (N_7361,In_1830,In_3447);
nor U7362 (N_7362,In_3374,In_1965);
or U7363 (N_7363,In_3848,In_1314);
nor U7364 (N_7364,In_4397,In_4509);
xor U7365 (N_7365,In_673,In_1794);
nand U7366 (N_7366,In_896,In_4330);
or U7367 (N_7367,In_370,In_2524);
nand U7368 (N_7368,In_1610,In_4522);
xnor U7369 (N_7369,In_2440,In_2244);
nand U7370 (N_7370,In_232,In_1893);
nor U7371 (N_7371,In_4818,In_2232);
nor U7372 (N_7372,In_832,In_1294);
nand U7373 (N_7373,In_60,In_3749);
nand U7374 (N_7374,In_2913,In_3586);
nor U7375 (N_7375,In_2915,In_3);
and U7376 (N_7376,In_148,In_527);
nand U7377 (N_7377,In_1297,In_1198);
nand U7378 (N_7378,In_3139,In_1125);
and U7379 (N_7379,In_3665,In_2024);
and U7380 (N_7380,In_4571,In_2122);
or U7381 (N_7381,In_180,In_3622);
nand U7382 (N_7382,In_3899,In_90);
xor U7383 (N_7383,In_449,In_4891);
and U7384 (N_7384,In_2301,In_2848);
nor U7385 (N_7385,In_171,In_2463);
nor U7386 (N_7386,In_296,In_3024);
nand U7387 (N_7387,In_1045,In_3781);
nand U7388 (N_7388,In_4461,In_519);
or U7389 (N_7389,In_4990,In_3901);
nand U7390 (N_7390,In_1635,In_4755);
and U7391 (N_7391,In_3614,In_2593);
nand U7392 (N_7392,In_4650,In_4461);
nand U7393 (N_7393,In_3891,In_1188);
nand U7394 (N_7394,In_1904,In_4050);
nor U7395 (N_7395,In_3166,In_3139);
nor U7396 (N_7396,In_2432,In_690);
nand U7397 (N_7397,In_3482,In_4012);
nand U7398 (N_7398,In_1626,In_2873);
and U7399 (N_7399,In_3893,In_2679);
nor U7400 (N_7400,In_4083,In_1766);
and U7401 (N_7401,In_482,In_2451);
and U7402 (N_7402,In_1208,In_2058);
or U7403 (N_7403,In_1619,In_749);
and U7404 (N_7404,In_3638,In_2790);
and U7405 (N_7405,In_2538,In_2731);
nand U7406 (N_7406,In_85,In_3577);
nand U7407 (N_7407,In_1758,In_4927);
xnor U7408 (N_7408,In_1461,In_2002);
or U7409 (N_7409,In_1445,In_160);
and U7410 (N_7410,In_1140,In_997);
nor U7411 (N_7411,In_4767,In_4962);
nand U7412 (N_7412,In_2078,In_1966);
nor U7413 (N_7413,In_2855,In_3385);
or U7414 (N_7414,In_4617,In_3757);
nor U7415 (N_7415,In_2613,In_2098);
nand U7416 (N_7416,In_4287,In_1150);
nor U7417 (N_7417,In_2449,In_1743);
xnor U7418 (N_7418,In_2923,In_3659);
and U7419 (N_7419,In_4714,In_4965);
xor U7420 (N_7420,In_4791,In_14);
and U7421 (N_7421,In_2031,In_3485);
nor U7422 (N_7422,In_928,In_2666);
xor U7423 (N_7423,In_2017,In_328);
and U7424 (N_7424,In_1119,In_2525);
nand U7425 (N_7425,In_408,In_4266);
or U7426 (N_7426,In_4412,In_773);
or U7427 (N_7427,In_1734,In_3);
xor U7428 (N_7428,In_515,In_1472);
and U7429 (N_7429,In_1910,In_1036);
nor U7430 (N_7430,In_3221,In_3621);
nand U7431 (N_7431,In_625,In_4867);
nor U7432 (N_7432,In_1093,In_4956);
and U7433 (N_7433,In_4754,In_502);
nand U7434 (N_7434,In_4383,In_1823);
or U7435 (N_7435,In_3761,In_3998);
or U7436 (N_7436,In_3559,In_4179);
xor U7437 (N_7437,In_340,In_3937);
nor U7438 (N_7438,In_4247,In_1271);
and U7439 (N_7439,In_3736,In_599);
or U7440 (N_7440,In_4828,In_3466);
nor U7441 (N_7441,In_156,In_4343);
xnor U7442 (N_7442,In_1368,In_1626);
nor U7443 (N_7443,In_4434,In_4037);
and U7444 (N_7444,In_1105,In_3409);
nand U7445 (N_7445,In_1054,In_4544);
nand U7446 (N_7446,In_2913,In_1963);
or U7447 (N_7447,In_1154,In_3400);
or U7448 (N_7448,In_4442,In_1134);
or U7449 (N_7449,In_2070,In_3155);
xnor U7450 (N_7450,In_3216,In_546);
nand U7451 (N_7451,In_120,In_2709);
xor U7452 (N_7452,In_394,In_2566);
nor U7453 (N_7453,In_1640,In_845);
nor U7454 (N_7454,In_1708,In_4691);
nand U7455 (N_7455,In_2390,In_4551);
xnor U7456 (N_7456,In_4750,In_2385);
nand U7457 (N_7457,In_2460,In_766);
nor U7458 (N_7458,In_1592,In_4905);
or U7459 (N_7459,In_707,In_1833);
and U7460 (N_7460,In_918,In_3158);
nand U7461 (N_7461,In_4610,In_445);
nor U7462 (N_7462,In_3019,In_2923);
xnor U7463 (N_7463,In_3525,In_559);
nand U7464 (N_7464,In_1662,In_1578);
or U7465 (N_7465,In_4642,In_461);
nor U7466 (N_7466,In_2742,In_3825);
nand U7467 (N_7467,In_3307,In_627);
xor U7468 (N_7468,In_3280,In_2868);
nand U7469 (N_7469,In_817,In_1200);
nand U7470 (N_7470,In_3918,In_3693);
nor U7471 (N_7471,In_2673,In_2803);
nand U7472 (N_7472,In_1338,In_4885);
and U7473 (N_7473,In_4739,In_807);
and U7474 (N_7474,In_1150,In_1058);
nand U7475 (N_7475,In_1533,In_1636);
or U7476 (N_7476,In_3589,In_3064);
and U7477 (N_7477,In_3704,In_4156);
or U7478 (N_7478,In_1369,In_3847);
or U7479 (N_7479,In_4121,In_2750);
nor U7480 (N_7480,In_1357,In_4670);
nand U7481 (N_7481,In_2977,In_837);
nand U7482 (N_7482,In_3654,In_3340);
nand U7483 (N_7483,In_4838,In_906);
or U7484 (N_7484,In_4747,In_1344);
nor U7485 (N_7485,In_3703,In_867);
nand U7486 (N_7486,In_144,In_1189);
nand U7487 (N_7487,In_4253,In_1521);
and U7488 (N_7488,In_3712,In_4989);
and U7489 (N_7489,In_3655,In_4673);
nor U7490 (N_7490,In_2766,In_1144);
nand U7491 (N_7491,In_2594,In_4760);
xor U7492 (N_7492,In_1508,In_4774);
or U7493 (N_7493,In_4461,In_3770);
nand U7494 (N_7494,In_553,In_600);
nor U7495 (N_7495,In_60,In_4273);
or U7496 (N_7496,In_3043,In_1907);
or U7497 (N_7497,In_3578,In_1825);
nand U7498 (N_7498,In_247,In_1193);
nor U7499 (N_7499,In_603,In_729);
nor U7500 (N_7500,In_1980,In_2502);
nor U7501 (N_7501,In_418,In_703);
nand U7502 (N_7502,In_929,In_2745);
and U7503 (N_7503,In_2114,In_2561);
nor U7504 (N_7504,In_4429,In_693);
nand U7505 (N_7505,In_2087,In_1227);
nand U7506 (N_7506,In_1319,In_3154);
nand U7507 (N_7507,In_3405,In_1029);
nor U7508 (N_7508,In_718,In_3529);
and U7509 (N_7509,In_126,In_1016);
nand U7510 (N_7510,In_3481,In_2662);
nor U7511 (N_7511,In_771,In_3137);
nor U7512 (N_7512,In_3962,In_2993);
nand U7513 (N_7513,In_1240,In_15);
nor U7514 (N_7514,In_3432,In_3262);
nor U7515 (N_7515,In_4527,In_3777);
nor U7516 (N_7516,In_17,In_1173);
xnor U7517 (N_7517,In_111,In_2322);
and U7518 (N_7518,In_2251,In_4133);
or U7519 (N_7519,In_974,In_166);
and U7520 (N_7520,In_2915,In_933);
nand U7521 (N_7521,In_3669,In_2203);
nor U7522 (N_7522,In_3161,In_3624);
or U7523 (N_7523,In_1181,In_768);
nand U7524 (N_7524,In_3603,In_984);
or U7525 (N_7525,In_1986,In_2631);
nor U7526 (N_7526,In_1747,In_2957);
xnor U7527 (N_7527,In_2492,In_2007);
nand U7528 (N_7528,In_34,In_3008);
nor U7529 (N_7529,In_2656,In_4054);
xnor U7530 (N_7530,In_213,In_4401);
nor U7531 (N_7531,In_113,In_3551);
or U7532 (N_7532,In_754,In_1908);
xor U7533 (N_7533,In_1844,In_4259);
nand U7534 (N_7534,In_2589,In_1049);
nor U7535 (N_7535,In_2635,In_4900);
and U7536 (N_7536,In_716,In_2752);
or U7537 (N_7537,In_2550,In_4174);
nor U7538 (N_7538,In_1588,In_2785);
or U7539 (N_7539,In_1208,In_3521);
or U7540 (N_7540,In_2987,In_2315);
nand U7541 (N_7541,In_500,In_489);
or U7542 (N_7542,In_1799,In_1337);
nand U7543 (N_7543,In_357,In_2445);
and U7544 (N_7544,In_4666,In_2908);
nor U7545 (N_7545,In_2585,In_4831);
and U7546 (N_7546,In_677,In_104);
or U7547 (N_7547,In_4610,In_1593);
nor U7548 (N_7548,In_986,In_4438);
and U7549 (N_7549,In_4314,In_2347);
nor U7550 (N_7550,In_2559,In_4330);
nand U7551 (N_7551,In_3015,In_4653);
nand U7552 (N_7552,In_4310,In_4271);
nand U7553 (N_7553,In_2151,In_4454);
or U7554 (N_7554,In_1237,In_4262);
or U7555 (N_7555,In_2684,In_282);
nor U7556 (N_7556,In_3265,In_4553);
nand U7557 (N_7557,In_2677,In_4554);
nor U7558 (N_7558,In_3067,In_4450);
and U7559 (N_7559,In_174,In_2699);
or U7560 (N_7560,In_4179,In_2173);
xnor U7561 (N_7561,In_1346,In_1026);
or U7562 (N_7562,In_1331,In_4579);
nor U7563 (N_7563,In_3560,In_2474);
and U7564 (N_7564,In_3015,In_209);
nor U7565 (N_7565,In_4785,In_1432);
nand U7566 (N_7566,In_2036,In_3504);
nor U7567 (N_7567,In_4044,In_898);
nand U7568 (N_7568,In_3426,In_4875);
and U7569 (N_7569,In_2673,In_4284);
or U7570 (N_7570,In_3425,In_1356);
nor U7571 (N_7571,In_904,In_4681);
and U7572 (N_7572,In_1447,In_3715);
and U7573 (N_7573,In_1536,In_4269);
xnor U7574 (N_7574,In_4450,In_1718);
nor U7575 (N_7575,In_4277,In_1872);
nor U7576 (N_7576,In_3245,In_1402);
and U7577 (N_7577,In_4710,In_3133);
nor U7578 (N_7578,In_3399,In_3950);
nor U7579 (N_7579,In_1640,In_4785);
or U7580 (N_7580,In_2811,In_19);
nand U7581 (N_7581,In_2815,In_2106);
or U7582 (N_7582,In_1733,In_2738);
and U7583 (N_7583,In_2691,In_4000);
nor U7584 (N_7584,In_2600,In_4819);
nand U7585 (N_7585,In_988,In_2937);
or U7586 (N_7586,In_3658,In_3424);
nand U7587 (N_7587,In_296,In_2050);
nand U7588 (N_7588,In_1099,In_598);
and U7589 (N_7589,In_13,In_2071);
nand U7590 (N_7590,In_3959,In_1181);
xor U7591 (N_7591,In_1463,In_3499);
or U7592 (N_7592,In_4418,In_4614);
and U7593 (N_7593,In_3802,In_226);
and U7594 (N_7594,In_4944,In_4854);
or U7595 (N_7595,In_201,In_4902);
nand U7596 (N_7596,In_4235,In_4202);
and U7597 (N_7597,In_365,In_4224);
or U7598 (N_7598,In_3643,In_2406);
xnor U7599 (N_7599,In_1929,In_2980);
nor U7600 (N_7600,In_1492,In_1130);
nand U7601 (N_7601,In_4024,In_4461);
or U7602 (N_7602,In_2803,In_147);
xor U7603 (N_7603,In_4264,In_2134);
nor U7604 (N_7604,In_2140,In_782);
or U7605 (N_7605,In_3279,In_4932);
and U7606 (N_7606,In_1566,In_508);
nor U7607 (N_7607,In_596,In_2007);
nand U7608 (N_7608,In_817,In_3172);
nand U7609 (N_7609,In_165,In_4945);
xor U7610 (N_7610,In_3441,In_3278);
nand U7611 (N_7611,In_90,In_4155);
xor U7612 (N_7612,In_137,In_1051);
nand U7613 (N_7613,In_1564,In_1616);
or U7614 (N_7614,In_2442,In_3570);
or U7615 (N_7615,In_1331,In_3588);
and U7616 (N_7616,In_4008,In_2746);
nand U7617 (N_7617,In_2611,In_4016);
nand U7618 (N_7618,In_1364,In_684);
nor U7619 (N_7619,In_4087,In_4951);
or U7620 (N_7620,In_2120,In_4324);
nand U7621 (N_7621,In_2882,In_2961);
and U7622 (N_7622,In_896,In_4931);
nor U7623 (N_7623,In_4793,In_2752);
nand U7624 (N_7624,In_630,In_2655);
xor U7625 (N_7625,In_3586,In_3556);
xnor U7626 (N_7626,In_207,In_272);
nand U7627 (N_7627,In_2791,In_1966);
nor U7628 (N_7628,In_2370,In_4246);
nand U7629 (N_7629,In_774,In_2739);
nor U7630 (N_7630,In_4375,In_490);
xnor U7631 (N_7631,In_3962,In_3651);
or U7632 (N_7632,In_1062,In_4033);
nor U7633 (N_7633,In_639,In_441);
xnor U7634 (N_7634,In_4217,In_540);
nor U7635 (N_7635,In_4424,In_3488);
and U7636 (N_7636,In_888,In_4961);
nand U7637 (N_7637,In_3610,In_1290);
nor U7638 (N_7638,In_3680,In_1781);
nor U7639 (N_7639,In_275,In_4008);
or U7640 (N_7640,In_759,In_1117);
nor U7641 (N_7641,In_4645,In_1459);
or U7642 (N_7642,In_4323,In_693);
nand U7643 (N_7643,In_170,In_1714);
nand U7644 (N_7644,In_1407,In_3729);
or U7645 (N_7645,In_3829,In_4377);
and U7646 (N_7646,In_697,In_4349);
and U7647 (N_7647,In_2119,In_301);
or U7648 (N_7648,In_1490,In_2893);
xnor U7649 (N_7649,In_3095,In_3666);
or U7650 (N_7650,In_4482,In_4759);
and U7651 (N_7651,In_1253,In_2285);
nand U7652 (N_7652,In_1882,In_4512);
and U7653 (N_7653,In_3525,In_178);
or U7654 (N_7654,In_3262,In_3137);
and U7655 (N_7655,In_1770,In_2462);
xnor U7656 (N_7656,In_1584,In_1497);
nand U7657 (N_7657,In_176,In_1629);
or U7658 (N_7658,In_2451,In_2186);
nand U7659 (N_7659,In_1858,In_3072);
xnor U7660 (N_7660,In_2832,In_1334);
and U7661 (N_7661,In_4997,In_653);
nand U7662 (N_7662,In_1217,In_3702);
nand U7663 (N_7663,In_2665,In_1006);
nand U7664 (N_7664,In_3298,In_2844);
or U7665 (N_7665,In_1074,In_4705);
nor U7666 (N_7666,In_1541,In_2847);
nand U7667 (N_7667,In_4653,In_4157);
and U7668 (N_7668,In_2085,In_884);
nand U7669 (N_7669,In_275,In_3166);
and U7670 (N_7670,In_2361,In_2334);
and U7671 (N_7671,In_3149,In_4755);
or U7672 (N_7672,In_4807,In_3263);
and U7673 (N_7673,In_1723,In_3585);
xor U7674 (N_7674,In_115,In_3776);
nand U7675 (N_7675,In_3883,In_2311);
nor U7676 (N_7676,In_3333,In_2928);
or U7677 (N_7677,In_1161,In_1348);
nand U7678 (N_7678,In_4631,In_4317);
nand U7679 (N_7679,In_2360,In_4591);
nor U7680 (N_7680,In_4105,In_2759);
or U7681 (N_7681,In_3949,In_309);
and U7682 (N_7682,In_1292,In_3053);
xnor U7683 (N_7683,In_3357,In_1863);
and U7684 (N_7684,In_1336,In_4363);
nand U7685 (N_7685,In_735,In_3907);
nor U7686 (N_7686,In_1040,In_4869);
nand U7687 (N_7687,In_2957,In_4161);
and U7688 (N_7688,In_560,In_4990);
nor U7689 (N_7689,In_3243,In_2766);
nand U7690 (N_7690,In_3251,In_4753);
and U7691 (N_7691,In_1247,In_3056);
xor U7692 (N_7692,In_3371,In_4653);
xnor U7693 (N_7693,In_2719,In_1972);
nor U7694 (N_7694,In_3955,In_1641);
and U7695 (N_7695,In_3807,In_479);
nor U7696 (N_7696,In_1357,In_3923);
nand U7697 (N_7697,In_4975,In_4427);
nor U7698 (N_7698,In_3602,In_753);
and U7699 (N_7699,In_536,In_4971);
nor U7700 (N_7700,In_4589,In_4968);
and U7701 (N_7701,In_1856,In_2249);
xnor U7702 (N_7702,In_4460,In_724);
and U7703 (N_7703,In_3632,In_1133);
and U7704 (N_7704,In_3148,In_4633);
nand U7705 (N_7705,In_1340,In_4254);
nand U7706 (N_7706,In_4844,In_284);
nand U7707 (N_7707,In_3284,In_596);
and U7708 (N_7708,In_4117,In_4720);
and U7709 (N_7709,In_635,In_517);
nand U7710 (N_7710,In_4571,In_3464);
nand U7711 (N_7711,In_4860,In_4584);
nand U7712 (N_7712,In_2572,In_1496);
nor U7713 (N_7713,In_1110,In_1940);
nor U7714 (N_7714,In_1505,In_873);
or U7715 (N_7715,In_2142,In_2305);
xor U7716 (N_7716,In_3049,In_3453);
nand U7717 (N_7717,In_2534,In_2667);
and U7718 (N_7718,In_4827,In_3977);
nand U7719 (N_7719,In_4255,In_1736);
and U7720 (N_7720,In_2182,In_4152);
or U7721 (N_7721,In_3931,In_3842);
or U7722 (N_7722,In_2153,In_1778);
or U7723 (N_7723,In_3454,In_4540);
and U7724 (N_7724,In_3918,In_4479);
nand U7725 (N_7725,In_3118,In_1748);
nand U7726 (N_7726,In_1170,In_1559);
and U7727 (N_7727,In_1654,In_4551);
nor U7728 (N_7728,In_2297,In_4451);
nand U7729 (N_7729,In_2416,In_3758);
or U7730 (N_7730,In_2985,In_4736);
and U7731 (N_7731,In_2658,In_2841);
xnor U7732 (N_7732,In_273,In_434);
or U7733 (N_7733,In_1179,In_4786);
or U7734 (N_7734,In_340,In_1289);
nor U7735 (N_7735,In_4850,In_318);
or U7736 (N_7736,In_3723,In_2557);
nor U7737 (N_7737,In_4499,In_1130);
xor U7738 (N_7738,In_2311,In_4637);
and U7739 (N_7739,In_2670,In_3072);
xor U7740 (N_7740,In_576,In_4147);
or U7741 (N_7741,In_2890,In_3249);
or U7742 (N_7742,In_1847,In_3084);
nor U7743 (N_7743,In_1895,In_4967);
and U7744 (N_7744,In_200,In_859);
nand U7745 (N_7745,In_98,In_4459);
nand U7746 (N_7746,In_1399,In_4642);
and U7747 (N_7747,In_3157,In_1774);
nor U7748 (N_7748,In_4956,In_1439);
nand U7749 (N_7749,In_528,In_3200);
xnor U7750 (N_7750,In_2456,In_2958);
nor U7751 (N_7751,In_2072,In_354);
nor U7752 (N_7752,In_371,In_1588);
nor U7753 (N_7753,In_17,In_2805);
nand U7754 (N_7754,In_13,In_1259);
or U7755 (N_7755,In_1133,In_768);
and U7756 (N_7756,In_2866,In_813);
xor U7757 (N_7757,In_1377,In_1161);
or U7758 (N_7758,In_3131,In_2657);
nor U7759 (N_7759,In_3609,In_676);
or U7760 (N_7760,In_2127,In_2539);
nand U7761 (N_7761,In_97,In_496);
and U7762 (N_7762,In_4572,In_3612);
or U7763 (N_7763,In_758,In_3279);
or U7764 (N_7764,In_4370,In_1588);
xnor U7765 (N_7765,In_4469,In_4292);
xnor U7766 (N_7766,In_1427,In_4755);
or U7767 (N_7767,In_2154,In_359);
nor U7768 (N_7768,In_4318,In_953);
and U7769 (N_7769,In_2961,In_2074);
nand U7770 (N_7770,In_2290,In_4529);
nor U7771 (N_7771,In_4358,In_531);
nand U7772 (N_7772,In_1979,In_4695);
nand U7773 (N_7773,In_1635,In_1342);
xor U7774 (N_7774,In_3465,In_934);
and U7775 (N_7775,In_4254,In_310);
xor U7776 (N_7776,In_1449,In_4377);
and U7777 (N_7777,In_863,In_351);
xnor U7778 (N_7778,In_2193,In_415);
nor U7779 (N_7779,In_4564,In_1371);
nor U7780 (N_7780,In_710,In_3220);
nor U7781 (N_7781,In_2827,In_1183);
nor U7782 (N_7782,In_1549,In_2789);
or U7783 (N_7783,In_4479,In_1400);
xnor U7784 (N_7784,In_2718,In_1121);
or U7785 (N_7785,In_4431,In_2141);
and U7786 (N_7786,In_2158,In_2164);
and U7787 (N_7787,In_1009,In_2741);
nor U7788 (N_7788,In_755,In_113);
nand U7789 (N_7789,In_1581,In_1742);
or U7790 (N_7790,In_3658,In_2187);
or U7791 (N_7791,In_1334,In_2263);
nand U7792 (N_7792,In_4206,In_2158);
nand U7793 (N_7793,In_2515,In_4228);
nor U7794 (N_7794,In_791,In_203);
nor U7795 (N_7795,In_2379,In_3909);
nor U7796 (N_7796,In_3138,In_1418);
nand U7797 (N_7797,In_2277,In_3689);
xnor U7798 (N_7798,In_3140,In_3542);
nand U7799 (N_7799,In_4054,In_2856);
and U7800 (N_7800,In_4361,In_2724);
nor U7801 (N_7801,In_4581,In_2528);
nor U7802 (N_7802,In_1289,In_4726);
xor U7803 (N_7803,In_4547,In_2758);
nand U7804 (N_7804,In_3628,In_4062);
or U7805 (N_7805,In_1938,In_1109);
or U7806 (N_7806,In_4898,In_580);
nor U7807 (N_7807,In_92,In_774);
and U7808 (N_7808,In_4596,In_1801);
or U7809 (N_7809,In_1651,In_1230);
or U7810 (N_7810,In_3123,In_4869);
nor U7811 (N_7811,In_1331,In_4008);
or U7812 (N_7812,In_3417,In_4302);
or U7813 (N_7813,In_203,In_667);
xnor U7814 (N_7814,In_11,In_2645);
or U7815 (N_7815,In_1758,In_4969);
xnor U7816 (N_7816,In_4601,In_2021);
or U7817 (N_7817,In_495,In_1835);
nor U7818 (N_7818,In_3231,In_1088);
or U7819 (N_7819,In_2016,In_3926);
nand U7820 (N_7820,In_3827,In_843);
or U7821 (N_7821,In_4418,In_3974);
xnor U7822 (N_7822,In_3423,In_1076);
xor U7823 (N_7823,In_1607,In_2743);
and U7824 (N_7824,In_4824,In_2325);
and U7825 (N_7825,In_424,In_3044);
nor U7826 (N_7826,In_418,In_1764);
or U7827 (N_7827,In_3603,In_2088);
xnor U7828 (N_7828,In_4460,In_1841);
and U7829 (N_7829,In_2047,In_3048);
xnor U7830 (N_7830,In_4225,In_4000);
or U7831 (N_7831,In_3696,In_2752);
and U7832 (N_7832,In_955,In_3797);
nor U7833 (N_7833,In_1336,In_2717);
and U7834 (N_7834,In_3104,In_1367);
xor U7835 (N_7835,In_1456,In_1174);
and U7836 (N_7836,In_2792,In_2411);
nor U7837 (N_7837,In_654,In_740);
nor U7838 (N_7838,In_3603,In_1400);
or U7839 (N_7839,In_3517,In_1654);
nor U7840 (N_7840,In_3107,In_2409);
nand U7841 (N_7841,In_323,In_2976);
nand U7842 (N_7842,In_1349,In_982);
nand U7843 (N_7843,In_2325,In_3946);
or U7844 (N_7844,In_3176,In_3811);
nand U7845 (N_7845,In_2042,In_3586);
and U7846 (N_7846,In_1907,In_231);
nor U7847 (N_7847,In_1297,In_2660);
nor U7848 (N_7848,In_83,In_1611);
or U7849 (N_7849,In_3487,In_4079);
and U7850 (N_7850,In_1008,In_1434);
and U7851 (N_7851,In_3159,In_237);
or U7852 (N_7852,In_1849,In_189);
and U7853 (N_7853,In_476,In_760);
or U7854 (N_7854,In_1115,In_1848);
and U7855 (N_7855,In_2446,In_2339);
and U7856 (N_7856,In_2200,In_2247);
or U7857 (N_7857,In_1220,In_564);
xnor U7858 (N_7858,In_2573,In_3664);
and U7859 (N_7859,In_4996,In_989);
and U7860 (N_7860,In_3793,In_1429);
or U7861 (N_7861,In_4847,In_3738);
nand U7862 (N_7862,In_3148,In_4033);
nand U7863 (N_7863,In_1016,In_4008);
nor U7864 (N_7864,In_1408,In_2347);
nand U7865 (N_7865,In_19,In_147);
nor U7866 (N_7866,In_2295,In_1179);
and U7867 (N_7867,In_182,In_3708);
nand U7868 (N_7868,In_4395,In_1278);
or U7869 (N_7869,In_705,In_3037);
or U7870 (N_7870,In_874,In_2050);
and U7871 (N_7871,In_2953,In_2033);
nand U7872 (N_7872,In_4309,In_3828);
or U7873 (N_7873,In_2253,In_3230);
nor U7874 (N_7874,In_3701,In_4294);
or U7875 (N_7875,In_3613,In_4709);
and U7876 (N_7876,In_3304,In_1709);
xor U7877 (N_7877,In_857,In_2835);
and U7878 (N_7878,In_325,In_3806);
and U7879 (N_7879,In_4845,In_4984);
or U7880 (N_7880,In_2306,In_4054);
xnor U7881 (N_7881,In_582,In_2616);
or U7882 (N_7882,In_1062,In_3775);
and U7883 (N_7883,In_1455,In_2724);
nand U7884 (N_7884,In_817,In_4477);
nand U7885 (N_7885,In_3857,In_3633);
nor U7886 (N_7886,In_1587,In_3620);
and U7887 (N_7887,In_956,In_2806);
xnor U7888 (N_7888,In_4171,In_1573);
nor U7889 (N_7889,In_2577,In_2842);
nor U7890 (N_7890,In_4187,In_2514);
or U7891 (N_7891,In_2318,In_1524);
or U7892 (N_7892,In_4328,In_4456);
and U7893 (N_7893,In_1908,In_3068);
nor U7894 (N_7894,In_4411,In_2019);
or U7895 (N_7895,In_2858,In_2881);
and U7896 (N_7896,In_3844,In_3267);
or U7897 (N_7897,In_2649,In_561);
or U7898 (N_7898,In_2994,In_150);
or U7899 (N_7899,In_3950,In_2296);
nand U7900 (N_7900,In_3378,In_2732);
nand U7901 (N_7901,In_4604,In_1908);
nor U7902 (N_7902,In_616,In_730);
nor U7903 (N_7903,In_4760,In_2191);
and U7904 (N_7904,In_3762,In_3080);
or U7905 (N_7905,In_2225,In_3003);
or U7906 (N_7906,In_482,In_3225);
nand U7907 (N_7907,In_2316,In_637);
nor U7908 (N_7908,In_3716,In_4488);
and U7909 (N_7909,In_4527,In_3954);
nor U7910 (N_7910,In_2906,In_4596);
or U7911 (N_7911,In_1275,In_2308);
nand U7912 (N_7912,In_2642,In_3449);
nand U7913 (N_7913,In_1416,In_1479);
nor U7914 (N_7914,In_3388,In_1235);
or U7915 (N_7915,In_3061,In_3064);
xnor U7916 (N_7916,In_2424,In_2724);
xor U7917 (N_7917,In_2246,In_4023);
or U7918 (N_7918,In_4988,In_211);
and U7919 (N_7919,In_149,In_2577);
xnor U7920 (N_7920,In_1603,In_562);
nand U7921 (N_7921,In_3025,In_4933);
nor U7922 (N_7922,In_3739,In_98);
nor U7923 (N_7923,In_3073,In_2196);
nor U7924 (N_7924,In_2094,In_1310);
xor U7925 (N_7925,In_2180,In_2248);
nor U7926 (N_7926,In_3174,In_3411);
and U7927 (N_7927,In_372,In_2545);
and U7928 (N_7928,In_3908,In_3502);
nand U7929 (N_7929,In_4323,In_531);
or U7930 (N_7930,In_691,In_451);
or U7931 (N_7931,In_2837,In_3620);
nand U7932 (N_7932,In_2013,In_475);
nor U7933 (N_7933,In_1739,In_3703);
nor U7934 (N_7934,In_194,In_2658);
or U7935 (N_7935,In_4072,In_979);
xor U7936 (N_7936,In_1457,In_3301);
and U7937 (N_7937,In_1694,In_4763);
or U7938 (N_7938,In_1614,In_3336);
or U7939 (N_7939,In_147,In_4735);
nand U7940 (N_7940,In_4416,In_1787);
and U7941 (N_7941,In_4458,In_4697);
nand U7942 (N_7942,In_1241,In_2978);
or U7943 (N_7943,In_651,In_532);
and U7944 (N_7944,In_4276,In_446);
nor U7945 (N_7945,In_3819,In_589);
nand U7946 (N_7946,In_3249,In_486);
or U7947 (N_7947,In_691,In_3270);
xnor U7948 (N_7948,In_3978,In_3578);
and U7949 (N_7949,In_2996,In_420);
nand U7950 (N_7950,In_2675,In_4221);
and U7951 (N_7951,In_1363,In_3885);
and U7952 (N_7952,In_714,In_1931);
nor U7953 (N_7953,In_2089,In_4695);
nor U7954 (N_7954,In_21,In_1849);
nor U7955 (N_7955,In_241,In_3010);
nand U7956 (N_7956,In_1612,In_4326);
or U7957 (N_7957,In_2008,In_1336);
and U7958 (N_7958,In_2602,In_2673);
and U7959 (N_7959,In_4364,In_2271);
or U7960 (N_7960,In_4164,In_2831);
and U7961 (N_7961,In_2722,In_625);
and U7962 (N_7962,In_4288,In_3779);
and U7963 (N_7963,In_4816,In_2274);
and U7964 (N_7964,In_4448,In_2972);
nand U7965 (N_7965,In_1558,In_4308);
and U7966 (N_7966,In_743,In_4799);
and U7967 (N_7967,In_2335,In_1838);
nand U7968 (N_7968,In_1628,In_2379);
or U7969 (N_7969,In_4971,In_2642);
nand U7970 (N_7970,In_240,In_2866);
nor U7971 (N_7971,In_2189,In_2263);
xnor U7972 (N_7972,In_1845,In_3229);
xor U7973 (N_7973,In_3027,In_4391);
nand U7974 (N_7974,In_4445,In_75);
or U7975 (N_7975,In_542,In_4521);
nand U7976 (N_7976,In_3928,In_4543);
or U7977 (N_7977,In_1183,In_450);
and U7978 (N_7978,In_3390,In_2865);
or U7979 (N_7979,In_4772,In_3360);
and U7980 (N_7980,In_2578,In_2205);
and U7981 (N_7981,In_3376,In_2262);
nand U7982 (N_7982,In_1789,In_2163);
and U7983 (N_7983,In_725,In_3359);
nand U7984 (N_7984,In_1391,In_2497);
or U7985 (N_7985,In_1550,In_4071);
or U7986 (N_7986,In_738,In_3149);
nand U7987 (N_7987,In_553,In_2785);
or U7988 (N_7988,In_3099,In_785);
or U7989 (N_7989,In_1172,In_4598);
nand U7990 (N_7990,In_2168,In_3270);
nand U7991 (N_7991,In_2894,In_267);
or U7992 (N_7992,In_25,In_940);
nor U7993 (N_7993,In_2837,In_2378);
or U7994 (N_7994,In_1343,In_222);
nand U7995 (N_7995,In_4644,In_2202);
nand U7996 (N_7996,In_804,In_831);
and U7997 (N_7997,In_4712,In_477);
nand U7998 (N_7998,In_803,In_4756);
nand U7999 (N_7999,In_3209,In_3016);
or U8000 (N_8000,In_4088,In_2862);
xor U8001 (N_8001,In_4669,In_4480);
or U8002 (N_8002,In_2760,In_1825);
or U8003 (N_8003,In_255,In_3459);
and U8004 (N_8004,In_3068,In_3901);
nand U8005 (N_8005,In_163,In_1719);
and U8006 (N_8006,In_449,In_4551);
xnor U8007 (N_8007,In_2695,In_92);
or U8008 (N_8008,In_3697,In_4664);
and U8009 (N_8009,In_2303,In_3107);
nor U8010 (N_8010,In_4745,In_1712);
xnor U8011 (N_8011,In_1312,In_4787);
nand U8012 (N_8012,In_609,In_2592);
xnor U8013 (N_8013,In_2804,In_392);
xnor U8014 (N_8014,In_1195,In_10);
or U8015 (N_8015,In_1060,In_2709);
xnor U8016 (N_8016,In_3607,In_1167);
and U8017 (N_8017,In_3183,In_1538);
and U8018 (N_8018,In_2492,In_2729);
nor U8019 (N_8019,In_2853,In_3775);
and U8020 (N_8020,In_4449,In_888);
or U8021 (N_8021,In_1783,In_4824);
nor U8022 (N_8022,In_1052,In_1818);
and U8023 (N_8023,In_1053,In_3458);
nor U8024 (N_8024,In_795,In_4543);
xnor U8025 (N_8025,In_3875,In_735);
nor U8026 (N_8026,In_261,In_1924);
nand U8027 (N_8027,In_1866,In_1244);
or U8028 (N_8028,In_2128,In_1219);
xor U8029 (N_8029,In_2879,In_2988);
xnor U8030 (N_8030,In_3727,In_3099);
xor U8031 (N_8031,In_1947,In_287);
nand U8032 (N_8032,In_3364,In_1783);
and U8033 (N_8033,In_4145,In_3720);
and U8034 (N_8034,In_3524,In_2941);
nor U8035 (N_8035,In_2907,In_635);
or U8036 (N_8036,In_2353,In_3379);
nand U8037 (N_8037,In_1921,In_708);
nor U8038 (N_8038,In_3086,In_4361);
nand U8039 (N_8039,In_2061,In_2506);
nor U8040 (N_8040,In_962,In_942);
nand U8041 (N_8041,In_3071,In_2369);
and U8042 (N_8042,In_130,In_1864);
or U8043 (N_8043,In_4950,In_3887);
and U8044 (N_8044,In_2203,In_4701);
and U8045 (N_8045,In_1317,In_2575);
nand U8046 (N_8046,In_779,In_4195);
nand U8047 (N_8047,In_1869,In_3642);
nor U8048 (N_8048,In_2212,In_646);
nand U8049 (N_8049,In_4844,In_3055);
nand U8050 (N_8050,In_2794,In_1154);
and U8051 (N_8051,In_304,In_2595);
nand U8052 (N_8052,In_2760,In_4579);
or U8053 (N_8053,In_1786,In_4054);
nor U8054 (N_8054,In_4919,In_4826);
or U8055 (N_8055,In_3826,In_1805);
nor U8056 (N_8056,In_3816,In_2925);
or U8057 (N_8057,In_3104,In_3737);
or U8058 (N_8058,In_255,In_1207);
or U8059 (N_8059,In_4203,In_4658);
nor U8060 (N_8060,In_3590,In_61);
nand U8061 (N_8061,In_612,In_1460);
nor U8062 (N_8062,In_1418,In_1369);
or U8063 (N_8063,In_0,In_2360);
nand U8064 (N_8064,In_1519,In_2880);
or U8065 (N_8065,In_284,In_577);
or U8066 (N_8066,In_1608,In_1773);
nor U8067 (N_8067,In_56,In_2176);
nor U8068 (N_8068,In_3918,In_4227);
nand U8069 (N_8069,In_970,In_2545);
nor U8070 (N_8070,In_1971,In_2398);
and U8071 (N_8071,In_2445,In_1327);
and U8072 (N_8072,In_4257,In_4431);
nand U8073 (N_8073,In_3228,In_1883);
or U8074 (N_8074,In_2586,In_3089);
or U8075 (N_8075,In_4459,In_4600);
nand U8076 (N_8076,In_24,In_4879);
or U8077 (N_8077,In_2732,In_3445);
and U8078 (N_8078,In_2828,In_3643);
nor U8079 (N_8079,In_954,In_1131);
xor U8080 (N_8080,In_2768,In_2166);
or U8081 (N_8081,In_623,In_2234);
and U8082 (N_8082,In_1702,In_4196);
nor U8083 (N_8083,In_239,In_2279);
nor U8084 (N_8084,In_513,In_1196);
and U8085 (N_8085,In_1931,In_136);
nor U8086 (N_8086,In_1183,In_300);
and U8087 (N_8087,In_2727,In_157);
or U8088 (N_8088,In_2066,In_4365);
xor U8089 (N_8089,In_3079,In_3404);
nand U8090 (N_8090,In_2768,In_1051);
nor U8091 (N_8091,In_3684,In_1708);
and U8092 (N_8092,In_507,In_4071);
nand U8093 (N_8093,In_4719,In_1231);
nor U8094 (N_8094,In_4754,In_1086);
nand U8095 (N_8095,In_210,In_710);
nand U8096 (N_8096,In_2143,In_965);
and U8097 (N_8097,In_4795,In_1441);
and U8098 (N_8098,In_3443,In_2093);
nor U8099 (N_8099,In_4503,In_1483);
and U8100 (N_8100,In_295,In_4790);
xor U8101 (N_8101,In_1396,In_1659);
or U8102 (N_8102,In_1735,In_2551);
and U8103 (N_8103,In_2868,In_4765);
nand U8104 (N_8104,In_2578,In_2796);
nand U8105 (N_8105,In_3252,In_4869);
nand U8106 (N_8106,In_4312,In_697);
and U8107 (N_8107,In_3905,In_4527);
nor U8108 (N_8108,In_339,In_1212);
and U8109 (N_8109,In_1266,In_1425);
nand U8110 (N_8110,In_2850,In_3474);
nand U8111 (N_8111,In_3192,In_2301);
xor U8112 (N_8112,In_221,In_3223);
and U8113 (N_8113,In_4308,In_240);
and U8114 (N_8114,In_1288,In_397);
or U8115 (N_8115,In_4237,In_700);
or U8116 (N_8116,In_1224,In_789);
nand U8117 (N_8117,In_1922,In_2949);
or U8118 (N_8118,In_1688,In_3090);
or U8119 (N_8119,In_2474,In_1101);
nand U8120 (N_8120,In_298,In_1286);
xor U8121 (N_8121,In_4591,In_1744);
and U8122 (N_8122,In_3781,In_516);
nor U8123 (N_8123,In_3242,In_4665);
nand U8124 (N_8124,In_1733,In_176);
nor U8125 (N_8125,In_3767,In_4857);
or U8126 (N_8126,In_2916,In_996);
nand U8127 (N_8127,In_1934,In_667);
and U8128 (N_8128,In_4549,In_2086);
nand U8129 (N_8129,In_2579,In_2052);
and U8130 (N_8130,In_4109,In_4023);
and U8131 (N_8131,In_501,In_1091);
nor U8132 (N_8132,In_1137,In_3270);
or U8133 (N_8133,In_4635,In_1064);
or U8134 (N_8134,In_4694,In_1787);
nor U8135 (N_8135,In_3356,In_2289);
nor U8136 (N_8136,In_4205,In_2533);
or U8137 (N_8137,In_4482,In_3929);
nand U8138 (N_8138,In_4275,In_4956);
or U8139 (N_8139,In_3466,In_369);
xnor U8140 (N_8140,In_2502,In_1656);
nand U8141 (N_8141,In_4065,In_3974);
or U8142 (N_8142,In_1960,In_3077);
or U8143 (N_8143,In_1036,In_4852);
nand U8144 (N_8144,In_311,In_876);
xor U8145 (N_8145,In_1446,In_1530);
nand U8146 (N_8146,In_2984,In_3830);
and U8147 (N_8147,In_2415,In_1485);
and U8148 (N_8148,In_18,In_4193);
nand U8149 (N_8149,In_1831,In_4571);
nand U8150 (N_8150,In_550,In_3353);
nand U8151 (N_8151,In_3776,In_4609);
nand U8152 (N_8152,In_759,In_178);
and U8153 (N_8153,In_1979,In_4092);
xnor U8154 (N_8154,In_4255,In_4001);
nand U8155 (N_8155,In_2639,In_3263);
nor U8156 (N_8156,In_212,In_4551);
nand U8157 (N_8157,In_4791,In_4141);
nor U8158 (N_8158,In_4321,In_2217);
and U8159 (N_8159,In_2385,In_996);
and U8160 (N_8160,In_251,In_4975);
and U8161 (N_8161,In_4588,In_4577);
xnor U8162 (N_8162,In_3960,In_3191);
nand U8163 (N_8163,In_3964,In_536);
or U8164 (N_8164,In_3160,In_2600);
nor U8165 (N_8165,In_4167,In_2712);
or U8166 (N_8166,In_3209,In_4038);
nor U8167 (N_8167,In_4474,In_27);
xnor U8168 (N_8168,In_1813,In_906);
or U8169 (N_8169,In_3400,In_2804);
and U8170 (N_8170,In_4088,In_2085);
or U8171 (N_8171,In_3192,In_4559);
or U8172 (N_8172,In_3079,In_3437);
or U8173 (N_8173,In_2035,In_238);
nor U8174 (N_8174,In_2649,In_4421);
xnor U8175 (N_8175,In_271,In_3391);
nor U8176 (N_8176,In_4268,In_4972);
nand U8177 (N_8177,In_2140,In_3991);
and U8178 (N_8178,In_3085,In_2112);
nand U8179 (N_8179,In_642,In_3671);
or U8180 (N_8180,In_3443,In_340);
or U8181 (N_8181,In_638,In_2707);
and U8182 (N_8182,In_2580,In_3695);
and U8183 (N_8183,In_1489,In_1808);
nor U8184 (N_8184,In_2939,In_3558);
nor U8185 (N_8185,In_4630,In_816);
nor U8186 (N_8186,In_3745,In_3828);
nand U8187 (N_8187,In_677,In_488);
nand U8188 (N_8188,In_999,In_467);
or U8189 (N_8189,In_1201,In_394);
nand U8190 (N_8190,In_3307,In_1992);
nand U8191 (N_8191,In_198,In_1599);
or U8192 (N_8192,In_153,In_169);
and U8193 (N_8193,In_140,In_3592);
or U8194 (N_8194,In_3814,In_1868);
nand U8195 (N_8195,In_2443,In_3071);
and U8196 (N_8196,In_3252,In_1035);
or U8197 (N_8197,In_2356,In_3069);
nand U8198 (N_8198,In_454,In_2535);
nor U8199 (N_8199,In_3265,In_466);
nand U8200 (N_8200,In_3074,In_2883);
or U8201 (N_8201,In_3320,In_599);
and U8202 (N_8202,In_3344,In_4027);
nor U8203 (N_8203,In_1891,In_233);
or U8204 (N_8204,In_3515,In_2531);
and U8205 (N_8205,In_2800,In_4866);
or U8206 (N_8206,In_1408,In_3175);
and U8207 (N_8207,In_167,In_988);
nand U8208 (N_8208,In_1113,In_886);
xor U8209 (N_8209,In_903,In_3546);
xor U8210 (N_8210,In_3291,In_594);
or U8211 (N_8211,In_1359,In_2073);
nor U8212 (N_8212,In_4333,In_502);
nand U8213 (N_8213,In_2929,In_4580);
nor U8214 (N_8214,In_4787,In_2514);
nand U8215 (N_8215,In_2935,In_1938);
nor U8216 (N_8216,In_2065,In_2144);
or U8217 (N_8217,In_2645,In_428);
or U8218 (N_8218,In_1679,In_1473);
or U8219 (N_8219,In_1702,In_4072);
nor U8220 (N_8220,In_2006,In_3572);
nor U8221 (N_8221,In_4699,In_2587);
or U8222 (N_8222,In_1012,In_3663);
or U8223 (N_8223,In_4431,In_1414);
xor U8224 (N_8224,In_2725,In_1472);
and U8225 (N_8225,In_113,In_2917);
and U8226 (N_8226,In_943,In_4511);
nor U8227 (N_8227,In_1940,In_3216);
or U8228 (N_8228,In_1889,In_4735);
nand U8229 (N_8229,In_3738,In_3963);
nor U8230 (N_8230,In_3696,In_3232);
nand U8231 (N_8231,In_475,In_622);
xor U8232 (N_8232,In_3537,In_3654);
or U8233 (N_8233,In_905,In_1473);
xor U8234 (N_8234,In_1493,In_3617);
and U8235 (N_8235,In_2762,In_1541);
or U8236 (N_8236,In_1116,In_4118);
nand U8237 (N_8237,In_4777,In_1993);
and U8238 (N_8238,In_2472,In_876);
nand U8239 (N_8239,In_2576,In_1121);
nor U8240 (N_8240,In_3692,In_88);
and U8241 (N_8241,In_340,In_2836);
nor U8242 (N_8242,In_1020,In_2182);
nand U8243 (N_8243,In_3355,In_3583);
and U8244 (N_8244,In_1971,In_4858);
nor U8245 (N_8245,In_1705,In_4169);
nand U8246 (N_8246,In_878,In_4623);
and U8247 (N_8247,In_2213,In_368);
nand U8248 (N_8248,In_2498,In_51);
nor U8249 (N_8249,In_3040,In_4074);
nand U8250 (N_8250,In_3946,In_584);
nand U8251 (N_8251,In_3265,In_2040);
nand U8252 (N_8252,In_1479,In_1864);
or U8253 (N_8253,In_3830,In_2182);
or U8254 (N_8254,In_3964,In_1298);
and U8255 (N_8255,In_3142,In_4134);
xnor U8256 (N_8256,In_2329,In_844);
or U8257 (N_8257,In_2690,In_2958);
or U8258 (N_8258,In_927,In_3556);
and U8259 (N_8259,In_4334,In_4591);
xor U8260 (N_8260,In_2894,In_4811);
and U8261 (N_8261,In_3304,In_2291);
nor U8262 (N_8262,In_3881,In_3635);
nand U8263 (N_8263,In_105,In_2512);
nand U8264 (N_8264,In_1915,In_4219);
or U8265 (N_8265,In_2663,In_4480);
nor U8266 (N_8266,In_4066,In_1281);
nand U8267 (N_8267,In_2859,In_3399);
and U8268 (N_8268,In_302,In_1751);
xor U8269 (N_8269,In_1329,In_1980);
or U8270 (N_8270,In_4063,In_576);
nor U8271 (N_8271,In_635,In_2294);
or U8272 (N_8272,In_958,In_1426);
or U8273 (N_8273,In_200,In_3221);
nor U8274 (N_8274,In_3637,In_649);
nor U8275 (N_8275,In_1370,In_3486);
nor U8276 (N_8276,In_1126,In_740);
nor U8277 (N_8277,In_4872,In_4912);
or U8278 (N_8278,In_4518,In_4737);
or U8279 (N_8279,In_2557,In_4138);
nor U8280 (N_8280,In_1990,In_2236);
nor U8281 (N_8281,In_1890,In_679);
nand U8282 (N_8282,In_4137,In_1558);
and U8283 (N_8283,In_162,In_3973);
xor U8284 (N_8284,In_83,In_478);
nor U8285 (N_8285,In_2575,In_2614);
nor U8286 (N_8286,In_3612,In_1154);
or U8287 (N_8287,In_842,In_771);
nand U8288 (N_8288,In_2077,In_3692);
or U8289 (N_8289,In_2858,In_3081);
and U8290 (N_8290,In_621,In_2132);
xnor U8291 (N_8291,In_416,In_1100);
nor U8292 (N_8292,In_2967,In_4666);
or U8293 (N_8293,In_1300,In_290);
and U8294 (N_8294,In_324,In_2372);
nor U8295 (N_8295,In_2749,In_4403);
nand U8296 (N_8296,In_3706,In_2772);
nand U8297 (N_8297,In_4088,In_200);
nor U8298 (N_8298,In_3395,In_4512);
or U8299 (N_8299,In_2243,In_737);
nand U8300 (N_8300,In_4666,In_1441);
nand U8301 (N_8301,In_3247,In_2498);
nor U8302 (N_8302,In_4824,In_1115);
or U8303 (N_8303,In_1507,In_1992);
nor U8304 (N_8304,In_126,In_3561);
and U8305 (N_8305,In_4121,In_1434);
nand U8306 (N_8306,In_3579,In_868);
and U8307 (N_8307,In_2286,In_4419);
nor U8308 (N_8308,In_3643,In_1197);
nor U8309 (N_8309,In_3612,In_537);
xor U8310 (N_8310,In_4973,In_213);
or U8311 (N_8311,In_4336,In_2352);
nand U8312 (N_8312,In_1015,In_3469);
nor U8313 (N_8313,In_3161,In_2099);
nor U8314 (N_8314,In_4004,In_396);
nor U8315 (N_8315,In_3002,In_1384);
nor U8316 (N_8316,In_2399,In_3182);
nor U8317 (N_8317,In_2929,In_1900);
xnor U8318 (N_8318,In_367,In_1577);
nand U8319 (N_8319,In_1042,In_3759);
and U8320 (N_8320,In_445,In_179);
and U8321 (N_8321,In_166,In_519);
nor U8322 (N_8322,In_4818,In_1079);
or U8323 (N_8323,In_1926,In_515);
xor U8324 (N_8324,In_4776,In_918);
or U8325 (N_8325,In_307,In_3187);
and U8326 (N_8326,In_947,In_1164);
nor U8327 (N_8327,In_458,In_4040);
nor U8328 (N_8328,In_4562,In_3802);
nand U8329 (N_8329,In_2664,In_4156);
nor U8330 (N_8330,In_2717,In_3670);
nor U8331 (N_8331,In_1999,In_3557);
xnor U8332 (N_8332,In_4621,In_4459);
and U8333 (N_8333,In_1496,In_2643);
nor U8334 (N_8334,In_3208,In_4412);
or U8335 (N_8335,In_4773,In_1132);
nand U8336 (N_8336,In_3724,In_4246);
nand U8337 (N_8337,In_1493,In_2363);
and U8338 (N_8338,In_1442,In_4745);
nor U8339 (N_8339,In_2188,In_3114);
nor U8340 (N_8340,In_1027,In_1428);
and U8341 (N_8341,In_1624,In_3958);
or U8342 (N_8342,In_3720,In_429);
nor U8343 (N_8343,In_1094,In_167);
and U8344 (N_8344,In_4450,In_1967);
nand U8345 (N_8345,In_541,In_2946);
and U8346 (N_8346,In_2905,In_2037);
nor U8347 (N_8347,In_958,In_4885);
nor U8348 (N_8348,In_3888,In_699);
nor U8349 (N_8349,In_205,In_2841);
nand U8350 (N_8350,In_4806,In_4027);
nor U8351 (N_8351,In_2565,In_1061);
and U8352 (N_8352,In_1416,In_1911);
nor U8353 (N_8353,In_37,In_1138);
nor U8354 (N_8354,In_1132,In_2558);
and U8355 (N_8355,In_2534,In_2652);
and U8356 (N_8356,In_4384,In_2);
nand U8357 (N_8357,In_4195,In_2512);
nor U8358 (N_8358,In_613,In_1421);
and U8359 (N_8359,In_3437,In_4511);
nand U8360 (N_8360,In_985,In_1163);
nand U8361 (N_8361,In_3418,In_4130);
and U8362 (N_8362,In_4078,In_1264);
nor U8363 (N_8363,In_2531,In_1895);
and U8364 (N_8364,In_4850,In_3098);
nor U8365 (N_8365,In_1653,In_1201);
or U8366 (N_8366,In_1102,In_2674);
and U8367 (N_8367,In_1216,In_2474);
or U8368 (N_8368,In_141,In_2883);
or U8369 (N_8369,In_2626,In_3949);
xor U8370 (N_8370,In_1532,In_4183);
xor U8371 (N_8371,In_767,In_2590);
nor U8372 (N_8372,In_3286,In_3953);
or U8373 (N_8373,In_3789,In_4255);
and U8374 (N_8374,In_4633,In_4470);
nand U8375 (N_8375,In_3388,In_2135);
nor U8376 (N_8376,In_2594,In_2595);
xnor U8377 (N_8377,In_2954,In_3658);
nor U8378 (N_8378,In_1017,In_3353);
or U8379 (N_8379,In_4578,In_2919);
and U8380 (N_8380,In_227,In_2986);
nor U8381 (N_8381,In_3573,In_1477);
or U8382 (N_8382,In_3077,In_3929);
and U8383 (N_8383,In_202,In_1482);
and U8384 (N_8384,In_2357,In_2203);
xnor U8385 (N_8385,In_4077,In_3966);
and U8386 (N_8386,In_939,In_1884);
nand U8387 (N_8387,In_2237,In_4764);
nand U8388 (N_8388,In_3421,In_4267);
nand U8389 (N_8389,In_2688,In_4545);
and U8390 (N_8390,In_4336,In_4838);
nor U8391 (N_8391,In_4524,In_4083);
nor U8392 (N_8392,In_2393,In_4072);
and U8393 (N_8393,In_4060,In_2813);
xnor U8394 (N_8394,In_4845,In_1213);
nor U8395 (N_8395,In_3564,In_3565);
or U8396 (N_8396,In_4175,In_3598);
or U8397 (N_8397,In_2911,In_4288);
or U8398 (N_8398,In_547,In_4895);
nand U8399 (N_8399,In_2485,In_4755);
nor U8400 (N_8400,In_1959,In_4149);
and U8401 (N_8401,In_1008,In_3130);
or U8402 (N_8402,In_4051,In_4385);
or U8403 (N_8403,In_1833,In_3986);
xor U8404 (N_8404,In_2289,In_282);
nand U8405 (N_8405,In_2800,In_444);
nor U8406 (N_8406,In_3098,In_1508);
nor U8407 (N_8407,In_1190,In_2372);
nor U8408 (N_8408,In_3914,In_1195);
and U8409 (N_8409,In_3527,In_3707);
or U8410 (N_8410,In_2868,In_1708);
or U8411 (N_8411,In_4875,In_3119);
or U8412 (N_8412,In_70,In_4784);
and U8413 (N_8413,In_3750,In_1684);
nand U8414 (N_8414,In_1572,In_3307);
nand U8415 (N_8415,In_1333,In_1241);
nor U8416 (N_8416,In_1223,In_1750);
and U8417 (N_8417,In_1252,In_811);
xor U8418 (N_8418,In_637,In_2599);
xnor U8419 (N_8419,In_4180,In_325);
or U8420 (N_8420,In_211,In_4438);
or U8421 (N_8421,In_1570,In_4207);
xor U8422 (N_8422,In_495,In_2325);
or U8423 (N_8423,In_3193,In_2729);
and U8424 (N_8424,In_608,In_3255);
nand U8425 (N_8425,In_2142,In_1429);
or U8426 (N_8426,In_1415,In_548);
nor U8427 (N_8427,In_3422,In_605);
nor U8428 (N_8428,In_1510,In_4320);
xor U8429 (N_8429,In_1255,In_4535);
or U8430 (N_8430,In_4438,In_658);
nand U8431 (N_8431,In_92,In_2274);
nand U8432 (N_8432,In_3798,In_3772);
nand U8433 (N_8433,In_2766,In_3000);
nand U8434 (N_8434,In_4250,In_2945);
nor U8435 (N_8435,In_3810,In_3410);
or U8436 (N_8436,In_4404,In_3590);
xnor U8437 (N_8437,In_984,In_2649);
or U8438 (N_8438,In_3484,In_1244);
nor U8439 (N_8439,In_3825,In_606);
or U8440 (N_8440,In_385,In_2055);
xnor U8441 (N_8441,In_4849,In_2258);
nor U8442 (N_8442,In_1176,In_4278);
or U8443 (N_8443,In_2655,In_1345);
nand U8444 (N_8444,In_1397,In_2011);
nor U8445 (N_8445,In_3998,In_734);
xor U8446 (N_8446,In_3727,In_741);
or U8447 (N_8447,In_3144,In_1399);
and U8448 (N_8448,In_3326,In_4796);
or U8449 (N_8449,In_1100,In_3506);
xnor U8450 (N_8450,In_2382,In_1654);
or U8451 (N_8451,In_2934,In_2992);
or U8452 (N_8452,In_2434,In_4451);
nor U8453 (N_8453,In_4209,In_3801);
xor U8454 (N_8454,In_143,In_1824);
nand U8455 (N_8455,In_1293,In_2313);
nand U8456 (N_8456,In_3001,In_513);
xnor U8457 (N_8457,In_3651,In_3881);
and U8458 (N_8458,In_1541,In_1241);
and U8459 (N_8459,In_4951,In_3612);
and U8460 (N_8460,In_2450,In_156);
and U8461 (N_8461,In_4061,In_1403);
nand U8462 (N_8462,In_784,In_2757);
xnor U8463 (N_8463,In_2942,In_2052);
xnor U8464 (N_8464,In_674,In_1313);
and U8465 (N_8465,In_3677,In_4537);
nor U8466 (N_8466,In_987,In_4144);
nand U8467 (N_8467,In_4608,In_356);
nor U8468 (N_8468,In_1550,In_3834);
or U8469 (N_8469,In_754,In_1694);
nor U8470 (N_8470,In_3189,In_733);
nand U8471 (N_8471,In_2039,In_2751);
nor U8472 (N_8472,In_2751,In_2201);
nand U8473 (N_8473,In_4613,In_4922);
or U8474 (N_8474,In_2073,In_4392);
and U8475 (N_8475,In_3541,In_1387);
or U8476 (N_8476,In_4681,In_1261);
or U8477 (N_8477,In_4837,In_3871);
nor U8478 (N_8478,In_1678,In_3515);
or U8479 (N_8479,In_2290,In_3435);
nand U8480 (N_8480,In_516,In_1095);
and U8481 (N_8481,In_1963,In_4391);
xor U8482 (N_8482,In_3989,In_4010);
xnor U8483 (N_8483,In_1804,In_3589);
nand U8484 (N_8484,In_1188,In_4088);
and U8485 (N_8485,In_2644,In_1499);
and U8486 (N_8486,In_2050,In_394);
and U8487 (N_8487,In_3212,In_791);
and U8488 (N_8488,In_1535,In_501);
nand U8489 (N_8489,In_1313,In_1816);
nor U8490 (N_8490,In_42,In_2240);
and U8491 (N_8491,In_4969,In_3813);
nor U8492 (N_8492,In_2879,In_4498);
nand U8493 (N_8493,In_535,In_4715);
nor U8494 (N_8494,In_4387,In_593);
or U8495 (N_8495,In_508,In_4398);
or U8496 (N_8496,In_2,In_4927);
and U8497 (N_8497,In_684,In_4641);
and U8498 (N_8498,In_4940,In_1096);
and U8499 (N_8499,In_430,In_4456);
and U8500 (N_8500,In_3983,In_4184);
nor U8501 (N_8501,In_4631,In_3363);
xor U8502 (N_8502,In_3511,In_2564);
xor U8503 (N_8503,In_2138,In_805);
nand U8504 (N_8504,In_1364,In_4781);
and U8505 (N_8505,In_2637,In_4086);
nand U8506 (N_8506,In_3018,In_440);
nor U8507 (N_8507,In_2748,In_4863);
nor U8508 (N_8508,In_2958,In_1894);
or U8509 (N_8509,In_444,In_4144);
xnor U8510 (N_8510,In_4628,In_2108);
nand U8511 (N_8511,In_604,In_2044);
and U8512 (N_8512,In_1622,In_2484);
or U8513 (N_8513,In_4127,In_40);
or U8514 (N_8514,In_4420,In_3307);
and U8515 (N_8515,In_355,In_1980);
or U8516 (N_8516,In_2072,In_1548);
and U8517 (N_8517,In_1226,In_3546);
nor U8518 (N_8518,In_3325,In_3819);
nand U8519 (N_8519,In_2452,In_4520);
nand U8520 (N_8520,In_3149,In_2611);
xor U8521 (N_8521,In_4418,In_4655);
and U8522 (N_8522,In_4926,In_4852);
or U8523 (N_8523,In_4483,In_4379);
nand U8524 (N_8524,In_549,In_1507);
nand U8525 (N_8525,In_2666,In_1734);
nand U8526 (N_8526,In_4718,In_1479);
nand U8527 (N_8527,In_4548,In_623);
xnor U8528 (N_8528,In_2380,In_110);
nor U8529 (N_8529,In_438,In_2292);
or U8530 (N_8530,In_3580,In_4084);
and U8531 (N_8531,In_4438,In_923);
nand U8532 (N_8532,In_2273,In_2599);
or U8533 (N_8533,In_4679,In_2455);
or U8534 (N_8534,In_1468,In_593);
and U8535 (N_8535,In_4082,In_2830);
xor U8536 (N_8536,In_4486,In_4286);
and U8537 (N_8537,In_2645,In_2719);
or U8538 (N_8538,In_2462,In_3092);
and U8539 (N_8539,In_3570,In_709);
nor U8540 (N_8540,In_2307,In_2826);
nand U8541 (N_8541,In_1577,In_86);
or U8542 (N_8542,In_3648,In_2657);
and U8543 (N_8543,In_4263,In_1931);
and U8544 (N_8544,In_1883,In_4170);
nor U8545 (N_8545,In_842,In_1468);
or U8546 (N_8546,In_4217,In_2175);
nor U8547 (N_8547,In_2310,In_4658);
and U8548 (N_8548,In_977,In_1755);
nand U8549 (N_8549,In_3744,In_62);
nand U8550 (N_8550,In_110,In_4394);
nand U8551 (N_8551,In_2056,In_3321);
nor U8552 (N_8552,In_1751,In_3506);
nor U8553 (N_8553,In_3088,In_2726);
and U8554 (N_8554,In_804,In_2806);
or U8555 (N_8555,In_1148,In_4538);
nand U8556 (N_8556,In_885,In_60);
xnor U8557 (N_8557,In_4348,In_4469);
nor U8558 (N_8558,In_1014,In_4345);
xor U8559 (N_8559,In_335,In_404);
nand U8560 (N_8560,In_2863,In_2966);
or U8561 (N_8561,In_4940,In_701);
and U8562 (N_8562,In_4,In_3890);
nor U8563 (N_8563,In_1213,In_2788);
nor U8564 (N_8564,In_2403,In_4764);
nand U8565 (N_8565,In_2658,In_2429);
nor U8566 (N_8566,In_4662,In_3568);
nand U8567 (N_8567,In_454,In_747);
or U8568 (N_8568,In_2479,In_3611);
xnor U8569 (N_8569,In_345,In_790);
nand U8570 (N_8570,In_2114,In_3523);
nor U8571 (N_8571,In_2022,In_860);
nand U8572 (N_8572,In_3809,In_1016);
nand U8573 (N_8573,In_4745,In_4257);
nor U8574 (N_8574,In_4569,In_368);
nand U8575 (N_8575,In_2840,In_2651);
or U8576 (N_8576,In_729,In_2239);
or U8577 (N_8577,In_328,In_1795);
and U8578 (N_8578,In_1722,In_1647);
or U8579 (N_8579,In_3862,In_1699);
or U8580 (N_8580,In_471,In_2957);
nand U8581 (N_8581,In_141,In_4573);
nand U8582 (N_8582,In_319,In_4080);
nand U8583 (N_8583,In_1732,In_1564);
xor U8584 (N_8584,In_2389,In_4509);
nor U8585 (N_8585,In_3589,In_4000);
or U8586 (N_8586,In_4810,In_4461);
and U8587 (N_8587,In_4296,In_2748);
nor U8588 (N_8588,In_3530,In_1953);
or U8589 (N_8589,In_999,In_3771);
nor U8590 (N_8590,In_1873,In_2842);
nor U8591 (N_8591,In_4900,In_4224);
and U8592 (N_8592,In_413,In_4978);
or U8593 (N_8593,In_1284,In_1341);
and U8594 (N_8594,In_1016,In_3602);
or U8595 (N_8595,In_3398,In_830);
or U8596 (N_8596,In_1909,In_1119);
or U8597 (N_8597,In_534,In_1385);
nor U8598 (N_8598,In_3576,In_3340);
or U8599 (N_8599,In_4080,In_530);
and U8600 (N_8600,In_4171,In_605);
nand U8601 (N_8601,In_1078,In_4290);
and U8602 (N_8602,In_4040,In_3290);
nand U8603 (N_8603,In_642,In_700);
nor U8604 (N_8604,In_1146,In_981);
nor U8605 (N_8605,In_3712,In_2292);
nor U8606 (N_8606,In_4212,In_1414);
xor U8607 (N_8607,In_3917,In_4508);
and U8608 (N_8608,In_1783,In_3069);
and U8609 (N_8609,In_3747,In_550);
nand U8610 (N_8610,In_1542,In_2289);
nand U8611 (N_8611,In_873,In_4076);
nand U8612 (N_8612,In_2580,In_1413);
and U8613 (N_8613,In_4644,In_1905);
or U8614 (N_8614,In_209,In_4373);
nand U8615 (N_8615,In_3123,In_1368);
nor U8616 (N_8616,In_2743,In_761);
nand U8617 (N_8617,In_4794,In_4574);
nand U8618 (N_8618,In_1247,In_3352);
nor U8619 (N_8619,In_1190,In_3668);
and U8620 (N_8620,In_1811,In_1810);
xnor U8621 (N_8621,In_1595,In_3957);
and U8622 (N_8622,In_4593,In_2824);
and U8623 (N_8623,In_2498,In_1419);
nor U8624 (N_8624,In_1583,In_4951);
nor U8625 (N_8625,In_580,In_2867);
nand U8626 (N_8626,In_4812,In_1802);
or U8627 (N_8627,In_2951,In_2414);
nor U8628 (N_8628,In_2831,In_2161);
or U8629 (N_8629,In_525,In_213);
nand U8630 (N_8630,In_56,In_58);
or U8631 (N_8631,In_3059,In_3481);
xor U8632 (N_8632,In_2683,In_410);
and U8633 (N_8633,In_2412,In_1898);
nand U8634 (N_8634,In_2777,In_839);
and U8635 (N_8635,In_4395,In_189);
nand U8636 (N_8636,In_388,In_4772);
nand U8637 (N_8637,In_1347,In_1464);
nand U8638 (N_8638,In_2750,In_1979);
and U8639 (N_8639,In_769,In_2450);
nor U8640 (N_8640,In_4847,In_2981);
nor U8641 (N_8641,In_3133,In_4993);
or U8642 (N_8642,In_113,In_490);
or U8643 (N_8643,In_2628,In_2321);
or U8644 (N_8644,In_88,In_1462);
or U8645 (N_8645,In_4709,In_3456);
and U8646 (N_8646,In_730,In_3037);
or U8647 (N_8647,In_2606,In_2207);
and U8648 (N_8648,In_2855,In_837);
and U8649 (N_8649,In_4718,In_2961);
xnor U8650 (N_8650,In_3118,In_4815);
or U8651 (N_8651,In_3880,In_3001);
nand U8652 (N_8652,In_2435,In_2696);
nand U8653 (N_8653,In_1201,In_2783);
or U8654 (N_8654,In_302,In_1007);
xnor U8655 (N_8655,In_637,In_2079);
and U8656 (N_8656,In_365,In_1857);
nor U8657 (N_8657,In_4868,In_4017);
nor U8658 (N_8658,In_1625,In_1219);
nand U8659 (N_8659,In_2586,In_4701);
and U8660 (N_8660,In_2874,In_2977);
nand U8661 (N_8661,In_2970,In_4472);
nor U8662 (N_8662,In_1444,In_3324);
nor U8663 (N_8663,In_2372,In_277);
nor U8664 (N_8664,In_14,In_1162);
and U8665 (N_8665,In_1323,In_1391);
nor U8666 (N_8666,In_3712,In_3411);
or U8667 (N_8667,In_936,In_1327);
nand U8668 (N_8668,In_1183,In_1014);
and U8669 (N_8669,In_3208,In_2532);
nor U8670 (N_8670,In_3110,In_4556);
or U8671 (N_8671,In_678,In_3883);
or U8672 (N_8672,In_4522,In_1702);
nand U8673 (N_8673,In_1371,In_1738);
nand U8674 (N_8674,In_3547,In_3795);
nand U8675 (N_8675,In_3597,In_2743);
or U8676 (N_8676,In_3752,In_3166);
and U8677 (N_8677,In_4692,In_2060);
or U8678 (N_8678,In_4944,In_3235);
nor U8679 (N_8679,In_4660,In_4359);
nor U8680 (N_8680,In_2528,In_4603);
nor U8681 (N_8681,In_499,In_4807);
nor U8682 (N_8682,In_2240,In_4574);
nand U8683 (N_8683,In_4510,In_3177);
and U8684 (N_8684,In_3837,In_2185);
nor U8685 (N_8685,In_1434,In_4262);
nor U8686 (N_8686,In_4021,In_1813);
nand U8687 (N_8687,In_2639,In_1714);
and U8688 (N_8688,In_103,In_3609);
nor U8689 (N_8689,In_3876,In_1330);
and U8690 (N_8690,In_4663,In_3892);
nand U8691 (N_8691,In_425,In_2605);
and U8692 (N_8692,In_4181,In_2458);
nand U8693 (N_8693,In_4803,In_3039);
xnor U8694 (N_8694,In_1122,In_1336);
or U8695 (N_8695,In_3509,In_4333);
nand U8696 (N_8696,In_1832,In_1741);
and U8697 (N_8697,In_3741,In_2203);
nor U8698 (N_8698,In_1149,In_927);
nand U8699 (N_8699,In_4625,In_1775);
and U8700 (N_8700,In_3540,In_2076);
xnor U8701 (N_8701,In_1736,In_4189);
nor U8702 (N_8702,In_3266,In_2084);
and U8703 (N_8703,In_389,In_3289);
nor U8704 (N_8704,In_3993,In_4525);
or U8705 (N_8705,In_888,In_1623);
or U8706 (N_8706,In_1845,In_4523);
or U8707 (N_8707,In_2735,In_1090);
or U8708 (N_8708,In_4726,In_4513);
nor U8709 (N_8709,In_351,In_3993);
xor U8710 (N_8710,In_1970,In_4978);
and U8711 (N_8711,In_219,In_3791);
nor U8712 (N_8712,In_980,In_419);
nor U8713 (N_8713,In_441,In_3766);
nor U8714 (N_8714,In_4160,In_1938);
nor U8715 (N_8715,In_4786,In_906);
nand U8716 (N_8716,In_1474,In_580);
nand U8717 (N_8717,In_419,In_240);
or U8718 (N_8718,In_3858,In_1511);
nor U8719 (N_8719,In_316,In_4799);
and U8720 (N_8720,In_2920,In_486);
nor U8721 (N_8721,In_2576,In_153);
nand U8722 (N_8722,In_2766,In_2641);
or U8723 (N_8723,In_4764,In_114);
or U8724 (N_8724,In_2788,In_4362);
xnor U8725 (N_8725,In_4376,In_3349);
or U8726 (N_8726,In_226,In_4244);
nor U8727 (N_8727,In_1427,In_1393);
nor U8728 (N_8728,In_84,In_670);
xor U8729 (N_8729,In_4984,In_1795);
nor U8730 (N_8730,In_78,In_2086);
or U8731 (N_8731,In_920,In_1976);
nor U8732 (N_8732,In_2336,In_3535);
nand U8733 (N_8733,In_1476,In_498);
or U8734 (N_8734,In_4364,In_4276);
nor U8735 (N_8735,In_941,In_4835);
nor U8736 (N_8736,In_3942,In_1232);
or U8737 (N_8737,In_1431,In_3701);
nand U8738 (N_8738,In_263,In_4721);
or U8739 (N_8739,In_1279,In_2113);
xor U8740 (N_8740,In_2468,In_2641);
nand U8741 (N_8741,In_4858,In_3477);
nor U8742 (N_8742,In_3793,In_474);
or U8743 (N_8743,In_1436,In_4819);
and U8744 (N_8744,In_1249,In_1170);
and U8745 (N_8745,In_2592,In_4219);
nand U8746 (N_8746,In_420,In_1984);
nor U8747 (N_8747,In_563,In_3144);
nor U8748 (N_8748,In_1681,In_3520);
or U8749 (N_8749,In_4460,In_3669);
and U8750 (N_8750,In_1614,In_3695);
and U8751 (N_8751,In_2459,In_492);
nor U8752 (N_8752,In_3082,In_2053);
or U8753 (N_8753,In_857,In_3012);
nand U8754 (N_8754,In_2098,In_266);
and U8755 (N_8755,In_3508,In_1073);
xnor U8756 (N_8756,In_1579,In_3799);
and U8757 (N_8757,In_2694,In_3004);
or U8758 (N_8758,In_1396,In_2452);
and U8759 (N_8759,In_4759,In_1231);
nor U8760 (N_8760,In_4741,In_4648);
nor U8761 (N_8761,In_60,In_3124);
nor U8762 (N_8762,In_4529,In_1666);
and U8763 (N_8763,In_4503,In_75);
nor U8764 (N_8764,In_3514,In_4222);
or U8765 (N_8765,In_4702,In_4990);
or U8766 (N_8766,In_4244,In_2978);
or U8767 (N_8767,In_1670,In_4944);
xnor U8768 (N_8768,In_1254,In_3795);
nand U8769 (N_8769,In_2505,In_2582);
nand U8770 (N_8770,In_3708,In_3784);
nand U8771 (N_8771,In_2927,In_871);
or U8772 (N_8772,In_317,In_3373);
nor U8773 (N_8773,In_2481,In_4469);
nand U8774 (N_8774,In_21,In_3801);
and U8775 (N_8775,In_3326,In_1153);
nand U8776 (N_8776,In_4100,In_4024);
or U8777 (N_8777,In_4882,In_1820);
and U8778 (N_8778,In_879,In_1627);
nand U8779 (N_8779,In_153,In_4855);
and U8780 (N_8780,In_1479,In_1458);
or U8781 (N_8781,In_4806,In_1433);
xor U8782 (N_8782,In_723,In_2221);
and U8783 (N_8783,In_3087,In_1854);
and U8784 (N_8784,In_4061,In_419);
xor U8785 (N_8785,In_4800,In_314);
and U8786 (N_8786,In_2717,In_2224);
and U8787 (N_8787,In_2478,In_4090);
nor U8788 (N_8788,In_3843,In_3971);
xor U8789 (N_8789,In_2769,In_1613);
nor U8790 (N_8790,In_4507,In_2922);
or U8791 (N_8791,In_63,In_4861);
nand U8792 (N_8792,In_1856,In_3497);
and U8793 (N_8793,In_3522,In_1281);
and U8794 (N_8794,In_3097,In_3658);
or U8795 (N_8795,In_2565,In_1837);
nor U8796 (N_8796,In_1999,In_4460);
and U8797 (N_8797,In_1551,In_2589);
nor U8798 (N_8798,In_4971,In_1253);
or U8799 (N_8799,In_1103,In_4501);
and U8800 (N_8800,In_472,In_3590);
xnor U8801 (N_8801,In_3607,In_4532);
nor U8802 (N_8802,In_197,In_1401);
nand U8803 (N_8803,In_1367,In_591);
or U8804 (N_8804,In_3759,In_856);
or U8805 (N_8805,In_2000,In_531);
and U8806 (N_8806,In_2368,In_2859);
nor U8807 (N_8807,In_2560,In_2518);
and U8808 (N_8808,In_104,In_4451);
nor U8809 (N_8809,In_2065,In_4339);
and U8810 (N_8810,In_279,In_1630);
nand U8811 (N_8811,In_4950,In_2123);
and U8812 (N_8812,In_318,In_4476);
nand U8813 (N_8813,In_972,In_3542);
or U8814 (N_8814,In_1183,In_1097);
or U8815 (N_8815,In_2990,In_4777);
nor U8816 (N_8816,In_2936,In_1094);
nand U8817 (N_8817,In_3015,In_2123);
nor U8818 (N_8818,In_3788,In_3375);
and U8819 (N_8819,In_2935,In_2541);
and U8820 (N_8820,In_3815,In_4213);
nor U8821 (N_8821,In_1205,In_1779);
or U8822 (N_8822,In_3189,In_4115);
and U8823 (N_8823,In_2282,In_1461);
nor U8824 (N_8824,In_2819,In_2657);
nand U8825 (N_8825,In_3790,In_391);
nand U8826 (N_8826,In_100,In_3562);
or U8827 (N_8827,In_4042,In_4568);
or U8828 (N_8828,In_2371,In_1333);
nor U8829 (N_8829,In_1338,In_3173);
or U8830 (N_8830,In_1702,In_981);
nor U8831 (N_8831,In_3188,In_3483);
nand U8832 (N_8832,In_798,In_4442);
nand U8833 (N_8833,In_0,In_2400);
nand U8834 (N_8834,In_4913,In_155);
and U8835 (N_8835,In_3036,In_2270);
nand U8836 (N_8836,In_3468,In_2748);
and U8837 (N_8837,In_2372,In_643);
nor U8838 (N_8838,In_2236,In_3484);
nor U8839 (N_8839,In_4783,In_1977);
xor U8840 (N_8840,In_1487,In_2804);
nor U8841 (N_8841,In_1617,In_3698);
nand U8842 (N_8842,In_1974,In_1202);
nor U8843 (N_8843,In_4170,In_3657);
and U8844 (N_8844,In_4878,In_4019);
or U8845 (N_8845,In_1011,In_3894);
or U8846 (N_8846,In_4702,In_3250);
xor U8847 (N_8847,In_2144,In_4351);
and U8848 (N_8848,In_3356,In_3910);
or U8849 (N_8849,In_3258,In_3861);
nand U8850 (N_8850,In_2716,In_3499);
or U8851 (N_8851,In_3951,In_1512);
nor U8852 (N_8852,In_156,In_121);
nor U8853 (N_8853,In_3405,In_3828);
and U8854 (N_8854,In_3148,In_1187);
and U8855 (N_8855,In_1564,In_1813);
and U8856 (N_8856,In_1698,In_3218);
nor U8857 (N_8857,In_4784,In_1001);
xnor U8858 (N_8858,In_1035,In_2334);
and U8859 (N_8859,In_2095,In_4565);
and U8860 (N_8860,In_4464,In_1179);
nand U8861 (N_8861,In_2235,In_495);
nand U8862 (N_8862,In_4547,In_3329);
xnor U8863 (N_8863,In_1098,In_504);
nand U8864 (N_8864,In_2769,In_2544);
nor U8865 (N_8865,In_292,In_358);
and U8866 (N_8866,In_1775,In_1212);
nor U8867 (N_8867,In_3513,In_3254);
or U8868 (N_8868,In_827,In_4696);
or U8869 (N_8869,In_3193,In_3036);
and U8870 (N_8870,In_97,In_510);
or U8871 (N_8871,In_4348,In_3191);
nand U8872 (N_8872,In_2812,In_1294);
nor U8873 (N_8873,In_245,In_2743);
or U8874 (N_8874,In_4046,In_1122);
nand U8875 (N_8875,In_4855,In_1848);
and U8876 (N_8876,In_322,In_1319);
and U8877 (N_8877,In_2675,In_423);
or U8878 (N_8878,In_3153,In_2727);
and U8879 (N_8879,In_2716,In_4331);
nor U8880 (N_8880,In_4746,In_3208);
nor U8881 (N_8881,In_4697,In_2505);
or U8882 (N_8882,In_1073,In_2640);
and U8883 (N_8883,In_1614,In_859);
nand U8884 (N_8884,In_2573,In_1422);
nor U8885 (N_8885,In_2318,In_3146);
or U8886 (N_8886,In_1960,In_2762);
nor U8887 (N_8887,In_3067,In_1);
nand U8888 (N_8888,In_4638,In_194);
and U8889 (N_8889,In_1507,In_1953);
nand U8890 (N_8890,In_4521,In_997);
nand U8891 (N_8891,In_4237,In_4976);
nand U8892 (N_8892,In_1962,In_455);
xnor U8893 (N_8893,In_3299,In_2279);
nand U8894 (N_8894,In_1511,In_4238);
and U8895 (N_8895,In_528,In_4494);
and U8896 (N_8896,In_1314,In_3637);
or U8897 (N_8897,In_1148,In_4321);
nor U8898 (N_8898,In_396,In_4807);
or U8899 (N_8899,In_2015,In_2372);
xnor U8900 (N_8900,In_3074,In_3321);
and U8901 (N_8901,In_2193,In_4687);
or U8902 (N_8902,In_4852,In_2449);
nand U8903 (N_8903,In_3393,In_327);
nor U8904 (N_8904,In_2738,In_2363);
nor U8905 (N_8905,In_60,In_2536);
and U8906 (N_8906,In_4456,In_39);
nand U8907 (N_8907,In_4579,In_3631);
and U8908 (N_8908,In_3474,In_1758);
nand U8909 (N_8909,In_1651,In_3507);
and U8910 (N_8910,In_2591,In_4469);
xnor U8911 (N_8911,In_1905,In_4525);
and U8912 (N_8912,In_3982,In_2824);
and U8913 (N_8913,In_2737,In_1943);
and U8914 (N_8914,In_3125,In_3893);
nand U8915 (N_8915,In_988,In_1879);
and U8916 (N_8916,In_2531,In_1024);
and U8917 (N_8917,In_234,In_2410);
nand U8918 (N_8918,In_3813,In_40);
and U8919 (N_8919,In_4135,In_3980);
or U8920 (N_8920,In_3669,In_4790);
nor U8921 (N_8921,In_935,In_4059);
nor U8922 (N_8922,In_3486,In_3346);
and U8923 (N_8923,In_4436,In_693);
or U8924 (N_8924,In_1409,In_3416);
and U8925 (N_8925,In_4847,In_479);
xnor U8926 (N_8926,In_4643,In_1570);
or U8927 (N_8927,In_4774,In_4456);
nand U8928 (N_8928,In_2848,In_1265);
nand U8929 (N_8929,In_120,In_3617);
or U8930 (N_8930,In_3317,In_2603);
or U8931 (N_8931,In_3433,In_1031);
xnor U8932 (N_8932,In_1258,In_3215);
or U8933 (N_8933,In_4187,In_2228);
or U8934 (N_8934,In_1315,In_3575);
or U8935 (N_8935,In_3624,In_3589);
and U8936 (N_8936,In_1847,In_2226);
xnor U8937 (N_8937,In_3699,In_1130);
and U8938 (N_8938,In_3279,In_1807);
nand U8939 (N_8939,In_707,In_3370);
nand U8940 (N_8940,In_3847,In_3901);
nor U8941 (N_8941,In_3408,In_3308);
and U8942 (N_8942,In_4592,In_938);
nand U8943 (N_8943,In_2241,In_437);
and U8944 (N_8944,In_3336,In_1195);
or U8945 (N_8945,In_3904,In_360);
nor U8946 (N_8946,In_2226,In_1443);
nor U8947 (N_8947,In_1501,In_3607);
and U8948 (N_8948,In_1215,In_279);
or U8949 (N_8949,In_1142,In_4775);
nor U8950 (N_8950,In_1376,In_1453);
or U8951 (N_8951,In_165,In_2666);
and U8952 (N_8952,In_2086,In_898);
or U8953 (N_8953,In_2964,In_2915);
and U8954 (N_8954,In_2952,In_4492);
xor U8955 (N_8955,In_1058,In_1829);
nand U8956 (N_8956,In_4368,In_2199);
nor U8957 (N_8957,In_1225,In_3591);
nor U8958 (N_8958,In_2884,In_410);
xor U8959 (N_8959,In_586,In_3757);
nor U8960 (N_8960,In_3483,In_4175);
and U8961 (N_8961,In_1395,In_2278);
nor U8962 (N_8962,In_242,In_3249);
or U8963 (N_8963,In_2032,In_4522);
nand U8964 (N_8964,In_1604,In_3823);
or U8965 (N_8965,In_2067,In_3066);
and U8966 (N_8966,In_1562,In_2376);
and U8967 (N_8967,In_4550,In_2917);
or U8968 (N_8968,In_4704,In_3993);
nor U8969 (N_8969,In_3459,In_4012);
xnor U8970 (N_8970,In_1400,In_3465);
or U8971 (N_8971,In_4715,In_3531);
and U8972 (N_8972,In_662,In_1624);
nand U8973 (N_8973,In_4899,In_1359);
xor U8974 (N_8974,In_745,In_4220);
nand U8975 (N_8975,In_985,In_464);
or U8976 (N_8976,In_2919,In_3176);
nand U8977 (N_8977,In_3022,In_4439);
and U8978 (N_8978,In_4958,In_131);
nor U8979 (N_8979,In_7,In_2445);
nor U8980 (N_8980,In_1184,In_1440);
nor U8981 (N_8981,In_1340,In_2005);
and U8982 (N_8982,In_3940,In_2914);
nand U8983 (N_8983,In_3660,In_4176);
or U8984 (N_8984,In_1115,In_3544);
and U8985 (N_8985,In_3957,In_1426);
nor U8986 (N_8986,In_4819,In_411);
and U8987 (N_8987,In_3440,In_3090);
nand U8988 (N_8988,In_2927,In_4556);
and U8989 (N_8989,In_117,In_2851);
nor U8990 (N_8990,In_4770,In_1087);
nand U8991 (N_8991,In_597,In_2301);
or U8992 (N_8992,In_1360,In_4645);
nand U8993 (N_8993,In_2665,In_1574);
or U8994 (N_8994,In_3621,In_2331);
nand U8995 (N_8995,In_1893,In_3227);
nand U8996 (N_8996,In_2670,In_1004);
xnor U8997 (N_8997,In_2104,In_127);
or U8998 (N_8998,In_456,In_4482);
nor U8999 (N_8999,In_794,In_3901);
xor U9000 (N_9000,In_1572,In_2968);
and U9001 (N_9001,In_3399,In_452);
and U9002 (N_9002,In_2699,In_123);
and U9003 (N_9003,In_4062,In_1878);
or U9004 (N_9004,In_2812,In_1712);
and U9005 (N_9005,In_1770,In_2997);
nand U9006 (N_9006,In_417,In_2035);
nand U9007 (N_9007,In_2895,In_3129);
xor U9008 (N_9008,In_2181,In_3535);
nand U9009 (N_9009,In_1200,In_368);
xnor U9010 (N_9010,In_203,In_4908);
xor U9011 (N_9011,In_2191,In_4641);
nand U9012 (N_9012,In_4210,In_2981);
and U9013 (N_9013,In_2455,In_413);
xnor U9014 (N_9014,In_2429,In_1293);
nor U9015 (N_9015,In_4083,In_2184);
and U9016 (N_9016,In_2251,In_454);
xnor U9017 (N_9017,In_4679,In_107);
or U9018 (N_9018,In_4229,In_4049);
nor U9019 (N_9019,In_4108,In_4002);
nor U9020 (N_9020,In_4525,In_489);
nor U9021 (N_9021,In_2493,In_1955);
nand U9022 (N_9022,In_2600,In_2785);
or U9023 (N_9023,In_2051,In_4562);
or U9024 (N_9024,In_556,In_2259);
nand U9025 (N_9025,In_2236,In_1827);
xnor U9026 (N_9026,In_2852,In_4741);
and U9027 (N_9027,In_956,In_4640);
and U9028 (N_9028,In_1327,In_4743);
nand U9029 (N_9029,In_2878,In_1971);
nand U9030 (N_9030,In_338,In_725);
nand U9031 (N_9031,In_3191,In_3317);
and U9032 (N_9032,In_709,In_4203);
xnor U9033 (N_9033,In_1622,In_2556);
or U9034 (N_9034,In_2059,In_2751);
nor U9035 (N_9035,In_3782,In_4848);
nor U9036 (N_9036,In_4729,In_4152);
xor U9037 (N_9037,In_1982,In_1509);
nor U9038 (N_9038,In_3594,In_1128);
nand U9039 (N_9039,In_1719,In_1805);
and U9040 (N_9040,In_4567,In_4407);
nor U9041 (N_9041,In_4162,In_2493);
or U9042 (N_9042,In_2629,In_1007);
or U9043 (N_9043,In_3459,In_4522);
nor U9044 (N_9044,In_3173,In_298);
or U9045 (N_9045,In_2572,In_2069);
nor U9046 (N_9046,In_1685,In_3734);
nor U9047 (N_9047,In_2634,In_318);
nor U9048 (N_9048,In_1418,In_4862);
xor U9049 (N_9049,In_4464,In_1103);
nand U9050 (N_9050,In_4439,In_4744);
and U9051 (N_9051,In_4410,In_4907);
nand U9052 (N_9052,In_3977,In_3934);
and U9053 (N_9053,In_3576,In_2242);
nand U9054 (N_9054,In_3334,In_1541);
or U9055 (N_9055,In_797,In_2671);
or U9056 (N_9056,In_3384,In_4029);
or U9057 (N_9057,In_3457,In_1579);
and U9058 (N_9058,In_3731,In_519);
xor U9059 (N_9059,In_711,In_552);
nor U9060 (N_9060,In_2227,In_4975);
and U9061 (N_9061,In_4012,In_1287);
or U9062 (N_9062,In_818,In_4827);
nor U9063 (N_9063,In_4531,In_3136);
and U9064 (N_9064,In_3354,In_1905);
or U9065 (N_9065,In_2693,In_3754);
and U9066 (N_9066,In_851,In_341);
and U9067 (N_9067,In_2712,In_4908);
and U9068 (N_9068,In_2491,In_3575);
nand U9069 (N_9069,In_1203,In_2599);
nand U9070 (N_9070,In_3496,In_4993);
nor U9071 (N_9071,In_4723,In_2702);
nand U9072 (N_9072,In_4880,In_2609);
nor U9073 (N_9073,In_86,In_2523);
or U9074 (N_9074,In_3614,In_2910);
or U9075 (N_9075,In_2253,In_979);
nand U9076 (N_9076,In_4505,In_2326);
and U9077 (N_9077,In_1130,In_3710);
nand U9078 (N_9078,In_2348,In_1235);
nor U9079 (N_9079,In_2072,In_4480);
nand U9080 (N_9080,In_1425,In_4031);
xor U9081 (N_9081,In_796,In_3160);
nor U9082 (N_9082,In_3820,In_2866);
nor U9083 (N_9083,In_1917,In_1014);
or U9084 (N_9084,In_3479,In_4158);
or U9085 (N_9085,In_874,In_2822);
and U9086 (N_9086,In_4223,In_847);
xor U9087 (N_9087,In_2632,In_1148);
nor U9088 (N_9088,In_1562,In_4958);
or U9089 (N_9089,In_2540,In_1052);
and U9090 (N_9090,In_3014,In_2770);
and U9091 (N_9091,In_3957,In_4361);
nand U9092 (N_9092,In_1313,In_1277);
or U9093 (N_9093,In_4567,In_1218);
and U9094 (N_9094,In_405,In_3339);
and U9095 (N_9095,In_3214,In_2603);
nor U9096 (N_9096,In_801,In_2618);
or U9097 (N_9097,In_3766,In_2625);
nor U9098 (N_9098,In_531,In_1804);
nand U9099 (N_9099,In_4745,In_2489);
or U9100 (N_9100,In_2043,In_4059);
nor U9101 (N_9101,In_3773,In_3656);
or U9102 (N_9102,In_3706,In_2855);
and U9103 (N_9103,In_4470,In_428);
nand U9104 (N_9104,In_1243,In_4452);
or U9105 (N_9105,In_3921,In_4354);
nor U9106 (N_9106,In_739,In_3358);
or U9107 (N_9107,In_1961,In_4300);
or U9108 (N_9108,In_1030,In_1756);
and U9109 (N_9109,In_1943,In_3151);
nand U9110 (N_9110,In_3119,In_2399);
and U9111 (N_9111,In_1378,In_1080);
and U9112 (N_9112,In_3769,In_3216);
or U9113 (N_9113,In_533,In_2971);
or U9114 (N_9114,In_3226,In_4489);
nand U9115 (N_9115,In_4734,In_2761);
or U9116 (N_9116,In_509,In_332);
nor U9117 (N_9117,In_38,In_4536);
and U9118 (N_9118,In_3141,In_513);
xor U9119 (N_9119,In_1978,In_2553);
nand U9120 (N_9120,In_805,In_1570);
and U9121 (N_9121,In_4306,In_3841);
and U9122 (N_9122,In_473,In_3926);
or U9123 (N_9123,In_2238,In_4225);
nand U9124 (N_9124,In_3100,In_124);
or U9125 (N_9125,In_1728,In_2071);
nand U9126 (N_9126,In_1026,In_4625);
or U9127 (N_9127,In_436,In_2114);
nor U9128 (N_9128,In_4850,In_2993);
or U9129 (N_9129,In_1814,In_1729);
or U9130 (N_9130,In_173,In_1449);
xor U9131 (N_9131,In_3279,In_4594);
and U9132 (N_9132,In_765,In_4732);
xnor U9133 (N_9133,In_3618,In_148);
or U9134 (N_9134,In_2779,In_1367);
and U9135 (N_9135,In_1973,In_483);
nor U9136 (N_9136,In_4322,In_1301);
xor U9137 (N_9137,In_3019,In_1000);
nand U9138 (N_9138,In_1384,In_973);
and U9139 (N_9139,In_1180,In_971);
or U9140 (N_9140,In_1963,In_3283);
or U9141 (N_9141,In_2589,In_2909);
or U9142 (N_9142,In_2647,In_3453);
and U9143 (N_9143,In_575,In_649);
or U9144 (N_9144,In_4638,In_2026);
nand U9145 (N_9145,In_2545,In_531);
nor U9146 (N_9146,In_2370,In_4127);
nand U9147 (N_9147,In_1625,In_2341);
xor U9148 (N_9148,In_3413,In_3689);
nand U9149 (N_9149,In_2339,In_1743);
nand U9150 (N_9150,In_299,In_1798);
or U9151 (N_9151,In_619,In_4322);
nor U9152 (N_9152,In_831,In_4592);
or U9153 (N_9153,In_4099,In_2959);
nor U9154 (N_9154,In_104,In_2027);
or U9155 (N_9155,In_126,In_2138);
and U9156 (N_9156,In_3613,In_1486);
xor U9157 (N_9157,In_620,In_3969);
and U9158 (N_9158,In_1429,In_2050);
nor U9159 (N_9159,In_3087,In_2178);
or U9160 (N_9160,In_2695,In_3286);
nand U9161 (N_9161,In_4787,In_3498);
nand U9162 (N_9162,In_306,In_384);
or U9163 (N_9163,In_630,In_3570);
or U9164 (N_9164,In_2137,In_138);
xnor U9165 (N_9165,In_2296,In_1609);
or U9166 (N_9166,In_1870,In_2680);
nor U9167 (N_9167,In_3330,In_898);
and U9168 (N_9168,In_4865,In_3830);
nor U9169 (N_9169,In_3235,In_2404);
or U9170 (N_9170,In_4831,In_1610);
and U9171 (N_9171,In_1716,In_1904);
and U9172 (N_9172,In_2951,In_373);
xnor U9173 (N_9173,In_1179,In_4343);
and U9174 (N_9174,In_2762,In_344);
nor U9175 (N_9175,In_1025,In_1374);
nor U9176 (N_9176,In_4773,In_4818);
xnor U9177 (N_9177,In_1906,In_4097);
and U9178 (N_9178,In_4458,In_2421);
and U9179 (N_9179,In_313,In_4);
and U9180 (N_9180,In_4760,In_2233);
nand U9181 (N_9181,In_686,In_3986);
xor U9182 (N_9182,In_2953,In_4055);
xor U9183 (N_9183,In_66,In_3116);
or U9184 (N_9184,In_2336,In_736);
nand U9185 (N_9185,In_3,In_4586);
nor U9186 (N_9186,In_4303,In_283);
nor U9187 (N_9187,In_582,In_3058);
nor U9188 (N_9188,In_2,In_4072);
or U9189 (N_9189,In_1700,In_4699);
nand U9190 (N_9190,In_1702,In_3935);
nand U9191 (N_9191,In_1239,In_4232);
nor U9192 (N_9192,In_1944,In_4720);
nand U9193 (N_9193,In_4118,In_4777);
nor U9194 (N_9194,In_3578,In_3401);
nor U9195 (N_9195,In_3962,In_2547);
nor U9196 (N_9196,In_2484,In_316);
nand U9197 (N_9197,In_2525,In_1477);
nand U9198 (N_9198,In_3216,In_3018);
xor U9199 (N_9199,In_979,In_365);
or U9200 (N_9200,In_2318,In_1880);
and U9201 (N_9201,In_777,In_3813);
xor U9202 (N_9202,In_372,In_1690);
or U9203 (N_9203,In_333,In_1233);
or U9204 (N_9204,In_3981,In_2915);
nand U9205 (N_9205,In_2862,In_4159);
xor U9206 (N_9206,In_1055,In_2181);
and U9207 (N_9207,In_1702,In_1689);
nor U9208 (N_9208,In_3303,In_1880);
or U9209 (N_9209,In_4727,In_3820);
nand U9210 (N_9210,In_4671,In_4492);
or U9211 (N_9211,In_3854,In_2760);
and U9212 (N_9212,In_504,In_1302);
nand U9213 (N_9213,In_2383,In_2071);
or U9214 (N_9214,In_2912,In_4677);
nor U9215 (N_9215,In_2916,In_1613);
or U9216 (N_9216,In_2114,In_943);
nor U9217 (N_9217,In_2096,In_4882);
and U9218 (N_9218,In_2988,In_3511);
xor U9219 (N_9219,In_4996,In_2805);
and U9220 (N_9220,In_2479,In_4283);
and U9221 (N_9221,In_205,In_3226);
nand U9222 (N_9222,In_3646,In_1043);
or U9223 (N_9223,In_2830,In_1069);
nand U9224 (N_9224,In_1783,In_469);
nor U9225 (N_9225,In_3136,In_4283);
or U9226 (N_9226,In_1854,In_1542);
nor U9227 (N_9227,In_3141,In_1470);
nor U9228 (N_9228,In_3917,In_2680);
nand U9229 (N_9229,In_2909,In_706);
and U9230 (N_9230,In_3798,In_1645);
nand U9231 (N_9231,In_4174,In_4362);
and U9232 (N_9232,In_364,In_1066);
nor U9233 (N_9233,In_1118,In_4722);
and U9234 (N_9234,In_3822,In_3017);
or U9235 (N_9235,In_2033,In_4323);
nand U9236 (N_9236,In_3648,In_1213);
nand U9237 (N_9237,In_2937,In_1629);
and U9238 (N_9238,In_2622,In_2819);
nand U9239 (N_9239,In_1015,In_4252);
or U9240 (N_9240,In_3127,In_1567);
or U9241 (N_9241,In_117,In_2488);
and U9242 (N_9242,In_1927,In_3858);
nor U9243 (N_9243,In_565,In_591);
nor U9244 (N_9244,In_3281,In_2409);
nand U9245 (N_9245,In_1010,In_908);
or U9246 (N_9246,In_1477,In_2116);
or U9247 (N_9247,In_3466,In_3698);
and U9248 (N_9248,In_390,In_96);
nand U9249 (N_9249,In_4570,In_3199);
or U9250 (N_9250,In_16,In_4755);
and U9251 (N_9251,In_2692,In_2780);
and U9252 (N_9252,In_2473,In_4733);
or U9253 (N_9253,In_100,In_1657);
nand U9254 (N_9254,In_1636,In_834);
or U9255 (N_9255,In_3923,In_1317);
nor U9256 (N_9256,In_2541,In_191);
nand U9257 (N_9257,In_2873,In_2912);
or U9258 (N_9258,In_1607,In_145);
nor U9259 (N_9259,In_254,In_2435);
xnor U9260 (N_9260,In_4297,In_2082);
and U9261 (N_9261,In_3559,In_3628);
or U9262 (N_9262,In_4565,In_1909);
or U9263 (N_9263,In_159,In_1214);
or U9264 (N_9264,In_1618,In_4495);
nand U9265 (N_9265,In_3842,In_4929);
or U9266 (N_9266,In_4807,In_4926);
or U9267 (N_9267,In_1501,In_2436);
nand U9268 (N_9268,In_794,In_1002);
nand U9269 (N_9269,In_2958,In_4890);
or U9270 (N_9270,In_2167,In_1802);
xor U9271 (N_9271,In_1314,In_3444);
nand U9272 (N_9272,In_4894,In_3787);
nor U9273 (N_9273,In_95,In_668);
or U9274 (N_9274,In_3130,In_1912);
nand U9275 (N_9275,In_3173,In_3965);
and U9276 (N_9276,In_1975,In_4553);
or U9277 (N_9277,In_2527,In_3073);
nor U9278 (N_9278,In_1685,In_1151);
nor U9279 (N_9279,In_1141,In_115);
or U9280 (N_9280,In_4058,In_2443);
xnor U9281 (N_9281,In_4369,In_2162);
xor U9282 (N_9282,In_795,In_321);
nand U9283 (N_9283,In_4900,In_772);
and U9284 (N_9284,In_2117,In_3654);
or U9285 (N_9285,In_1077,In_3454);
or U9286 (N_9286,In_930,In_4741);
and U9287 (N_9287,In_2616,In_1620);
and U9288 (N_9288,In_3793,In_102);
nand U9289 (N_9289,In_3951,In_4381);
and U9290 (N_9290,In_1300,In_2595);
or U9291 (N_9291,In_2577,In_1361);
xnor U9292 (N_9292,In_1037,In_3070);
nand U9293 (N_9293,In_1624,In_4059);
xor U9294 (N_9294,In_1841,In_3318);
and U9295 (N_9295,In_1561,In_1595);
and U9296 (N_9296,In_4495,In_4303);
and U9297 (N_9297,In_919,In_2489);
or U9298 (N_9298,In_821,In_2969);
and U9299 (N_9299,In_305,In_4340);
or U9300 (N_9300,In_3848,In_2467);
xor U9301 (N_9301,In_3004,In_2407);
nand U9302 (N_9302,In_2254,In_2496);
or U9303 (N_9303,In_3491,In_4635);
nor U9304 (N_9304,In_1083,In_1890);
and U9305 (N_9305,In_4510,In_1475);
or U9306 (N_9306,In_4360,In_4983);
or U9307 (N_9307,In_1961,In_1307);
and U9308 (N_9308,In_1296,In_4845);
xor U9309 (N_9309,In_3099,In_1805);
or U9310 (N_9310,In_2334,In_3108);
nand U9311 (N_9311,In_2635,In_3114);
or U9312 (N_9312,In_4900,In_903);
or U9313 (N_9313,In_4210,In_3207);
nand U9314 (N_9314,In_3159,In_2749);
and U9315 (N_9315,In_4160,In_1649);
and U9316 (N_9316,In_4732,In_1763);
and U9317 (N_9317,In_719,In_2890);
nor U9318 (N_9318,In_471,In_334);
or U9319 (N_9319,In_1740,In_1829);
nand U9320 (N_9320,In_2609,In_3814);
xor U9321 (N_9321,In_3712,In_1812);
or U9322 (N_9322,In_4851,In_3478);
nor U9323 (N_9323,In_2505,In_3688);
nand U9324 (N_9324,In_1663,In_108);
and U9325 (N_9325,In_4916,In_3757);
and U9326 (N_9326,In_1163,In_232);
xor U9327 (N_9327,In_1557,In_4163);
nor U9328 (N_9328,In_2575,In_1010);
nand U9329 (N_9329,In_1378,In_2756);
or U9330 (N_9330,In_957,In_1501);
or U9331 (N_9331,In_1939,In_1231);
nand U9332 (N_9332,In_810,In_2372);
xnor U9333 (N_9333,In_3527,In_2724);
or U9334 (N_9334,In_1268,In_3596);
nor U9335 (N_9335,In_4922,In_1515);
or U9336 (N_9336,In_1738,In_3223);
nor U9337 (N_9337,In_3445,In_3983);
xor U9338 (N_9338,In_2662,In_2992);
nand U9339 (N_9339,In_2058,In_2029);
and U9340 (N_9340,In_2739,In_1481);
and U9341 (N_9341,In_4139,In_2496);
nand U9342 (N_9342,In_4288,In_3381);
nand U9343 (N_9343,In_3015,In_4547);
nor U9344 (N_9344,In_2051,In_1169);
and U9345 (N_9345,In_2507,In_2176);
nand U9346 (N_9346,In_3222,In_1891);
or U9347 (N_9347,In_803,In_70);
and U9348 (N_9348,In_4533,In_402);
nor U9349 (N_9349,In_1275,In_2354);
or U9350 (N_9350,In_1478,In_3907);
nand U9351 (N_9351,In_4449,In_787);
nand U9352 (N_9352,In_1415,In_935);
or U9353 (N_9353,In_4319,In_1953);
xnor U9354 (N_9354,In_1815,In_4231);
nor U9355 (N_9355,In_2377,In_149);
and U9356 (N_9356,In_2721,In_2173);
or U9357 (N_9357,In_553,In_2452);
nor U9358 (N_9358,In_2194,In_1347);
nand U9359 (N_9359,In_1858,In_4689);
nand U9360 (N_9360,In_4939,In_4594);
and U9361 (N_9361,In_4655,In_312);
nand U9362 (N_9362,In_4662,In_4032);
nor U9363 (N_9363,In_15,In_458);
xnor U9364 (N_9364,In_690,In_3846);
xnor U9365 (N_9365,In_419,In_992);
nor U9366 (N_9366,In_540,In_1085);
nor U9367 (N_9367,In_1223,In_941);
and U9368 (N_9368,In_1871,In_3242);
nor U9369 (N_9369,In_387,In_3531);
or U9370 (N_9370,In_3315,In_4105);
xnor U9371 (N_9371,In_139,In_89);
nor U9372 (N_9372,In_2002,In_3082);
nor U9373 (N_9373,In_4867,In_3339);
nand U9374 (N_9374,In_1047,In_989);
and U9375 (N_9375,In_214,In_2888);
and U9376 (N_9376,In_2715,In_2434);
nor U9377 (N_9377,In_4004,In_2401);
nor U9378 (N_9378,In_1015,In_3945);
nor U9379 (N_9379,In_2407,In_2311);
nor U9380 (N_9380,In_4545,In_2946);
nand U9381 (N_9381,In_4769,In_2109);
nor U9382 (N_9382,In_1036,In_3974);
or U9383 (N_9383,In_1949,In_3151);
nand U9384 (N_9384,In_2683,In_807);
or U9385 (N_9385,In_3697,In_603);
or U9386 (N_9386,In_2630,In_4319);
or U9387 (N_9387,In_2326,In_1042);
or U9388 (N_9388,In_4744,In_3757);
or U9389 (N_9389,In_2595,In_2973);
and U9390 (N_9390,In_4778,In_2016);
and U9391 (N_9391,In_2865,In_3443);
xnor U9392 (N_9392,In_1982,In_489);
xor U9393 (N_9393,In_2537,In_2631);
nand U9394 (N_9394,In_3452,In_4304);
nand U9395 (N_9395,In_3492,In_641);
nor U9396 (N_9396,In_4966,In_4786);
xnor U9397 (N_9397,In_3683,In_2845);
or U9398 (N_9398,In_25,In_3264);
and U9399 (N_9399,In_1718,In_1413);
nand U9400 (N_9400,In_1109,In_1340);
nand U9401 (N_9401,In_3949,In_3086);
and U9402 (N_9402,In_1875,In_878);
and U9403 (N_9403,In_77,In_443);
or U9404 (N_9404,In_3603,In_3853);
nand U9405 (N_9405,In_1704,In_305);
or U9406 (N_9406,In_4137,In_1109);
nor U9407 (N_9407,In_3247,In_1016);
and U9408 (N_9408,In_4094,In_769);
nand U9409 (N_9409,In_682,In_1776);
and U9410 (N_9410,In_539,In_2328);
nor U9411 (N_9411,In_4290,In_2159);
and U9412 (N_9412,In_3977,In_3478);
nor U9413 (N_9413,In_2756,In_2560);
nor U9414 (N_9414,In_4461,In_262);
and U9415 (N_9415,In_4709,In_654);
and U9416 (N_9416,In_1560,In_3017);
nor U9417 (N_9417,In_1880,In_4681);
nand U9418 (N_9418,In_58,In_4080);
nor U9419 (N_9419,In_874,In_1024);
and U9420 (N_9420,In_3919,In_3038);
or U9421 (N_9421,In_2527,In_346);
and U9422 (N_9422,In_3704,In_2927);
nor U9423 (N_9423,In_1012,In_3385);
nor U9424 (N_9424,In_3285,In_1019);
and U9425 (N_9425,In_1668,In_1915);
nand U9426 (N_9426,In_3272,In_3138);
nor U9427 (N_9427,In_1455,In_2561);
nand U9428 (N_9428,In_1174,In_1856);
nor U9429 (N_9429,In_643,In_4988);
and U9430 (N_9430,In_4312,In_4296);
nand U9431 (N_9431,In_3437,In_1153);
nand U9432 (N_9432,In_1894,In_2496);
nor U9433 (N_9433,In_353,In_1273);
or U9434 (N_9434,In_5,In_1180);
nor U9435 (N_9435,In_2868,In_791);
nand U9436 (N_9436,In_3054,In_1754);
or U9437 (N_9437,In_2573,In_1022);
nand U9438 (N_9438,In_3003,In_2332);
or U9439 (N_9439,In_2692,In_334);
nand U9440 (N_9440,In_4435,In_808);
xor U9441 (N_9441,In_2270,In_210);
nand U9442 (N_9442,In_3931,In_75);
xnor U9443 (N_9443,In_422,In_4993);
and U9444 (N_9444,In_1204,In_4398);
xor U9445 (N_9445,In_1892,In_1112);
and U9446 (N_9446,In_2545,In_3083);
and U9447 (N_9447,In_4397,In_2163);
and U9448 (N_9448,In_4645,In_4797);
nand U9449 (N_9449,In_4668,In_236);
xnor U9450 (N_9450,In_1892,In_763);
or U9451 (N_9451,In_2671,In_45);
or U9452 (N_9452,In_4811,In_2238);
nor U9453 (N_9453,In_4579,In_159);
nor U9454 (N_9454,In_1105,In_1895);
nand U9455 (N_9455,In_2402,In_3816);
nor U9456 (N_9456,In_695,In_3108);
nor U9457 (N_9457,In_2214,In_4054);
and U9458 (N_9458,In_1741,In_332);
nor U9459 (N_9459,In_4405,In_3302);
nand U9460 (N_9460,In_4931,In_555);
xnor U9461 (N_9461,In_1020,In_1491);
xnor U9462 (N_9462,In_2056,In_3407);
xor U9463 (N_9463,In_1991,In_2834);
nor U9464 (N_9464,In_1879,In_1902);
and U9465 (N_9465,In_465,In_2277);
and U9466 (N_9466,In_4884,In_3413);
xor U9467 (N_9467,In_2974,In_2921);
and U9468 (N_9468,In_639,In_3777);
or U9469 (N_9469,In_713,In_1567);
nor U9470 (N_9470,In_241,In_2522);
xor U9471 (N_9471,In_2508,In_151);
or U9472 (N_9472,In_883,In_1932);
nand U9473 (N_9473,In_1440,In_1533);
and U9474 (N_9474,In_2089,In_2455);
and U9475 (N_9475,In_4721,In_2240);
or U9476 (N_9476,In_1747,In_1147);
nand U9477 (N_9477,In_1059,In_2744);
and U9478 (N_9478,In_4922,In_4039);
nand U9479 (N_9479,In_2666,In_1221);
or U9480 (N_9480,In_660,In_2812);
nand U9481 (N_9481,In_4499,In_4713);
nand U9482 (N_9482,In_1279,In_1686);
or U9483 (N_9483,In_273,In_3336);
and U9484 (N_9484,In_123,In_2560);
nand U9485 (N_9485,In_593,In_1333);
nand U9486 (N_9486,In_641,In_3534);
nor U9487 (N_9487,In_4581,In_2685);
or U9488 (N_9488,In_4712,In_700);
nand U9489 (N_9489,In_332,In_423);
nor U9490 (N_9490,In_3257,In_1022);
and U9491 (N_9491,In_4204,In_3330);
nand U9492 (N_9492,In_4061,In_4531);
xor U9493 (N_9493,In_2875,In_3676);
and U9494 (N_9494,In_4752,In_2917);
nand U9495 (N_9495,In_1259,In_4195);
nand U9496 (N_9496,In_481,In_4162);
and U9497 (N_9497,In_2110,In_235);
or U9498 (N_9498,In_3043,In_2094);
and U9499 (N_9499,In_2757,In_2593);
nor U9500 (N_9500,In_4520,In_2967);
nor U9501 (N_9501,In_2837,In_2277);
nand U9502 (N_9502,In_590,In_4698);
or U9503 (N_9503,In_4871,In_4590);
xor U9504 (N_9504,In_3033,In_3064);
nand U9505 (N_9505,In_4764,In_2553);
xor U9506 (N_9506,In_2762,In_690);
nor U9507 (N_9507,In_4177,In_4423);
nor U9508 (N_9508,In_3546,In_2781);
nor U9509 (N_9509,In_171,In_4499);
nand U9510 (N_9510,In_1279,In_1344);
or U9511 (N_9511,In_3089,In_3944);
nor U9512 (N_9512,In_2998,In_3471);
nor U9513 (N_9513,In_2950,In_2538);
and U9514 (N_9514,In_3093,In_3536);
nor U9515 (N_9515,In_20,In_2716);
and U9516 (N_9516,In_4254,In_407);
or U9517 (N_9517,In_3598,In_3635);
or U9518 (N_9518,In_2016,In_4211);
nand U9519 (N_9519,In_4698,In_2789);
or U9520 (N_9520,In_318,In_3195);
and U9521 (N_9521,In_266,In_39);
and U9522 (N_9522,In_2122,In_2362);
xor U9523 (N_9523,In_4059,In_2820);
xnor U9524 (N_9524,In_1078,In_2512);
nor U9525 (N_9525,In_1509,In_1634);
or U9526 (N_9526,In_3600,In_1064);
and U9527 (N_9527,In_40,In_2451);
xnor U9528 (N_9528,In_4812,In_2026);
nor U9529 (N_9529,In_1298,In_3340);
nand U9530 (N_9530,In_4487,In_4311);
and U9531 (N_9531,In_2118,In_3211);
or U9532 (N_9532,In_806,In_2370);
and U9533 (N_9533,In_4645,In_4362);
xor U9534 (N_9534,In_1369,In_1573);
nand U9535 (N_9535,In_405,In_87);
and U9536 (N_9536,In_4361,In_1575);
and U9537 (N_9537,In_1113,In_1475);
and U9538 (N_9538,In_4384,In_887);
nand U9539 (N_9539,In_4068,In_3058);
nand U9540 (N_9540,In_2990,In_3921);
and U9541 (N_9541,In_4391,In_3611);
nand U9542 (N_9542,In_1318,In_1313);
and U9543 (N_9543,In_319,In_4457);
nor U9544 (N_9544,In_2506,In_2263);
nand U9545 (N_9545,In_4733,In_3605);
nand U9546 (N_9546,In_920,In_1107);
and U9547 (N_9547,In_576,In_4488);
xor U9548 (N_9548,In_1373,In_4071);
and U9549 (N_9549,In_3958,In_336);
and U9550 (N_9550,In_4554,In_3041);
nand U9551 (N_9551,In_4615,In_2667);
nor U9552 (N_9552,In_4892,In_223);
or U9553 (N_9553,In_531,In_1326);
nand U9554 (N_9554,In_2863,In_2152);
or U9555 (N_9555,In_4951,In_3036);
and U9556 (N_9556,In_3349,In_4556);
nand U9557 (N_9557,In_4836,In_776);
xnor U9558 (N_9558,In_1205,In_2022);
or U9559 (N_9559,In_1607,In_3465);
or U9560 (N_9560,In_4096,In_2309);
nand U9561 (N_9561,In_4306,In_3080);
nor U9562 (N_9562,In_1873,In_283);
and U9563 (N_9563,In_4241,In_4521);
nor U9564 (N_9564,In_2515,In_1463);
and U9565 (N_9565,In_2228,In_2963);
or U9566 (N_9566,In_4855,In_1398);
nand U9567 (N_9567,In_4024,In_4044);
nor U9568 (N_9568,In_1415,In_3268);
nor U9569 (N_9569,In_952,In_1593);
or U9570 (N_9570,In_3747,In_4758);
xnor U9571 (N_9571,In_2646,In_2359);
or U9572 (N_9572,In_3546,In_1935);
nor U9573 (N_9573,In_4156,In_4619);
or U9574 (N_9574,In_716,In_3976);
nor U9575 (N_9575,In_780,In_150);
or U9576 (N_9576,In_1957,In_1034);
nor U9577 (N_9577,In_4682,In_2016);
nor U9578 (N_9578,In_2535,In_2397);
nand U9579 (N_9579,In_835,In_3450);
xor U9580 (N_9580,In_4022,In_2356);
nand U9581 (N_9581,In_381,In_4788);
or U9582 (N_9582,In_4889,In_2186);
nand U9583 (N_9583,In_2260,In_3936);
and U9584 (N_9584,In_2324,In_950);
nand U9585 (N_9585,In_3121,In_4329);
nor U9586 (N_9586,In_4461,In_628);
and U9587 (N_9587,In_2761,In_601);
and U9588 (N_9588,In_1504,In_3815);
nand U9589 (N_9589,In_222,In_2837);
nand U9590 (N_9590,In_2433,In_4679);
xnor U9591 (N_9591,In_1281,In_3621);
nand U9592 (N_9592,In_429,In_4890);
nor U9593 (N_9593,In_4147,In_2155);
and U9594 (N_9594,In_3632,In_4028);
and U9595 (N_9595,In_2455,In_3810);
nand U9596 (N_9596,In_3453,In_1483);
nand U9597 (N_9597,In_1228,In_4684);
nor U9598 (N_9598,In_2987,In_3608);
nor U9599 (N_9599,In_187,In_3975);
and U9600 (N_9600,In_1918,In_4494);
nand U9601 (N_9601,In_2730,In_454);
nand U9602 (N_9602,In_3126,In_430);
and U9603 (N_9603,In_1104,In_323);
and U9604 (N_9604,In_254,In_2227);
or U9605 (N_9605,In_1801,In_2822);
nor U9606 (N_9606,In_4726,In_134);
and U9607 (N_9607,In_1321,In_3877);
or U9608 (N_9608,In_1745,In_244);
nor U9609 (N_9609,In_3070,In_2745);
nand U9610 (N_9610,In_530,In_2667);
nor U9611 (N_9611,In_426,In_1597);
nand U9612 (N_9612,In_1040,In_663);
nand U9613 (N_9613,In_2037,In_3698);
and U9614 (N_9614,In_2124,In_163);
and U9615 (N_9615,In_4500,In_1605);
nor U9616 (N_9616,In_4672,In_1192);
or U9617 (N_9617,In_2117,In_4514);
nand U9618 (N_9618,In_280,In_98);
and U9619 (N_9619,In_1113,In_4527);
xor U9620 (N_9620,In_856,In_1809);
and U9621 (N_9621,In_4246,In_964);
and U9622 (N_9622,In_4848,In_3217);
and U9623 (N_9623,In_4390,In_891);
or U9624 (N_9624,In_3245,In_91);
nand U9625 (N_9625,In_150,In_1828);
nand U9626 (N_9626,In_4832,In_4951);
and U9627 (N_9627,In_3970,In_1481);
nand U9628 (N_9628,In_3685,In_4924);
and U9629 (N_9629,In_3309,In_3066);
nor U9630 (N_9630,In_4992,In_4267);
or U9631 (N_9631,In_4586,In_3048);
xnor U9632 (N_9632,In_2169,In_4229);
xnor U9633 (N_9633,In_1580,In_1533);
nor U9634 (N_9634,In_1561,In_2660);
or U9635 (N_9635,In_4626,In_4592);
or U9636 (N_9636,In_2854,In_72);
xor U9637 (N_9637,In_2270,In_4657);
nand U9638 (N_9638,In_2295,In_1406);
nand U9639 (N_9639,In_722,In_4761);
or U9640 (N_9640,In_1864,In_3616);
or U9641 (N_9641,In_2420,In_3433);
or U9642 (N_9642,In_2275,In_4495);
nand U9643 (N_9643,In_1844,In_1110);
or U9644 (N_9644,In_2837,In_1819);
and U9645 (N_9645,In_912,In_1082);
nand U9646 (N_9646,In_1878,In_2666);
and U9647 (N_9647,In_3710,In_4560);
or U9648 (N_9648,In_2095,In_3436);
nand U9649 (N_9649,In_4260,In_1125);
nor U9650 (N_9650,In_2113,In_220);
xnor U9651 (N_9651,In_2432,In_2998);
nor U9652 (N_9652,In_1705,In_3915);
or U9653 (N_9653,In_2785,In_4630);
or U9654 (N_9654,In_958,In_6);
nand U9655 (N_9655,In_3447,In_4706);
nand U9656 (N_9656,In_4086,In_2846);
or U9657 (N_9657,In_587,In_3238);
nand U9658 (N_9658,In_3248,In_2339);
nor U9659 (N_9659,In_230,In_2873);
and U9660 (N_9660,In_3179,In_4149);
or U9661 (N_9661,In_518,In_4439);
or U9662 (N_9662,In_3289,In_1546);
and U9663 (N_9663,In_3875,In_1058);
and U9664 (N_9664,In_3731,In_2398);
xor U9665 (N_9665,In_1564,In_4385);
or U9666 (N_9666,In_2930,In_4423);
and U9667 (N_9667,In_1781,In_2393);
nor U9668 (N_9668,In_411,In_3735);
nand U9669 (N_9669,In_4378,In_39);
or U9670 (N_9670,In_3032,In_3584);
nand U9671 (N_9671,In_4841,In_84);
or U9672 (N_9672,In_4665,In_2354);
nor U9673 (N_9673,In_1919,In_3648);
and U9674 (N_9674,In_679,In_893);
and U9675 (N_9675,In_3048,In_4666);
and U9676 (N_9676,In_2307,In_2320);
nand U9677 (N_9677,In_725,In_3014);
and U9678 (N_9678,In_4087,In_4906);
nor U9679 (N_9679,In_3437,In_1212);
and U9680 (N_9680,In_3463,In_3822);
or U9681 (N_9681,In_2536,In_615);
or U9682 (N_9682,In_2139,In_2682);
and U9683 (N_9683,In_2417,In_2226);
nand U9684 (N_9684,In_425,In_1897);
or U9685 (N_9685,In_3540,In_1633);
nor U9686 (N_9686,In_4633,In_4024);
nand U9687 (N_9687,In_3926,In_4219);
nand U9688 (N_9688,In_951,In_4537);
nand U9689 (N_9689,In_4340,In_3354);
xor U9690 (N_9690,In_2257,In_4179);
nand U9691 (N_9691,In_319,In_1265);
or U9692 (N_9692,In_4365,In_4906);
and U9693 (N_9693,In_1895,In_1657);
or U9694 (N_9694,In_1346,In_1672);
nor U9695 (N_9695,In_1690,In_4948);
or U9696 (N_9696,In_865,In_1052);
and U9697 (N_9697,In_1451,In_3775);
nand U9698 (N_9698,In_1520,In_3003);
nand U9699 (N_9699,In_3004,In_354);
and U9700 (N_9700,In_259,In_4936);
nand U9701 (N_9701,In_4937,In_3838);
or U9702 (N_9702,In_398,In_4723);
or U9703 (N_9703,In_1327,In_4784);
and U9704 (N_9704,In_376,In_980);
nor U9705 (N_9705,In_1271,In_611);
and U9706 (N_9706,In_3317,In_112);
or U9707 (N_9707,In_3372,In_2358);
nand U9708 (N_9708,In_4848,In_3487);
nor U9709 (N_9709,In_4821,In_2418);
nor U9710 (N_9710,In_4842,In_4221);
and U9711 (N_9711,In_3979,In_3480);
nor U9712 (N_9712,In_3409,In_4778);
or U9713 (N_9713,In_3564,In_848);
or U9714 (N_9714,In_3732,In_2897);
nand U9715 (N_9715,In_1212,In_1720);
nand U9716 (N_9716,In_3678,In_1200);
or U9717 (N_9717,In_1192,In_4464);
and U9718 (N_9718,In_222,In_2615);
nor U9719 (N_9719,In_1746,In_4744);
or U9720 (N_9720,In_3772,In_2064);
and U9721 (N_9721,In_859,In_242);
and U9722 (N_9722,In_4153,In_1311);
or U9723 (N_9723,In_3578,In_4891);
nand U9724 (N_9724,In_4764,In_1571);
nor U9725 (N_9725,In_4542,In_2826);
nand U9726 (N_9726,In_1468,In_3651);
and U9727 (N_9727,In_4241,In_849);
xnor U9728 (N_9728,In_4443,In_1698);
nor U9729 (N_9729,In_1885,In_3995);
nand U9730 (N_9730,In_2949,In_602);
nor U9731 (N_9731,In_2934,In_2723);
or U9732 (N_9732,In_794,In_4811);
and U9733 (N_9733,In_204,In_3907);
nand U9734 (N_9734,In_1262,In_1842);
nor U9735 (N_9735,In_3690,In_2510);
or U9736 (N_9736,In_2312,In_1481);
nor U9737 (N_9737,In_3365,In_92);
xnor U9738 (N_9738,In_204,In_1745);
nor U9739 (N_9739,In_594,In_3800);
and U9740 (N_9740,In_4253,In_2903);
nor U9741 (N_9741,In_4912,In_4739);
and U9742 (N_9742,In_3857,In_3566);
nor U9743 (N_9743,In_3027,In_645);
or U9744 (N_9744,In_2275,In_1805);
xnor U9745 (N_9745,In_3439,In_1646);
nand U9746 (N_9746,In_3550,In_3826);
xnor U9747 (N_9747,In_1350,In_4550);
or U9748 (N_9748,In_292,In_1378);
nor U9749 (N_9749,In_3505,In_1878);
xnor U9750 (N_9750,In_3577,In_4788);
or U9751 (N_9751,In_4468,In_4437);
nor U9752 (N_9752,In_190,In_2375);
xor U9753 (N_9753,In_25,In_713);
or U9754 (N_9754,In_1256,In_3989);
xnor U9755 (N_9755,In_2828,In_906);
nand U9756 (N_9756,In_552,In_4387);
nand U9757 (N_9757,In_4299,In_1750);
or U9758 (N_9758,In_439,In_1453);
nor U9759 (N_9759,In_4175,In_3197);
nor U9760 (N_9760,In_2101,In_3995);
or U9761 (N_9761,In_3982,In_1060);
and U9762 (N_9762,In_2311,In_2545);
or U9763 (N_9763,In_1350,In_4752);
or U9764 (N_9764,In_4234,In_3572);
nand U9765 (N_9765,In_310,In_897);
and U9766 (N_9766,In_490,In_3479);
nor U9767 (N_9767,In_4979,In_3473);
or U9768 (N_9768,In_618,In_634);
nand U9769 (N_9769,In_421,In_4292);
nor U9770 (N_9770,In_2015,In_1969);
nand U9771 (N_9771,In_176,In_2154);
and U9772 (N_9772,In_785,In_4071);
xnor U9773 (N_9773,In_4425,In_2523);
or U9774 (N_9774,In_461,In_465);
nand U9775 (N_9775,In_3820,In_767);
nand U9776 (N_9776,In_1842,In_3109);
nor U9777 (N_9777,In_2905,In_3882);
and U9778 (N_9778,In_4831,In_2373);
or U9779 (N_9779,In_2812,In_591);
nand U9780 (N_9780,In_2354,In_569);
nor U9781 (N_9781,In_3416,In_4711);
nor U9782 (N_9782,In_990,In_655);
and U9783 (N_9783,In_3964,In_2494);
nor U9784 (N_9784,In_2678,In_4102);
nand U9785 (N_9785,In_3372,In_4496);
or U9786 (N_9786,In_1620,In_4846);
nand U9787 (N_9787,In_1910,In_1865);
nor U9788 (N_9788,In_2746,In_2083);
xor U9789 (N_9789,In_933,In_2972);
and U9790 (N_9790,In_2252,In_1108);
xnor U9791 (N_9791,In_1841,In_2681);
nand U9792 (N_9792,In_1385,In_2073);
nor U9793 (N_9793,In_820,In_2238);
nand U9794 (N_9794,In_2003,In_1908);
and U9795 (N_9795,In_4982,In_3386);
or U9796 (N_9796,In_4582,In_3187);
nand U9797 (N_9797,In_410,In_2375);
nand U9798 (N_9798,In_4603,In_3116);
and U9799 (N_9799,In_2457,In_1524);
or U9800 (N_9800,In_4700,In_3165);
and U9801 (N_9801,In_1070,In_4351);
and U9802 (N_9802,In_1667,In_2066);
nor U9803 (N_9803,In_3137,In_373);
nor U9804 (N_9804,In_1794,In_1325);
and U9805 (N_9805,In_993,In_2915);
nor U9806 (N_9806,In_2726,In_4250);
nand U9807 (N_9807,In_3549,In_2063);
and U9808 (N_9808,In_500,In_1641);
nor U9809 (N_9809,In_1284,In_4615);
nor U9810 (N_9810,In_101,In_4959);
or U9811 (N_9811,In_1779,In_2166);
nor U9812 (N_9812,In_1804,In_945);
nor U9813 (N_9813,In_2156,In_4914);
or U9814 (N_9814,In_1525,In_4569);
and U9815 (N_9815,In_2386,In_577);
or U9816 (N_9816,In_2085,In_4968);
nor U9817 (N_9817,In_4045,In_2549);
xor U9818 (N_9818,In_58,In_2722);
xor U9819 (N_9819,In_2358,In_2482);
xor U9820 (N_9820,In_474,In_351);
and U9821 (N_9821,In_1958,In_4800);
xor U9822 (N_9822,In_3182,In_881);
and U9823 (N_9823,In_2672,In_4757);
nor U9824 (N_9824,In_4845,In_575);
nand U9825 (N_9825,In_2051,In_3136);
nor U9826 (N_9826,In_4622,In_578);
nand U9827 (N_9827,In_3518,In_547);
nor U9828 (N_9828,In_3215,In_2378);
and U9829 (N_9829,In_673,In_2744);
xnor U9830 (N_9830,In_3065,In_1299);
nor U9831 (N_9831,In_3018,In_3101);
and U9832 (N_9832,In_2228,In_1983);
nand U9833 (N_9833,In_3358,In_4440);
or U9834 (N_9834,In_2096,In_1124);
or U9835 (N_9835,In_1361,In_3619);
nand U9836 (N_9836,In_4982,In_1000);
or U9837 (N_9837,In_4445,In_1845);
nand U9838 (N_9838,In_2711,In_1552);
and U9839 (N_9839,In_536,In_1431);
nor U9840 (N_9840,In_4878,In_3139);
or U9841 (N_9841,In_1296,In_2734);
xnor U9842 (N_9842,In_874,In_3399);
nor U9843 (N_9843,In_4017,In_1381);
and U9844 (N_9844,In_214,In_2913);
nor U9845 (N_9845,In_915,In_2452);
or U9846 (N_9846,In_2360,In_593);
and U9847 (N_9847,In_4519,In_3713);
nor U9848 (N_9848,In_1187,In_2150);
nor U9849 (N_9849,In_2764,In_3301);
nand U9850 (N_9850,In_300,In_3457);
and U9851 (N_9851,In_3271,In_2057);
nor U9852 (N_9852,In_443,In_2858);
nor U9853 (N_9853,In_3368,In_2880);
or U9854 (N_9854,In_2155,In_2777);
and U9855 (N_9855,In_1903,In_2585);
nor U9856 (N_9856,In_85,In_2074);
nor U9857 (N_9857,In_3826,In_3832);
and U9858 (N_9858,In_58,In_4004);
nand U9859 (N_9859,In_2481,In_785);
or U9860 (N_9860,In_418,In_2095);
or U9861 (N_9861,In_4549,In_3388);
and U9862 (N_9862,In_3670,In_1908);
xnor U9863 (N_9863,In_632,In_2618);
and U9864 (N_9864,In_877,In_3639);
or U9865 (N_9865,In_520,In_393);
and U9866 (N_9866,In_573,In_438);
nand U9867 (N_9867,In_2890,In_610);
and U9868 (N_9868,In_3436,In_2533);
nor U9869 (N_9869,In_4029,In_2077);
nor U9870 (N_9870,In_4392,In_636);
or U9871 (N_9871,In_554,In_1380);
nor U9872 (N_9872,In_4993,In_1742);
and U9873 (N_9873,In_3217,In_1759);
nand U9874 (N_9874,In_1598,In_2715);
and U9875 (N_9875,In_3219,In_286);
and U9876 (N_9876,In_1840,In_2004);
or U9877 (N_9877,In_3964,In_954);
and U9878 (N_9878,In_2932,In_1150);
or U9879 (N_9879,In_2841,In_267);
nand U9880 (N_9880,In_2808,In_215);
nor U9881 (N_9881,In_2523,In_604);
xnor U9882 (N_9882,In_3620,In_2032);
nand U9883 (N_9883,In_3816,In_3127);
nor U9884 (N_9884,In_1864,In_429);
nand U9885 (N_9885,In_3145,In_2629);
and U9886 (N_9886,In_2478,In_3687);
and U9887 (N_9887,In_1342,In_2506);
or U9888 (N_9888,In_2822,In_966);
or U9889 (N_9889,In_2872,In_2116);
nand U9890 (N_9890,In_1405,In_3705);
nand U9891 (N_9891,In_1787,In_940);
nand U9892 (N_9892,In_2429,In_415);
or U9893 (N_9893,In_2252,In_4669);
or U9894 (N_9894,In_742,In_2905);
and U9895 (N_9895,In_45,In_2923);
or U9896 (N_9896,In_475,In_3569);
nor U9897 (N_9897,In_2755,In_2055);
and U9898 (N_9898,In_2163,In_581);
or U9899 (N_9899,In_3470,In_171);
nand U9900 (N_9900,In_1667,In_3075);
xnor U9901 (N_9901,In_21,In_4754);
nand U9902 (N_9902,In_4276,In_2196);
nand U9903 (N_9903,In_3439,In_1736);
nor U9904 (N_9904,In_728,In_4461);
or U9905 (N_9905,In_845,In_4147);
nor U9906 (N_9906,In_3827,In_3145);
and U9907 (N_9907,In_4614,In_4529);
nand U9908 (N_9908,In_1395,In_247);
nor U9909 (N_9909,In_482,In_3430);
nor U9910 (N_9910,In_1849,In_666);
xnor U9911 (N_9911,In_3064,In_1520);
xor U9912 (N_9912,In_917,In_1882);
or U9913 (N_9913,In_2722,In_508);
nor U9914 (N_9914,In_3808,In_4817);
and U9915 (N_9915,In_647,In_4423);
or U9916 (N_9916,In_4634,In_441);
nor U9917 (N_9917,In_636,In_4926);
xnor U9918 (N_9918,In_4580,In_1373);
nand U9919 (N_9919,In_3410,In_4679);
nand U9920 (N_9920,In_1110,In_3303);
nand U9921 (N_9921,In_3013,In_3903);
xor U9922 (N_9922,In_2603,In_2024);
or U9923 (N_9923,In_1054,In_1138);
nor U9924 (N_9924,In_1677,In_4471);
xor U9925 (N_9925,In_1365,In_192);
or U9926 (N_9926,In_2025,In_1986);
nor U9927 (N_9927,In_1507,In_4563);
nor U9928 (N_9928,In_872,In_2967);
or U9929 (N_9929,In_3849,In_2727);
or U9930 (N_9930,In_3502,In_543);
or U9931 (N_9931,In_290,In_2691);
nand U9932 (N_9932,In_3539,In_2390);
nor U9933 (N_9933,In_3924,In_2994);
nand U9934 (N_9934,In_3821,In_3418);
nand U9935 (N_9935,In_2764,In_1360);
or U9936 (N_9936,In_1681,In_294);
nor U9937 (N_9937,In_3441,In_4391);
and U9938 (N_9938,In_941,In_2407);
and U9939 (N_9939,In_2407,In_2234);
nand U9940 (N_9940,In_2246,In_3121);
xnor U9941 (N_9941,In_971,In_2755);
nor U9942 (N_9942,In_1088,In_3424);
nand U9943 (N_9943,In_2161,In_256);
and U9944 (N_9944,In_681,In_3886);
nor U9945 (N_9945,In_2771,In_1153);
or U9946 (N_9946,In_2011,In_4610);
xor U9947 (N_9947,In_1272,In_4894);
or U9948 (N_9948,In_4070,In_4569);
nor U9949 (N_9949,In_4335,In_3965);
nand U9950 (N_9950,In_308,In_856);
or U9951 (N_9951,In_143,In_2505);
nand U9952 (N_9952,In_4496,In_4348);
nor U9953 (N_9953,In_4248,In_4599);
or U9954 (N_9954,In_776,In_273);
and U9955 (N_9955,In_1546,In_4747);
and U9956 (N_9956,In_3060,In_2219);
nand U9957 (N_9957,In_3168,In_250);
nor U9958 (N_9958,In_502,In_4957);
nor U9959 (N_9959,In_4905,In_945);
and U9960 (N_9960,In_1245,In_3248);
nand U9961 (N_9961,In_182,In_3000);
xnor U9962 (N_9962,In_236,In_1044);
nor U9963 (N_9963,In_2340,In_596);
or U9964 (N_9964,In_2809,In_4186);
nor U9965 (N_9965,In_715,In_1849);
nand U9966 (N_9966,In_1076,In_2196);
nand U9967 (N_9967,In_3279,In_373);
and U9968 (N_9968,In_1938,In_2359);
or U9969 (N_9969,In_3555,In_2727);
and U9970 (N_9970,In_557,In_259);
nor U9971 (N_9971,In_2452,In_3297);
nor U9972 (N_9972,In_1046,In_3190);
or U9973 (N_9973,In_92,In_3871);
xnor U9974 (N_9974,In_1766,In_2939);
nor U9975 (N_9975,In_4281,In_4863);
nand U9976 (N_9976,In_4017,In_1006);
nor U9977 (N_9977,In_1381,In_383);
or U9978 (N_9978,In_3938,In_3005);
nand U9979 (N_9979,In_2707,In_1768);
or U9980 (N_9980,In_2767,In_2142);
nand U9981 (N_9981,In_4535,In_4443);
xnor U9982 (N_9982,In_2532,In_3040);
nand U9983 (N_9983,In_1171,In_2274);
nand U9984 (N_9984,In_627,In_1401);
nand U9985 (N_9985,In_2249,In_2643);
nor U9986 (N_9986,In_1891,In_1928);
or U9987 (N_9987,In_1203,In_1246);
nand U9988 (N_9988,In_4724,In_3860);
or U9989 (N_9989,In_4285,In_1268);
nor U9990 (N_9990,In_524,In_545);
or U9991 (N_9991,In_3705,In_3994);
or U9992 (N_9992,In_4108,In_4032);
or U9993 (N_9993,In_3793,In_3971);
nor U9994 (N_9994,In_2796,In_4596);
and U9995 (N_9995,In_1070,In_4876);
nand U9996 (N_9996,In_3603,In_2713);
or U9997 (N_9997,In_696,In_3621);
nor U9998 (N_9998,In_387,In_1532);
nand U9999 (N_9999,In_249,In_1776);
or U10000 (N_10000,N_1864,N_4061);
nand U10001 (N_10001,N_3557,N_211);
nor U10002 (N_10002,N_4325,N_4955);
or U10003 (N_10003,N_2007,N_3150);
nor U10004 (N_10004,N_2672,N_7405);
nand U10005 (N_10005,N_7922,N_8509);
xor U10006 (N_10006,N_220,N_9681);
nor U10007 (N_10007,N_2079,N_7102);
and U10008 (N_10008,N_9075,N_6520);
xor U10009 (N_10009,N_2429,N_9602);
or U10010 (N_10010,N_573,N_8761);
or U10011 (N_10011,N_7403,N_5595);
nor U10012 (N_10012,N_1998,N_5217);
nor U10013 (N_10013,N_1621,N_7663);
nand U10014 (N_10014,N_9528,N_6595);
and U10015 (N_10015,N_8964,N_3298);
nand U10016 (N_10016,N_4039,N_3674);
nand U10017 (N_10017,N_6835,N_1775);
nand U10018 (N_10018,N_2633,N_7618);
nor U10019 (N_10019,N_6429,N_9105);
nand U10020 (N_10020,N_4978,N_927);
nand U10021 (N_10021,N_5293,N_4040);
xor U10022 (N_10022,N_9680,N_7038);
nor U10023 (N_10023,N_5508,N_4048);
nor U10024 (N_10024,N_1988,N_4683);
and U10025 (N_10025,N_8565,N_527);
or U10026 (N_10026,N_3481,N_5505);
and U10027 (N_10027,N_3086,N_7068);
nand U10028 (N_10028,N_3068,N_2221);
nor U10029 (N_10029,N_592,N_7932);
nand U10030 (N_10030,N_1206,N_8474);
nor U10031 (N_10031,N_2226,N_8040);
nor U10032 (N_10032,N_1924,N_9840);
nor U10033 (N_10033,N_2062,N_9863);
nand U10034 (N_10034,N_6091,N_2494);
or U10035 (N_10035,N_4499,N_5283);
and U10036 (N_10036,N_9821,N_6965);
or U10037 (N_10037,N_7937,N_6395);
nor U10038 (N_10038,N_2823,N_6304);
and U10039 (N_10039,N_4666,N_585);
nand U10040 (N_10040,N_3616,N_284);
nand U10041 (N_10041,N_4989,N_6352);
nand U10042 (N_10042,N_3853,N_6857);
and U10043 (N_10043,N_7796,N_5710);
xor U10044 (N_10044,N_4654,N_8163);
nand U10045 (N_10045,N_2511,N_5430);
nor U10046 (N_10046,N_3098,N_4923);
or U10047 (N_10047,N_9456,N_5821);
nor U10048 (N_10048,N_9768,N_5754);
nor U10049 (N_10049,N_730,N_7779);
and U10050 (N_10050,N_8347,N_778);
and U10051 (N_10051,N_3726,N_1535);
or U10052 (N_10052,N_8870,N_7020);
and U10053 (N_10053,N_8937,N_8805);
xor U10054 (N_10054,N_290,N_2994);
and U10055 (N_10055,N_3882,N_9799);
or U10056 (N_10056,N_1235,N_3408);
or U10057 (N_10057,N_9123,N_5998);
and U10058 (N_10058,N_551,N_6126);
nand U10059 (N_10059,N_2924,N_3862);
nor U10060 (N_10060,N_7889,N_6828);
or U10061 (N_10061,N_323,N_7564);
and U10062 (N_10062,N_6206,N_3015);
or U10063 (N_10063,N_5145,N_9995);
or U10064 (N_10064,N_727,N_63);
nor U10065 (N_10065,N_6462,N_6087);
nand U10066 (N_10066,N_7621,N_2840);
nand U10067 (N_10067,N_1728,N_2655);
nand U10068 (N_10068,N_2100,N_2235);
and U10069 (N_10069,N_4276,N_675);
nand U10070 (N_10070,N_1428,N_7416);
xor U10071 (N_10071,N_2454,N_8437);
and U10072 (N_10072,N_1909,N_2019);
nand U10073 (N_10073,N_1501,N_3736);
nor U10074 (N_10074,N_6711,N_4672);
and U10075 (N_10075,N_4475,N_2264);
and U10076 (N_10076,N_1510,N_4364);
or U10077 (N_10077,N_4434,N_7085);
nand U10078 (N_10078,N_1450,N_8592);
nor U10079 (N_10079,N_106,N_3076);
and U10080 (N_10080,N_6930,N_9145);
nand U10081 (N_10081,N_4793,N_6513);
or U10082 (N_10082,N_5352,N_6209);
or U10083 (N_10083,N_3701,N_6474);
or U10084 (N_10084,N_8914,N_2613);
nand U10085 (N_10085,N_5102,N_2066);
nor U10086 (N_10086,N_7311,N_7241);
or U10087 (N_10087,N_6690,N_2940);
nand U10088 (N_10088,N_3484,N_2905);
nor U10089 (N_10089,N_785,N_854);
and U10090 (N_10090,N_4304,N_5785);
nand U10091 (N_10091,N_6191,N_4412);
or U10092 (N_10092,N_6421,N_9174);
nand U10093 (N_10093,N_3125,N_8485);
nor U10094 (N_10094,N_756,N_2350);
or U10095 (N_10095,N_8164,N_9429);
and U10096 (N_10096,N_6005,N_7256);
nor U10097 (N_10097,N_2039,N_2992);
nand U10098 (N_10098,N_7099,N_6457);
nand U10099 (N_10099,N_5668,N_8323);
nand U10100 (N_10100,N_8907,N_1805);
nor U10101 (N_10101,N_2509,N_4707);
or U10102 (N_10102,N_9857,N_8793);
nand U10103 (N_10103,N_8380,N_4881);
nand U10104 (N_10104,N_5651,N_4222);
nor U10105 (N_10105,N_5959,N_5611);
nand U10106 (N_10106,N_2964,N_7856);
nor U10107 (N_10107,N_2484,N_8117);
and U10108 (N_10108,N_5432,N_5697);
nand U10109 (N_10109,N_2304,N_7673);
nand U10110 (N_10110,N_7142,N_2579);
nor U10111 (N_10111,N_1761,N_217);
nor U10112 (N_10112,N_9848,N_5187);
nand U10113 (N_10113,N_7630,N_8458);
nand U10114 (N_10114,N_3929,N_5439);
xor U10115 (N_10115,N_8528,N_5367);
and U10116 (N_10116,N_5490,N_8095);
and U10117 (N_10117,N_3091,N_51);
or U10118 (N_10118,N_8419,N_640);
and U10119 (N_10119,N_5847,N_7827);
nor U10120 (N_10120,N_8846,N_7198);
nand U10121 (N_10121,N_2929,N_2174);
or U10122 (N_10122,N_5342,N_4336);
nor U10123 (N_10123,N_2841,N_7975);
or U10124 (N_10124,N_3516,N_5245);
nor U10125 (N_10125,N_6406,N_6879);
nor U10126 (N_10126,N_4252,N_131);
and U10127 (N_10127,N_1973,N_5506);
nor U10128 (N_10128,N_6233,N_3887);
nor U10129 (N_10129,N_9153,N_8316);
xor U10130 (N_10130,N_1222,N_2391);
nor U10131 (N_10131,N_1242,N_3467);
or U10132 (N_10132,N_6533,N_7036);
and U10133 (N_10133,N_2734,N_7331);
nor U10134 (N_10134,N_6010,N_9779);
or U10135 (N_10135,N_5377,N_1368);
nor U10136 (N_10136,N_2786,N_5023);
and U10137 (N_10137,N_6459,N_6725);
or U10138 (N_10138,N_2289,N_6441);
nand U10139 (N_10139,N_1611,N_2510);
nor U10140 (N_10140,N_8886,N_6150);
and U10141 (N_10141,N_8058,N_8029);
xnor U10142 (N_10142,N_6167,N_9638);
nor U10143 (N_10143,N_6756,N_2206);
nand U10144 (N_10144,N_3375,N_9362);
nor U10145 (N_10145,N_6733,N_5330);
nor U10146 (N_10146,N_9233,N_7516);
nand U10147 (N_10147,N_1599,N_9138);
nor U10148 (N_10148,N_4709,N_9319);
and U10149 (N_10149,N_9802,N_5376);
and U10150 (N_10150,N_9500,N_1332);
nand U10151 (N_10151,N_4952,N_6743);
nand U10152 (N_10152,N_6407,N_219);
and U10153 (N_10153,N_6840,N_5464);
nor U10154 (N_10154,N_9028,N_7603);
nor U10155 (N_10155,N_7137,N_9795);
nand U10156 (N_10156,N_2738,N_8839);
nand U10157 (N_10157,N_4441,N_8531);
nand U10158 (N_10158,N_1796,N_5573);
or U10159 (N_10159,N_3707,N_4067);
nor U10160 (N_10160,N_1936,N_8219);
nor U10161 (N_10161,N_981,N_2588);
nor U10162 (N_10162,N_7177,N_8307);
nor U10163 (N_10163,N_1361,N_133);
and U10164 (N_10164,N_918,N_1978);
nand U10165 (N_10165,N_6214,N_3020);
nor U10166 (N_10166,N_9399,N_4278);
xor U10167 (N_10167,N_6850,N_5876);
nand U10168 (N_10168,N_9055,N_8411);
nand U10169 (N_10169,N_777,N_8660);
nand U10170 (N_10170,N_8157,N_1549);
or U10171 (N_10171,N_6548,N_4381);
and U10172 (N_10172,N_2227,N_5445);
xnor U10173 (N_10173,N_1119,N_8972);
or U10174 (N_10174,N_3040,N_8653);
nor U10175 (N_10175,N_8470,N_7696);
or U10176 (N_10176,N_729,N_8535);
xnor U10177 (N_10177,N_3850,N_7491);
nand U10178 (N_10178,N_6668,N_424);
or U10179 (N_10179,N_5219,N_2159);
nor U10180 (N_10180,N_9828,N_2694);
nand U10181 (N_10181,N_4894,N_7118);
nand U10182 (N_10182,N_4423,N_410);
nor U10183 (N_10183,N_5979,N_4349);
nor U10184 (N_10184,N_2351,N_4257);
nand U10185 (N_10185,N_3838,N_2461);
nor U10186 (N_10186,N_6859,N_3498);
nor U10187 (N_10187,N_4795,N_1769);
xor U10188 (N_10188,N_2747,N_3160);
or U10189 (N_10189,N_1228,N_3695);
xnor U10190 (N_10190,N_9482,N_2946);
and U10191 (N_10191,N_1388,N_6175);
xnor U10192 (N_10192,N_1096,N_8467);
and U10193 (N_10193,N_5924,N_5486);
and U10194 (N_10194,N_2233,N_2933);
nand U10195 (N_10195,N_3019,N_9214);
and U10196 (N_10196,N_6931,N_3818);
or U10197 (N_10197,N_2186,N_3947);
nand U10198 (N_10198,N_9958,N_2054);
and U10199 (N_10199,N_1462,N_3170);
nand U10200 (N_10200,N_7034,N_3956);
nand U10201 (N_10201,N_721,N_5570);
nand U10202 (N_10202,N_4600,N_4689);
nand U10203 (N_10203,N_1317,N_1932);
xor U10204 (N_10204,N_9240,N_8971);
and U10205 (N_10205,N_781,N_9310);
or U10206 (N_10206,N_5538,N_4047);
and U10207 (N_10207,N_293,N_1406);
nand U10208 (N_10208,N_6076,N_6526);
or U10209 (N_10209,N_4416,N_9235);
or U10210 (N_10210,N_5348,N_4258);
nor U10211 (N_10211,N_5662,N_3851);
or U10212 (N_10212,N_92,N_7968);
and U10213 (N_10213,N_4831,N_9659);
nor U10214 (N_10214,N_3789,N_3051);
nand U10215 (N_10215,N_226,N_628);
and U10216 (N_10216,N_1327,N_1068);
and U10217 (N_10217,N_3366,N_9307);
and U10218 (N_10218,N_8506,N_7866);
or U10219 (N_10219,N_9020,N_4291);
xnor U10220 (N_10220,N_8208,N_1420);
nand U10221 (N_10221,N_7386,N_4663);
or U10222 (N_10222,N_906,N_8717);
nand U10223 (N_10223,N_9062,N_4757);
nand U10224 (N_10224,N_4467,N_8065);
xnor U10225 (N_10225,N_5967,N_3566);
or U10226 (N_10226,N_2348,N_3801);
or U10227 (N_10227,N_5406,N_6278);
and U10228 (N_10228,N_2121,N_975);
and U10229 (N_10229,N_3510,N_1548);
nor U10230 (N_10230,N_9364,N_6146);
xor U10231 (N_10231,N_7329,N_2377);
and U10232 (N_10232,N_3356,N_2498);
xnor U10233 (N_10233,N_3799,N_9041);
nand U10234 (N_10234,N_8477,N_3286);
nor U10235 (N_10235,N_1118,N_6266);
and U10236 (N_10236,N_8744,N_3447);
or U10237 (N_10237,N_7053,N_5246);
or U10238 (N_10238,N_8178,N_1140);
or U10239 (N_10239,N_2139,N_6774);
and U10240 (N_10240,N_4588,N_2947);
and U10241 (N_10241,N_1070,N_4010);
xnor U10242 (N_10242,N_6242,N_701);
xor U10243 (N_10243,N_7307,N_2251);
nor U10244 (N_10244,N_1677,N_6168);
and U10245 (N_10245,N_4229,N_4386);
xnor U10246 (N_10246,N_1861,N_7362);
nor U10247 (N_10247,N_6614,N_2867);
nand U10248 (N_10248,N_9895,N_1733);
xnor U10249 (N_10249,N_222,N_142);
nand U10250 (N_10250,N_6306,N_6020);
and U10251 (N_10251,N_475,N_5032);
nor U10252 (N_10252,N_7836,N_3796);
or U10253 (N_10253,N_8772,N_4315);
and U10254 (N_10254,N_9612,N_5534);
nand U10255 (N_10255,N_2599,N_365);
nor U10256 (N_10256,N_8913,N_9172);
nor U10257 (N_10257,N_3392,N_4995);
nor U10258 (N_10258,N_2175,N_5333);
or U10259 (N_10259,N_4368,N_3834);
nand U10260 (N_10260,N_3774,N_6435);
nand U10261 (N_10261,N_1706,N_3045);
nand U10262 (N_10262,N_8328,N_5412);
xnor U10263 (N_10263,N_3655,N_2667);
nand U10264 (N_10264,N_4908,N_8071);
or U10265 (N_10265,N_2312,N_9609);
and U10266 (N_10266,N_2874,N_3275);
or U10267 (N_10267,N_3176,N_5122);
nor U10268 (N_10268,N_9427,N_2600);
or U10269 (N_10269,N_3438,N_9639);
xnor U10270 (N_10270,N_8083,N_3415);
nor U10271 (N_10271,N_5263,N_1987);
nor U10272 (N_10272,N_180,N_4904);
nand U10273 (N_10273,N_9941,N_1562);
and U10274 (N_10274,N_8089,N_8657);
nor U10275 (N_10275,N_1930,N_2369);
nor U10276 (N_10276,N_8946,N_5203);
or U10277 (N_10277,N_5626,N_9739);
and U10278 (N_10278,N_5907,N_2883);
nand U10279 (N_10279,N_4376,N_6463);
nand U10280 (N_10280,N_5489,N_9730);
nand U10281 (N_10281,N_2154,N_6186);
and U10282 (N_10282,N_3752,N_7125);
or U10283 (N_10283,N_2355,N_689);
or U10284 (N_10284,N_8500,N_3431);
nor U10285 (N_10285,N_2288,N_3270);
and U10286 (N_10286,N_2758,N_5653);
nand U10287 (N_10287,N_7052,N_5807);
nor U10288 (N_10288,N_1486,N_6361);
and U10289 (N_10289,N_7724,N_977);
nand U10290 (N_10290,N_4074,N_5119);
or U10291 (N_10291,N_8568,N_6517);
nor U10292 (N_10292,N_7272,N_7711);
or U10293 (N_10293,N_3363,N_3478);
xor U10294 (N_10294,N_4549,N_3300);
and U10295 (N_10295,N_3224,N_563);
and U10296 (N_10296,N_2257,N_4629);
nand U10297 (N_10297,N_4266,N_4275);
nor U10298 (N_10298,N_2056,N_4158);
or U10299 (N_10299,N_3221,N_4993);
and U10300 (N_10300,N_4311,N_1597);
and U10301 (N_10301,N_1750,N_7749);
or U10302 (N_10302,N_4591,N_9564);
xor U10303 (N_10303,N_7801,N_8879);
nand U10304 (N_10304,N_4250,N_5005);
and U10305 (N_10305,N_6716,N_1715);
or U10306 (N_10306,N_909,N_8200);
nor U10307 (N_10307,N_9261,N_7222);
xor U10308 (N_10308,N_8041,N_6764);
or U10309 (N_10309,N_202,N_8986);
nor U10310 (N_10310,N_4122,N_4938);
or U10311 (N_10311,N_5992,N_3546);
xnor U10312 (N_10312,N_5658,N_5084);
nand U10313 (N_10313,N_2036,N_7953);
nor U10314 (N_10314,N_1095,N_5628);
nand U10315 (N_10315,N_768,N_4263);
or U10316 (N_10316,N_3021,N_4976);
and U10317 (N_10317,N_7905,N_4410);
nand U10318 (N_10318,N_1204,N_3564);
or U10319 (N_10319,N_4283,N_4969);
nand U10320 (N_10320,N_8424,N_9098);
and U10321 (N_10321,N_1665,N_8862);
and U10322 (N_10322,N_6867,N_8202);
or U10323 (N_10323,N_513,N_8782);
or U10324 (N_10324,N_7651,N_8514);
nor U10325 (N_10325,N_9245,N_898);
nand U10326 (N_10326,N_9589,N_3713);
and U10327 (N_10327,N_2853,N_490);
or U10328 (N_10328,N_3833,N_1069);
nor U10329 (N_10329,N_6874,N_7352);
and U10330 (N_10330,N_6094,N_8698);
xor U10331 (N_10331,N_5047,N_9443);
nor U10332 (N_10332,N_6993,N_8350);
nand U10333 (N_10333,N_6040,N_3211);
or U10334 (N_10334,N_8300,N_4430);
nand U10335 (N_10335,N_3374,N_9994);
nand U10336 (N_10336,N_8126,N_39);
nand U10337 (N_10337,N_8712,N_9263);
or U10338 (N_10338,N_8413,N_8962);
and U10339 (N_10339,N_741,N_7738);
nor U10340 (N_10340,N_9853,N_1057);
and U10341 (N_10341,N_8222,N_808);
xor U10342 (N_10342,N_8230,N_8161);
xnor U10343 (N_10343,N_4713,N_6964);
nand U10344 (N_10344,N_4457,N_7167);
nand U10345 (N_10345,N_7989,N_4830);
nor U10346 (N_10346,N_1638,N_5606);
nand U10347 (N_10347,N_2106,N_5780);
or U10348 (N_10348,N_2172,N_1359);
nand U10349 (N_10349,N_8808,N_8194);
and U10350 (N_10350,N_4882,N_9552);
nand U10351 (N_10351,N_6316,N_2602);
nor U10352 (N_10352,N_2373,N_6638);
nor U10353 (N_10353,N_5418,N_739);
xnor U10354 (N_10354,N_7141,N_3372);
nand U10355 (N_10355,N_8724,N_1410);
nor U10356 (N_10356,N_4554,N_4699);
nand U10357 (N_10357,N_912,N_9773);
nand U10358 (N_10358,N_2088,N_8261);
nor U10359 (N_10359,N_7424,N_5116);
nand U10360 (N_10360,N_172,N_6344);
nor U10361 (N_10361,N_5537,N_9143);
nor U10362 (N_10362,N_7410,N_382);
and U10363 (N_10363,N_9081,N_6499);
and U10364 (N_10364,N_3642,N_1871);
or U10365 (N_10365,N_5727,N_3760);
or U10366 (N_10366,N_7443,N_1591);
and U10367 (N_10367,N_8461,N_578);
xnor U10368 (N_10368,N_7124,N_2732);
and U10369 (N_10369,N_597,N_1732);
or U10370 (N_10370,N_8439,N_5331);
nor U10371 (N_10371,N_7452,N_3639);
nand U10372 (N_10372,N_2024,N_3964);
nor U10373 (N_10373,N_3756,N_3696);
and U10374 (N_10374,N_8850,N_6476);
and U10375 (N_10375,N_6443,N_8688);
nor U10376 (N_10376,N_154,N_6641);
nor U10377 (N_10377,N_7148,N_8158);
nand U10378 (N_10378,N_197,N_5533);
and U10379 (N_10379,N_6080,N_2870);
nand U10380 (N_10380,N_548,N_7004);
xnor U10381 (N_10381,N_2899,N_224);
nand U10382 (N_10382,N_3603,N_901);
and U10383 (N_10383,N_1485,N_1033);
nand U10384 (N_10384,N_890,N_7128);
nand U10385 (N_10385,N_5080,N_9400);
nor U10386 (N_10386,N_614,N_6885);
nand U10387 (N_10387,N_4806,N_5918);
or U10388 (N_10388,N_4178,N_926);
nor U10389 (N_10389,N_3663,N_6360);
xor U10390 (N_10390,N_9865,N_2959);
nand U10391 (N_10391,N_7981,N_2656);
nor U10392 (N_10392,N_8129,N_249);
nand U10393 (N_10393,N_6095,N_564);
and U10394 (N_10394,N_4975,N_2966);
nor U10395 (N_10395,N_4023,N_8109);
nand U10396 (N_10396,N_4119,N_6410);
xor U10397 (N_10397,N_3120,N_7652);
nor U10398 (N_10398,N_7186,N_1633);
xnor U10399 (N_10399,N_8220,N_1085);
nor U10400 (N_10400,N_1121,N_5101);
nor U10401 (N_10401,N_5070,N_5273);
or U10402 (N_10402,N_4347,N_4747);
or U10403 (N_10403,N_6502,N_8948);
nor U10404 (N_10404,N_4928,N_4021);
nor U10405 (N_10405,N_6500,N_7464);
or U10406 (N_10406,N_5878,N_8750);
nand U10407 (N_10407,N_6710,N_7617);
and U10408 (N_10408,N_2128,N_5737);
nor U10409 (N_10409,N_6114,N_878);
nand U10410 (N_10410,N_3317,N_9499);
xor U10411 (N_10411,N_4450,N_3138);
nand U10412 (N_10412,N_8557,N_1514);
xnor U10413 (N_10413,N_2240,N_9571);
or U10414 (N_10414,N_6032,N_3400);
or U10415 (N_10415,N_1594,N_3458);
nand U10416 (N_10416,N_9112,N_8049);
nor U10417 (N_10417,N_3991,N_6207);
and U10418 (N_10418,N_5511,N_8436);
nor U10419 (N_10419,N_2217,N_1505);
and U10420 (N_10420,N_4986,N_4334);
nand U10421 (N_10421,N_5623,N_8050);
and U10422 (N_10422,N_5451,N_7132);
or U10423 (N_10423,N_1040,N_3876);
nor U10424 (N_10424,N_9069,N_1739);
nor U10425 (N_10425,N_4319,N_4162);
xor U10426 (N_10426,N_5207,N_2135);
nand U10427 (N_10427,N_539,N_3675);
xor U10428 (N_10428,N_8920,N_5151);
and U10429 (N_10429,N_9371,N_3858);
nand U10430 (N_10430,N_9824,N_5220);
or U10431 (N_10431,N_3683,N_1602);
xor U10432 (N_10432,N_6848,N_1282);
nor U10433 (N_10433,N_7037,N_2204);
and U10434 (N_10434,N_1376,N_9598);
nor U10435 (N_10435,N_7248,N_9226);
or U10436 (N_10436,N_2029,N_5747);
nand U10437 (N_10437,N_2469,N_3217);
nor U10438 (N_10438,N_2497,N_7457);
and U10439 (N_10439,N_4157,N_268);
and U10440 (N_10440,N_838,N_3029);
and U10441 (N_10441,N_6324,N_3377);
and U10442 (N_10442,N_4286,N_449);
or U10443 (N_10443,N_1903,N_9619);
nor U10444 (N_10444,N_1295,N_5684);
or U10445 (N_10445,N_704,N_103);
xor U10446 (N_10446,N_521,N_123);
nor U10447 (N_10447,N_5456,N_9260);
nand U10448 (N_10448,N_5788,N_457);
nand U10449 (N_10449,N_8926,N_4584);
and U10450 (N_10450,N_2714,N_4687);
or U10451 (N_10451,N_7016,N_7829);
and U10452 (N_10452,N_8517,N_6388);
nor U10453 (N_10453,N_793,N_1371);
or U10454 (N_10454,N_3247,N_2665);
nand U10455 (N_10455,N_2418,N_9666);
or U10456 (N_10456,N_3805,N_7494);
or U10457 (N_10457,N_1567,N_1011);
nor U10458 (N_10458,N_1253,N_4863);
nand U10459 (N_10459,N_9288,N_398);
xor U10460 (N_10460,N_2532,N_7730);
and U10461 (N_10461,N_7861,N_427);
and U10462 (N_10462,N_1669,N_4848);
nor U10463 (N_10463,N_3283,N_1720);
nor U10464 (N_10464,N_6546,N_9373);
nand U10465 (N_10465,N_9911,N_4660);
or U10466 (N_10466,N_1647,N_8365);
or U10467 (N_10467,N_2094,N_2863);
xor U10468 (N_10468,N_9032,N_8824);
and U10469 (N_10469,N_2210,N_3548);
nand U10470 (N_10470,N_1673,N_772);
xnor U10471 (N_10471,N_1067,N_7288);
and U10472 (N_10472,N_3089,N_943);
or U10473 (N_10473,N_7558,N_1251);
nor U10474 (N_10474,N_9338,N_8973);
or U10475 (N_10475,N_7276,N_8234);
nand U10476 (N_10476,N_7971,N_3233);
and U10477 (N_10477,N_1280,N_8735);
or U10478 (N_10478,N_6059,N_6704);
nor U10479 (N_10479,N_4179,N_1565);
or U10480 (N_10480,N_8369,N_2344);
and U10481 (N_10481,N_4072,N_7458);
nor U10482 (N_10482,N_3759,N_3689);
nor U10483 (N_10483,N_4332,N_437);
nand U10484 (N_10484,N_4890,N_8575);
nor U10485 (N_10485,N_7316,N_4384);
or U10486 (N_10486,N_6724,N_2698);
xor U10487 (N_10487,N_4740,N_2857);
and U10488 (N_10488,N_1048,N_4697);
or U10489 (N_10489,N_798,N_1897);
and U10490 (N_10490,N_56,N_4615);
xnor U10491 (N_10491,N_7964,N_9108);
nor U10492 (N_10492,N_3631,N_4069);
nor U10493 (N_10493,N_742,N_7297);
nor U10494 (N_10494,N_5209,N_9925);
and U10495 (N_10495,N_6853,N_9737);
or U10496 (N_10496,N_2646,N_5676);
nor U10497 (N_10497,N_1303,N_3096);
and U10498 (N_10498,N_581,N_9933);
or U10499 (N_10499,N_4572,N_2382);
or U10500 (N_10500,N_6414,N_1062);
or U10501 (N_10501,N_413,N_5086);
or U10502 (N_10502,N_8822,N_8449);
or U10503 (N_10503,N_3575,N_1823);
nor U10504 (N_10504,N_40,N_1702);
nor U10505 (N_10505,N_8943,N_1224);
nand U10506 (N_10506,N_2360,N_6776);
or U10507 (N_10507,N_2424,N_8645);
nand U10508 (N_10508,N_8902,N_6107);
xor U10509 (N_10509,N_4324,N_1425);
or U10510 (N_10510,N_1137,N_4136);
nor U10511 (N_10511,N_112,N_402);
nand U10512 (N_10512,N_6612,N_227);
xor U10513 (N_10513,N_6149,N_9056);
nor U10514 (N_10514,N_6054,N_5458);
or U10515 (N_10515,N_3900,N_2459);
nor U10516 (N_10516,N_5756,N_9517);
or U10517 (N_10517,N_9337,N_1946);
nor U10518 (N_10518,N_7298,N_6078);
and U10519 (N_10519,N_1185,N_8582);
and U10520 (N_10520,N_7456,N_5251);
nor U10521 (N_10521,N_5558,N_455);
and U10522 (N_10522,N_8327,N_6022);
nor U10523 (N_10523,N_6026,N_7449);
nor U10524 (N_10524,N_7355,N_7781);
or U10525 (N_10525,N_2290,N_8001);
nand U10526 (N_10526,N_4695,N_8229);
xnor U10527 (N_10527,N_8415,N_6392);
and U10528 (N_10528,N_8919,N_5774);
nand U10529 (N_10529,N_1618,N_2089);
and U10530 (N_10530,N_231,N_8105);
or U10531 (N_10531,N_9635,N_5819);
nand U10532 (N_10532,N_4285,N_5477);
nor U10533 (N_10533,N_4026,N_1446);
nand U10534 (N_10534,N_8099,N_8726);
or U10535 (N_10535,N_7755,N_5279);
nor U10536 (N_10536,N_1949,N_2409);
and U10537 (N_10537,N_6093,N_7302);
nor U10538 (N_10538,N_212,N_5284);
nor U10539 (N_10539,N_4561,N_8799);
nand U10540 (N_10540,N_359,N_3079);
or U10541 (N_10541,N_7235,N_8252);
or U10542 (N_10542,N_6315,N_4132);
nor U10543 (N_10543,N_8664,N_4842);
nand U10544 (N_10544,N_9721,N_2025);
nor U10545 (N_10545,N_1955,N_4634);
and U10546 (N_10546,N_2146,N_5372);
nand U10547 (N_10547,N_2456,N_1168);
nand U10548 (N_10548,N_2142,N_7442);
nand U10549 (N_10549,N_2075,N_662);
xnor U10550 (N_10550,N_2620,N_7303);
nor U10551 (N_10551,N_3733,N_6112);
or U10552 (N_10552,N_2445,N_1850);
or U10553 (N_10553,N_1487,N_5859);
nand U10554 (N_10554,N_5519,N_1499);
and U10555 (N_10555,N_2414,N_579);
and U10556 (N_10556,N_478,N_2679);
and U10557 (N_10557,N_4333,N_7013);
nor U10558 (N_10558,N_3556,N_4407);
nor U10559 (N_10559,N_8954,N_532);
xnor U10560 (N_10560,N_7268,N_1001);
nor U10561 (N_10561,N_4148,N_1176);
nor U10562 (N_10562,N_6851,N_5641);
nor U10563 (N_10563,N_5928,N_5385);
nand U10564 (N_10564,N_9496,N_4300);
and U10565 (N_10565,N_6855,N_4828);
nor U10566 (N_10566,N_5180,N_2622);
nand U10567 (N_10567,N_5848,N_9054);
or U10568 (N_10568,N_9408,N_7219);
xnor U10569 (N_10569,N_3457,N_627);
or U10570 (N_10570,N_6789,N_3416);
or U10571 (N_10571,N_8275,N_3816);
nand U10572 (N_10572,N_5223,N_10);
nor U10573 (N_10573,N_8221,N_2157);
and U10574 (N_10574,N_6652,N_5725);
and U10575 (N_10575,N_8996,N_5485);
nand U10576 (N_10576,N_1679,N_9284);
nand U10577 (N_10577,N_2298,N_104);
and U10578 (N_10578,N_9280,N_6);
and U10579 (N_10579,N_8418,N_6148);
or U10580 (N_10580,N_3378,N_905);
and U10581 (N_10581,N_2650,N_7419);
and U10582 (N_10582,N_6356,N_7096);
and U10583 (N_10583,N_4338,N_8279);
nor U10584 (N_10584,N_5340,N_6050);
and U10585 (N_10585,N_5699,N_2155);
nand U10586 (N_10586,N_23,N_74);
and U10587 (N_10587,N_2671,N_4515);
nor U10588 (N_10588,N_5488,N_4429);
and U10589 (N_10589,N_3196,N_5995);
xnor U10590 (N_10590,N_294,N_7660);
nand U10591 (N_10591,N_3972,N_9565);
or U10592 (N_10592,N_1701,N_6385);
or U10593 (N_10593,N_8240,N_2560);
nand U10594 (N_10594,N_238,N_5875);
nor U10595 (N_10595,N_630,N_395);
nand U10596 (N_10596,N_7845,N_6173);
and U10597 (N_10597,N_2542,N_1925);
or U10598 (N_10598,N_260,N_683);
or U10599 (N_10599,N_2518,N_5896);
nor U10600 (N_10600,N_9436,N_7940);
nand U10601 (N_10601,N_1540,N_3108);
nor U10602 (N_10602,N_3017,N_7933);
and U10603 (N_10603,N_7474,N_8810);
nor U10604 (N_10604,N_3856,N_3920);
nor U10605 (N_10605,N_3931,N_4223);
nor U10606 (N_10606,N_8465,N_1666);
nor U10607 (N_10607,N_5973,N_6484);
nand U10608 (N_10608,N_6454,N_4502);
and U10609 (N_10609,N_266,N_7205);
and U10610 (N_10610,N_9606,N_8878);
nand U10611 (N_10611,N_6210,N_8423);
nand U10612 (N_10612,N_8137,N_9175);
or U10613 (N_10613,N_9996,N_2504);
or U10614 (N_10614,N_7566,N_2681);
or U10615 (N_10615,N_6524,N_2624);
and U10616 (N_10616,N_6493,N_8315);
nor U10617 (N_10617,N_5500,N_8250);
and U10618 (N_10618,N_7338,N_6376);
or U10619 (N_10619,N_372,N_3382);
or U10620 (N_10620,N_9579,N_3992);
xnor U10621 (N_10621,N_5769,N_218);
nor U10622 (N_10622,N_691,N_5336);
or U10623 (N_10623,N_3102,N_6829);
nor U10624 (N_10624,N_8039,N_6051);
nor U10625 (N_10625,N_8897,N_6019);
nand U10626 (N_10626,N_4034,N_1742);
or U10627 (N_10627,N_5686,N_1792);
nand U10628 (N_10628,N_9404,N_3832);
nor U10629 (N_10629,N_3734,N_2628);
xor U10630 (N_10630,N_6129,N_3323);
xor U10631 (N_10631,N_3396,N_1972);
nor U10632 (N_10632,N_3188,N_888);
nor U10633 (N_10633,N_8237,N_3448);
nand U10634 (N_10634,N_9184,N_4284);
and U10635 (N_10635,N_1258,N_4789);
xnor U10636 (N_10636,N_1890,N_612);
nor U10637 (N_10637,N_6773,N_765);
or U10638 (N_10638,N_273,N_2366);
and U10639 (N_10639,N_2854,N_7250);
nand U10640 (N_10640,N_5585,N_8668);
nand U10641 (N_10641,N_2611,N_6115);
or U10642 (N_10642,N_3231,N_7106);
xnor U10643 (N_10643,N_481,N_9734);
or U10644 (N_10644,N_6813,N_5692);
and U10645 (N_10645,N_3249,N_8044);
or U10646 (N_10646,N_7155,N_5711);
or U10647 (N_10647,N_7522,N_1804);
nand U10648 (N_10648,N_5343,N_5132);
nand U10649 (N_10649,N_3973,N_2191);
nor U10650 (N_10650,N_2197,N_1010);
nor U10651 (N_10651,N_9438,N_5578);
or U10652 (N_10652,N_7616,N_9544);
or U10653 (N_10653,N_47,N_1417);
nor U10654 (N_10654,N_451,N_7091);
or U10655 (N_10655,N_2358,N_4811);
nor U10656 (N_10656,N_7469,N_4988);
and U10657 (N_10657,N_9113,N_6506);
and U10658 (N_10658,N_5624,N_762);
nand U10659 (N_10659,N_2741,N_2192);
xnor U10660 (N_10660,N_7418,N_1697);
and U10661 (N_10661,N_5698,N_7070);
nor U10662 (N_10662,N_7342,N_5137);
nor U10663 (N_10663,N_6760,N_8613);
nor U10664 (N_10664,N_1883,N_5262);
and U10665 (N_10665,N_687,N_6491);
or U10666 (N_10666,N_4130,N_4611);
nor U10667 (N_10667,N_2769,N_9208);
or U10668 (N_10668,N_4290,N_7340);
or U10669 (N_10669,N_6968,N_8409);
nand U10670 (N_10670,N_835,N_9128);
xor U10671 (N_10671,N_9199,N_8454);
xor U10672 (N_10672,N_6063,N_6714);
and U10673 (N_10673,N_8579,N_7804);
and U10674 (N_10674,N_8608,N_2984);
or U10675 (N_10675,N_3933,N_9881);
nor U10676 (N_10676,N_4785,N_6923);
xnor U10677 (N_10677,N_7642,N_7299);
xor U10678 (N_10678,N_7479,N_5017);
and U10679 (N_10679,N_6925,N_176);
or U10680 (N_10680,N_1477,N_3026);
and U10681 (N_10681,N_328,N_9396);
and U10682 (N_10682,N_4809,N_6831);
and U10683 (N_10683,N_1414,N_7899);
or U10684 (N_10684,N_9167,N_7502);
nand U10685 (N_10685,N_7669,N_6057);
nand U10686 (N_10686,N_6470,N_7394);
nor U10687 (N_10687,N_9883,N_9039);
or U10688 (N_10688,N_5645,N_9715);
nor U10689 (N_10689,N_5362,N_2040);
or U10690 (N_10690,N_6064,N_1034);
and U10691 (N_10691,N_6975,N_8056);
nand U10692 (N_10692,N_3879,N_2353);
nand U10693 (N_10693,N_5947,N_3343);
and U10694 (N_10694,N_1421,N_1056);
nand U10695 (N_10695,N_2879,N_9074);
and U10696 (N_10696,N_2031,N_8671);
or U10697 (N_10697,N_6619,N_2876);
nand U10698 (N_10698,N_7705,N_4182);
nand U10699 (N_10699,N_7440,N_8706);
or U10700 (N_10700,N_3335,N_8923);
and U10701 (N_10701,N_4929,N_5083);
or U10702 (N_10702,N_2880,N_9000);
and U10703 (N_10703,N_2829,N_5073);
xnor U10704 (N_10704,N_7935,N_7117);
or U10705 (N_10705,N_5112,N_6265);
nand U10706 (N_10706,N_9931,N_4339);
nand U10707 (N_10707,N_5289,N_3877);
or U10708 (N_10708,N_8272,N_3280);
nand U10709 (N_10709,N_3672,N_1210);
and U10710 (N_10710,N_8938,N_2093);
nand U10711 (N_10711,N_6213,N_8806);
or U10712 (N_10712,N_8478,N_2711);
nand U10713 (N_10713,N_7619,N_2387);
nor U10714 (N_10714,N_7415,N_6037);
and U10715 (N_10715,N_8741,N_7743);
nand U10716 (N_10716,N_1777,N_3646);
and U10717 (N_10717,N_1498,N_1325);
nor U10718 (N_10718,N_3487,N_4471);
and U10719 (N_10719,N_8597,N_1993);
nor U10720 (N_10720,N_2915,N_6246);
or U10721 (N_10721,N_7314,N_1213);
and U10722 (N_10722,N_8792,N_9851);
and U10723 (N_10723,N_9586,N_165);
or U10724 (N_10724,N_3907,N_375);
nor U10725 (N_10725,N_8652,N_7086);
nand U10726 (N_10726,N_8410,N_1866);
and U10727 (N_10727,N_4980,N_5571);
or U10728 (N_10728,N_1826,N_6738);
nor U10729 (N_10729,N_1401,N_2950);
nor U10730 (N_10730,N_9807,N_8103);
nand U10731 (N_10731,N_6818,N_4055);
nand U10732 (N_10732,N_6646,N_3077);
and U10733 (N_10733,N_80,N_7757);
or U10734 (N_10734,N_556,N_1339);
or U10735 (N_10735,N_5746,N_1482);
xor U10736 (N_10736,N_1541,N_7654);
or U10737 (N_10737,N_2496,N_5905);
and U10738 (N_10738,N_5517,N_5433);
xnor U10739 (N_10739,N_3295,N_1392);
and U10740 (N_10740,N_8860,N_9176);
nand U10741 (N_10741,N_6066,N_9223);
or U10742 (N_10742,N_2678,N_8807);
xor U10743 (N_10743,N_4551,N_3513);
or U10744 (N_10744,N_5481,N_8329);
and U10745 (N_10745,N_7728,N_6323);
and U10746 (N_10746,N_3797,N_2400);
nor U10747 (N_10747,N_1617,N_1324);
xor U10748 (N_10748,N_8654,N_3656);
nand U10749 (N_10749,N_2285,N_9888);
and U10750 (N_10750,N_9467,N_6481);
nand U10751 (N_10751,N_6926,N_9358);
or U10752 (N_10752,N_9109,N_2952);
nand U10753 (N_10753,N_7625,N_9470);
or U10754 (N_10754,N_1267,N_5357);
nor U10755 (N_10755,N_468,N_1971);
nand U10756 (N_10756,N_9256,N_7546);
or U10757 (N_10757,N_1246,N_3267);
and U10758 (N_10758,N_2383,N_1538);
xor U10759 (N_10759,N_7389,N_9027);
or U10760 (N_10760,N_7523,N_942);
and U10761 (N_10761,N_9965,N_2858);
xor U10762 (N_10762,N_971,N_2453);
and U10763 (N_10763,N_6294,N_5665);
and U10764 (N_10764,N_6179,N_9006);
nand U10765 (N_10765,N_2169,N_4254);
nand U10766 (N_10766,N_6348,N_4954);
nand U10767 (N_10767,N_620,N_2828);
or U10768 (N_10768,N_6883,N_5194);
nand U10769 (N_10769,N_9516,N_7461);
nand U10770 (N_10770,N_8317,N_9596);
or U10771 (N_10771,N_3745,N_2277);
and U10772 (N_10772,N_6287,N_9146);
xor U10773 (N_10773,N_8764,N_4650);
and U10774 (N_10774,N_1716,N_2814);
nand U10775 (N_10775,N_2606,N_4873);
nand U10776 (N_10776,N_1227,N_8881);
nor U10777 (N_10777,N_9423,N_6586);
and U10778 (N_10778,N_5022,N_5654);
nand U10779 (N_10779,N_9908,N_2381);
nand U10780 (N_10780,N_4534,N_1380);
nand U10781 (N_10781,N_9543,N_3025);
xnor U10782 (N_10782,N_9121,N_2941);
nor U10783 (N_10783,N_964,N_6569);
nand U10784 (N_10784,N_241,N_5404);
and U10785 (N_10785,N_5643,N_4739);
nor U10786 (N_10786,N_1608,N_5764);
nand U10787 (N_10787,N_3321,N_9633);
nand U10788 (N_10788,N_1887,N_8885);
or U10789 (N_10789,N_6942,N_1526);
nor U10790 (N_10790,N_3167,N_7098);
and U10791 (N_10791,N_5447,N_1846);
nand U10792 (N_10792,N_7735,N_4060);
nand U10793 (N_10793,N_5031,N_7707);
and U10794 (N_10794,N_317,N_3845);
or U10795 (N_10795,N_1680,N_6881);
xnor U10796 (N_10796,N_3899,N_2713);
nor U10797 (N_10797,N_2975,N_8730);
or U10798 (N_10798,N_7466,N_903);
or U10799 (N_10799,N_760,N_7994);
or U10800 (N_10800,N_8112,N_8615);
or U10801 (N_10801,N_4271,N_7472);
nand U10802 (N_10802,N_9024,N_6559);
nand U10803 (N_10803,N_3934,N_507);
and U10804 (N_10804,N_5354,N_526);
nor U10805 (N_10805,N_3894,N_5494);
and U10806 (N_10806,N_8958,N_815);
and U10807 (N_10807,N_9416,N_9707);
nand U10808 (N_10808,N_9561,N_1179);
nor U10809 (N_10809,N_9577,N_3331);
nand U10810 (N_10810,N_8023,N_7151);
or U10811 (N_10811,N_1226,N_1928);
xor U10812 (N_10812,N_7844,N_7513);
and U10813 (N_10813,N_915,N_3380);
and U10814 (N_10814,N_8268,N_6661);
xnor U10815 (N_10815,N_6343,N_5523);
nor U10816 (N_10816,N_9262,N_1374);
or U10817 (N_10817,N_1120,N_645);
xnor U10818 (N_10818,N_6911,N_682);
nor U10819 (N_10819,N_8511,N_8346);
or U10820 (N_10820,N_5379,N_3953);
and U10821 (N_10821,N_7279,N_5422);
nand U10822 (N_10822,N_2203,N_3579);
nor U10823 (N_10823,N_4891,N_3868);
nand U10824 (N_10824,N_4896,N_799);
nand U10825 (N_10825,N_665,N_8856);
and U10826 (N_10826,N_5256,N_2402);
xnor U10827 (N_10827,N_1997,N_4218);
nand U10828 (N_10828,N_8728,N_5827);
nand U10829 (N_10829,N_162,N_4418);
and U10830 (N_10830,N_1014,N_8495);
nand U10831 (N_10831,N_71,N_907);
nand U10832 (N_10832,N_9660,N_1212);
or U10833 (N_10833,N_6819,N_6650);
xnor U10834 (N_10834,N_1326,N_8732);
and U10835 (N_10835,N_7487,N_9053);
or U10836 (N_10836,N_2844,N_3038);
or U10837 (N_10837,N_7780,N_3054);
and U10838 (N_10838,N_6550,N_9978);
or U10839 (N_10839,N_7896,N_9290);
nor U10840 (N_10840,N_7908,N_8929);
nor U10841 (N_10841,N_2049,N_6717);
nand U10842 (N_10842,N_8270,N_3619);
nor U10843 (N_10843,N_3388,N_7139);
and U10844 (N_10844,N_3234,N_672);
or U10845 (N_10845,N_6418,N_1705);
or U10846 (N_10846,N_5163,N_3936);
nor U10847 (N_10847,N_9114,N_2804);
nand U10848 (N_10848,N_4009,N_9385);
nand U10849 (N_10849,N_5814,N_8925);
and U10850 (N_10850,N_1797,N_5791);
or U10851 (N_10851,N_2378,N_8714);
nor U10852 (N_10852,N_883,N_8059);
xor U10853 (N_10853,N_5365,N_2485);
nand U10854 (N_10854,N_436,N_9445);
and U10855 (N_10855,N_666,N_2011);
nand U10856 (N_10856,N_2115,N_6109);
and U10857 (N_10857,N_9079,N_4744);
xor U10858 (N_10858,N_7526,N_4770);
or U10859 (N_10859,N_1751,N_9649);
and U10860 (N_10860,N_9010,N_2520);
nand U10861 (N_10861,N_7613,N_1035);
xor U10862 (N_10862,N_9775,N_1683);
or U10863 (N_10863,N_5610,N_1723);
and U10864 (N_10864,N_4327,N_2683);
xor U10865 (N_10865,N_8721,N_8293);
or U10866 (N_10866,N_5039,N_7807);
and U10867 (N_10867,N_1223,N_974);
nand U10868 (N_10868,N_1824,N_7670);
or U10869 (N_10869,N_334,N_2376);
nand U10870 (N_10870,N_7172,N_5425);
nor U10871 (N_10871,N_2607,N_997);
nor U10872 (N_10872,N_8989,N_951);
and U10873 (N_10873,N_9361,N_4079);
nand U10874 (N_10874,N_7278,N_590);
xnor U10875 (N_10875,N_4552,N_3178);
nor U10876 (N_10876,N_8874,N_8944);
nor U10877 (N_10877,N_4175,N_8507);
and U10878 (N_10878,N_431,N_4606);
nand U10879 (N_10879,N_9519,N_5879);
and U10880 (N_10880,N_5190,N_7143);
and U10881 (N_10881,N_2760,N_9525);
nand U10882 (N_10882,N_6354,N_9814);
xnor U10883 (N_10883,N_4571,N_2307);
and U10884 (N_10884,N_1908,N_2849);
or U10885 (N_10885,N_1911,N_9902);
or U10886 (N_10886,N_7697,N_9204);
nor U10887 (N_10887,N_8468,N_9647);
or U10888 (N_10888,N_6479,N_9489);
and U10889 (N_10889,N_5491,N_3337);
nand U10890 (N_10890,N_6539,N_3769);
nand U10891 (N_10891,N_836,N_1736);
nand U10892 (N_10892,N_3764,N_986);
and U10893 (N_10893,N_3618,N_6887);
nand U10894 (N_10894,N_6592,N_6528);
and U10895 (N_10895,N_6399,N_4613);
nor U10896 (N_10896,N_1610,N_8102);
and U10897 (N_10897,N_1442,N_4580);
and U10898 (N_10898,N_2906,N_4367);
or U10899 (N_10899,N_8785,N_8945);
and U10900 (N_10900,N_4121,N_8298);
or U10901 (N_10901,N_4595,N_924);
nor U10902 (N_10902,N_2750,N_7061);
and U10903 (N_10903,N_2183,N_9880);
and U10904 (N_10904,N_9894,N_9272);
nand U10905 (N_10905,N_5099,N_4961);
and U10906 (N_10906,N_8754,N_9227);
or U10907 (N_10907,N_4244,N_5723);
and U10908 (N_10908,N_1172,N_6644);
or U10909 (N_10909,N_5014,N_8683);
nor U10910 (N_10910,N_6632,N_3078);
and U10911 (N_10911,N_6041,N_265);
nor U10912 (N_10912,N_2102,N_9754);
and U10913 (N_10913,N_6686,N_8703);
and U10914 (N_10914,N_9046,N_6336);
or U10915 (N_10915,N_5750,N_7097);
nand U10916 (N_10916,N_1128,N_4833);
xnor U10917 (N_10917,N_5646,N_7265);
or U10918 (N_10918,N_9507,N_1496);
nor U10919 (N_10919,N_9700,N_1171);
nand U10920 (N_10920,N_694,N_2914);
nor U10921 (N_10921,N_8064,N_3140);
nor U10922 (N_10922,N_8430,N_6071);
nand U10923 (N_10923,N_8643,N_7812);
or U10924 (N_10924,N_9243,N_1013);
and U10925 (N_10925,N_2466,N_4421);
or U10926 (N_10926,N_8713,N_6890);
nor U10927 (N_10927,N_8864,N_9934);
xnor U10928 (N_10928,N_7524,N_9780);
nand U10929 (N_10929,N_9181,N_2153);
and U10930 (N_10930,N_4042,N_6688);
or U10931 (N_10931,N_6511,N_4799);
nand U10932 (N_10932,N_4779,N_7344);
and U10933 (N_10933,N_5553,N_8243);
nor U10934 (N_10934,N_4589,N_271);
nand U10935 (N_10935,N_6159,N_1793);
nor U10936 (N_10936,N_5984,N_6861);
nand U10937 (N_10937,N_1533,N_3885);
or U10938 (N_10938,N_4560,N_1310);
and U10939 (N_10939,N_4612,N_1849);
and U10940 (N_10940,N_2927,N_4630);
nor U10941 (N_10941,N_5064,N_4721);
or U10942 (N_10942,N_495,N_7088);
nor U10943 (N_10943,N_1475,N_1187);
and U10944 (N_10944,N_9330,N_6358);
or U10945 (N_10945,N_5546,N_9678);
and U10946 (N_10946,N_852,N_7426);
and U10947 (N_10947,N_9225,N_3387);
or U10948 (N_10948,N_1808,N_1994);
or U10949 (N_10949,N_2675,N_6139);
nor U10950 (N_10950,N_8536,N_2803);
or U10951 (N_10951,N_6475,N_6140);
or U10952 (N_10952,N_2774,N_8667);
xnor U10953 (N_10953,N_2269,N_6355);
and U10954 (N_10954,N_7511,N_7886);
and U10955 (N_10955,N_5753,N_2208);
nand U10956 (N_10956,N_5890,N_1660);
or U10957 (N_10957,N_9209,N_2616);
and U10958 (N_10958,N_1344,N_5994);
nand U10959 (N_10959,N_7351,N_9798);
or U10960 (N_10960,N_9023,N_5198);
nor U10961 (N_10961,N_1416,N_4918);
xnor U10962 (N_10962,N_3524,N_6643);
and U10963 (N_10963,N_2649,N_301);
nor U10964 (N_10964,N_8160,N_1902);
and U10965 (N_10965,N_5884,N_3539);
xor U10966 (N_10966,N_2703,N_4262);
and U10967 (N_10967,N_4395,N_6183);
nor U10968 (N_10968,N_6804,N_6204);
and U10969 (N_10969,N_7719,N_2822);
xor U10970 (N_10970,N_4722,N_6468);
and U10971 (N_10971,N_5166,N_1620);
nor U10972 (N_10972,N_9778,N_710);
nor U10973 (N_10973,N_5666,N_5154);
nand U10974 (N_10974,N_3499,N_3011);
nor U10975 (N_10975,N_4897,N_6518);
nor U10976 (N_10976,N_2364,N_1078);
and U10977 (N_10977,N_2287,N_1757);
nor U10978 (N_10978,N_7328,N_2795);
and U10979 (N_10979,N_287,N_7242);
nand U10980 (N_10980,N_6969,N_5378);
and U10981 (N_10981,N_6894,N_5233);
or U10982 (N_10982,N_392,N_6618);
nor U10983 (N_10983,N_6283,N_6918);
xor U10984 (N_10984,N_2481,N_9884);
xnor U10985 (N_10985,N_4926,N_7123);
and U10986 (N_10986,N_6043,N_779);
nand U10987 (N_10987,N_8191,N_8333);
or U10988 (N_10988,N_2572,N_8666);
nor U10989 (N_10989,N_1189,N_6318);
nor U10990 (N_10990,N_1145,N_11);
nand U10991 (N_10991,N_189,N_3857);
nand U10992 (N_10992,N_2697,N_1127);
nand U10993 (N_10993,N_6345,N_3169);
and U10994 (N_10994,N_3703,N_2826);
and U10995 (N_10995,N_4731,N_167);
nor U10996 (N_10996,N_64,N_9165);
nor U10997 (N_10997,N_9465,N_6123);
nor U10998 (N_10998,N_538,N_4702);
or U10999 (N_10999,N_346,N_8673);
xor U11000 (N_11000,N_8723,N_2654);
nor U11001 (N_11001,N_4193,N_9951);
nor U11002 (N_11002,N_5146,N_7783);
nor U11003 (N_11003,N_5745,N_7951);
xnor U11004 (N_11004,N_724,N_6557);
or U11005 (N_11005,N_3978,N_7820);
or U11006 (N_11006,N_8656,N_9695);
nand U11007 (N_11007,N_8104,N_2258);
or U11008 (N_11008,N_3721,N_7924);
nand U11009 (N_11009,N_2352,N_6729);
or U11010 (N_11010,N_6927,N_3118);
or U11011 (N_11011,N_1232,N_3358);
nor U11012 (N_11012,N_5803,N_8444);
nand U11013 (N_11013,N_8483,N_4313);
nand U11014 (N_11014,N_1693,N_6015);
and U11015 (N_11015,N_7050,N_5679);
nand U11016 (N_11016,N_8147,N_4865);
or U11017 (N_11017,N_7562,N_4104);
nor U11018 (N_11018,N_3154,N_8060);
and U11019 (N_11019,N_5936,N_3840);
and U11020 (N_11020,N_2733,N_9834);
nand U11021 (N_11021,N_2095,N_7778);
and U11022 (N_11022,N_321,N_324);
nand U11023 (N_11023,N_185,N_7614);
nand U11024 (N_11024,N_8453,N_2593);
and U11025 (N_11025,N_4922,N_5693);
xor U11026 (N_11026,N_2869,N_2877);
or U11027 (N_11027,N_2640,N_6560);
nor U11028 (N_11028,N_8276,N_8387);
xor U11029 (N_11029,N_6237,N_2603);
nor U11030 (N_11030,N_2918,N_6383);
and U11031 (N_11031,N_613,N_7769);
and U11032 (N_11032,N_1787,N_3889);
nor U11033 (N_11033,N_6446,N_6180);
nand U11034 (N_11034,N_1916,N_5888);
nor U11035 (N_11035,N_887,N_7764);
or U11036 (N_11036,N_2850,N_22);
nor U11037 (N_11037,N_7582,N_9491);
and U11038 (N_11038,N_4363,N_343);
and U11039 (N_11039,N_987,N_1954);
nand U11040 (N_11040,N_4951,N_8400);
or U11041 (N_11041,N_595,N_9328);
nand U11042 (N_11042,N_2404,N_6527);
and U11043 (N_11043,N_9530,N_849);
and U11044 (N_11044,N_2735,N_2792);
nor U11045 (N_11045,N_2586,N_9375);
xor U11046 (N_11046,N_749,N_726);
nor U11047 (N_11047,N_2815,N_6631);
nand U11048 (N_11048,N_8566,N_4083);
nor U11049 (N_11049,N_4196,N_6268);
nor U11050 (N_11050,N_2612,N_8835);
and U11051 (N_11051,N_5269,N_1012);
and U11052 (N_11052,N_5287,N_6703);
nand U11053 (N_11053,N_8185,N_3391);
nand U11054 (N_11054,N_5431,N_2263);
nand U11055 (N_11055,N_1939,N_955);
or U11056 (N_11056,N_8767,N_6537);
nor U11057 (N_11057,N_150,N_3268);
nand U11058 (N_11058,N_8576,N_9915);
and U11059 (N_11059,N_4850,N_5627);
nand U11060 (N_11060,N_7869,N_8915);
nor U11061 (N_11061,N_6980,N_952);
nor U11062 (N_11062,N_3864,N_580);
nand U11063 (N_11063,N_4726,N_6254);
xor U11064 (N_11064,N_500,N_2207);
xnor U11065 (N_11065,N_1134,N_7628);
xnor U11066 (N_11066,N_6145,N_8890);
xnor U11067 (N_11067,N_4464,N_2081);
or U11068 (N_11068,N_8007,N_95);
nor U11069 (N_11069,N_5794,N_3635);
nor U11070 (N_11070,N_6671,N_2027);
nand U11071 (N_11071,N_3273,N_6033);
xor U11072 (N_11072,N_4264,N_1377);
nor U11073 (N_11073,N_3403,N_6162);
and U11074 (N_11074,N_8691,N_70);
nor U11075 (N_11075,N_6437,N_2338);
and U11076 (N_11076,N_6390,N_2618);
or U11077 (N_11077,N_3861,N_124);
or U11078 (N_11078,N_6515,N_7865);
and U11079 (N_11079,N_3620,N_1200);
or U11080 (N_11080,N_7715,N_61);
nor U11081 (N_11081,N_5469,N_59);
or U11082 (N_11082,N_6320,N_8155);
and U11083 (N_11083,N_2775,N_8233);
xnor U11084 (N_11084,N_7206,N_2225);
nor U11085 (N_11085,N_6611,N_4308);
and U11086 (N_11086,N_2662,N_8857);
or U11087 (N_11087,N_4465,N_7026);
nand U11088 (N_11088,N_4781,N_9663);
nand U11089 (N_11089,N_4489,N_2322);
and U11090 (N_11090,N_8641,N_4797);
nand U11091 (N_11091,N_3727,N_3640);
or U11092 (N_11092,N_4703,N_2785);
nor U11093 (N_11093,N_4631,N_4968);
nand U11094 (N_11094,N_966,N_745);
and U11095 (N_11095,N_2479,N_8784);
nor U11096 (N_11096,N_4394,N_281);
and U11097 (N_11097,N_8378,N_6889);
nor U11098 (N_11098,N_9104,N_7110);
nor U11099 (N_11099,N_6275,N_3636);
or U11100 (N_11100,N_3723,N_4415);
nor U11101 (N_11101,N_928,N_6284);
nor U11102 (N_11102,N_634,N_2546);
nand U11103 (N_11103,N_9089,N_6884);
nand U11104 (N_11104,N_8238,N_8223);
or U11105 (N_11105,N_7832,N_5178);
or U11106 (N_11106,N_4657,N_7902);
nand U11107 (N_11107,N_2147,N_2016);
nor U11108 (N_11108,N_9670,N_5976);
xor U11109 (N_11109,N_9449,N_4135);
or U11110 (N_11110,N_4825,N_7404);
nor U11111 (N_11111,N_3783,N_239);
and U11112 (N_11112,N_7508,N_1828);
or U11113 (N_11113,N_8282,N_6232);
nor U11114 (N_11114,N_3753,N_7929);
and U11115 (N_11115,N_3472,N_6006);
or U11116 (N_11116,N_3626,N_5424);
nand U11117 (N_11117,N_4780,N_4451);
or U11118 (N_11118,N_330,N_3767);
or U11119 (N_11119,N_3208,N_7658);
nand U11120 (N_11120,N_6563,N_1965);
and U11121 (N_11121,N_5366,N_5415);
xor U11122 (N_11122,N_235,N_9581);
nand U11123 (N_11123,N_8503,N_6967);
and U11124 (N_11124,N_351,N_5391);
or U11125 (N_11125,N_5276,N_4764);
nand U11126 (N_11126,N_369,N_3315);
xor U11127 (N_11127,N_8357,N_58);
xnor U11128 (N_11128,N_855,N_6245);
or U11129 (N_11129,N_110,N_1947);
nor U11130 (N_11130,N_782,N_3711);
and U11131 (N_11131,N_7539,N_5999);
nor U11132 (N_11132,N_5428,N_2597);
xnor U11133 (N_11133,N_4115,N_7638);
or U11134 (N_11134,N_99,N_6705);
nand U11135 (N_11135,N_3665,N_6654);
xnor U11136 (N_11136,N_3257,N_8828);
nand U11137 (N_11137,N_759,N_5471);
or U11138 (N_11138,N_9878,N_512);
xnor U11139 (N_11139,N_1016,N_8816);
nand U11140 (N_11140,N_102,N_1876);
and U11141 (N_11141,N_9761,N_5800);
nor U11142 (N_11142,N_8348,N_2818);
nor U11143 (N_11143,N_8534,N_9992);
or U11144 (N_11144,N_2308,N_9159);
or U11145 (N_11145,N_801,N_3515);
nor U11146 (N_11146,N_9689,N_8475);
and U11147 (N_11147,N_9106,N_5707);
and U11148 (N_11148,N_8210,N_7170);
and U11149 (N_11149,N_3318,N_680);
and U11150 (N_11150,N_8700,N_5057);
xnor U11151 (N_11151,N_699,N_1529);
nor U11152 (N_11152,N_2759,N_7754);
nor U11153 (N_11153,N_4563,N_3624);
xor U11154 (N_11154,N_5260,N_9258);
and U11155 (N_11155,N_8076,N_1970);
nor U11156 (N_11156,N_4466,N_5837);
nand U11157 (N_11157,N_3027,N_3811);
or U11158 (N_11158,N_9418,N_9325);
nand U11159 (N_11159,N_8077,N_1240);
or U11160 (N_11160,N_7484,N_8770);
and U11161 (N_11161,N_6296,N_2891);
nor U11162 (N_11162,N_1682,N_2965);
or U11163 (N_11163,N_6937,N_84);
or U11164 (N_11164,N_3164,N_7277);
and U11165 (N_11165,N_5140,N_8283);
or U11166 (N_11166,N_2087,N_1825);
xnor U11167 (N_11167,N_3195,N_1030);
and U11168 (N_11168,N_2638,N_5660);
or U11169 (N_11169,N_6286,N_5141);
and U11170 (N_11170,N_8189,N_435);
nand U11171 (N_11171,N_2799,N_3052);
and U11172 (N_11172,N_6042,N_3495);
nor U11173 (N_11173,N_1402,N_9394);
or U11174 (N_11174,N_3336,N_1275);
or U11175 (N_11175,N_9158,N_8355);
or U11176 (N_11176,N_7420,N_5714);
and U11177 (N_11177,N_2467,N_4678);
or U11178 (N_11178,N_4877,N_3126);
nand U11179 (N_11179,N_6753,N_3456);
nand U11180 (N_11180,N_3730,N_5719);
nand U11181 (N_11181,N_270,N_6849);
nand U11182 (N_11182,N_8975,N_3686);
and U11183 (N_11183,N_6397,N_416);
and U11184 (N_11184,N_9825,N_6778);
or U11185 (N_11185,N_1348,N_5824);
and U11186 (N_11186,N_1430,N_667);
nor U11187 (N_11187,N_2416,N_7002);
nor U11188 (N_11188,N_8809,N_3305);
nand U11189 (N_11189,N_315,N_984);
nand U11190 (N_11190,N_1927,N_1363);
nand U11191 (N_11191,N_6699,N_9407);
nand U11192 (N_11192,N_4374,N_8019);
nor U11193 (N_11193,N_3148,N_4117);
nor U11194 (N_11194,N_6369,N_1473);
nand U11195 (N_11195,N_161,N_2576);
nor U11196 (N_11196,N_8088,N_3360);
or U11197 (N_11197,N_2099,N_3048);
or U11198 (N_11198,N_9987,N_5117);
nand U11199 (N_11199,N_591,N_9440);
and U11200 (N_11200,N_7263,N_6978);
and U11201 (N_11201,N_9472,N_1968);
nor U11202 (N_11202,N_5765,N_6282);
or U11203 (N_11203,N_4259,N_6674);
and U11204 (N_11204,N_6578,N_7401);
nand U11205 (N_11205,N_4971,N_8833);
nand U11206 (N_11206,N_363,N_8108);
or U11207 (N_11207,N_5885,N_2149);
nand U11208 (N_11208,N_4603,N_7467);
nand U11209 (N_11209,N_3813,N_3041);
nor U11210 (N_11210,N_1452,N_3692);
xor U11211 (N_11211,N_8281,N_9398);
or U11212 (N_11212,N_9531,N_1749);
and U11213 (N_11213,N_2051,N_5804);
nor U11214 (N_11214,N_3507,N_8931);
or U11215 (N_11215,N_9651,N_8867);
nand U11216 (N_11216,N_2575,N_4474);
nor U11217 (N_11217,N_9813,N_6846);
or U11218 (N_11218,N_9305,N_2820);
or U11219 (N_11219,N_7656,N_8226);
and U11220 (N_11220,N_1195,N_5594);
or U11221 (N_11221,N_1833,N_1741);
and U11222 (N_11222,N_2173,N_9559);
xor U11223 (N_11223,N_6331,N_6074);
or U11224 (N_11224,N_7583,N_264);
and U11225 (N_11225,N_5954,N_2955);
or U11226 (N_11226,N_1982,N_2581);
or U11227 (N_11227,N_9211,N_688);
or U11228 (N_11228,N_1521,N_8128);
and U11229 (N_11229,N_3659,N_3847);
nand U11230 (N_11230,N_6313,N_7931);
nor U11231 (N_11231,N_3612,N_5906);
nor U11232 (N_11232,N_9605,N_3757);
nor U11233 (N_11233,N_7029,N_2556);
nor U11234 (N_11234,N_4506,N_1717);
or U11235 (N_11235,N_9535,N_3716);
nand U11236 (N_11236,N_3093,N_5387);
nor U11237 (N_11237,N_3386,N_6953);
nand U11238 (N_11238,N_1130,N_4330);
or U11239 (N_11239,N_6239,N_5760);
and U11240 (N_11240,N_3547,N_8132);
xor U11241 (N_11241,N_5559,N_9835);
and U11242 (N_11242,N_5313,N_6445);
nor U11243 (N_11243,N_1215,N_6172);
and U11244 (N_11244,N_8841,N_1516);
and U11245 (N_11245,N_2437,N_9194);
nand U11246 (N_11246,N_5839,N_5739);
nor U11247 (N_11247,N_3798,N_9665);
and U11248 (N_11248,N_1509,N_9435);
nand U11249 (N_11249,N_8199,N_8426);
and U11250 (N_11250,N_4216,N_8322);
xor U11251 (N_11251,N_3187,N_7051);
and U11252 (N_11252,N_3867,N_6256);
xnor U11253 (N_11253,N_4574,N_1297);
and U11254 (N_11254,N_2110,N_7048);
nand U11255 (N_11255,N_8288,N_1900);
and U11256 (N_11256,N_5640,N_2657);
or U11257 (N_11257,N_7159,N_8353);
nand U11258 (N_11258,N_5937,N_53);
xor U11259 (N_11259,N_4628,N_1933);
and U11260 (N_11260,N_26,N_100);
xnor U11261 (N_11261,N_1584,N_4905);
xor U11262 (N_11262,N_5531,N_6943);
xnor U11263 (N_11263,N_2427,N_9215);
and U11264 (N_11264,N_5569,N_776);
and U11265 (N_11265,N_8896,N_3528);
nand U11266 (N_11266,N_3504,N_1357);
xnor U11267 (N_11267,N_383,N_9206);
nand U11268 (N_11268,N_9073,N_6983);
nor U11269 (N_11269,N_8581,N_2327);
nand U11270 (N_11270,N_6083,N_2141);
nand U11271 (N_11271,N_3142,N_5089);
nand U11272 (N_11272,N_5515,N_5619);
and U11273 (N_11273,N_6409,N_2428);
nor U11274 (N_11274,N_6166,N_2824);
xor U11275 (N_11275,N_7800,N_1216);
or U11276 (N_11276,N_8520,N_4556);
nand U11277 (N_11277,N_7259,N_6900);
and U11278 (N_11278,N_476,N_9827);
and U11279 (N_11279,N_5854,N_1587);
nor U11280 (N_11280,N_5724,N_4843);
and U11281 (N_11281,N_2328,N_4151);
and U11282 (N_11282,N_356,N_8616);
nand U11283 (N_11283,N_7903,N_6417);
nand U11284 (N_11284,N_276,N_2990);
nand U11285 (N_11285,N_4340,N_3144);
or U11286 (N_11286,N_8107,N_4567);
and U11287 (N_11287,N_8670,N_2847);
nor U11288 (N_11288,N_6349,N_1114);
and U11289 (N_11289,N_5136,N_9464);
nor U11290 (N_11290,N_5373,N_9593);
and U11291 (N_11291,N_5715,N_842);
nor U11292 (N_11292,N_352,N_6373);
or U11293 (N_11293,N_2425,N_5688);
or U11294 (N_11294,N_1588,N_2911);
nand U11295 (N_11295,N_9186,N_1379);
nand U11296 (N_11296,N_1330,N_6744);
and U11297 (N_11297,N_1891,N_4127);
nand U11298 (N_11298,N_9064,N_4751);
and U11299 (N_11299,N_7154,N_9236);
and U11300 (N_11300,N_5630,N_651);
xnor U11301 (N_11301,N_8980,N_3819);
nor U11302 (N_11302,N_1197,N_5041);
or U11303 (N_11303,N_170,N_7689);
and U11304 (N_11304,N_3121,N_2349);
or U11305 (N_11305,N_1064,N_1886);
nand U11306 (N_11306,N_4526,N_4211);
or U11307 (N_11307,N_2047,N_9022);
or U11308 (N_11308,N_206,N_2232);
xnor U11309 (N_11309,N_638,N_4609);
xnor U11310 (N_11310,N_215,N_9771);
or U11311 (N_11311,N_2442,N_4879);
nor U11312 (N_11312,N_8829,N_7934);
xnor U11313 (N_11313,N_6224,N_4733);
xnor U11314 (N_11314,N_3585,N_32);
nor U11315 (N_11315,N_3945,N_9860);
and U11316 (N_11316,N_1545,N_4982);
or U11317 (N_11317,N_3028,N_4443);
xnor U11318 (N_11318,N_1653,N_2659);
nand U11319 (N_11319,N_1830,N_9584);
nand U11320 (N_11320,N_9794,N_5740);
and U11321 (N_11321,N_6453,N_5394);
nand U11322 (N_11322,N_1208,N_979);
and U11323 (N_11323,N_4003,N_7774);
nor U11324 (N_11324,N_6805,N_7432);
or U11325 (N_11325,N_1302,N_9202);
nand U11326 (N_11326,N_8247,N_705);
nor U11327 (N_11327,N_9276,N_3974);
nor U11328 (N_11328,N_1857,N_1350);
nand U11329 (N_11329,N_4579,N_3251);
or U11330 (N_11330,N_775,N_9891);
or U11331 (N_11331,N_6796,N_6873);
nor U11332 (N_11332,N_7232,N_5013);
or U11333 (N_11333,N_5034,N_9162);
nand U11334 (N_11334,N_5749,N_8979);
nand U11335 (N_11335,N_8802,N_8967);
or U11336 (N_11336,N_5539,N_1352);
and U11337 (N_11337,N_832,N_8359);
nand U11338 (N_11338,N_1300,N_1532);
or U11339 (N_11339,N_6800,N_2617);
and U11340 (N_11340,N_1507,N_3037);
and U11341 (N_11341,N_6761,N_9546);
or U11342 (N_11342,N_2045,N_9576);
nand U11343 (N_11343,N_1307,N_2790);
or U11344 (N_11344,N_313,N_1845);
nand U11345 (N_11345,N_4619,N_5257);
and U11346 (N_11346,N_973,N_6335);
xnor U11347 (N_11347,N_7168,N_746);
nor U11348 (N_11348,N_130,N_8351);
and U11349 (N_11349,N_2365,N_9921);
and U11350 (N_11350,N_3264,N_6427);
nor U11351 (N_11351,N_3591,N_5656);
xnor U11352 (N_11352,N_1087,N_2550);
nor U11353 (N_11353,N_6067,N_9566);
or U11354 (N_11354,N_4249,N_2363);
nor U11355 (N_11355,N_3135,N_7175);
and U11356 (N_11356,N_1559,N_1957);
nor U11357 (N_11357,N_4623,N_7791);
and U11358 (N_11358,N_8647,N_1585);
or U11359 (N_11359,N_4640,N_9580);
nor U11360 (N_11360,N_8603,N_8273);
or U11361 (N_11361,N_4679,N_3219);
xor U11362 (N_11362,N_8617,N_5734);
and U11363 (N_11363,N_713,N_3239);
nand U11364 (N_11364,N_1413,N_7817);
nor U11365 (N_11365,N_5761,N_1776);
nand U11366 (N_11366,N_1435,N_2052);
nand U11367 (N_11367,N_2222,N_4845);
and U11368 (N_11368,N_9541,N_2449);
nand U11369 (N_11369,N_6769,N_8604);
or U11370 (N_11370,N_7412,N_8290);
or U11371 (N_11371,N_5901,N_2499);
nor U11372 (N_11372,N_4573,N_9002);
and U11373 (N_11373,N_1996,N_7101);
nand U11374 (N_11374,N_8285,N_840);
nor U11375 (N_11375,N_303,N_1768);
nand U11376 (N_11376,N_5700,N_5453);
and U11377 (N_11377,N_3737,N_1451);
nor U11378 (N_11378,N_8087,N_497);
and U11379 (N_11379,N_6334,N_3697);
nand U11380 (N_11380,N_7356,N_379);
nand U11381 (N_11381,N_4245,N_9882);
and U11382 (N_11382,N_2046,N_1695);
or U11383 (N_11383,N_2527,N_9823);
nor U11384 (N_11384,N_2006,N_135);
or U11385 (N_11385,N_9765,N_9932);
or U11386 (N_11386,N_6000,N_3773);
and U11387 (N_11387,N_5296,N_439);
nand U11388 (N_11388,N_4427,N_7021);
nor U11389 (N_11389,N_6046,N_2165);
nor U11390 (N_11390,N_6241,N_5522);
nor U11391 (N_11391,N_4198,N_3937);
and U11392 (N_11392,N_7542,N_1433);
nor U11393 (N_11393,N_2687,N_5674);
nor U11394 (N_11394,N_1301,N_7047);
nor U11395 (N_11395,N_9692,N_3615);
and U11396 (N_11396,N_8788,N_5782);
or U11397 (N_11397,N_8245,N_94);
and U11398 (N_11398,N_7750,N_2451);
nor U11399 (N_11399,N_2598,N_1320);
and U11400 (N_11400,N_9237,N_5673);
nor U11401 (N_11401,N_1774,N_8335);
nand U11402 (N_11402,N_4002,N_2343);
nand U11403 (N_11403,N_2636,N_4032);
and U11404 (N_11404,N_4050,N_3766);
and U11405 (N_11405,N_9191,N_9406);
or U11406 (N_11406,N_401,N_8260);
nor U11407 (N_11407,N_3735,N_3576);
nor U11408 (N_11408,N_3500,N_2696);
nand U11409 (N_11409,N_505,N_1553);
nor U11410 (N_11410,N_7439,N_8241);
or U11411 (N_11411,N_1575,N_3359);
and U11412 (N_11412,N_7686,N_3080);
and U11413 (N_11413,N_4826,N_5474);
nand U11414 (N_11414,N_8206,N_8861);
xor U11415 (N_11415,N_8947,N_2777);
or U11416 (N_11416,N_6424,N_7114);
or U11417 (N_11417,N_4052,N_5095);
or U11418 (N_11418,N_7435,N_3662);
and U11419 (N_11419,N_2114,N_163);
nand U11420 (N_11420,N_990,N_3097);
or U11421 (N_11421,N_7109,N_7438);
and U11422 (N_11422,N_8325,N_2910);
nand U11423 (N_11423,N_522,N_4228);
nor U11424 (N_11424,N_9421,N_3824);
xor U11425 (N_11425,N_3404,N_1073);
nor U11426 (N_11426,N_3146,N_3808);
nor U11427 (N_11427,N_6396,N_9147);
nor U11428 (N_11428,N_2073,N_9623);
nand U11429 (N_11429,N_9629,N_6721);
nand U11430 (N_11430,N_7985,N_5195);
and U11431 (N_11431,N_9311,N_3560);
and U11432 (N_11432,N_5871,N_8135);
nand U11433 (N_11433,N_8801,N_1688);
nor U11434 (N_11434,N_508,N_253);
xnor U11435 (N_11435,N_6990,N_3152);
nor U11436 (N_11436,N_2570,N_2478);
nand U11437 (N_11437,N_7881,N_1203);
xnor U11438 (N_11438,N_7397,N_639);
and U11439 (N_11439,N_2033,N_4839);
and U11440 (N_11440,N_2158,N_5002);
nor U11441 (N_11441,N_8898,N_7343);
xnor U11442 (N_11442,N_8924,N_2105);
and U11443 (N_11443,N_9164,N_8115);
nand U11444 (N_11444,N_6347,N_4933);
or U11445 (N_11445,N_8110,N_7761);
or U11446 (N_11446,N_9461,N_8432);
nor U11447 (N_11447,N_2262,N_8354);
nand U11448 (N_11448,N_6862,N_7649);
nand U11449 (N_11449,N_8532,N_6258);
or U11450 (N_11450,N_1563,N_8685);
nand U11451 (N_11451,N_6575,N_5403);
and U11452 (N_11452,N_5614,N_6247);
nand U11453 (N_11453,N_339,N_6583);
nand U11454 (N_11454,N_7577,N_5621);
or U11455 (N_11455,N_186,N_3477);
or U11456 (N_11456,N_3468,N_9833);
or U11457 (N_11457,N_1488,N_9955);
or U11458 (N_11458,N_2241,N_295);
or U11459 (N_11459,N_214,N_8882);
and U11460 (N_11460,N_9896,N_5316);
nand U11461 (N_11461,N_5701,N_1094);
or U11462 (N_11462,N_4710,N_2720);
nand U11463 (N_11463,N_9460,N_6877);
and U11464 (N_11464,N_7510,N_279);
or U11465 (N_11465,N_3892,N_930);
nor U11466 (N_11466,N_9266,N_8533);
nor U11467 (N_11467,N_555,N_5599);
nand U11468 (N_11468,N_12,N_143);
nor U11469 (N_11469,N_3288,N_4593);
and U11470 (N_11470,N_5856,N_2893);
nor U11471 (N_11471,N_6430,N_5206);
and U11472 (N_11472,N_8677,N_5130);
or U11473 (N_11473,N_8114,N_9981);
nor U11474 (N_11474,N_4642,N_1129);
nand U11475 (N_11475,N_5133,N_9636);
or U11476 (N_11476,N_2243,N_4390);
nor U11477 (N_11477,N_2072,N_4436);
and U11478 (N_11478,N_1556,N_9850);
nor U11479 (N_11479,N_3561,N_1583);
nand U11480 (N_11480,N_5337,N_6561);
nand U11481 (N_11481,N_190,N_1494);
or U11482 (N_11482,N_2978,N_9140);
or U11483 (N_11483,N_4355,N_7848);
and U11484 (N_11484,N_4207,N_4299);
or U11485 (N_11485,N_6713,N_2944);
nand U11486 (N_11486,N_9287,N_3454);
nor U11487 (N_11487,N_2313,N_3417);
and U11488 (N_11488,N_5392,N_5922);
nand U11489 (N_11489,N_4798,N_2717);
and U11490 (N_11490,N_9522,N_1589);
nor U11491 (N_11491,N_2491,N_9553);
or U11492 (N_11492,N_7309,N_8872);
and U11493 (N_11493,N_1875,N_7831);
nor U11494 (N_11494,N_9976,N_9216);
or U11495 (N_11495,N_8524,N_8081);
and U11496 (N_11496,N_3055,N_9899);
or U11497 (N_11497,N_7145,N_5963);
and U11498 (N_11498,N_1773,N_471);
nor U11499 (N_11499,N_491,N_6948);
xnor U11500 (N_11500,N_894,N_822);
xnor U11501 (N_11501,N_7319,N_1552);
or U11502 (N_11502,N_6825,N_1093);
or U11503 (N_11503,N_2274,N_5410);
or U11504 (N_11504,N_1101,N_3145);
nand U11505 (N_11505,N_2074,N_3439);
nand U11506 (N_11506,N_7382,N_2917);
nand U11507 (N_11507,N_994,N_4569);
nand U11508 (N_11508,N_3475,N_5582);
and U11509 (N_11509,N_5597,N_6133);
nor U11510 (N_11510,N_4231,N_7597);
nand U11511 (N_11511,N_4166,N_3425);
and U11512 (N_11512,N_3944,N_921);
nor U11513 (N_11513,N_7204,N_6817);
and U11514 (N_11514,N_9205,N_8883);
or U11515 (N_11515,N_706,N_3531);
and U11516 (N_11516,N_3722,N_9190);
and U11517 (N_11517,N_3890,N_8588);
nor U11518 (N_11518,N_4329,N_3810);
and U11519 (N_11519,N_2634,N_2118);
and U11520 (N_11520,N_1152,N_3238);
xor U11521 (N_11521,N_1572,N_5452);
nor U11522 (N_11522,N_4456,N_5230);
nor U11523 (N_11523,N_8969,N_6875);
nor U11524 (N_11524,N_4004,N_9129);
nand U11525 (N_11525,N_1622,N_4140);
nand U11526 (N_11526,N_9862,N_5556);
or U11527 (N_11527,N_1960,N_7296);
or U11528 (N_11528,N_9763,N_7445);
or U11529 (N_11529,N_7966,N_3066);
or U11530 (N_11530,N_9050,N_9120);
nor U11531 (N_11531,N_1645,N_900);
or U11532 (N_11532,N_1178,N_4790);
nor U11533 (N_11533,N_5858,N_8564);
or U11534 (N_11534,N_1694,N_6989);
xnor U11535 (N_11535,N_8448,N_5895);
nor U11536 (N_11536,N_2188,N_4507);
nand U11537 (N_11537,N_2044,N_3252);
or U11538 (N_11538,N_1182,N_4816);
xor U11539 (N_11539,N_7810,N_2700);
nand U11540 (N_11540,N_9662,N_3225);
and U11541 (N_11541,N_9906,N_5100);
nand U11542 (N_11542,N_8768,N_7979);
and U11543 (N_11543,N_9711,N_209);
and U11544 (N_11544,N_7722,N_1218);
and U11545 (N_11545,N_8074,N_5016);
or U11546 (N_11546,N_6553,N_743);
nand U11547 (N_11547,N_7990,N_8722);
or U11548 (N_11548,N_6073,N_5993);
nand U11549 (N_11549,N_423,N_4511);
nand U11550 (N_11550,N_7112,N_1765);
nand U11551 (N_11551,N_65,N_5577);
and U11552 (N_11552,N_3693,N_6860);
xor U11553 (N_11553,N_6762,N_8842);
nand U11554 (N_11554,N_517,N_9781);
nand U11555 (N_11555,N_9136,N_7568);
nand U11556 (N_11556,N_5437,N_9038);
nor U11557 (N_11557,N_9968,N_4183);
nand U11558 (N_11558,N_9196,N_7927);
or U11559 (N_11559,N_3302,N_9043);
or U11560 (N_11560,N_9603,N_6116);
or U11561 (N_11561,N_9241,N_2048);
or U11562 (N_11562,N_2539,N_8627);
nand U11563 (N_11563,N_5395,N_3694);
or U11564 (N_11564,N_2224,N_3159);
and U11565 (N_11565,N_1806,N_7153);
nand U11566 (N_11566,N_4760,N_1250);
nand U11567 (N_11567,N_2673,N_3975);
nand U11568 (N_11568,N_6090,N_3990);
nand U11569 (N_11569,N_3775,N_3657);
nand U11570 (N_11570,N_5593,N_656);
nand U11571 (N_11571,N_1382,N_5499);
nand U11572 (N_11572,N_5286,N_3222);
nor U11573 (N_11573,N_7236,N_6264);
or U11574 (N_11574,N_4440,N_1351);
and U11575 (N_11575,N_6127,N_9433);
nor U11576 (N_11576,N_4337,N_9877);
or U11577 (N_11577,N_1265,N_6216);
or U11578 (N_11578,N_201,N_2340);
and U11579 (N_11579,N_5498,N_8909);
xor U11580 (N_11580,N_1193,N_8552);
nor U11581 (N_11581,N_4187,N_9547);
nand U11582 (N_11582,N_488,N_2872);
nor U11583 (N_11583,N_1298,N_2137);
xor U11584 (N_11584,N_9299,N_8366);
xor U11585 (N_11585,N_9866,N_4847);
nor U11586 (N_11586,N_5910,N_8580);
nor U11587 (N_11587,N_7211,N_7149);
and U11588 (N_11588,N_1667,N_3201);
nand U11589 (N_11589,N_9297,N_7253);
or U11590 (N_11590,N_501,N_7327);
and U11591 (N_11591,N_2101,N_2901);
and U11592 (N_11592,N_9514,N_4147);
or U11593 (N_11593,N_7398,N_7368);
and U11594 (N_11594,N_4888,N_473);
and U11595 (N_11595,N_9591,N_4131);
and U11596 (N_11596,N_7495,N_6372);
nor U11597 (N_11597,N_2886,N_1158);
nand U11598 (N_11598,N_8812,N_4765);
xnor U11599 (N_11599,N_5191,N_8469);
nand U11600 (N_11600,N_3771,N_2943);
nand U11601 (N_11601,N_5098,N_327);
or U11602 (N_11602,N_896,N_9447);
nand U11603 (N_11603,N_7906,N_2156);
nand U11604 (N_11604,N_9124,N_1306);
xnor U11605 (N_11605,N_6904,N_4596);
and U11606 (N_11606,N_9182,N_2133);
nand U11607 (N_11607,N_7079,N_1175);
xnor U11608 (N_11608,N_6434,N_4761);
nand U11609 (N_11609,N_3293,N_250);
nor U11610 (N_11610,N_5617,N_7916);
xor U11611 (N_11611,N_3873,N_9637);
and U11612 (N_11612,N_6300,N_5955);
and U11613 (N_11613,N_516,N_875);
nand U11614 (N_11614,N_8186,N_9193);
nor U11615 (N_11615,N_9698,N_3869);
nor U11616 (N_11616,N_1089,N_4840);
nand U11617 (N_11617,N_5160,N_354);
and U11618 (N_11618,N_2736,N_1631);
nor U11619 (N_11619,N_7207,N_1657);
and U11620 (N_11620,N_7766,N_2117);
or U11621 (N_11621,N_7729,N_5855);
or U11622 (N_11622,N_7842,N_3084);
nand U11623 (N_11623,N_5501,N_809);
nand U11624 (N_11624,N_582,N_2396);
or U11625 (N_11625,N_1123,N_7907);
xor U11626 (N_11626,N_4916,N_9057);
or U11627 (N_11627,N_5282,N_3042);
xor U11628 (N_11628,N_7771,N_326);
or U11629 (N_11629,N_2330,N_5938);
or U11630 (N_11630,N_4025,N_5171);
nand U11631 (N_11631,N_1579,N_3968);
or U11632 (N_11632,N_2669,N_8037);
or U11633 (N_11633,N_9327,N_2998);
nand U11634 (N_11634,N_6623,N_2168);
nor U11635 (N_11635,N_4082,N_98);
and U11636 (N_11636,N_4965,N_3994);
or U11637 (N_11637,N_3986,N_3117);
nor U11638 (N_11638,N_1400,N_2907);
and U11639 (N_11639,N_5528,N_6119);
and U11640 (N_11640,N_9696,N_6645);
xor U11641 (N_11641,N_2987,N_7395);
nor U11642 (N_11642,N_3923,N_5703);
or U11643 (N_11643,N_5648,N_9685);
xnor U11644 (N_11644,N_377,N_2514);
and U11645 (N_11645,N_4044,N_2764);
nor U11646 (N_11646,N_9760,N_9248);
and U11647 (N_11647,N_7627,N_5825);
and U11648 (N_11648,N_7997,N_3649);
and U11649 (N_11649,N_348,N_9026);
and U11650 (N_11650,N_6332,N_2500);
nor U11651 (N_11651,N_2756,N_8692);
and U11652 (N_11652,N_4717,N_652);
and U11653 (N_11653,N_8496,N_5338);
xnor U11654 (N_11654,N_3568,N_8217);
or U11655 (N_11655,N_8181,N_3901);
and U11656 (N_11656,N_1905,N_3272);
or U11657 (N_11657,N_3310,N_6420);
and U11658 (N_11658,N_8168,N_342);
nand U11659 (N_11659,N_4205,N_6072);
nand U11660 (N_11660,N_8619,N_3328);
and U11661 (N_11661,N_4753,N_6700);
xnor U11662 (N_11662,N_6267,N_1008);
or U11663 (N_11663,N_4967,N_8762);
or U11664 (N_11664,N_3580,N_7486);
nand U11665 (N_11665,N_8638,N_9151);
or U11666 (N_11666,N_4870,N_2722);
or U11667 (N_11667,N_4225,N_7983);
nor U11668 (N_11668,N_1525,N_7364);
nand U11669 (N_11669,N_118,N_1710);
nor U11670 (N_11670,N_2845,N_8124);
and U11671 (N_11671,N_9348,N_9007);
nand U11672 (N_11672,N_5264,N_1704);
nand U11673 (N_11673,N_1279,N_5449);
xnor U11674 (N_11674,N_4667,N_2580);
and U11675 (N_11675,N_8120,N_2782);
nor U11676 (N_11676,N_3610,N_8292);
nand U11677 (N_11677,N_2923,N_8471);
nand U11678 (N_11678,N_18,N_1811);
nor U11679 (N_11679,N_6944,N_1133);
and U11680 (N_11680,N_1619,N_8725);
or U11681 (N_11681,N_6728,N_5368);
and U11682 (N_11682,N_6188,N_3112);
nor U11683 (N_11683,N_6202,N_247);
nor U11684 (N_11684,N_3888,N_5835);
and U11685 (N_11685,N_4306,N_9986);
and U11686 (N_11686,N_7645,N_3898);
xor U11687 (N_11687,N_5254,N_4592);
nor U11688 (N_11688,N_4163,N_4658);
and U11689 (N_11689,N_3241,N_9127);
nor U11690 (N_11690,N_2077,N_216);
or U11691 (N_11691,N_8940,N_4479);
nor U11692 (N_11692,N_2920,N_2004);
xor U11693 (N_11693,N_9558,N_1854);
nand U11694 (N_11694,N_5426,N_8457);
and U11695 (N_11695,N_1985,N_795);
or U11696 (N_11696,N_6924,N_3878);
xnor U11697 (N_11697,N_2120,N_6143);
nor U11698 (N_11698,N_9772,N_1429);
nor U11699 (N_11699,N_7411,N_6687);
or U11700 (N_11700,N_9210,N_6598);
xor U11701 (N_11701,N_1198,N_6582);
nand U11702 (N_11702,N_5843,N_7767);
nand U11703 (N_11703,N_3389,N_3967);
or U11704 (N_11704,N_441,N_357);
nor U11705 (N_11705,N_2900,N_9390);
nand U11706 (N_11706,N_6752,N_4756);
or U11707 (N_11707,N_2545,N_5833);
and U11708 (N_11708,N_7503,N_8640);
xor U11709 (N_11709,N_8876,N_5520);
nand U11710 (N_11710,N_1060,N_5078);
nand U11711 (N_11711,N_8729,N_3872);
or U11712 (N_11712,N_7482,N_668);
or U11713 (N_11713,N_9861,N_5423);
and U11714 (N_11714,N_6036,N_8367);
nor U11715 (N_11715,N_5374,N_9203);
nor U11716 (N_11716,N_1885,N_751);
and U11717 (N_11717,N_5787,N_9141);
or U11718 (N_11718,N_1386,N_4370);
or U11719 (N_11719,N_3821,N_8242);
and U11720 (N_11720,N_3202,N_109);
nor U11721 (N_11721,N_8609,N_4114);
nand U11722 (N_11722,N_6995,N_2017);
or U11723 (N_11723,N_2026,N_6442);
nor U11724 (N_11724,N_4420,N_7723);
xor U11725 (N_11725,N_9937,N_5808);
nand U11726 (N_11726,N_5741,N_6821);
nor U11727 (N_11727,N_7626,N_3009);
or U11728 (N_11728,N_2757,N_9843);
nor U11729 (N_11729,N_4874,N_6426);
nor U11730 (N_11730,N_719,N_9321);
or U11731 (N_11731,N_5204,N_7518);
nand U11732 (N_11732,N_9957,N_4902);
and U11733 (N_11733,N_8570,N_7600);
and U11734 (N_11734,N_3637,N_486);
or U11735 (N_11735,N_3595,N_69);
nor U11736 (N_11736,N_8538,N_6251);
xor U11737 (N_11737,N_7950,N_2032);
nor U11738 (N_11738,N_834,N_7147);
and U11739 (N_11739,N_2386,N_7631);
nand U11740 (N_11740,N_4066,N_720);
nor U11741 (N_11741,N_5721,N_3002);
and U11742 (N_11742,N_1025,N_3537);
nor U11743 (N_11743,N_6408,N_6415);
nor U11744 (N_11744,N_4484,N_6494);
nand U11745 (N_11745,N_6836,N_9086);
or U11746 (N_11746,N_2060,N_8574);
xnor U11747 (N_11747,N_5530,N_1277);
and U11748 (N_11748,N_8573,N_6621);
nor U11749 (N_11749,N_6322,N_6272);
and U11750 (N_11750,N_9336,N_1409);
nor U11751 (N_11751,N_7910,N_7679);
and U11752 (N_11752,N_4538,N_8963);
nand U11753 (N_11753,N_7160,N_4895);
or U11754 (N_11754,N_152,N_9420);
and U11755 (N_11755,N_5574,N_2384);
or U11756 (N_11756,N_3488,N_5434);
nand U11757 (N_11757,N_1116,N_2432);
or U11758 (N_11758,N_1393,N_3827);
or U11759 (N_11759,N_5613,N_5135);
or U11760 (N_11760,N_5033,N_1904);
nor U11761 (N_11761,N_4610,N_3237);
nor U11762 (N_11762,N_577,N_9372);
or U11763 (N_11763,N_5303,N_4644);
nand U11764 (N_11764,N_2888,N_1674);
or U11765 (N_11765,N_1369,N_5898);
nor U11766 (N_11766,N_6630,N_7992);
nand U11767 (N_11767,N_6403,N_1943);
nand U11768 (N_11768,N_366,N_3156);
xnor U11769 (N_11769,N_7239,N_7606);
xor U11770 (N_11770,N_7726,N_1260);
and U11771 (N_11771,N_7453,N_2273);
nand U11772 (N_11772,N_2682,N_4195);
or U11773 (N_11773,N_9962,N_2776);
xnor U11774 (N_11774,N_2807,N_1098);
nor U11775 (N_11775,N_4555,N_9320);
nand U11776 (N_11776,N_3806,N_2670);
and U11777 (N_11777,N_9234,N_3836);
and U11778 (N_11778,N_6858,N_2468);
nor U11779 (N_11779,N_3032,N_5309);
nor U11780 (N_11780,N_9837,N_5988);
nand U11781 (N_11781,N_4627,N_1153);
nor U11782 (N_11782,N_1383,N_6053);
or U11783 (N_11783,N_8035,N_8745);
or U11784 (N_11784,N_3459,N_1117);
nor U11785 (N_11785,N_8593,N_7744);
nand U11786 (N_11786,N_9756,N_812);
xnor U11787 (N_11787,N_877,N_3518);
or U11788 (N_11788,N_8296,N_8278);
and U11789 (N_11789,N_995,N_5393);
nor U11790 (N_11790,N_2904,N_1831);
nand U11791 (N_11791,N_5510,N_5650);
and U11792 (N_11792,N_3804,N_4169);
xor U11793 (N_11793,N_6255,N_5736);
nor U11794 (N_11794,N_5138,N_5167);
xnor U11795 (N_11795,N_6697,N_9539);
nor U11796 (N_11796,N_4716,N_7959);
nor U11797 (N_11797,N_380,N_7323);
xor U11798 (N_11798,N_528,N_9556);
or U11799 (N_11799,N_6240,N_2170);
or U11800 (N_11800,N_3823,N_4449);
or U11801 (N_11801,N_4827,N_1719);
or U11802 (N_11802,N_3828,N_3555);
nand U11803 (N_11803,N_673,N_6508);
xnor U11804 (N_11804,N_8061,N_2968);
nor U11805 (N_11805,N_3294,N_6593);
or U11806 (N_11806,N_3197,N_2297);
nor U11807 (N_11807,N_6489,N_7354);
nand U11808 (N_11808,N_8257,N_1713);
or U11809 (N_11809,N_5127,N_1799);
and U11810 (N_11810,N_1314,N_4460);
xor U11811 (N_11811,N_5708,N_4803);
and U11812 (N_11812,N_8749,N_2301);
or U11813 (N_11813,N_8256,N_608);
nor U11814 (N_11814,N_4046,N_7740);
xnor U11815 (N_11815,N_6554,N_5790);
xnor U11816 (N_11816,N_9486,N_3627);
and U11817 (N_11817,N_6712,N_3309);
nor U11818 (N_11818,N_886,N_9613);
nand U11819 (N_11819,N_7830,N_7609);
nand U11820 (N_11820,N_3136,N_3299);
and U11821 (N_11821,N_7702,N_9393);
or U11822 (N_11822,N_6936,N_8267);
nor U11823 (N_11823,N_6498,N_7882);
and U11824 (N_11824,N_1984,N_1220);
nand U11825 (N_11825,N_9126,N_6155);
or U11826 (N_11826,N_7813,N_6428);
or U11827 (N_11827,N_2420,N_9004);
nand U11828 (N_11828,N_9178,N_7647);
or U11829 (N_11829,N_2326,N_6549);
and U11830 (N_11830,N_2806,N_2522);
and U11831 (N_11831,N_4161,N_9274);
or U11832 (N_11832,N_5889,N_3926);
and U11833 (N_11833,N_594,N_5306);
or U11834 (N_11834,N_3554,N_5308);
nor U11835 (N_11835,N_8383,N_9401);
nor U11836 (N_11836,N_4230,N_5689);
or U11837 (N_11837,N_9228,N_7231);
and U11838 (N_11838,N_1391,N_5751);
or U11839 (N_11839,N_5239,N_605);
and U11840 (N_11840,N_1399,N_1043);
and U11841 (N_11841,N_9379,N_9907);
nand U11842 (N_11842,N_7273,N_1138);
nand U11843 (N_11843,N_3092,N_2283);
nor U11844 (N_11844,N_5629,N_5717);
and U11845 (N_11845,N_2855,N_766);
and U11846 (N_11846,N_2571,N_258);
and U11847 (N_11847,N_5043,N_7324);
nand U11848 (N_11848,N_7745,N_1142);
nand U11849 (N_11849,N_409,N_8910);
nor U11850 (N_11850,N_2512,N_5265);
nor U11851 (N_11851,N_5588,N_9597);
or U11852 (N_11852,N_461,N_6220);
nand U11853 (N_11853,N_965,N_4453);
nor U11854 (N_11854,N_2271,N_8501);
nor U11855 (N_11855,N_2064,N_1560);
and U11856 (N_11856,N_6979,N_8539);
or U11857 (N_11857,N_4045,N_8004);
and U11858 (N_11858,N_7262,N_3660);
or U11859 (N_11859,N_1041,N_4860);
nand U11860 (N_11860,N_3039,N_5409);
nand U11861 (N_11861,N_3732,N_6048);
or U11862 (N_11862,N_8486,N_5532);
nand U11863 (N_11863,N_5450,N_7332);
or U11864 (N_11864,N_3218,N_7634);
nor U11865 (N_11865,N_5672,N_670);
and U11866 (N_11866,N_1547,N_8779);
or U11867 (N_11867,N_8034,N_9156);
nor U11868 (N_11868,N_4817,N_1434);
and U11869 (N_11869,N_5019,N_8214);
and U11870 (N_11870,N_998,N_8277);
nand U11871 (N_11871,N_7492,N_9219);
nor U11872 (N_11872,N_7379,N_4698);
nor U11873 (N_11873,N_6610,N_8399);
nor U11874 (N_11874,N_9611,N_4766);
xnor U11875 (N_11875,N_9419,N_261);
and U11876 (N_11876,N_8602,N_8066);
nor U11877 (N_11877,N_57,N_7874);
and U11878 (N_11878,N_4235,N_4788);
nand U11879 (N_11879,N_6972,N_647);
nand U11880 (N_11880,N_4585,N_6755);
nor U11881 (N_11881,N_2836,N_6455);
and U11882 (N_11882,N_467,N_6591);
nand U11883 (N_11883,N_9326,N_3433);
or U11884 (N_11884,N_6707,N_2825);
and U11885 (N_11885,N_2787,N_8414);
nor U11886 (N_11886,N_7434,N_1503);
or U11887 (N_11887,N_8459,N_5631);
xnor U11888 (N_11888,N_9757,N_8984);
nand U11889 (N_11889,N_944,N_8309);
nand U11890 (N_11890,N_9229,N_1934);
and U11891 (N_11891,N_3213,N_9725);
nand U11892 (N_11892,N_6842,N_7387);
nand U11893 (N_11893,N_3114,N_7760);
nor U11894 (N_11894,N_7659,N_7814);
and U11895 (N_11895,N_2686,N_9077);
nand U11896 (N_11896,N_870,N_2446);
nand U11897 (N_11897,N_4068,N_4800);
and U11898 (N_11898,N_2055,N_1851);
and U11899 (N_11899,N_9842,N_9776);
nand U11900 (N_11900,N_550,N_2144);
nand U11901 (N_11901,N_52,N_1921);
or U11902 (N_11902,N_50,N_923);
nor U11903 (N_11903,N_1819,N_121);
nor U11904 (N_11904,N_2658,N_4274);
nor U11905 (N_11905,N_7212,N_1415);
nand U11906 (N_11906,N_4059,N_9977);
or U11907 (N_11907,N_8512,N_1343);
and U11908 (N_11908,N_1319,N_3536);
and U11909 (N_11909,N_7381,N_8769);
xor U11910 (N_11910,N_6413,N_817);
nor U11911 (N_11911,N_7246,N_4016);
or U11912 (N_11912,N_2808,N_7489);
nor U11913 (N_11913,N_2300,N_4985);
or U11914 (N_11914,N_9332,N_6031);
or U11915 (N_11915,N_79,N_8678);
or U11916 (N_11916,N_9084,N_2119);
nand U11917 (N_11917,N_8146,N_9030);
xnor U11918 (N_11918,N_6198,N_2552);
nor U11919 (N_11919,N_2529,N_1445);
and U11920 (N_11920,N_1847,N_2767);
and U11921 (N_11921,N_4553,N_7875);
nor U11922 (N_11922,N_5090,N_3645);
nor U11923 (N_11923,N_1989,N_7883);
nand U11924 (N_11924,N_9082,N_9083);
nor U11925 (N_11925,N_4885,N_134);
xor U11926 (N_11926,N_4139,N_1199);
or U11927 (N_11927,N_1456,N_4035);
or U11928 (N_11928,N_4373,N_5969);
nor U11929 (N_11929,N_8368,N_5866);
and U11930 (N_11930,N_3795,N_1606);
xnor U11931 (N_11931,N_3330,N_9573);
xnor U11932 (N_11932,N_9035,N_7731);
or U11933 (N_11933,N_6966,N_5655);
or U11934 (N_11934,N_8655,N_4749);
or U11935 (N_11935,N_4419,N_7089);
nand U11936 (N_11936,N_259,N_4185);
or U11937 (N_11937,N_8804,N_2495);
xor U11938 (N_11938,N_5529,N_5175);
and U11939 (N_11939,N_3578,N_8968);
or U11940 (N_11940,N_3053,N_3719);
or U11941 (N_11941,N_2648,N_204);
nand U11942 (N_11942,N_7824,N_7826);
nand U11943 (N_11943,N_8452,N_6512);
xnor U11944 (N_11944,N_4693,N_1502);
and U11945 (N_11945,N_240,N_7015);
or U11946 (N_11946,N_7370,N_1573);
and U11947 (N_11947,N_5479,N_1637);
and U11948 (N_11948,N_4784,N_2134);
and U11949 (N_11949,N_6667,N_7218);
or U11950 (N_11950,N_9805,N_3407);
nand U11951 (N_11951,N_4084,N_1966);
nand U11952 (N_11952,N_6807,N_8086);
nand U11953 (N_11953,N_3061,N_4768);
and U11954 (N_11954,N_5681,N_5632);
and U11955 (N_11955,N_4810,N_7635);
or U11956 (N_11956,N_3229,N_624);
xnor U11957 (N_11957,N_602,N_7185);
nand U11958 (N_11958,N_2131,N_968);
xor U11959 (N_11959,N_6492,N_5236);
nand U11960 (N_11960,N_7233,N_7165);
xor U11961 (N_11961,N_5744,N_6869);
or U11962 (N_11962,N_2689,N_2521);
xnor U11963 (N_11963,N_9324,N_2557);
nand U11964 (N_11964,N_8708,N_9568);
or U11965 (N_11965,N_3432,N_676);
or U11966 (N_11966,N_9758,N_4899);
nor U11967 (N_11967,N_148,N_2286);
xor U11968 (N_11968,N_6649,N_4622);
or U11969 (N_11969,N_8489,N_7984);
or U11970 (N_11970,N_1853,N_8048);
nor U11971 (N_11971,N_2417,N_3932);
or U11972 (N_11972,N_7530,N_9115);
and U11973 (N_11973,N_9676,N_6701);
and U11974 (N_11974,N_2660,N_2666);
nor U11975 (N_11975,N_8858,N_7939);
and U11976 (N_11976,N_3911,N_2037);
nand U11977 (N_11977,N_9133,N_9451);
and U11978 (N_11978,N_8264,N_1953);
or U11979 (N_11979,N_802,N_4598);
nand U11980 (N_11980,N_5011,N_4536);
or U11981 (N_11981,N_6400,N_8999);
nor U11982 (N_11982,N_4391,N_6234);
nand U11983 (N_11983,N_1323,N_648);
nor U11984 (N_11984,N_8031,N_4528);
nand U11985 (N_11985,N_6330,N_2986);
nor U11986 (N_11986,N_8499,N_1727);
nand U11987 (N_11987,N_3509,N_4065);
xnor U11988 (N_11988,N_5586,N_129);
nand U11989 (N_11989,N_8676,N_300);
and U11990 (N_11990,N_9770,N_7688);
and U11991 (N_11991,N_9509,N_6160);
nor U11992 (N_11992,N_9950,N_5012);
or U11993 (N_11993,N_7747,N_1523);
nand U11994 (N_11994,N_2766,N_6117);
nor U11995 (N_11995,N_2187,N_1937);
nor U11996 (N_11996,N_4531,N_6747);
and U11997 (N_11997,N_5923,N_9434);
and U11998 (N_11998,N_2553,N_8791);
nor U11999 (N_11999,N_5817,N_3897);
nor U12000 (N_12000,N_9471,N_2791);
or U12001 (N_12001,N_4684,N_5350);
or U12002 (N_12002,N_9483,N_4647);
or U12003 (N_12003,N_3463,N_2068);
and U12004 (N_12004,N_8547,N_5869);
and U12005 (N_12005,N_6439,N_8375);
nor U12006 (N_12006,N_4316,N_5705);
or U12007 (N_12007,N_8877,N_558);
or U12008 (N_12008,N_5775,N_7825);
nand U12009 (N_12009,N_2536,N_5278);
or U12010 (N_12010,N_3577,N_9642);
xor U12011 (N_12011,N_6634,N_5344);
xnor U12012 (N_12012,N_6854,N_6541);
nand U12013 (N_12013,N_7772,N_8445);
or U12014 (N_12014,N_1007,N_252);
or U12015 (N_12015,N_2234,N_2030);
nor U12016 (N_12016,N_4098,N_4282);
nor U12017 (N_12017,N_7610,N_7062);
or U12018 (N_12018,N_2800,N_7803);
nor U12019 (N_12019,N_8393,N_5359);
xor U12020 (N_12020,N_7075,N_7620);
or U12021 (N_12021,N_9257,N_6106);
xor U12022 (N_12022,N_7925,N_5927);
nor U12023 (N_12023,N_9116,N_7948);
or U12024 (N_12024,N_7682,N_4815);
or U12025 (N_12025,N_2058,N_1173);
nand U12026 (N_12026,N_406,N_9016);
or U12027 (N_12027,N_9879,N_9346);
nand U12028 (N_12028,N_8429,N_7789);
nor U12029 (N_12029,N_4167,N_6030);
or U12030 (N_12030,N_1600,N_9694);
nand U12031 (N_12031,N_7035,N_5874);
nor U12032 (N_12032,N_7468,N_9875);
nand U12033 (N_12033,N_1807,N_430);
or U12034 (N_12034,N_6416,N_6135);
or U12035 (N_12035,N_8985,N_3005);
xor U12036 (N_12036,N_6727,N_9555);
nor U12037 (N_12037,N_1241,N_7341);
nor U12038 (N_12038,N_257,N_9679);
nor U12039 (N_12039,N_5237,N_2176);
and U12040 (N_12040,N_1459,N_5958);
nor U12041 (N_12041,N_7692,N_9021);
and U12042 (N_12042,N_7197,N_879);
or U12043 (N_12043,N_1225,N_3099);
or U12044 (N_12044,N_1813,N_7873);
nor U12045 (N_12045,N_4214,N_6908);
nor U12046 (N_12046,N_4087,N_4635);
nor U12047 (N_12047,N_8600,N_3313);
nand U12048 (N_12048,N_8253,N_6876);
nor U12049 (N_12049,N_6509,N_9474);
and U12050 (N_12050,N_5000,N_5168);
nor U12051 (N_12051,N_1780,N_2082);
nor U12052 (N_12052,N_1840,N_5156);
nor U12053 (N_12053,N_1233,N_7244);
xor U12054 (N_12054,N_5980,N_913);
or U12055 (N_12055,N_5638,N_4480);
nand U12056 (N_12056,N_4064,N_4676);
and U12057 (N_12057,N_6052,N_5369);
xor U12058 (N_12058,N_4208,N_4156);
nor U12059 (N_12059,N_4509,N_7287);
or U12060 (N_12060,N_4901,N_4296);
nand U12061 (N_12061,N_5916,N_8541);
nand U12062 (N_12062,N_9410,N_9991);
nor U12063 (N_12063,N_8950,N_3307);
nand U12064 (N_12064,N_9777,N_7847);
nor U12065 (N_12065,N_8391,N_5429);
and U12066 (N_12066,N_8358,N_3691);
or U12067 (N_12067,N_8571,N_1190);
xnor U12068 (N_12068,N_603,N_7898);
nand U12069 (N_12069,N_7912,N_7121);
or U12070 (N_12070,N_4215,N_789);
nand U12071 (N_12071,N_8663,N_9615);
nor U12072 (N_12072,N_525,N_8851);
nand U12073 (N_12073,N_6138,N_7592);
nand U12074 (N_12074,N_8422,N_2256);
nand U12075 (N_12075,N_2113,N_139);
nand U12076 (N_12076,N_4294,N_1696);
and U12077 (N_12077,N_671,N_5126);
xor U12078 (N_12078,N_1926,N_96);
nor U12079 (N_12079,N_7664,N_3141);
nor U12080 (N_12080,N_735,N_5767);
or U12081 (N_12081,N_3132,N_2063);
nor U12082 (N_12082,N_344,N_3482);
nand U12083 (N_12083,N_9333,N_606);
and U12084 (N_12084,N_1605,N_8618);
nor U12085 (N_12085,N_8711,N_8304);
or U12086 (N_12086,N_4671,N_6193);
nor U12087 (N_12087,N_4071,N_1626);
nand U12088 (N_12088,N_1958,N_2294);
or U12089 (N_12089,N_9343,N_3951);
and U12090 (N_12090,N_8738,N_353);
and U12091 (N_12091,N_3050,N_5675);
and U12092 (N_12092,N_3963,N_9458);
or U12093 (N_12093,N_9265,N_7535);
and U12094 (N_12094,N_9997,N_7040);
and U12095 (N_12095,N_8142,N_2647);
and U12096 (N_12096,N_1698,N_6035);
nor U12097 (N_12097,N_3914,N_320);
or U12098 (N_12098,N_9632,N_3702);
nor U12099 (N_12099,N_5221,N_3246);
nand U12100 (N_12100,N_151,N_9684);
nor U12101 (N_12101,N_5547,N_9815);
or U12102 (N_12102,N_2331,N_8798);
nand U12103 (N_12103,N_1465,N_3746);
nand U12104 (N_12104,N_2568,N_2569);
nand U12105 (N_12105,N_5815,N_5894);
nand U12106 (N_12106,N_3446,N_4668);
and U12107 (N_12107,N_2544,N_6872);
and U12108 (N_12108,N_9351,N_1478);
nor U12109 (N_12109,N_4483,N_2866);
nand U12110 (N_12110,N_8908,N_4106);
or U12111 (N_12111,N_8661,N_6693);
nand U12112 (N_12112,N_2245,N_722);
xor U12113 (N_12113,N_5472,N_786);
xor U12114 (N_12114,N_654,N_583);
or U12115 (N_12115,N_5870,N_2531);
or U12116 (N_12116,N_196,N_7460);
or U12117 (N_12117,N_4369,N_7926);
and U12118 (N_12118,N_1881,N_4936);
and U12119 (N_12119,N_4539,N_4516);
nor U12120 (N_12120,N_7039,N_5526);
and U12121 (N_12121,N_7960,N_5799);
nor U12122 (N_12122,N_6961,N_72);
nor U12123 (N_12123,N_8697,N_499);
or U12124 (N_12124,N_5419,N_256);
or U12125 (N_12125,N_6775,N_7714);
nand U12126 (N_12126,N_5478,N_5052);
nor U12127 (N_12127,N_3712,N_8055);
and U12128 (N_12128,N_5259,N_3203);
and U12129 (N_12129,N_4637,N_2282);
and U12130 (N_12130,N_4900,N_3259);
xnor U12131 (N_12131,N_282,N_3846);
xnor U12132 (N_12132,N_1157,N_7695);
nor U12133 (N_12133,N_2067,N_2249);
xor U12134 (N_12134,N_1230,N_78);
and U12135 (N_12135,N_5040,N_2465);
and U12136 (N_12136,N_484,N_8844);
nand U12137 (N_12137,N_1125,N_9250);
nand U12138 (N_12138,N_5010,N_1051);
or U12139 (N_12139,N_554,N_8052);
or U12140 (N_12140,N_1355,N_681);
and U12141 (N_12141,N_6963,N_7593);
xnor U12142 (N_12142,N_4688,N_1512);
nor U12143 (N_12143,N_9090,N_1655);
nor U12144 (N_12144,N_4153,N_3445);
and U12145 (N_12145,N_7756,N_5053);
or U12146 (N_12146,N_9664,N_8679);
and U12147 (N_12147,N_9783,N_5820);
and U12148 (N_12148,N_7601,N_9809);
or U12149 (N_12149,N_200,N_9161);
xor U12150 (N_12150,N_9139,N_7551);
and U12151 (N_12151,N_283,N_2621);
or U12152 (N_12152,N_4889,N_8020);
nor U12153 (N_12153,N_3643,N_6367);
nor U12154 (N_12154,N_6731,N_9709);
or U12155 (N_12155,N_1255,N_5081);
and U12156 (N_12156,N_7904,N_8412);
xor U12157 (N_12157,N_4947,N_4213);
nand U12158 (N_12158,N_2401,N_9557);
nor U12159 (N_12159,N_2260,N_8092);
and U12160 (N_12160,N_5197,N_1729);
and U12161 (N_12161,N_8709,N_4491);
nor U12162 (N_12162,N_6982,N_6536);
nor U12163 (N_12163,N_5037,N_1601);
and U12164 (N_12164,N_3162,N_2839);
nor U12165 (N_12165,N_8073,N_6572);
and U12166 (N_12166,N_653,N_763);
nand U12167 (N_12167,N_559,N_5291);
or U12168 (N_12168,N_3699,N_2411);
or U12169 (N_12169,N_2357,N_576);
nor U12170 (N_12170,N_2455,N_8758);
nand U12171 (N_12171,N_2015,N_4240);
and U12172 (N_12172,N_4149,N_1690);
and U12173 (N_12173,N_1646,N_9599);
nand U12174 (N_12174,N_2489,N_2985);
xnor U12175 (N_12175,N_7557,N_5075);
nand U12176 (N_12176,N_6456,N_2614);
and U12177 (N_12177,N_2699,N_7131);
nor U12178 (N_12178,N_9668,N_3634);
or U12179 (N_12179,N_6432,N_1345);
nor U12180 (N_12180,N_3952,N_3839);
nand U12181 (N_12181,N_9318,N_6708);
or U12182 (N_12182,N_9785,N_9859);
or U12183 (N_12183,N_8196,N_4232);
nand U12184 (N_12184,N_5544,N_6389);
nor U12185 (N_12185,N_4331,N_3849);
nor U12186 (N_12186,N_9088,N_7776);
nand U12187 (N_12187,N_8390,N_4819);
or U12188 (N_12188,N_2043,N_9293);
nor U12189 (N_12189,N_7853,N_4729);
xnor U12190 (N_12190,N_6750,N_7104);
or U12191 (N_12191,N_5568,N_1438);
nor U12192 (N_12192,N_1356,N_7952);
and U12193 (N_12193,N_9501,N_462);
or U12194 (N_12194,N_1917,N_6244);
or U12195 (N_12195,N_248,N_828);
nor U12196 (N_12196,N_5968,N_9197);
nand U12197 (N_12197,N_7427,N_5069);
or U12198 (N_12198,N_3780,N_4846);
and U12199 (N_12199,N_1289,N_9431);
nand U12200 (N_12200,N_2314,N_3409);
or U12201 (N_12201,N_9047,N_1272);
or U12202 (N_12202,N_4514,N_7365);
or U12203 (N_12203,N_3903,N_9003);
or U12204 (N_12204,N_4089,N_1770);
and U12205 (N_12205,N_7135,N_6897);
nand U12206 (N_12206,N_4737,N_3065);
nand U12207 (N_12207,N_7019,N_6531);
nor U12208 (N_12208,N_1671,N_3543);
nand U12209 (N_12209,N_9110,N_7119);
or U12210 (N_12210,N_2761,N_5465);
or U12211 (N_12211,N_6100,N_2922);
xor U12212 (N_12212,N_8933,N_4523);
nor U12213 (N_12213,N_2706,N_4248);
or U12214 (N_12214,N_2723,N_1625);
nand U12215 (N_12215,N_8787,N_5590);
or U12216 (N_12216,N_1219,N_5805);
nand U12217 (N_12217,N_2817,N_6636);
nor U12218 (N_12218,N_6709,N_8978);
and U12219 (N_12219,N_5953,N_9487);
and U12220 (N_12220,N_1126,N_7708);
nor U12221 (N_12221,N_6307,N_7164);
or U12222 (N_12222,N_2038,N_347);
or U12223 (N_12223,N_7894,N_4020);
or U12224 (N_12224,N_4382,N_2961);
nand U12225 (N_12225,N_4876,N_684);
or U12226 (N_12226,N_6274,N_3935);
and U12227 (N_12227,N_1568,N_9774);
nor U12228 (N_12228,N_3479,N_8111);
and U12229 (N_12229,N_6219,N_3460);
or U12230 (N_12230,N_1328,N_2213);
xor U12231 (N_12231,N_4461,N_9425);
or U12232 (N_12232,N_1148,N_9923);
and U12233 (N_12233,N_7093,N_9452);
or U12234 (N_12234,N_5892,N_1919);
xor U12235 (N_12235,N_969,N_4287);
nand U12236 (N_12236,N_9493,N_6949);
and U12237 (N_12237,N_5784,N_5563);
nand U12238 (N_12238,N_1044,N_771);
nor U12239 (N_12239,N_6128,N_9412);
and U12240 (N_12240,N_9570,N_4018);
nor U12241 (N_12241,N_7376,N_2230);
nand U12242 (N_12242,N_5224,N_5375);
or U12243 (N_12243,N_2889,N_6603);
nor U12244 (N_12244,N_3186,N_4173);
nor U12245 (N_12245,N_549,N_8786);
or U12246 (N_12246,N_4625,N_1296);
and U12247 (N_12247,N_7919,N_2151);
nor U12248 (N_12248,N_1155,N_8562);
nand U12249 (N_12249,N_1270,N_4142);
and U12250 (N_12250,N_7633,N_159);
nand U12251 (N_12251,N_7891,N_8149);
and U12252 (N_12252,N_3334,N_1809);
and U12253 (N_12253,N_9961,N_2926);
or U12254 (N_12254,N_5974,N_7377);
xnor U12255 (N_12255,N_1318,N_6505);
nor U12256 (N_12256,N_45,N_27);
nand U12257 (N_12257,N_7739,N_8320);
and U12258 (N_12258,N_7174,N_6401);
or U12259 (N_12259,N_1059,N_6152);
nand U12260 (N_12260,N_9345,N_207);
or U12261 (N_12261,N_8134,N_3390);
nand U12262 (N_12262,N_8821,N_3284);
and U12263 (N_12263,N_8720,N_8294);
xor U12264 (N_12264,N_1107,N_2012);
nand U12265 (N_12265,N_4512,N_4399);
nor U12266 (N_12266,N_1439,N_9369);
nand U12267 (N_12267,N_9607,N_862);
nand U12268 (N_12268,N_3841,N_8912);
xor U12269 (N_12269,N_1192,N_669);
nor U12270 (N_12270,N_8463,N_5179);
nor U12271 (N_12271,N_378,N_9578);
nand U12272 (N_12272,N_1844,N_2972);
and U12273 (N_12273,N_5056,N_245);
and U12274 (N_12274,N_872,N_992);
xnor U12275 (N_12275,N_4724,N_544);
nand U12276 (N_12276,N_8982,N_8731);
or U12277 (N_12277,N_2997,N_5322);
nand U12278 (N_12278,N_2279,N_9097);
nand U12279 (N_12279,N_6958,N_2333);
nand U12280 (N_12280,N_5509,N_8727);
nor U12281 (N_12281,N_3704,N_8892);
nor U12282 (N_12282,N_7230,N_3115);
or U12283 (N_12283,N_707,N_535);
xor U12284 (N_12284,N_6893,N_9353);
or U12285 (N_12285,N_3122,N_5731);
or U12286 (N_12286,N_458,N_7346);
xnor U12287 (N_12287,N_2626,N_5771);
or U12288 (N_12288,N_469,N_7284);
or U12289 (N_12289,N_306,N_4614);
or U12290 (N_12290,N_2630,N_2543);
nand U12291 (N_12291,N_8521,N_1593);
or U12292 (N_12292,N_4385,N_2623);
nor U12293 (N_12293,N_5776,N_3058);
nand U12294 (N_12294,N_1273,N_1291);
nand U12295 (N_12295,N_4727,N_2359);
xnor U12296 (N_12296,N_4432,N_6986);
and U12297 (N_12297,N_9454,N_2583);
xnor U12298 (N_12298,N_482,N_9391);
xnor U12299 (N_12299,N_9554,N_6217);
xnor U12300 (N_12300,N_5770,N_9657);
nand U12301 (N_12301,N_9826,N_2909);
and U12302 (N_12302,N_8421,N_9490);
and U12303 (N_12303,N_1484,N_7005);
nor U12304 (N_12304,N_21,N_1358);
nand U12305 (N_12305,N_4620,N_3608);
nand U12306 (N_12306,N_7388,N_8525);
nand U12307 (N_12307,N_8513,N_9269);
or U12308 (N_12308,N_1848,N_9008);
nand U12309 (N_12309,N_6176,N_2948);
nand U12310 (N_12310,N_8096,N_8386);
and U12311 (N_12311,N_7996,N_7685);
and U12312 (N_12312,N_6921,N_4049);
xnor U12313 (N_12313,N_4298,N_1472);
nor U12314 (N_12314,N_3332,N_574);
and U12315 (N_12315,N_9973,N_81);
nand U12316 (N_12316,N_1061,N_686);
or U12317 (N_12317,N_571,N_2490);
nand U12318 (N_12318,N_2524,N_6599);
or U12319 (N_12319,N_4582,N_3344);
or U12320 (N_12320,N_3049,N_9900);
and U12321 (N_12321,N_7209,N_8596);
nor U12322 (N_12322,N_632,N_659);
or U12323 (N_12323,N_3254,N_6892);
nor U12324 (N_12324,N_4448,N_8203);
nor U12325 (N_12325,N_5364,N_4808);
and U12326 (N_12326,N_794,N_3749);
nor U12327 (N_12327,N_2185,N_86);
or U12328 (N_12328,N_7493,N_5581);
nor U12329 (N_12329,N_2674,N_2516);
or U12330 (N_12330,N_839,N_1896);
or U12331 (N_12331,N_417,N_4518);
nor U12332 (N_12332,N_1333,N_568);
or U12333 (N_12333,N_1286,N_696);
or U12334 (N_12334,N_2116,N_1245);
and U12335 (N_12335,N_8054,N_8490);
and U12336 (N_12336,N_7507,N_5779);
xnor U12337 (N_12337,N_1546,N_9298);
nor U12338 (N_12338,N_5399,N_7430);
xnor U12339 (N_12339,N_3308,N_8930);
and U12340 (N_12340,N_1868,N_3083);
and U12341 (N_12341,N_8344,N_7958);
and U12342 (N_12342,N_7913,N_7544);
and U12343 (N_12343,N_8662,N_4288);
nor U12344 (N_12344,N_9847,N_7488);
nor U12345 (N_12345,N_2784,N_5691);
or U12346 (N_12346,N_1590,N_4387);
nand U12347 (N_12347,N_8036,N_636);
nor U12348 (N_12348,N_1058,N_5841);
nor U12349 (N_12349,N_8397,N_6302);
or U12350 (N_12350,N_4675,N_3248);
and U12351 (N_12351,N_6405,N_8611);
or U12352 (N_12352,N_7120,N_8190);
nand U12353 (N_12353,N_2003,N_3685);
xor U12354 (N_12354,N_2949,N_937);
or U12355 (N_12355,N_2896,N_9268);
or U12356 (N_12356,N_5956,N_4354);
or U12357 (N_12357,N_7258,N_1878);
nand U12358 (N_12358,N_7330,N_8819);
nand U12359 (N_12359,N_4859,N_9157);
nor U12360 (N_12360,N_7214,N_596);
nor U12361 (N_12361,N_9303,N_3802);
nor U12362 (N_12362,N_7144,N_7727);
xor U12363 (N_12363,N_1668,N_9512);
nor U12364 (N_12364,N_2125,N_3614);
xnor U12365 (N_12365,N_3430,N_1923);
and U12366 (N_12366,N_4,N_3787);
or U12367 (N_12367,N_7643,N_8699);
and U12368 (N_12368,N_3373,N_7129);
and U12369 (N_12369,N_7423,N_3422);
and U12370 (N_12370,N_9943,N_6951);
and U12371 (N_12371,N_9091,N_6698);
nand U12372 (N_12372,N_6038,N_9505);
nor U12373 (N_12373,N_1159,N_5729);
and U12374 (N_12374,N_1642,N_6791);
and U12375 (N_12375,N_7208,N_1046);
nor U12376 (N_12376,N_6552,N_8934);
nand U12377 (N_12377,N_2770,N_1017);
nand U12378 (N_12378,N_1530,N_113);
nand U12379 (N_12379,N_6802,N_3669);
nor U12380 (N_12380,N_4513,N_7561);
nand U12381 (N_12381,N_5934,N_991);
nor U12382 (N_12382,N_9646,N_6120);
and U12383 (N_12383,N_2302,N_7369);
nor U12384 (N_12384,N_2960,N_2229);
nor U12385 (N_12385,N_5545,N_8295);
nand U12386 (N_12386,N_6665,N_6540);
nor U12387 (N_12387,N_9366,N_4492);
nor U12388 (N_12388,N_5045,N_9316);
and U12389 (N_12389,N_7018,N_6039);
xnor U12390 (N_12390,N_9856,N_3982);
and U12391 (N_12391,N_7852,N_5288);
or U12392 (N_12392,N_3987,N_4583);
and U12393 (N_12393,N_4587,N_5493);
and U12394 (N_12394,N_5652,N_2164);
nor U12395 (N_12395,N_1551,N_91);
xor U12396 (N_12396,N_9437,N_1888);
nand U12397 (N_12397,N_3279,N_6662);
nor U12398 (N_12398,N_9645,N_2528);
xnor U12399 (N_12399,N_3220,N_438);
and U12400 (N_12400,N_6034,N_6624);
and U12401 (N_12401,N_9339,N_5332);
or U12402 (N_12402,N_1316,N_8381);
nand U12403 (N_12403,N_2337,N_1839);
xnor U12404 (N_12404,N_4822,N_6780);
and U12405 (N_12405,N_335,N_6534);
nor U12406 (N_12406,N_3747,N_7210);
or U12407 (N_12407,N_7612,N_8094);
and U12408 (N_12408,N_678,N_736);
or U12409 (N_12409,N_9044,N_5783);
xor U12410 (N_12410,N_1084,N_9914);
or U12411 (N_12411,N_1422,N_9051);
or U12412 (N_12412,N_8299,N_9005);
and U12413 (N_12413,N_6199,N_9731);
nand U12414 (N_12414,N_7977,N_5612);
nor U12415 (N_12415,N_7173,N_8905);
or U12416 (N_12416,N_6933,N_8342);
nand U12417 (N_12417,N_3644,N_5860);
or U12418 (N_12418,N_7179,N_1092);
nor U12419 (N_12419,N_3177,N_2743);
and U12420 (N_12420,N_8122,N_2291);
and U12421 (N_12421,N_7359,N_194);
and U12422 (N_12422,N_5696,N_4677);
and U12423 (N_12423,N_4836,N_128);
or U12424 (N_12424,N_9929,N_769);
nand U12425 (N_12425,N_6449,N_4442);
nor U12426 (N_12426,N_1284,N_2838);
or U12427 (N_12427,N_4562,N_2779);
xnor U12428 (N_12428,N_4849,N_4269);
nand U12429 (N_12429,N_4972,N_1266);
nand U12430 (N_12430,N_7531,N_9149);
nor U12431 (N_12431,N_6084,N_3611);
nor U12432 (N_12432,N_9854,N_5521);
nor U12433 (N_12433,N_9253,N_7585);
nand U12434 (N_12434,N_464,N_3107);
and U12435 (N_12435,N_7260,N_8051);
or U12436 (N_12436,N_2143,N_4138);
nor U12437 (N_12437,N_1052,N_2772);
nor U12438 (N_12438,N_7006,N_3301);
nand U12439 (N_12439,N_9988,N_5353);
and U12440 (N_12440,N_3204,N_8310);
xnor U12441 (N_12441,N_122,N_2443);
xnor U12442 (N_12442,N_3742,N_5961);
nor U12443 (N_12443,N_1209,N_203);
xnor U12444 (N_12444,N_5082,N_322);
xor U12445 (N_12445,N_4191,N_2707);
nor U12446 (N_12446,N_8605,N_3012);
or U12447 (N_12447,N_520,N_6847);
and U12448 (N_12448,N_2730,N_4792);
nor U12449 (N_12449,N_2719,N_1500);
and U12450 (N_12450,N_6564,N_3979);
nor U12451 (N_12451,N_2092,N_7676);
or U12452 (N_12452,N_5446,N_9315);
or U12453 (N_12453,N_565,N_7417);
nor U12454 (N_12454,N_753,N_3075);
nand U12455 (N_12455,N_1746,N_7213);
or U12456 (N_12456,N_4550,N_8183);
xnor U12457 (N_12457,N_4123,N_5038);
or U12458 (N_12458,N_4041,N_4281);
or U12459 (N_12459,N_7169,N_6976);
nand U12460 (N_12460,N_2013,N_8651);
nor U12461 (N_12461,N_1508,N_5828);
nor U12462 (N_12462,N_5060,N_8995);
and U12463 (N_12463,N_841,N_6337);
and U12464 (N_12464,N_1942,N_685);
nor U12465 (N_12465,N_6888,N_9655);
or U12466 (N_12466,N_6469,N_7274);
nand U12467 (N_12467,N_641,N_1181);
or U12468 (N_12468,N_38,N_8939);
nor U12469 (N_12469,N_3965,N_6105);
xnor U12470 (N_12470,N_816,N_572);
and U12471 (N_12471,N_8783,N_1271);
nor U12472 (N_12472,N_7501,N_6289);
or U12473 (N_12473,N_4024,N_2963);
nor U12474 (N_12474,N_6765,N_8466);
and U12475 (N_12475,N_1969,N_1238);
and U12476 (N_12476,N_2332,N_7270);
nand U12477 (N_12477,N_107,N_5561);
nor U12478 (N_12478,N_893,N_8888);
and U12479 (N_12479,N_1053,N_4165);
or U12480 (N_12480,N_7944,N_144);
xnor U12481 (N_12481,N_6832,N_8918);
and U12482 (N_12482,N_1513,N_3584);
or U12483 (N_12483,N_3688,N_1879);
and U12484 (N_12484,N_860,N_8401);
and U12485 (N_12485,N_770,N_7753);
and U12486 (N_12486,N_7459,N_892);
nand U12487 (N_12487,N_3471,N_5601);
or U12488 (N_12488,N_1763,N_2439);
nor U12489 (N_12489,N_567,N_8209);
or U12490 (N_12490,N_4820,N_6912);
nor U12491 (N_12491,N_7361,N_3501);
nor U12492 (N_12492,N_6338,N_650);
nand U12493 (N_12493,N_9381,N_6974);
and U12494 (N_12494,N_237,N_6288);
or U12495 (N_12495,N_8957,N_8431);
and U12496 (N_12496,N_2393,N_4725);
nor U12497 (N_12497,N_9094,N_867);
and U12498 (N_12498,N_4154,N_5694);
nand U12499 (N_12499,N_868,N_5483);
or U12500 (N_12500,N_3215,N_2005);
nor U12501 (N_12501,N_5872,N_3127);
and U12502 (N_12502,N_7785,N_5390);
or U12503 (N_12503,N_5742,N_9868);
nand U12504 (N_12504,N_9125,N_4102);
nand U12505 (N_12505,N_29,N_5920);
and U12506 (N_12506,N_4358,N_9103);
nor U12507 (N_12507,N_2995,N_4012);
xnor U12508 (N_12508,N_8584,N_9819);
or U12509 (N_12509,N_4498,N_6436);
nor U12510 (N_12510,N_4608,N_8815);
or U12511 (N_12511,N_716,N_7451);
nand U12512 (N_12512,N_2768,N_7146);
xor U12513 (N_12513,N_4454,N_9949);
nand U12514 (N_12514,N_5781,N_2436);
or U12515 (N_12515,N_4261,N_7108);
nand U12516 (N_12516,N_6749,N_2680);
and U12517 (N_12517,N_1712,N_3399);
or U12518 (N_12518,N_8631,N_452);
nand U12519 (N_12519,N_6833,N_2009);
or U12520 (N_12520,N_2368,N_2716);
nor U12521 (N_12521,N_4307,N_174);
nor U12522 (N_12522,N_6864,N_2642);
and U12523 (N_12523,N_6447,N_3553);
nor U12524 (N_12524,N_2843,N_169);
and U12525 (N_12525,N_1684,N_889);
and U12526 (N_12526,N_9520,N_4458);
nor U12527 (N_12527,N_9762,N_8684);
nand U12528 (N_12528,N_7639,N_7312);
nand U12529 (N_12529,N_2293,N_9017);
or U12530 (N_12530,N_4126,N_734);
or U12531 (N_12531,N_1364,N_3880);
xor U12532 (N_12532,N_820,N_9446);
or U12533 (N_12533,N_7741,N_5663);
nor U12534 (N_12534,N_2605,N_6303);
and U12535 (N_12535,N_3534,N_856);
and U12536 (N_12536,N_8659,N_1453);
nor U12537 (N_12537,N_6788,N_3629);
and U12538 (N_12538,N_6574,N_6011);
nand U12539 (N_12539,N_1948,N_7318);
nor U12540 (N_12540,N_3227,N_5173);
or U12541 (N_12541,N_7793,N_2802);
or U12542 (N_12542,N_9426,N_8205);
nand U12543 (N_12543,N_2980,N_3320);
nand U12544 (N_12544,N_3976,N_1537);
or U12545 (N_12545,N_7527,N_2894);
and U12546 (N_12546,N_7509,N_7868);
nand U12547 (N_12547,N_7806,N_2515);
nand U12548 (N_12548,N_2691,N_7182);
or U12549 (N_12549,N_3398,N_4070);
or U12550 (N_12550,N_3244,N_9627);
nor U12551 (N_12551,N_8024,N_2083);
and U12552 (N_12552,N_957,N_9616);
nor U12553 (N_12553,N_6935,N_2200);
and U12554 (N_12554,N_6218,N_5863);
nor U12555 (N_12555,N_2212,N_4624);
and U12556 (N_12556,N_7862,N_6811);
and U12557 (N_12557,N_8204,N_9494);
and U12558 (N_12558,N_7802,N_3924);
nor U12559 (N_12559,N_1162,N_447);
nor U12560 (N_12560,N_9144,N_6916);
xor U12561 (N_12561,N_6223,N_2195);
xor U12562 (N_12562,N_2712,N_4062);
and U12563 (N_12563,N_114,N_4017);
xnor U12564 (N_12564,N_6058,N_2254);
nor U12565 (N_12565,N_1354,N_5068);
or U12566 (N_12566,N_2718,N_4931);
or U12567 (N_12567,N_9295,N_4309);
nor U12568 (N_12568,N_4007,N_2582);
xnor U12569 (N_12569,N_8090,N_3668);
or U12570 (N_12570,N_9808,N_7374);
nor U12571 (N_12571,N_7962,N_6629);
or U12572 (N_12572,N_3362,N_6799);
or U12573 (N_12573,N_428,N_4527);
or U12574 (N_12574,N_4648,N_8075);
nand U12575 (N_12575,N_7537,N_9849);
nand U12576 (N_12576,N_4520,N_561);
nor U12577 (N_12577,N_5942,N_4197);
and U12578 (N_12578,N_302,N_7402);
nand U12579 (N_12579,N_9484,N_9797);
and U12580 (N_12580,N_6365,N_4712);
nand U12581 (N_12581,N_5042,N_740);
and U12582 (N_12582,N_1353,N_3942);
nor U12583 (N_12583,N_6393,N_6746);
or U12584 (N_12584,N_2988,N_2482);
and U12585 (N_12585,N_8789,N_7547);
nor U12586 (N_12586,N_1308,N_7269);
or U12587 (N_12587,N_4305,N_6845);
and U12588 (N_12588,N_1961,N_8556);
nor U12589 (N_12589,N_7199,N_8121);
and U12590 (N_12590,N_9791,N_1340);
and U12591 (N_12591,N_5158,N_7194);
or U12592 (N_12592,N_9476,N_3355);
and U12593 (N_12593,N_9967,N_1981);
and U12594 (N_12594,N_7063,N_8377);
xnor U12595 (N_12595,N_8022,N_4979);
and U12596 (N_12596,N_4618,N_9166);
and U12597 (N_12597,N_9107,N_5608);
nand U12598 (N_12598,N_3520,N_9705);
or U12599 (N_12599,N_3064,N_5261);
nand U12600 (N_12600,N_1561,N_5164);
nand U12601 (N_12601,N_3606,N_8990);
nand U12602 (N_12602,N_7957,N_3223);
xor U12603 (N_12603,N_160,N_8935);
xor U12604 (N_12604,N_7321,N_2473);
or U12605 (N_12605,N_800,N_2129);
nor U12606 (N_12606,N_8686,N_2193);
nand U12607 (N_12607,N_1628,N_2577);
nand U12608 (N_12608,N_5738,N_7022);
nand U12609 (N_12609,N_6742,N_3287);
or U12610 (N_12610,N_4535,N_8953);
nor U12611 (N_12611,N_4107,N_9463);
nor U12612 (N_12612,N_7000,N_2441);
xor U12613 (N_12613,N_1370,N_1648);
xnor U12614 (N_12614,N_1338,N_5165);
xnor U12615 (N_12615,N_2852,N_7107);
nand U12616 (N_12616,N_493,N_5268);
nor U12617 (N_12617,N_6682,N_9102);
xnor U12618 (N_12618,N_8133,N_5982);
or U12619 (N_12619,N_9746,N_4377);
nand U12620 (N_12620,N_5971,N_6501);
nor U12621 (N_12621,N_8955,N_6556);
nor U12622 (N_12622,N_175,N_5495);
or U12623 (N_12623,N_4917,N_1191);
nand U12624 (N_12624,N_8991,N_1229);
and U12625 (N_12625,N_4008,N_2201);
nand U12626 (N_12626,N_5381,N_7017);
nor U12627 (N_12627,N_2913,N_2317);
nor U12628 (N_12628,N_8817,N_4265);
and U12629 (N_12629,N_429,N_5189);
nor U12630 (N_12630,N_1144,N_9183);
nor U12631 (N_12631,N_6865,N_3381);
and U12632 (N_12632,N_5664,N_904);
xnor U12633 (N_12633,N_7437,N_2549);
and U12634 (N_12634,N_6955,N_8026);
and U12635 (N_12635,N_1758,N_1945);
or U12636 (N_12636,N_3896,N_4431);
nand U12637 (N_12637,N_4829,N_1419);
nand U12638 (N_12638,N_1,N_895);
and U12639 (N_12639,N_9656,N_850);
nand U12640 (N_12640,N_4481,N_1863);
nand U12641 (N_12641,N_3163,N_3104);
xnor U12642 (N_12642,N_7462,N_4878);
or U12643 (N_12643,N_643,N_5838);
nand U12644 (N_12644,N_7163,N_6440);
nand U12645 (N_12645,N_2644,N_3441);
and U12646 (N_12646,N_4241,N_593);
and U12647 (N_12647,N_1407,N_4468);
nand U12648 (N_12648,N_2034,N_2324);
nand U12649 (N_12649,N_8826,N_4958);
nand U12650 (N_12650,N_3476,N_9745);
and U12651 (N_12651,N_364,N_7476);
and U12652 (N_12652,N_1755,N_5200);
nor U12653 (N_12653,N_8665,N_6023);
nor U12654 (N_12654,N_9001,N_9222);
or U12655 (N_12655,N_4348,N_2540);
or U12656 (N_12656,N_3128,N_2458);
and U12657 (N_12657,N_773,N_6226);
and U12658 (N_12658,N_4192,N_619);
nand U12659 (N_12659,N_1870,N_3519);
or U12660 (N_12660,N_2250,N_8182);
nor U12661 (N_12661,N_54,N_3158);
and U12662 (N_12662,N_6008,N_8130);
nand U12663 (N_12663,N_1708,N_9395);
or U12664 (N_12664,N_421,N_1906);
nand U12665 (N_12665,N_5728,N_9751);
nor U12666 (N_12666,N_4547,N_4759);
nand U12667 (N_12667,N_4234,N_2042);
xor U12668 (N_12668,N_5851,N_5118);
nor U12669 (N_12669,N_2762,N_1744);
or U12670 (N_12670,N_6227,N_9909);
nor U12671 (N_12671,N_4425,N_644);
or U12672 (N_12672,N_3256,N_2989);
or U12673 (N_12673,N_845,N_9453);
nand U12674 (N_12674,N_2567,N_4557);
xor U12675 (N_12675,N_4472,N_4973);
or U12676 (N_12676,N_5826,N_1254);
xnor U12677 (N_12677,N_4108,N_3670);
and U12678 (N_12678,N_1737,N_3185);
and U12679 (N_12679,N_2475,N_950);
or U12680 (N_12680,N_3414,N_5105);
xnor U12681 (N_12681,N_9155,N_7407);
or U12682 (N_12682,N_2320,N_7703);
nand U12683 (N_12683,N_1731,N_3893);
nor U12684 (N_12684,N_4920,N_9286);
and U12685 (N_12685,N_7012,N_6394);
xnor U12686 (N_12686,N_5921,N_9289);
and U12687 (N_12687,N_1976,N_6402);
or U12688 (N_12688,N_2138,N_7782);
and U12689 (N_12689,N_3700,N_8869);
nand U12690 (N_12690,N_2939,N_916);
xnor U12691 (N_12691,N_6607,N_8165);
nor U12692 (N_12692,N_3181,N_2347);
or U12693 (N_12693,N_1834,N_7573);
or U12694 (N_12694,N_6997,N_164);
or U12695 (N_12695,N_3420,N_8398);
nand U12696 (N_12696,N_2403,N_8498);
xnor U12697 (N_12697,N_2591,N_3296);
and U12698 (N_12698,N_6482,N_4341);
nor U12699 (N_12699,N_963,N_9804);
and U12700 (N_12700,N_5125,N_9803);
and U12701 (N_12701,N_2281,N_6871);
and U12702 (N_12702,N_9365,N_3916);
and U12703 (N_12703,N_9590,N_6786);
nor U12704 (N_12704,N_6734,N_2601);
xnor U12705 (N_12705,N_480,N_6141);
nand U12706 (N_12706,N_7936,N_2684);
nand U12707 (N_12707,N_3003,N_7748);
or U12708 (N_12708,N_5797,N_5948);
or U12709 (N_12709,N_8062,N_6909);
and U12710 (N_12710,N_2935,N_6996);
xor U12711 (N_12711,N_4943,N_6960);
xor U12712 (N_12712,N_2296,N_6060);
and U12713 (N_12713,N_5904,N_3397);
or U12714 (N_12714,N_3623,N_2181);
nand U12715 (N_12715,N_7786,N_3035);
nor U12716 (N_12716,N_6691,N_1239);
xor U12717 (N_12717,N_2280,N_9898);
xor U12718 (N_12718,N_4267,N_5468);
nand U12719 (N_12719,N_4867,N_4720);
and U12720 (N_12720,N_5349,N_3303);
or U12721 (N_12721,N_6615,N_1495);
or U12722 (N_12722,N_8384,N_7885);
and U12723 (N_12723,N_8016,N_7245);
or U12724 (N_12724,N_7928,N_6252);
nor U12725 (N_12725,N_5020,N_9224);
or U12726 (N_12726,N_8803,N_9200);
or U12727 (N_12727,N_3072,N_6451);
nand U12728 (N_12728,N_1841,N_7060);
nand U12729 (N_12729,N_358,N_9220);
nand U12730 (N_12730,N_5229,N_1527);
and U12731 (N_12731,N_7014,N_3324);
xor U12732 (N_12732,N_5913,N_2323);
or U12733 (N_12733,N_7220,N_1149);
nand U12734 (N_12734,N_55,N_1243);
nor U12735 (N_12735,N_333,N_7955);
nand U12736 (N_12736,N_7353,N_6521);
nor U12737 (N_12737,N_9592,N_8274);
and U12738 (N_12738,N_5400,N_621);
xor U12739 (N_12739,N_1196,N_1517);
and U12740 (N_12740,N_8742,N_4058);
or U12741 (N_12741,N_2413,N_8266);
nor U12742 (N_12742,N_1026,N_1347);
or U12743 (N_12743,N_5305,N_534);
nand U12744 (N_12744,N_7588,N_4393);
and U12745 (N_12745,N_4855,N_9930);
nor U12746 (N_12746,N_7556,N_292);
nand U12747 (N_12747,N_7675,N_1659);
and U12748 (N_12748,N_403,N_8629);
nor U12749 (N_12749,N_9699,N_229);
nand U12750 (N_12750,N_2463,N_7751);
or U12751 (N_12751,N_7092,N_7506);
and U12752 (N_12752,N_9755,N_3314);
and U12753 (N_12753,N_4360,N_4372);
nor U12754 (N_12754,N_7072,N_4200);
and U12755 (N_12755,N_2435,N_2127);
nor U12756 (N_12756,N_1141,N_5713);
and U12757 (N_12757,N_93,N_1263);
xor U12758 (N_12758,N_5908,N_8873);
or U12759 (N_12759,N_5830,N_9912);
nand U12760 (N_12760,N_6271,N_4019);
or U12761 (N_12761,N_2887,N_360);
nor U12762 (N_12762,N_1336,N_7650);
and U12763 (N_12763,N_6386,N_5903);
xnor U12764 (N_12764,N_7095,N_9551);
and U12765 (N_12765,N_8630,N_1944);
or U12766 (N_12766,N_6971,N_5321);
and U12767 (N_12767,N_4977,N_8349);
nand U12768 (N_12768,N_2223,N_8974);
or U12769 (N_12769,N_2652,N_664);
nor U12770 (N_12770,N_6118,N_4912);
and U12771 (N_12771,N_8911,N_6101);
nand U12772 (N_12772,N_25,N_6514);
nand U12773 (N_12773,N_6628,N_1718);
and U12774 (N_12774,N_24,N_9259);
or U12775 (N_12775,N_7280,N_8734);
xor U12776 (N_12776,N_1920,N_6069);
and U12777 (N_12777,N_9363,N_2755);
xnor U12778 (N_12778,N_5292,N_6458);
and U12779 (N_12779,N_3842,N_9972);
nor U12780 (N_12780,N_1009,N_1493);
nor U12781 (N_12781,N_1629,N_5706);
nand U12782 (N_12782,N_5798,N_6171);
nor U12783 (N_12783,N_2780,N_4401);
nand U12784 (N_12784,N_5566,N_9644);
and U12785 (N_12785,N_5810,N_3119);
and U12786 (N_12786,N_8227,N_4866);
or U12787 (N_12787,N_7196,N_8);
nor U12788 (N_12788,N_4963,N_6154);
nand U12789 (N_12789,N_1423,N_8301);
nor U12790 (N_12790,N_5996,N_9195);
nor U12791 (N_12791,N_9481,N_6308);
or U12792 (N_12792,N_4160,N_9317);
xnor U12793 (N_12793,N_9631,N_2819);
nor U12794 (N_12794,N_483,N_4129);
and U12795 (N_12795,N_1991,N_1632);
or U12796 (N_12796,N_2835,N_7661);
or U12797 (N_12797,N_7901,N_2751);
or U12798 (N_12798,N_6962,N_4029);
nor U12799 (N_12799,N_7515,N_7765);
nand U12800 (N_12800,N_3044,N_5304);
xor U12801 (N_12801,N_2239,N_1820);
and U12802 (N_12802,N_4704,N_8837);
nand U12803 (N_12803,N_8402,N_7301);
nand U12804 (N_12804,N_7181,N_8405);
nand U12805 (N_12805,N_8451,N_6525);
nand U12806 (N_12806,N_7595,N_8747);
or U12807 (N_12807,N_4380,N_9998);
nand U12808 (N_12808,N_8994,N_5066);
xnor U12809 (N_12809,N_5877,N_2295);
nand U12810 (N_12810,N_2881,N_1664);
xor U12811 (N_12811,N_2846,N_5846);
and U12812 (N_12812,N_4924,N_3583);
nor U12813 (N_12813,N_2405,N_9067);
or U12814 (N_12814,N_7481,N_7275);
or U12815 (N_12815,N_487,N_5065);
and U12816 (N_12816,N_2423,N_1076);
and U12817 (N_12817,N_9722,N_4422);
xor U12818 (N_12818,N_8894,N_6680);
nor U12819 (N_12819,N_7725,N_8753);
and U12820 (N_12820,N_9111,N_8101);
nand U12821 (N_12821,N_9713,N_1234);
nand U12822 (N_12822,N_510,N_285);
nor U12823 (N_12823,N_8763,N_8895);
nand U12824 (N_12824,N_19,N_5185);
nand U12825 (N_12825,N_2558,N_8063);
or U12826 (N_12826,N_3777,N_4043);
nor U12827 (N_12827,N_9641,N_7243);
and U12828 (N_12828,N_7993,N_1935);
nand U12829 (N_12829,N_1700,N_2255);
nand U12830 (N_12830,N_5355,N_4812);
xor U12831 (N_12831,N_7790,N_4312);
nand U12832 (N_12832,N_3717,N_9885);
nor U12833 (N_12833,N_2919,N_4559);
nand U12834 (N_12834,N_4174,N_1248);
nor U12835 (N_12835,N_5272,N_7295);
nand U12836 (N_12836,N_1237,N_9686);
nand U12837 (N_12837,N_5677,N_7822);
and U12838 (N_12838,N_111,N_9993);
or U12839 (N_12839,N_4326,N_2765);
nor U12840 (N_12840,N_7819,N_1740);
nand U12841 (N_12841,N_9920,N_5540);
nand U12842 (N_12842,N_7066,N_1999);
or U12843 (N_12843,N_8009,N_504);
nand U12844 (N_12844,N_8977,N_5044);
nand U12845 (N_12845,N_976,N_6249);
xnor U12846 (N_12846,N_3904,N_2130);
or U12847 (N_12847,N_3768,N_5657);
and U12848 (N_12848,N_728,N_537);
nor U12849 (N_12849,N_1170,N_6657);
or U12850 (N_12850,N_2104,N_933);
nand U12851 (N_12851,N_3529,N_3434);
or U12852 (N_12852,N_6243,N_5148);
and U12853 (N_12853,N_4201,N_1817);
xnor U12854 (N_12854,N_6941,N_7350);
xor U12855 (N_12855,N_7974,N_5560);
or U12856 (N_12856,N_267,N_9600);
nor U12857 (N_12857,N_6659,N_4813);
nor U12858 (N_12858,N_4056,N_2921);
or U12859 (N_12859,N_4314,N_6792);
nor U12860 (N_12860,N_1794,N_3748);
nand U12861 (N_12861,N_6012,N_5792);
xor U12862 (N_12862,N_1315,N_3329);
and U12863 (N_12863,N_1362,N_1236);
and U12864 (N_12864,N_5030,N_374);
nor U12865 (N_12865,N_3449,N_9703);
nand U12866 (N_12866,N_2596,N_5997);
and U12867 (N_12867,N_853,N_5036);
xnor U12868 (N_12868,N_2252,N_4540);
or U12869 (N_12869,N_3676,N_3350);
or U12870 (N_12870,N_1884,N_4805);
nand U12871 (N_12871,N_9723,N_1146);
nor U12872 (N_12872,N_4659,N_1036);
and U12873 (N_12873,N_6411,N_661);
or U12874 (N_12874,N_3172,N_1135);
or U12875 (N_12875,N_16,N_2861);
or U12876 (N_12876,N_2574,N_5926);
or U12877 (N_12877,N_7704,N_1778);
or U12878 (N_12878,N_5919,N_6551);
and U12879 (N_12879,N_2163,N_6024);
or U12880 (N_12880,N_8042,N_4134);
nor U12881 (N_12881,N_5049,N_2908);
or U12882 (N_12882,N_7264,N_2471);
or U12883 (N_12883,N_7736,N_2789);
and U12884 (N_12884,N_9354,N_2014);
and U12885 (N_12885,N_1867,N_8006);
nand U12886 (N_12886,N_4455,N_2050);
nor U12887 (N_12887,N_7215,N_8417);
nor U12888 (N_12888,N_394,N_9065);
nor U12889 (N_12889,N_9357,N_9131);
nor U12890 (N_12890,N_8820,N_2395);
nand U12891 (N_12891,N_2752,N_5182);
or U12892 (N_12892,N_8443,N_7100);
nand U12893 (N_12893,N_4164,N_4077);
and U12894 (N_12894,N_4723,N_5360);
and U12895 (N_12895,N_5986,N_6685);
or U12896 (N_12896,N_6545,N_2731);
nand U12897 (N_12897,N_3492,N_5382);
and U12898 (N_12898,N_345,N_9706);
and U12899 (N_12899,N_299,N_2783);
and U12900 (N_12900,N_8636,N_5188);
nand U12901 (N_12901,N_6543,N_4544);
and U12902 (N_12902,N_3338,N_7653);
nor U12903 (N_12903,N_6581,N_922);
nand U12904 (N_12904,N_586,N_6142);
nor U12905 (N_12905,N_1426,N_8863);
nor U12906 (N_12906,N_970,N_2809);
nor U12907 (N_12907,N_3709,N_6675);
nor U12908 (N_12908,N_5622,N_2090);
nand U12909 (N_12909,N_3306,N_3462);
and U12910 (N_12910,N_1461,N_1091);
or U12911 (N_12911,N_5440,N_7191);
nand U12912 (N_12912,N_6273,N_6672);
or U12913 (N_12913,N_615,N_5202);
nand U12914 (N_12914,N_456,N_8287);
nor U12915 (N_12915,N_8983,N_3654);
xor U12916 (N_12916,N_1412,N_3948);
or U12917 (N_12917,N_4256,N_6810);
and U12918 (N_12918,N_9405,N_6816);
nor U12919 (N_12919,N_8563,N_6404);
nor U12920 (N_12920,N_5864,N_9738);
or U12921 (N_12921,N_5964,N_4342);
or U12922 (N_12922,N_5290,N_6902);
nor U12923 (N_12923,N_4586,N_560);
nor U12924 (N_12924,N_4210,N_8790);
or U12925 (N_12925,N_2,N_3018);
or U12926 (N_12926,N_1373,N_3073);
or U12927 (N_12927,N_5176,N_6906);
and U12928 (N_12928,N_4636,N_178);
and U12929 (N_12929,N_8689,N_9526);
or U12930 (N_12930,N_3129,N_7282);
nor U12931 (N_12931,N_2619,N_3725);
and U12932 (N_12932,N_3870,N_1570);
and U12933 (N_12933,N_5502,N_2827);
and U12934 (N_12934,N_1614,N_9359);
or U12935 (N_12935,N_6261,N_3532);
or U12936 (N_12936,N_6111,N_3776);
nand U12937 (N_12937,N_7033,N_649);
or U12938 (N_12938,N_7833,N_6156);
xnor U12939 (N_12939,N_7286,N_9279);
nor U12940 (N_12940,N_6605,N_2078);
nor U12941 (N_12941,N_7366,N_6782);
and U12942 (N_12942,N_2057,N_7768);
nand U12943 (N_12943,N_7193,N_3088);
or U12944 (N_12944,N_8921,N_4260);
and U12945 (N_12945,N_9300,N_6212);
nor U12946 (N_12946,N_7077,N_6580);
nor U12947 (N_12947,N_4097,N_3913);
nand U12948 (N_12948,N_9306,N_3511);
or U12949 (N_12949,N_8481,N_6597);
and U12950 (N_12950,N_5659,N_4404);
xor U12951 (N_12951,N_2122,N_712);
nor U12952 (N_12952,N_988,N_4884);
nand U12953 (N_12953,N_2661,N_5315);
nor U12954 (N_12954,N_243,N_9034);
and U12955 (N_12955,N_338,N_7023);
or U12956 (N_12956,N_3682,N_5318);
and U12957 (N_12957,N_7667,N_4680);
nand U12958 (N_12958,N_4118,N_5882);
xnor U12959 (N_12959,N_3989,N_5270);
or U12960 (N_12960,N_2111,N_6736);
nand U12961 (N_12961,N_8705,N_6827);
or U12962 (N_12962,N_3922,N_3677);
xnor U12963 (N_12963,N_4398,N_8635);
or U12964 (N_12964,N_3572,N_8586);
nor U12965 (N_12965,N_1786,N_6814);
and U12966 (N_12966,N_5297,N_2983);
nor U12967 (N_12967,N_764,N_1907);
nor U12968 (N_12968,N_4594,N_5607);
nor U12969 (N_12969,N_3276,N_633);
xor U12970 (N_12970,N_960,N_3781);
nor U12971 (N_12971,N_8162,N_7863);
nor U12972 (N_12972,N_2953,N_5361);
nand U12973 (N_12973,N_7305,N_8097);
nand U12974 (N_12974,N_6604,N_9011);
and U12975 (N_12975,N_2868,N_6824);
or U12976 (N_12976,N_8834,N_4621);
nor U12977 (N_12977,N_2336,N_3232);
and U12978 (N_12978,N_8244,N_8032);
nand U12979 (N_12979,N_7914,N_6577);
nor U12980 (N_12980,N_1651,N_7310);
and U12981 (N_12981,N_5326,N_5444);
nand U12982 (N_12982,N_7690,N_2999);
xor U12983 (N_12983,N_2394,N_5405);
and U12984 (N_12984,N_1558,N_2564);
xor U12985 (N_12985,N_6250,N_2956);
nand U12986 (N_12986,N_7565,N_2928);
xor U12987 (N_12987,N_3800,N_5718);
nand U12988 (N_12988,N_2270,N_4769);
nor U12989 (N_12989,N_7267,N_6516);
or U12990 (N_12990,N_4941,N_3772);
xor U12991 (N_12991,N_3207,N_5467);
and U12992 (N_12992,N_4705,N_4937);
nor U12993 (N_12993,N_7828,N_5549);
nor U12994 (N_12994,N_7887,N_9867);
or U12995 (N_12995,N_3592,N_2096);
or U12996 (N_12996,N_5059,N_138);
nand U12997 (N_12997,N_7313,N_426);
and U12998 (N_12998,N_4073,N_9985);
and U12999 (N_12999,N_3406,N_4396);
nand U13000 (N_13000,N_3628,N_8338);
nand U13001 (N_13001,N_9185,N_5225);
nor U13002 (N_13002,N_6766,N_319);
and U13003 (N_13003,N_4389,N_5462);
nor U13004 (N_13004,N_715,N_695);
and U13005 (N_13005,N_9594,N_8634);
nor U13006 (N_13006,N_5842,N_1518);
or U13007 (N_13007,N_7087,N_814);
or U13008 (N_13008,N_8526,N_4758);
nor U13009 (N_13009,N_4869,N_7300);
nor U13010 (N_13010,N_1766,N_9654);
or U13011 (N_13011,N_6891,N_3428);
and U13012 (N_13012,N_4883,N_7308);
xnor U13013 (N_13013,N_5473,N_1385);
or U13014 (N_13014,N_7247,N_9192);
nand U13015 (N_13015,N_3226,N_663);
nand U13016 (N_13016,N_3782,N_5442);
nand U13017 (N_13017,N_9890,N_2008);
nor U13018 (N_13018,N_4774,N_4542);
xor U13019 (N_13019,N_8519,N_6384);
or U13020 (N_13020,N_6666,N_8100);
nor U13021 (N_13021,N_4279,N_697);
nor U13022 (N_13022,N_4383,N_3405);
and U13023 (N_13023,N_6992,N_6452);
xor U13024 (N_13024,N_7255,N_8494);
nand U13025 (N_13025,N_2517,N_9990);
nand U13026 (N_13026,N_2957,N_9959);
nand U13027 (N_13027,N_1217,N_5680);
nand U13028 (N_13028,N_9506,N_4771);
and U13029 (N_13029,N_3261,N_89);
and U13030 (N_13030,N_7422,N_9267);
xnor U13031 (N_13031,N_502,N_8614);
nor U13032 (N_13032,N_562,N_3173);
nand U13033 (N_13033,N_9495,N_9322);
nor U13034 (N_13034,N_2916,N_2493);
and U13035 (N_13035,N_8195,N_3007);
and U13036 (N_13036,N_9488,N_1464);
nand U13037 (N_13037,N_4495,N_1801);
and U13038 (N_13038,N_6444,N_9148);
or U13039 (N_13039,N_8549,N_1099);
nand U13040 (N_13040,N_3681,N_6959);
nor U13041 (N_13041,N_4145,N_1468);
nor U13042 (N_13042,N_3790,N_1252);
and U13043 (N_13043,N_7602,N_9980);
nand U13044 (N_13044,N_8216,N_7238);
and U13045 (N_13045,N_3043,N_7157);
nand U13046 (N_13046,N_848,N_9924);
xnor U13047 (N_13047,N_3199,N_8187);
and U13048 (N_13048,N_7918,N_9740);
or U13049 (N_13049,N_1045,N_723);
and U13050 (N_13050,N_7956,N_1615);
and U13051 (N_13051,N_33,N_3470);
or U13052 (N_13052,N_5818,N_3527);
or U13053 (N_13053,N_3761,N_6770);
and U13054 (N_13054,N_3367,N_4778);
xnor U13055 (N_13055,N_177,N_7161);
nand U13056 (N_13056,N_7525,N_954);
nor U13057 (N_13057,N_6450,N_1342);
and U13058 (N_13058,N_9549,N_7949);
nand U13059 (N_13059,N_6625,N_6181);
nand U13060 (N_13060,N_8392,N_1975);
or U13061 (N_13061,N_7158,N_2339);
or U13062 (N_13062,N_1603,N_6719);
nand U13063 (N_13063,N_2228,N_8553);
xor U13064 (N_13064,N_9413,N_6905);
xor U13065 (N_13065,N_4085,N_1404);
and U13066 (N_13066,N_3886,N_9661);
or U13067 (N_13067,N_5247,N_8116);
nor U13068 (N_13068,N_4206,N_7666);
nand U13069 (N_13069,N_4786,N_6673);
and U13070 (N_13070,N_1536,N_4558);
or U13071 (N_13071,N_3429,N_9749);
and U13072 (N_13072,N_5580,N_7293);
and U13073 (N_13073,N_6723,N_4293);
xor U13074 (N_13074,N_6663,N_5960);
xor U13075 (N_13075,N_540,N_8993);
nor U13076 (N_13076,N_4546,N_3322);
nand U13077 (N_13077,N_7413,N_6419);
nand U13078 (N_13078,N_857,N_4113);
or U13079 (N_13079,N_5850,N_6616);
nand U13080 (N_13080,N_8396,N_6478);
nand U13081 (N_13081,N_3541,N_2177);
nand U13082 (N_13082,N_5949,N_7471);
or U13083 (N_13083,N_8932,N_9409);
or U13084 (N_13084,N_9122,N_6679);
or U13085 (N_13085,N_4932,N_5345);
xnor U13086 (N_13086,N_1707,N_3959);
nand U13087 (N_13087,N_796,N_7594);
and U13088 (N_13088,N_3059,N_9389);
nand U13089 (N_13089,N_1842,N_9845);
nand U13090 (N_13090,N_7657,N_6928);
and U13091 (N_13091,N_5455,N_5829);
xor U13092 (N_13092,N_4133,N_5192);
nand U13093 (N_13093,N_6433,N_3980);
nor U13094 (N_13094,N_3523,N_3212);
nand U13095 (N_13095,N_4238,N_8047);
nand U13096 (N_13096,N_4392,N_3327);
nor U13097 (N_13097,N_4220,N_953);
xnor U13098 (N_13098,N_2022,N_7553);
nand U13099 (N_13099,N_3418,N_4124);
nor U13100 (N_13100,N_6655,N_2632);
nand U13101 (N_13101,N_4037,N_5584);
nor U13102 (N_13102,N_2216,N_2346);
nor U13103 (N_13103,N_4907,N_2584);
and U13104 (N_13104,N_5900,N_5944);
or U13105 (N_13105,N_9308,N_1483);
or U13106 (N_13106,N_3739,N_2535);
and U13107 (N_13107,N_4463,N_3194);
xnor U13108 (N_13108,N_2375,N_4638);
nor U13109 (N_13109,N_6754,N_1122);
nor U13110 (N_13110,N_5067,N_7041);
or U13111 (N_13111,N_9852,N_9231);
nand U13112 (N_13112,N_7436,N_6748);
and U13113 (N_13113,N_9344,N_1054);
or U13114 (N_13114,N_7991,N_1372);
nand U13115 (N_13115,N_8752,N_7560);
nor U13116 (N_13116,N_6185,N_5542);
and U13117 (N_13117,N_6945,N_1418);
and U13118 (N_13118,N_6787,N_6882);
nand U13119 (N_13119,N_6310,N_2310);
and U13120 (N_13120,N_7687,N_8291);
nor U13121 (N_13121,N_2573,N_1542);
and U13122 (N_13122,N_6382,N_7409);
nor U13123 (N_13123,N_7534,N_7967);
and U13124 (N_13124,N_1165,N_5111);
xor U13125 (N_13125,N_5548,N_8308);
xnor U13126 (N_13126,N_2259,N_1440);
or U13127 (N_13127,N_6190,N_8623);
nand U13128 (N_13128,N_5743,N_5687);
and U13129 (N_13129,N_3444,N_350);
or U13130 (N_13130,N_8658,N_714);
and U13131 (N_13131,N_1366,N_6838);
and U13132 (N_13132,N_5768,N_9690);
nand U13133 (N_13133,N_7201,N_3602);
or U13134 (N_13134,N_8068,N_8175);
and U13135 (N_13135,N_149,N_1479);
nand U13136 (N_13136,N_6028,N_8961);
nor U13137 (N_13137,N_9397,N_251);
nand U13138 (N_13138,N_5671,N_6522);
and U13139 (N_13139,N_8030,N_4752);
and U13140 (N_13140,N_6333,N_7792);
xnor U13141 (N_13141,N_7641,N_9836);
or U13142 (N_13142,N_9403,N_7784);
nand U13143 (N_13143,N_3630,N_980);
and U13144 (N_13144,N_787,N_825);
nor U13145 (N_13145,N_914,N_3192);
or U13146 (N_13146,N_5074,N_4566);
nor U13147 (N_13147,N_9901,N_5564);
xor U13148 (N_13148,N_7454,N_6200);
or U13149 (N_13149,N_1476,N_8868);
and U13150 (N_13150,N_7941,N_158);
or U13151 (N_13151,N_8389,N_1023);
xor U13152 (N_13152,N_7030,N_3031);
nand U13153 (N_13153,N_7622,N_1375);
or U13154 (N_13154,N_2329,N_6225);
nand U13155 (N_13155,N_4095,N_8690);
nor U13156 (N_13156,N_9759,N_7683);
and U13157 (N_13157,N_9455,N_5408);
nand U13158 (N_13158,N_5796,N_2166);
nor U13159 (N_13159,N_547,N_6485);
nor U13160 (N_13160,N_9518,N_5618);
and U13161 (N_13161,N_931,N_7465);
or U13162 (N_13162,N_2541,N_7042);
nor U13163 (N_13163,N_5335,N_2566);
and U13164 (N_13164,N_8070,N_9430);
xor U13165 (N_13165,N_304,N_5356);
nand U13166 (N_13166,N_738,N_6490);
and U13167 (N_13167,N_4875,N_3483);
nor U13168 (N_13168,N_6826,N_6973);
or U13169 (N_13169,N_4303,N_8456);
xnor U13170 (N_13170,N_5880,N_8831);
nor U13171 (N_13171,N_391,N_946);
nor U13172 (N_13172,N_9538,N_5945);
and U13173 (N_13173,N_1520,N_3814);
nand U13174 (N_13174,N_9905,N_3069);
and U13175 (N_13175,N_8601,N_8248);
and U13176 (N_13176,N_8067,N_1454);
nor U13177 (N_13177,N_2969,N_7064);
nor U13178 (N_13178,N_6425,N_2813);
and U13179 (N_13179,N_858,N_8644);
nand U13180 (N_13180,N_6182,N_9744);
nand U13181 (N_13181,N_7880,N_2801);
or U13182 (N_13182,N_297,N_9677);
nand U13183 (N_13183,N_7608,N_6984);
nor U13184 (N_13184,N_9693,N_1047);
nand U13185 (N_13185,N_3036,N_557);
nand U13186 (N_13186,N_6544,N_7590);
or U13187 (N_13187,N_2215,N_8771);
xnor U13188 (N_13188,N_8904,N_325);
xor U13189 (N_13189,N_1003,N_7672);
and U13190 (N_13190,N_9812,N_5401);
or U13191 (N_13191,N_5142,N_5018);
and U13192 (N_13192,N_7045,N_6783);
nand U13193 (N_13193,N_2211,N_7032);
and U13194 (N_13194,N_3930,N_9524);
nor U13195 (N_13195,N_1675,N_6049);
or U13196 (N_13196,N_4366,N_7065);
nand U13197 (N_13197,N_8780,N_5008);
and U13198 (N_13198,N_7227,N_9683);
nand U13199 (N_13199,N_5380,N_3573);
or U13200 (N_13200,N_5214,N_7483);
nand U13201 (N_13201,N_2267,N_198);
and U13202 (N_13202,N_9788,N_8716);
and U13203 (N_13203,N_6542,N_2590);
or U13204 (N_13204,N_2641,N_9273);
or U13205 (N_13205,N_2374,N_6466);
nor U13206 (N_13206,N_1724,N_9085);
nor U13207 (N_13207,N_2315,N_5294);
nor U13208 (N_13208,N_6327,N_3133);
and U13209 (N_13209,N_5386,N_9903);
nor U13210 (N_13210,N_8695,N_4190);
nand U13211 (N_13211,N_3770,N_9171);
and U13212 (N_13212,N_2859,N_7576);
or U13213 (N_13213,N_7963,N_3791);
and U13214 (N_13214,N_9787,N_847);
nor U13215 (N_13215,N_6137,N_5518);
xor U13216 (N_13216,N_3860,N_7854);
nor U13217 (N_13217,N_6627,N_5735);
and U13218 (N_13218,N_3153,N_3750);
nand U13219 (N_13219,N_8737,N_5097);
xor U13220 (N_13220,N_1578,N_4081);
and U13221 (N_13221,N_7773,N_5121);
or U13222 (N_13222,N_625,N_6319);
nor U13223 (N_13223,N_4517,N_6571);
nand U13224 (N_13224,N_3057,N_7532);
nor U13225 (N_13225,N_1721,N_938);
and U13226 (N_13226,N_2123,N_355);
nand U13227 (N_13227,N_1261,N_5891);
nand U13228 (N_13228,N_3490,N_184);
or U13229 (N_13229,N_7775,N_8098);
nand U13230 (N_13230,N_3506,N_3648);
nor U13231 (N_13231,N_3785,N_5152);
xor U13232 (N_13232,N_2444,N_9697);
or U13233 (N_13233,N_8172,N_4692);
or U13234 (N_13234,N_2334,N_6658);
or U13235 (N_13235,N_5172,N_3687);
nor U13236 (N_13236,N_6312,N_1544);
nor U13237 (N_13237,N_7271,N_7252);
xnor U13238 (N_13238,N_5004,N_9750);
nor U13239 (N_13239,N_2749,N_8356);
nand U13240 (N_13240,N_9063,N_698);
or U13241 (N_13241,N_4170,N_5339);
xor U13242 (N_13242,N_9076,N_1735);
nand U13243 (N_13243,N_8345,N_9444);
nand U13244 (N_13244,N_9916,N_3137);
or U13245 (N_13245,N_444,N_4864);
or U13246 (N_13246,N_4643,N_5307);
xor U13247 (N_13247,N_5726,N_7221);
and U13248 (N_13248,N_4014,N_3533);
and U13249 (N_13249,N_1151,N_7694);
or U13250 (N_13250,N_4400,N_533);
nor U13251 (N_13251,N_2202,N_7046);
and U13252 (N_13252,N_2305,N_4011);
nand U13253 (N_13253,N_9729,N_3106);
or U13254 (N_13254,N_9134,N_8302);
and U13255 (N_13255,N_8669,N_4934);
nor U13256 (N_13256,N_9717,N_3228);
nand U13257 (N_13257,N_9887,N_6785);
or U13258 (N_13258,N_7203,N_9189);
nor U13259 (N_13259,N_2167,N_4359);
or U13260 (N_13260,N_8297,N_610);
nand U13261 (N_13261,N_2196,N_1818);
nor U13262 (N_13262,N_7541,N_8675);
and U13263 (N_13263,N_983,N_3902);
nor U13264 (N_13264,N_5129,N_5881);
nand U13265 (N_13265,N_5050,N_7699);
xnor U13266 (N_13266,N_3671,N_7431);
and U13267 (N_13267,N_489,N_7917);
or U13268 (N_13268,N_9275,N_4473);
nor U13269 (N_13269,N_5930,N_4948);
or U13270 (N_13270,N_3912,N_6617);
nand U13271 (N_13271,N_1398,N_7138);
or U13272 (N_13272,N_6422,N_7360);
nand U13273 (N_13273,N_4935,N_7973);
nor U13274 (N_13274,N_9982,N_7392);
nor U13275 (N_13275,N_993,N_9417);
nor U13276 (N_13276,N_4949,N_414);
nand U13277 (N_13277,N_6939,N_9442);
or U13278 (N_13278,N_3792,N_3940);
or U13279 (N_13279,N_1396,N_2925);
xor U13280 (N_13280,N_5772,N_7116);
or U13281 (N_13281,N_2981,N_1082);
nand U13282 (N_13282,N_5255,N_146);
or U13283 (N_13283,N_8154,N_3090);
and U13284 (N_13284,N_7947,N_4787);
and U13285 (N_13285,N_4804,N_8271);
nand U13286 (N_13286,N_1039,N_5983);
nor U13287 (N_13287,N_7027,N_6295);
or U13288 (N_13288,N_8544,N_7821);
and U13289 (N_13289,N_8649,N_7391);
nor U13290 (N_13290,N_7010,N_7872);
nor U13291 (N_13291,N_8903,N_1915);
nand U13292 (N_13292,N_6375,N_3401);
and U13293 (N_13293,N_8352,N_14);
nand U13294 (N_13294,N_2882,N_4796);
or U13295 (N_13295,N_6588,N_1832);
and U13296 (N_13296,N_972,N_7497);
or U13297 (N_13297,N_7946,N_9675);
and U13298 (N_13298,N_748,N_4219);
or U13299 (N_13299,N_978,N_4379);
or U13300 (N_13300,N_5320,N_4031);
xnor U13301 (N_13301,N_4930,N_2214);
xor U13302 (N_13302,N_8693,N_8545);
or U13303 (N_13303,N_6177,N_882);
nand U13304 (N_13304,N_7446,N_4143);
nand U13305 (N_13305,N_3046,N_3060);
or U13306 (N_13306,N_1110,N_3200);
nand U13307 (N_13307,N_7496,N_552);
and U13308 (N_13308,N_1147,N_296);
nor U13309 (N_13309,N_8951,N_3371);
or U13310 (N_13310,N_8249,N_9601);
and U13311 (N_13311,N_472,N_8487);
xor U13312 (N_13312,N_4565,N_8113);
or U13313 (N_13313,N_9350,N_4776);
nor U13314 (N_13314,N_3852,N_4202);
xor U13315 (N_13315,N_1381,N_9796);
and U13316 (N_13316,N_2629,N_4577);
and U13317 (N_13317,N_7860,N_7073);
or U13318 (N_13318,N_2028,N_8988);
nor U13319 (N_13319,N_3710,N_4088);
xnor U13320 (N_13320,N_404,N_9278);
nand U13321 (N_13321,N_7815,N_3357);
nand U13322 (N_13322,N_9871,N_4105);
nor U13323 (N_13323,N_1967,N_4957);
nand U13324 (N_13324,N_7763,N_5535);
or U13325 (N_13325,N_1188,N_9302);
xor U13326 (N_13326,N_7290,N_7797);
or U13327 (N_13327,N_4128,N_1661);
and U13328 (N_13328,N_1467,N_7945);
or U13329 (N_13329,N_5438,N_7521);
nor U13330 (N_13330,N_7140,N_3714);
and U13331 (N_13331,N_5778,N_7188);
or U13332 (N_13332,N_2136,N_1709);
and U13333 (N_13333,N_2021,N_996);
and U13334 (N_13334,N_1489,N_498);
and U13335 (N_13335,N_5484,N_76);
nor U13336 (N_13336,N_3452,N_5716);
or U13337 (N_13337,N_9154,N_9748);
or U13338 (N_13338,N_4177,N_8170);
nor U13339 (N_13339,N_9630,N_9960);
nor U13340 (N_13340,N_1576,N_6339);
nor U13341 (N_13341,N_1113,N_8516);
nand U13342 (N_13342,N_4477,N_2851);
or U13343 (N_13343,N_6896,N_117);
and U13344 (N_13344,N_6203,N_8502);
and U13345 (N_13345,N_1687,N_2609);
or U13346 (N_13346,N_6299,N_611);
xor U13347 (N_13347,N_3393,N_1767);
nor U13348 (N_13348,N_2725,N_2190);
nand U13349 (N_13349,N_6689,N_210);
nor U13350 (N_13350,N_9092,N_4001);
and U13351 (N_13351,N_4832,N_7178);
nand U13352 (N_13352,N_837,N_8005);
and U13353 (N_13353,N_7183,N_4446);
nor U13354 (N_13354,N_9688,N_1894);
and U13355 (N_13355,N_8797,N_8085);
nor U13356 (N_13356,N_9264,N_2507);
and U13357 (N_13357,N_5212,N_8840);
and U13358 (N_13358,N_485,N_182);
nand U13359 (N_13359,N_87,N_2268);
nor U13360 (N_13360,N_8642,N_3230);
or U13361 (N_13361,N_2069,N_6192);
and U13362 (N_13362,N_1397,N_5492);
or U13363 (N_13363,N_3014,N_336);
or U13364 (N_13364,N_5435,N_8952);
nand U13365 (N_13365,N_8442,N_272);
nor U13366 (N_13366,N_5587,N_885);
or U13367 (N_13367,N_5647,N_5417);
and U13368 (N_13368,N_9876,N_7475);
nand U13369 (N_13369,N_6637,N_9741);
and U13370 (N_13370,N_737,N_7632);
or U13371 (N_13371,N_600,N_4868);
nor U13372 (N_13372,N_3101,N_5912);
nor U13373 (N_13373,N_5897,N_3346);
nand U13374 (N_13374,N_157,N_8374);
or U13375 (N_13375,N_4110,N_7289);
or U13376 (N_13376,N_4852,N_9301);
and U13377 (N_13377,N_1365,N_223);
and U13378 (N_13378,N_6899,N_4639);
or U13379 (N_13379,N_3803,N_3352);
nor U13380 (N_13380,N_8871,N_4243);
or U13381 (N_13381,N_9617,N_7171);
nand U13382 (N_13382,N_8774,N_2161);
nand U13383 (N_13383,N_5989,N_1798);
or U13384 (N_13384,N_2422,N_1950);
and U13385 (N_13385,N_8084,N_518);
nor U13386 (N_13386,N_1055,N_7292);
nor U13387 (N_13387,N_1105,N_8014);
xor U13388 (N_13388,N_7837,N_5443);
nor U13389 (N_13389,N_985,N_8899);
or U13390 (N_13390,N_9667,N_631);
or U13391 (N_13391,N_3884,N_9479);
or U13392 (N_13392,N_9368,N_8225);
nor U13393 (N_13393,N_4962,N_2954);
nor U13394 (N_13394,N_1836,N_7448);
nand U13395 (N_13395,N_3744,N_6460);
and U13396 (N_13396,N_7291,N_6640);
nand U13397 (N_13397,N_1595,N_9072);
nand U13398 (N_13398,N_8548,N_2341);
nor U13399 (N_13399,N_8370,N_4906);
and U13400 (N_13400,N_8976,N_5285);
nand U13401 (N_13401,N_4176,N_5421);
nand U13402 (N_13402,N_7976,N_8906);
nand U13403 (N_13403,N_8427,N_7809);
and U13404 (N_13404,N_4530,N_4590);
nor U13405 (N_13405,N_5383,N_3465);
nand U13406 (N_13406,N_7980,N_7587);
and U13407 (N_13407,N_2748,N_3116);
or U13408 (N_13408,N_492,N_1004);
nor U13409 (N_13409,N_1952,N_7081);
nor U13410 (N_13410,N_2871,N_7480);
nor U13411 (N_13411,N_9415,N_4028);
and U13412 (N_13412,N_5670,N_5169);
nand U13413 (N_13413,N_8928,N_4150);
nor U13414 (N_13414,N_3034,N_1285);
nand U13415 (N_13415,N_9294,N_5857);
or U13416 (N_13416,N_8585,N_8326);
or U13417 (N_13417,N_9830,N_2325);
nand U13418 (N_13418,N_1910,N_4837);
and U13419 (N_13419,N_3082,N_4681);
and U13420 (N_13420,N_1470,N_37);
nand U13421 (N_13421,N_1027,N_8997);
nor U13422 (N_13422,N_3641,N_3999);
nand U13423 (N_13423,N_3741,N_2371);
xor U13424 (N_13424,N_8003,N_6027);
and U13425 (N_13425,N_2645,N_2728);
nor U13426 (N_13426,N_4927,N_3718);
and U13427 (N_13427,N_2421,N_8966);
nand U13428 (N_13428,N_3794,N_8311);
xnor U13429 (N_13429,N_9033,N_2321);
and U13430 (N_13430,N_332,N_8518);
xor U13431 (N_13431,N_1281,N_314);
nand U13432 (N_13432,N_4365,N_8460);
nand U13433 (N_13433,N_752,N_588);
nand U13434 (N_13434,N_9137,N_8000);
xor U13435 (N_13435,N_2724,N_8140);
nand U13436 (N_13436,N_658,N_7396);
or U13437 (N_13437,N_2367,N_5244);
nand U13438 (N_13438,N_5932,N_8382);
nand U13439 (N_13439,N_8587,N_6608);
or U13440 (N_13440,N_3410,N_718);
and U13441 (N_13441,N_8332,N_3960);
and U13442 (N_13442,N_1015,N_2318);
or U13443 (N_13443,N_9806,N_2862);
nand U13444 (N_13444,N_2875,N_7127);
xnor U13445 (N_13445,N_731,N_4414);
nand U13446 (N_13446,N_5106,N_3758);
nand U13447 (N_13447,N_8078,N_2991);
or U13448 (N_13448,N_3013,N_2071);
or U13449 (N_13449,N_5755,N_8038);
nor U13450 (N_13450,N_4903,N_6326);
nand U13451 (N_13451,N_5720,N_4273);
or U13452 (N_13452,N_5181,N_7304);
and U13453 (N_13453,N_8255,N_7373);
nor U13454 (N_13454,N_2086,N_6158);
or U13455 (N_13455,N_7543,N_368);
and U13456 (N_13456,N_6483,N_2392);
nor U13457 (N_13457,N_8145,N_8598);
nor U13458 (N_13458,N_4537,N_1511);
or U13459 (N_13459,N_6683,N_5314);
and U13460 (N_13460,N_3915,N_1360);
and U13461 (N_13461,N_5371,N_8607);
xnor U13462 (N_13462,N_73,N_3609);
and U13463 (N_13463,N_7752,N_6653);
or U13464 (N_13464,N_62,N_4944);
and U13465 (N_13465,N_9388,N_7615);
nand U13466 (N_13466,N_618,N_6269);
nand U13467 (N_13467,N_8505,N_7069);
nor U13468 (N_13468,N_3395,N_5865);
or U13469 (N_13469,N_3333,N_5862);
and U13470 (N_13470,N_9935,N_8473);
nand U13471 (N_13471,N_7189,N_5370);
nor U13472 (N_13472,N_8696,N_6529);
and U13473 (N_13473,N_4834,N_8893);
or U13474 (N_13474,N_2474,N_6003);
or U13475 (N_13475,N_8118,N_5834);
and U13476 (N_13476,N_145,N_9095);
nor U13477 (N_13477,N_6157,N_1156);
and U13478 (N_13478,N_5211,N_6045);
xnor U13479 (N_13479,N_833,N_4452);
and U13480 (N_13480,N_5216,N_8303);
nand U13481 (N_13481,N_8916,N_804);
and U13482 (N_13482,N_7978,N_8231);
nand U13483 (N_13483,N_1221,N_8324);
nor U13484 (N_13484,N_6798,N_3290);
nor U13485 (N_13485,N_9238,N_7536);
or U13486 (N_13486,N_1874,N_7732);
or U13487 (N_13487,N_9492,N_8127);
or U13488 (N_13488,N_3216,N_4872);
and U13489 (N_13489,N_1109,N_1080);
and U13490 (N_13490,N_4736,N_5507);
nand U13491 (N_13491,N_5266,N_8560);
nand U13492 (N_13492,N_1745,N_8228);
xnor U13493 (N_13493,N_7986,N_4251);
nor U13494 (N_13494,N_2431,N_8866);
or U13495 (N_13495,N_308,N_179);
or U13496 (N_13496,N_541,N_1963);
and U13497 (N_13497,N_2526,N_3243);
or U13498 (N_13498,N_2753,N_2085);
and U13499 (N_13499,N_9671,N_2931);
or U13500 (N_13500,N_5836,N_8577);
and U13501 (N_13501,N_7049,N_4092);
nor U13502 (N_13502,N_6253,N_1211);
nor U13503 (N_13503,N_6170,N_3349);
nor U13504 (N_13504,N_9971,N_4743);
and U13505 (N_13505,N_3412,N_3413);
and U13506 (N_13506,N_9247,N_316);
nor U13507 (N_13507,N_1106,N_7668);
nor U13508 (N_13508,N_5077,N_8239);
nand U13509 (N_13509,N_3526,N_4478);
nor U13510 (N_13510,N_373,N_3793);
nand U13511 (N_13511,N_4227,N_9334);
and U13512 (N_13512,N_8595,N_6878);
and U13513 (N_13513,N_232,N_246);
nor U13514 (N_13514,N_4990,N_6856);
nand U13515 (N_13515,N_8033,N_1466);
and U13516 (N_13516,N_1313,N_8259);
nor U13517 (N_13517,N_7850,N_8599);
nor U13518 (N_13518,N_7152,N_1782);
nand U13519 (N_13519,N_1424,N_2690);
nor U13520 (N_13520,N_6311,N_1543);
and U13521 (N_13521,N_6380,N_9801);
and U13522 (N_13522,N_2834,N_5591);
nand U13523 (N_13523,N_8628,N_9251);
xor U13524 (N_13524,N_4357,N_3552);
nand U13525 (N_13525,N_8847,N_1959);
nand U13526 (N_13526,N_6669,N_9180);
nand U13527 (N_13527,N_9569,N_1772);
nor U13528 (N_13528,N_8136,N_2788);
nand U13529 (N_13529,N_1880,N_1815);
xnor U13530 (N_13530,N_9428,N_5470);
nand U13531 (N_13531,N_432,N_9527);
nor U13532 (N_13532,N_4898,N_5232);
and U13533 (N_13533,N_1931,N_9281);
or U13534 (N_13534,N_4486,N_8959);
nand U13535 (N_13535,N_9822,N_6263);
and U13536 (N_13536,N_3551,N_7598);
and U13537 (N_13537,N_9291,N_4735);
or U13538 (N_13538,N_4433,N_4459);
nand U13539 (N_13539,N_629,N_1460);
xnor U13540 (N_13540,N_940,N_2974);
or U13541 (N_13541,N_1882,N_7581);
and U13542 (N_13542,N_5873,N_7969);
xor U13543 (N_13543,N_7134,N_5454);
nand U13544 (N_13544,N_1032,N_2362);
and U13545 (N_13545,N_1335,N_2236);
and U13546 (N_13546,N_3474,N_1859);
and U13547 (N_13547,N_3939,N_278);
or U13548 (N_13548,N_5554,N_1309);
or U13549 (N_13549,N_7838,N_5777);
or U13550 (N_13550,N_5667,N_9059);
nor U13551 (N_13551,N_9523,N_897);
or U13552 (N_13552,N_5242,N_7322);
and U13553 (N_13553,N_5604,N_7624);
and U13554 (N_13554,N_3599,N_6364);
nand U13555 (N_13555,N_2721,N_8394);
nor U13556 (N_13556,N_7216,N_9727);
and U13557 (N_13557,N_1747,N_3147);
or U13558 (N_13558,N_183,N_1898);
and U13559 (N_13559,N_1205,N_4510);
nand U13560 (N_13560,N_4255,N_925);
nand U13561 (N_13561,N_826,N_6751);
nand U13562 (N_13562,N_2811,N_9872);
nor U13563 (N_13563,N_407,N_3905);
and U13564 (N_13564,N_9719,N_3423);
and U13565 (N_13565,N_8373,N_2508);
nand U13566 (N_13566,N_5552,N_4437);
or U13567 (N_13567,N_4732,N_1892);
and U13568 (N_13568,N_9710,N_7574);
xnor U13569 (N_13569,N_3100,N_1169);
nand U13570 (N_13570,N_9386,N_4750);
or U13571 (N_13571,N_5388,N_5063);
and U13572 (N_13572,N_3394,N_1534);
or U13573 (N_13573,N_2218,N_4435);
nor U13574 (N_13574,N_3652,N_7762);
nand U13575 (N_13575,N_5249,N_2589);
and U13576 (N_13576,N_1557,N_677);
and U13577 (N_13577,N_1784,N_2460);
xor U13578 (N_13578,N_4892,N_7533);
xnor U13579 (N_13579,N_7799,N_2247);
nor U13580 (N_13580,N_1000,N_4661);
or U13581 (N_13581,N_2710,N_3209);
or U13582 (N_13582,N_3666,N_8148);
nand U13583 (N_13583,N_3312,N_5402);
nand U13584 (N_13584,N_876,N_8215);
or U13585 (N_13585,N_657,N_8053);
nor U13586 (N_13586,N_7571,N_1469);
nor U13587 (N_13587,N_1789,N_5295);
nor U13588 (N_13588,N_3993,N_8289);
nor U13589 (N_13589,N_810,N_7758);
and U13590 (N_13590,N_1929,N_9682);
and U13591 (N_13591,N_3559,N_1506);
and U13592 (N_13592,N_9503,N_1790);
nand U13593 (N_13593,N_6573,N_3450);
nor U13594 (N_13594,N_873,N_3997);
and U13595 (N_13595,N_2292,N_3326);
or U13596 (N_13596,N_4155,N_3728);
or U13597 (N_13597,N_7226,N_7540);
nor U13598 (N_13598,N_7133,N_6387);
nor U13599 (N_13599,N_3925,N_7988);
and U13600 (N_13600,N_1912,N_213);
nor U13601 (N_13601,N_4545,N_5861);
or U13602 (N_13602,N_5398,N_655);
or U13603 (N_13603,N_9534,N_6448);
nor U13604 (N_13604,N_4246,N_4321);
xnor U13605 (N_13605,N_9829,N_5240);
and U13606 (N_13606,N_1812,N_4485);
nor U13607 (N_13607,N_3517,N_6321);
or U13608 (N_13608,N_807,N_4690);
or U13609 (N_13609,N_1066,N_7234);
or U13610 (N_13610,N_2635,N_5222);
nor U13611 (N_13611,N_7795,N_7257);
and U13612 (N_13612,N_6279,N_8838);
nand U13613 (N_13613,N_9009,N_7136);
or U13614 (N_13614,N_9874,N_9515);
and U13615 (N_13615,N_1139,N_9720);
and U13616 (N_13616,N_3544,N_1791);
xor U13617 (N_13617,N_3855,N_1829);
nand U13618 (N_13618,N_5420,N_6082);
and U13619 (N_13619,N_6301,N_1293);
nor U13620 (N_13620,N_9387,N_1641);
nor U13621 (N_13621,N_5551,N_6779);
nor U13622 (N_13622,N_1581,N_6431);
nor U13623 (N_13623,N_7954,N_7640);
nor U13624 (N_13624,N_9477,N_956);
and U13625 (N_13625,N_9432,N_8794);
and U13626 (N_13626,N_3651,N_9537);
nand U13627 (N_13627,N_6530,N_4543);
nand U13628 (N_13628,N_4413,N_3193);
xor U13629 (N_13629,N_7057,N_5550);
nor U13630 (N_13630,N_8012,N_733);
or U13631 (N_13631,N_891,N_3464);
and U13632 (N_13632,N_8010,N_4746);
nand U13633 (N_13633,N_8610,N_6584);
nand U13634 (N_13634,N_8425,N_2930);
nor U13635 (N_13635,N_3525,N_6532);
or U13636 (N_13636,N_9271,N_3497);
or U13637 (N_13637,N_242,N_4607);
nor U13638 (N_13638,N_3062,N_5683);
nor U13639 (N_13639,N_7846,N_711);
nor U13640 (N_13640,N_1609,N_5461);
nor U13641 (N_13641,N_3921,N_2503);
nand U13642 (N_13642,N_6757,N_6837);
or U13643 (N_13643,N_2715,N_6913);
or U13644 (N_13644,N_4221,N_9844);
and U13645 (N_13645,N_7578,N_6238);
or U13646 (N_13646,N_1689,N_5174);
or U13647 (N_13647,N_4172,N_156);
nor U13648 (N_13648,N_3485,N_3617);
nand U13649 (N_13649,N_4651,N_9718);
nand U13650 (N_13650,N_2109,N_443);
xor U13651 (N_13651,N_999,N_155);
nand U13652 (N_13652,N_9708,N_5813);
nor U13653 (N_13653,N_3807,N_2303);
nor U13654 (N_13654,N_3023,N_2440);
or U13655 (N_13655,N_3995,N_5917);
or U13656 (N_13656,N_6229,N_8201);
or U13657 (N_13657,N_8420,N_3139);
xnor U13658 (N_13658,N_1858,N_5235);
nand U13659 (N_13659,N_3698,N_2937);
nor U13660 (N_13660,N_5527,N_8091);
or U13661 (N_13661,N_8235,N_5009);
or U13662 (N_13662,N_193,N_1922);
nand U13663 (N_13663,N_4239,N_9691);
nor U13664 (N_13664,N_7266,N_4998);
and U13665 (N_13665,N_1654,N_9989);
xor U13666 (N_13666,N_4838,N_7998);
and U13667 (N_13667,N_7084,N_4950);
nand U13668 (N_13668,N_5001,N_7794);
nand U13669 (N_13669,N_307,N_2668);
xnor U13670 (N_13670,N_3113,N_5411);
nand U13671 (N_13671,N_747,N_1899);
or U13672 (N_13672,N_7372,N_7150);
nor U13673 (N_13673,N_4674,N_6794);
nand U13674 (N_13674,N_9212,N_5902);
nor U13675 (N_13675,N_570,N_6670);
nor U13676 (N_13676,N_6793,N_9742);
and U13677 (N_13677,N_6795,N_546);
nand U13678 (N_13678,N_6122,N_6221);
or U13679 (N_13679,N_3653,N_4691);
and U13680 (N_13680,N_7528,N_9701);
or U13681 (N_13681,N_2112,N_8045);
and U13682 (N_13682,N_8621,N_8438);
nor U13683 (N_13683,N_4807,N_1384);
and U13684 (N_13684,N_3124,N_9648);
or U13685 (N_13685,N_7334,N_4773);
and U13686 (N_13686,N_7915,N_4741);
and U13687 (N_13687,N_5061,N_6732);
xnor U13688 (N_13688,N_3919,N_9846);
or U13689 (N_13689,N_1431,N_5363);
nor U13690 (N_13690,N_6377,N_3340);
and U13691 (N_13691,N_362,N_1893);
nand U13692 (N_13692,N_7103,N_4343);
nor U13693 (N_13693,N_3316,N_9747);
nor U13694 (N_13694,N_5226,N_4893);
nor U13695 (N_13695,N_7554,N_9239);
nand U13696 (N_13696,N_9947,N_7876);
xor U13697 (N_13697,N_4604,N_2335);
xnor U13698 (N_13698,N_8674,N_6952);
and U13699 (N_13699,N_3587,N_8795);
nand U13700 (N_13700,N_9687,N_6013);
and U13701 (N_13701,N_5840,N_8093);
and U13702 (N_13702,N_5812,N_7054);
or U13703 (N_13703,N_7911,N_1143);
or U13704 (N_13704,N_5605,N_6379);
nand U13705 (N_13705,N_4051,N_389);
or U13706 (N_13706,N_5103,N_9360);
and U13707 (N_13707,N_6852,N_1703);
nand U13708 (N_13708,N_767,N_5);
nor U13709 (N_13709,N_1531,N_1131);
or U13710 (N_13710,N_7893,N_3242);
nand U13711 (N_13711,N_5952,N_4212);
nand U13712 (N_13712,N_1639,N_8480);
nand U13713 (N_13713,N_2993,N_3521);
and U13714 (N_13714,N_2041,N_5929);
or U13715 (N_13715,N_9545,N_6153);
xor U13716 (N_13716,N_7433,N_225);
nor U13717 (N_13717,N_8949,N_9604);
xor U13718 (N_13718,N_6555,N_289);
nand U13719 (N_13719,N_7080,N_6276);
or U13720 (N_13720,N_9475,N_9540);
nand U13721 (N_13721,N_7078,N_2627);
nor U13722 (N_13722,N_2884,N_4099);
nor U13723 (N_13723,N_1759,N_6567);
xor U13724 (N_13724,N_519,N_4696);
or U13725 (N_13725,N_2299,N_3661);
nand U13726 (N_13726,N_3788,N_4006);
or U13727 (N_13727,N_5695,N_6329);
and U13728 (N_13728,N_9170,N_6351);
or U13729 (N_13729,N_5427,N_5476);
or U13730 (N_13730,N_3491,N_4960);
nor U13731 (N_13731,N_318,N_8583);
nor U13732 (N_13732,N_9733,N_7805);
xor U13733 (N_13733,N_8551,N_6737);
and U13734 (N_13734,N_8262,N_6099);
nand U13735 (N_13735,N_8701,N_4686);
nor U13736 (N_13736,N_7363,N_8082);
and U13737 (N_13737,N_3180,N_4493);
xor U13738 (N_13738,N_1132,N_9766);
nand U13739 (N_13739,N_6362,N_7879);
and U13740 (N_13740,N_3835,N_42);
nor U13741 (N_13741,N_6438,N_7008);
or U13742 (N_13742,N_7425,N_3786);
and U13743 (N_13743,N_4519,N_6702);
nor U13744 (N_13744,N_4921,N_9100);
nand U13745 (N_13745,N_341,N_7470);
or U13746 (N_13746,N_9058,N_187);
and U13747 (N_13747,N_7871,N_8212);
or U13748 (N_13748,N_494,N_2124);
xor U13749 (N_13749,N_8718,N_7345);
and U13750 (N_13750,N_4103,N_6062);
nand U13751 (N_13751,N_7878,N_8434);
nor U13752 (N_13752,N_2832,N_8639);
and U13753 (N_13753,N_4730,N_309);
or U13754 (N_13754,N_2316,N_6088);
nor U13755 (N_13755,N_6342,N_8340);
xnor U13756 (N_13756,N_2483,N_7200);
nand U13757 (N_13757,N_8433,N_8845);
nor U13758 (N_13758,N_7083,N_3155);
nor U13759 (N_13759,N_3440,N_101);
xor U13760 (N_13760,N_4966,N_5328);
and U13761 (N_13761,N_5931,N_9789);
nand U13762 (N_13762,N_7225,N_4237);
nor U13763 (N_13763,N_3998,N_7399);
nand U13764 (N_13764,N_7584,N_2979);
and U13765 (N_13765,N_5823,N_3738);
nor U13766 (N_13766,N_3809,N_5007);
and U13767 (N_13767,N_8589,N_9411);
nand U13768 (N_13768,N_1992,N_2171);
nand U13769 (N_13769,N_2663,N_8002);
and U13770 (N_13770,N_6309,N_9218);
and U13771 (N_13771,N_9614,N_9066);
nor U13772 (N_13772,N_9669,N_7115);
and U13773 (N_13773,N_1803,N_503);
nand U13774 (N_13774,N_7961,N_2492);
and U13775 (N_13775,N_1024,N_1408);
nand U13776 (N_13776,N_5603,N_4887);
and U13777 (N_13777,N_465,N_2695);
or U13778 (N_13778,N_408,N_6290);
and U13779 (N_13779,N_7995,N_2438);
or U13780 (N_13780,N_6194,N_792);
xor U13781 (N_13781,N_8633,N_3198);
or U13782 (N_13782,N_4469,N_791);
nand U13783 (N_13783,N_7390,N_7900);
nand U13784 (N_13784,N_8760,N_6472);
nand U13785 (N_13785,N_3731,N_3508);
nand U13786 (N_13786,N_3085,N_4652);
and U13787 (N_13787,N_5384,N_6678);
nand U13788 (N_13788,N_3161,N_7623);
or U13789 (N_13789,N_5215,N_3074);
nor U13790 (N_13790,N_5459,N_3589);
xnor U13791 (N_13791,N_3512,N_6589);
xnor U13792 (N_13792,N_399,N_2231);
and U13793 (N_13793,N_9764,N_5965);
and U13794 (N_13794,N_3109,N_6510);
or U13795 (N_13795,N_1995,N_5329);
nand U13796 (N_13796,N_843,N_1481);
or U13797 (N_13797,N_2426,N_3236);
or U13798 (N_13798,N_4646,N_6130);
xor U13799 (N_13799,N_2472,N_8756);
and U13800 (N_13800,N_6730,N_5143);
nand U13801 (N_13801,N_6061,N_2379);
and U13802 (N_13802,N_5806,N_1022);
nand U13803 (N_13803,N_9312,N_5025);
nor U13804 (N_13804,N_9037,N_5503);
nand U13805 (N_13805,N_6722,N_9658);
xnor U13806 (N_13806,N_4204,N_1329);
nor U13807 (N_13807,N_917,N_5883);
nand U13808 (N_13808,N_3131,N_6790);
or U13809 (N_13809,N_5981,N_1028);
and U13810 (N_13810,N_1071,N_7839);
nand U13811 (N_13811,N_5054,N_7192);
and U13812 (N_13812,N_2934,N_1449);
or U13813 (N_13813,N_1754,N_702);
and U13814 (N_13814,N_2864,N_1856);
xnor U13815 (N_13815,N_4533,N_2578);
or U13816 (N_13816,N_2744,N_7552);
and U13817 (N_13817,N_9936,N_9948);
and U13818 (N_13818,N_5341,N_8687);
and U13819 (N_13819,N_5972,N_7224);
or U13820 (N_13820,N_5620,N_3949);
and U13821 (N_13821,N_7463,N_8150);
and U13822 (N_13822,N_8258,N_3496);
nor U13823 (N_13823,N_1111,N_3277);
and U13824 (N_13824,N_757,N_9588);
or U13825 (N_13825,N_2525,N_3817);
or U13826 (N_13826,N_8956,N_1290);
nand U13827 (N_13827,N_9704,N_7357);
and U13828 (N_13828,N_1604,N_2275);
nor U13829 (N_13829,N_5702,N_646);
and U13830 (N_13830,N_6587,N_153);
and U13831 (N_13831,N_6767,N_1872);
nand U13832 (N_13832,N_3988,N_1186);
or U13833 (N_13833,N_7176,N_5463);
nor U13834 (N_13834,N_7130,N_3110);
or U13835 (N_13835,N_9314,N_4821);
and U13836 (N_13836,N_9414,N_1835);
xnor U13837 (N_13837,N_1202,N_31);
xnor U13838 (N_13838,N_7569,N_3825);
and U13839 (N_13839,N_9839,N_4706);
or U13840 (N_13840,N_6165,N_105);
or U13841 (N_13841,N_1738,N_5252);
and U13842 (N_13842,N_9620,N_1771);
nand U13843 (N_13843,N_288,N_3540);
and U13844 (N_13844,N_9508,N_7428);
nor U13845 (N_13845,N_9347,N_361);
or U13846 (N_13846,N_3690,N_6314);
or U13847 (N_13847,N_4038,N_5943);
or U13848 (N_13848,N_2958,N_4100);
or U13849 (N_13849,N_4280,N_1072);
nor U13850 (N_13850,N_8650,N_1161);
nor U13851 (N_13851,N_1574,N_587);
and U13852 (N_13852,N_5565,N_9036);
and U13853 (N_13853,N_2182,N_5978);
nand U13854 (N_13854,N_2538,N_7770);
or U13855 (N_13855,N_4983,N_2010);
nor U13856 (N_13856,N_9653,N_8376);
xor U13857 (N_13857,N_4335,N_496);
and U13858 (N_13858,N_5093,N_9610);
nor U13859 (N_13859,N_9031,N_1288);
nor U13860 (N_13860,N_4101,N_7823);
nand U13861 (N_13861,N_6001,N_7071);
and U13862 (N_13862,N_9533,N_4292);
nand U13863 (N_13863,N_8119,N_3010);
and U13864 (N_13864,N_2704,N_8286);
and U13865 (N_13865,N_9953,N_2150);
nand U13866 (N_13866,N_9942,N_1662);
xnor U13867 (N_13867,N_8265,N_7681);
or U13868 (N_13868,N_6999,N_8284);
and U13869 (N_13869,N_824,N_8777);
or U13870 (N_13870,N_367,N_2865);
or U13871 (N_13871,N_9060,N_2608);
xnor U13872 (N_13872,N_8236,N_7567);
or U13873 (N_13873,N_9201,N_1005);
and U13874 (N_13874,N_1441,N_7604);
or U13875 (N_13875,N_2796,N_6841);
and U13876 (N_13876,N_8192,N_3274);
and U13877 (N_13877,N_140,N_1607);
nand U13878 (N_13878,N_9869,N_5228);
nand U13879 (N_13879,N_4532,N_6695);
xnor U13880 (N_13880,N_8141,N_2434);
nor U13881 (N_13881,N_6594,N_4524);
and U13882 (N_13882,N_4945,N_2194);
or U13883 (N_13883,N_6558,N_7646);
nor U13884 (N_13884,N_6901,N_9292);
and U13885 (N_13885,N_4080,N_9910);
or U13886 (N_13886,N_2537,N_9904);
and U13887 (N_13887,N_2000,N_692);
nand U13888 (N_13888,N_7261,N_6317);
and U13889 (N_13889,N_3385,N_7254);
or U13890 (N_13890,N_454,N_4428);
nand U13891 (N_13891,N_4120,N_2996);
xor U13892 (N_13892,N_523,N_8550);
nor U13893 (N_13893,N_376,N_9282);
nor U13894 (N_13894,N_7337,N_2554);
or U13895 (N_13895,N_3361,N_388);
xor U13896 (N_13896,N_4005,N_8567);
or U13897 (N_13897,N_1437,N_6985);
nand U13898 (N_13898,N_4981,N_7444);
xor U13899 (N_13899,N_8331,N_4991);
or U13900 (N_13900,N_2830,N_1577);
nor U13901 (N_13901,N_4152,N_4911);
or U13902 (N_13902,N_1627,N_6259);
and U13903 (N_13903,N_5685,N_7162);
or U13904 (N_13904,N_6370,N_7281);
nor U13905 (N_13905,N_803,N_1491);
or U13906 (N_13906,N_7499,N_967);
nor U13907 (N_13907,N_2464,N_3558);
and U13908 (N_13908,N_7811,N_8942);
nor U13909 (N_13909,N_6739,N_3253);
nor U13910 (N_13910,N_5128,N_8362);
nand U13911 (N_13911,N_6231,N_9831);
xnor U13912 (N_13912,N_9575,N_3190);
xor U13913 (N_13913,N_2523,N_6480);
nand U13914 (N_13914,N_4984,N_2615);
nand U13915 (N_13915,N_1037,N_6602);
or U13916 (N_13916,N_4525,N_6745);
xnor U13917 (N_13917,N_8151,N_8337);
and U13918 (N_13918,N_2053,N_5319);
or U13919 (N_13919,N_5514,N_1299);
and U13920 (N_13920,N_7895,N_1331);
nor U13921 (N_13921,N_5759,N_6922);
xnor U13922 (N_13922,N_3971,N_5914);
nand U13923 (N_13923,N_7237,N_8766);
nor U13924 (N_13924,N_6622,N_2148);
nand U13925 (N_13925,N_7798,N_7294);
xnor U13926 (N_13926,N_7999,N_8488);
nor U13927 (N_13927,N_4682,N_8395);
nor U13928 (N_13928,N_2860,N_1802);
and U13929 (N_13929,N_2548,N_9712);
and U13930 (N_13930,N_6085,N_3351);
and U13931 (N_13931,N_5046,N_783);
xor U13932 (N_13932,N_6797,N_2594);
or U13933 (N_13933,N_228,N_7111);
and U13934 (N_13934,N_9252,N_166);
or U13935 (N_13935,N_830,N_2140);
nand U13936 (N_13936,N_1322,N_4616);
nand U13937 (N_13937,N_6880,N_1102);
nand U13938 (N_13938,N_5193,N_2220);
and U13939 (N_13939,N_2878,N_5149);
xor U13940 (N_13940,N_4402,N_7636);
nand U13941 (N_13941,N_1088,N_1726);
nor U13942 (N_13942,N_2253,N_466);
and U13943 (N_13943,N_4503,N_3966);
nand U13944 (N_13944,N_8143,N_4086);
or U13945 (N_13945,N_6065,N_9207);
nand U13946 (N_13946,N_6381,N_6363);
nor U13947 (N_13947,N_1405,N_5567);
nand U13948 (N_13948,N_4953,N_7777);
nor U13949 (N_13949,N_6047,N_7113);
or U13950 (N_13950,N_8218,N_8529);
and U13951 (N_13951,N_6248,N_3962);
or U13952 (N_13952,N_7228,N_5757);
or U13953 (N_13953,N_8998,N_1515);
or U13954 (N_13954,N_2242,N_3969);
nor U13955 (N_13955,N_4987,N_4728);
nand U13956 (N_13956,N_7400,N_8646);
nor U13957 (N_13957,N_7024,N_864);
or U13958 (N_13958,N_929,N_6538);
nor U13959 (N_13959,N_3961,N_3436);
xor U13960 (N_13960,N_1079,N_6570);
nor U13961 (N_13961,N_1029,N_5970);
or U13962 (N_13962,N_9529,N_8572);
and U13963 (N_13963,N_2107,N_5789);
or U13964 (N_13964,N_7718,N_3183);
and U13965 (N_13965,N_4913,N_902);
and U13966 (N_13966,N_8330,N_2407);
nand U13967 (N_13967,N_1063,N_8493);
nor U13968 (N_13968,N_7166,N_4669);
xnor U13969 (N_13969,N_6056,N_7347);
nor U13970 (N_13970,N_6477,N_5669);
or U13971 (N_13971,N_3565,N_5557);
nand U13972 (N_13972,N_2126,N_2533);
nor U13973 (N_13973,N_1843,N_6886);
xnor U13974 (N_13974,N_7717,N_8970);
nor U13975 (N_13975,N_8880,N_7393);
nand U13976 (N_13976,N_6772,N_1305);
or U13977 (N_13977,N_3958,N_4180);
and U13978 (N_13978,N_9974,N_4438);
and U13979 (N_13979,N_3291,N_8169);
and U13980 (N_13980,N_4125,N_9230);
or U13981 (N_13981,N_2797,N_9015);
or U13982 (N_13982,N_5196,N_4871);
nand U13983 (N_13983,N_2132,N_6504);
and U13984 (N_13984,N_2061,N_5300);
or U13985 (N_13985,N_7835,N_5637);
or U13986 (N_13986,N_4318,N_3269);
nor U13987 (N_13987,N_3001,N_7884);
xnor U13988 (N_13988,N_254,N_6325);
nor U13989 (N_13989,N_6938,N_147);
and U13990 (N_13990,N_5583,N_7970);
nor U13991 (N_13991,N_8537,N_2103);
and U13992 (N_13992,N_4632,N_2184);
nand U13993 (N_13993,N_4748,N_3235);
and U13994 (N_13994,N_34,N_5572);
nor U13995 (N_13995,N_9562,N_536);
or U13996 (N_13996,N_9270,N_5991);
nor U13997 (N_13997,N_543,N_5497);
nor U13998 (N_13998,N_7512,N_5576);
nand U13999 (N_13999,N_1656,N_5475);
nor U14000 (N_14000,N_460,N_6096);
and U14001 (N_14001,N_9767,N_6771);
xor U14002 (N_14002,N_6784,N_7938);
or U14003 (N_14003,N_199,N_2284);
nor U14004 (N_14004,N_8887,N_9587);
nand U14005 (N_14005,N_1103,N_3859);
or U14006 (N_14006,N_8981,N_2705);
nor U14007 (N_14007,N_5975,N_8197);
xor U14008 (N_14008,N_5946,N_3263);
xnor U14009 (N_14009,N_8527,N_9244);
nor U14010 (N_14010,N_3588,N_9025);
and U14011 (N_14011,N_8917,N_3265);
nor U14012 (N_14012,N_3622,N_8681);
and U14013 (N_14013,N_9309,N_6189);
and U14014 (N_14014,N_1065,N_3865);
nor U14015 (N_14015,N_5161,N_5592);
or U14016 (N_14016,N_7473,N_7184);
nor U14017 (N_14017,N_865,N_9096);
and U14018 (N_14018,N_5091,N_2530);
or U14019 (N_14019,N_5512,N_949);
or U14020 (N_14020,N_3593,N_125);
and U14021 (N_14021,N_8371,N_7575);
nand U14022 (N_14022,N_6726,N_5915);
nand U14023 (N_14023,N_2902,N_9886);
nor U14024 (N_14024,N_4649,N_3684);
and U14025 (N_14025,N_4378,N_3826);
or U14026 (N_14026,N_6487,N_3679);
nor U14027 (N_14027,N_8057,N_9567);
nor U14028 (N_14028,N_312,N_7545);
or U14029 (N_14029,N_5275,N_3442);
and U14030 (N_14030,N_453,N_5933);
nand U14031 (N_14031,N_8530,N_2639);
and U14032 (N_14032,N_3285,N_7500);
xor U14033 (N_14033,N_6366,N_4078);
nor U14034 (N_14034,N_8743,N_7477);
and U14035 (N_14035,N_823,N_8884);
xnor U14036 (N_14036,N_5334,N_1002);
nand U14037 (N_14037,N_1566,N_8755);
and U14038 (N_14038,N_6741,N_2209);
nand U14039 (N_14039,N_9459,N_851);
or U14040 (N_14040,N_7478,N_2345);
and U14041 (N_14041,N_6684,N_1497);
xor U14042 (N_14042,N_9897,N_2447);
nor U14043 (N_14043,N_4835,N_6147);
or U14044 (N_14044,N_4488,N_3545);
nand U14045 (N_14045,N_1714,N_7788);
and U14046 (N_14046,N_7504,N_910);
xor U14047 (N_14047,N_8672,N_5642);
and U14048 (N_14048,N_4289,N_4411);
nand U14049 (N_14049,N_5123,N_1580);
nor U14050 (N_14050,N_3281,N_1166);
and U14051 (N_14051,N_3105,N_8251);
or U14052 (N_14052,N_6486,N_8021);
nand U14053 (N_14053,N_1436,N_8341);
nor U14054 (N_14054,N_5109,N_1334);
nand U14055 (N_14055,N_1136,N_6297);
nor U14056 (N_14056,N_4910,N_1349);
nand U14057 (N_14057,N_6098,N_2237);
nor U14058 (N_14058,N_6075,N_8733);
and U14059 (N_14059,N_9918,N_6423);
nor U14060 (N_14060,N_3650,N_1760);
or U14061 (N_14061,N_5346,N_2080);
and U14062 (N_14062,N_7589,N_8504);
nor U14063 (N_14063,N_8173,N_4992);
nor U14064 (N_14064,N_9542,N_2763);
nand U14065 (N_14065,N_7864,N_8854);
xor U14066 (N_14066,N_5358,N_3348);
and U14067 (N_14067,N_4091,N_2771);
or U14068 (N_14068,N_3673,N_119);
and U14069 (N_14069,N_8263,N_9117);
nor U14070 (N_14070,N_8778,N_1018);
nor U14071 (N_14071,N_6178,N_7285);
nand U14072 (N_14072,N_8491,N_8865);
xor U14073 (N_14073,N_1644,N_5579);
or U14074 (N_14074,N_9254,N_4013);
and U14075 (N_14075,N_6018,N_1346);
nand U14076 (N_14076,N_1865,N_1031);
or U14077 (N_14077,N_2198,N_9979);
and U14078 (N_14078,N_829,N_9583);
nor U14079 (N_14079,N_3891,N_4823);
nor U14080 (N_14080,N_1167,N_9130);
nand U14081 (N_14081,N_4734,N_8334);
and U14082 (N_14082,N_3240,N_945);
nand U14083 (N_14083,N_7414,N_5795);
xnor U14084 (N_14084,N_4209,N_9944);
nor U14085 (N_14085,N_6201,N_6647);
and U14086 (N_14086,N_9335,N_1214);
and U14087 (N_14087,N_9382,N_1986);
and U14088 (N_14088,N_8715,N_506);
nor U14089 (N_14089,N_4656,N_3165);
nor U14090 (N_14090,N_4578,N_6461);
and U14091 (N_14091,N_419,N_7529);
nand U14092 (N_14092,N_393,N_6017);
or U14093 (N_14093,N_3908,N_9946);
nand U14094 (N_14094,N_8522,N_381);
or U14095 (N_14095,N_3597,N_1670);
nand U14096 (N_14096,N_9439,N_9532);
nor U14097 (N_14097,N_2798,N_1571);
or U14098 (N_14098,N_8211,N_3647);
or U14099 (N_14099,N_35,N_3255);
and U14100 (N_14100,N_5302,N_584);
nor U14101 (N_14101,N_755,N_6077);
nor U14102 (N_14102,N_642,N_6917);
and U14103 (N_14103,N_6002,N_9945);
xnor U14104 (N_14104,N_1550,N_116);
and U14105 (N_14105,N_9277,N_6565);
nand U14106 (N_14106,N_5055,N_6124);
nor U14107 (N_14107,N_370,N_1860);
or U14108 (N_14108,N_8339,N_8836);
and U14109 (N_14109,N_9793,N_9498);
and U14110 (N_14110,N_9536,N_1177);
nor U14111 (N_14111,N_2726,N_4424);
nand U14112 (N_14112,N_459,N_1471);
xor U14113 (N_14113,N_4494,N_2592);
nor U14114 (N_14114,N_6919,N_8179);
nor U14115 (N_14115,N_2970,N_6412);
nor U14116 (N_14116,N_5555,N_4576);
nand U14117 (N_14117,N_8406,N_1490);
nand U14118 (N_14118,N_9466,N_859);
nor U14119 (N_14119,N_831,N_3954);
xor U14120 (N_14120,N_8015,N_4783);
or U14121 (N_14121,N_947,N_3875);
or U14122 (N_14122,N_9061,N_1569);
nand U14123 (N_14123,N_7421,N_3779);
nor U14124 (N_14124,N_6823,N_871);
nor U14125 (N_14125,N_5277,N_7942);
or U14126 (N_14126,N_4295,N_2701);
nand U14127 (N_14127,N_5951,N_2501);
and U14128 (N_14128,N_181,N_2415);
nand U14129 (N_14129,N_7843,N_221);
nand U14130 (N_14130,N_6132,N_6230);
or U14131 (N_14131,N_693,N_5110);
nand U14132 (N_14132,N_9018,N_7384);
nand U14133 (N_14133,N_4886,N_2476);
or U14134 (N_14134,N_1596,N_5389);
and U14135 (N_14135,N_6694,N_6473);
nand U14136 (N_14136,N_8167,N_8818);
or U14137 (N_14137,N_6898,N_3720);
and U14138 (N_14138,N_4186,N_6280);
or U14139 (N_14139,N_7987,N_4508);
nand U14140 (N_14140,N_2805,N_626);
nand U14141 (N_14141,N_8207,N_8612);
and U14142 (N_14142,N_8682,N_4447);
nor U14143 (N_14143,N_9724,N_4268);
nand U14144 (N_14144,N_6535,N_7375);
nand U14145 (N_14145,N_3134,N_3184);
nand U14146 (N_14146,N_1652,N_8796);
nor U14147 (N_14147,N_230,N_4504);
and U14148 (N_14148,N_2276,N_9048);
xor U14149 (N_14149,N_8482,N_1913);
and U14150 (N_14150,N_919,N_6523);
and U14151 (N_14151,N_9087,N_7067);
and U14152 (N_14152,N_2895,N_531);
nor U14153 (N_14153,N_8620,N_6113);
xor U14154 (N_14154,N_412,N_3754);
and U14155 (N_14155,N_4763,N_2179);
or U14156 (N_14156,N_8455,N_8843);
or U14157 (N_14157,N_5155,N_9249);
xor U14158 (N_14158,N_1685,N_1049);
and U14159 (N_14159,N_9168,N_6467);
and U14160 (N_14160,N_415,N_609);
and U14161 (N_14161,N_5088,N_6222);
nor U14162 (N_14162,N_4094,N_5153);
or U14163 (N_14163,N_6131,N_8025);
or U14164 (N_14164,N_3245,N_6371);
nand U14165 (N_14165,N_6987,N_4184);
nand U14166 (N_14166,N_9999,N_5317);
or U14167 (N_14167,N_6981,N_1100);
nor U14168 (N_14168,N_1734,N_7698);
nand U14169 (N_14169,N_440,N_6692);
nor U14170 (N_14170,N_1914,N_1616);
and U14171 (N_14171,N_1184,N_6391);
or U14172 (N_14172,N_5615,N_8138);
and U14173 (N_14173,N_5238,N_2604);
nand U14174 (N_14174,N_9485,N_9217);
nor U14175 (N_14175,N_1524,N_6929);
nand U14176 (N_14176,N_7859,N_3918);
or U14177 (N_14177,N_5661,N_422);
and U14178 (N_14178,N_2189,N_690);
and U14179 (N_14179,N_9521,N_9013);
nand U14180 (N_14180,N_3569,N_7548);
or U14181 (N_14181,N_9150,N_7498);
nand U14182 (N_14182,N_5600,N_5844);
nand U14183 (N_14183,N_5940,N_3562);
nand U14184 (N_14184,N_1394,N_1457);
xor U14185 (N_14185,N_5482,N_5441);
and U14186 (N_14186,N_8416,N_3345);
and U14187 (N_14187,N_529,N_6496);
or U14188 (N_14188,N_575,N_9329);
nor U14189 (N_14189,N_9504,N_3182);
nand U14190 (N_14190,N_233,N_6633);
nand U14191 (N_14191,N_2936,N_2018);
nand U14192 (N_14192,N_2419,N_8941);
nand U14193 (N_14193,N_8428,N_3443);
nand U14194 (N_14194,N_9342,N_3022);
xor U14195 (N_14195,N_9198,N_8312);
and U14196 (N_14196,N_6257,N_5763);
nand U14197 (N_14197,N_6104,N_3871);
nor U14198 (N_14198,N_6021,N_9817);
and U14199 (N_14199,N_236,N_9511);
and U14200 (N_14200,N_5966,N_8008);
nand U14201 (N_14201,N_5301,N_9939);
nor U14202 (N_14202,N_6293,N_2152);
and U14203 (N_14203,N_4242,N_188);
xor U14204 (N_14204,N_6735,N_7490);
and U14205 (N_14205,N_709,N_9983);
nor U14206 (N_14206,N_8578,N_2462);
nand U14207 (N_14207,N_3278,N_9769);
or U14208 (N_14208,N_7930,N_2932);
nand U14209 (N_14209,N_1367,N_4665);
xor U14210 (N_14210,N_3175,N_9550);
or U14211 (N_14211,N_7559,N_1432);
nor U14212 (N_14212,N_6102,N_3461);
nand U14213 (N_14213,N_3384,N_3081);
nand U14214 (N_14214,N_5990,N_9790);
nor U14215 (N_14215,N_8927,N_598);
or U14216 (N_14216,N_337,N_8702);
nand U14217 (N_14217,N_5006,N_9101);
nand U14218 (N_14218,N_6009,N_4715);
nor U14219 (N_14219,N_7890,N_4328);
nor U14220 (N_14220,N_3567,N_2433);
or U14221 (N_14221,N_41,N_6374);
nor U14222 (N_14222,N_3844,N_2702);
xor U14223 (N_14223,N_6007,N_4445);
or U14224 (N_14224,N_1940,N_3755);
or U14225 (N_14225,N_9650,N_8306);
nor U14226 (N_14226,N_6956,N_9732);
nand U14227 (N_14227,N_6808,N_9913);
or U14228 (N_14228,N_6092,N_936);
or U14229 (N_14229,N_2065,N_9728);
or U14230 (N_14230,N_7,N_7734);
or U14231 (N_14231,N_5536,N_6004);
xor U14232 (N_14232,N_4854,N_7580);
and U14233 (N_14233,N_8704,N_4673);
and U14234 (N_14234,N_545,N_6471);
and U14235 (N_14235,N_3815,N_2001);
and U14236 (N_14236,N_1006,N_5644);
and U14237 (N_14237,N_6070,N_8781);
or U14238 (N_14238,N_3621,N_3455);
xnor U14239 (N_14239,N_5253,N_9963);
and U14240 (N_14240,N_8901,N_8852);
nor U14241 (N_14241,N_275,N_2410);
nand U14242 (N_14242,N_863,N_3604);
nor U14243 (N_14243,N_4036,N_1762);
nand U14244 (N_14244,N_7684,N_4168);
xnor U14245 (N_14245,N_5985,N_8800);
nor U14246 (N_14246,N_3970,N_2020);
or U14247 (N_14247,N_5177,N_6298);
or U14248 (N_14248,N_7126,N_3130);
nand U14249 (N_14249,N_3996,N_9019);
and U14250 (N_14250,N_6609,N_5325);
nand U14251 (N_14251,N_396,N_2108);
nor U14252 (N_14252,N_4403,N_514);
xor U14253 (N_14253,N_9810,N_5347);
nor U14254 (N_14254,N_7855,N_9938);
nor U14255 (N_14255,N_6164,N_7348);
or U14256 (N_14256,N_8379,N_1077);
or U14257 (N_14257,N_679,N_3955);
and U14258 (N_14258,N_384,N_7972);
nand U14259 (N_14259,N_1264,N_8017);
and U14260 (N_14260,N_4470,N_2178);
nor U14261 (N_14261,N_4236,N_4851);
or U14262 (N_14262,N_8922,N_132);
or U14263 (N_14263,N_8759,N_4701);
xor U14264 (N_14264,N_311,N_7025);
nand U14265 (N_14265,N_7637,N_6579);
and U14266 (N_14266,N_2180,N_6988);
xnor U14267 (N_14267,N_3632,N_1681);
nand U14268 (N_14268,N_269,N_4645);
nand U14269 (N_14269,N_1564,N_4974);
or U14270 (N_14270,N_3370,N_8622);
nand U14271 (N_14271,N_6208,N_8144);
or U14272 (N_14272,N_5234,N_9450);
xnor U14273 (N_14273,N_4063,N_3437);
nand U14274 (N_14274,N_7336,N_173);
or U14275 (N_14275,N_7555,N_6806);
and U14276 (N_14276,N_4694,N_5124);
or U14277 (N_14277,N_7385,N_7455);
and U14278 (N_14278,N_4137,N_48);
nand U14279 (N_14279,N_1519,N_405);
and U14280 (N_14280,N_708,N_3103);
and U14281 (N_14281,N_5939,N_2506);
xor U14282 (N_14282,N_2962,N_3486);
or U14283 (N_14283,N_6870,N_7306);
xor U14284 (N_14284,N_5035,N_3191);
nor U14285 (N_14285,N_3928,N_2585);
nor U14286 (N_14286,N_6235,N_5396);
nand U14287 (N_14287,N_7611,N_5241);
or U14288 (N_14288,N_3339,N_3582);
and U14289 (N_14289,N_9702,N_1636);
nand U14290 (N_14290,N_2278,N_599);
or U14291 (N_14291,N_5733,N_5280);
or U14292 (N_14292,N_3883,N_6025);
nand U14293 (N_14293,N_5575,N_5071);
xnor U14294 (N_14294,N_5351,N_784);
xnor U14295 (N_14295,N_36,N_2945);
xnor U14296 (N_14296,N_7520,N_637);
nor U14297 (N_14297,N_790,N_8407);
and U14298 (N_14298,N_3067,N_1480);
nor U14299 (N_14299,N_4653,N_589);
and U14300 (N_14300,N_6097,N_2246);
and U14301 (N_14301,N_8403,N_2967);
nand U14302 (N_14302,N_5822,N_5909);
nand U14303 (N_14303,N_30,N_7358);
or U14304 (N_14304,N_7058,N_1827);
nand U14305 (N_14305,N_7094,N_3522);
nor U14306 (N_14306,N_1201,N_8773);
or U14307 (N_14307,N_7550,N_819);
and U14308 (N_14308,N_8546,N_5058);
nand U14309 (N_14309,N_4181,N_8813);
nor U14310 (N_14310,N_1781,N_4346);
xnor U14311 (N_14311,N_6108,N_1624);
or U14312 (N_14312,N_7011,N_2488);
xor U14313 (N_14313,N_2070,N_1612);
nor U14314 (N_14314,N_9283,N_126);
and U14315 (N_14315,N_6681,N_9628);
or U14316 (N_14316,N_7317,N_3341);
nor U14317 (N_14317,N_2833,N_6205);
nor U14318 (N_14318,N_509,N_6368);
nand U14319 (N_14319,N_8152,N_8710);
nor U14320 (N_14320,N_1278,N_6340);
or U14321 (N_14321,N_3658,N_3535);
xor U14322 (N_14322,N_1822,N_2685);
nor U14323 (N_14323,N_9672,N_1980);
and U14324 (N_14324,N_5682,N_6656);
nor U14325 (N_14325,N_5831,N_4940);
nor U14326 (N_14326,N_43,N_1081);
or U14327 (N_14327,N_3033,N_3590);
or U14328 (N_14328,N_7187,N_8018);
or U14329 (N_14329,N_3094,N_9497);
and U14330 (N_14330,N_7982,N_7059);
and U14331 (N_14331,N_4199,N_4841);
and U14332 (N_14332,N_9634,N_5773);
nand U14333 (N_14333,N_8739,N_920);
or U14334 (N_14334,N_2982,N_5911);
or U14335 (N_14335,N_2873,N_4320);
and U14336 (N_14336,N_82,N_8305);
xor U14337 (N_14337,N_1658,N_3166);
and U14338 (N_14338,N_3304,N_7678);
and U14339 (N_14339,N_385,N_7599);
xor U14340 (N_14340,N_7712,N_3095);
nor U14341 (N_14341,N_1692,N_6341);
nand U14342 (N_14342,N_2781,N_5108);
or U14343 (N_14343,N_3740,N_5397);
nand U14344 (N_14344,N_5048,N_2406);
nand U14345 (N_14345,N_6281,N_5250);
or U14346 (N_14346,N_4189,N_5015);
or U14347 (N_14347,N_8224,N_7315);
and U14348 (N_14348,N_6768,N_3784);
nor U14349 (N_14349,N_948,N_5144);
and U14350 (N_14350,N_3411,N_3325);
xnor U14351 (N_14351,N_5199,N_4476);
or U14352 (N_14352,N_1207,N_7857);
or U14353 (N_14353,N_3743,N_8848);
or U14354 (N_14354,N_1678,N_4755);
or U14355 (N_14355,N_6055,N_280);
and U14356 (N_14356,N_8936,N_1274);
nor U14357 (N_14357,N_750,N_4075);
nand U14358 (N_14358,N_3983,N_4159);
xor U14359 (N_14359,N_8069,N_9132);
and U14360 (N_14360,N_1256,N_1124);
nand U14361 (N_14361,N_2693,N_5957);
or U14362 (N_14362,N_6305,N_9356);
xor U14363 (N_14363,N_4053,N_4767);
or U14364 (N_14364,N_108,N_542);
and U14365 (N_14365,N_1287,N_6947);
or U14366 (N_14366,N_8159,N_7009);
nand U14367 (N_14367,N_1837,N_7383);
and U14368 (N_14368,N_1623,N_5635);
nand U14369 (N_14369,N_4188,N_5298);
or U14370 (N_14370,N_8748,N_4297);
xor U14371 (N_14371,N_7408,N_4345);
nor U14372 (N_14372,N_3607,N_137);
nand U14373 (N_14373,N_2643,N_2810);
nor U14374 (N_14374,N_9,N_1643);
and U14375 (N_14375,N_880,N_2547);
nor U14376 (N_14376,N_1180,N_2470);
nand U14377 (N_14377,N_7349,N_4581);
and U14378 (N_14378,N_411,N_5457);
nor U14379 (N_14379,N_8472,N_5413);
or U14380 (N_14380,N_3664,N_9858);
nor U14381 (N_14381,N_8625,N_9752);
nor U14382 (N_14382,N_8280,N_5312);
nand U14383 (N_14383,N_5184,N_9173);
or U14384 (N_14384,N_9377,N_3149);
or U14385 (N_14385,N_7156,N_1764);
nand U14386 (N_14386,N_8484,N_932);
xnor U14387 (N_14387,N_6081,N_9040);
nand U14388 (N_14388,N_8830,N_9068);
nor U14389 (N_14389,N_1231,N_2587);
nor U14390 (N_14390,N_90,N_7105);
nand U14391 (N_14391,N_5678,N_7733);
xnor U14392 (N_14392,N_9352,N_1630);
and U14393 (N_14393,N_6740,N_6350);
xor U14394 (N_14394,N_9782,N_6914);
or U14395 (N_14395,N_3047,N_4497);
and U14396 (N_14396,N_7759,N_9392);
and U14397 (N_14397,N_5480,N_6907);
xnor U14398 (N_14398,N_7447,N_3353);
nand U14399 (N_14399,N_4856,N_9966);
and U14400 (N_14400,N_5026,N_3571);
nor U14401 (N_14401,N_8336,N_8542);
nor U14402 (N_14402,N_5802,N_4344);
or U14403 (N_14403,N_2754,N_6596);
and U14404 (N_14404,N_1276,N_1395);
and U14405 (N_14405,N_3210,N_7677);
and U14406 (N_14406,N_9816,N_6291);
and U14407 (N_14407,N_821,N_4956);
and U14408 (N_14408,N_7240,N_305);
nand U14409 (N_14409,N_8889,N_6606);
nand U14410 (N_14410,N_9160,N_7629);
nand U14411 (N_14411,N_8523,N_9582);
xor U14412 (N_14412,N_5589,N_1691);
nor U14413 (N_14413,N_4738,N_2513);
xnor U14414 (N_14414,N_4939,N_5062);
nand U14415 (N_14415,N_2502,N_7867);
and U14416 (N_14416,N_3030,N_4791);
and U14417 (N_14417,N_5868,N_8198);
and U14418 (N_14418,N_1262,N_5636);
or U14419 (N_14419,N_1311,N_4057);
xor U14420 (N_14420,N_8184,N_28);
nor U14421 (N_14421,N_2942,N_5893);
or U14422 (N_14422,N_1962,N_7920);
nand U14423 (N_14423,N_2976,N_4915);
and U14424 (N_14424,N_2370,N_420);
nor U14425 (N_14425,N_7648,N_5852);
nor U14426 (N_14426,N_553,N_3895);
and U14427 (N_14427,N_2551,N_8360);
and U14428 (N_14428,N_4353,N_5114);
or U14429 (N_14429,N_1269,N_4925);
or U14430 (N_14430,N_2708,N_9855);
nand U14431 (N_14431,N_9070,N_2477);
xor U14432 (N_14432,N_3680,N_3421);
or U14433 (N_14433,N_7514,N_8590);
or U14434 (N_14434,N_3708,N_6777);
and U14435 (N_14435,N_7691,N_3289);
and U14436 (N_14436,N_4762,N_5925);
and U14437 (N_14437,N_5732,N_1555);
and U14438 (N_14438,N_3402,N_5609);
xor U14439 (N_14439,N_7283,N_1390);
xnor U14440 (N_14440,N_9674,N_4317);
and U14441 (N_14441,N_9621,N_744);
nand U14442 (N_14442,N_1640,N_9370);
nor U14443 (N_14443,N_8188,N_3910);
nand U14444 (N_14444,N_4711,N_3514);
or U14445 (N_14445,N_329,N_2319);
or U14446 (N_14446,N_1725,N_2162);
nand U14447 (N_14447,N_46,N_6187);
nor U14448 (N_14448,N_8765,N_2973);
nor U14449 (N_14449,N_1294,N_7716);
nand U14450 (N_14450,N_9246,N_3505);
nand U14451 (N_14451,N_1821,N_604);
nand U14452 (N_14452,N_6613,N_291);
nand U14453 (N_14453,N_7519,N_3633);
nor U14454 (N_14454,N_4203,N_6270);
or U14455 (N_14455,N_1528,N_4397);
xnor U14456 (N_14456,N_1115,N_8680);
or U14457 (N_14457,N_5596,N_3179);
or U14458 (N_14458,N_6957,N_6357);
nor U14459 (N_14459,N_4857,N_3596);
and U14460 (N_14460,N_8719,N_9163);
and U14461 (N_14461,N_3008,N_2519);
nor U14462 (N_14462,N_8694,N_7406);
and U14463 (N_14463,N_3369,N_2565);
xnor U14464 (N_14464,N_7870,N_806);
nand U14465 (N_14465,N_5150,N_3613);
xor U14466 (N_14466,N_4708,N_6262);
and U14467 (N_14467,N_2812,N_3342);
or U14468 (N_14468,N_2023,N_3379);
and U14469 (N_14469,N_9340,N_1097);
and U14470 (N_14470,N_2397,N_7229);
or U14471 (N_14471,N_4626,N_4272);
nand U14472 (N_14472,N_2898,N_2559);
or U14473 (N_14473,N_1816,N_4853);
nor U14474 (N_14474,N_2486,N_9753);
or U14475 (N_14475,N_5853,N_5310);
nand U14476 (N_14476,N_7043,N_725);
and U14477 (N_14477,N_3909,N_617);
and U14478 (N_14478,N_3667,N_2084);
nor U14479 (N_14479,N_5816,N_4794);
or U14480 (N_14480,N_8153,N_8319);
nor U14481 (N_14481,N_5704,N_4599);
nand U14482 (N_14482,N_4444,N_1613);
and U14483 (N_14483,N_2737,N_7706);
nor U14484 (N_14484,N_3943,N_6676);
nand U14485 (N_14485,N_4568,N_2892);
nand U14486 (N_14486,N_3311,N_6706);
nand U14487 (N_14487,N_1838,N_349);
or U14488 (N_14488,N_9892,N_8648);
and U14489 (N_14489,N_6915,N_1249);
nor U14490 (N_14490,N_4522,N_8776);
nand U14491 (N_14491,N_2244,N_8814);
nand U14492 (N_14492,N_7671,N_3258);
nor U14493 (N_14493,N_7607,N_6547);
nor U14494 (N_14494,N_881,N_935);
nor U14495 (N_14495,N_8131,N_1877);
or U14496 (N_14496,N_2361,N_5157);
nor U14497 (N_14497,N_6620,N_8363);
nand U14498 (N_14498,N_1873,N_8246);
nor U14499 (N_14499,N_2676,N_4914);
nand U14500 (N_14500,N_7909,N_5258);
and U14501 (N_14501,N_75,N_1086);
and U14502 (N_14502,N_5935,N_208);
nand U14503 (N_14503,N_4310,N_5748);
xnor U14504 (N_14504,N_7709,N_15);
xor U14505 (N_14505,N_77,N_7665);
nand U14506 (N_14506,N_5162,N_5113);
xnor U14507 (N_14507,N_5205,N_6236);
nor U14508 (N_14508,N_9864,N_4641);
or U14509 (N_14509,N_1711,N_3123);
or U14510 (N_14510,N_9784,N_44);
or U14511 (N_14511,N_3016,N_7326);
and U14512 (N_14512,N_5414,N_397);
xor U14513 (N_14513,N_400,N_4548);
or U14514 (N_14514,N_4775,N_566);
or U14515 (N_14515,N_3260,N_3004);
nor U14516 (N_14516,N_4662,N_5147);
xnor U14517 (N_14517,N_4490,N_8960);
or U14518 (N_14518,N_5639,N_939);
nand U14519 (N_14519,N_371,N_1889);
xor U14520 (N_14520,N_1964,N_2002);
and U14521 (N_14521,N_68,N_3354);
or U14522 (N_14522,N_1592,N_3946);
and U14523 (N_14523,N_5186,N_6977);
nand U14524 (N_14524,N_2848,N_827);
nor U14525 (N_14525,N_861,N_3365);
xor U14526 (N_14526,N_9119,N_8388);
and U14527 (N_14527,N_9374,N_8028);
and U14528 (N_14528,N_3751,N_4405);
nand U14529 (N_14529,N_6839,N_1586);
nand U14530 (N_14530,N_9296,N_1941);
and U14531 (N_14531,N_5028,N_6211);
and U14532 (N_14532,N_8313,N_9585);
xor U14533 (N_14533,N_3,N_7320);
nand U14534 (N_14534,N_445,N_5271);
and U14535 (N_14535,N_1090,N_7001);
nand U14536 (N_14536,N_9468,N_8404);
and U14537 (N_14537,N_5274,N_5886);
nor U14538 (N_14538,N_3724,N_5170);
or U14539 (N_14539,N_1337,N_1785);
or U14540 (N_14540,N_9626,N_3297);
and U14541 (N_14541,N_8775,N_3469);
nand U14542 (N_14542,N_6696,N_7897);
or U14543 (N_14543,N_9574,N_9331);
and U14544 (N_14544,N_3549,N_4301);
or U14545 (N_14545,N_141,N_340);
nor U14546 (N_14546,N_2842,N_1259);
and U14547 (N_14547,N_5183,N_911);
nand U14548 (N_14548,N_2098,N_7834);
nor U14549 (N_14549,N_780,N_9873);
nor U14550 (N_14550,N_6720,N_2097);
or U14551 (N_14551,N_3000,N_3594);
nand U14552 (N_14552,N_4247,N_4323);
and U14553 (N_14553,N_3143,N_2856);
or U14554 (N_14554,N_2272,N_7693);
or U14555 (N_14555,N_524,N_3550);
nand U14556 (N_14556,N_4909,N_5616);
and U14557 (N_14557,N_9818,N_9618);
nand U14558 (N_14558,N_5513,N_277);
or U14559 (N_14559,N_934,N_3984);
or U14560 (N_14560,N_5448,N_5120);
or U14561 (N_14561,N_4719,N_8707);
or U14562 (N_14562,N_3473,N_9478);
or U14563 (N_14563,N_5466,N_9640);
or U14564 (N_14564,N_6285,N_6903);
and U14565 (N_14565,N_9323,N_7586);
or U14566 (N_14566,N_6184,N_6497);
and U14567 (N_14567,N_7591,N_5524);
nand U14568 (N_14568,N_5562,N_797);
and U14569 (N_14569,N_6260,N_9383);
nor U14570 (N_14570,N_3881,N_7563);
or U14571 (N_14571,N_4664,N_3715);
nor U14572 (N_14572,N_2059,N_7333);
or U14573 (N_14573,N_1020,N_8046);
nor U14574 (N_14574,N_6763,N_9469);
and U14575 (N_14575,N_9349,N_3111);
nor U14576 (N_14576,N_8992,N_5281);
nand U14577 (N_14577,N_7943,N_7028);
and U14578 (N_14578,N_4226,N_7190);
or U14579 (N_14579,N_9029,N_60);
nor U14580 (N_14580,N_2448,N_1458);
nor U14581 (N_14581,N_7055,N_5021);
or U14582 (N_14582,N_9889,N_4919);
or U14583 (N_14583,N_4745,N_2746);
and U14584 (N_14584,N_6197,N_1598);
nand U14585 (N_14585,N_7849,N_1504);
nor U14586 (N_14586,N_6151,N_8746);
or U14587 (N_14587,N_5076,N_8321);
xnor U14588 (N_14588,N_7674,N_2306);
nor U14589 (N_14589,N_2430,N_3950);
xnor U14590 (N_14590,N_6086,N_4194);
xnor U14591 (N_14591,N_6651,N_5072);
or U14592 (N_14592,N_448,N_5094);
and U14593 (N_14593,N_3070,N_5722);
and U14594 (N_14594,N_1672,N_9441);
nand U14595 (N_14595,N_4997,N_9652);
and U14596 (N_14596,N_6863,N_8441);
or U14597 (N_14597,N_869,N_6759);
nor U14598 (N_14598,N_6809,N_3778);
nand U14599 (N_14599,N_5096,N_4814);
or U14600 (N_14600,N_7007,N_2727);
nor U14601 (N_14601,N_6079,N_5845);
nand U14602 (N_14602,N_2610,N_908);
and U14603 (N_14603,N_1783,N_9956);
nor U14604 (N_14604,N_9049,N_5525);
nor U14605 (N_14605,N_1444,N_5987);
xnor U14606 (N_14606,N_4501,N_2534);
nand U14607 (N_14607,N_6398,N_7787);
and U14608 (N_14608,N_8343,N_7579);
nand U14609 (N_14609,N_1649,N_6169);
or U14610 (N_14610,N_7335,N_4417);
nand U14611 (N_14611,N_4233,N_1183);
nand U14612 (N_14612,N_4777,N_1788);
nand U14613 (N_14613,N_3364,N_8254);
or U14614 (N_14614,N_4408,N_9462);
xnor U14615 (N_14615,N_1443,N_5243);
and U14616 (N_14616,N_3854,N_5487);
xnor U14617 (N_14617,N_9255,N_1539);
nor U14618 (N_14618,N_1163,N_298);
or U14619 (N_14619,N_4112,N_4111);
nand U14620 (N_14620,N_6950,N_5208);
nand U14621 (N_14621,N_9595,N_6163);
xor U14622 (N_14622,N_5950,N_4824);
nand U14623 (N_14623,N_4371,N_2977);
and U14624 (N_14624,N_13,N_6196);
and U14625 (N_14625,N_3538,N_2342);
nand U14626 (N_14626,N_6016,N_6822);
or U14627 (N_14627,N_1075,N_9093);
nand U14628 (N_14628,N_2356,N_9786);
or U14629 (N_14629,N_8559,N_3292);
or U14630 (N_14630,N_8632,N_6954);
nor U14631 (N_14631,N_6590,N_2265);
nor U14632 (N_14632,N_8811,N_3638);
or U14633 (N_14633,N_4714,N_4141);
or U14634 (N_14634,N_3087,N_4818);
nor U14635 (N_14635,N_1663,N_660);
xnor U14636 (N_14636,N_5416,N_1800);
or U14637 (N_14637,N_9940,N_7223);
or U14638 (N_14638,N_8624,N_6576);
nand U14639 (N_14639,N_6121,N_9625);
or U14640 (N_14640,N_9743,N_8832);
or U14641 (N_14641,N_3822,N_9135);
nand U14642 (N_14642,N_9811,N_8440);
nand U14643 (N_14643,N_7339,N_1974);
or U14644 (N_14644,N_7713,N_3763);
nand U14645 (N_14645,N_2399,N_4406);
or U14646 (N_14646,N_9502,N_286);
nand U14647 (N_14647,N_1448,N_1341);
nor U14648 (N_14648,N_1554,N_310);
xor U14649 (N_14649,N_9142,N_4351);
and U14650 (N_14650,N_2729,N_732);
and U14651 (N_14651,N_9622,N_1194);
nand U14652 (N_14652,N_2664,N_274);
and U14653 (N_14653,N_127,N_5625);
nor U14654 (N_14654,N_5115,N_7485);
nor U14655 (N_14655,N_2035,N_387);
nor U14656 (N_14656,N_3941,N_9984);
nor U14657 (N_14657,N_4270,N_3848);
nand U14658 (N_14658,N_5227,N_7044);
and U14659 (N_14659,N_7090,N_1635);
xnor U14660 (N_14660,N_8314,N_3368);
or U14661 (N_14661,N_6718,N_6503);
nor U14662 (N_14662,N_5633,N_9673);
or U14663 (N_14663,N_9964,N_8987);
nand U14664 (N_14664,N_2380,N_1154);
nand U14665 (N_14665,N_811,N_9969);
nor U14666 (N_14666,N_9042,N_1522);
or U14667 (N_14667,N_5598,N_7710);
nand U14668 (N_14668,N_8447,N_2631);
nor U14669 (N_14669,N_8408,N_3600);
xor U14670 (N_14670,N_2390,N_2457);
nor U14671 (N_14671,N_8591,N_8827);
xnor U14672 (N_14672,N_2778,N_3581);
or U14673 (N_14673,N_6465,N_818);
and U14674 (N_14674,N_6868,N_7505);
nand U14675 (N_14675,N_5087,N_6144);
or U14676 (N_14676,N_8106,N_7858);
or U14677 (N_14677,N_4564,N_3006);
nand U14678 (N_14678,N_1403,N_3957);
xnor U14679 (N_14679,N_3563,N_6600);
and U14680 (N_14680,N_5267,N_331);
or U14681 (N_14681,N_3830,N_6626);
or U14682 (N_14682,N_4022,N_9380);
nor U14683 (N_14683,N_4361,N_5516);
nand U14684 (N_14684,N_234,N_2563);
nand U14685 (N_14685,N_4054,N_8072);
nor U14686 (N_14686,N_4529,N_8177);
and U14687 (N_14687,N_7082,N_8232);
and U14688 (N_14688,N_6815,N_4718);
or U14689 (N_14689,N_9919,N_6946);
xnor U14690 (N_14690,N_9563,N_4015);
or U14691 (N_14691,N_4942,N_1676);
or U14692 (N_14692,N_6228,N_4999);
nor U14693 (N_14693,N_5504,N_4964);
nor U14694 (N_14694,N_6089,N_7888);
nor U14695 (N_14695,N_1582,N_8027);
and U14696 (N_14696,N_9367,N_479);
and U14697 (N_14697,N_941,N_2897);
nor U14698 (N_14698,N_3466,N_3024);
and U14699 (N_14699,N_6195,N_4754);
and U14700 (N_14700,N_7450,N_3347);
nor U14701 (N_14701,N_6134,N_8364);
nor U14702 (N_14702,N_2831,N_4782);
and U14703 (N_14703,N_2653,N_4880);
nor U14704 (N_14704,N_8043,N_8013);
or U14705 (N_14705,N_5867,N_4601);
nor U14706 (N_14706,N_9510,N_7517);
and U14707 (N_14707,N_9927,N_899);
and U14708 (N_14708,N_390,N_4409);
nor U14709 (N_14709,N_9402,N_255);
and U14710 (N_14710,N_601,N_1722);
and U14711 (N_14711,N_3985,N_2219);
nor U14712 (N_14712,N_2951,N_9376);
nor U14713 (N_14713,N_7031,N_3729);
or U14714 (N_14714,N_8736,N_8875);
and U14715 (N_14715,N_8450,N_8464);
or U14716 (N_14716,N_6029,N_8079);
or U14717 (N_14717,N_9378,N_6664);
xor U14718 (N_14718,N_7737,N_2837);
and U14719 (N_14719,N_4861,N_8166);
or U14720 (N_14720,N_6103,N_9422);
nor U14721 (N_14721,N_3493,N_2450);
and U14722 (N_14722,N_6866,N_4350);
nand U14723 (N_14723,N_9179,N_1938);
and U14724 (N_14724,N_6642,N_2487);
xnor U14725 (N_14725,N_4090,N_2261);
xor U14726 (N_14726,N_7076,N_5762);
or U14727 (N_14727,N_6812,N_6353);
nor U14728 (N_14728,N_6161,N_205);
nor U14729 (N_14729,N_3829,N_8561);
xnor U14730 (N_14730,N_2562,N_3205);
nand U14731 (N_14731,N_1244,N_2688);
nand U14732 (N_14732,N_8125,N_4146);
and U14733 (N_14733,N_1474,N_67);
nor U14734 (N_14734,N_1038,N_1895);
and U14735 (N_14735,N_9548,N_4302);
and U14736 (N_14736,N_8193,N_418);
xnor U14737 (N_14737,N_8849,N_1083);
and U14738 (N_14738,N_2388,N_2452);
nor U14739 (N_14739,N_9560,N_2692);
and U14740 (N_14740,N_1492,N_3451);
or U14741 (N_14741,N_1455,N_9071);
nor U14742 (N_14742,N_7605,N_4521);
or U14743 (N_14743,N_5758,N_3489);
and U14744 (N_14744,N_5634,N_5299);
and U14745 (N_14745,N_7965,N_1748);
nand U14746 (N_14746,N_3271,N_2971);
nand U14747 (N_14747,N_9355,N_4602);
xor U14748 (N_14748,N_9118,N_9624);
nand U14749 (N_14749,N_8446,N_4116);
nand U14750 (N_14750,N_7816,N_7721);
or U14751 (N_14751,N_1387,N_2912);
and U14752 (N_14752,N_9341,N_2651);
nor U14753 (N_14753,N_8853,N_4352);
nand U14754 (N_14754,N_8156,N_2890);
nor U14755 (N_14755,N_3174,N_9014);
and U14756 (N_14756,N_386,N_7325);
or U14757 (N_14757,N_9012,N_8080);
and U14758 (N_14758,N_989,N_474);
nor U14759 (N_14759,N_2311,N_1108);
nand U14760 (N_14760,N_4000,N_3705);
or U14761 (N_14761,N_3419,N_4109);
nand U14762 (N_14762,N_2821,N_4033);
nand U14763 (N_14763,N_6801,N_3453);
nand U14764 (N_14764,N_5709,N_3837);
nand U14765 (N_14765,N_2561,N_6844);
or U14766 (N_14766,N_9714,N_2205);
nand U14767 (N_14767,N_7367,N_433);
nor U14768 (N_14768,N_4700,N_5899);
nand U14769 (N_14769,N_17,N_4426);
nor U14770 (N_14770,N_3168,N_3214);
nor U14771 (N_14771,N_1752,N_8176);
and U14772 (N_14772,N_8965,N_3424);
and U14773 (N_14773,N_5801,N_2740);
nor U14774 (N_14774,N_9304,N_3625);
nor U14775 (N_14775,N_1795,N_8855);
and U14776 (N_14776,N_3157,N_6488);
xnor U14777 (N_14777,N_3426,N_1869);
or U14778 (N_14778,N_5730,N_7429);
or U14779 (N_14779,N_6660,N_8476);
nand U14780 (N_14780,N_6601,N_515);
nor U14781 (N_14781,N_2742,N_6359);
or U14782 (N_14782,N_5849,N_9870);
and U14783 (N_14783,N_9838,N_3601);
nor U14784 (N_14784,N_6495,N_5766);
nand U14785 (N_14785,N_7923,N_846);
nor U14786 (N_14786,N_7549,N_6346);
nor U14787 (N_14787,N_6562,N_9285);
nand U14788 (N_14788,N_1283,N_9152);
nand U14789 (N_14789,N_3502,N_5085);
nor U14790 (N_14790,N_7877,N_3282);
and U14791 (N_14791,N_1951,N_1862);
or U14792 (N_14792,N_8555,N_3874);
and U14793 (N_14793,N_2555,N_8740);
nor U14794 (N_14794,N_700,N_9736);
nor U14795 (N_14795,N_9975,N_6568);
or U14796 (N_14796,N_962,N_7700);
nand U14797 (N_14797,N_9052,N_6648);
or U14798 (N_14798,N_8213,N_4356);
nor U14799 (N_14799,N_8606,N_4030);
and U14800 (N_14800,N_8510,N_4496);
xor U14801 (N_14801,N_9926,N_1268);
or U14802 (N_14802,N_115,N_9800);
xor U14803 (N_14803,N_6998,N_7701);
nand U14804 (N_14804,N_2145,N_7921);
xor U14805 (N_14805,N_1411,N_8492);
and U14806 (N_14806,N_1650,N_5793);
nand U14807 (N_14807,N_4597,N_1150);
nand U14808 (N_14808,N_192,N_6566);
and U14809 (N_14809,N_6635,N_6378);
xor U14810 (N_14810,N_3435,N_7056);
nor U14811 (N_14811,N_4388,N_5131);
and U14812 (N_14812,N_6932,N_7441);
or U14813 (N_14813,N_2709,N_9177);
nand U14814 (N_14814,N_9954,N_7074);
or U14815 (N_14815,N_3927,N_191);
nand U14816 (N_14816,N_6519,N_717);
and U14817 (N_14817,N_8891,N_5323);
or U14818 (N_14818,N_9572,N_6068);
xor U14819 (N_14819,N_8757,N_2938);
nand U14820 (N_14820,N_2885,N_7892);
nand U14821 (N_14821,N_5104,N_9384);
or U14822 (N_14822,N_7840,N_959);
and U14823 (N_14823,N_7570,N_3570);
and U14824 (N_14824,N_6940,N_6991);
nand U14825 (N_14825,N_8180,N_9928);
or U14826 (N_14826,N_2816,N_9313);
or U14827 (N_14827,N_2745,N_788);
nor U14828 (N_14828,N_5649,N_4742);
nand U14829 (N_14829,N_6136,N_530);
or U14830 (N_14830,N_66,N_6934);
or U14831 (N_14831,N_3262,N_9221);
or U14832 (N_14832,N_4027,N_3266);
and U14833 (N_14833,N_3319,N_8361);
nand U14834 (N_14834,N_5977,N_1901);
or U14835 (N_14835,N_3843,N_7596);
nor U14836 (N_14836,N_8497,N_9726);
nor U14837 (N_14837,N_4996,N_2794);
xor U14838 (N_14838,N_754,N_6044);
or U14839 (N_14839,N_5024,N_8637);
and U14840 (N_14840,N_5941,N_7251);
or U14841 (N_14841,N_88,N_4505);
and U14842 (N_14842,N_2076,N_874);
nor U14843 (N_14843,N_6677,N_5602);
or U14844 (N_14844,N_6830,N_168);
and U14845 (N_14845,N_5231,N_1634);
nor U14846 (N_14846,N_477,N_8011);
xnor U14847 (N_14847,N_6843,N_4655);
nor U14848 (N_14848,N_97,N_9922);
or U14849 (N_14849,N_6328,N_8385);
nor U14850 (N_14850,N_4500,N_9917);
nand U14851 (N_14851,N_1918,N_1447);
nor U14852 (N_14852,N_5029,N_2773);
and U14853 (N_14853,N_9792,N_3938);
nor U14854 (N_14854,N_4487,N_5460);
nor U14855 (N_14855,N_1292,N_6910);
nand U14856 (N_14856,N_6895,N_1743);
or U14857 (N_14857,N_9045,N_3542);
nor U14858 (N_14858,N_5027,N_5159);
or U14859 (N_14859,N_4375,N_6920);
nor U14860 (N_14860,N_7202,N_1427);
or U14861 (N_14861,N_3574,N_1112);
or U14862 (N_14862,N_4994,N_6820);
nand U14863 (N_14863,N_470,N_9952);
and U14864 (N_14864,N_8174,N_2625);
and U14865 (N_14865,N_263,N_1699);
nand U14866 (N_14866,N_9457,N_2160);
nor U14867 (N_14867,N_3863,N_2238);
nor U14868 (N_14868,N_4959,N_6834);
xor U14869 (N_14869,N_2091,N_8462);
or U14870 (N_14870,N_3376,N_3678);
nand U14871 (N_14871,N_83,N_5092);
xor U14872 (N_14872,N_9832,N_1814);
and U14873 (N_14873,N_4970,N_5811);
nor U14874 (N_14874,N_7662,N_7644);
or U14875 (N_14875,N_9841,N_3427);
and U14876 (N_14876,N_4858,N_9893);
xnor U14877 (N_14877,N_4617,N_8900);
or U14878 (N_14878,N_85,N_3917);
xnor U14879 (N_14879,N_5543,N_3977);
nor U14880 (N_14880,N_6781,N_703);
or U14881 (N_14881,N_4217,N_6994);
or U14882 (N_14882,N_7378,N_1312);
and U14883 (N_14883,N_5712,N_434);
nand U14884 (N_14884,N_6758,N_5139);
and U14885 (N_14885,N_3598,N_622);
nand U14886 (N_14886,N_5311,N_3906);
and U14887 (N_14887,N_4802,N_8859);
nand U14888 (N_14888,N_7841,N_8171);
nor U14889 (N_14889,N_2903,N_4772);
nor U14890 (N_14890,N_5436,N_3056);
nor U14891 (N_14891,N_3480,N_9716);
or U14892 (N_14892,N_1756,N_5832);
or U14893 (N_14893,N_616,N_49);
and U14894 (N_14894,N_5248,N_9424);
or U14895 (N_14895,N_1050,N_3071);
and U14896 (N_14896,N_4670,N_3063);
or U14897 (N_14897,N_6292,N_1979);
or U14898 (N_14898,N_3762,N_635);
or U14899 (N_14899,N_4570,N_425);
nand U14900 (N_14900,N_5107,N_961);
xor U14901 (N_14901,N_6585,N_262);
and U14902 (N_14902,N_607,N_7818);
and U14903 (N_14903,N_4862,N_2389);
and U14904 (N_14904,N_5752,N_8626);
nor U14905 (N_14905,N_3250,N_1378);
and U14906 (N_14906,N_8540,N_7371);
nand U14907 (N_14907,N_1042,N_244);
nor U14908 (N_14908,N_195,N_2266);
xor U14909 (N_14909,N_5327,N_884);
nor U14910 (N_14910,N_8139,N_1686);
or U14911 (N_14911,N_4541,N_3189);
nor U14912 (N_14912,N_9643,N_4946);
and U14913 (N_14913,N_8515,N_6507);
xnor U14914 (N_14914,N_9820,N_9473);
nand U14915 (N_14915,N_6174,N_8318);
or U14916 (N_14916,N_1164,N_9448);
and U14917 (N_14917,N_7217,N_8508);
and U14918 (N_14918,N_6110,N_5003);
and U14919 (N_14919,N_8554,N_5962);
nor U14920 (N_14920,N_4093,N_1810);
or U14921 (N_14921,N_2793,N_805);
and U14922 (N_14922,N_8543,N_4575);
and U14923 (N_14923,N_1463,N_6277);
nor U14924 (N_14924,N_1983,N_5690);
nand U14925 (N_14925,N_7851,N_7808);
nor U14926 (N_14926,N_569,N_4277);
and U14927 (N_14927,N_450,N_5407);
xor U14928 (N_14928,N_774,N_7720);
xor U14929 (N_14929,N_2677,N_7249);
xor U14930 (N_14930,N_7746,N_8269);
and U14931 (N_14931,N_866,N_3586);
xor U14932 (N_14932,N_7742,N_4322);
and U14933 (N_14933,N_463,N_7572);
and U14934 (N_14934,N_3171,N_5134);
nand U14935 (N_14935,N_446,N_758);
nor U14936 (N_14936,N_171,N_8751);
nand U14937 (N_14937,N_5051,N_5079);
and U14938 (N_14938,N_4224,N_2309);
or U14939 (N_14939,N_1104,N_9735);
nor U14940 (N_14940,N_8558,N_6215);
or U14941 (N_14941,N_9188,N_1304);
nor U14942 (N_14942,N_8825,N_2505);
xnor U14943 (N_14943,N_7680,N_2412);
and U14944 (N_14944,N_511,N_4462);
or U14945 (N_14945,N_1257,N_5809);
and U14946 (N_14946,N_2408,N_442);
nor U14947 (N_14947,N_1247,N_2480);
and U14948 (N_14948,N_7655,N_3503);
nor U14949 (N_14949,N_120,N_1730);
and U14950 (N_14950,N_4144,N_9232);
and U14951 (N_14951,N_5786,N_7195);
nor U14952 (N_14952,N_2199,N_4439);
xnor U14953 (N_14953,N_8823,N_6715);
and U14954 (N_14954,N_2354,N_2595);
nor U14955 (N_14955,N_7003,N_9169);
and U14956 (N_14956,N_5213,N_8479);
and U14957 (N_14957,N_623,N_1753);
and U14958 (N_14958,N_9608,N_9187);
nor U14959 (N_14959,N_1977,N_2372);
xor U14960 (N_14960,N_2248,N_1852);
nor U14961 (N_14961,N_5201,N_3151);
nand U14962 (N_14962,N_6464,N_3866);
or U14963 (N_14963,N_3812,N_4096);
and U14964 (N_14964,N_4253,N_2637);
nor U14965 (N_14965,N_2385,N_4076);
nand U14966 (N_14966,N_8569,N_7180);
and U14967 (N_14967,N_3706,N_982);
nor U14968 (N_14968,N_761,N_1990);
or U14969 (N_14969,N_4171,N_1019);
nor U14970 (N_14970,N_813,N_9480);
nor U14971 (N_14971,N_3605,N_7122);
xor U14972 (N_14972,N_1389,N_9099);
and U14973 (N_14973,N_1174,N_958);
and U14974 (N_14974,N_2398,N_7538);
nor U14975 (N_14975,N_6639,N_5887);
nor U14976 (N_14976,N_1021,N_1321);
xor U14977 (N_14977,N_8123,N_7380);
and U14978 (N_14978,N_1956,N_4482);
or U14979 (N_14979,N_4685,N_4801);
and U14980 (N_14980,N_3981,N_1160);
nor U14981 (N_14981,N_8435,N_9080);
and U14982 (N_14982,N_8372,N_3765);
nand U14983 (N_14983,N_5218,N_9213);
and U14984 (N_14984,N_9513,N_674);
or U14985 (N_14985,N_0,N_9242);
nand U14986 (N_14986,N_9078,N_6125);
nor U14987 (N_14987,N_20,N_844);
nor U14988 (N_14988,N_3383,N_1855);
nand U14989 (N_14989,N_3820,N_5541);
nor U14990 (N_14990,N_4633,N_1779);
or U14991 (N_14991,N_2739,N_3206);
nand U14992 (N_14992,N_3831,N_6803);
and U14993 (N_14993,N_5324,N_5496);
nand U14994 (N_14994,N_1074,N_3494);
nand U14995 (N_14995,N_4844,N_4362);
and U14996 (N_14996,N_5210,N_136);
xor U14997 (N_14997,N_4605,N_9970);
xor U14998 (N_14998,N_3530,N_8594);
or U14999 (N_14999,N_6014,N_6970);
and U15000 (N_15000,N_8093,N_8037);
nor U15001 (N_15001,N_8145,N_4591);
or U15002 (N_15002,N_8520,N_118);
nand U15003 (N_15003,N_8666,N_1934);
and U15004 (N_15004,N_5471,N_6369);
nor U15005 (N_15005,N_7897,N_3061);
or U15006 (N_15006,N_9013,N_124);
or U15007 (N_15007,N_763,N_3785);
nor U15008 (N_15008,N_1010,N_3249);
and U15009 (N_15009,N_1145,N_6333);
or U15010 (N_15010,N_4816,N_8917);
nor U15011 (N_15011,N_9326,N_1226);
or U15012 (N_15012,N_9039,N_3422);
or U15013 (N_15013,N_5658,N_4023);
nand U15014 (N_15014,N_3531,N_7790);
or U15015 (N_15015,N_3503,N_2445);
nor U15016 (N_15016,N_7595,N_4136);
xnor U15017 (N_15017,N_2407,N_556);
nand U15018 (N_15018,N_1528,N_8134);
and U15019 (N_15019,N_4765,N_6315);
and U15020 (N_15020,N_7683,N_9186);
and U15021 (N_15021,N_8499,N_1990);
and U15022 (N_15022,N_6317,N_9834);
nor U15023 (N_15023,N_5752,N_9011);
nor U15024 (N_15024,N_7467,N_1830);
or U15025 (N_15025,N_5328,N_5214);
nor U15026 (N_15026,N_4000,N_6750);
and U15027 (N_15027,N_1499,N_6663);
and U15028 (N_15028,N_4696,N_2846);
and U15029 (N_15029,N_6840,N_4400);
xor U15030 (N_15030,N_7869,N_3199);
or U15031 (N_15031,N_5256,N_5772);
nand U15032 (N_15032,N_5123,N_6340);
and U15033 (N_15033,N_9926,N_5188);
nand U15034 (N_15034,N_7372,N_9344);
nand U15035 (N_15035,N_3980,N_8141);
nand U15036 (N_15036,N_1015,N_317);
nor U15037 (N_15037,N_7516,N_1577);
and U15038 (N_15038,N_3021,N_5181);
or U15039 (N_15039,N_5472,N_54);
nor U15040 (N_15040,N_4564,N_1630);
nand U15041 (N_15041,N_3174,N_9269);
and U15042 (N_15042,N_7327,N_9154);
nor U15043 (N_15043,N_2271,N_1721);
and U15044 (N_15044,N_1570,N_4266);
nand U15045 (N_15045,N_3065,N_2029);
nand U15046 (N_15046,N_6269,N_4933);
or U15047 (N_15047,N_2605,N_4311);
xor U15048 (N_15048,N_3250,N_7643);
or U15049 (N_15049,N_6937,N_5406);
nor U15050 (N_15050,N_3411,N_3708);
or U15051 (N_15051,N_7309,N_2439);
xnor U15052 (N_15052,N_30,N_2439);
or U15053 (N_15053,N_6492,N_3657);
nand U15054 (N_15054,N_1789,N_1167);
xor U15055 (N_15055,N_6117,N_9382);
nand U15056 (N_15056,N_4644,N_3250);
nand U15057 (N_15057,N_684,N_8049);
and U15058 (N_15058,N_7271,N_5741);
or U15059 (N_15059,N_8432,N_7658);
and U15060 (N_15060,N_2049,N_6833);
nor U15061 (N_15061,N_2641,N_2532);
and U15062 (N_15062,N_5597,N_9103);
and U15063 (N_15063,N_2696,N_6513);
xnor U15064 (N_15064,N_6891,N_1292);
or U15065 (N_15065,N_173,N_6371);
nand U15066 (N_15066,N_5019,N_684);
nand U15067 (N_15067,N_3917,N_3367);
and U15068 (N_15068,N_8369,N_1246);
nor U15069 (N_15069,N_911,N_9949);
xnor U15070 (N_15070,N_2290,N_7816);
and U15071 (N_15071,N_4039,N_5421);
and U15072 (N_15072,N_2782,N_1068);
nand U15073 (N_15073,N_7331,N_4351);
or U15074 (N_15074,N_3912,N_5586);
and U15075 (N_15075,N_8125,N_7746);
and U15076 (N_15076,N_6741,N_1456);
and U15077 (N_15077,N_8288,N_5040);
or U15078 (N_15078,N_563,N_2883);
or U15079 (N_15079,N_7891,N_2440);
nor U15080 (N_15080,N_6183,N_1009);
nand U15081 (N_15081,N_1643,N_2462);
nand U15082 (N_15082,N_1915,N_8388);
and U15083 (N_15083,N_8779,N_8011);
nor U15084 (N_15084,N_2693,N_6792);
nand U15085 (N_15085,N_4883,N_7173);
or U15086 (N_15086,N_5790,N_4731);
nand U15087 (N_15087,N_3718,N_5716);
nor U15088 (N_15088,N_7568,N_1789);
xor U15089 (N_15089,N_7912,N_6805);
or U15090 (N_15090,N_8962,N_9426);
nor U15091 (N_15091,N_2712,N_2243);
nand U15092 (N_15092,N_1140,N_7880);
nor U15093 (N_15093,N_4135,N_8880);
nor U15094 (N_15094,N_5704,N_5372);
or U15095 (N_15095,N_4022,N_7872);
xnor U15096 (N_15096,N_5587,N_8551);
and U15097 (N_15097,N_761,N_870);
nand U15098 (N_15098,N_7647,N_356);
nand U15099 (N_15099,N_1360,N_6929);
nor U15100 (N_15100,N_8919,N_7430);
and U15101 (N_15101,N_1203,N_1099);
nand U15102 (N_15102,N_1352,N_3975);
nor U15103 (N_15103,N_8947,N_6933);
and U15104 (N_15104,N_3384,N_6642);
and U15105 (N_15105,N_8469,N_5895);
nand U15106 (N_15106,N_973,N_4164);
or U15107 (N_15107,N_2543,N_3067);
and U15108 (N_15108,N_9425,N_4287);
and U15109 (N_15109,N_2884,N_8620);
and U15110 (N_15110,N_189,N_9299);
and U15111 (N_15111,N_9581,N_5130);
xor U15112 (N_15112,N_5681,N_6659);
nand U15113 (N_15113,N_6370,N_2478);
nor U15114 (N_15114,N_5265,N_8737);
nor U15115 (N_15115,N_2439,N_8235);
nand U15116 (N_15116,N_2880,N_1519);
or U15117 (N_15117,N_9962,N_1566);
and U15118 (N_15118,N_7077,N_2544);
and U15119 (N_15119,N_7425,N_5293);
and U15120 (N_15120,N_9511,N_8782);
or U15121 (N_15121,N_9560,N_5835);
nor U15122 (N_15122,N_5345,N_2922);
nor U15123 (N_15123,N_3150,N_4440);
nor U15124 (N_15124,N_2315,N_8265);
and U15125 (N_15125,N_4382,N_7953);
nor U15126 (N_15126,N_3290,N_6519);
and U15127 (N_15127,N_7965,N_3882);
and U15128 (N_15128,N_5417,N_97);
or U15129 (N_15129,N_1055,N_5741);
or U15130 (N_15130,N_8680,N_9049);
nor U15131 (N_15131,N_4048,N_5906);
and U15132 (N_15132,N_5038,N_5145);
nor U15133 (N_15133,N_6917,N_5749);
xor U15134 (N_15134,N_5982,N_5027);
or U15135 (N_15135,N_1894,N_8733);
and U15136 (N_15136,N_4498,N_337);
or U15137 (N_15137,N_5170,N_3139);
and U15138 (N_15138,N_4141,N_2675);
nor U15139 (N_15139,N_8734,N_9010);
nand U15140 (N_15140,N_4308,N_6822);
nand U15141 (N_15141,N_3039,N_9011);
or U15142 (N_15142,N_162,N_8332);
nand U15143 (N_15143,N_5183,N_5746);
xor U15144 (N_15144,N_828,N_9831);
or U15145 (N_15145,N_6858,N_5428);
nand U15146 (N_15146,N_51,N_6215);
and U15147 (N_15147,N_1840,N_6023);
and U15148 (N_15148,N_4101,N_5161);
nand U15149 (N_15149,N_6858,N_2686);
xnor U15150 (N_15150,N_5772,N_3602);
nor U15151 (N_15151,N_3187,N_562);
nor U15152 (N_15152,N_7818,N_1935);
nor U15153 (N_15153,N_5586,N_553);
nor U15154 (N_15154,N_7401,N_3502);
nand U15155 (N_15155,N_5115,N_5087);
nor U15156 (N_15156,N_1025,N_1003);
and U15157 (N_15157,N_5789,N_3636);
or U15158 (N_15158,N_537,N_7556);
and U15159 (N_15159,N_929,N_4271);
nand U15160 (N_15160,N_6085,N_3792);
or U15161 (N_15161,N_5293,N_6919);
xor U15162 (N_15162,N_2501,N_2237);
and U15163 (N_15163,N_484,N_1756);
nand U15164 (N_15164,N_4063,N_9272);
nor U15165 (N_15165,N_6983,N_4804);
nand U15166 (N_15166,N_8430,N_4089);
or U15167 (N_15167,N_8846,N_4104);
xor U15168 (N_15168,N_4983,N_945);
nand U15169 (N_15169,N_176,N_5257);
or U15170 (N_15170,N_8506,N_7165);
nand U15171 (N_15171,N_4838,N_1127);
nor U15172 (N_15172,N_5467,N_145);
nand U15173 (N_15173,N_1055,N_7537);
nor U15174 (N_15174,N_9112,N_7791);
nor U15175 (N_15175,N_7431,N_1406);
nor U15176 (N_15176,N_2601,N_2972);
or U15177 (N_15177,N_150,N_7636);
xor U15178 (N_15178,N_2869,N_6346);
nand U15179 (N_15179,N_5497,N_9540);
and U15180 (N_15180,N_9516,N_5666);
or U15181 (N_15181,N_5775,N_8614);
nand U15182 (N_15182,N_9886,N_1510);
and U15183 (N_15183,N_9385,N_5787);
nor U15184 (N_15184,N_3235,N_4781);
or U15185 (N_15185,N_2480,N_6690);
nand U15186 (N_15186,N_8939,N_7750);
nand U15187 (N_15187,N_3396,N_5004);
nand U15188 (N_15188,N_1788,N_2276);
nand U15189 (N_15189,N_3967,N_8554);
or U15190 (N_15190,N_3849,N_5707);
xnor U15191 (N_15191,N_6701,N_8364);
xnor U15192 (N_15192,N_3824,N_6140);
nand U15193 (N_15193,N_3264,N_9869);
and U15194 (N_15194,N_1615,N_4819);
nor U15195 (N_15195,N_6561,N_3490);
nand U15196 (N_15196,N_503,N_3255);
nor U15197 (N_15197,N_2235,N_1901);
nor U15198 (N_15198,N_6556,N_4512);
or U15199 (N_15199,N_7045,N_4495);
or U15200 (N_15200,N_6083,N_70);
and U15201 (N_15201,N_4193,N_2952);
nor U15202 (N_15202,N_1315,N_2410);
and U15203 (N_15203,N_5100,N_7707);
nand U15204 (N_15204,N_9941,N_2569);
nor U15205 (N_15205,N_7027,N_5134);
nand U15206 (N_15206,N_2501,N_1491);
and U15207 (N_15207,N_658,N_4640);
or U15208 (N_15208,N_6567,N_2601);
and U15209 (N_15209,N_2468,N_7487);
and U15210 (N_15210,N_7100,N_1582);
and U15211 (N_15211,N_6276,N_3319);
or U15212 (N_15212,N_9513,N_6516);
and U15213 (N_15213,N_9070,N_8065);
nor U15214 (N_15214,N_3727,N_7146);
or U15215 (N_15215,N_7251,N_669);
xor U15216 (N_15216,N_5531,N_1762);
nand U15217 (N_15217,N_7775,N_5566);
and U15218 (N_15218,N_6332,N_9672);
nand U15219 (N_15219,N_7908,N_4604);
nand U15220 (N_15220,N_5565,N_6983);
and U15221 (N_15221,N_6841,N_1696);
nor U15222 (N_15222,N_8666,N_5078);
nor U15223 (N_15223,N_4818,N_1423);
nand U15224 (N_15224,N_7966,N_6204);
nand U15225 (N_15225,N_2888,N_4881);
nand U15226 (N_15226,N_7379,N_7142);
and U15227 (N_15227,N_6985,N_6783);
or U15228 (N_15228,N_9241,N_9228);
or U15229 (N_15229,N_4431,N_3801);
nor U15230 (N_15230,N_9389,N_8053);
nor U15231 (N_15231,N_6931,N_525);
or U15232 (N_15232,N_7282,N_2242);
nor U15233 (N_15233,N_9094,N_2399);
nor U15234 (N_15234,N_7721,N_8654);
and U15235 (N_15235,N_1670,N_5280);
or U15236 (N_15236,N_9705,N_6485);
nand U15237 (N_15237,N_2744,N_5965);
or U15238 (N_15238,N_5418,N_3116);
nand U15239 (N_15239,N_8800,N_6182);
nand U15240 (N_15240,N_2977,N_1920);
or U15241 (N_15241,N_6311,N_8035);
nand U15242 (N_15242,N_4802,N_729);
or U15243 (N_15243,N_3137,N_6674);
or U15244 (N_15244,N_7266,N_1100);
or U15245 (N_15245,N_5360,N_4370);
or U15246 (N_15246,N_8935,N_6640);
or U15247 (N_15247,N_5765,N_1624);
or U15248 (N_15248,N_5689,N_2443);
nor U15249 (N_15249,N_8835,N_8671);
nand U15250 (N_15250,N_1552,N_2354);
and U15251 (N_15251,N_4009,N_1137);
and U15252 (N_15252,N_439,N_9059);
nand U15253 (N_15253,N_8793,N_6184);
nor U15254 (N_15254,N_6480,N_4143);
and U15255 (N_15255,N_2058,N_1149);
and U15256 (N_15256,N_1802,N_6864);
and U15257 (N_15257,N_9478,N_6238);
nand U15258 (N_15258,N_1549,N_6852);
nor U15259 (N_15259,N_7550,N_1282);
nor U15260 (N_15260,N_6293,N_1272);
nor U15261 (N_15261,N_1237,N_5061);
nand U15262 (N_15262,N_9781,N_2893);
nand U15263 (N_15263,N_5379,N_8839);
nand U15264 (N_15264,N_751,N_5171);
nand U15265 (N_15265,N_5499,N_454);
or U15266 (N_15266,N_2527,N_5402);
nand U15267 (N_15267,N_7405,N_8235);
and U15268 (N_15268,N_9687,N_4937);
or U15269 (N_15269,N_1201,N_5927);
and U15270 (N_15270,N_1371,N_5443);
nand U15271 (N_15271,N_8628,N_4058);
and U15272 (N_15272,N_9996,N_4297);
nand U15273 (N_15273,N_7057,N_7521);
nand U15274 (N_15274,N_9873,N_7803);
and U15275 (N_15275,N_85,N_3542);
nand U15276 (N_15276,N_9306,N_1195);
nand U15277 (N_15277,N_2730,N_4636);
or U15278 (N_15278,N_5850,N_8790);
xnor U15279 (N_15279,N_8721,N_4164);
nand U15280 (N_15280,N_5894,N_2918);
nand U15281 (N_15281,N_2887,N_1289);
or U15282 (N_15282,N_4585,N_3380);
or U15283 (N_15283,N_9282,N_663);
xnor U15284 (N_15284,N_9330,N_4815);
nand U15285 (N_15285,N_6306,N_8729);
or U15286 (N_15286,N_8940,N_6932);
or U15287 (N_15287,N_1703,N_5917);
and U15288 (N_15288,N_5389,N_2481);
nand U15289 (N_15289,N_5774,N_9335);
nand U15290 (N_15290,N_6903,N_5329);
and U15291 (N_15291,N_1253,N_5529);
and U15292 (N_15292,N_6033,N_9234);
and U15293 (N_15293,N_1334,N_8133);
nor U15294 (N_15294,N_5222,N_1132);
and U15295 (N_15295,N_6852,N_6860);
nand U15296 (N_15296,N_8028,N_3433);
or U15297 (N_15297,N_8471,N_9773);
or U15298 (N_15298,N_5640,N_8587);
or U15299 (N_15299,N_3201,N_4504);
xor U15300 (N_15300,N_3262,N_2534);
nand U15301 (N_15301,N_4746,N_3900);
xnor U15302 (N_15302,N_8205,N_6917);
nand U15303 (N_15303,N_973,N_1176);
or U15304 (N_15304,N_1,N_5755);
nand U15305 (N_15305,N_2580,N_4284);
or U15306 (N_15306,N_8794,N_5874);
and U15307 (N_15307,N_9157,N_9403);
nor U15308 (N_15308,N_3864,N_3258);
nor U15309 (N_15309,N_9176,N_8026);
or U15310 (N_15310,N_6886,N_8416);
nor U15311 (N_15311,N_6465,N_6401);
and U15312 (N_15312,N_4119,N_1996);
or U15313 (N_15313,N_9954,N_3461);
or U15314 (N_15314,N_2559,N_4164);
nor U15315 (N_15315,N_7557,N_2500);
and U15316 (N_15316,N_8964,N_2895);
xnor U15317 (N_15317,N_5887,N_928);
xor U15318 (N_15318,N_6727,N_8527);
and U15319 (N_15319,N_2268,N_3479);
nand U15320 (N_15320,N_1775,N_5906);
or U15321 (N_15321,N_6104,N_590);
nand U15322 (N_15322,N_2420,N_8467);
or U15323 (N_15323,N_9490,N_1733);
nand U15324 (N_15324,N_4283,N_9719);
nand U15325 (N_15325,N_8620,N_4449);
or U15326 (N_15326,N_7737,N_8931);
or U15327 (N_15327,N_2857,N_9722);
nor U15328 (N_15328,N_6117,N_8267);
or U15329 (N_15329,N_7800,N_4987);
xor U15330 (N_15330,N_265,N_2601);
nand U15331 (N_15331,N_5903,N_7685);
nand U15332 (N_15332,N_4757,N_3410);
nor U15333 (N_15333,N_2284,N_1017);
nor U15334 (N_15334,N_4248,N_9922);
xnor U15335 (N_15335,N_2634,N_5078);
nor U15336 (N_15336,N_3358,N_1392);
or U15337 (N_15337,N_221,N_8762);
and U15338 (N_15338,N_6497,N_1725);
or U15339 (N_15339,N_6777,N_6093);
and U15340 (N_15340,N_9089,N_3352);
or U15341 (N_15341,N_2129,N_1594);
nand U15342 (N_15342,N_1707,N_1015);
and U15343 (N_15343,N_4417,N_295);
or U15344 (N_15344,N_3864,N_1490);
and U15345 (N_15345,N_5598,N_7535);
nor U15346 (N_15346,N_8074,N_2906);
and U15347 (N_15347,N_1026,N_1973);
nand U15348 (N_15348,N_966,N_5111);
nand U15349 (N_15349,N_2827,N_8761);
and U15350 (N_15350,N_7,N_5029);
or U15351 (N_15351,N_8675,N_9131);
nor U15352 (N_15352,N_2469,N_7754);
and U15353 (N_15353,N_4208,N_2999);
nor U15354 (N_15354,N_7707,N_1184);
nand U15355 (N_15355,N_2276,N_3067);
nand U15356 (N_15356,N_3101,N_8321);
and U15357 (N_15357,N_7916,N_7511);
or U15358 (N_15358,N_3193,N_3244);
nand U15359 (N_15359,N_9548,N_3673);
nor U15360 (N_15360,N_5785,N_5933);
or U15361 (N_15361,N_3425,N_195);
nor U15362 (N_15362,N_6281,N_5525);
nor U15363 (N_15363,N_4649,N_1711);
nor U15364 (N_15364,N_5550,N_9494);
xor U15365 (N_15365,N_5127,N_3261);
and U15366 (N_15366,N_9280,N_7773);
nand U15367 (N_15367,N_9264,N_3527);
nor U15368 (N_15368,N_4582,N_591);
nor U15369 (N_15369,N_5583,N_6850);
or U15370 (N_15370,N_5625,N_147);
or U15371 (N_15371,N_6728,N_4211);
nand U15372 (N_15372,N_7667,N_718);
nand U15373 (N_15373,N_1578,N_3182);
nand U15374 (N_15374,N_7297,N_402);
and U15375 (N_15375,N_1019,N_6580);
or U15376 (N_15376,N_6675,N_8374);
xor U15377 (N_15377,N_4253,N_2198);
nand U15378 (N_15378,N_2158,N_5945);
nor U15379 (N_15379,N_1912,N_657);
nor U15380 (N_15380,N_7212,N_2289);
nand U15381 (N_15381,N_3441,N_2263);
and U15382 (N_15382,N_3227,N_4319);
nand U15383 (N_15383,N_1608,N_5873);
xnor U15384 (N_15384,N_7963,N_6830);
or U15385 (N_15385,N_6212,N_6567);
and U15386 (N_15386,N_8648,N_4425);
nand U15387 (N_15387,N_1775,N_9614);
xnor U15388 (N_15388,N_2355,N_5318);
and U15389 (N_15389,N_5153,N_6775);
or U15390 (N_15390,N_3739,N_4631);
or U15391 (N_15391,N_7639,N_1886);
and U15392 (N_15392,N_7405,N_923);
and U15393 (N_15393,N_1725,N_2636);
and U15394 (N_15394,N_3074,N_6895);
and U15395 (N_15395,N_7105,N_320);
nand U15396 (N_15396,N_4885,N_4309);
nand U15397 (N_15397,N_1945,N_5757);
nor U15398 (N_15398,N_1067,N_6738);
or U15399 (N_15399,N_1368,N_723);
nor U15400 (N_15400,N_5156,N_9054);
nor U15401 (N_15401,N_2363,N_1493);
xnor U15402 (N_15402,N_914,N_7256);
or U15403 (N_15403,N_4574,N_3624);
or U15404 (N_15404,N_3596,N_8510);
nand U15405 (N_15405,N_2795,N_6697);
nor U15406 (N_15406,N_9343,N_5568);
or U15407 (N_15407,N_151,N_4651);
nor U15408 (N_15408,N_2589,N_6440);
xor U15409 (N_15409,N_5937,N_4579);
nand U15410 (N_15410,N_9358,N_5601);
or U15411 (N_15411,N_3071,N_4423);
xor U15412 (N_15412,N_5268,N_9475);
and U15413 (N_15413,N_6358,N_6027);
xor U15414 (N_15414,N_1031,N_7849);
or U15415 (N_15415,N_2711,N_9113);
nor U15416 (N_15416,N_966,N_8943);
nor U15417 (N_15417,N_9252,N_7449);
nand U15418 (N_15418,N_5303,N_8930);
and U15419 (N_15419,N_8629,N_3662);
or U15420 (N_15420,N_1467,N_2441);
nor U15421 (N_15421,N_3304,N_1356);
and U15422 (N_15422,N_1541,N_224);
xnor U15423 (N_15423,N_9348,N_2110);
nor U15424 (N_15424,N_8945,N_902);
nand U15425 (N_15425,N_4463,N_3088);
nor U15426 (N_15426,N_7383,N_3102);
xor U15427 (N_15427,N_7468,N_4050);
xnor U15428 (N_15428,N_5977,N_7914);
nor U15429 (N_15429,N_3227,N_8863);
nor U15430 (N_15430,N_222,N_9232);
nand U15431 (N_15431,N_8907,N_7572);
xnor U15432 (N_15432,N_1104,N_5567);
or U15433 (N_15433,N_714,N_8204);
or U15434 (N_15434,N_8565,N_4667);
nor U15435 (N_15435,N_7970,N_2960);
nor U15436 (N_15436,N_4301,N_1900);
nand U15437 (N_15437,N_6395,N_7703);
xnor U15438 (N_15438,N_3939,N_1500);
nand U15439 (N_15439,N_9138,N_2466);
and U15440 (N_15440,N_8981,N_1115);
or U15441 (N_15441,N_2300,N_9743);
nor U15442 (N_15442,N_5964,N_2867);
nand U15443 (N_15443,N_1104,N_1063);
xnor U15444 (N_15444,N_9544,N_967);
or U15445 (N_15445,N_3255,N_1099);
nand U15446 (N_15446,N_1426,N_7887);
nor U15447 (N_15447,N_8989,N_7666);
nor U15448 (N_15448,N_8487,N_8386);
nor U15449 (N_15449,N_6366,N_4385);
and U15450 (N_15450,N_2489,N_6595);
and U15451 (N_15451,N_7775,N_25);
or U15452 (N_15452,N_4901,N_4346);
or U15453 (N_15453,N_1137,N_7771);
nor U15454 (N_15454,N_8039,N_8990);
and U15455 (N_15455,N_694,N_9164);
nor U15456 (N_15456,N_7396,N_1703);
xor U15457 (N_15457,N_9972,N_260);
nand U15458 (N_15458,N_6219,N_687);
nand U15459 (N_15459,N_177,N_116);
and U15460 (N_15460,N_931,N_925);
nor U15461 (N_15461,N_9516,N_3418);
nor U15462 (N_15462,N_7625,N_6778);
nor U15463 (N_15463,N_4984,N_2706);
or U15464 (N_15464,N_7655,N_1112);
and U15465 (N_15465,N_5891,N_1477);
nor U15466 (N_15466,N_3205,N_2619);
and U15467 (N_15467,N_8362,N_7805);
xor U15468 (N_15468,N_239,N_445);
nor U15469 (N_15469,N_8309,N_6240);
or U15470 (N_15470,N_8483,N_2087);
nor U15471 (N_15471,N_417,N_1963);
xnor U15472 (N_15472,N_4398,N_7647);
nor U15473 (N_15473,N_5094,N_8202);
or U15474 (N_15474,N_3245,N_4391);
and U15475 (N_15475,N_9337,N_1685);
and U15476 (N_15476,N_707,N_6631);
nand U15477 (N_15477,N_3629,N_520);
nand U15478 (N_15478,N_3833,N_4713);
and U15479 (N_15479,N_1543,N_7916);
and U15480 (N_15480,N_7136,N_4302);
or U15481 (N_15481,N_1564,N_3045);
and U15482 (N_15482,N_210,N_6568);
nor U15483 (N_15483,N_424,N_1189);
nand U15484 (N_15484,N_5246,N_4494);
nor U15485 (N_15485,N_5488,N_6134);
and U15486 (N_15486,N_1345,N_3200);
or U15487 (N_15487,N_3144,N_8445);
xnor U15488 (N_15488,N_7817,N_2554);
and U15489 (N_15489,N_107,N_9865);
or U15490 (N_15490,N_8157,N_6183);
or U15491 (N_15491,N_8738,N_5277);
nor U15492 (N_15492,N_2658,N_9908);
or U15493 (N_15493,N_1240,N_2761);
nor U15494 (N_15494,N_5572,N_6706);
xnor U15495 (N_15495,N_6495,N_1650);
and U15496 (N_15496,N_5916,N_5452);
nor U15497 (N_15497,N_8075,N_1671);
or U15498 (N_15498,N_4572,N_8187);
and U15499 (N_15499,N_8932,N_9696);
or U15500 (N_15500,N_3590,N_37);
or U15501 (N_15501,N_9541,N_9832);
or U15502 (N_15502,N_5465,N_2600);
nor U15503 (N_15503,N_2850,N_6134);
nor U15504 (N_15504,N_4325,N_5950);
nor U15505 (N_15505,N_3642,N_6918);
nand U15506 (N_15506,N_5843,N_5800);
nand U15507 (N_15507,N_3182,N_1814);
or U15508 (N_15508,N_6901,N_2370);
nand U15509 (N_15509,N_3053,N_8863);
or U15510 (N_15510,N_3566,N_6389);
nor U15511 (N_15511,N_209,N_207);
nor U15512 (N_15512,N_3456,N_328);
or U15513 (N_15513,N_378,N_1655);
or U15514 (N_15514,N_2636,N_693);
xnor U15515 (N_15515,N_4693,N_4073);
nand U15516 (N_15516,N_7098,N_8803);
nor U15517 (N_15517,N_6020,N_7987);
and U15518 (N_15518,N_3066,N_9679);
and U15519 (N_15519,N_8225,N_6747);
nand U15520 (N_15520,N_3993,N_6794);
nor U15521 (N_15521,N_9013,N_2019);
nand U15522 (N_15522,N_3248,N_3375);
nor U15523 (N_15523,N_7990,N_6386);
and U15524 (N_15524,N_2731,N_2435);
nand U15525 (N_15525,N_7217,N_1297);
xor U15526 (N_15526,N_3602,N_881);
or U15527 (N_15527,N_849,N_14);
or U15528 (N_15528,N_212,N_3390);
nand U15529 (N_15529,N_4412,N_6118);
nor U15530 (N_15530,N_3170,N_3480);
nor U15531 (N_15531,N_8076,N_5783);
or U15532 (N_15532,N_9369,N_5162);
or U15533 (N_15533,N_9316,N_3226);
nor U15534 (N_15534,N_917,N_8075);
and U15535 (N_15535,N_6398,N_164);
and U15536 (N_15536,N_5855,N_5777);
nor U15537 (N_15537,N_1513,N_8422);
nor U15538 (N_15538,N_9590,N_2684);
nor U15539 (N_15539,N_9951,N_6600);
nand U15540 (N_15540,N_6295,N_2344);
nand U15541 (N_15541,N_1666,N_574);
and U15542 (N_15542,N_7942,N_6712);
or U15543 (N_15543,N_8553,N_8025);
or U15544 (N_15544,N_4147,N_1355);
or U15545 (N_15545,N_2489,N_6488);
nor U15546 (N_15546,N_702,N_4347);
or U15547 (N_15547,N_3433,N_1939);
or U15548 (N_15548,N_112,N_9423);
nor U15549 (N_15549,N_480,N_8983);
or U15550 (N_15550,N_4005,N_4822);
and U15551 (N_15551,N_5495,N_7665);
or U15552 (N_15552,N_9697,N_5974);
nor U15553 (N_15553,N_8251,N_8594);
nor U15554 (N_15554,N_4141,N_3477);
xor U15555 (N_15555,N_7058,N_1349);
and U15556 (N_15556,N_3826,N_6827);
and U15557 (N_15557,N_1856,N_7201);
or U15558 (N_15558,N_6595,N_638);
or U15559 (N_15559,N_5472,N_5020);
xor U15560 (N_15560,N_6585,N_5186);
or U15561 (N_15561,N_8229,N_6284);
nand U15562 (N_15562,N_5492,N_1132);
or U15563 (N_15563,N_9797,N_4091);
or U15564 (N_15564,N_3344,N_8561);
xnor U15565 (N_15565,N_7947,N_5048);
or U15566 (N_15566,N_5163,N_7426);
and U15567 (N_15567,N_9307,N_6583);
or U15568 (N_15568,N_4121,N_8817);
and U15569 (N_15569,N_2675,N_6297);
and U15570 (N_15570,N_7857,N_1569);
and U15571 (N_15571,N_3111,N_9064);
or U15572 (N_15572,N_280,N_4983);
or U15573 (N_15573,N_7082,N_7468);
nand U15574 (N_15574,N_3021,N_5994);
nor U15575 (N_15575,N_3866,N_7734);
nor U15576 (N_15576,N_4214,N_7501);
nor U15577 (N_15577,N_283,N_8353);
and U15578 (N_15578,N_9271,N_8340);
and U15579 (N_15579,N_1007,N_5581);
and U15580 (N_15580,N_1047,N_6991);
nand U15581 (N_15581,N_1395,N_1253);
or U15582 (N_15582,N_6550,N_917);
or U15583 (N_15583,N_8119,N_907);
nor U15584 (N_15584,N_7691,N_7593);
nor U15585 (N_15585,N_3011,N_1499);
or U15586 (N_15586,N_5550,N_6257);
nor U15587 (N_15587,N_5175,N_8766);
or U15588 (N_15588,N_5468,N_7202);
or U15589 (N_15589,N_8374,N_1602);
nor U15590 (N_15590,N_7579,N_4341);
nor U15591 (N_15591,N_475,N_4049);
or U15592 (N_15592,N_6759,N_1289);
or U15593 (N_15593,N_4320,N_3571);
nor U15594 (N_15594,N_6612,N_2810);
nand U15595 (N_15595,N_2343,N_8);
and U15596 (N_15596,N_7037,N_7606);
nor U15597 (N_15597,N_4114,N_5263);
or U15598 (N_15598,N_3797,N_7788);
xnor U15599 (N_15599,N_7895,N_4172);
nand U15600 (N_15600,N_8133,N_6471);
nor U15601 (N_15601,N_8662,N_5941);
nor U15602 (N_15602,N_4430,N_4762);
or U15603 (N_15603,N_6007,N_7266);
nor U15604 (N_15604,N_2250,N_1577);
nand U15605 (N_15605,N_3846,N_3149);
xnor U15606 (N_15606,N_4781,N_8441);
nand U15607 (N_15607,N_8821,N_8167);
or U15608 (N_15608,N_4676,N_315);
nand U15609 (N_15609,N_191,N_6704);
or U15610 (N_15610,N_4793,N_1010);
nand U15611 (N_15611,N_4377,N_5631);
xor U15612 (N_15612,N_9731,N_1686);
or U15613 (N_15613,N_633,N_2527);
nand U15614 (N_15614,N_9659,N_5269);
or U15615 (N_15615,N_6860,N_867);
and U15616 (N_15616,N_6755,N_5030);
nor U15617 (N_15617,N_1247,N_6764);
and U15618 (N_15618,N_1314,N_7206);
nor U15619 (N_15619,N_8515,N_9099);
xnor U15620 (N_15620,N_6820,N_423);
or U15621 (N_15621,N_2081,N_5415);
nand U15622 (N_15622,N_7792,N_2489);
nand U15623 (N_15623,N_1532,N_1945);
and U15624 (N_15624,N_2588,N_590);
nand U15625 (N_15625,N_603,N_8326);
and U15626 (N_15626,N_4700,N_5655);
nor U15627 (N_15627,N_9225,N_4502);
xnor U15628 (N_15628,N_4531,N_7311);
and U15629 (N_15629,N_8076,N_1275);
nand U15630 (N_15630,N_6437,N_7740);
or U15631 (N_15631,N_9799,N_6086);
nand U15632 (N_15632,N_8999,N_6129);
nor U15633 (N_15633,N_4743,N_6630);
nor U15634 (N_15634,N_4159,N_2645);
or U15635 (N_15635,N_3243,N_8684);
xnor U15636 (N_15636,N_6345,N_6434);
nor U15637 (N_15637,N_7511,N_924);
or U15638 (N_15638,N_2192,N_6690);
and U15639 (N_15639,N_5423,N_7110);
and U15640 (N_15640,N_2533,N_9584);
and U15641 (N_15641,N_1271,N_2758);
and U15642 (N_15642,N_1304,N_2504);
and U15643 (N_15643,N_3086,N_6307);
xor U15644 (N_15644,N_8647,N_6354);
nand U15645 (N_15645,N_3173,N_1307);
or U15646 (N_15646,N_537,N_1034);
or U15647 (N_15647,N_2833,N_2388);
nand U15648 (N_15648,N_1207,N_876);
or U15649 (N_15649,N_7023,N_1894);
nand U15650 (N_15650,N_5606,N_390);
nor U15651 (N_15651,N_9337,N_2438);
and U15652 (N_15652,N_6086,N_7716);
or U15653 (N_15653,N_5175,N_7181);
and U15654 (N_15654,N_9529,N_2539);
nand U15655 (N_15655,N_738,N_8894);
xor U15656 (N_15656,N_756,N_7454);
or U15657 (N_15657,N_4814,N_7966);
nor U15658 (N_15658,N_6943,N_5197);
nor U15659 (N_15659,N_2371,N_1784);
nor U15660 (N_15660,N_4408,N_8385);
nor U15661 (N_15661,N_3691,N_1023);
and U15662 (N_15662,N_9766,N_3935);
nor U15663 (N_15663,N_9360,N_6139);
and U15664 (N_15664,N_6876,N_1727);
or U15665 (N_15665,N_5004,N_3551);
and U15666 (N_15666,N_1559,N_7888);
nand U15667 (N_15667,N_5705,N_9448);
and U15668 (N_15668,N_1147,N_1428);
nand U15669 (N_15669,N_9654,N_4903);
and U15670 (N_15670,N_8945,N_7764);
and U15671 (N_15671,N_5686,N_68);
nor U15672 (N_15672,N_1833,N_9797);
xnor U15673 (N_15673,N_739,N_8457);
and U15674 (N_15674,N_9232,N_8443);
nand U15675 (N_15675,N_7814,N_9306);
nor U15676 (N_15676,N_4549,N_9230);
and U15677 (N_15677,N_7200,N_3460);
nor U15678 (N_15678,N_3928,N_5842);
nand U15679 (N_15679,N_5544,N_9617);
xnor U15680 (N_15680,N_3621,N_4602);
nand U15681 (N_15681,N_5239,N_2867);
nand U15682 (N_15682,N_6691,N_5392);
nor U15683 (N_15683,N_6840,N_9762);
and U15684 (N_15684,N_5391,N_3115);
and U15685 (N_15685,N_2751,N_7592);
and U15686 (N_15686,N_6599,N_8501);
nand U15687 (N_15687,N_3004,N_4069);
or U15688 (N_15688,N_3858,N_3751);
nor U15689 (N_15689,N_1678,N_1219);
xnor U15690 (N_15690,N_3907,N_2383);
and U15691 (N_15691,N_262,N_3939);
or U15692 (N_15692,N_6652,N_3867);
and U15693 (N_15693,N_4640,N_8269);
nor U15694 (N_15694,N_5525,N_8312);
and U15695 (N_15695,N_9403,N_4892);
and U15696 (N_15696,N_424,N_786);
or U15697 (N_15697,N_8398,N_6687);
xor U15698 (N_15698,N_7757,N_6633);
nor U15699 (N_15699,N_7567,N_4671);
or U15700 (N_15700,N_3065,N_2432);
or U15701 (N_15701,N_7472,N_7551);
xnor U15702 (N_15702,N_8843,N_3819);
nand U15703 (N_15703,N_6648,N_1196);
or U15704 (N_15704,N_6076,N_9233);
nor U15705 (N_15705,N_3518,N_5883);
and U15706 (N_15706,N_3129,N_8221);
nor U15707 (N_15707,N_1604,N_9275);
nand U15708 (N_15708,N_1862,N_7165);
xor U15709 (N_15709,N_5081,N_3744);
nor U15710 (N_15710,N_6059,N_8682);
nand U15711 (N_15711,N_6385,N_7310);
and U15712 (N_15712,N_3727,N_1249);
nor U15713 (N_15713,N_676,N_5366);
nor U15714 (N_15714,N_2527,N_1538);
and U15715 (N_15715,N_9560,N_4434);
nor U15716 (N_15716,N_2045,N_2020);
and U15717 (N_15717,N_5319,N_7807);
or U15718 (N_15718,N_7016,N_3161);
or U15719 (N_15719,N_4366,N_4088);
nor U15720 (N_15720,N_9240,N_1401);
and U15721 (N_15721,N_385,N_6271);
nor U15722 (N_15722,N_904,N_5613);
xnor U15723 (N_15723,N_7090,N_3715);
and U15724 (N_15724,N_3638,N_8137);
and U15725 (N_15725,N_8469,N_1208);
or U15726 (N_15726,N_1995,N_416);
nand U15727 (N_15727,N_8893,N_8179);
nand U15728 (N_15728,N_9356,N_5926);
xor U15729 (N_15729,N_8656,N_8692);
or U15730 (N_15730,N_65,N_365);
or U15731 (N_15731,N_4239,N_1675);
or U15732 (N_15732,N_6672,N_3193);
xnor U15733 (N_15733,N_9264,N_3692);
or U15734 (N_15734,N_4998,N_5043);
nor U15735 (N_15735,N_9414,N_3671);
nor U15736 (N_15736,N_9610,N_3581);
and U15737 (N_15737,N_4188,N_5116);
and U15738 (N_15738,N_8075,N_9366);
or U15739 (N_15739,N_3672,N_4106);
nand U15740 (N_15740,N_6540,N_2872);
or U15741 (N_15741,N_5519,N_2880);
or U15742 (N_15742,N_704,N_8337);
and U15743 (N_15743,N_2337,N_1068);
and U15744 (N_15744,N_9503,N_3592);
nor U15745 (N_15745,N_6309,N_4730);
or U15746 (N_15746,N_284,N_8824);
nor U15747 (N_15747,N_1185,N_1646);
or U15748 (N_15748,N_4848,N_8200);
or U15749 (N_15749,N_100,N_6929);
nor U15750 (N_15750,N_4213,N_1650);
nor U15751 (N_15751,N_3096,N_5753);
nand U15752 (N_15752,N_6872,N_2231);
nor U15753 (N_15753,N_5106,N_169);
nand U15754 (N_15754,N_2712,N_1392);
and U15755 (N_15755,N_1123,N_2581);
nand U15756 (N_15756,N_2378,N_4367);
and U15757 (N_15757,N_8338,N_7980);
and U15758 (N_15758,N_2179,N_4142);
xor U15759 (N_15759,N_8144,N_3391);
nand U15760 (N_15760,N_8125,N_1505);
nor U15761 (N_15761,N_9207,N_2041);
and U15762 (N_15762,N_3315,N_3135);
nor U15763 (N_15763,N_920,N_7657);
nand U15764 (N_15764,N_2941,N_4412);
nand U15765 (N_15765,N_6592,N_5022);
and U15766 (N_15766,N_2325,N_3121);
or U15767 (N_15767,N_8413,N_6864);
or U15768 (N_15768,N_6536,N_8788);
nand U15769 (N_15769,N_2553,N_7335);
nor U15770 (N_15770,N_4553,N_8316);
and U15771 (N_15771,N_4511,N_1526);
and U15772 (N_15772,N_4430,N_7402);
xor U15773 (N_15773,N_3900,N_9689);
or U15774 (N_15774,N_6589,N_1528);
or U15775 (N_15775,N_4960,N_5833);
nand U15776 (N_15776,N_9258,N_1477);
or U15777 (N_15777,N_4650,N_3180);
nor U15778 (N_15778,N_8466,N_8230);
and U15779 (N_15779,N_9849,N_1779);
nor U15780 (N_15780,N_5429,N_1836);
and U15781 (N_15781,N_9001,N_7236);
nor U15782 (N_15782,N_4871,N_8165);
and U15783 (N_15783,N_2716,N_8588);
or U15784 (N_15784,N_1506,N_4009);
and U15785 (N_15785,N_2997,N_199);
or U15786 (N_15786,N_4336,N_2577);
nand U15787 (N_15787,N_2880,N_7932);
or U15788 (N_15788,N_2245,N_6399);
or U15789 (N_15789,N_8645,N_4010);
nand U15790 (N_15790,N_3586,N_6675);
or U15791 (N_15791,N_9305,N_8336);
nor U15792 (N_15792,N_2086,N_4674);
and U15793 (N_15793,N_8731,N_802);
nand U15794 (N_15794,N_9719,N_128);
nand U15795 (N_15795,N_3466,N_1851);
and U15796 (N_15796,N_1858,N_8394);
or U15797 (N_15797,N_2641,N_7372);
and U15798 (N_15798,N_8070,N_7752);
and U15799 (N_15799,N_7658,N_6156);
xor U15800 (N_15800,N_410,N_47);
nand U15801 (N_15801,N_1535,N_3390);
and U15802 (N_15802,N_3766,N_5801);
and U15803 (N_15803,N_5260,N_2299);
nor U15804 (N_15804,N_7927,N_6143);
nand U15805 (N_15805,N_1119,N_4932);
or U15806 (N_15806,N_7488,N_2306);
and U15807 (N_15807,N_477,N_535);
or U15808 (N_15808,N_7337,N_4573);
nor U15809 (N_15809,N_2511,N_6217);
xor U15810 (N_15810,N_5006,N_9849);
nand U15811 (N_15811,N_6966,N_7586);
or U15812 (N_15812,N_6345,N_7179);
nor U15813 (N_15813,N_295,N_3518);
and U15814 (N_15814,N_6767,N_4199);
nor U15815 (N_15815,N_278,N_3886);
or U15816 (N_15816,N_9015,N_2536);
and U15817 (N_15817,N_2023,N_4403);
nand U15818 (N_15818,N_8331,N_1082);
nand U15819 (N_15819,N_229,N_5285);
nand U15820 (N_15820,N_3084,N_5757);
nand U15821 (N_15821,N_9995,N_4728);
nor U15822 (N_15822,N_3719,N_5155);
nand U15823 (N_15823,N_8563,N_108);
or U15824 (N_15824,N_9738,N_2487);
or U15825 (N_15825,N_3403,N_8013);
nand U15826 (N_15826,N_1431,N_2632);
or U15827 (N_15827,N_4769,N_8447);
and U15828 (N_15828,N_4352,N_3804);
nand U15829 (N_15829,N_1228,N_6527);
and U15830 (N_15830,N_889,N_6161);
nand U15831 (N_15831,N_7500,N_6215);
and U15832 (N_15832,N_4900,N_3433);
or U15833 (N_15833,N_569,N_7218);
xnor U15834 (N_15834,N_8663,N_7153);
nor U15835 (N_15835,N_4123,N_2313);
nand U15836 (N_15836,N_2832,N_8039);
nand U15837 (N_15837,N_5164,N_9210);
nand U15838 (N_15838,N_509,N_2065);
xor U15839 (N_15839,N_363,N_6193);
and U15840 (N_15840,N_7132,N_7413);
nand U15841 (N_15841,N_1101,N_1483);
nor U15842 (N_15842,N_3657,N_860);
nand U15843 (N_15843,N_4433,N_1810);
nand U15844 (N_15844,N_6276,N_461);
nand U15845 (N_15845,N_3323,N_4422);
or U15846 (N_15846,N_6142,N_7613);
xor U15847 (N_15847,N_23,N_590);
nor U15848 (N_15848,N_1991,N_2398);
nor U15849 (N_15849,N_2125,N_7256);
nor U15850 (N_15850,N_6465,N_4253);
and U15851 (N_15851,N_6461,N_9063);
or U15852 (N_15852,N_6548,N_8239);
nand U15853 (N_15853,N_6629,N_1349);
or U15854 (N_15854,N_7584,N_3096);
or U15855 (N_15855,N_5530,N_4152);
xnor U15856 (N_15856,N_4569,N_6841);
nor U15857 (N_15857,N_5576,N_5412);
or U15858 (N_15858,N_707,N_4242);
and U15859 (N_15859,N_9839,N_7826);
nand U15860 (N_15860,N_2185,N_8119);
or U15861 (N_15861,N_6461,N_6602);
nand U15862 (N_15862,N_6640,N_3598);
nor U15863 (N_15863,N_5501,N_4282);
and U15864 (N_15864,N_3190,N_3014);
or U15865 (N_15865,N_1969,N_825);
xor U15866 (N_15866,N_4180,N_3694);
xor U15867 (N_15867,N_9121,N_5568);
and U15868 (N_15868,N_2771,N_3583);
nand U15869 (N_15869,N_3884,N_9950);
xor U15870 (N_15870,N_9787,N_1607);
nand U15871 (N_15871,N_7290,N_8914);
nor U15872 (N_15872,N_1832,N_896);
nand U15873 (N_15873,N_9443,N_4639);
xnor U15874 (N_15874,N_3888,N_3237);
xor U15875 (N_15875,N_4361,N_1390);
nand U15876 (N_15876,N_7095,N_2872);
xnor U15877 (N_15877,N_9015,N_9156);
or U15878 (N_15878,N_4385,N_1604);
and U15879 (N_15879,N_5679,N_1964);
nand U15880 (N_15880,N_8810,N_3419);
or U15881 (N_15881,N_6563,N_5858);
and U15882 (N_15882,N_4116,N_6327);
xor U15883 (N_15883,N_6024,N_4350);
nor U15884 (N_15884,N_9801,N_176);
or U15885 (N_15885,N_4414,N_7022);
nand U15886 (N_15886,N_4360,N_9358);
or U15887 (N_15887,N_7615,N_3455);
nor U15888 (N_15888,N_2057,N_3515);
or U15889 (N_15889,N_7350,N_5826);
and U15890 (N_15890,N_9934,N_3238);
or U15891 (N_15891,N_6838,N_8911);
xor U15892 (N_15892,N_2701,N_7749);
xor U15893 (N_15893,N_5139,N_1264);
or U15894 (N_15894,N_198,N_3938);
or U15895 (N_15895,N_3900,N_3984);
nand U15896 (N_15896,N_6102,N_6146);
xnor U15897 (N_15897,N_8376,N_2086);
and U15898 (N_15898,N_7945,N_1064);
nand U15899 (N_15899,N_5688,N_244);
and U15900 (N_15900,N_6441,N_4296);
or U15901 (N_15901,N_3491,N_8630);
nor U15902 (N_15902,N_5876,N_763);
or U15903 (N_15903,N_3550,N_9304);
xnor U15904 (N_15904,N_934,N_6608);
or U15905 (N_15905,N_3118,N_2660);
or U15906 (N_15906,N_2884,N_8234);
nor U15907 (N_15907,N_758,N_7905);
or U15908 (N_15908,N_6013,N_3281);
nand U15909 (N_15909,N_5140,N_3242);
or U15910 (N_15910,N_2941,N_3407);
or U15911 (N_15911,N_6207,N_8572);
and U15912 (N_15912,N_5432,N_6497);
or U15913 (N_15913,N_4178,N_6432);
nor U15914 (N_15914,N_8217,N_9502);
or U15915 (N_15915,N_4642,N_8285);
and U15916 (N_15916,N_5504,N_9785);
and U15917 (N_15917,N_7317,N_8442);
or U15918 (N_15918,N_4027,N_1096);
and U15919 (N_15919,N_7522,N_5927);
nand U15920 (N_15920,N_8600,N_2439);
or U15921 (N_15921,N_6656,N_3594);
nor U15922 (N_15922,N_2,N_276);
nand U15923 (N_15923,N_12,N_6778);
or U15924 (N_15924,N_2685,N_2237);
and U15925 (N_15925,N_9990,N_2815);
xor U15926 (N_15926,N_9604,N_9660);
or U15927 (N_15927,N_4906,N_8210);
xor U15928 (N_15928,N_7548,N_9797);
and U15929 (N_15929,N_9405,N_2975);
nor U15930 (N_15930,N_7571,N_3620);
nor U15931 (N_15931,N_1403,N_135);
nand U15932 (N_15932,N_3427,N_1626);
nand U15933 (N_15933,N_393,N_7294);
and U15934 (N_15934,N_4146,N_1712);
nand U15935 (N_15935,N_6659,N_9316);
nor U15936 (N_15936,N_2990,N_4129);
and U15937 (N_15937,N_3419,N_9624);
and U15938 (N_15938,N_9840,N_9307);
or U15939 (N_15939,N_9541,N_1793);
and U15940 (N_15940,N_553,N_2342);
nand U15941 (N_15941,N_577,N_2912);
or U15942 (N_15942,N_7299,N_6798);
and U15943 (N_15943,N_6744,N_9569);
nand U15944 (N_15944,N_4551,N_6259);
or U15945 (N_15945,N_77,N_8076);
nor U15946 (N_15946,N_7770,N_9091);
nor U15947 (N_15947,N_6538,N_9653);
nand U15948 (N_15948,N_5362,N_8148);
and U15949 (N_15949,N_7332,N_1023);
or U15950 (N_15950,N_5698,N_371);
nand U15951 (N_15951,N_1155,N_9451);
and U15952 (N_15952,N_5893,N_3354);
and U15953 (N_15953,N_100,N_8238);
or U15954 (N_15954,N_8551,N_6166);
nand U15955 (N_15955,N_6466,N_4766);
nor U15956 (N_15956,N_6709,N_4865);
xor U15957 (N_15957,N_8943,N_8843);
nand U15958 (N_15958,N_4774,N_5317);
and U15959 (N_15959,N_6882,N_2352);
or U15960 (N_15960,N_4134,N_5176);
and U15961 (N_15961,N_8372,N_3737);
and U15962 (N_15962,N_3633,N_5829);
nand U15963 (N_15963,N_1984,N_8307);
and U15964 (N_15964,N_5725,N_4110);
nand U15965 (N_15965,N_9238,N_2523);
or U15966 (N_15966,N_1190,N_3669);
xnor U15967 (N_15967,N_2015,N_1741);
nand U15968 (N_15968,N_3305,N_2591);
nor U15969 (N_15969,N_9012,N_594);
and U15970 (N_15970,N_808,N_3022);
or U15971 (N_15971,N_1257,N_1900);
nor U15972 (N_15972,N_2947,N_6258);
nor U15973 (N_15973,N_5743,N_8621);
nor U15974 (N_15974,N_3566,N_3511);
xnor U15975 (N_15975,N_2595,N_6528);
nand U15976 (N_15976,N_5772,N_9700);
nor U15977 (N_15977,N_901,N_5640);
nand U15978 (N_15978,N_4151,N_6066);
nor U15979 (N_15979,N_3998,N_5396);
nand U15980 (N_15980,N_8652,N_2107);
xnor U15981 (N_15981,N_5395,N_2991);
and U15982 (N_15982,N_3743,N_5321);
nor U15983 (N_15983,N_7405,N_9714);
nor U15984 (N_15984,N_4324,N_110);
or U15985 (N_15985,N_7800,N_2352);
nand U15986 (N_15986,N_2227,N_3994);
or U15987 (N_15987,N_4077,N_9063);
or U15988 (N_15988,N_200,N_2048);
or U15989 (N_15989,N_764,N_5643);
and U15990 (N_15990,N_5292,N_6935);
nand U15991 (N_15991,N_1638,N_7958);
nor U15992 (N_15992,N_6012,N_5331);
or U15993 (N_15993,N_7455,N_6826);
nor U15994 (N_15994,N_9964,N_488);
and U15995 (N_15995,N_7721,N_845);
and U15996 (N_15996,N_4923,N_471);
nand U15997 (N_15997,N_1964,N_9783);
nor U15998 (N_15998,N_9993,N_4793);
xnor U15999 (N_15999,N_6928,N_5555);
nand U16000 (N_16000,N_234,N_1294);
or U16001 (N_16001,N_2526,N_8250);
or U16002 (N_16002,N_3920,N_6273);
nand U16003 (N_16003,N_9510,N_3560);
or U16004 (N_16004,N_522,N_7622);
and U16005 (N_16005,N_4004,N_5220);
or U16006 (N_16006,N_4601,N_9400);
nand U16007 (N_16007,N_1494,N_7379);
and U16008 (N_16008,N_228,N_2602);
and U16009 (N_16009,N_9393,N_6712);
nor U16010 (N_16010,N_411,N_8241);
nor U16011 (N_16011,N_1433,N_3574);
nand U16012 (N_16012,N_7920,N_4337);
nor U16013 (N_16013,N_101,N_1856);
or U16014 (N_16014,N_4128,N_5136);
nand U16015 (N_16015,N_4924,N_5520);
nor U16016 (N_16016,N_6365,N_328);
nor U16017 (N_16017,N_73,N_4318);
nand U16018 (N_16018,N_7994,N_371);
or U16019 (N_16019,N_3409,N_3870);
nand U16020 (N_16020,N_8308,N_3140);
nand U16021 (N_16021,N_7592,N_3423);
and U16022 (N_16022,N_5283,N_3084);
nor U16023 (N_16023,N_6088,N_5609);
nand U16024 (N_16024,N_1583,N_9432);
nor U16025 (N_16025,N_4075,N_1131);
or U16026 (N_16026,N_4548,N_3594);
nor U16027 (N_16027,N_1517,N_7394);
and U16028 (N_16028,N_4056,N_7508);
and U16029 (N_16029,N_4892,N_9015);
and U16030 (N_16030,N_5735,N_4316);
and U16031 (N_16031,N_2414,N_8529);
xor U16032 (N_16032,N_3211,N_7910);
nor U16033 (N_16033,N_6684,N_988);
or U16034 (N_16034,N_6063,N_7493);
nand U16035 (N_16035,N_2005,N_5037);
nor U16036 (N_16036,N_7597,N_3197);
xor U16037 (N_16037,N_6577,N_2078);
nor U16038 (N_16038,N_8802,N_2764);
xor U16039 (N_16039,N_4463,N_582);
nor U16040 (N_16040,N_615,N_7839);
nor U16041 (N_16041,N_4629,N_7128);
xor U16042 (N_16042,N_7125,N_285);
or U16043 (N_16043,N_6422,N_6290);
nand U16044 (N_16044,N_7932,N_4713);
nor U16045 (N_16045,N_6428,N_6457);
nand U16046 (N_16046,N_6308,N_3585);
nand U16047 (N_16047,N_2478,N_2492);
nand U16048 (N_16048,N_6166,N_1498);
and U16049 (N_16049,N_9449,N_3279);
nand U16050 (N_16050,N_3212,N_1102);
xor U16051 (N_16051,N_6376,N_3234);
nor U16052 (N_16052,N_6264,N_4443);
and U16053 (N_16053,N_4574,N_7232);
nand U16054 (N_16054,N_4556,N_6580);
nand U16055 (N_16055,N_4769,N_9702);
xnor U16056 (N_16056,N_8250,N_5974);
xnor U16057 (N_16057,N_9227,N_419);
nand U16058 (N_16058,N_5555,N_1149);
nand U16059 (N_16059,N_1467,N_2097);
or U16060 (N_16060,N_9463,N_7537);
nand U16061 (N_16061,N_1384,N_3966);
and U16062 (N_16062,N_2216,N_2392);
and U16063 (N_16063,N_1009,N_6971);
or U16064 (N_16064,N_3301,N_609);
or U16065 (N_16065,N_6627,N_6483);
nor U16066 (N_16066,N_7176,N_2138);
nor U16067 (N_16067,N_3030,N_3335);
and U16068 (N_16068,N_4607,N_9615);
nand U16069 (N_16069,N_4056,N_2099);
and U16070 (N_16070,N_7355,N_9171);
and U16071 (N_16071,N_1892,N_8684);
xor U16072 (N_16072,N_4449,N_577);
or U16073 (N_16073,N_6903,N_4945);
nand U16074 (N_16074,N_6833,N_5082);
and U16075 (N_16075,N_6907,N_6487);
and U16076 (N_16076,N_9013,N_712);
xor U16077 (N_16077,N_3922,N_3340);
nand U16078 (N_16078,N_4232,N_9639);
and U16079 (N_16079,N_147,N_6992);
or U16080 (N_16080,N_4103,N_7350);
xnor U16081 (N_16081,N_7326,N_8468);
nand U16082 (N_16082,N_1946,N_3563);
nor U16083 (N_16083,N_2252,N_260);
nand U16084 (N_16084,N_3908,N_8350);
xnor U16085 (N_16085,N_9461,N_8753);
nor U16086 (N_16086,N_4396,N_1636);
nand U16087 (N_16087,N_2160,N_1999);
or U16088 (N_16088,N_4425,N_2691);
or U16089 (N_16089,N_5686,N_9789);
and U16090 (N_16090,N_4827,N_4789);
and U16091 (N_16091,N_3697,N_7083);
or U16092 (N_16092,N_324,N_9315);
or U16093 (N_16093,N_7205,N_6987);
or U16094 (N_16094,N_3483,N_6970);
nand U16095 (N_16095,N_965,N_5986);
and U16096 (N_16096,N_5456,N_4871);
xor U16097 (N_16097,N_6310,N_1593);
xnor U16098 (N_16098,N_5648,N_3801);
and U16099 (N_16099,N_5812,N_2913);
nand U16100 (N_16100,N_7087,N_9087);
xor U16101 (N_16101,N_7130,N_9743);
or U16102 (N_16102,N_4631,N_7545);
nor U16103 (N_16103,N_2223,N_9798);
xnor U16104 (N_16104,N_1086,N_7544);
nand U16105 (N_16105,N_1795,N_6208);
nand U16106 (N_16106,N_8006,N_4267);
or U16107 (N_16107,N_5742,N_3477);
or U16108 (N_16108,N_5361,N_3066);
nand U16109 (N_16109,N_7193,N_5297);
and U16110 (N_16110,N_2484,N_6872);
xor U16111 (N_16111,N_5575,N_4448);
nand U16112 (N_16112,N_4267,N_6053);
nand U16113 (N_16113,N_16,N_9333);
and U16114 (N_16114,N_2377,N_2023);
or U16115 (N_16115,N_2865,N_4191);
nand U16116 (N_16116,N_5586,N_199);
xnor U16117 (N_16117,N_9794,N_7463);
nor U16118 (N_16118,N_9498,N_4260);
or U16119 (N_16119,N_1499,N_286);
or U16120 (N_16120,N_6577,N_4281);
nand U16121 (N_16121,N_6123,N_7838);
and U16122 (N_16122,N_171,N_9320);
nor U16123 (N_16123,N_6086,N_9793);
and U16124 (N_16124,N_1600,N_8576);
nor U16125 (N_16125,N_1050,N_3209);
nor U16126 (N_16126,N_9465,N_4516);
and U16127 (N_16127,N_1855,N_5187);
or U16128 (N_16128,N_4231,N_3019);
or U16129 (N_16129,N_8807,N_3383);
nor U16130 (N_16130,N_2043,N_4104);
or U16131 (N_16131,N_3869,N_3969);
or U16132 (N_16132,N_3580,N_8841);
or U16133 (N_16133,N_713,N_5805);
nand U16134 (N_16134,N_7230,N_5760);
xnor U16135 (N_16135,N_5326,N_2108);
and U16136 (N_16136,N_1380,N_4158);
and U16137 (N_16137,N_9619,N_9614);
and U16138 (N_16138,N_7527,N_3304);
or U16139 (N_16139,N_3955,N_2704);
nand U16140 (N_16140,N_802,N_4510);
or U16141 (N_16141,N_5636,N_1187);
nor U16142 (N_16142,N_1512,N_1719);
or U16143 (N_16143,N_2429,N_2055);
nand U16144 (N_16144,N_8654,N_2376);
nand U16145 (N_16145,N_3120,N_838);
nor U16146 (N_16146,N_3839,N_7423);
or U16147 (N_16147,N_3061,N_1244);
nor U16148 (N_16148,N_4182,N_8836);
nor U16149 (N_16149,N_855,N_2650);
or U16150 (N_16150,N_3228,N_755);
or U16151 (N_16151,N_2256,N_6440);
nor U16152 (N_16152,N_3657,N_5945);
and U16153 (N_16153,N_4468,N_3402);
and U16154 (N_16154,N_994,N_638);
or U16155 (N_16155,N_7376,N_542);
nand U16156 (N_16156,N_2848,N_1247);
nor U16157 (N_16157,N_23,N_4213);
or U16158 (N_16158,N_334,N_292);
and U16159 (N_16159,N_4613,N_1281);
nand U16160 (N_16160,N_2794,N_8773);
nand U16161 (N_16161,N_7861,N_2689);
nand U16162 (N_16162,N_2114,N_9694);
or U16163 (N_16163,N_9597,N_8252);
and U16164 (N_16164,N_783,N_200);
xnor U16165 (N_16165,N_5352,N_6454);
and U16166 (N_16166,N_9940,N_2384);
xor U16167 (N_16167,N_639,N_8067);
nor U16168 (N_16168,N_7466,N_1688);
or U16169 (N_16169,N_6607,N_8649);
nor U16170 (N_16170,N_6951,N_3924);
nand U16171 (N_16171,N_9344,N_7451);
or U16172 (N_16172,N_5051,N_8525);
or U16173 (N_16173,N_9304,N_1725);
xnor U16174 (N_16174,N_8381,N_1574);
or U16175 (N_16175,N_2236,N_5487);
nor U16176 (N_16176,N_4236,N_2301);
nor U16177 (N_16177,N_8662,N_5793);
nor U16178 (N_16178,N_9271,N_3587);
nand U16179 (N_16179,N_7113,N_474);
xnor U16180 (N_16180,N_4889,N_4137);
and U16181 (N_16181,N_1597,N_1862);
or U16182 (N_16182,N_7087,N_5525);
and U16183 (N_16183,N_6972,N_4971);
nand U16184 (N_16184,N_2886,N_921);
and U16185 (N_16185,N_829,N_4743);
or U16186 (N_16186,N_8711,N_3903);
nor U16187 (N_16187,N_3274,N_3358);
nand U16188 (N_16188,N_417,N_7933);
and U16189 (N_16189,N_7890,N_6503);
nor U16190 (N_16190,N_8647,N_4025);
and U16191 (N_16191,N_9641,N_4845);
nor U16192 (N_16192,N_1048,N_5466);
nand U16193 (N_16193,N_4666,N_9625);
or U16194 (N_16194,N_9891,N_29);
nand U16195 (N_16195,N_3776,N_9802);
or U16196 (N_16196,N_5017,N_3587);
nor U16197 (N_16197,N_4470,N_7779);
nor U16198 (N_16198,N_1162,N_8900);
nand U16199 (N_16199,N_2787,N_7156);
nor U16200 (N_16200,N_8792,N_9427);
nand U16201 (N_16201,N_964,N_2350);
and U16202 (N_16202,N_1885,N_316);
or U16203 (N_16203,N_5942,N_1329);
nor U16204 (N_16204,N_1553,N_721);
and U16205 (N_16205,N_4207,N_8324);
nand U16206 (N_16206,N_8531,N_449);
nor U16207 (N_16207,N_9850,N_1342);
nand U16208 (N_16208,N_2286,N_93);
xnor U16209 (N_16209,N_3331,N_7801);
or U16210 (N_16210,N_7104,N_6165);
or U16211 (N_16211,N_5114,N_3441);
nand U16212 (N_16212,N_5984,N_6890);
nor U16213 (N_16213,N_5185,N_2684);
nand U16214 (N_16214,N_9587,N_5295);
or U16215 (N_16215,N_2892,N_3157);
and U16216 (N_16216,N_622,N_9262);
and U16217 (N_16217,N_571,N_1901);
nor U16218 (N_16218,N_4076,N_1889);
nor U16219 (N_16219,N_389,N_6447);
or U16220 (N_16220,N_2705,N_966);
and U16221 (N_16221,N_6926,N_9599);
and U16222 (N_16222,N_7192,N_2316);
nor U16223 (N_16223,N_4176,N_4124);
and U16224 (N_16224,N_8851,N_9362);
and U16225 (N_16225,N_7213,N_8103);
or U16226 (N_16226,N_6129,N_3575);
nor U16227 (N_16227,N_1180,N_3603);
nand U16228 (N_16228,N_847,N_8486);
nor U16229 (N_16229,N_1352,N_9395);
or U16230 (N_16230,N_9016,N_6152);
or U16231 (N_16231,N_2215,N_7707);
nand U16232 (N_16232,N_5082,N_4628);
or U16233 (N_16233,N_6176,N_6655);
and U16234 (N_16234,N_4541,N_5436);
and U16235 (N_16235,N_7943,N_8424);
or U16236 (N_16236,N_5736,N_4703);
nand U16237 (N_16237,N_9954,N_5475);
or U16238 (N_16238,N_6392,N_2914);
and U16239 (N_16239,N_3296,N_9120);
and U16240 (N_16240,N_5045,N_8383);
nand U16241 (N_16241,N_4390,N_6697);
and U16242 (N_16242,N_2776,N_8414);
nor U16243 (N_16243,N_8110,N_310);
and U16244 (N_16244,N_4472,N_9734);
nor U16245 (N_16245,N_9969,N_212);
nand U16246 (N_16246,N_7249,N_4515);
nand U16247 (N_16247,N_2740,N_2750);
nor U16248 (N_16248,N_1343,N_9483);
and U16249 (N_16249,N_9669,N_3399);
nor U16250 (N_16250,N_8245,N_9055);
xnor U16251 (N_16251,N_7856,N_2040);
and U16252 (N_16252,N_351,N_3942);
and U16253 (N_16253,N_7680,N_3832);
xor U16254 (N_16254,N_9601,N_4941);
or U16255 (N_16255,N_743,N_4000);
or U16256 (N_16256,N_8771,N_4711);
or U16257 (N_16257,N_4158,N_4299);
nand U16258 (N_16258,N_3381,N_7618);
or U16259 (N_16259,N_2860,N_3093);
xor U16260 (N_16260,N_8649,N_4146);
nor U16261 (N_16261,N_1624,N_5718);
nor U16262 (N_16262,N_4051,N_3804);
and U16263 (N_16263,N_3723,N_9153);
or U16264 (N_16264,N_5091,N_7448);
nand U16265 (N_16265,N_1059,N_9869);
and U16266 (N_16266,N_4916,N_228);
or U16267 (N_16267,N_5373,N_391);
and U16268 (N_16268,N_6368,N_3677);
or U16269 (N_16269,N_8940,N_5016);
or U16270 (N_16270,N_3691,N_409);
nor U16271 (N_16271,N_7782,N_6140);
or U16272 (N_16272,N_7412,N_1511);
nand U16273 (N_16273,N_9019,N_7966);
and U16274 (N_16274,N_7495,N_1708);
nand U16275 (N_16275,N_2212,N_3569);
nor U16276 (N_16276,N_6677,N_4101);
or U16277 (N_16277,N_7754,N_351);
or U16278 (N_16278,N_7759,N_8714);
nor U16279 (N_16279,N_1790,N_9774);
and U16280 (N_16280,N_4031,N_4238);
nand U16281 (N_16281,N_5522,N_7916);
or U16282 (N_16282,N_1835,N_9359);
and U16283 (N_16283,N_2313,N_3668);
and U16284 (N_16284,N_7115,N_5304);
nand U16285 (N_16285,N_8488,N_1917);
or U16286 (N_16286,N_6681,N_7938);
and U16287 (N_16287,N_5678,N_8811);
nand U16288 (N_16288,N_9843,N_4613);
or U16289 (N_16289,N_8980,N_8569);
or U16290 (N_16290,N_352,N_3030);
or U16291 (N_16291,N_1060,N_5186);
and U16292 (N_16292,N_8052,N_6022);
and U16293 (N_16293,N_2960,N_5242);
or U16294 (N_16294,N_1877,N_1224);
or U16295 (N_16295,N_9297,N_9338);
or U16296 (N_16296,N_1014,N_2349);
nor U16297 (N_16297,N_5181,N_4343);
and U16298 (N_16298,N_8408,N_1800);
nand U16299 (N_16299,N_8302,N_2231);
or U16300 (N_16300,N_5232,N_9757);
xor U16301 (N_16301,N_6169,N_8967);
and U16302 (N_16302,N_332,N_1592);
nand U16303 (N_16303,N_7098,N_1766);
and U16304 (N_16304,N_2860,N_8809);
and U16305 (N_16305,N_4076,N_2862);
nand U16306 (N_16306,N_702,N_9127);
nand U16307 (N_16307,N_894,N_2848);
or U16308 (N_16308,N_9422,N_3591);
and U16309 (N_16309,N_7724,N_6744);
or U16310 (N_16310,N_4018,N_9211);
or U16311 (N_16311,N_1916,N_4579);
and U16312 (N_16312,N_8292,N_1832);
and U16313 (N_16313,N_2364,N_3733);
nand U16314 (N_16314,N_7642,N_1569);
xor U16315 (N_16315,N_9922,N_5339);
nand U16316 (N_16316,N_8331,N_4769);
xor U16317 (N_16317,N_5817,N_886);
or U16318 (N_16318,N_9291,N_4845);
nand U16319 (N_16319,N_8932,N_5495);
nor U16320 (N_16320,N_663,N_4492);
nor U16321 (N_16321,N_9716,N_7902);
or U16322 (N_16322,N_5378,N_4903);
and U16323 (N_16323,N_5116,N_6765);
nor U16324 (N_16324,N_785,N_5591);
nor U16325 (N_16325,N_3098,N_5391);
or U16326 (N_16326,N_2602,N_6526);
nand U16327 (N_16327,N_931,N_5913);
or U16328 (N_16328,N_9290,N_273);
or U16329 (N_16329,N_9700,N_426);
and U16330 (N_16330,N_6837,N_7559);
or U16331 (N_16331,N_7583,N_6005);
xnor U16332 (N_16332,N_5583,N_1291);
nor U16333 (N_16333,N_3238,N_7958);
xor U16334 (N_16334,N_7214,N_8659);
nand U16335 (N_16335,N_8946,N_7895);
xnor U16336 (N_16336,N_8691,N_3705);
or U16337 (N_16337,N_3174,N_3839);
and U16338 (N_16338,N_2866,N_5502);
or U16339 (N_16339,N_3594,N_6320);
xor U16340 (N_16340,N_7193,N_2901);
and U16341 (N_16341,N_7069,N_7601);
nand U16342 (N_16342,N_1881,N_8169);
nor U16343 (N_16343,N_1953,N_4811);
nand U16344 (N_16344,N_9024,N_7848);
nand U16345 (N_16345,N_4950,N_6985);
nor U16346 (N_16346,N_2312,N_7540);
and U16347 (N_16347,N_2482,N_8360);
nor U16348 (N_16348,N_7064,N_6768);
and U16349 (N_16349,N_4960,N_4232);
or U16350 (N_16350,N_1675,N_3904);
nor U16351 (N_16351,N_9888,N_6417);
and U16352 (N_16352,N_1620,N_5612);
and U16353 (N_16353,N_3473,N_3438);
and U16354 (N_16354,N_6119,N_5446);
nand U16355 (N_16355,N_3251,N_6347);
and U16356 (N_16356,N_1263,N_1722);
nor U16357 (N_16357,N_8119,N_98);
nor U16358 (N_16358,N_2042,N_563);
or U16359 (N_16359,N_8152,N_5423);
nand U16360 (N_16360,N_5487,N_2753);
and U16361 (N_16361,N_2460,N_3135);
and U16362 (N_16362,N_5020,N_4491);
and U16363 (N_16363,N_3403,N_2726);
and U16364 (N_16364,N_8562,N_7982);
or U16365 (N_16365,N_8847,N_43);
xor U16366 (N_16366,N_6231,N_3228);
nand U16367 (N_16367,N_9970,N_3066);
nand U16368 (N_16368,N_5421,N_8934);
and U16369 (N_16369,N_7755,N_398);
nand U16370 (N_16370,N_9353,N_808);
and U16371 (N_16371,N_8465,N_951);
and U16372 (N_16372,N_9325,N_2832);
or U16373 (N_16373,N_3584,N_3150);
and U16374 (N_16374,N_7415,N_7815);
nand U16375 (N_16375,N_5090,N_6272);
nor U16376 (N_16376,N_9157,N_5233);
nand U16377 (N_16377,N_1114,N_168);
and U16378 (N_16378,N_8418,N_1693);
xnor U16379 (N_16379,N_8270,N_4437);
or U16380 (N_16380,N_2338,N_5129);
nand U16381 (N_16381,N_1422,N_7911);
xnor U16382 (N_16382,N_1895,N_199);
xor U16383 (N_16383,N_7183,N_6084);
or U16384 (N_16384,N_6998,N_5002);
or U16385 (N_16385,N_2187,N_3630);
and U16386 (N_16386,N_1395,N_1889);
and U16387 (N_16387,N_1928,N_2124);
nand U16388 (N_16388,N_555,N_2366);
nand U16389 (N_16389,N_3056,N_2504);
or U16390 (N_16390,N_4226,N_1639);
or U16391 (N_16391,N_6941,N_9026);
nand U16392 (N_16392,N_2713,N_8211);
or U16393 (N_16393,N_7888,N_8418);
nor U16394 (N_16394,N_2329,N_5438);
nor U16395 (N_16395,N_8362,N_4278);
xor U16396 (N_16396,N_3205,N_238);
nand U16397 (N_16397,N_5583,N_5248);
and U16398 (N_16398,N_9022,N_9110);
xor U16399 (N_16399,N_1043,N_6713);
nand U16400 (N_16400,N_4449,N_7307);
nor U16401 (N_16401,N_8286,N_2438);
nand U16402 (N_16402,N_4208,N_2608);
xor U16403 (N_16403,N_6978,N_6960);
nand U16404 (N_16404,N_568,N_8936);
xnor U16405 (N_16405,N_1960,N_7999);
xor U16406 (N_16406,N_5025,N_8435);
nor U16407 (N_16407,N_4762,N_1114);
xor U16408 (N_16408,N_1154,N_8906);
xnor U16409 (N_16409,N_1938,N_1194);
nor U16410 (N_16410,N_699,N_6127);
nor U16411 (N_16411,N_9819,N_2490);
or U16412 (N_16412,N_4825,N_5815);
or U16413 (N_16413,N_7622,N_7275);
nor U16414 (N_16414,N_1623,N_7328);
nand U16415 (N_16415,N_8602,N_348);
nand U16416 (N_16416,N_6503,N_4562);
nor U16417 (N_16417,N_5512,N_4606);
nand U16418 (N_16418,N_983,N_7888);
xor U16419 (N_16419,N_7480,N_7926);
nor U16420 (N_16420,N_421,N_4312);
and U16421 (N_16421,N_3202,N_9424);
and U16422 (N_16422,N_9493,N_6167);
nor U16423 (N_16423,N_8060,N_3441);
xor U16424 (N_16424,N_8791,N_5433);
and U16425 (N_16425,N_7375,N_6916);
and U16426 (N_16426,N_4974,N_8081);
or U16427 (N_16427,N_9180,N_6741);
nand U16428 (N_16428,N_4672,N_6062);
and U16429 (N_16429,N_3107,N_1631);
or U16430 (N_16430,N_9860,N_1159);
xor U16431 (N_16431,N_6429,N_9726);
and U16432 (N_16432,N_4238,N_7114);
and U16433 (N_16433,N_7433,N_2227);
nand U16434 (N_16434,N_3938,N_1314);
and U16435 (N_16435,N_4449,N_227);
and U16436 (N_16436,N_6716,N_6537);
or U16437 (N_16437,N_1475,N_5324);
nor U16438 (N_16438,N_4896,N_6712);
or U16439 (N_16439,N_2703,N_451);
nor U16440 (N_16440,N_9107,N_6930);
or U16441 (N_16441,N_3465,N_1986);
or U16442 (N_16442,N_5458,N_8061);
nor U16443 (N_16443,N_5841,N_1681);
nand U16444 (N_16444,N_3875,N_1195);
nor U16445 (N_16445,N_9404,N_3544);
and U16446 (N_16446,N_9091,N_1452);
nand U16447 (N_16447,N_823,N_8801);
nand U16448 (N_16448,N_2627,N_6095);
or U16449 (N_16449,N_3586,N_11);
or U16450 (N_16450,N_4798,N_8308);
or U16451 (N_16451,N_1141,N_7424);
and U16452 (N_16452,N_6080,N_5558);
nor U16453 (N_16453,N_5801,N_3824);
nand U16454 (N_16454,N_734,N_1257);
or U16455 (N_16455,N_9409,N_4226);
or U16456 (N_16456,N_7824,N_6422);
nand U16457 (N_16457,N_2858,N_3545);
nand U16458 (N_16458,N_7774,N_7455);
or U16459 (N_16459,N_6011,N_1754);
nor U16460 (N_16460,N_2514,N_508);
or U16461 (N_16461,N_885,N_3605);
or U16462 (N_16462,N_2379,N_9489);
nor U16463 (N_16463,N_4980,N_6745);
and U16464 (N_16464,N_3077,N_1063);
or U16465 (N_16465,N_3709,N_3582);
or U16466 (N_16466,N_8501,N_3558);
or U16467 (N_16467,N_7427,N_7572);
nand U16468 (N_16468,N_9243,N_7975);
or U16469 (N_16469,N_5609,N_5376);
and U16470 (N_16470,N_3795,N_8308);
and U16471 (N_16471,N_1321,N_5346);
nand U16472 (N_16472,N_6442,N_6961);
or U16473 (N_16473,N_6751,N_3550);
or U16474 (N_16474,N_8593,N_8295);
nand U16475 (N_16475,N_2900,N_5335);
or U16476 (N_16476,N_8401,N_9448);
and U16477 (N_16477,N_3003,N_2496);
or U16478 (N_16478,N_7829,N_5083);
or U16479 (N_16479,N_5838,N_4070);
xnor U16480 (N_16480,N_4480,N_3604);
and U16481 (N_16481,N_2263,N_1530);
nor U16482 (N_16482,N_2273,N_4477);
and U16483 (N_16483,N_5751,N_9120);
nor U16484 (N_16484,N_2389,N_2936);
nand U16485 (N_16485,N_2291,N_7274);
nor U16486 (N_16486,N_9295,N_6850);
and U16487 (N_16487,N_7555,N_5410);
and U16488 (N_16488,N_3197,N_8260);
or U16489 (N_16489,N_5616,N_2451);
nand U16490 (N_16490,N_5662,N_2550);
or U16491 (N_16491,N_2608,N_7634);
nand U16492 (N_16492,N_6686,N_4197);
nor U16493 (N_16493,N_2637,N_57);
or U16494 (N_16494,N_6307,N_7581);
and U16495 (N_16495,N_1308,N_2555);
nand U16496 (N_16496,N_3376,N_5811);
or U16497 (N_16497,N_321,N_919);
nand U16498 (N_16498,N_4012,N_6502);
nand U16499 (N_16499,N_1567,N_7431);
nand U16500 (N_16500,N_8304,N_1897);
or U16501 (N_16501,N_3560,N_5486);
or U16502 (N_16502,N_8551,N_2193);
nor U16503 (N_16503,N_8646,N_4109);
nand U16504 (N_16504,N_7116,N_7531);
nor U16505 (N_16505,N_865,N_4940);
nor U16506 (N_16506,N_2717,N_2148);
nand U16507 (N_16507,N_2553,N_2708);
and U16508 (N_16508,N_8263,N_7515);
or U16509 (N_16509,N_9864,N_2564);
nor U16510 (N_16510,N_7948,N_3335);
nand U16511 (N_16511,N_4415,N_8384);
or U16512 (N_16512,N_8082,N_8065);
xor U16513 (N_16513,N_8427,N_7669);
nand U16514 (N_16514,N_4571,N_3374);
or U16515 (N_16515,N_1770,N_3063);
and U16516 (N_16516,N_1969,N_6677);
and U16517 (N_16517,N_3584,N_8332);
nand U16518 (N_16518,N_4311,N_7303);
nor U16519 (N_16519,N_4066,N_4737);
or U16520 (N_16520,N_6168,N_2787);
and U16521 (N_16521,N_4127,N_8451);
or U16522 (N_16522,N_20,N_1172);
xnor U16523 (N_16523,N_4532,N_9459);
nor U16524 (N_16524,N_1627,N_8287);
nand U16525 (N_16525,N_4651,N_4483);
or U16526 (N_16526,N_2626,N_1678);
nand U16527 (N_16527,N_7879,N_5007);
or U16528 (N_16528,N_606,N_3094);
nor U16529 (N_16529,N_1039,N_4536);
and U16530 (N_16530,N_5678,N_2244);
xor U16531 (N_16531,N_5297,N_896);
or U16532 (N_16532,N_9901,N_1674);
or U16533 (N_16533,N_4876,N_1810);
or U16534 (N_16534,N_4049,N_6805);
nor U16535 (N_16535,N_8693,N_8100);
or U16536 (N_16536,N_5453,N_8972);
nand U16537 (N_16537,N_9319,N_7697);
xor U16538 (N_16538,N_8243,N_7904);
nand U16539 (N_16539,N_3924,N_4494);
nor U16540 (N_16540,N_8271,N_5787);
or U16541 (N_16541,N_6197,N_7740);
nor U16542 (N_16542,N_3098,N_8040);
or U16543 (N_16543,N_1966,N_633);
and U16544 (N_16544,N_7558,N_5347);
nor U16545 (N_16545,N_8263,N_6066);
xnor U16546 (N_16546,N_8961,N_4544);
or U16547 (N_16547,N_8698,N_3407);
or U16548 (N_16548,N_9637,N_7088);
nor U16549 (N_16549,N_1911,N_5865);
nor U16550 (N_16550,N_7006,N_3446);
or U16551 (N_16551,N_2746,N_3800);
or U16552 (N_16552,N_4522,N_8921);
nor U16553 (N_16553,N_940,N_2222);
and U16554 (N_16554,N_5985,N_1795);
xor U16555 (N_16555,N_1990,N_7009);
and U16556 (N_16556,N_8183,N_4661);
xnor U16557 (N_16557,N_8436,N_3129);
xnor U16558 (N_16558,N_8934,N_7903);
nor U16559 (N_16559,N_1434,N_8904);
nand U16560 (N_16560,N_534,N_3723);
nor U16561 (N_16561,N_3811,N_8888);
nand U16562 (N_16562,N_8490,N_4625);
nor U16563 (N_16563,N_6948,N_4769);
and U16564 (N_16564,N_3548,N_3278);
nand U16565 (N_16565,N_5842,N_4955);
and U16566 (N_16566,N_8113,N_7104);
nor U16567 (N_16567,N_7045,N_5905);
xnor U16568 (N_16568,N_5765,N_744);
xor U16569 (N_16569,N_9216,N_1061);
and U16570 (N_16570,N_5069,N_9636);
or U16571 (N_16571,N_764,N_197);
nand U16572 (N_16572,N_7358,N_6261);
nand U16573 (N_16573,N_5633,N_6784);
or U16574 (N_16574,N_8278,N_4865);
or U16575 (N_16575,N_8824,N_2233);
nor U16576 (N_16576,N_8362,N_6512);
xnor U16577 (N_16577,N_7298,N_1900);
nand U16578 (N_16578,N_8066,N_8685);
and U16579 (N_16579,N_25,N_2090);
and U16580 (N_16580,N_7826,N_787);
or U16581 (N_16581,N_149,N_3392);
nor U16582 (N_16582,N_824,N_7071);
or U16583 (N_16583,N_86,N_2009);
and U16584 (N_16584,N_8056,N_1281);
nor U16585 (N_16585,N_6160,N_8407);
or U16586 (N_16586,N_4615,N_9816);
or U16587 (N_16587,N_9050,N_3630);
or U16588 (N_16588,N_6896,N_4386);
nor U16589 (N_16589,N_5432,N_3692);
and U16590 (N_16590,N_7023,N_3297);
nand U16591 (N_16591,N_1286,N_8272);
nand U16592 (N_16592,N_158,N_8186);
or U16593 (N_16593,N_2987,N_8911);
nor U16594 (N_16594,N_8942,N_6545);
or U16595 (N_16595,N_536,N_8466);
or U16596 (N_16596,N_7954,N_1560);
xnor U16597 (N_16597,N_6236,N_9203);
and U16598 (N_16598,N_8707,N_5766);
and U16599 (N_16599,N_4506,N_7113);
nor U16600 (N_16600,N_4392,N_8087);
or U16601 (N_16601,N_1258,N_2956);
nand U16602 (N_16602,N_3388,N_1598);
or U16603 (N_16603,N_1467,N_5912);
nor U16604 (N_16604,N_9375,N_9416);
nand U16605 (N_16605,N_2851,N_6328);
nand U16606 (N_16606,N_6305,N_7039);
and U16607 (N_16607,N_9188,N_632);
nor U16608 (N_16608,N_4668,N_4080);
xnor U16609 (N_16609,N_9343,N_1621);
nand U16610 (N_16610,N_1287,N_9678);
nand U16611 (N_16611,N_9968,N_9777);
or U16612 (N_16612,N_5379,N_5752);
nor U16613 (N_16613,N_1349,N_5202);
nor U16614 (N_16614,N_2769,N_8525);
xnor U16615 (N_16615,N_1980,N_5333);
xor U16616 (N_16616,N_463,N_3832);
and U16617 (N_16617,N_7424,N_5153);
nand U16618 (N_16618,N_505,N_595);
xor U16619 (N_16619,N_0,N_9182);
nand U16620 (N_16620,N_324,N_5198);
nand U16621 (N_16621,N_5280,N_4417);
nor U16622 (N_16622,N_2843,N_3050);
nor U16623 (N_16623,N_3405,N_9546);
or U16624 (N_16624,N_5746,N_5461);
xor U16625 (N_16625,N_580,N_6332);
or U16626 (N_16626,N_4884,N_9528);
or U16627 (N_16627,N_3614,N_2840);
nor U16628 (N_16628,N_4382,N_6229);
nor U16629 (N_16629,N_9544,N_8);
or U16630 (N_16630,N_2002,N_5530);
xor U16631 (N_16631,N_1317,N_3219);
nor U16632 (N_16632,N_2955,N_3929);
or U16633 (N_16633,N_4583,N_3211);
nor U16634 (N_16634,N_8104,N_2456);
nor U16635 (N_16635,N_2302,N_788);
nand U16636 (N_16636,N_9061,N_5321);
or U16637 (N_16637,N_6372,N_9031);
and U16638 (N_16638,N_332,N_2212);
nor U16639 (N_16639,N_3262,N_2978);
or U16640 (N_16640,N_5299,N_3024);
xnor U16641 (N_16641,N_7592,N_1500);
nor U16642 (N_16642,N_2765,N_6092);
xnor U16643 (N_16643,N_8766,N_7329);
and U16644 (N_16644,N_436,N_1176);
nand U16645 (N_16645,N_6865,N_7543);
nand U16646 (N_16646,N_9988,N_3206);
or U16647 (N_16647,N_5876,N_438);
or U16648 (N_16648,N_8424,N_1056);
and U16649 (N_16649,N_8794,N_5918);
nand U16650 (N_16650,N_3043,N_5910);
nor U16651 (N_16651,N_9382,N_2556);
and U16652 (N_16652,N_2598,N_7839);
or U16653 (N_16653,N_7478,N_3718);
nor U16654 (N_16654,N_5197,N_2745);
and U16655 (N_16655,N_5563,N_5808);
nand U16656 (N_16656,N_6741,N_5102);
and U16657 (N_16657,N_6554,N_8896);
or U16658 (N_16658,N_9511,N_5287);
nor U16659 (N_16659,N_9578,N_9243);
or U16660 (N_16660,N_4679,N_2085);
xor U16661 (N_16661,N_9881,N_5225);
and U16662 (N_16662,N_9660,N_5889);
nor U16663 (N_16663,N_7373,N_2342);
xor U16664 (N_16664,N_5463,N_8061);
nor U16665 (N_16665,N_4409,N_6315);
or U16666 (N_16666,N_4095,N_8888);
and U16667 (N_16667,N_1077,N_8054);
nand U16668 (N_16668,N_1031,N_2503);
nand U16669 (N_16669,N_4403,N_6792);
nor U16670 (N_16670,N_3584,N_5596);
nand U16671 (N_16671,N_6659,N_5936);
nand U16672 (N_16672,N_4729,N_4100);
nor U16673 (N_16673,N_761,N_1561);
or U16674 (N_16674,N_1768,N_7733);
xor U16675 (N_16675,N_3611,N_2574);
or U16676 (N_16676,N_2705,N_9577);
or U16677 (N_16677,N_9935,N_9941);
and U16678 (N_16678,N_7550,N_972);
nand U16679 (N_16679,N_5205,N_7304);
and U16680 (N_16680,N_1099,N_9555);
and U16681 (N_16681,N_310,N_4531);
nor U16682 (N_16682,N_7802,N_8753);
or U16683 (N_16683,N_1508,N_1567);
nand U16684 (N_16684,N_706,N_1273);
or U16685 (N_16685,N_5058,N_9660);
nand U16686 (N_16686,N_1289,N_1602);
or U16687 (N_16687,N_2063,N_2492);
xnor U16688 (N_16688,N_7220,N_1999);
xnor U16689 (N_16689,N_8797,N_8891);
nand U16690 (N_16690,N_3759,N_2150);
or U16691 (N_16691,N_7232,N_1263);
nor U16692 (N_16692,N_924,N_9802);
or U16693 (N_16693,N_2400,N_7709);
nor U16694 (N_16694,N_4497,N_4696);
or U16695 (N_16695,N_7177,N_607);
and U16696 (N_16696,N_3857,N_7559);
or U16697 (N_16697,N_8457,N_8085);
or U16698 (N_16698,N_8438,N_5557);
or U16699 (N_16699,N_2514,N_2924);
and U16700 (N_16700,N_7569,N_3383);
nand U16701 (N_16701,N_1041,N_2568);
or U16702 (N_16702,N_606,N_3083);
nor U16703 (N_16703,N_981,N_1289);
nor U16704 (N_16704,N_941,N_7641);
and U16705 (N_16705,N_8896,N_9789);
nor U16706 (N_16706,N_8411,N_378);
xor U16707 (N_16707,N_1526,N_3794);
or U16708 (N_16708,N_5788,N_6834);
and U16709 (N_16709,N_2675,N_8776);
or U16710 (N_16710,N_4324,N_8192);
and U16711 (N_16711,N_4259,N_3544);
nand U16712 (N_16712,N_8243,N_3816);
xor U16713 (N_16713,N_1407,N_7884);
and U16714 (N_16714,N_4903,N_3399);
nand U16715 (N_16715,N_3317,N_7471);
nand U16716 (N_16716,N_4222,N_3190);
or U16717 (N_16717,N_4824,N_9130);
xor U16718 (N_16718,N_2356,N_7798);
nor U16719 (N_16719,N_2549,N_245);
and U16720 (N_16720,N_6495,N_4589);
or U16721 (N_16721,N_3009,N_5590);
xor U16722 (N_16722,N_6770,N_9773);
nor U16723 (N_16723,N_4454,N_5994);
nand U16724 (N_16724,N_6170,N_9060);
or U16725 (N_16725,N_7580,N_5286);
nand U16726 (N_16726,N_2999,N_6076);
xor U16727 (N_16727,N_1425,N_9337);
nor U16728 (N_16728,N_605,N_8230);
xnor U16729 (N_16729,N_201,N_6121);
nand U16730 (N_16730,N_4671,N_4397);
nand U16731 (N_16731,N_8145,N_838);
nor U16732 (N_16732,N_9003,N_9610);
and U16733 (N_16733,N_4263,N_4325);
and U16734 (N_16734,N_119,N_1388);
nor U16735 (N_16735,N_1521,N_1771);
nand U16736 (N_16736,N_2510,N_1203);
nor U16737 (N_16737,N_1662,N_8070);
nor U16738 (N_16738,N_4486,N_9718);
or U16739 (N_16739,N_5016,N_2351);
nor U16740 (N_16740,N_1339,N_5371);
and U16741 (N_16741,N_2556,N_4475);
and U16742 (N_16742,N_7342,N_2680);
and U16743 (N_16743,N_7672,N_381);
or U16744 (N_16744,N_396,N_1451);
nand U16745 (N_16745,N_5411,N_2125);
xnor U16746 (N_16746,N_5437,N_260);
and U16747 (N_16747,N_1689,N_3811);
and U16748 (N_16748,N_5881,N_2062);
nor U16749 (N_16749,N_1347,N_4581);
xnor U16750 (N_16750,N_8821,N_6605);
xor U16751 (N_16751,N_504,N_8325);
and U16752 (N_16752,N_389,N_6575);
or U16753 (N_16753,N_8048,N_5317);
nand U16754 (N_16754,N_2615,N_474);
nor U16755 (N_16755,N_3167,N_2882);
and U16756 (N_16756,N_7539,N_8221);
or U16757 (N_16757,N_4543,N_5356);
xor U16758 (N_16758,N_9562,N_9012);
xor U16759 (N_16759,N_315,N_1018);
or U16760 (N_16760,N_2863,N_4400);
xor U16761 (N_16761,N_6949,N_741);
and U16762 (N_16762,N_233,N_2908);
and U16763 (N_16763,N_652,N_82);
nand U16764 (N_16764,N_7013,N_4318);
or U16765 (N_16765,N_9218,N_6756);
and U16766 (N_16766,N_1236,N_8531);
nor U16767 (N_16767,N_8550,N_3606);
nand U16768 (N_16768,N_8038,N_8333);
or U16769 (N_16769,N_4713,N_3213);
nand U16770 (N_16770,N_2182,N_7623);
and U16771 (N_16771,N_4014,N_8890);
and U16772 (N_16772,N_5736,N_620);
and U16773 (N_16773,N_4136,N_5362);
xnor U16774 (N_16774,N_6593,N_5726);
and U16775 (N_16775,N_347,N_5875);
or U16776 (N_16776,N_3311,N_4287);
and U16777 (N_16777,N_6141,N_9110);
xor U16778 (N_16778,N_6675,N_938);
or U16779 (N_16779,N_6655,N_867);
or U16780 (N_16780,N_7846,N_4198);
or U16781 (N_16781,N_1643,N_4401);
or U16782 (N_16782,N_8422,N_2770);
nor U16783 (N_16783,N_7641,N_5063);
and U16784 (N_16784,N_2438,N_5377);
nand U16785 (N_16785,N_5028,N_3465);
nand U16786 (N_16786,N_4111,N_6076);
or U16787 (N_16787,N_7301,N_3112);
and U16788 (N_16788,N_7555,N_885);
or U16789 (N_16789,N_4234,N_6933);
nor U16790 (N_16790,N_8755,N_8070);
and U16791 (N_16791,N_6691,N_342);
nand U16792 (N_16792,N_7620,N_5208);
nor U16793 (N_16793,N_6415,N_3302);
nand U16794 (N_16794,N_3647,N_1236);
nor U16795 (N_16795,N_4791,N_3040);
nand U16796 (N_16796,N_1118,N_4099);
nor U16797 (N_16797,N_1310,N_946);
nor U16798 (N_16798,N_3410,N_491);
and U16799 (N_16799,N_5001,N_6184);
and U16800 (N_16800,N_4269,N_7102);
nor U16801 (N_16801,N_5369,N_6418);
nand U16802 (N_16802,N_1648,N_7984);
or U16803 (N_16803,N_3478,N_9174);
and U16804 (N_16804,N_8498,N_2915);
xor U16805 (N_16805,N_5518,N_460);
or U16806 (N_16806,N_810,N_596);
xnor U16807 (N_16807,N_6202,N_5146);
or U16808 (N_16808,N_2298,N_7019);
nor U16809 (N_16809,N_2977,N_5426);
nand U16810 (N_16810,N_8803,N_4276);
or U16811 (N_16811,N_4664,N_7127);
and U16812 (N_16812,N_8479,N_2250);
nand U16813 (N_16813,N_2254,N_8370);
and U16814 (N_16814,N_4454,N_3875);
and U16815 (N_16815,N_8355,N_9744);
nor U16816 (N_16816,N_7113,N_7415);
nor U16817 (N_16817,N_1852,N_8059);
and U16818 (N_16818,N_9531,N_2831);
nand U16819 (N_16819,N_6339,N_5726);
or U16820 (N_16820,N_4241,N_5020);
nand U16821 (N_16821,N_5375,N_1376);
xnor U16822 (N_16822,N_3839,N_8650);
or U16823 (N_16823,N_974,N_2682);
or U16824 (N_16824,N_4490,N_8898);
nor U16825 (N_16825,N_7293,N_2208);
or U16826 (N_16826,N_2020,N_5076);
xor U16827 (N_16827,N_4968,N_6780);
and U16828 (N_16828,N_3076,N_3456);
nand U16829 (N_16829,N_5194,N_2693);
nor U16830 (N_16830,N_1720,N_8159);
xnor U16831 (N_16831,N_4423,N_2622);
and U16832 (N_16832,N_5219,N_8731);
and U16833 (N_16833,N_3947,N_5728);
or U16834 (N_16834,N_1947,N_8036);
or U16835 (N_16835,N_1075,N_4102);
or U16836 (N_16836,N_7392,N_2368);
nor U16837 (N_16837,N_5643,N_6850);
and U16838 (N_16838,N_6228,N_3010);
nand U16839 (N_16839,N_7227,N_6100);
nand U16840 (N_16840,N_1830,N_8417);
nand U16841 (N_16841,N_8060,N_7228);
nor U16842 (N_16842,N_6609,N_4915);
xor U16843 (N_16843,N_7056,N_2057);
or U16844 (N_16844,N_1610,N_7534);
nand U16845 (N_16845,N_9566,N_4048);
and U16846 (N_16846,N_3270,N_5562);
xor U16847 (N_16847,N_1185,N_8373);
nor U16848 (N_16848,N_8468,N_1565);
nand U16849 (N_16849,N_3456,N_8041);
and U16850 (N_16850,N_5011,N_4906);
nand U16851 (N_16851,N_3275,N_7374);
and U16852 (N_16852,N_7172,N_516);
and U16853 (N_16853,N_9852,N_7216);
xnor U16854 (N_16854,N_1473,N_6863);
xnor U16855 (N_16855,N_7865,N_7434);
and U16856 (N_16856,N_2982,N_3835);
nand U16857 (N_16857,N_1907,N_5239);
nand U16858 (N_16858,N_8943,N_1719);
xor U16859 (N_16859,N_1382,N_2163);
or U16860 (N_16860,N_6695,N_5288);
and U16861 (N_16861,N_9703,N_1666);
xor U16862 (N_16862,N_2874,N_6470);
nand U16863 (N_16863,N_5910,N_1106);
nand U16864 (N_16864,N_3840,N_5027);
nand U16865 (N_16865,N_9553,N_5675);
or U16866 (N_16866,N_1861,N_7730);
nor U16867 (N_16867,N_9966,N_2192);
or U16868 (N_16868,N_1077,N_6376);
and U16869 (N_16869,N_2380,N_4288);
and U16870 (N_16870,N_8984,N_9055);
nor U16871 (N_16871,N_2083,N_6525);
xor U16872 (N_16872,N_8477,N_3643);
or U16873 (N_16873,N_8886,N_7138);
or U16874 (N_16874,N_1191,N_4403);
or U16875 (N_16875,N_270,N_189);
and U16876 (N_16876,N_6815,N_3391);
xnor U16877 (N_16877,N_9930,N_2898);
and U16878 (N_16878,N_4931,N_3898);
nor U16879 (N_16879,N_1078,N_9165);
nand U16880 (N_16880,N_3768,N_4029);
nand U16881 (N_16881,N_6284,N_6877);
or U16882 (N_16882,N_5932,N_1765);
and U16883 (N_16883,N_5374,N_2204);
nand U16884 (N_16884,N_8910,N_8596);
or U16885 (N_16885,N_7947,N_2054);
nand U16886 (N_16886,N_107,N_8247);
or U16887 (N_16887,N_2957,N_7132);
or U16888 (N_16888,N_6093,N_8098);
and U16889 (N_16889,N_440,N_3420);
nor U16890 (N_16890,N_4687,N_3903);
and U16891 (N_16891,N_9826,N_5823);
xor U16892 (N_16892,N_6298,N_3263);
or U16893 (N_16893,N_7727,N_8922);
nand U16894 (N_16894,N_3526,N_1049);
nand U16895 (N_16895,N_4622,N_6734);
or U16896 (N_16896,N_228,N_1704);
nor U16897 (N_16897,N_1948,N_1611);
and U16898 (N_16898,N_8627,N_6200);
nand U16899 (N_16899,N_1204,N_1602);
nand U16900 (N_16900,N_3100,N_6769);
and U16901 (N_16901,N_5057,N_5406);
or U16902 (N_16902,N_3109,N_9595);
nor U16903 (N_16903,N_5727,N_6875);
or U16904 (N_16904,N_3425,N_4933);
or U16905 (N_16905,N_2888,N_6408);
or U16906 (N_16906,N_5171,N_6254);
nor U16907 (N_16907,N_7168,N_7943);
nor U16908 (N_16908,N_453,N_6818);
nand U16909 (N_16909,N_8048,N_9519);
and U16910 (N_16910,N_1721,N_7466);
and U16911 (N_16911,N_6686,N_6981);
and U16912 (N_16912,N_1228,N_4685);
or U16913 (N_16913,N_3893,N_43);
and U16914 (N_16914,N_6111,N_854);
xnor U16915 (N_16915,N_4071,N_8609);
and U16916 (N_16916,N_5855,N_7727);
or U16917 (N_16917,N_5158,N_8307);
and U16918 (N_16918,N_9944,N_4914);
nand U16919 (N_16919,N_725,N_9374);
and U16920 (N_16920,N_3440,N_4517);
nor U16921 (N_16921,N_9722,N_324);
and U16922 (N_16922,N_5724,N_2678);
and U16923 (N_16923,N_4267,N_4032);
and U16924 (N_16924,N_5951,N_2547);
or U16925 (N_16925,N_7513,N_5510);
or U16926 (N_16926,N_8171,N_7925);
nor U16927 (N_16927,N_9368,N_7924);
or U16928 (N_16928,N_909,N_5077);
or U16929 (N_16929,N_5560,N_5114);
nor U16930 (N_16930,N_2277,N_1036);
nor U16931 (N_16931,N_9117,N_4792);
xor U16932 (N_16932,N_325,N_265);
nand U16933 (N_16933,N_2730,N_6814);
nor U16934 (N_16934,N_700,N_6894);
nand U16935 (N_16935,N_5924,N_661);
nor U16936 (N_16936,N_8932,N_1924);
and U16937 (N_16937,N_3402,N_4034);
and U16938 (N_16938,N_1427,N_4885);
and U16939 (N_16939,N_8764,N_832);
nor U16940 (N_16940,N_2811,N_9);
or U16941 (N_16941,N_8952,N_7336);
and U16942 (N_16942,N_8466,N_5674);
or U16943 (N_16943,N_5582,N_6322);
nor U16944 (N_16944,N_4637,N_181);
nor U16945 (N_16945,N_728,N_4015);
xnor U16946 (N_16946,N_758,N_1812);
nor U16947 (N_16947,N_1950,N_9425);
and U16948 (N_16948,N_6787,N_772);
nor U16949 (N_16949,N_6353,N_2144);
or U16950 (N_16950,N_8593,N_8458);
or U16951 (N_16951,N_8828,N_4660);
or U16952 (N_16952,N_516,N_9923);
and U16953 (N_16953,N_4099,N_7406);
or U16954 (N_16954,N_7133,N_1147);
nor U16955 (N_16955,N_192,N_3849);
nand U16956 (N_16956,N_960,N_7896);
nor U16957 (N_16957,N_9005,N_9762);
and U16958 (N_16958,N_4461,N_4154);
and U16959 (N_16959,N_7095,N_9785);
and U16960 (N_16960,N_1749,N_2113);
or U16961 (N_16961,N_1817,N_6296);
nand U16962 (N_16962,N_9222,N_7678);
and U16963 (N_16963,N_8543,N_4020);
xor U16964 (N_16964,N_6554,N_4649);
nand U16965 (N_16965,N_663,N_8920);
or U16966 (N_16966,N_476,N_2264);
or U16967 (N_16967,N_8298,N_8882);
nor U16968 (N_16968,N_6760,N_7927);
and U16969 (N_16969,N_2723,N_4917);
xnor U16970 (N_16970,N_7879,N_6814);
or U16971 (N_16971,N_2093,N_7220);
nand U16972 (N_16972,N_8465,N_1060);
or U16973 (N_16973,N_6508,N_3267);
or U16974 (N_16974,N_5113,N_6081);
and U16975 (N_16975,N_3573,N_482);
or U16976 (N_16976,N_3848,N_9658);
nand U16977 (N_16977,N_6784,N_1901);
or U16978 (N_16978,N_5457,N_1618);
nor U16979 (N_16979,N_5040,N_7956);
nor U16980 (N_16980,N_5020,N_4262);
nor U16981 (N_16981,N_738,N_8484);
and U16982 (N_16982,N_4418,N_89);
nand U16983 (N_16983,N_907,N_645);
nor U16984 (N_16984,N_9854,N_5248);
and U16985 (N_16985,N_4899,N_1786);
nor U16986 (N_16986,N_2082,N_4545);
or U16987 (N_16987,N_1420,N_8987);
and U16988 (N_16988,N_5776,N_3284);
xnor U16989 (N_16989,N_7870,N_8151);
or U16990 (N_16990,N_8958,N_4169);
nand U16991 (N_16991,N_9688,N_8276);
nand U16992 (N_16992,N_2666,N_5960);
and U16993 (N_16993,N_6732,N_9103);
or U16994 (N_16994,N_4712,N_9805);
nand U16995 (N_16995,N_1678,N_1466);
or U16996 (N_16996,N_8714,N_7681);
and U16997 (N_16997,N_7732,N_3445);
and U16998 (N_16998,N_2634,N_8318);
nor U16999 (N_16999,N_7243,N_8672);
and U17000 (N_17000,N_9407,N_2699);
nor U17001 (N_17001,N_1746,N_3678);
nand U17002 (N_17002,N_6376,N_2058);
or U17003 (N_17003,N_9072,N_988);
or U17004 (N_17004,N_8142,N_5898);
nor U17005 (N_17005,N_4908,N_9212);
and U17006 (N_17006,N_784,N_4188);
and U17007 (N_17007,N_4183,N_8999);
or U17008 (N_17008,N_8416,N_9548);
nor U17009 (N_17009,N_2655,N_4815);
xnor U17010 (N_17010,N_1842,N_8705);
and U17011 (N_17011,N_1972,N_7201);
or U17012 (N_17012,N_8612,N_9375);
or U17013 (N_17013,N_2030,N_6019);
and U17014 (N_17014,N_4145,N_6006);
nor U17015 (N_17015,N_4386,N_6069);
and U17016 (N_17016,N_787,N_7742);
nand U17017 (N_17017,N_3506,N_9039);
or U17018 (N_17018,N_5436,N_5746);
and U17019 (N_17019,N_5818,N_1455);
nand U17020 (N_17020,N_8645,N_413);
nand U17021 (N_17021,N_2181,N_6946);
or U17022 (N_17022,N_3024,N_9364);
xnor U17023 (N_17023,N_5111,N_4974);
nand U17024 (N_17024,N_8415,N_9629);
and U17025 (N_17025,N_219,N_1257);
or U17026 (N_17026,N_7600,N_729);
and U17027 (N_17027,N_1706,N_637);
nand U17028 (N_17028,N_5247,N_6178);
nand U17029 (N_17029,N_8742,N_96);
nor U17030 (N_17030,N_740,N_8691);
and U17031 (N_17031,N_3873,N_5102);
or U17032 (N_17032,N_136,N_9768);
xnor U17033 (N_17033,N_4669,N_8900);
nand U17034 (N_17034,N_199,N_8617);
nor U17035 (N_17035,N_9917,N_7062);
and U17036 (N_17036,N_688,N_9266);
and U17037 (N_17037,N_9298,N_2903);
nand U17038 (N_17038,N_6777,N_6117);
or U17039 (N_17039,N_5313,N_8534);
nand U17040 (N_17040,N_886,N_4828);
and U17041 (N_17041,N_9984,N_2306);
nand U17042 (N_17042,N_2731,N_6140);
or U17043 (N_17043,N_2040,N_2054);
and U17044 (N_17044,N_8301,N_7835);
nand U17045 (N_17045,N_1634,N_8194);
nor U17046 (N_17046,N_6984,N_8338);
nand U17047 (N_17047,N_5465,N_1624);
and U17048 (N_17048,N_8674,N_1273);
and U17049 (N_17049,N_44,N_959);
or U17050 (N_17050,N_9403,N_8101);
or U17051 (N_17051,N_4111,N_5662);
nand U17052 (N_17052,N_5544,N_4438);
nor U17053 (N_17053,N_3730,N_6747);
nand U17054 (N_17054,N_3017,N_2632);
nand U17055 (N_17055,N_1697,N_283);
xor U17056 (N_17056,N_9182,N_2394);
nand U17057 (N_17057,N_8210,N_3171);
nand U17058 (N_17058,N_2516,N_5607);
nand U17059 (N_17059,N_2287,N_9507);
nor U17060 (N_17060,N_6716,N_9927);
nor U17061 (N_17061,N_3521,N_2739);
nor U17062 (N_17062,N_3817,N_4655);
and U17063 (N_17063,N_144,N_4281);
nand U17064 (N_17064,N_4516,N_4610);
and U17065 (N_17065,N_9324,N_9645);
nor U17066 (N_17066,N_5813,N_8204);
nor U17067 (N_17067,N_5128,N_9869);
nor U17068 (N_17068,N_9688,N_2203);
or U17069 (N_17069,N_1673,N_310);
nand U17070 (N_17070,N_3485,N_7700);
xnor U17071 (N_17071,N_9677,N_524);
nor U17072 (N_17072,N_3353,N_6085);
or U17073 (N_17073,N_6686,N_4393);
nor U17074 (N_17074,N_140,N_2763);
and U17075 (N_17075,N_1837,N_3014);
nand U17076 (N_17076,N_147,N_8244);
or U17077 (N_17077,N_4855,N_9236);
and U17078 (N_17078,N_8979,N_2685);
nor U17079 (N_17079,N_382,N_825);
or U17080 (N_17080,N_5841,N_203);
xor U17081 (N_17081,N_5934,N_4387);
and U17082 (N_17082,N_9088,N_1408);
nor U17083 (N_17083,N_1840,N_8902);
nand U17084 (N_17084,N_6698,N_5850);
nor U17085 (N_17085,N_8184,N_2698);
and U17086 (N_17086,N_7180,N_8034);
and U17087 (N_17087,N_6256,N_3442);
nor U17088 (N_17088,N_6222,N_319);
and U17089 (N_17089,N_1308,N_1793);
and U17090 (N_17090,N_3370,N_8849);
nor U17091 (N_17091,N_6165,N_3632);
nand U17092 (N_17092,N_3390,N_5978);
and U17093 (N_17093,N_5614,N_9919);
nor U17094 (N_17094,N_1037,N_6069);
nand U17095 (N_17095,N_4276,N_3180);
nor U17096 (N_17096,N_3120,N_7597);
or U17097 (N_17097,N_2500,N_9153);
or U17098 (N_17098,N_9578,N_5640);
xnor U17099 (N_17099,N_3355,N_4002);
or U17100 (N_17100,N_1690,N_7773);
xor U17101 (N_17101,N_8317,N_5241);
nor U17102 (N_17102,N_8323,N_3295);
and U17103 (N_17103,N_1204,N_1100);
nor U17104 (N_17104,N_728,N_723);
and U17105 (N_17105,N_8079,N_2284);
xor U17106 (N_17106,N_9454,N_3696);
nor U17107 (N_17107,N_5967,N_9342);
or U17108 (N_17108,N_3842,N_6415);
nor U17109 (N_17109,N_8342,N_6125);
nand U17110 (N_17110,N_9891,N_1990);
nor U17111 (N_17111,N_4862,N_4333);
nor U17112 (N_17112,N_9300,N_7284);
nor U17113 (N_17113,N_4290,N_7159);
nand U17114 (N_17114,N_3915,N_389);
and U17115 (N_17115,N_3695,N_7029);
nor U17116 (N_17116,N_73,N_9733);
nand U17117 (N_17117,N_8211,N_5804);
or U17118 (N_17118,N_3999,N_1293);
nor U17119 (N_17119,N_6423,N_4508);
nand U17120 (N_17120,N_6240,N_5137);
nor U17121 (N_17121,N_2687,N_1673);
nand U17122 (N_17122,N_9054,N_4944);
nor U17123 (N_17123,N_8340,N_9863);
nor U17124 (N_17124,N_5411,N_7511);
or U17125 (N_17125,N_4489,N_7063);
nand U17126 (N_17126,N_7781,N_6506);
xor U17127 (N_17127,N_3620,N_7488);
xor U17128 (N_17128,N_2007,N_436);
or U17129 (N_17129,N_918,N_5638);
and U17130 (N_17130,N_1060,N_5423);
nor U17131 (N_17131,N_2464,N_9182);
nand U17132 (N_17132,N_1647,N_1902);
and U17133 (N_17133,N_1650,N_4636);
nand U17134 (N_17134,N_1276,N_7000);
or U17135 (N_17135,N_921,N_6839);
or U17136 (N_17136,N_8895,N_9125);
or U17137 (N_17137,N_27,N_3576);
and U17138 (N_17138,N_8874,N_8869);
nand U17139 (N_17139,N_336,N_6728);
nand U17140 (N_17140,N_7647,N_2563);
or U17141 (N_17141,N_7777,N_6249);
or U17142 (N_17142,N_7541,N_1618);
and U17143 (N_17143,N_5003,N_6893);
or U17144 (N_17144,N_8423,N_3993);
nor U17145 (N_17145,N_8235,N_8995);
xor U17146 (N_17146,N_7341,N_1285);
xnor U17147 (N_17147,N_9129,N_6073);
nand U17148 (N_17148,N_3943,N_7463);
nor U17149 (N_17149,N_5208,N_3398);
and U17150 (N_17150,N_5918,N_3183);
nor U17151 (N_17151,N_2468,N_1649);
nand U17152 (N_17152,N_2790,N_6081);
or U17153 (N_17153,N_3846,N_4659);
nand U17154 (N_17154,N_2532,N_3348);
or U17155 (N_17155,N_4217,N_9573);
nor U17156 (N_17156,N_6145,N_7062);
nor U17157 (N_17157,N_6820,N_2246);
nand U17158 (N_17158,N_7612,N_5275);
nand U17159 (N_17159,N_9697,N_465);
xnor U17160 (N_17160,N_5913,N_6045);
nor U17161 (N_17161,N_1367,N_5733);
and U17162 (N_17162,N_6614,N_4779);
nor U17163 (N_17163,N_3514,N_2894);
xnor U17164 (N_17164,N_8193,N_2406);
nand U17165 (N_17165,N_6092,N_2141);
and U17166 (N_17166,N_8384,N_8967);
and U17167 (N_17167,N_1262,N_838);
nor U17168 (N_17168,N_6985,N_1366);
and U17169 (N_17169,N_8399,N_4715);
nand U17170 (N_17170,N_8282,N_9137);
and U17171 (N_17171,N_5010,N_3623);
nor U17172 (N_17172,N_2542,N_8738);
and U17173 (N_17173,N_2188,N_3404);
or U17174 (N_17174,N_9295,N_524);
nor U17175 (N_17175,N_1011,N_3720);
nor U17176 (N_17176,N_9192,N_9417);
nand U17177 (N_17177,N_1150,N_4687);
nor U17178 (N_17178,N_5728,N_1259);
nand U17179 (N_17179,N_7344,N_6822);
nand U17180 (N_17180,N_7025,N_3152);
and U17181 (N_17181,N_6190,N_3283);
nor U17182 (N_17182,N_9571,N_9515);
nand U17183 (N_17183,N_3652,N_5801);
nand U17184 (N_17184,N_2976,N_7381);
or U17185 (N_17185,N_8179,N_1962);
or U17186 (N_17186,N_1301,N_3522);
xor U17187 (N_17187,N_5853,N_6176);
or U17188 (N_17188,N_3431,N_636);
nor U17189 (N_17189,N_7477,N_8721);
and U17190 (N_17190,N_8611,N_5175);
xor U17191 (N_17191,N_2069,N_7673);
nand U17192 (N_17192,N_9381,N_9960);
nor U17193 (N_17193,N_9293,N_855);
nand U17194 (N_17194,N_2830,N_112);
or U17195 (N_17195,N_970,N_6451);
or U17196 (N_17196,N_7890,N_4055);
nand U17197 (N_17197,N_8191,N_2651);
or U17198 (N_17198,N_118,N_6668);
nand U17199 (N_17199,N_4034,N_6012);
or U17200 (N_17200,N_7067,N_2870);
nand U17201 (N_17201,N_2105,N_8399);
or U17202 (N_17202,N_2078,N_8568);
and U17203 (N_17203,N_7673,N_3231);
xnor U17204 (N_17204,N_6107,N_8498);
nand U17205 (N_17205,N_9617,N_8425);
nand U17206 (N_17206,N_3158,N_1545);
and U17207 (N_17207,N_8950,N_4764);
xnor U17208 (N_17208,N_7656,N_1872);
nor U17209 (N_17209,N_391,N_9492);
and U17210 (N_17210,N_179,N_5246);
and U17211 (N_17211,N_4137,N_9442);
or U17212 (N_17212,N_7492,N_5478);
or U17213 (N_17213,N_2979,N_4874);
nor U17214 (N_17214,N_8851,N_7617);
nor U17215 (N_17215,N_5270,N_5817);
nor U17216 (N_17216,N_147,N_2459);
and U17217 (N_17217,N_4921,N_8170);
and U17218 (N_17218,N_8452,N_8367);
xor U17219 (N_17219,N_3146,N_6874);
xor U17220 (N_17220,N_6610,N_8697);
nor U17221 (N_17221,N_4730,N_6381);
or U17222 (N_17222,N_2521,N_5377);
and U17223 (N_17223,N_8988,N_7254);
or U17224 (N_17224,N_1630,N_2743);
or U17225 (N_17225,N_7129,N_1310);
nand U17226 (N_17226,N_4058,N_8231);
nand U17227 (N_17227,N_9965,N_3241);
and U17228 (N_17228,N_4570,N_9740);
xnor U17229 (N_17229,N_533,N_3303);
nand U17230 (N_17230,N_1850,N_4209);
xnor U17231 (N_17231,N_6335,N_4974);
and U17232 (N_17232,N_5477,N_6793);
and U17233 (N_17233,N_5733,N_2806);
and U17234 (N_17234,N_1048,N_6641);
nand U17235 (N_17235,N_9854,N_6505);
nand U17236 (N_17236,N_6035,N_1442);
and U17237 (N_17237,N_8707,N_4013);
xor U17238 (N_17238,N_8503,N_9687);
and U17239 (N_17239,N_7591,N_1108);
and U17240 (N_17240,N_9686,N_222);
and U17241 (N_17241,N_3218,N_5042);
and U17242 (N_17242,N_4743,N_698);
nor U17243 (N_17243,N_9071,N_6665);
and U17244 (N_17244,N_4974,N_7784);
or U17245 (N_17245,N_7359,N_8206);
nor U17246 (N_17246,N_8074,N_1050);
nand U17247 (N_17247,N_4307,N_7476);
and U17248 (N_17248,N_9532,N_9741);
and U17249 (N_17249,N_6133,N_849);
or U17250 (N_17250,N_7340,N_2463);
and U17251 (N_17251,N_876,N_1067);
nor U17252 (N_17252,N_496,N_1753);
or U17253 (N_17253,N_1580,N_6820);
nand U17254 (N_17254,N_2220,N_42);
and U17255 (N_17255,N_1086,N_2292);
nor U17256 (N_17256,N_9186,N_247);
or U17257 (N_17257,N_1494,N_7190);
nand U17258 (N_17258,N_1363,N_9562);
xnor U17259 (N_17259,N_7742,N_8714);
and U17260 (N_17260,N_2658,N_9597);
or U17261 (N_17261,N_988,N_9752);
nand U17262 (N_17262,N_7497,N_626);
nor U17263 (N_17263,N_5676,N_613);
xnor U17264 (N_17264,N_6376,N_5863);
and U17265 (N_17265,N_3652,N_1561);
and U17266 (N_17266,N_687,N_1903);
or U17267 (N_17267,N_6588,N_814);
nand U17268 (N_17268,N_1647,N_2132);
nand U17269 (N_17269,N_1354,N_5373);
nor U17270 (N_17270,N_5607,N_9858);
nor U17271 (N_17271,N_6362,N_301);
nand U17272 (N_17272,N_7107,N_5262);
or U17273 (N_17273,N_1465,N_3348);
nand U17274 (N_17274,N_8454,N_36);
or U17275 (N_17275,N_1293,N_4379);
and U17276 (N_17276,N_1578,N_3219);
or U17277 (N_17277,N_3629,N_9661);
nand U17278 (N_17278,N_7722,N_2008);
nand U17279 (N_17279,N_6828,N_4593);
nand U17280 (N_17280,N_8407,N_4961);
nand U17281 (N_17281,N_1747,N_6472);
and U17282 (N_17282,N_5939,N_4001);
and U17283 (N_17283,N_120,N_777);
and U17284 (N_17284,N_6158,N_82);
nor U17285 (N_17285,N_4185,N_5086);
or U17286 (N_17286,N_1250,N_8056);
nor U17287 (N_17287,N_3380,N_7462);
and U17288 (N_17288,N_2870,N_4374);
xnor U17289 (N_17289,N_3969,N_4197);
nand U17290 (N_17290,N_3460,N_6828);
nand U17291 (N_17291,N_6723,N_8596);
nand U17292 (N_17292,N_9704,N_9205);
nor U17293 (N_17293,N_2232,N_3814);
nand U17294 (N_17294,N_9318,N_5335);
and U17295 (N_17295,N_4048,N_5582);
or U17296 (N_17296,N_5814,N_8551);
or U17297 (N_17297,N_6850,N_2513);
nor U17298 (N_17298,N_5586,N_4274);
nand U17299 (N_17299,N_9562,N_8863);
or U17300 (N_17300,N_8628,N_9244);
and U17301 (N_17301,N_309,N_9720);
and U17302 (N_17302,N_2670,N_718);
or U17303 (N_17303,N_5749,N_7470);
xnor U17304 (N_17304,N_731,N_9979);
xnor U17305 (N_17305,N_5011,N_8420);
or U17306 (N_17306,N_7437,N_1760);
nor U17307 (N_17307,N_9196,N_2923);
nand U17308 (N_17308,N_5815,N_2690);
nand U17309 (N_17309,N_4881,N_6530);
and U17310 (N_17310,N_3120,N_4659);
or U17311 (N_17311,N_7701,N_6665);
xnor U17312 (N_17312,N_2755,N_3753);
and U17313 (N_17313,N_5872,N_4896);
nand U17314 (N_17314,N_158,N_8439);
and U17315 (N_17315,N_7454,N_9530);
nor U17316 (N_17316,N_8739,N_4197);
nor U17317 (N_17317,N_3174,N_1810);
or U17318 (N_17318,N_3387,N_7967);
and U17319 (N_17319,N_7223,N_7192);
nor U17320 (N_17320,N_369,N_7615);
nand U17321 (N_17321,N_7102,N_9325);
or U17322 (N_17322,N_6207,N_3233);
or U17323 (N_17323,N_5352,N_296);
and U17324 (N_17324,N_9171,N_6894);
nor U17325 (N_17325,N_159,N_6082);
or U17326 (N_17326,N_8612,N_8965);
nand U17327 (N_17327,N_9717,N_237);
or U17328 (N_17328,N_9896,N_7154);
xor U17329 (N_17329,N_1479,N_1687);
nor U17330 (N_17330,N_9445,N_7380);
or U17331 (N_17331,N_687,N_6400);
nor U17332 (N_17332,N_2983,N_5343);
nor U17333 (N_17333,N_7587,N_1301);
and U17334 (N_17334,N_5564,N_719);
or U17335 (N_17335,N_9148,N_5874);
nor U17336 (N_17336,N_4733,N_6080);
or U17337 (N_17337,N_6612,N_2725);
nor U17338 (N_17338,N_7773,N_8112);
nor U17339 (N_17339,N_7007,N_1967);
nor U17340 (N_17340,N_407,N_9198);
nand U17341 (N_17341,N_72,N_1789);
nor U17342 (N_17342,N_9532,N_1271);
or U17343 (N_17343,N_2880,N_636);
and U17344 (N_17344,N_8287,N_4937);
nand U17345 (N_17345,N_9397,N_651);
and U17346 (N_17346,N_8662,N_3206);
nor U17347 (N_17347,N_8354,N_1112);
nor U17348 (N_17348,N_3902,N_1751);
and U17349 (N_17349,N_2289,N_4888);
and U17350 (N_17350,N_9443,N_4742);
and U17351 (N_17351,N_7413,N_9245);
or U17352 (N_17352,N_6955,N_6437);
nor U17353 (N_17353,N_9123,N_9549);
nor U17354 (N_17354,N_8425,N_6405);
nand U17355 (N_17355,N_2424,N_6506);
nand U17356 (N_17356,N_3458,N_2620);
nand U17357 (N_17357,N_7620,N_8648);
nand U17358 (N_17358,N_9990,N_3687);
nor U17359 (N_17359,N_6378,N_6320);
or U17360 (N_17360,N_1747,N_4883);
or U17361 (N_17361,N_5319,N_5571);
and U17362 (N_17362,N_9306,N_752);
nand U17363 (N_17363,N_3926,N_3043);
or U17364 (N_17364,N_5730,N_4451);
nand U17365 (N_17365,N_8132,N_4010);
nor U17366 (N_17366,N_5866,N_751);
or U17367 (N_17367,N_2184,N_1666);
and U17368 (N_17368,N_4197,N_3386);
and U17369 (N_17369,N_550,N_7537);
nor U17370 (N_17370,N_4224,N_873);
nor U17371 (N_17371,N_3763,N_4638);
or U17372 (N_17372,N_3768,N_1178);
nand U17373 (N_17373,N_3435,N_4661);
nand U17374 (N_17374,N_2607,N_5337);
nor U17375 (N_17375,N_8175,N_5089);
xnor U17376 (N_17376,N_2905,N_108);
nand U17377 (N_17377,N_7781,N_4791);
or U17378 (N_17378,N_8506,N_8830);
nor U17379 (N_17379,N_1819,N_6829);
or U17380 (N_17380,N_4445,N_5078);
and U17381 (N_17381,N_1783,N_9471);
xor U17382 (N_17382,N_1676,N_3686);
and U17383 (N_17383,N_6434,N_1541);
and U17384 (N_17384,N_5942,N_5623);
nand U17385 (N_17385,N_4911,N_9589);
nand U17386 (N_17386,N_9417,N_2693);
or U17387 (N_17387,N_9389,N_1157);
or U17388 (N_17388,N_603,N_7849);
xnor U17389 (N_17389,N_2788,N_5481);
and U17390 (N_17390,N_9824,N_2558);
and U17391 (N_17391,N_9712,N_3459);
nand U17392 (N_17392,N_8883,N_2973);
nor U17393 (N_17393,N_9968,N_5265);
or U17394 (N_17394,N_3505,N_9499);
nor U17395 (N_17395,N_3955,N_1390);
and U17396 (N_17396,N_2819,N_7596);
nand U17397 (N_17397,N_6668,N_2056);
xor U17398 (N_17398,N_5478,N_6977);
nor U17399 (N_17399,N_8550,N_2446);
and U17400 (N_17400,N_1866,N_6114);
nand U17401 (N_17401,N_8445,N_9157);
or U17402 (N_17402,N_8205,N_7392);
or U17403 (N_17403,N_6688,N_1829);
and U17404 (N_17404,N_7613,N_5711);
nor U17405 (N_17405,N_7055,N_3626);
nand U17406 (N_17406,N_4612,N_8765);
or U17407 (N_17407,N_699,N_1685);
nand U17408 (N_17408,N_6514,N_9696);
and U17409 (N_17409,N_9930,N_7598);
nand U17410 (N_17410,N_7857,N_9172);
nor U17411 (N_17411,N_4415,N_8761);
or U17412 (N_17412,N_110,N_579);
nor U17413 (N_17413,N_7002,N_2237);
or U17414 (N_17414,N_5031,N_3544);
nand U17415 (N_17415,N_7458,N_7965);
or U17416 (N_17416,N_9373,N_3396);
nand U17417 (N_17417,N_1282,N_8538);
or U17418 (N_17418,N_5995,N_1290);
nor U17419 (N_17419,N_5409,N_4959);
or U17420 (N_17420,N_7166,N_3295);
nand U17421 (N_17421,N_3587,N_6325);
or U17422 (N_17422,N_1574,N_932);
nand U17423 (N_17423,N_2044,N_6396);
or U17424 (N_17424,N_8196,N_1611);
and U17425 (N_17425,N_3315,N_6991);
nor U17426 (N_17426,N_9831,N_19);
and U17427 (N_17427,N_5273,N_5297);
and U17428 (N_17428,N_6605,N_1003);
and U17429 (N_17429,N_8068,N_6547);
nand U17430 (N_17430,N_9698,N_6802);
nor U17431 (N_17431,N_6715,N_7829);
or U17432 (N_17432,N_4523,N_8452);
nand U17433 (N_17433,N_8005,N_3467);
or U17434 (N_17434,N_8180,N_4431);
nand U17435 (N_17435,N_2800,N_1516);
nor U17436 (N_17436,N_7303,N_2830);
nor U17437 (N_17437,N_3433,N_170);
and U17438 (N_17438,N_8338,N_8595);
nor U17439 (N_17439,N_1725,N_1784);
nand U17440 (N_17440,N_4350,N_3314);
nor U17441 (N_17441,N_6384,N_2840);
nor U17442 (N_17442,N_6935,N_1144);
and U17443 (N_17443,N_6277,N_1177);
or U17444 (N_17444,N_7513,N_1281);
and U17445 (N_17445,N_5462,N_7424);
nand U17446 (N_17446,N_9479,N_7467);
xor U17447 (N_17447,N_7214,N_3652);
nor U17448 (N_17448,N_1962,N_5319);
nor U17449 (N_17449,N_4511,N_2170);
xnor U17450 (N_17450,N_1716,N_8377);
xnor U17451 (N_17451,N_1898,N_3802);
or U17452 (N_17452,N_901,N_1814);
xnor U17453 (N_17453,N_9975,N_268);
nand U17454 (N_17454,N_9719,N_8745);
nor U17455 (N_17455,N_537,N_2062);
and U17456 (N_17456,N_112,N_2649);
and U17457 (N_17457,N_2033,N_602);
and U17458 (N_17458,N_9187,N_2375);
nor U17459 (N_17459,N_2250,N_9256);
nand U17460 (N_17460,N_1209,N_7691);
xor U17461 (N_17461,N_7769,N_1499);
nand U17462 (N_17462,N_6476,N_1376);
nand U17463 (N_17463,N_4488,N_2514);
or U17464 (N_17464,N_2467,N_5589);
or U17465 (N_17465,N_7872,N_7153);
nand U17466 (N_17466,N_3369,N_4357);
nand U17467 (N_17467,N_225,N_3845);
or U17468 (N_17468,N_8336,N_6085);
xor U17469 (N_17469,N_9115,N_8186);
or U17470 (N_17470,N_9530,N_7250);
or U17471 (N_17471,N_9510,N_923);
nand U17472 (N_17472,N_174,N_9411);
and U17473 (N_17473,N_684,N_6017);
nor U17474 (N_17474,N_234,N_5402);
nand U17475 (N_17475,N_9422,N_3014);
or U17476 (N_17476,N_5105,N_5451);
or U17477 (N_17477,N_427,N_6099);
or U17478 (N_17478,N_4020,N_4683);
or U17479 (N_17479,N_3493,N_8307);
and U17480 (N_17480,N_6490,N_5074);
nand U17481 (N_17481,N_4809,N_5029);
or U17482 (N_17482,N_7584,N_5260);
nor U17483 (N_17483,N_978,N_3191);
or U17484 (N_17484,N_4393,N_5428);
and U17485 (N_17485,N_3054,N_3360);
nor U17486 (N_17486,N_3726,N_6920);
nor U17487 (N_17487,N_3284,N_5406);
nor U17488 (N_17488,N_6668,N_7763);
nor U17489 (N_17489,N_4017,N_891);
and U17490 (N_17490,N_1818,N_5536);
xor U17491 (N_17491,N_2140,N_5462);
or U17492 (N_17492,N_5485,N_4113);
nor U17493 (N_17493,N_4227,N_2966);
nor U17494 (N_17494,N_3769,N_9155);
and U17495 (N_17495,N_4728,N_3560);
xnor U17496 (N_17496,N_1251,N_5493);
xor U17497 (N_17497,N_4625,N_4555);
and U17498 (N_17498,N_5546,N_2874);
nand U17499 (N_17499,N_8226,N_5372);
nor U17500 (N_17500,N_3875,N_127);
and U17501 (N_17501,N_9475,N_2012);
and U17502 (N_17502,N_2031,N_6802);
nor U17503 (N_17503,N_7511,N_6506);
nor U17504 (N_17504,N_6378,N_1388);
nand U17505 (N_17505,N_9387,N_859);
nand U17506 (N_17506,N_7254,N_3784);
or U17507 (N_17507,N_6035,N_4256);
nand U17508 (N_17508,N_9109,N_549);
or U17509 (N_17509,N_2212,N_1187);
or U17510 (N_17510,N_8136,N_4657);
and U17511 (N_17511,N_9285,N_613);
nor U17512 (N_17512,N_4921,N_3684);
or U17513 (N_17513,N_8070,N_4053);
or U17514 (N_17514,N_159,N_7449);
and U17515 (N_17515,N_4295,N_8241);
xor U17516 (N_17516,N_9525,N_1245);
nand U17517 (N_17517,N_4784,N_704);
xor U17518 (N_17518,N_1208,N_8286);
nand U17519 (N_17519,N_3129,N_866);
or U17520 (N_17520,N_701,N_6732);
nand U17521 (N_17521,N_7551,N_3433);
or U17522 (N_17522,N_861,N_1463);
nand U17523 (N_17523,N_3120,N_7922);
xor U17524 (N_17524,N_6822,N_3980);
nand U17525 (N_17525,N_8870,N_8021);
and U17526 (N_17526,N_5356,N_1175);
nor U17527 (N_17527,N_2218,N_9268);
nand U17528 (N_17528,N_9092,N_8894);
and U17529 (N_17529,N_4525,N_2341);
and U17530 (N_17530,N_5571,N_1095);
and U17531 (N_17531,N_149,N_8894);
nor U17532 (N_17532,N_4438,N_4199);
and U17533 (N_17533,N_4258,N_3018);
or U17534 (N_17534,N_1404,N_504);
nand U17535 (N_17535,N_360,N_9610);
or U17536 (N_17536,N_6733,N_383);
or U17537 (N_17537,N_2519,N_6697);
nand U17538 (N_17538,N_4317,N_2974);
and U17539 (N_17539,N_2325,N_1335);
or U17540 (N_17540,N_4882,N_499);
or U17541 (N_17541,N_2422,N_9682);
or U17542 (N_17542,N_2543,N_8414);
and U17543 (N_17543,N_549,N_2227);
or U17544 (N_17544,N_4625,N_514);
nand U17545 (N_17545,N_9465,N_8074);
nor U17546 (N_17546,N_9010,N_755);
nor U17547 (N_17547,N_3215,N_1004);
nor U17548 (N_17548,N_693,N_5121);
nand U17549 (N_17549,N_8184,N_5989);
and U17550 (N_17550,N_4136,N_104);
and U17551 (N_17551,N_372,N_9750);
nor U17552 (N_17552,N_1903,N_6483);
nor U17553 (N_17553,N_8550,N_7533);
nand U17554 (N_17554,N_306,N_5935);
nand U17555 (N_17555,N_1676,N_1277);
or U17556 (N_17556,N_1871,N_4872);
nand U17557 (N_17557,N_4146,N_5332);
and U17558 (N_17558,N_6809,N_8245);
nand U17559 (N_17559,N_6472,N_5705);
or U17560 (N_17560,N_8713,N_3764);
nor U17561 (N_17561,N_3328,N_3572);
nand U17562 (N_17562,N_3076,N_5797);
nand U17563 (N_17563,N_3397,N_3568);
or U17564 (N_17564,N_1943,N_6848);
nand U17565 (N_17565,N_5980,N_9359);
and U17566 (N_17566,N_7182,N_4424);
nor U17567 (N_17567,N_9599,N_6615);
nand U17568 (N_17568,N_6133,N_4120);
nor U17569 (N_17569,N_6647,N_5340);
and U17570 (N_17570,N_3942,N_7482);
xnor U17571 (N_17571,N_9042,N_2510);
or U17572 (N_17572,N_2795,N_772);
nand U17573 (N_17573,N_6040,N_1995);
nand U17574 (N_17574,N_2332,N_4605);
and U17575 (N_17575,N_6629,N_8382);
nor U17576 (N_17576,N_8266,N_8661);
nand U17577 (N_17577,N_3328,N_4648);
or U17578 (N_17578,N_6376,N_1919);
or U17579 (N_17579,N_9919,N_7286);
or U17580 (N_17580,N_2149,N_1492);
xor U17581 (N_17581,N_2321,N_8854);
or U17582 (N_17582,N_1131,N_7319);
or U17583 (N_17583,N_8773,N_719);
nand U17584 (N_17584,N_5448,N_5955);
nor U17585 (N_17585,N_1053,N_1361);
nor U17586 (N_17586,N_7508,N_1464);
xnor U17587 (N_17587,N_2642,N_6720);
and U17588 (N_17588,N_87,N_5407);
xor U17589 (N_17589,N_2722,N_5576);
nor U17590 (N_17590,N_5952,N_1149);
or U17591 (N_17591,N_3480,N_7483);
nor U17592 (N_17592,N_5368,N_9257);
or U17593 (N_17593,N_9815,N_331);
xnor U17594 (N_17594,N_9146,N_807);
nor U17595 (N_17595,N_7943,N_9503);
nand U17596 (N_17596,N_137,N_9634);
nand U17597 (N_17597,N_5120,N_7696);
and U17598 (N_17598,N_7095,N_8462);
or U17599 (N_17599,N_6274,N_6108);
nand U17600 (N_17600,N_8599,N_3608);
nand U17601 (N_17601,N_3278,N_6286);
or U17602 (N_17602,N_3481,N_1576);
nand U17603 (N_17603,N_3711,N_7216);
or U17604 (N_17604,N_1164,N_9455);
nor U17605 (N_17605,N_2688,N_4601);
and U17606 (N_17606,N_2313,N_7495);
nor U17607 (N_17607,N_2413,N_6662);
and U17608 (N_17608,N_657,N_457);
nor U17609 (N_17609,N_6827,N_4401);
and U17610 (N_17610,N_5472,N_4722);
and U17611 (N_17611,N_1252,N_4899);
or U17612 (N_17612,N_8149,N_8251);
nor U17613 (N_17613,N_2009,N_4457);
nand U17614 (N_17614,N_7017,N_6172);
or U17615 (N_17615,N_8436,N_2182);
nor U17616 (N_17616,N_2468,N_7879);
xor U17617 (N_17617,N_9126,N_7853);
and U17618 (N_17618,N_5503,N_8312);
nand U17619 (N_17619,N_6103,N_9159);
and U17620 (N_17620,N_1290,N_9319);
or U17621 (N_17621,N_5474,N_9546);
nand U17622 (N_17622,N_9752,N_4785);
or U17623 (N_17623,N_1092,N_4168);
xor U17624 (N_17624,N_1343,N_3569);
and U17625 (N_17625,N_6667,N_2458);
and U17626 (N_17626,N_5763,N_602);
and U17627 (N_17627,N_5125,N_5893);
nor U17628 (N_17628,N_4016,N_5461);
nor U17629 (N_17629,N_8429,N_7133);
and U17630 (N_17630,N_2462,N_4064);
xnor U17631 (N_17631,N_4432,N_6911);
nor U17632 (N_17632,N_7627,N_241);
and U17633 (N_17633,N_2007,N_667);
nor U17634 (N_17634,N_7144,N_9070);
and U17635 (N_17635,N_4881,N_3630);
and U17636 (N_17636,N_1097,N_9588);
nand U17637 (N_17637,N_4749,N_6547);
xnor U17638 (N_17638,N_1817,N_4353);
xnor U17639 (N_17639,N_3499,N_5400);
nor U17640 (N_17640,N_3741,N_3170);
or U17641 (N_17641,N_3074,N_5501);
nand U17642 (N_17642,N_654,N_9708);
or U17643 (N_17643,N_5393,N_8435);
xnor U17644 (N_17644,N_601,N_6547);
nor U17645 (N_17645,N_1984,N_2051);
or U17646 (N_17646,N_676,N_5226);
nand U17647 (N_17647,N_6748,N_6570);
nor U17648 (N_17648,N_2837,N_7782);
nor U17649 (N_17649,N_5580,N_144);
nor U17650 (N_17650,N_4118,N_1847);
nand U17651 (N_17651,N_9244,N_2117);
nand U17652 (N_17652,N_4010,N_6114);
and U17653 (N_17653,N_1203,N_9035);
and U17654 (N_17654,N_3799,N_3415);
nand U17655 (N_17655,N_4356,N_4956);
or U17656 (N_17656,N_7639,N_7591);
and U17657 (N_17657,N_6326,N_1357);
or U17658 (N_17658,N_26,N_1287);
nor U17659 (N_17659,N_5379,N_9598);
or U17660 (N_17660,N_2395,N_2853);
nor U17661 (N_17661,N_537,N_5754);
xor U17662 (N_17662,N_9400,N_1084);
nor U17663 (N_17663,N_8905,N_869);
nand U17664 (N_17664,N_5544,N_1619);
or U17665 (N_17665,N_9427,N_2699);
and U17666 (N_17666,N_5540,N_438);
or U17667 (N_17667,N_1983,N_4347);
xor U17668 (N_17668,N_5619,N_3068);
nand U17669 (N_17669,N_4388,N_1619);
nor U17670 (N_17670,N_5718,N_270);
nand U17671 (N_17671,N_3432,N_4787);
and U17672 (N_17672,N_2821,N_8161);
and U17673 (N_17673,N_3827,N_5327);
or U17674 (N_17674,N_1365,N_394);
and U17675 (N_17675,N_9079,N_6646);
nor U17676 (N_17676,N_9481,N_6252);
or U17677 (N_17677,N_3417,N_1461);
nand U17678 (N_17678,N_1659,N_9647);
nor U17679 (N_17679,N_3681,N_5734);
or U17680 (N_17680,N_1116,N_2225);
nand U17681 (N_17681,N_7430,N_7912);
or U17682 (N_17682,N_4295,N_8305);
or U17683 (N_17683,N_7193,N_5932);
or U17684 (N_17684,N_7243,N_2207);
xnor U17685 (N_17685,N_1842,N_6508);
nand U17686 (N_17686,N_2815,N_257);
nor U17687 (N_17687,N_672,N_7977);
and U17688 (N_17688,N_9438,N_3528);
nand U17689 (N_17689,N_6077,N_6764);
xor U17690 (N_17690,N_1020,N_7134);
nand U17691 (N_17691,N_80,N_5651);
or U17692 (N_17692,N_6097,N_9382);
or U17693 (N_17693,N_3456,N_9156);
and U17694 (N_17694,N_224,N_8332);
or U17695 (N_17695,N_4981,N_5007);
nor U17696 (N_17696,N_1459,N_9935);
nand U17697 (N_17697,N_2814,N_7698);
nand U17698 (N_17698,N_1580,N_395);
or U17699 (N_17699,N_1661,N_5180);
nor U17700 (N_17700,N_829,N_8647);
or U17701 (N_17701,N_4318,N_9940);
nor U17702 (N_17702,N_8157,N_8505);
xor U17703 (N_17703,N_6321,N_5947);
nand U17704 (N_17704,N_8918,N_2781);
and U17705 (N_17705,N_4320,N_3962);
or U17706 (N_17706,N_630,N_6417);
or U17707 (N_17707,N_9228,N_7600);
xnor U17708 (N_17708,N_5670,N_8458);
nand U17709 (N_17709,N_867,N_3569);
nor U17710 (N_17710,N_1986,N_2321);
nand U17711 (N_17711,N_6627,N_7792);
nor U17712 (N_17712,N_677,N_8042);
nor U17713 (N_17713,N_8088,N_7806);
or U17714 (N_17714,N_9465,N_6778);
or U17715 (N_17715,N_8102,N_52);
or U17716 (N_17716,N_8665,N_4709);
nand U17717 (N_17717,N_9096,N_5463);
nand U17718 (N_17718,N_9740,N_4874);
or U17719 (N_17719,N_7064,N_1681);
nand U17720 (N_17720,N_796,N_6509);
or U17721 (N_17721,N_1826,N_7886);
xor U17722 (N_17722,N_3077,N_9094);
and U17723 (N_17723,N_943,N_9299);
or U17724 (N_17724,N_7853,N_835);
xor U17725 (N_17725,N_5981,N_6498);
nor U17726 (N_17726,N_4220,N_5667);
nor U17727 (N_17727,N_6724,N_3032);
or U17728 (N_17728,N_6109,N_3602);
nor U17729 (N_17729,N_9711,N_6049);
and U17730 (N_17730,N_7597,N_8855);
or U17731 (N_17731,N_1054,N_8124);
or U17732 (N_17732,N_2724,N_2371);
or U17733 (N_17733,N_8741,N_820);
nand U17734 (N_17734,N_8036,N_4438);
nand U17735 (N_17735,N_3576,N_7038);
nand U17736 (N_17736,N_3625,N_9355);
nor U17737 (N_17737,N_776,N_5717);
xnor U17738 (N_17738,N_9799,N_7644);
xor U17739 (N_17739,N_3376,N_6159);
or U17740 (N_17740,N_5475,N_4312);
nor U17741 (N_17741,N_3838,N_9769);
and U17742 (N_17742,N_5262,N_3453);
nor U17743 (N_17743,N_4675,N_8739);
nor U17744 (N_17744,N_5291,N_8746);
and U17745 (N_17745,N_2488,N_4866);
nand U17746 (N_17746,N_1980,N_728);
or U17747 (N_17747,N_2613,N_9470);
or U17748 (N_17748,N_4912,N_205);
nand U17749 (N_17749,N_3010,N_2440);
nand U17750 (N_17750,N_2393,N_8391);
and U17751 (N_17751,N_3083,N_1609);
nand U17752 (N_17752,N_1470,N_7369);
xor U17753 (N_17753,N_1961,N_4823);
nand U17754 (N_17754,N_8864,N_8352);
or U17755 (N_17755,N_5536,N_2119);
nand U17756 (N_17756,N_3713,N_1418);
nor U17757 (N_17757,N_9916,N_6446);
nand U17758 (N_17758,N_3621,N_8068);
or U17759 (N_17759,N_6672,N_9134);
or U17760 (N_17760,N_6654,N_7478);
and U17761 (N_17761,N_4933,N_6019);
and U17762 (N_17762,N_3128,N_3156);
nor U17763 (N_17763,N_544,N_8253);
xnor U17764 (N_17764,N_3001,N_6639);
and U17765 (N_17765,N_3768,N_1803);
and U17766 (N_17766,N_4072,N_9132);
and U17767 (N_17767,N_4876,N_6515);
nand U17768 (N_17768,N_602,N_5473);
and U17769 (N_17769,N_1206,N_7484);
or U17770 (N_17770,N_9831,N_3839);
and U17771 (N_17771,N_6628,N_7099);
or U17772 (N_17772,N_6689,N_8434);
xor U17773 (N_17773,N_5622,N_1268);
nor U17774 (N_17774,N_5265,N_4435);
or U17775 (N_17775,N_8053,N_7605);
or U17776 (N_17776,N_6236,N_6099);
nand U17777 (N_17777,N_86,N_1340);
or U17778 (N_17778,N_139,N_6216);
and U17779 (N_17779,N_4876,N_1742);
nor U17780 (N_17780,N_3286,N_6866);
nor U17781 (N_17781,N_7605,N_6198);
nand U17782 (N_17782,N_5433,N_8833);
or U17783 (N_17783,N_3413,N_8602);
nand U17784 (N_17784,N_8698,N_3253);
nor U17785 (N_17785,N_2737,N_4110);
and U17786 (N_17786,N_6872,N_6945);
nand U17787 (N_17787,N_3730,N_5519);
nand U17788 (N_17788,N_5605,N_6013);
nor U17789 (N_17789,N_1355,N_3171);
or U17790 (N_17790,N_6640,N_9670);
nand U17791 (N_17791,N_5880,N_4816);
and U17792 (N_17792,N_407,N_4290);
nand U17793 (N_17793,N_647,N_8184);
nor U17794 (N_17794,N_9049,N_5260);
nand U17795 (N_17795,N_1509,N_463);
nor U17796 (N_17796,N_6939,N_130);
nand U17797 (N_17797,N_8449,N_8416);
and U17798 (N_17798,N_6430,N_9707);
nand U17799 (N_17799,N_4003,N_9884);
or U17800 (N_17800,N_5770,N_1845);
or U17801 (N_17801,N_4305,N_5101);
xnor U17802 (N_17802,N_473,N_4205);
and U17803 (N_17803,N_7343,N_1449);
and U17804 (N_17804,N_8148,N_6569);
nand U17805 (N_17805,N_3665,N_4352);
xnor U17806 (N_17806,N_8385,N_4101);
or U17807 (N_17807,N_4743,N_980);
nor U17808 (N_17808,N_6663,N_7323);
and U17809 (N_17809,N_5135,N_5712);
nor U17810 (N_17810,N_6191,N_2733);
nor U17811 (N_17811,N_8162,N_5504);
nor U17812 (N_17812,N_7979,N_6579);
and U17813 (N_17813,N_7721,N_9115);
nand U17814 (N_17814,N_7533,N_8555);
nand U17815 (N_17815,N_5390,N_8248);
or U17816 (N_17816,N_787,N_9881);
and U17817 (N_17817,N_4517,N_5050);
and U17818 (N_17818,N_6037,N_8985);
and U17819 (N_17819,N_651,N_3003);
nor U17820 (N_17820,N_3508,N_861);
and U17821 (N_17821,N_3707,N_6625);
nand U17822 (N_17822,N_7808,N_9959);
xor U17823 (N_17823,N_7963,N_7411);
xnor U17824 (N_17824,N_7582,N_3629);
nand U17825 (N_17825,N_6929,N_6980);
and U17826 (N_17826,N_284,N_1056);
and U17827 (N_17827,N_3658,N_7803);
nand U17828 (N_17828,N_1052,N_6992);
and U17829 (N_17829,N_5539,N_2200);
nor U17830 (N_17830,N_4960,N_1338);
or U17831 (N_17831,N_3986,N_7341);
and U17832 (N_17832,N_59,N_1797);
xnor U17833 (N_17833,N_3367,N_6520);
nor U17834 (N_17834,N_348,N_7281);
xnor U17835 (N_17835,N_6133,N_598);
or U17836 (N_17836,N_4555,N_5752);
xnor U17837 (N_17837,N_4683,N_8904);
or U17838 (N_17838,N_3400,N_8607);
or U17839 (N_17839,N_3332,N_1421);
and U17840 (N_17840,N_3567,N_1875);
or U17841 (N_17841,N_1862,N_1059);
and U17842 (N_17842,N_1009,N_9911);
nor U17843 (N_17843,N_5411,N_9304);
nand U17844 (N_17844,N_4915,N_5261);
or U17845 (N_17845,N_9289,N_3008);
and U17846 (N_17846,N_2381,N_2959);
nor U17847 (N_17847,N_2135,N_107);
xor U17848 (N_17848,N_9557,N_8536);
nor U17849 (N_17849,N_1189,N_643);
xnor U17850 (N_17850,N_1664,N_4754);
xor U17851 (N_17851,N_5570,N_4704);
or U17852 (N_17852,N_8618,N_5558);
nor U17853 (N_17853,N_3602,N_8192);
and U17854 (N_17854,N_1569,N_5778);
nand U17855 (N_17855,N_5863,N_4434);
or U17856 (N_17856,N_1888,N_3079);
and U17857 (N_17857,N_8422,N_4373);
nor U17858 (N_17858,N_7407,N_2263);
xnor U17859 (N_17859,N_4353,N_8801);
and U17860 (N_17860,N_2211,N_5588);
nor U17861 (N_17861,N_4790,N_6168);
xnor U17862 (N_17862,N_502,N_3821);
and U17863 (N_17863,N_7585,N_7987);
and U17864 (N_17864,N_885,N_6340);
or U17865 (N_17865,N_3071,N_9768);
or U17866 (N_17866,N_4681,N_5659);
and U17867 (N_17867,N_2795,N_1167);
nand U17868 (N_17868,N_9246,N_7161);
xor U17869 (N_17869,N_6687,N_1253);
or U17870 (N_17870,N_7035,N_1245);
and U17871 (N_17871,N_1397,N_8308);
nand U17872 (N_17872,N_5990,N_6103);
nor U17873 (N_17873,N_6795,N_6601);
and U17874 (N_17874,N_807,N_891);
xor U17875 (N_17875,N_2341,N_5940);
xor U17876 (N_17876,N_1213,N_156);
nor U17877 (N_17877,N_2508,N_5066);
and U17878 (N_17878,N_4067,N_1029);
nor U17879 (N_17879,N_3249,N_9632);
xor U17880 (N_17880,N_1199,N_7722);
nand U17881 (N_17881,N_3287,N_2804);
or U17882 (N_17882,N_5300,N_7455);
or U17883 (N_17883,N_812,N_744);
and U17884 (N_17884,N_3394,N_5572);
nor U17885 (N_17885,N_5389,N_2485);
xor U17886 (N_17886,N_8211,N_2295);
nor U17887 (N_17887,N_342,N_7436);
and U17888 (N_17888,N_9163,N_9977);
or U17889 (N_17889,N_4138,N_1894);
xnor U17890 (N_17890,N_2144,N_5447);
nor U17891 (N_17891,N_3475,N_5107);
xnor U17892 (N_17892,N_2903,N_8251);
nor U17893 (N_17893,N_317,N_9144);
and U17894 (N_17894,N_6712,N_5846);
or U17895 (N_17895,N_6443,N_9511);
and U17896 (N_17896,N_7120,N_3500);
xor U17897 (N_17897,N_4224,N_8053);
or U17898 (N_17898,N_5967,N_209);
and U17899 (N_17899,N_6597,N_2404);
nand U17900 (N_17900,N_3598,N_6936);
nand U17901 (N_17901,N_1704,N_8961);
and U17902 (N_17902,N_590,N_6129);
nand U17903 (N_17903,N_634,N_4391);
or U17904 (N_17904,N_9250,N_290);
nand U17905 (N_17905,N_3502,N_778);
and U17906 (N_17906,N_2361,N_4860);
nand U17907 (N_17907,N_707,N_5085);
nor U17908 (N_17908,N_3127,N_177);
and U17909 (N_17909,N_2330,N_8117);
nand U17910 (N_17910,N_2772,N_3504);
nand U17911 (N_17911,N_3216,N_3548);
or U17912 (N_17912,N_2678,N_2528);
nor U17913 (N_17913,N_6057,N_5587);
or U17914 (N_17914,N_3923,N_6447);
nor U17915 (N_17915,N_5158,N_5975);
or U17916 (N_17916,N_3080,N_3295);
and U17917 (N_17917,N_3508,N_4405);
or U17918 (N_17918,N_7048,N_1501);
nand U17919 (N_17919,N_5738,N_3266);
nor U17920 (N_17920,N_3914,N_4533);
or U17921 (N_17921,N_6094,N_879);
and U17922 (N_17922,N_8896,N_1610);
and U17923 (N_17923,N_2484,N_7637);
and U17924 (N_17924,N_7020,N_8306);
and U17925 (N_17925,N_6088,N_2119);
nand U17926 (N_17926,N_7597,N_8893);
or U17927 (N_17927,N_300,N_137);
nand U17928 (N_17928,N_6429,N_1707);
or U17929 (N_17929,N_8654,N_3729);
and U17930 (N_17930,N_6688,N_8399);
nor U17931 (N_17931,N_4254,N_2020);
and U17932 (N_17932,N_7495,N_7435);
nor U17933 (N_17933,N_593,N_6188);
or U17934 (N_17934,N_416,N_7286);
nor U17935 (N_17935,N_4042,N_1479);
nand U17936 (N_17936,N_146,N_1921);
and U17937 (N_17937,N_9932,N_3042);
and U17938 (N_17938,N_5229,N_2701);
nor U17939 (N_17939,N_1981,N_9771);
nor U17940 (N_17940,N_1994,N_8692);
and U17941 (N_17941,N_3515,N_1944);
nand U17942 (N_17942,N_5916,N_5197);
nor U17943 (N_17943,N_4051,N_8907);
or U17944 (N_17944,N_4488,N_4899);
xnor U17945 (N_17945,N_5584,N_4397);
and U17946 (N_17946,N_2829,N_8514);
nand U17947 (N_17947,N_8385,N_8870);
nand U17948 (N_17948,N_4788,N_449);
or U17949 (N_17949,N_8982,N_3224);
and U17950 (N_17950,N_333,N_9079);
or U17951 (N_17951,N_5620,N_5974);
or U17952 (N_17952,N_5278,N_8395);
nor U17953 (N_17953,N_3520,N_4045);
and U17954 (N_17954,N_5906,N_3509);
nor U17955 (N_17955,N_7990,N_7739);
or U17956 (N_17956,N_4336,N_7535);
nand U17957 (N_17957,N_8412,N_4261);
or U17958 (N_17958,N_5058,N_3004);
nand U17959 (N_17959,N_7986,N_8418);
or U17960 (N_17960,N_4499,N_6510);
nand U17961 (N_17961,N_5518,N_4253);
nand U17962 (N_17962,N_6815,N_8742);
and U17963 (N_17963,N_878,N_642);
or U17964 (N_17964,N_4998,N_2550);
nand U17965 (N_17965,N_9701,N_151);
nand U17966 (N_17966,N_1996,N_6350);
nand U17967 (N_17967,N_3490,N_3589);
and U17968 (N_17968,N_2435,N_6762);
nand U17969 (N_17969,N_2340,N_6257);
nand U17970 (N_17970,N_2255,N_9764);
or U17971 (N_17971,N_8667,N_4600);
nor U17972 (N_17972,N_4862,N_4760);
and U17973 (N_17973,N_1467,N_9952);
nand U17974 (N_17974,N_2154,N_9301);
or U17975 (N_17975,N_1227,N_7060);
and U17976 (N_17976,N_5161,N_9448);
or U17977 (N_17977,N_9340,N_1364);
or U17978 (N_17978,N_8480,N_7766);
nor U17979 (N_17979,N_9655,N_568);
or U17980 (N_17980,N_6451,N_7755);
and U17981 (N_17981,N_7091,N_7875);
nand U17982 (N_17982,N_417,N_2258);
and U17983 (N_17983,N_1674,N_4248);
or U17984 (N_17984,N_8982,N_7290);
or U17985 (N_17985,N_2309,N_3742);
and U17986 (N_17986,N_7133,N_6439);
and U17987 (N_17987,N_6865,N_3004);
and U17988 (N_17988,N_329,N_1972);
or U17989 (N_17989,N_317,N_8977);
xor U17990 (N_17990,N_4854,N_9599);
or U17991 (N_17991,N_4118,N_2630);
nor U17992 (N_17992,N_4273,N_1826);
or U17993 (N_17993,N_6118,N_9357);
and U17994 (N_17994,N_5938,N_2262);
nand U17995 (N_17995,N_1795,N_5173);
and U17996 (N_17996,N_7138,N_2228);
xor U17997 (N_17997,N_3226,N_5566);
or U17998 (N_17998,N_7491,N_2234);
or U17999 (N_17999,N_7874,N_4206);
nand U18000 (N_18000,N_7232,N_3425);
nor U18001 (N_18001,N_4372,N_4719);
nor U18002 (N_18002,N_1339,N_8956);
or U18003 (N_18003,N_7125,N_7333);
and U18004 (N_18004,N_6718,N_156);
and U18005 (N_18005,N_7033,N_4319);
nor U18006 (N_18006,N_9965,N_9024);
nor U18007 (N_18007,N_4246,N_4737);
and U18008 (N_18008,N_6331,N_2814);
and U18009 (N_18009,N_5792,N_7325);
xnor U18010 (N_18010,N_3031,N_7371);
nor U18011 (N_18011,N_7757,N_3492);
or U18012 (N_18012,N_4258,N_583);
nor U18013 (N_18013,N_5365,N_1000);
nand U18014 (N_18014,N_1064,N_273);
or U18015 (N_18015,N_3223,N_7010);
nor U18016 (N_18016,N_6016,N_1730);
or U18017 (N_18017,N_4912,N_1485);
and U18018 (N_18018,N_1190,N_2105);
nor U18019 (N_18019,N_7565,N_4301);
nand U18020 (N_18020,N_4756,N_2605);
and U18021 (N_18021,N_8789,N_2459);
nand U18022 (N_18022,N_1240,N_4368);
nand U18023 (N_18023,N_9578,N_7998);
xor U18024 (N_18024,N_9301,N_9466);
or U18025 (N_18025,N_9793,N_9198);
nor U18026 (N_18026,N_8562,N_5940);
nand U18027 (N_18027,N_4346,N_2324);
nor U18028 (N_18028,N_1219,N_4520);
nand U18029 (N_18029,N_5260,N_7389);
xnor U18030 (N_18030,N_3018,N_4635);
or U18031 (N_18031,N_994,N_8624);
xnor U18032 (N_18032,N_4729,N_628);
nand U18033 (N_18033,N_1076,N_329);
or U18034 (N_18034,N_5617,N_8891);
and U18035 (N_18035,N_6265,N_2179);
nand U18036 (N_18036,N_8944,N_9386);
and U18037 (N_18037,N_4735,N_7433);
xor U18038 (N_18038,N_4513,N_3670);
and U18039 (N_18039,N_6300,N_4386);
nand U18040 (N_18040,N_565,N_2801);
and U18041 (N_18041,N_2456,N_6987);
nand U18042 (N_18042,N_1174,N_7780);
nor U18043 (N_18043,N_7694,N_2127);
and U18044 (N_18044,N_543,N_8003);
or U18045 (N_18045,N_2480,N_3950);
or U18046 (N_18046,N_8882,N_9303);
nor U18047 (N_18047,N_7202,N_5667);
nor U18048 (N_18048,N_5180,N_6774);
xor U18049 (N_18049,N_9288,N_3202);
and U18050 (N_18050,N_4742,N_9136);
or U18051 (N_18051,N_9205,N_6358);
or U18052 (N_18052,N_1469,N_5402);
xnor U18053 (N_18053,N_3692,N_1958);
and U18054 (N_18054,N_7942,N_2461);
nor U18055 (N_18055,N_980,N_7973);
and U18056 (N_18056,N_906,N_8599);
nor U18057 (N_18057,N_1985,N_4851);
xor U18058 (N_18058,N_9828,N_8998);
or U18059 (N_18059,N_403,N_3520);
xor U18060 (N_18060,N_8351,N_3329);
nor U18061 (N_18061,N_8119,N_5542);
nand U18062 (N_18062,N_422,N_1044);
and U18063 (N_18063,N_7693,N_6349);
or U18064 (N_18064,N_3837,N_3052);
nor U18065 (N_18065,N_8131,N_864);
and U18066 (N_18066,N_9914,N_2552);
nor U18067 (N_18067,N_5028,N_3452);
nor U18068 (N_18068,N_8436,N_867);
nand U18069 (N_18069,N_3136,N_8685);
or U18070 (N_18070,N_8678,N_724);
and U18071 (N_18071,N_9690,N_9466);
and U18072 (N_18072,N_5099,N_5091);
and U18073 (N_18073,N_854,N_9680);
and U18074 (N_18074,N_7702,N_7866);
and U18075 (N_18075,N_924,N_1690);
or U18076 (N_18076,N_3428,N_6931);
or U18077 (N_18077,N_6589,N_9389);
xor U18078 (N_18078,N_8352,N_7502);
xor U18079 (N_18079,N_8403,N_9139);
and U18080 (N_18080,N_3346,N_8438);
or U18081 (N_18081,N_7167,N_5579);
or U18082 (N_18082,N_5049,N_8785);
nor U18083 (N_18083,N_6083,N_3014);
and U18084 (N_18084,N_8427,N_8374);
nor U18085 (N_18085,N_3818,N_6666);
and U18086 (N_18086,N_6253,N_5990);
nor U18087 (N_18087,N_1717,N_1813);
nand U18088 (N_18088,N_5740,N_6116);
xor U18089 (N_18089,N_5864,N_5863);
nor U18090 (N_18090,N_8038,N_2884);
nand U18091 (N_18091,N_9348,N_2363);
and U18092 (N_18092,N_1226,N_8320);
nor U18093 (N_18093,N_8188,N_7623);
nand U18094 (N_18094,N_3877,N_6017);
or U18095 (N_18095,N_9048,N_5530);
nor U18096 (N_18096,N_7402,N_4734);
or U18097 (N_18097,N_5767,N_1228);
or U18098 (N_18098,N_2203,N_7100);
and U18099 (N_18099,N_6846,N_6678);
nand U18100 (N_18100,N_688,N_5591);
and U18101 (N_18101,N_5261,N_4776);
and U18102 (N_18102,N_9465,N_8634);
or U18103 (N_18103,N_8184,N_9694);
nor U18104 (N_18104,N_627,N_8409);
nand U18105 (N_18105,N_402,N_1034);
xor U18106 (N_18106,N_324,N_609);
xnor U18107 (N_18107,N_7712,N_1049);
nand U18108 (N_18108,N_7410,N_4049);
or U18109 (N_18109,N_3771,N_7145);
nor U18110 (N_18110,N_2398,N_978);
and U18111 (N_18111,N_1561,N_5968);
nand U18112 (N_18112,N_1179,N_4922);
nand U18113 (N_18113,N_265,N_4104);
nand U18114 (N_18114,N_1865,N_1677);
and U18115 (N_18115,N_2383,N_2739);
and U18116 (N_18116,N_2082,N_6124);
xor U18117 (N_18117,N_5337,N_2768);
nor U18118 (N_18118,N_2934,N_7056);
or U18119 (N_18119,N_6846,N_3272);
xnor U18120 (N_18120,N_4845,N_3647);
or U18121 (N_18121,N_6389,N_4373);
and U18122 (N_18122,N_8954,N_2794);
and U18123 (N_18123,N_687,N_2907);
xor U18124 (N_18124,N_35,N_8097);
nor U18125 (N_18125,N_8146,N_6800);
or U18126 (N_18126,N_117,N_2925);
or U18127 (N_18127,N_6277,N_3217);
nor U18128 (N_18128,N_6521,N_1032);
or U18129 (N_18129,N_2340,N_479);
nor U18130 (N_18130,N_8117,N_3144);
nand U18131 (N_18131,N_5945,N_9735);
and U18132 (N_18132,N_7016,N_9981);
nor U18133 (N_18133,N_7982,N_8592);
xor U18134 (N_18134,N_9259,N_1016);
nor U18135 (N_18135,N_1544,N_1446);
xnor U18136 (N_18136,N_8179,N_482);
or U18137 (N_18137,N_2970,N_3281);
nand U18138 (N_18138,N_9639,N_4523);
and U18139 (N_18139,N_695,N_7301);
or U18140 (N_18140,N_4556,N_9228);
xor U18141 (N_18141,N_1000,N_5053);
or U18142 (N_18142,N_1367,N_5177);
or U18143 (N_18143,N_7540,N_2166);
nor U18144 (N_18144,N_1404,N_7971);
and U18145 (N_18145,N_3145,N_1904);
nor U18146 (N_18146,N_4618,N_7032);
xnor U18147 (N_18147,N_5897,N_5029);
nand U18148 (N_18148,N_6309,N_8974);
nor U18149 (N_18149,N_405,N_5519);
nor U18150 (N_18150,N_3244,N_7298);
nand U18151 (N_18151,N_7511,N_7182);
or U18152 (N_18152,N_3970,N_6929);
xor U18153 (N_18153,N_8721,N_1596);
xor U18154 (N_18154,N_2844,N_9998);
nand U18155 (N_18155,N_1201,N_2753);
and U18156 (N_18156,N_3858,N_6974);
nor U18157 (N_18157,N_972,N_8394);
and U18158 (N_18158,N_1379,N_4799);
or U18159 (N_18159,N_1255,N_2431);
nor U18160 (N_18160,N_2901,N_6902);
nor U18161 (N_18161,N_4711,N_8353);
nor U18162 (N_18162,N_8903,N_8740);
nor U18163 (N_18163,N_7827,N_9297);
nor U18164 (N_18164,N_3072,N_3089);
nand U18165 (N_18165,N_16,N_6018);
or U18166 (N_18166,N_9130,N_2507);
or U18167 (N_18167,N_7800,N_4877);
nor U18168 (N_18168,N_5593,N_6405);
nor U18169 (N_18169,N_4022,N_5409);
nor U18170 (N_18170,N_6077,N_5085);
xnor U18171 (N_18171,N_7366,N_4948);
and U18172 (N_18172,N_3701,N_3036);
nor U18173 (N_18173,N_4830,N_369);
nor U18174 (N_18174,N_9318,N_153);
or U18175 (N_18175,N_6816,N_1837);
and U18176 (N_18176,N_6769,N_1269);
nand U18177 (N_18177,N_4798,N_43);
or U18178 (N_18178,N_8840,N_5558);
or U18179 (N_18179,N_7098,N_2100);
or U18180 (N_18180,N_1131,N_8903);
or U18181 (N_18181,N_9999,N_8902);
xnor U18182 (N_18182,N_715,N_6024);
or U18183 (N_18183,N_9959,N_1824);
or U18184 (N_18184,N_1641,N_6465);
and U18185 (N_18185,N_4225,N_1996);
xnor U18186 (N_18186,N_2019,N_9262);
nand U18187 (N_18187,N_8649,N_9509);
nor U18188 (N_18188,N_3872,N_3063);
xor U18189 (N_18189,N_9408,N_4650);
and U18190 (N_18190,N_8288,N_8037);
nand U18191 (N_18191,N_9675,N_3182);
nand U18192 (N_18192,N_2792,N_8086);
and U18193 (N_18193,N_7514,N_5668);
or U18194 (N_18194,N_5396,N_2272);
and U18195 (N_18195,N_5623,N_9721);
xor U18196 (N_18196,N_6902,N_1963);
nand U18197 (N_18197,N_2120,N_2699);
or U18198 (N_18198,N_1955,N_6721);
nor U18199 (N_18199,N_1775,N_8902);
nor U18200 (N_18200,N_823,N_2009);
and U18201 (N_18201,N_7621,N_1740);
or U18202 (N_18202,N_9118,N_2831);
xor U18203 (N_18203,N_2443,N_5744);
and U18204 (N_18204,N_7693,N_7576);
nand U18205 (N_18205,N_111,N_1028);
nor U18206 (N_18206,N_1862,N_615);
and U18207 (N_18207,N_6533,N_5455);
nor U18208 (N_18208,N_7503,N_6698);
nand U18209 (N_18209,N_7809,N_3280);
nand U18210 (N_18210,N_7659,N_6003);
nand U18211 (N_18211,N_7495,N_4683);
nor U18212 (N_18212,N_7000,N_5998);
nand U18213 (N_18213,N_6406,N_342);
and U18214 (N_18214,N_2696,N_8627);
nand U18215 (N_18215,N_106,N_585);
or U18216 (N_18216,N_2165,N_2295);
or U18217 (N_18217,N_9369,N_3328);
and U18218 (N_18218,N_3292,N_5440);
nand U18219 (N_18219,N_525,N_6347);
xor U18220 (N_18220,N_458,N_4471);
nand U18221 (N_18221,N_7033,N_447);
nand U18222 (N_18222,N_961,N_7038);
or U18223 (N_18223,N_8405,N_72);
nor U18224 (N_18224,N_4814,N_8562);
nor U18225 (N_18225,N_2200,N_4837);
nor U18226 (N_18226,N_1293,N_3571);
or U18227 (N_18227,N_5395,N_8019);
nor U18228 (N_18228,N_3117,N_5437);
nor U18229 (N_18229,N_3962,N_5278);
nand U18230 (N_18230,N_3649,N_6266);
nand U18231 (N_18231,N_1879,N_6639);
and U18232 (N_18232,N_4416,N_5418);
or U18233 (N_18233,N_1729,N_9272);
xor U18234 (N_18234,N_9002,N_8302);
nor U18235 (N_18235,N_9905,N_76);
nand U18236 (N_18236,N_151,N_5921);
xnor U18237 (N_18237,N_1450,N_354);
or U18238 (N_18238,N_5276,N_5775);
nand U18239 (N_18239,N_4465,N_1624);
and U18240 (N_18240,N_3594,N_8500);
nand U18241 (N_18241,N_1588,N_3219);
and U18242 (N_18242,N_1325,N_4066);
or U18243 (N_18243,N_6233,N_807);
or U18244 (N_18244,N_7647,N_3975);
nand U18245 (N_18245,N_1070,N_2544);
or U18246 (N_18246,N_9090,N_3146);
xnor U18247 (N_18247,N_1975,N_7057);
nor U18248 (N_18248,N_7457,N_3060);
and U18249 (N_18249,N_2726,N_543);
nand U18250 (N_18250,N_5789,N_8921);
nor U18251 (N_18251,N_5011,N_6596);
nor U18252 (N_18252,N_2791,N_968);
nor U18253 (N_18253,N_8310,N_7616);
xnor U18254 (N_18254,N_7334,N_1283);
xnor U18255 (N_18255,N_6633,N_2062);
nor U18256 (N_18256,N_7355,N_6130);
nor U18257 (N_18257,N_9379,N_8783);
xor U18258 (N_18258,N_4951,N_4579);
or U18259 (N_18259,N_8141,N_7484);
nor U18260 (N_18260,N_8755,N_1743);
or U18261 (N_18261,N_930,N_3578);
xnor U18262 (N_18262,N_6030,N_9694);
nor U18263 (N_18263,N_479,N_1282);
and U18264 (N_18264,N_361,N_2937);
nand U18265 (N_18265,N_4107,N_6825);
nand U18266 (N_18266,N_4071,N_3552);
nand U18267 (N_18267,N_4030,N_9755);
nor U18268 (N_18268,N_3987,N_29);
nor U18269 (N_18269,N_4097,N_9763);
and U18270 (N_18270,N_147,N_2056);
and U18271 (N_18271,N_5647,N_4681);
nor U18272 (N_18272,N_4249,N_4257);
and U18273 (N_18273,N_7106,N_6367);
and U18274 (N_18274,N_4160,N_8417);
or U18275 (N_18275,N_6831,N_4466);
xnor U18276 (N_18276,N_7703,N_6800);
nand U18277 (N_18277,N_6572,N_2576);
or U18278 (N_18278,N_2808,N_6098);
xor U18279 (N_18279,N_1346,N_5212);
and U18280 (N_18280,N_2339,N_3772);
xor U18281 (N_18281,N_7156,N_472);
and U18282 (N_18282,N_5403,N_4010);
nor U18283 (N_18283,N_4698,N_7253);
nor U18284 (N_18284,N_1216,N_2910);
nor U18285 (N_18285,N_1515,N_6990);
or U18286 (N_18286,N_3817,N_2262);
nor U18287 (N_18287,N_2233,N_9872);
or U18288 (N_18288,N_1272,N_7308);
and U18289 (N_18289,N_1705,N_3110);
nor U18290 (N_18290,N_3761,N_6802);
nor U18291 (N_18291,N_5657,N_7135);
nand U18292 (N_18292,N_5977,N_2634);
or U18293 (N_18293,N_6025,N_2248);
nand U18294 (N_18294,N_9661,N_5479);
and U18295 (N_18295,N_7355,N_9615);
nor U18296 (N_18296,N_1684,N_2752);
nor U18297 (N_18297,N_3813,N_9340);
and U18298 (N_18298,N_7302,N_8024);
nand U18299 (N_18299,N_5230,N_7228);
nand U18300 (N_18300,N_1007,N_4416);
nand U18301 (N_18301,N_4255,N_5367);
nand U18302 (N_18302,N_77,N_255);
nand U18303 (N_18303,N_9824,N_4541);
xor U18304 (N_18304,N_3303,N_5498);
nor U18305 (N_18305,N_7405,N_2573);
and U18306 (N_18306,N_5681,N_7643);
or U18307 (N_18307,N_9006,N_9467);
nor U18308 (N_18308,N_9485,N_2339);
xor U18309 (N_18309,N_4219,N_5386);
nor U18310 (N_18310,N_1928,N_3782);
xnor U18311 (N_18311,N_3308,N_5315);
nand U18312 (N_18312,N_6467,N_9652);
xnor U18313 (N_18313,N_4397,N_3838);
or U18314 (N_18314,N_2952,N_7825);
nand U18315 (N_18315,N_3476,N_5898);
nor U18316 (N_18316,N_8580,N_3888);
nand U18317 (N_18317,N_7111,N_536);
nand U18318 (N_18318,N_5036,N_4057);
or U18319 (N_18319,N_8007,N_1076);
nand U18320 (N_18320,N_8723,N_9518);
or U18321 (N_18321,N_79,N_5509);
nor U18322 (N_18322,N_7541,N_297);
nand U18323 (N_18323,N_9351,N_9051);
nor U18324 (N_18324,N_654,N_8614);
and U18325 (N_18325,N_2879,N_9126);
xnor U18326 (N_18326,N_2067,N_4348);
nor U18327 (N_18327,N_41,N_9171);
nand U18328 (N_18328,N_3259,N_7146);
nor U18329 (N_18329,N_3890,N_5258);
nand U18330 (N_18330,N_5649,N_9805);
and U18331 (N_18331,N_4680,N_3245);
and U18332 (N_18332,N_356,N_341);
or U18333 (N_18333,N_2753,N_7694);
nand U18334 (N_18334,N_3745,N_8048);
xnor U18335 (N_18335,N_8227,N_922);
nand U18336 (N_18336,N_9854,N_7607);
nor U18337 (N_18337,N_5973,N_4931);
nor U18338 (N_18338,N_588,N_5032);
and U18339 (N_18339,N_1395,N_6627);
nor U18340 (N_18340,N_5848,N_9449);
or U18341 (N_18341,N_5168,N_4682);
xor U18342 (N_18342,N_581,N_7979);
nand U18343 (N_18343,N_5173,N_3001);
nor U18344 (N_18344,N_9217,N_621);
nor U18345 (N_18345,N_3951,N_8686);
nor U18346 (N_18346,N_4903,N_8922);
and U18347 (N_18347,N_7930,N_4158);
or U18348 (N_18348,N_9451,N_3885);
or U18349 (N_18349,N_7816,N_3085);
nand U18350 (N_18350,N_6696,N_1273);
nor U18351 (N_18351,N_9957,N_938);
nand U18352 (N_18352,N_3221,N_5871);
and U18353 (N_18353,N_1696,N_9839);
nor U18354 (N_18354,N_7007,N_7285);
xor U18355 (N_18355,N_3431,N_6591);
or U18356 (N_18356,N_1266,N_2739);
or U18357 (N_18357,N_1980,N_2989);
and U18358 (N_18358,N_3711,N_9334);
and U18359 (N_18359,N_1131,N_6775);
nor U18360 (N_18360,N_9117,N_3568);
or U18361 (N_18361,N_9059,N_1290);
xnor U18362 (N_18362,N_6123,N_7263);
or U18363 (N_18363,N_6829,N_5950);
nor U18364 (N_18364,N_7603,N_871);
nor U18365 (N_18365,N_8919,N_3722);
nand U18366 (N_18366,N_9994,N_2438);
and U18367 (N_18367,N_2718,N_4346);
nand U18368 (N_18368,N_1375,N_4234);
and U18369 (N_18369,N_2641,N_1575);
or U18370 (N_18370,N_2122,N_2272);
nand U18371 (N_18371,N_8322,N_1832);
nand U18372 (N_18372,N_338,N_2716);
nand U18373 (N_18373,N_6043,N_4349);
xor U18374 (N_18374,N_1350,N_7408);
and U18375 (N_18375,N_6462,N_2398);
or U18376 (N_18376,N_8297,N_3963);
nand U18377 (N_18377,N_8226,N_7037);
and U18378 (N_18378,N_308,N_1246);
and U18379 (N_18379,N_6329,N_7243);
nand U18380 (N_18380,N_1929,N_3655);
and U18381 (N_18381,N_1853,N_9063);
and U18382 (N_18382,N_9897,N_167);
and U18383 (N_18383,N_7378,N_2749);
nor U18384 (N_18384,N_5865,N_9525);
and U18385 (N_18385,N_6180,N_2217);
or U18386 (N_18386,N_5507,N_4591);
or U18387 (N_18387,N_4551,N_5887);
and U18388 (N_18388,N_2859,N_7666);
nand U18389 (N_18389,N_8264,N_1841);
xor U18390 (N_18390,N_6073,N_428);
nor U18391 (N_18391,N_1101,N_4606);
nor U18392 (N_18392,N_8438,N_8747);
nand U18393 (N_18393,N_8846,N_9485);
nor U18394 (N_18394,N_3698,N_6279);
or U18395 (N_18395,N_6858,N_3428);
and U18396 (N_18396,N_521,N_7584);
or U18397 (N_18397,N_3552,N_2294);
or U18398 (N_18398,N_6744,N_295);
nand U18399 (N_18399,N_8686,N_1877);
or U18400 (N_18400,N_3058,N_5871);
xor U18401 (N_18401,N_5660,N_416);
and U18402 (N_18402,N_5671,N_6731);
and U18403 (N_18403,N_903,N_5320);
and U18404 (N_18404,N_4234,N_9899);
or U18405 (N_18405,N_7844,N_8164);
xnor U18406 (N_18406,N_2300,N_9773);
nand U18407 (N_18407,N_6225,N_3800);
nor U18408 (N_18408,N_1638,N_6941);
nand U18409 (N_18409,N_8065,N_568);
or U18410 (N_18410,N_6023,N_9503);
and U18411 (N_18411,N_9747,N_9625);
nor U18412 (N_18412,N_4042,N_2214);
and U18413 (N_18413,N_6357,N_5932);
and U18414 (N_18414,N_1107,N_2096);
or U18415 (N_18415,N_708,N_6602);
nand U18416 (N_18416,N_4992,N_8802);
or U18417 (N_18417,N_1790,N_2254);
and U18418 (N_18418,N_174,N_5133);
nand U18419 (N_18419,N_9182,N_1427);
and U18420 (N_18420,N_7417,N_4086);
nand U18421 (N_18421,N_7831,N_1801);
or U18422 (N_18422,N_1798,N_5675);
and U18423 (N_18423,N_5332,N_8948);
nor U18424 (N_18424,N_2934,N_6883);
and U18425 (N_18425,N_668,N_2929);
nor U18426 (N_18426,N_7573,N_3164);
nand U18427 (N_18427,N_4522,N_7137);
and U18428 (N_18428,N_3268,N_7112);
nand U18429 (N_18429,N_4816,N_5823);
nand U18430 (N_18430,N_387,N_3381);
xnor U18431 (N_18431,N_2458,N_3745);
nor U18432 (N_18432,N_7163,N_151);
xnor U18433 (N_18433,N_6465,N_5278);
or U18434 (N_18434,N_3529,N_8429);
nor U18435 (N_18435,N_3496,N_9449);
and U18436 (N_18436,N_9244,N_939);
nand U18437 (N_18437,N_4295,N_8345);
nand U18438 (N_18438,N_8216,N_9770);
and U18439 (N_18439,N_7776,N_9136);
nand U18440 (N_18440,N_4518,N_5715);
xnor U18441 (N_18441,N_4496,N_8121);
or U18442 (N_18442,N_7575,N_8924);
or U18443 (N_18443,N_9396,N_277);
and U18444 (N_18444,N_3952,N_4113);
nor U18445 (N_18445,N_3595,N_1635);
nand U18446 (N_18446,N_1357,N_6756);
xor U18447 (N_18447,N_940,N_441);
nand U18448 (N_18448,N_4975,N_4514);
nand U18449 (N_18449,N_5121,N_6516);
nand U18450 (N_18450,N_3072,N_5164);
or U18451 (N_18451,N_1938,N_8243);
nor U18452 (N_18452,N_2682,N_7030);
or U18453 (N_18453,N_6104,N_6524);
or U18454 (N_18454,N_8774,N_5635);
nor U18455 (N_18455,N_3311,N_7381);
and U18456 (N_18456,N_8659,N_809);
and U18457 (N_18457,N_5484,N_1739);
or U18458 (N_18458,N_594,N_6708);
nand U18459 (N_18459,N_8966,N_4290);
and U18460 (N_18460,N_2547,N_2700);
or U18461 (N_18461,N_5089,N_8862);
or U18462 (N_18462,N_216,N_6024);
nor U18463 (N_18463,N_6414,N_2675);
nor U18464 (N_18464,N_9610,N_6928);
nand U18465 (N_18465,N_1979,N_3934);
or U18466 (N_18466,N_4613,N_4790);
xnor U18467 (N_18467,N_9646,N_22);
nor U18468 (N_18468,N_2749,N_1303);
and U18469 (N_18469,N_5196,N_1793);
nor U18470 (N_18470,N_3340,N_9827);
nand U18471 (N_18471,N_945,N_710);
and U18472 (N_18472,N_696,N_328);
nand U18473 (N_18473,N_8666,N_5974);
or U18474 (N_18474,N_340,N_44);
xor U18475 (N_18475,N_8647,N_6449);
and U18476 (N_18476,N_3422,N_5345);
or U18477 (N_18477,N_6979,N_9389);
nand U18478 (N_18478,N_3489,N_7301);
or U18479 (N_18479,N_4787,N_6171);
and U18480 (N_18480,N_6983,N_220);
or U18481 (N_18481,N_1574,N_8630);
nand U18482 (N_18482,N_1278,N_8700);
or U18483 (N_18483,N_1350,N_7131);
and U18484 (N_18484,N_1560,N_3184);
and U18485 (N_18485,N_6409,N_5476);
or U18486 (N_18486,N_9911,N_3206);
nor U18487 (N_18487,N_3798,N_5273);
and U18488 (N_18488,N_3518,N_2440);
or U18489 (N_18489,N_3899,N_7407);
nor U18490 (N_18490,N_9274,N_3248);
nand U18491 (N_18491,N_3949,N_2501);
nand U18492 (N_18492,N_1451,N_4536);
and U18493 (N_18493,N_6010,N_7560);
or U18494 (N_18494,N_4335,N_6331);
nor U18495 (N_18495,N_1731,N_8201);
or U18496 (N_18496,N_5101,N_2604);
nor U18497 (N_18497,N_9672,N_9026);
and U18498 (N_18498,N_6117,N_3074);
nor U18499 (N_18499,N_7642,N_5172);
nor U18500 (N_18500,N_8996,N_4371);
nor U18501 (N_18501,N_889,N_9983);
nor U18502 (N_18502,N_8645,N_7757);
or U18503 (N_18503,N_8063,N_2111);
nor U18504 (N_18504,N_6924,N_8041);
or U18505 (N_18505,N_117,N_523);
nor U18506 (N_18506,N_8062,N_4452);
nor U18507 (N_18507,N_1900,N_5208);
nor U18508 (N_18508,N_443,N_4273);
nand U18509 (N_18509,N_5827,N_5809);
or U18510 (N_18510,N_2290,N_829);
nor U18511 (N_18511,N_4840,N_653);
xnor U18512 (N_18512,N_1309,N_2254);
or U18513 (N_18513,N_6566,N_249);
nand U18514 (N_18514,N_97,N_2713);
nand U18515 (N_18515,N_8018,N_8224);
xnor U18516 (N_18516,N_8450,N_867);
nand U18517 (N_18517,N_8995,N_2834);
or U18518 (N_18518,N_6980,N_484);
nand U18519 (N_18519,N_6565,N_2566);
xnor U18520 (N_18520,N_3634,N_2699);
and U18521 (N_18521,N_7130,N_5307);
and U18522 (N_18522,N_3560,N_8566);
and U18523 (N_18523,N_2190,N_5222);
and U18524 (N_18524,N_6131,N_6616);
nand U18525 (N_18525,N_2436,N_2980);
xor U18526 (N_18526,N_1875,N_5000);
and U18527 (N_18527,N_2884,N_3732);
nand U18528 (N_18528,N_2300,N_2660);
nor U18529 (N_18529,N_3167,N_9973);
nand U18530 (N_18530,N_386,N_5166);
or U18531 (N_18531,N_7887,N_5572);
nand U18532 (N_18532,N_6503,N_667);
xor U18533 (N_18533,N_418,N_7577);
nor U18534 (N_18534,N_4558,N_5708);
nand U18535 (N_18535,N_8296,N_5139);
or U18536 (N_18536,N_1116,N_3674);
or U18537 (N_18537,N_5559,N_5756);
nor U18538 (N_18538,N_1103,N_7117);
or U18539 (N_18539,N_5244,N_2431);
or U18540 (N_18540,N_5113,N_744);
nand U18541 (N_18541,N_130,N_2546);
and U18542 (N_18542,N_4213,N_2499);
nor U18543 (N_18543,N_17,N_9149);
xor U18544 (N_18544,N_1980,N_5785);
or U18545 (N_18545,N_7793,N_5746);
or U18546 (N_18546,N_5023,N_7785);
nor U18547 (N_18547,N_2909,N_70);
or U18548 (N_18548,N_6844,N_1804);
xor U18549 (N_18549,N_3055,N_2708);
nand U18550 (N_18550,N_9087,N_7005);
or U18551 (N_18551,N_7728,N_9598);
or U18552 (N_18552,N_9008,N_320);
and U18553 (N_18553,N_8687,N_2088);
nand U18554 (N_18554,N_2765,N_9431);
or U18555 (N_18555,N_2896,N_952);
nor U18556 (N_18556,N_3950,N_3126);
and U18557 (N_18557,N_8918,N_4665);
xnor U18558 (N_18558,N_9919,N_9256);
and U18559 (N_18559,N_1019,N_4267);
nor U18560 (N_18560,N_7268,N_4493);
nor U18561 (N_18561,N_7921,N_6302);
and U18562 (N_18562,N_5808,N_3421);
nand U18563 (N_18563,N_1361,N_168);
and U18564 (N_18564,N_9457,N_1651);
nand U18565 (N_18565,N_6804,N_5401);
and U18566 (N_18566,N_4719,N_9887);
nor U18567 (N_18567,N_3057,N_3138);
nand U18568 (N_18568,N_7410,N_2482);
nand U18569 (N_18569,N_4663,N_7803);
or U18570 (N_18570,N_4783,N_2968);
and U18571 (N_18571,N_3733,N_5110);
or U18572 (N_18572,N_5505,N_4860);
nor U18573 (N_18573,N_1304,N_7004);
or U18574 (N_18574,N_9265,N_6801);
and U18575 (N_18575,N_2338,N_4619);
nor U18576 (N_18576,N_4009,N_6117);
nor U18577 (N_18577,N_3412,N_8072);
nor U18578 (N_18578,N_1550,N_1332);
and U18579 (N_18579,N_9396,N_1039);
xor U18580 (N_18580,N_9721,N_2642);
nor U18581 (N_18581,N_2697,N_9349);
xnor U18582 (N_18582,N_9735,N_1849);
xor U18583 (N_18583,N_3303,N_7601);
or U18584 (N_18584,N_9107,N_4301);
or U18585 (N_18585,N_9445,N_8494);
and U18586 (N_18586,N_8889,N_591);
and U18587 (N_18587,N_6080,N_5534);
nand U18588 (N_18588,N_4103,N_9025);
or U18589 (N_18589,N_6536,N_4490);
or U18590 (N_18590,N_4601,N_3639);
nand U18591 (N_18591,N_1952,N_9486);
and U18592 (N_18592,N_84,N_7582);
nand U18593 (N_18593,N_7278,N_9541);
nand U18594 (N_18594,N_3541,N_5788);
or U18595 (N_18595,N_2652,N_183);
or U18596 (N_18596,N_1571,N_158);
nor U18597 (N_18597,N_4808,N_7292);
nand U18598 (N_18598,N_5028,N_8592);
nand U18599 (N_18599,N_3929,N_2640);
nand U18600 (N_18600,N_1210,N_9695);
nand U18601 (N_18601,N_212,N_5997);
nand U18602 (N_18602,N_8212,N_1472);
and U18603 (N_18603,N_2184,N_7766);
nand U18604 (N_18604,N_3386,N_7591);
xor U18605 (N_18605,N_9052,N_9165);
or U18606 (N_18606,N_6241,N_3795);
and U18607 (N_18607,N_6622,N_3561);
and U18608 (N_18608,N_6821,N_3996);
or U18609 (N_18609,N_2681,N_8804);
or U18610 (N_18610,N_5350,N_333);
and U18611 (N_18611,N_1234,N_8026);
nor U18612 (N_18612,N_9697,N_5921);
xor U18613 (N_18613,N_9038,N_3715);
and U18614 (N_18614,N_7513,N_8754);
xnor U18615 (N_18615,N_2399,N_6609);
nor U18616 (N_18616,N_3368,N_7312);
or U18617 (N_18617,N_7835,N_6019);
xor U18618 (N_18618,N_4969,N_8998);
xnor U18619 (N_18619,N_3296,N_8818);
or U18620 (N_18620,N_1834,N_592);
or U18621 (N_18621,N_7810,N_6657);
xor U18622 (N_18622,N_4557,N_6403);
and U18623 (N_18623,N_268,N_3902);
nor U18624 (N_18624,N_6219,N_3109);
nand U18625 (N_18625,N_9425,N_7120);
or U18626 (N_18626,N_9294,N_409);
and U18627 (N_18627,N_7724,N_2934);
and U18628 (N_18628,N_325,N_3253);
nor U18629 (N_18629,N_7099,N_3528);
nor U18630 (N_18630,N_7764,N_8789);
nand U18631 (N_18631,N_5860,N_2320);
or U18632 (N_18632,N_8428,N_4237);
and U18633 (N_18633,N_9056,N_8197);
xor U18634 (N_18634,N_1846,N_3745);
nor U18635 (N_18635,N_7030,N_7092);
nand U18636 (N_18636,N_7063,N_4271);
and U18637 (N_18637,N_2076,N_662);
and U18638 (N_18638,N_4068,N_2396);
and U18639 (N_18639,N_4410,N_2551);
nor U18640 (N_18640,N_2092,N_2646);
xor U18641 (N_18641,N_246,N_465);
and U18642 (N_18642,N_8461,N_1275);
nor U18643 (N_18643,N_3829,N_3452);
and U18644 (N_18644,N_2909,N_5862);
nand U18645 (N_18645,N_9045,N_7431);
nor U18646 (N_18646,N_5926,N_7214);
and U18647 (N_18647,N_8251,N_7031);
or U18648 (N_18648,N_5045,N_2018);
and U18649 (N_18649,N_7019,N_370);
nand U18650 (N_18650,N_5632,N_9457);
or U18651 (N_18651,N_7391,N_4427);
or U18652 (N_18652,N_8829,N_7434);
nand U18653 (N_18653,N_1404,N_3317);
nor U18654 (N_18654,N_3855,N_5363);
and U18655 (N_18655,N_6644,N_7451);
nor U18656 (N_18656,N_4133,N_2935);
nand U18657 (N_18657,N_1387,N_9721);
or U18658 (N_18658,N_3617,N_1015);
nor U18659 (N_18659,N_2381,N_3365);
nand U18660 (N_18660,N_3985,N_1979);
nand U18661 (N_18661,N_5078,N_2019);
nand U18662 (N_18662,N_568,N_5519);
xor U18663 (N_18663,N_1401,N_9800);
nand U18664 (N_18664,N_2818,N_8952);
and U18665 (N_18665,N_2478,N_4753);
and U18666 (N_18666,N_3497,N_7457);
xnor U18667 (N_18667,N_9649,N_3658);
nand U18668 (N_18668,N_3081,N_3770);
and U18669 (N_18669,N_4662,N_1747);
nand U18670 (N_18670,N_6042,N_4496);
nor U18671 (N_18671,N_8981,N_2653);
and U18672 (N_18672,N_7155,N_7326);
or U18673 (N_18673,N_4701,N_1590);
nand U18674 (N_18674,N_6327,N_5636);
nand U18675 (N_18675,N_4962,N_6412);
xnor U18676 (N_18676,N_9535,N_2918);
xnor U18677 (N_18677,N_6227,N_1127);
and U18678 (N_18678,N_4547,N_7368);
or U18679 (N_18679,N_7943,N_533);
nor U18680 (N_18680,N_7394,N_2733);
and U18681 (N_18681,N_8872,N_9762);
nand U18682 (N_18682,N_9758,N_61);
or U18683 (N_18683,N_6075,N_3886);
nand U18684 (N_18684,N_3236,N_177);
nand U18685 (N_18685,N_8070,N_6466);
or U18686 (N_18686,N_3797,N_1316);
or U18687 (N_18687,N_7783,N_7453);
xnor U18688 (N_18688,N_1813,N_9311);
or U18689 (N_18689,N_1225,N_1072);
nor U18690 (N_18690,N_2603,N_4105);
nand U18691 (N_18691,N_7195,N_5157);
nor U18692 (N_18692,N_366,N_4736);
and U18693 (N_18693,N_1772,N_3316);
or U18694 (N_18694,N_2435,N_7970);
nand U18695 (N_18695,N_3021,N_1911);
nand U18696 (N_18696,N_3944,N_2604);
and U18697 (N_18697,N_6693,N_9801);
xnor U18698 (N_18698,N_3937,N_8191);
nand U18699 (N_18699,N_8178,N_1149);
and U18700 (N_18700,N_717,N_2698);
and U18701 (N_18701,N_1302,N_1237);
or U18702 (N_18702,N_2507,N_7404);
nor U18703 (N_18703,N_2667,N_979);
or U18704 (N_18704,N_6291,N_6740);
nand U18705 (N_18705,N_3548,N_2288);
or U18706 (N_18706,N_7352,N_6298);
or U18707 (N_18707,N_3532,N_9845);
nor U18708 (N_18708,N_3519,N_9701);
nor U18709 (N_18709,N_3476,N_1181);
nand U18710 (N_18710,N_5830,N_5847);
or U18711 (N_18711,N_7311,N_8798);
or U18712 (N_18712,N_9202,N_337);
or U18713 (N_18713,N_4269,N_137);
xor U18714 (N_18714,N_3507,N_4243);
xnor U18715 (N_18715,N_1330,N_4954);
nand U18716 (N_18716,N_6324,N_2420);
nand U18717 (N_18717,N_9830,N_1705);
and U18718 (N_18718,N_5919,N_2428);
nor U18719 (N_18719,N_5492,N_5265);
nand U18720 (N_18720,N_3706,N_2247);
or U18721 (N_18721,N_412,N_3286);
and U18722 (N_18722,N_2535,N_8303);
and U18723 (N_18723,N_5629,N_4032);
nor U18724 (N_18724,N_6752,N_2861);
or U18725 (N_18725,N_8070,N_4296);
and U18726 (N_18726,N_3801,N_5419);
nor U18727 (N_18727,N_8266,N_4726);
nor U18728 (N_18728,N_9566,N_1524);
and U18729 (N_18729,N_5902,N_4457);
xor U18730 (N_18730,N_5364,N_1926);
or U18731 (N_18731,N_5707,N_5479);
or U18732 (N_18732,N_9376,N_304);
or U18733 (N_18733,N_1981,N_7832);
and U18734 (N_18734,N_1821,N_1857);
and U18735 (N_18735,N_3835,N_3888);
nand U18736 (N_18736,N_6254,N_4826);
and U18737 (N_18737,N_724,N_8684);
and U18738 (N_18738,N_151,N_639);
and U18739 (N_18739,N_3284,N_7270);
nand U18740 (N_18740,N_6149,N_4752);
nand U18741 (N_18741,N_3058,N_2183);
and U18742 (N_18742,N_7646,N_6846);
nand U18743 (N_18743,N_1358,N_1951);
xor U18744 (N_18744,N_4232,N_3836);
and U18745 (N_18745,N_7572,N_2808);
and U18746 (N_18746,N_6213,N_3668);
and U18747 (N_18747,N_1698,N_1437);
nand U18748 (N_18748,N_1467,N_9965);
nand U18749 (N_18749,N_3,N_6479);
nand U18750 (N_18750,N_9942,N_8125);
nand U18751 (N_18751,N_127,N_3136);
nor U18752 (N_18752,N_7367,N_1837);
nor U18753 (N_18753,N_8985,N_6705);
and U18754 (N_18754,N_4449,N_231);
and U18755 (N_18755,N_8492,N_1258);
nor U18756 (N_18756,N_853,N_5020);
nor U18757 (N_18757,N_7235,N_5703);
nand U18758 (N_18758,N_7450,N_7161);
nand U18759 (N_18759,N_8806,N_288);
xor U18760 (N_18760,N_1497,N_1808);
or U18761 (N_18761,N_3551,N_5084);
xor U18762 (N_18762,N_3146,N_8646);
nor U18763 (N_18763,N_6023,N_1906);
xor U18764 (N_18764,N_6411,N_923);
nand U18765 (N_18765,N_4430,N_2926);
xor U18766 (N_18766,N_3611,N_3367);
or U18767 (N_18767,N_8762,N_7649);
or U18768 (N_18768,N_4352,N_8557);
nand U18769 (N_18769,N_7953,N_2234);
or U18770 (N_18770,N_2597,N_9404);
nor U18771 (N_18771,N_8162,N_5773);
and U18772 (N_18772,N_2722,N_7500);
nand U18773 (N_18773,N_2265,N_1111);
xor U18774 (N_18774,N_8533,N_9505);
and U18775 (N_18775,N_8250,N_9390);
xnor U18776 (N_18776,N_7297,N_9779);
nor U18777 (N_18777,N_7894,N_1624);
nor U18778 (N_18778,N_9977,N_2330);
or U18779 (N_18779,N_5031,N_1307);
nor U18780 (N_18780,N_1973,N_2016);
nand U18781 (N_18781,N_2985,N_3397);
and U18782 (N_18782,N_5740,N_4289);
nand U18783 (N_18783,N_5171,N_6399);
nor U18784 (N_18784,N_8560,N_2111);
nand U18785 (N_18785,N_969,N_7580);
and U18786 (N_18786,N_5936,N_3749);
xor U18787 (N_18787,N_7467,N_936);
or U18788 (N_18788,N_299,N_8341);
and U18789 (N_18789,N_566,N_7398);
or U18790 (N_18790,N_38,N_2215);
and U18791 (N_18791,N_6732,N_597);
nor U18792 (N_18792,N_2169,N_4665);
nor U18793 (N_18793,N_5730,N_4173);
nand U18794 (N_18794,N_2684,N_8342);
and U18795 (N_18795,N_9424,N_1055);
nor U18796 (N_18796,N_1307,N_5365);
nand U18797 (N_18797,N_1659,N_1491);
nor U18798 (N_18798,N_4469,N_5066);
and U18799 (N_18799,N_7759,N_2373);
nor U18800 (N_18800,N_3801,N_7068);
nor U18801 (N_18801,N_9633,N_5384);
nor U18802 (N_18802,N_4231,N_7116);
or U18803 (N_18803,N_2115,N_692);
or U18804 (N_18804,N_5537,N_8975);
nand U18805 (N_18805,N_2529,N_6926);
nand U18806 (N_18806,N_5589,N_2304);
or U18807 (N_18807,N_6519,N_6629);
and U18808 (N_18808,N_3706,N_4017);
and U18809 (N_18809,N_6292,N_3363);
nand U18810 (N_18810,N_7421,N_5205);
and U18811 (N_18811,N_366,N_9996);
or U18812 (N_18812,N_2385,N_1209);
nand U18813 (N_18813,N_7612,N_4756);
nand U18814 (N_18814,N_712,N_5591);
and U18815 (N_18815,N_9424,N_1562);
nand U18816 (N_18816,N_9211,N_7405);
xor U18817 (N_18817,N_1755,N_5425);
nand U18818 (N_18818,N_6060,N_8973);
nor U18819 (N_18819,N_1077,N_1107);
and U18820 (N_18820,N_75,N_7681);
or U18821 (N_18821,N_7165,N_9366);
nand U18822 (N_18822,N_2913,N_8929);
nor U18823 (N_18823,N_8782,N_5317);
and U18824 (N_18824,N_5523,N_6779);
and U18825 (N_18825,N_4686,N_249);
xor U18826 (N_18826,N_8057,N_6293);
nand U18827 (N_18827,N_7631,N_2940);
nand U18828 (N_18828,N_856,N_4246);
nand U18829 (N_18829,N_6789,N_3816);
nor U18830 (N_18830,N_7140,N_8523);
nor U18831 (N_18831,N_9180,N_4868);
nor U18832 (N_18832,N_6453,N_1975);
or U18833 (N_18833,N_5783,N_6308);
nor U18834 (N_18834,N_1936,N_7150);
nand U18835 (N_18835,N_4727,N_3070);
and U18836 (N_18836,N_3868,N_1019);
nor U18837 (N_18837,N_7103,N_8201);
or U18838 (N_18838,N_5839,N_1549);
nand U18839 (N_18839,N_1694,N_4515);
xor U18840 (N_18840,N_4901,N_3698);
or U18841 (N_18841,N_1478,N_8109);
nand U18842 (N_18842,N_5428,N_3468);
nor U18843 (N_18843,N_737,N_5287);
or U18844 (N_18844,N_4991,N_9524);
or U18845 (N_18845,N_4907,N_5936);
nor U18846 (N_18846,N_2051,N_629);
nand U18847 (N_18847,N_3196,N_5155);
nor U18848 (N_18848,N_1303,N_8991);
nand U18849 (N_18849,N_4271,N_2762);
or U18850 (N_18850,N_162,N_4812);
and U18851 (N_18851,N_3137,N_3873);
xnor U18852 (N_18852,N_8847,N_2553);
and U18853 (N_18853,N_5365,N_4611);
nand U18854 (N_18854,N_5280,N_9209);
nand U18855 (N_18855,N_1287,N_7823);
or U18856 (N_18856,N_6972,N_6145);
and U18857 (N_18857,N_86,N_9571);
nand U18858 (N_18858,N_2756,N_6007);
nand U18859 (N_18859,N_9758,N_7492);
or U18860 (N_18860,N_5442,N_4350);
nand U18861 (N_18861,N_4114,N_4376);
and U18862 (N_18862,N_5450,N_2945);
nand U18863 (N_18863,N_289,N_6009);
and U18864 (N_18864,N_1859,N_1305);
nor U18865 (N_18865,N_8841,N_7962);
or U18866 (N_18866,N_7612,N_404);
nand U18867 (N_18867,N_9,N_5441);
nand U18868 (N_18868,N_1872,N_9099);
or U18869 (N_18869,N_8572,N_3351);
and U18870 (N_18870,N_4457,N_8050);
and U18871 (N_18871,N_4730,N_872);
or U18872 (N_18872,N_6575,N_6822);
and U18873 (N_18873,N_9451,N_5637);
xor U18874 (N_18874,N_9937,N_5433);
and U18875 (N_18875,N_2501,N_8657);
nand U18876 (N_18876,N_1633,N_8432);
or U18877 (N_18877,N_1008,N_1508);
nand U18878 (N_18878,N_3615,N_8341);
and U18879 (N_18879,N_5117,N_8974);
nand U18880 (N_18880,N_7565,N_4750);
and U18881 (N_18881,N_8009,N_375);
nor U18882 (N_18882,N_2768,N_5124);
nor U18883 (N_18883,N_2584,N_2545);
nor U18884 (N_18884,N_9053,N_748);
nor U18885 (N_18885,N_6415,N_2660);
and U18886 (N_18886,N_5421,N_104);
nor U18887 (N_18887,N_9331,N_431);
and U18888 (N_18888,N_8811,N_1492);
nand U18889 (N_18889,N_2545,N_5972);
nor U18890 (N_18890,N_4951,N_6636);
nor U18891 (N_18891,N_5565,N_8423);
nand U18892 (N_18892,N_6045,N_3276);
or U18893 (N_18893,N_2966,N_8388);
nor U18894 (N_18894,N_2092,N_5351);
and U18895 (N_18895,N_873,N_8118);
nand U18896 (N_18896,N_8981,N_7807);
and U18897 (N_18897,N_8236,N_2235);
or U18898 (N_18898,N_6413,N_5215);
and U18899 (N_18899,N_2484,N_6566);
nor U18900 (N_18900,N_4598,N_933);
nand U18901 (N_18901,N_710,N_7481);
or U18902 (N_18902,N_7661,N_7721);
and U18903 (N_18903,N_6377,N_1375);
or U18904 (N_18904,N_7150,N_7295);
and U18905 (N_18905,N_1698,N_9726);
or U18906 (N_18906,N_4836,N_517);
nor U18907 (N_18907,N_2240,N_4499);
xnor U18908 (N_18908,N_5358,N_6917);
and U18909 (N_18909,N_8582,N_9013);
and U18910 (N_18910,N_2948,N_2207);
nand U18911 (N_18911,N_8222,N_6944);
or U18912 (N_18912,N_5723,N_8534);
nand U18913 (N_18913,N_6350,N_9460);
or U18914 (N_18914,N_6590,N_4498);
nor U18915 (N_18915,N_4116,N_9536);
xnor U18916 (N_18916,N_6949,N_2340);
nand U18917 (N_18917,N_1450,N_3186);
and U18918 (N_18918,N_5523,N_6724);
or U18919 (N_18919,N_8252,N_737);
or U18920 (N_18920,N_9234,N_2448);
nor U18921 (N_18921,N_6327,N_5425);
or U18922 (N_18922,N_4898,N_7561);
and U18923 (N_18923,N_470,N_6835);
xor U18924 (N_18924,N_6935,N_8547);
nand U18925 (N_18925,N_3520,N_3484);
nor U18926 (N_18926,N_4052,N_6221);
and U18927 (N_18927,N_5340,N_9510);
or U18928 (N_18928,N_3976,N_3302);
xnor U18929 (N_18929,N_4597,N_713);
or U18930 (N_18930,N_5810,N_2111);
nor U18931 (N_18931,N_9257,N_4983);
nor U18932 (N_18932,N_8634,N_7081);
or U18933 (N_18933,N_5600,N_9311);
nor U18934 (N_18934,N_4118,N_9255);
nand U18935 (N_18935,N_5439,N_9174);
xnor U18936 (N_18936,N_2014,N_210);
and U18937 (N_18937,N_2705,N_7855);
xor U18938 (N_18938,N_4701,N_842);
nand U18939 (N_18939,N_4938,N_3054);
or U18940 (N_18940,N_2935,N_5902);
or U18941 (N_18941,N_9614,N_215);
nor U18942 (N_18942,N_9500,N_7750);
or U18943 (N_18943,N_9154,N_940);
nand U18944 (N_18944,N_5696,N_9891);
nor U18945 (N_18945,N_3971,N_1585);
and U18946 (N_18946,N_9166,N_1206);
or U18947 (N_18947,N_1988,N_4372);
and U18948 (N_18948,N_5415,N_3819);
nor U18949 (N_18949,N_5133,N_9525);
or U18950 (N_18950,N_3659,N_428);
nand U18951 (N_18951,N_2832,N_8878);
or U18952 (N_18952,N_1599,N_7392);
and U18953 (N_18953,N_3503,N_9619);
and U18954 (N_18954,N_1362,N_299);
and U18955 (N_18955,N_4227,N_5453);
and U18956 (N_18956,N_1037,N_3002);
nor U18957 (N_18957,N_9319,N_7009);
and U18958 (N_18958,N_8853,N_8134);
and U18959 (N_18959,N_2507,N_8119);
nand U18960 (N_18960,N_4846,N_123);
and U18961 (N_18961,N_5577,N_3619);
nor U18962 (N_18962,N_1932,N_2457);
nand U18963 (N_18963,N_5059,N_4868);
nor U18964 (N_18964,N_4393,N_5060);
or U18965 (N_18965,N_1809,N_5040);
and U18966 (N_18966,N_5076,N_7872);
xnor U18967 (N_18967,N_8831,N_9863);
nor U18968 (N_18968,N_8754,N_3404);
or U18969 (N_18969,N_2860,N_7301);
and U18970 (N_18970,N_6916,N_4572);
and U18971 (N_18971,N_5549,N_649);
or U18972 (N_18972,N_2012,N_6934);
or U18973 (N_18973,N_7289,N_8340);
or U18974 (N_18974,N_1010,N_8730);
and U18975 (N_18975,N_8437,N_7810);
xnor U18976 (N_18976,N_9911,N_3319);
nand U18977 (N_18977,N_7472,N_8637);
nand U18978 (N_18978,N_1962,N_4320);
nand U18979 (N_18979,N_1224,N_8248);
and U18980 (N_18980,N_6812,N_1156);
xnor U18981 (N_18981,N_6800,N_6875);
or U18982 (N_18982,N_493,N_5529);
nand U18983 (N_18983,N_6244,N_7046);
or U18984 (N_18984,N_3457,N_8318);
nand U18985 (N_18985,N_3559,N_6690);
nor U18986 (N_18986,N_6016,N_3581);
and U18987 (N_18987,N_7529,N_7439);
nand U18988 (N_18988,N_2875,N_6520);
or U18989 (N_18989,N_6991,N_6205);
xnor U18990 (N_18990,N_4750,N_2879);
nand U18991 (N_18991,N_2079,N_9925);
or U18992 (N_18992,N_5265,N_6751);
or U18993 (N_18993,N_4411,N_673);
and U18994 (N_18994,N_7385,N_2001);
nor U18995 (N_18995,N_4981,N_7240);
nor U18996 (N_18996,N_6235,N_9348);
or U18997 (N_18997,N_8407,N_9379);
and U18998 (N_18998,N_8473,N_4927);
or U18999 (N_18999,N_2898,N_6663);
nor U19000 (N_19000,N_7719,N_5784);
or U19001 (N_19001,N_5061,N_2330);
or U19002 (N_19002,N_9542,N_8964);
xor U19003 (N_19003,N_9982,N_7728);
and U19004 (N_19004,N_9817,N_3133);
xor U19005 (N_19005,N_5108,N_4355);
and U19006 (N_19006,N_6300,N_3310);
and U19007 (N_19007,N_927,N_5786);
nor U19008 (N_19008,N_5584,N_9310);
nand U19009 (N_19009,N_7871,N_8530);
or U19010 (N_19010,N_3522,N_480);
nor U19011 (N_19011,N_8675,N_8016);
or U19012 (N_19012,N_8341,N_7035);
nor U19013 (N_19013,N_3098,N_1065);
and U19014 (N_19014,N_5332,N_2725);
nand U19015 (N_19015,N_8599,N_5813);
nand U19016 (N_19016,N_7757,N_200);
or U19017 (N_19017,N_6804,N_5056);
and U19018 (N_19018,N_3126,N_3823);
nand U19019 (N_19019,N_4264,N_3324);
and U19020 (N_19020,N_5895,N_2318);
or U19021 (N_19021,N_1732,N_9938);
nand U19022 (N_19022,N_9393,N_4825);
nand U19023 (N_19023,N_7446,N_8550);
and U19024 (N_19024,N_9225,N_3401);
nor U19025 (N_19025,N_6833,N_4158);
or U19026 (N_19026,N_4145,N_3543);
xor U19027 (N_19027,N_1994,N_8412);
nand U19028 (N_19028,N_6956,N_9122);
or U19029 (N_19029,N_2724,N_5641);
or U19030 (N_19030,N_7483,N_1806);
or U19031 (N_19031,N_4210,N_9962);
or U19032 (N_19032,N_7260,N_3291);
nor U19033 (N_19033,N_2028,N_2615);
nor U19034 (N_19034,N_3549,N_1259);
nor U19035 (N_19035,N_5136,N_9315);
nand U19036 (N_19036,N_1434,N_9299);
nand U19037 (N_19037,N_4232,N_9500);
or U19038 (N_19038,N_928,N_2348);
or U19039 (N_19039,N_382,N_1620);
nor U19040 (N_19040,N_4084,N_9324);
nor U19041 (N_19041,N_6309,N_268);
and U19042 (N_19042,N_6846,N_4870);
and U19043 (N_19043,N_3965,N_6873);
or U19044 (N_19044,N_5046,N_3827);
or U19045 (N_19045,N_6455,N_3840);
nor U19046 (N_19046,N_431,N_383);
nor U19047 (N_19047,N_7710,N_1933);
or U19048 (N_19048,N_2878,N_9159);
nand U19049 (N_19049,N_6228,N_5386);
nor U19050 (N_19050,N_7401,N_568);
nand U19051 (N_19051,N_4757,N_9711);
or U19052 (N_19052,N_4123,N_1875);
nor U19053 (N_19053,N_6391,N_6627);
nand U19054 (N_19054,N_9389,N_6949);
and U19055 (N_19055,N_372,N_9648);
nor U19056 (N_19056,N_5273,N_8645);
and U19057 (N_19057,N_9915,N_2394);
nand U19058 (N_19058,N_2919,N_9681);
nor U19059 (N_19059,N_5106,N_2434);
or U19060 (N_19060,N_9866,N_3007);
or U19061 (N_19061,N_8643,N_127);
nor U19062 (N_19062,N_3559,N_7884);
or U19063 (N_19063,N_7462,N_206);
nand U19064 (N_19064,N_3828,N_4789);
nor U19065 (N_19065,N_2213,N_5161);
and U19066 (N_19066,N_2088,N_435);
and U19067 (N_19067,N_2606,N_8085);
or U19068 (N_19068,N_7691,N_4476);
nor U19069 (N_19069,N_6378,N_5574);
and U19070 (N_19070,N_2871,N_8649);
and U19071 (N_19071,N_2585,N_5169);
nand U19072 (N_19072,N_9871,N_2952);
xor U19073 (N_19073,N_2672,N_4434);
xnor U19074 (N_19074,N_578,N_4031);
nand U19075 (N_19075,N_109,N_5171);
or U19076 (N_19076,N_6597,N_3813);
nand U19077 (N_19077,N_5249,N_2805);
and U19078 (N_19078,N_4536,N_2935);
or U19079 (N_19079,N_5510,N_6880);
nand U19080 (N_19080,N_3963,N_5853);
or U19081 (N_19081,N_3244,N_9540);
nor U19082 (N_19082,N_854,N_234);
nor U19083 (N_19083,N_3628,N_7230);
and U19084 (N_19084,N_6450,N_3639);
or U19085 (N_19085,N_918,N_8335);
or U19086 (N_19086,N_2513,N_344);
or U19087 (N_19087,N_1414,N_9185);
and U19088 (N_19088,N_6741,N_7524);
or U19089 (N_19089,N_7042,N_1813);
or U19090 (N_19090,N_3239,N_6912);
and U19091 (N_19091,N_2519,N_1171);
nor U19092 (N_19092,N_8953,N_9296);
and U19093 (N_19093,N_8720,N_9961);
nand U19094 (N_19094,N_5421,N_5322);
and U19095 (N_19095,N_266,N_9919);
nor U19096 (N_19096,N_9526,N_8083);
or U19097 (N_19097,N_6639,N_238);
or U19098 (N_19098,N_1273,N_6758);
or U19099 (N_19099,N_4041,N_5756);
nor U19100 (N_19100,N_380,N_5753);
nand U19101 (N_19101,N_5832,N_1581);
nor U19102 (N_19102,N_554,N_3479);
or U19103 (N_19103,N_8356,N_2370);
nor U19104 (N_19104,N_7167,N_8841);
or U19105 (N_19105,N_5838,N_7962);
nand U19106 (N_19106,N_4053,N_4602);
nand U19107 (N_19107,N_5867,N_2079);
nand U19108 (N_19108,N_9121,N_5178);
and U19109 (N_19109,N_5522,N_3686);
nor U19110 (N_19110,N_132,N_977);
nand U19111 (N_19111,N_3175,N_9187);
nor U19112 (N_19112,N_9266,N_7030);
or U19113 (N_19113,N_4969,N_2869);
nand U19114 (N_19114,N_7544,N_8292);
or U19115 (N_19115,N_566,N_6204);
or U19116 (N_19116,N_334,N_8871);
and U19117 (N_19117,N_7962,N_8441);
and U19118 (N_19118,N_4424,N_4756);
and U19119 (N_19119,N_7059,N_7804);
and U19120 (N_19120,N_7959,N_3579);
nand U19121 (N_19121,N_9734,N_6892);
nor U19122 (N_19122,N_5753,N_1012);
nor U19123 (N_19123,N_1097,N_8335);
and U19124 (N_19124,N_7271,N_1722);
or U19125 (N_19125,N_7619,N_3375);
and U19126 (N_19126,N_819,N_9582);
xor U19127 (N_19127,N_2668,N_3060);
or U19128 (N_19128,N_6636,N_5399);
and U19129 (N_19129,N_2055,N_906);
nor U19130 (N_19130,N_3240,N_5089);
nor U19131 (N_19131,N_7385,N_5631);
and U19132 (N_19132,N_8155,N_4467);
nor U19133 (N_19133,N_491,N_9531);
or U19134 (N_19134,N_5726,N_6468);
and U19135 (N_19135,N_4412,N_4667);
nand U19136 (N_19136,N_737,N_9544);
nor U19137 (N_19137,N_9563,N_2591);
nand U19138 (N_19138,N_8508,N_9271);
nand U19139 (N_19139,N_3237,N_3742);
xnor U19140 (N_19140,N_7156,N_5617);
and U19141 (N_19141,N_2179,N_3808);
nand U19142 (N_19142,N_741,N_6814);
nor U19143 (N_19143,N_2311,N_8826);
or U19144 (N_19144,N_3741,N_6418);
nor U19145 (N_19145,N_5300,N_6637);
or U19146 (N_19146,N_5936,N_9700);
and U19147 (N_19147,N_3701,N_6631);
and U19148 (N_19148,N_4150,N_503);
or U19149 (N_19149,N_5409,N_6409);
xor U19150 (N_19150,N_2922,N_6104);
and U19151 (N_19151,N_8947,N_6807);
or U19152 (N_19152,N_8467,N_8760);
nand U19153 (N_19153,N_4852,N_6791);
or U19154 (N_19154,N_6742,N_7430);
xor U19155 (N_19155,N_5414,N_3170);
or U19156 (N_19156,N_9755,N_2319);
or U19157 (N_19157,N_2977,N_4529);
xor U19158 (N_19158,N_5800,N_380);
nand U19159 (N_19159,N_6251,N_4477);
nand U19160 (N_19160,N_3571,N_9343);
nand U19161 (N_19161,N_4478,N_9640);
xor U19162 (N_19162,N_6444,N_8950);
or U19163 (N_19163,N_7775,N_158);
or U19164 (N_19164,N_8263,N_8716);
or U19165 (N_19165,N_8881,N_4430);
nor U19166 (N_19166,N_9145,N_8584);
or U19167 (N_19167,N_9229,N_5328);
nor U19168 (N_19168,N_4848,N_8978);
nand U19169 (N_19169,N_7433,N_9519);
and U19170 (N_19170,N_3557,N_8904);
xnor U19171 (N_19171,N_3892,N_7087);
nor U19172 (N_19172,N_5758,N_5355);
nor U19173 (N_19173,N_897,N_9463);
nand U19174 (N_19174,N_6796,N_56);
nand U19175 (N_19175,N_3719,N_4893);
and U19176 (N_19176,N_671,N_4419);
nand U19177 (N_19177,N_5923,N_1965);
nand U19178 (N_19178,N_685,N_9894);
or U19179 (N_19179,N_7480,N_5686);
nor U19180 (N_19180,N_6418,N_2783);
or U19181 (N_19181,N_7946,N_677);
and U19182 (N_19182,N_2684,N_2757);
and U19183 (N_19183,N_3630,N_9705);
nor U19184 (N_19184,N_7850,N_2338);
and U19185 (N_19185,N_6163,N_6808);
nor U19186 (N_19186,N_6229,N_6682);
nand U19187 (N_19187,N_8208,N_1942);
and U19188 (N_19188,N_789,N_6891);
nor U19189 (N_19189,N_4870,N_1173);
and U19190 (N_19190,N_4170,N_8115);
and U19191 (N_19191,N_8296,N_1693);
nor U19192 (N_19192,N_4861,N_2880);
nor U19193 (N_19193,N_4375,N_3447);
or U19194 (N_19194,N_5862,N_1442);
nand U19195 (N_19195,N_8362,N_5520);
nor U19196 (N_19196,N_1367,N_5483);
xor U19197 (N_19197,N_9281,N_1855);
xnor U19198 (N_19198,N_8581,N_5662);
and U19199 (N_19199,N_3242,N_8126);
xor U19200 (N_19200,N_4161,N_1532);
and U19201 (N_19201,N_3478,N_5769);
nand U19202 (N_19202,N_361,N_6978);
and U19203 (N_19203,N_5440,N_9152);
xor U19204 (N_19204,N_3857,N_9234);
xnor U19205 (N_19205,N_5763,N_1092);
xnor U19206 (N_19206,N_172,N_3113);
nor U19207 (N_19207,N_8438,N_2411);
nand U19208 (N_19208,N_6534,N_7320);
nor U19209 (N_19209,N_2656,N_9938);
and U19210 (N_19210,N_955,N_6129);
nor U19211 (N_19211,N_1624,N_6800);
or U19212 (N_19212,N_9511,N_1360);
nor U19213 (N_19213,N_3655,N_7952);
or U19214 (N_19214,N_8317,N_2972);
nand U19215 (N_19215,N_4811,N_5854);
nor U19216 (N_19216,N_4912,N_1711);
nand U19217 (N_19217,N_3287,N_7913);
nor U19218 (N_19218,N_8314,N_6881);
and U19219 (N_19219,N_7626,N_8350);
nand U19220 (N_19220,N_4629,N_9351);
or U19221 (N_19221,N_5605,N_3693);
or U19222 (N_19222,N_6345,N_5353);
and U19223 (N_19223,N_1649,N_2779);
or U19224 (N_19224,N_1355,N_2016);
or U19225 (N_19225,N_3128,N_8984);
nand U19226 (N_19226,N_4709,N_257);
and U19227 (N_19227,N_9016,N_8304);
or U19228 (N_19228,N_4703,N_5626);
and U19229 (N_19229,N_3069,N_9405);
nor U19230 (N_19230,N_3213,N_7131);
or U19231 (N_19231,N_8200,N_2295);
and U19232 (N_19232,N_1781,N_3999);
nand U19233 (N_19233,N_9799,N_9242);
nor U19234 (N_19234,N_6346,N_5851);
or U19235 (N_19235,N_8339,N_2669);
nand U19236 (N_19236,N_996,N_6083);
nand U19237 (N_19237,N_6752,N_5496);
xnor U19238 (N_19238,N_94,N_2758);
nand U19239 (N_19239,N_8884,N_6421);
and U19240 (N_19240,N_3798,N_42);
nand U19241 (N_19241,N_2918,N_7176);
nand U19242 (N_19242,N_637,N_2629);
and U19243 (N_19243,N_1999,N_7713);
or U19244 (N_19244,N_6699,N_4607);
or U19245 (N_19245,N_7911,N_7757);
nand U19246 (N_19246,N_2791,N_4804);
nand U19247 (N_19247,N_5067,N_7617);
nor U19248 (N_19248,N_5775,N_8772);
xor U19249 (N_19249,N_3939,N_3255);
xor U19250 (N_19250,N_9584,N_5985);
or U19251 (N_19251,N_8443,N_6849);
nand U19252 (N_19252,N_3859,N_2975);
or U19253 (N_19253,N_6282,N_488);
and U19254 (N_19254,N_4184,N_2197);
and U19255 (N_19255,N_7173,N_591);
and U19256 (N_19256,N_153,N_9369);
nor U19257 (N_19257,N_6411,N_9463);
and U19258 (N_19258,N_5877,N_2595);
nand U19259 (N_19259,N_7682,N_8837);
nand U19260 (N_19260,N_5649,N_9345);
nor U19261 (N_19261,N_9749,N_5916);
or U19262 (N_19262,N_2295,N_8554);
or U19263 (N_19263,N_8300,N_7814);
nand U19264 (N_19264,N_915,N_7216);
nand U19265 (N_19265,N_771,N_1436);
and U19266 (N_19266,N_3171,N_2299);
nor U19267 (N_19267,N_1455,N_9369);
nor U19268 (N_19268,N_9831,N_9317);
or U19269 (N_19269,N_4501,N_6462);
or U19270 (N_19270,N_9199,N_5330);
and U19271 (N_19271,N_5087,N_3947);
nand U19272 (N_19272,N_8356,N_7579);
or U19273 (N_19273,N_2809,N_5379);
or U19274 (N_19274,N_2065,N_3680);
nor U19275 (N_19275,N_3168,N_6514);
or U19276 (N_19276,N_2685,N_693);
nor U19277 (N_19277,N_9578,N_2875);
and U19278 (N_19278,N_505,N_6701);
and U19279 (N_19279,N_5652,N_1427);
nor U19280 (N_19280,N_9224,N_3256);
and U19281 (N_19281,N_1499,N_7040);
and U19282 (N_19282,N_1553,N_7900);
nand U19283 (N_19283,N_583,N_3899);
nor U19284 (N_19284,N_9323,N_8438);
and U19285 (N_19285,N_4817,N_8971);
xnor U19286 (N_19286,N_5929,N_8191);
or U19287 (N_19287,N_3955,N_4165);
and U19288 (N_19288,N_6307,N_9224);
and U19289 (N_19289,N_7905,N_9067);
xnor U19290 (N_19290,N_6282,N_2628);
nand U19291 (N_19291,N_6178,N_7020);
or U19292 (N_19292,N_3290,N_6693);
nor U19293 (N_19293,N_6435,N_840);
nand U19294 (N_19294,N_31,N_7875);
nor U19295 (N_19295,N_4125,N_2787);
or U19296 (N_19296,N_5588,N_1117);
and U19297 (N_19297,N_1912,N_2529);
xnor U19298 (N_19298,N_895,N_4068);
nand U19299 (N_19299,N_9440,N_3139);
nor U19300 (N_19300,N_5588,N_638);
and U19301 (N_19301,N_2238,N_7134);
nand U19302 (N_19302,N_5453,N_7455);
and U19303 (N_19303,N_4110,N_3383);
nand U19304 (N_19304,N_1655,N_9047);
and U19305 (N_19305,N_4599,N_518);
or U19306 (N_19306,N_6720,N_3726);
and U19307 (N_19307,N_7808,N_5066);
and U19308 (N_19308,N_3929,N_1401);
and U19309 (N_19309,N_3121,N_4129);
nor U19310 (N_19310,N_7950,N_3578);
nor U19311 (N_19311,N_7964,N_2766);
xor U19312 (N_19312,N_6826,N_1796);
and U19313 (N_19313,N_6351,N_9150);
nor U19314 (N_19314,N_8907,N_9911);
or U19315 (N_19315,N_711,N_8787);
or U19316 (N_19316,N_6455,N_7167);
or U19317 (N_19317,N_9326,N_1208);
nand U19318 (N_19318,N_8899,N_3696);
nor U19319 (N_19319,N_6135,N_3838);
and U19320 (N_19320,N_2306,N_605);
and U19321 (N_19321,N_4536,N_918);
or U19322 (N_19322,N_533,N_5685);
and U19323 (N_19323,N_5038,N_8103);
and U19324 (N_19324,N_569,N_5655);
or U19325 (N_19325,N_5109,N_5558);
nand U19326 (N_19326,N_396,N_3440);
nor U19327 (N_19327,N_289,N_4614);
nor U19328 (N_19328,N_9300,N_6615);
and U19329 (N_19329,N_9959,N_4752);
or U19330 (N_19330,N_1348,N_1410);
nand U19331 (N_19331,N_8868,N_8982);
or U19332 (N_19332,N_5401,N_270);
and U19333 (N_19333,N_9816,N_6094);
nor U19334 (N_19334,N_4833,N_8294);
nand U19335 (N_19335,N_662,N_564);
and U19336 (N_19336,N_5212,N_8231);
or U19337 (N_19337,N_2496,N_8748);
nor U19338 (N_19338,N_5633,N_4644);
or U19339 (N_19339,N_3984,N_5505);
or U19340 (N_19340,N_6786,N_4184);
and U19341 (N_19341,N_8097,N_6606);
and U19342 (N_19342,N_1928,N_628);
xor U19343 (N_19343,N_1394,N_4253);
nand U19344 (N_19344,N_8219,N_8943);
xor U19345 (N_19345,N_6655,N_4921);
nor U19346 (N_19346,N_9146,N_8399);
and U19347 (N_19347,N_8474,N_1983);
nand U19348 (N_19348,N_9413,N_2136);
or U19349 (N_19349,N_2406,N_9592);
or U19350 (N_19350,N_8467,N_2459);
nand U19351 (N_19351,N_3181,N_3629);
or U19352 (N_19352,N_5236,N_5768);
or U19353 (N_19353,N_6576,N_2735);
xnor U19354 (N_19354,N_8055,N_8143);
nor U19355 (N_19355,N_457,N_489);
or U19356 (N_19356,N_2162,N_4564);
and U19357 (N_19357,N_6018,N_4041);
xor U19358 (N_19358,N_3328,N_6522);
nand U19359 (N_19359,N_6323,N_7442);
nand U19360 (N_19360,N_3081,N_4194);
or U19361 (N_19361,N_2033,N_4414);
nand U19362 (N_19362,N_567,N_3695);
or U19363 (N_19363,N_8879,N_6601);
xor U19364 (N_19364,N_2480,N_5594);
nor U19365 (N_19365,N_8889,N_8347);
and U19366 (N_19366,N_5295,N_5194);
nand U19367 (N_19367,N_2031,N_2279);
or U19368 (N_19368,N_9952,N_3919);
nor U19369 (N_19369,N_7052,N_4693);
nand U19370 (N_19370,N_3318,N_466);
and U19371 (N_19371,N_5092,N_2126);
or U19372 (N_19372,N_7524,N_8446);
nor U19373 (N_19373,N_1878,N_296);
xor U19374 (N_19374,N_9985,N_790);
and U19375 (N_19375,N_7147,N_3213);
or U19376 (N_19376,N_7034,N_4471);
or U19377 (N_19377,N_5863,N_4582);
or U19378 (N_19378,N_6411,N_4758);
or U19379 (N_19379,N_4895,N_5975);
nor U19380 (N_19380,N_9238,N_5697);
nor U19381 (N_19381,N_5158,N_5351);
nand U19382 (N_19382,N_3027,N_8816);
xnor U19383 (N_19383,N_6724,N_4595);
and U19384 (N_19384,N_7497,N_179);
and U19385 (N_19385,N_611,N_7711);
nand U19386 (N_19386,N_6143,N_1228);
nor U19387 (N_19387,N_3341,N_4883);
nor U19388 (N_19388,N_9063,N_998);
and U19389 (N_19389,N_1171,N_498);
nand U19390 (N_19390,N_1714,N_3516);
and U19391 (N_19391,N_967,N_8374);
nand U19392 (N_19392,N_8533,N_4451);
nand U19393 (N_19393,N_5761,N_4863);
nor U19394 (N_19394,N_5436,N_8099);
nand U19395 (N_19395,N_4876,N_755);
nand U19396 (N_19396,N_2407,N_7165);
xnor U19397 (N_19397,N_8128,N_3544);
and U19398 (N_19398,N_7108,N_5648);
nor U19399 (N_19399,N_5224,N_8477);
nand U19400 (N_19400,N_7015,N_450);
nor U19401 (N_19401,N_1791,N_7428);
nor U19402 (N_19402,N_4611,N_2194);
nor U19403 (N_19403,N_87,N_3542);
and U19404 (N_19404,N_1734,N_1119);
nand U19405 (N_19405,N_2850,N_6679);
nor U19406 (N_19406,N_7535,N_3332);
nand U19407 (N_19407,N_2940,N_6318);
nand U19408 (N_19408,N_8543,N_548);
or U19409 (N_19409,N_6293,N_1890);
and U19410 (N_19410,N_2476,N_4724);
or U19411 (N_19411,N_2391,N_9871);
and U19412 (N_19412,N_9263,N_7106);
or U19413 (N_19413,N_2094,N_9284);
or U19414 (N_19414,N_7228,N_9495);
nor U19415 (N_19415,N_8270,N_7689);
or U19416 (N_19416,N_9702,N_2946);
or U19417 (N_19417,N_7767,N_2482);
and U19418 (N_19418,N_1876,N_1189);
nor U19419 (N_19419,N_6112,N_6648);
nand U19420 (N_19420,N_7591,N_3795);
xor U19421 (N_19421,N_3615,N_9932);
nand U19422 (N_19422,N_4699,N_8353);
nor U19423 (N_19423,N_120,N_9009);
nand U19424 (N_19424,N_2355,N_7870);
or U19425 (N_19425,N_5165,N_2251);
or U19426 (N_19426,N_5718,N_28);
or U19427 (N_19427,N_9649,N_561);
nand U19428 (N_19428,N_4011,N_9023);
or U19429 (N_19429,N_8511,N_6894);
nor U19430 (N_19430,N_619,N_6190);
or U19431 (N_19431,N_9494,N_9322);
nor U19432 (N_19432,N_2230,N_9045);
nand U19433 (N_19433,N_912,N_2951);
nand U19434 (N_19434,N_480,N_3046);
xnor U19435 (N_19435,N_45,N_5219);
nor U19436 (N_19436,N_1474,N_7713);
and U19437 (N_19437,N_6426,N_7535);
nand U19438 (N_19438,N_6258,N_7463);
and U19439 (N_19439,N_7722,N_4533);
nand U19440 (N_19440,N_8725,N_6307);
nand U19441 (N_19441,N_6170,N_1999);
or U19442 (N_19442,N_8074,N_8222);
or U19443 (N_19443,N_8565,N_3026);
nand U19444 (N_19444,N_8725,N_1514);
or U19445 (N_19445,N_2328,N_3811);
and U19446 (N_19446,N_4073,N_283);
and U19447 (N_19447,N_6475,N_6401);
and U19448 (N_19448,N_8485,N_5960);
or U19449 (N_19449,N_152,N_3954);
or U19450 (N_19450,N_6879,N_7886);
xnor U19451 (N_19451,N_7140,N_4696);
or U19452 (N_19452,N_650,N_5832);
and U19453 (N_19453,N_9257,N_2651);
xnor U19454 (N_19454,N_5698,N_2749);
nand U19455 (N_19455,N_5302,N_9392);
nor U19456 (N_19456,N_8394,N_3334);
or U19457 (N_19457,N_2726,N_6451);
and U19458 (N_19458,N_4429,N_972);
nor U19459 (N_19459,N_435,N_1087);
or U19460 (N_19460,N_3877,N_2704);
xor U19461 (N_19461,N_2801,N_3427);
or U19462 (N_19462,N_8373,N_8962);
nand U19463 (N_19463,N_7071,N_8062);
nand U19464 (N_19464,N_6241,N_443);
nor U19465 (N_19465,N_9066,N_8261);
or U19466 (N_19466,N_1995,N_855);
nor U19467 (N_19467,N_8108,N_8014);
xnor U19468 (N_19468,N_6756,N_1974);
or U19469 (N_19469,N_4769,N_6612);
nor U19470 (N_19470,N_7389,N_3565);
and U19471 (N_19471,N_8190,N_2910);
or U19472 (N_19472,N_2119,N_6327);
nor U19473 (N_19473,N_109,N_8794);
nor U19474 (N_19474,N_9325,N_743);
nor U19475 (N_19475,N_7265,N_3987);
nor U19476 (N_19476,N_5020,N_7922);
or U19477 (N_19477,N_8393,N_8627);
nor U19478 (N_19478,N_7873,N_3399);
nor U19479 (N_19479,N_6684,N_1409);
and U19480 (N_19480,N_7977,N_4396);
and U19481 (N_19481,N_2886,N_1923);
or U19482 (N_19482,N_6929,N_9863);
nor U19483 (N_19483,N_5221,N_3554);
and U19484 (N_19484,N_9973,N_4317);
nand U19485 (N_19485,N_878,N_7190);
or U19486 (N_19486,N_7303,N_1962);
xnor U19487 (N_19487,N_1382,N_7136);
nand U19488 (N_19488,N_6421,N_9389);
nor U19489 (N_19489,N_1012,N_4194);
or U19490 (N_19490,N_685,N_9279);
and U19491 (N_19491,N_744,N_7842);
nand U19492 (N_19492,N_8742,N_5941);
nand U19493 (N_19493,N_4049,N_5094);
nand U19494 (N_19494,N_2030,N_8989);
nand U19495 (N_19495,N_6753,N_3357);
and U19496 (N_19496,N_4818,N_6724);
nand U19497 (N_19497,N_7138,N_461);
or U19498 (N_19498,N_7565,N_5854);
nor U19499 (N_19499,N_799,N_341);
nor U19500 (N_19500,N_2136,N_3280);
or U19501 (N_19501,N_1502,N_5036);
xor U19502 (N_19502,N_9440,N_1915);
and U19503 (N_19503,N_2274,N_5128);
nor U19504 (N_19504,N_2891,N_5030);
and U19505 (N_19505,N_4085,N_6558);
and U19506 (N_19506,N_555,N_8934);
nor U19507 (N_19507,N_4859,N_6921);
nor U19508 (N_19508,N_2201,N_944);
or U19509 (N_19509,N_7501,N_1109);
or U19510 (N_19510,N_2089,N_3609);
and U19511 (N_19511,N_8175,N_5955);
nand U19512 (N_19512,N_6596,N_5700);
nand U19513 (N_19513,N_305,N_9796);
and U19514 (N_19514,N_2835,N_4968);
nor U19515 (N_19515,N_9614,N_2862);
nand U19516 (N_19516,N_9395,N_8272);
or U19517 (N_19517,N_516,N_1307);
and U19518 (N_19518,N_8173,N_5660);
and U19519 (N_19519,N_7164,N_6262);
and U19520 (N_19520,N_8476,N_577);
nor U19521 (N_19521,N_5295,N_4838);
or U19522 (N_19522,N_9965,N_885);
and U19523 (N_19523,N_2868,N_7937);
xnor U19524 (N_19524,N_897,N_4733);
or U19525 (N_19525,N_1003,N_4682);
and U19526 (N_19526,N_2062,N_7529);
or U19527 (N_19527,N_4938,N_486);
nor U19528 (N_19528,N_7943,N_6303);
or U19529 (N_19529,N_4274,N_2166);
or U19530 (N_19530,N_2212,N_407);
nor U19531 (N_19531,N_591,N_4230);
and U19532 (N_19532,N_466,N_6864);
or U19533 (N_19533,N_9086,N_531);
nand U19534 (N_19534,N_885,N_9487);
and U19535 (N_19535,N_9863,N_5035);
xor U19536 (N_19536,N_2129,N_126);
and U19537 (N_19537,N_8139,N_7201);
and U19538 (N_19538,N_737,N_1712);
nand U19539 (N_19539,N_5653,N_1656);
and U19540 (N_19540,N_3078,N_3361);
and U19541 (N_19541,N_2325,N_702);
nor U19542 (N_19542,N_4576,N_9191);
nand U19543 (N_19543,N_1233,N_3187);
and U19544 (N_19544,N_4301,N_7782);
nor U19545 (N_19545,N_2831,N_5154);
nand U19546 (N_19546,N_2646,N_3018);
and U19547 (N_19547,N_5576,N_9367);
nor U19548 (N_19548,N_2220,N_7856);
nand U19549 (N_19549,N_7668,N_1793);
or U19550 (N_19550,N_9795,N_6734);
or U19551 (N_19551,N_9607,N_8598);
nor U19552 (N_19552,N_4217,N_2767);
nand U19553 (N_19553,N_5986,N_8552);
and U19554 (N_19554,N_2082,N_4767);
nor U19555 (N_19555,N_4616,N_823);
nor U19556 (N_19556,N_4502,N_2490);
or U19557 (N_19557,N_2785,N_7991);
or U19558 (N_19558,N_9308,N_6367);
and U19559 (N_19559,N_7792,N_939);
xnor U19560 (N_19560,N_6346,N_3619);
nor U19561 (N_19561,N_9178,N_911);
nor U19562 (N_19562,N_5630,N_9527);
or U19563 (N_19563,N_3312,N_5494);
or U19564 (N_19564,N_4327,N_6516);
or U19565 (N_19565,N_1441,N_6828);
or U19566 (N_19566,N_8147,N_4882);
or U19567 (N_19567,N_6044,N_6190);
and U19568 (N_19568,N_815,N_719);
xnor U19569 (N_19569,N_5005,N_4314);
xnor U19570 (N_19570,N_1259,N_4620);
or U19571 (N_19571,N_2477,N_8386);
nand U19572 (N_19572,N_6333,N_220);
nor U19573 (N_19573,N_6823,N_5058);
and U19574 (N_19574,N_8752,N_3904);
nand U19575 (N_19575,N_6181,N_9534);
nor U19576 (N_19576,N_1599,N_3115);
nor U19577 (N_19577,N_1727,N_387);
nor U19578 (N_19578,N_9538,N_4067);
nand U19579 (N_19579,N_5259,N_5747);
nor U19580 (N_19580,N_8251,N_7252);
nor U19581 (N_19581,N_2168,N_9977);
or U19582 (N_19582,N_9669,N_472);
nand U19583 (N_19583,N_4984,N_475);
nor U19584 (N_19584,N_3143,N_2404);
and U19585 (N_19585,N_9667,N_3706);
nor U19586 (N_19586,N_6627,N_5285);
xor U19587 (N_19587,N_3382,N_2900);
nor U19588 (N_19588,N_9740,N_8732);
nor U19589 (N_19589,N_7384,N_4987);
nand U19590 (N_19590,N_8703,N_6817);
nand U19591 (N_19591,N_6435,N_1511);
xor U19592 (N_19592,N_6504,N_1176);
nand U19593 (N_19593,N_9125,N_5101);
or U19594 (N_19594,N_2938,N_3431);
or U19595 (N_19595,N_7749,N_6811);
and U19596 (N_19596,N_6560,N_4427);
nand U19597 (N_19597,N_6201,N_2317);
or U19598 (N_19598,N_6552,N_6329);
nor U19599 (N_19599,N_1555,N_2443);
xnor U19600 (N_19600,N_4267,N_200);
and U19601 (N_19601,N_9430,N_291);
xnor U19602 (N_19602,N_711,N_5266);
nand U19603 (N_19603,N_8932,N_6290);
nand U19604 (N_19604,N_3452,N_3641);
and U19605 (N_19605,N_4772,N_6491);
nand U19606 (N_19606,N_3425,N_2664);
or U19607 (N_19607,N_6436,N_7931);
or U19608 (N_19608,N_9138,N_5536);
or U19609 (N_19609,N_7177,N_1678);
and U19610 (N_19610,N_6934,N_729);
nor U19611 (N_19611,N_7096,N_2750);
nor U19612 (N_19612,N_4282,N_2560);
nand U19613 (N_19613,N_5453,N_8417);
and U19614 (N_19614,N_3971,N_5603);
nand U19615 (N_19615,N_5083,N_7395);
xnor U19616 (N_19616,N_5301,N_3246);
nand U19617 (N_19617,N_6935,N_2459);
and U19618 (N_19618,N_9048,N_832);
xnor U19619 (N_19619,N_7686,N_3618);
and U19620 (N_19620,N_6589,N_8565);
and U19621 (N_19621,N_2074,N_1354);
xor U19622 (N_19622,N_6709,N_6874);
nand U19623 (N_19623,N_5252,N_8635);
nor U19624 (N_19624,N_4959,N_371);
nand U19625 (N_19625,N_2029,N_8033);
and U19626 (N_19626,N_7469,N_6268);
nand U19627 (N_19627,N_560,N_4908);
xor U19628 (N_19628,N_2538,N_7261);
and U19629 (N_19629,N_3716,N_5668);
nand U19630 (N_19630,N_122,N_9605);
or U19631 (N_19631,N_1156,N_598);
or U19632 (N_19632,N_7642,N_1497);
or U19633 (N_19633,N_6719,N_8105);
nand U19634 (N_19634,N_6001,N_3342);
or U19635 (N_19635,N_3080,N_8716);
nor U19636 (N_19636,N_7002,N_9452);
nand U19637 (N_19637,N_8743,N_3967);
nand U19638 (N_19638,N_7894,N_4039);
xor U19639 (N_19639,N_7479,N_658);
or U19640 (N_19640,N_2162,N_7243);
xor U19641 (N_19641,N_8097,N_3269);
nand U19642 (N_19642,N_3695,N_3335);
nand U19643 (N_19643,N_4987,N_8368);
or U19644 (N_19644,N_5042,N_4033);
and U19645 (N_19645,N_9536,N_5178);
and U19646 (N_19646,N_6111,N_6067);
nor U19647 (N_19647,N_5446,N_7672);
nor U19648 (N_19648,N_6000,N_3248);
xnor U19649 (N_19649,N_158,N_8125);
nand U19650 (N_19650,N_7711,N_99);
nand U19651 (N_19651,N_4679,N_1404);
xnor U19652 (N_19652,N_5610,N_6268);
and U19653 (N_19653,N_9405,N_5631);
nor U19654 (N_19654,N_9831,N_3931);
or U19655 (N_19655,N_3543,N_3394);
and U19656 (N_19656,N_8113,N_322);
and U19657 (N_19657,N_4684,N_3642);
or U19658 (N_19658,N_6012,N_7129);
or U19659 (N_19659,N_6919,N_5685);
nand U19660 (N_19660,N_6538,N_8612);
nand U19661 (N_19661,N_9508,N_5407);
xnor U19662 (N_19662,N_1514,N_8617);
nor U19663 (N_19663,N_3148,N_4047);
nor U19664 (N_19664,N_8468,N_7986);
and U19665 (N_19665,N_7917,N_442);
nand U19666 (N_19666,N_6927,N_8625);
and U19667 (N_19667,N_8194,N_5497);
nand U19668 (N_19668,N_7135,N_846);
nor U19669 (N_19669,N_4169,N_339);
or U19670 (N_19670,N_6349,N_6168);
xnor U19671 (N_19671,N_992,N_1933);
nand U19672 (N_19672,N_953,N_4);
nand U19673 (N_19673,N_546,N_5348);
xor U19674 (N_19674,N_2813,N_642);
nor U19675 (N_19675,N_492,N_6838);
nor U19676 (N_19676,N_2643,N_2324);
nor U19677 (N_19677,N_829,N_6907);
or U19678 (N_19678,N_5218,N_6433);
or U19679 (N_19679,N_525,N_4133);
and U19680 (N_19680,N_4571,N_6351);
nand U19681 (N_19681,N_5271,N_46);
or U19682 (N_19682,N_8150,N_3056);
nand U19683 (N_19683,N_5505,N_4341);
nand U19684 (N_19684,N_8621,N_1688);
nor U19685 (N_19685,N_3229,N_1099);
nor U19686 (N_19686,N_4711,N_4860);
and U19687 (N_19687,N_2528,N_6325);
nand U19688 (N_19688,N_1535,N_3753);
nand U19689 (N_19689,N_9929,N_9977);
nand U19690 (N_19690,N_8083,N_8102);
nand U19691 (N_19691,N_7214,N_7458);
nor U19692 (N_19692,N_4021,N_7593);
and U19693 (N_19693,N_2973,N_1119);
or U19694 (N_19694,N_2245,N_4137);
and U19695 (N_19695,N_2435,N_358);
nor U19696 (N_19696,N_5796,N_2788);
and U19697 (N_19697,N_6656,N_1342);
and U19698 (N_19698,N_3403,N_978);
or U19699 (N_19699,N_747,N_8759);
nor U19700 (N_19700,N_9551,N_9331);
or U19701 (N_19701,N_3960,N_1513);
nor U19702 (N_19702,N_2467,N_7724);
or U19703 (N_19703,N_574,N_617);
nand U19704 (N_19704,N_1030,N_6758);
nor U19705 (N_19705,N_1048,N_7546);
nor U19706 (N_19706,N_7231,N_2531);
or U19707 (N_19707,N_8502,N_9336);
nor U19708 (N_19708,N_6575,N_5956);
nand U19709 (N_19709,N_1381,N_3620);
nor U19710 (N_19710,N_6855,N_4158);
or U19711 (N_19711,N_7110,N_2598);
xnor U19712 (N_19712,N_9725,N_4375);
and U19713 (N_19713,N_1204,N_596);
and U19714 (N_19714,N_7644,N_3769);
or U19715 (N_19715,N_6370,N_3996);
nand U19716 (N_19716,N_5538,N_4901);
or U19717 (N_19717,N_1191,N_85);
nand U19718 (N_19718,N_254,N_8952);
nand U19719 (N_19719,N_2538,N_9919);
and U19720 (N_19720,N_7151,N_2925);
and U19721 (N_19721,N_172,N_2606);
nand U19722 (N_19722,N_7650,N_7478);
and U19723 (N_19723,N_9693,N_736);
or U19724 (N_19724,N_9511,N_1477);
and U19725 (N_19725,N_7213,N_9556);
nand U19726 (N_19726,N_1327,N_6214);
and U19727 (N_19727,N_1531,N_6119);
nand U19728 (N_19728,N_7948,N_5919);
nand U19729 (N_19729,N_6616,N_2312);
and U19730 (N_19730,N_3091,N_8908);
or U19731 (N_19731,N_7300,N_7474);
nor U19732 (N_19732,N_7355,N_7657);
nand U19733 (N_19733,N_5889,N_2901);
or U19734 (N_19734,N_8421,N_2166);
or U19735 (N_19735,N_169,N_3931);
and U19736 (N_19736,N_2003,N_9491);
nor U19737 (N_19737,N_1157,N_2933);
and U19738 (N_19738,N_9821,N_6233);
nor U19739 (N_19739,N_7970,N_7222);
nor U19740 (N_19740,N_5869,N_9885);
nor U19741 (N_19741,N_8326,N_1447);
or U19742 (N_19742,N_5746,N_2293);
and U19743 (N_19743,N_182,N_4472);
xor U19744 (N_19744,N_9496,N_2380);
nor U19745 (N_19745,N_2007,N_5584);
nor U19746 (N_19746,N_8812,N_9682);
and U19747 (N_19747,N_8414,N_9522);
nand U19748 (N_19748,N_6414,N_1391);
xnor U19749 (N_19749,N_475,N_2383);
xor U19750 (N_19750,N_9847,N_4086);
and U19751 (N_19751,N_7140,N_5172);
nand U19752 (N_19752,N_1486,N_723);
or U19753 (N_19753,N_4792,N_4607);
and U19754 (N_19754,N_7235,N_4671);
xnor U19755 (N_19755,N_9530,N_8542);
nor U19756 (N_19756,N_4064,N_8005);
nor U19757 (N_19757,N_4527,N_7599);
or U19758 (N_19758,N_6077,N_7331);
nor U19759 (N_19759,N_5892,N_2756);
nor U19760 (N_19760,N_3390,N_2309);
nor U19761 (N_19761,N_789,N_8464);
nand U19762 (N_19762,N_666,N_8338);
or U19763 (N_19763,N_9922,N_5326);
nand U19764 (N_19764,N_3292,N_2286);
and U19765 (N_19765,N_6283,N_2626);
nor U19766 (N_19766,N_8934,N_1499);
or U19767 (N_19767,N_9455,N_7584);
and U19768 (N_19768,N_3543,N_4120);
nand U19769 (N_19769,N_6035,N_6031);
nand U19770 (N_19770,N_5204,N_8906);
nor U19771 (N_19771,N_7870,N_5078);
and U19772 (N_19772,N_5458,N_9778);
nor U19773 (N_19773,N_4106,N_830);
nor U19774 (N_19774,N_6936,N_6569);
xor U19775 (N_19775,N_6235,N_6102);
nand U19776 (N_19776,N_7820,N_6490);
and U19777 (N_19777,N_8298,N_6973);
or U19778 (N_19778,N_5279,N_5222);
and U19779 (N_19779,N_2550,N_191);
or U19780 (N_19780,N_5216,N_473);
and U19781 (N_19781,N_9549,N_8740);
and U19782 (N_19782,N_624,N_783);
and U19783 (N_19783,N_9104,N_1686);
or U19784 (N_19784,N_2445,N_6119);
or U19785 (N_19785,N_4266,N_9619);
and U19786 (N_19786,N_6315,N_8634);
nand U19787 (N_19787,N_2327,N_1297);
nor U19788 (N_19788,N_5007,N_5995);
or U19789 (N_19789,N_5463,N_244);
and U19790 (N_19790,N_1459,N_7633);
xnor U19791 (N_19791,N_8470,N_5681);
or U19792 (N_19792,N_6116,N_1314);
nor U19793 (N_19793,N_3673,N_3154);
nor U19794 (N_19794,N_3070,N_732);
and U19795 (N_19795,N_4766,N_3083);
nor U19796 (N_19796,N_2257,N_7142);
and U19797 (N_19797,N_5269,N_450);
nand U19798 (N_19798,N_5962,N_5415);
xor U19799 (N_19799,N_8927,N_9524);
and U19800 (N_19800,N_1801,N_5633);
or U19801 (N_19801,N_3128,N_7346);
nand U19802 (N_19802,N_2913,N_4149);
and U19803 (N_19803,N_9323,N_9584);
or U19804 (N_19804,N_2368,N_5053);
nand U19805 (N_19805,N_803,N_1418);
nor U19806 (N_19806,N_4953,N_3063);
xnor U19807 (N_19807,N_5018,N_3407);
or U19808 (N_19808,N_4013,N_9554);
nand U19809 (N_19809,N_2243,N_3671);
nand U19810 (N_19810,N_761,N_2324);
nand U19811 (N_19811,N_8290,N_8992);
or U19812 (N_19812,N_8063,N_7561);
nor U19813 (N_19813,N_4478,N_7960);
nand U19814 (N_19814,N_5782,N_478);
nand U19815 (N_19815,N_6006,N_6602);
or U19816 (N_19816,N_4312,N_4035);
nor U19817 (N_19817,N_5935,N_9319);
nand U19818 (N_19818,N_4955,N_3188);
or U19819 (N_19819,N_9563,N_3191);
or U19820 (N_19820,N_4642,N_6173);
nor U19821 (N_19821,N_7665,N_8444);
or U19822 (N_19822,N_3819,N_183);
nor U19823 (N_19823,N_9202,N_5930);
and U19824 (N_19824,N_5491,N_6999);
nor U19825 (N_19825,N_7111,N_5861);
and U19826 (N_19826,N_813,N_3300);
or U19827 (N_19827,N_8672,N_4110);
nor U19828 (N_19828,N_732,N_9806);
nand U19829 (N_19829,N_8359,N_7408);
nand U19830 (N_19830,N_669,N_3460);
nand U19831 (N_19831,N_1621,N_801);
nand U19832 (N_19832,N_9859,N_5406);
and U19833 (N_19833,N_2248,N_680);
and U19834 (N_19834,N_5648,N_7643);
nor U19835 (N_19835,N_3507,N_1212);
or U19836 (N_19836,N_1567,N_2069);
and U19837 (N_19837,N_4386,N_3898);
nor U19838 (N_19838,N_8271,N_8612);
nor U19839 (N_19839,N_8848,N_4666);
nor U19840 (N_19840,N_1833,N_4649);
and U19841 (N_19841,N_2749,N_3052);
and U19842 (N_19842,N_7021,N_8324);
nand U19843 (N_19843,N_4511,N_1443);
nor U19844 (N_19844,N_4471,N_8159);
xnor U19845 (N_19845,N_8099,N_4209);
nand U19846 (N_19846,N_3644,N_5780);
and U19847 (N_19847,N_1661,N_1310);
nand U19848 (N_19848,N_6607,N_8029);
or U19849 (N_19849,N_2389,N_255);
or U19850 (N_19850,N_2775,N_9384);
nor U19851 (N_19851,N_2477,N_6477);
nor U19852 (N_19852,N_4065,N_1039);
or U19853 (N_19853,N_508,N_6661);
xor U19854 (N_19854,N_6986,N_5185);
nor U19855 (N_19855,N_5266,N_5035);
nand U19856 (N_19856,N_825,N_6712);
nor U19857 (N_19857,N_8557,N_2399);
and U19858 (N_19858,N_631,N_3991);
nor U19859 (N_19859,N_9294,N_1620);
nand U19860 (N_19860,N_5327,N_9700);
and U19861 (N_19861,N_7954,N_1673);
nor U19862 (N_19862,N_2013,N_7573);
nand U19863 (N_19863,N_5838,N_6496);
nor U19864 (N_19864,N_7085,N_8414);
or U19865 (N_19865,N_5815,N_1889);
nand U19866 (N_19866,N_751,N_1603);
and U19867 (N_19867,N_2742,N_4555);
nand U19868 (N_19868,N_6411,N_9967);
xor U19869 (N_19869,N_971,N_8563);
and U19870 (N_19870,N_694,N_9955);
nand U19871 (N_19871,N_8798,N_9554);
and U19872 (N_19872,N_4494,N_2594);
nor U19873 (N_19873,N_8400,N_8476);
or U19874 (N_19874,N_9480,N_4031);
and U19875 (N_19875,N_1719,N_7700);
or U19876 (N_19876,N_8370,N_2091);
nor U19877 (N_19877,N_9671,N_20);
and U19878 (N_19878,N_9276,N_9672);
nor U19879 (N_19879,N_3309,N_6740);
and U19880 (N_19880,N_5432,N_1840);
nor U19881 (N_19881,N_7242,N_9790);
nor U19882 (N_19882,N_1215,N_2992);
and U19883 (N_19883,N_9962,N_5263);
nor U19884 (N_19884,N_5836,N_6774);
nor U19885 (N_19885,N_9768,N_342);
nand U19886 (N_19886,N_1501,N_8400);
nor U19887 (N_19887,N_3091,N_6265);
nand U19888 (N_19888,N_7147,N_503);
or U19889 (N_19889,N_2440,N_7646);
and U19890 (N_19890,N_8949,N_9033);
or U19891 (N_19891,N_8050,N_8356);
or U19892 (N_19892,N_7853,N_7737);
nor U19893 (N_19893,N_6198,N_2339);
xor U19894 (N_19894,N_9873,N_3001);
nor U19895 (N_19895,N_3526,N_3790);
nor U19896 (N_19896,N_1440,N_7891);
nand U19897 (N_19897,N_3310,N_5755);
or U19898 (N_19898,N_4366,N_3789);
and U19899 (N_19899,N_2341,N_3264);
or U19900 (N_19900,N_1818,N_8039);
nor U19901 (N_19901,N_244,N_7053);
xnor U19902 (N_19902,N_6867,N_6422);
nand U19903 (N_19903,N_9023,N_6974);
xnor U19904 (N_19904,N_9270,N_1120);
and U19905 (N_19905,N_4451,N_3335);
or U19906 (N_19906,N_8946,N_4136);
nor U19907 (N_19907,N_2297,N_8797);
nand U19908 (N_19908,N_6121,N_3507);
or U19909 (N_19909,N_6789,N_1993);
nor U19910 (N_19910,N_9645,N_4191);
nand U19911 (N_19911,N_3877,N_9875);
nand U19912 (N_19912,N_3920,N_5504);
or U19913 (N_19913,N_8683,N_1305);
nand U19914 (N_19914,N_949,N_1880);
nor U19915 (N_19915,N_2277,N_5845);
or U19916 (N_19916,N_1911,N_5153);
nand U19917 (N_19917,N_7793,N_3768);
or U19918 (N_19918,N_1795,N_5997);
or U19919 (N_19919,N_5,N_4979);
nand U19920 (N_19920,N_6246,N_49);
and U19921 (N_19921,N_3848,N_4824);
and U19922 (N_19922,N_7533,N_7297);
and U19923 (N_19923,N_5123,N_8425);
nand U19924 (N_19924,N_2567,N_1350);
nand U19925 (N_19925,N_3618,N_5614);
xnor U19926 (N_19926,N_1898,N_2515);
nand U19927 (N_19927,N_2972,N_7110);
nor U19928 (N_19928,N_4462,N_1442);
or U19929 (N_19929,N_5866,N_9299);
nand U19930 (N_19930,N_9233,N_312);
nand U19931 (N_19931,N_5403,N_1955);
nand U19932 (N_19932,N_4815,N_4217);
and U19933 (N_19933,N_8534,N_7090);
and U19934 (N_19934,N_4275,N_1845);
nand U19935 (N_19935,N_8580,N_4175);
nand U19936 (N_19936,N_9602,N_1134);
or U19937 (N_19937,N_933,N_9423);
nor U19938 (N_19938,N_9579,N_5804);
and U19939 (N_19939,N_4230,N_2189);
or U19940 (N_19940,N_4779,N_7837);
or U19941 (N_19941,N_7545,N_7313);
and U19942 (N_19942,N_5506,N_7005);
nand U19943 (N_19943,N_8575,N_476);
xnor U19944 (N_19944,N_3491,N_3371);
or U19945 (N_19945,N_2124,N_533);
or U19946 (N_19946,N_5223,N_5232);
xor U19947 (N_19947,N_9459,N_7153);
nor U19948 (N_19948,N_1037,N_519);
or U19949 (N_19949,N_1814,N_4446);
nand U19950 (N_19950,N_3089,N_200);
or U19951 (N_19951,N_7004,N_2011);
and U19952 (N_19952,N_1995,N_4144);
and U19953 (N_19953,N_2872,N_6207);
nor U19954 (N_19954,N_8617,N_8315);
nand U19955 (N_19955,N_587,N_4048);
nand U19956 (N_19956,N_3030,N_2667);
and U19957 (N_19957,N_1531,N_5052);
nor U19958 (N_19958,N_4851,N_5326);
nor U19959 (N_19959,N_5252,N_5988);
or U19960 (N_19960,N_9436,N_4628);
or U19961 (N_19961,N_7676,N_8003);
nand U19962 (N_19962,N_3692,N_6800);
nand U19963 (N_19963,N_1147,N_7145);
and U19964 (N_19964,N_8029,N_2123);
nand U19965 (N_19965,N_7000,N_8107);
nand U19966 (N_19966,N_6386,N_9505);
or U19967 (N_19967,N_44,N_5466);
nor U19968 (N_19968,N_2283,N_1466);
xor U19969 (N_19969,N_6502,N_4745);
and U19970 (N_19970,N_6163,N_1321);
or U19971 (N_19971,N_4385,N_6299);
or U19972 (N_19972,N_6881,N_4690);
nor U19973 (N_19973,N_2183,N_8275);
xor U19974 (N_19974,N_2147,N_1106);
xor U19975 (N_19975,N_7802,N_9687);
xnor U19976 (N_19976,N_1672,N_7228);
or U19977 (N_19977,N_7376,N_350);
or U19978 (N_19978,N_40,N_7105);
and U19979 (N_19979,N_212,N_3011);
xor U19980 (N_19980,N_2849,N_4491);
nand U19981 (N_19981,N_4790,N_506);
and U19982 (N_19982,N_7772,N_6998);
or U19983 (N_19983,N_1929,N_3267);
nand U19984 (N_19984,N_6798,N_5894);
and U19985 (N_19985,N_8980,N_2726);
and U19986 (N_19986,N_4767,N_557);
nand U19987 (N_19987,N_9944,N_1119);
or U19988 (N_19988,N_7173,N_1470);
and U19989 (N_19989,N_5135,N_5943);
nand U19990 (N_19990,N_8178,N_9146);
or U19991 (N_19991,N_8694,N_7597);
nor U19992 (N_19992,N_1754,N_5107);
nor U19993 (N_19993,N_3662,N_5417);
or U19994 (N_19994,N_3519,N_7719);
nor U19995 (N_19995,N_3102,N_6220);
and U19996 (N_19996,N_8989,N_8438);
or U19997 (N_19997,N_1733,N_3389);
nand U19998 (N_19998,N_1830,N_922);
or U19999 (N_19999,N_4041,N_6862);
and U20000 (N_20000,N_17270,N_10535);
xnor U20001 (N_20001,N_13006,N_16573);
or U20002 (N_20002,N_19548,N_19204);
nor U20003 (N_20003,N_14320,N_12231);
or U20004 (N_20004,N_15560,N_17957);
and U20005 (N_20005,N_11470,N_11937);
and U20006 (N_20006,N_10259,N_13255);
and U20007 (N_20007,N_14960,N_19950);
xnor U20008 (N_20008,N_13955,N_15771);
nand U20009 (N_20009,N_10609,N_10919);
and U20010 (N_20010,N_12644,N_11133);
and U20011 (N_20011,N_10487,N_15868);
nand U20012 (N_20012,N_11434,N_15787);
and U20013 (N_20013,N_12692,N_12397);
nand U20014 (N_20014,N_12713,N_13726);
and U20015 (N_20015,N_19186,N_16632);
nand U20016 (N_20016,N_15334,N_15869);
or U20017 (N_20017,N_12089,N_15275);
nand U20018 (N_20018,N_13404,N_14902);
xnor U20019 (N_20019,N_17639,N_12969);
nand U20020 (N_20020,N_18921,N_19367);
nand U20021 (N_20021,N_17812,N_17493);
nor U20022 (N_20022,N_19954,N_12457);
xor U20023 (N_20023,N_13502,N_16120);
nor U20024 (N_20024,N_17326,N_14394);
and U20025 (N_20025,N_14113,N_14488);
nand U20026 (N_20026,N_12765,N_11376);
and U20027 (N_20027,N_12774,N_14035);
nor U20028 (N_20028,N_14012,N_19257);
or U20029 (N_20029,N_13801,N_12389);
nand U20030 (N_20030,N_16646,N_18665);
nand U20031 (N_20031,N_18409,N_16637);
nand U20032 (N_20032,N_19565,N_19205);
nand U20033 (N_20033,N_14596,N_13062);
nand U20034 (N_20034,N_16558,N_17168);
nand U20035 (N_20035,N_15059,N_10087);
and U20036 (N_20036,N_14690,N_17414);
or U20037 (N_20037,N_13492,N_17693);
and U20038 (N_20038,N_18649,N_11509);
or U20039 (N_20039,N_17701,N_18795);
and U20040 (N_20040,N_15429,N_19721);
xnor U20041 (N_20041,N_17296,N_16955);
or U20042 (N_20042,N_15746,N_13626);
or U20043 (N_20043,N_11419,N_13760);
nor U20044 (N_20044,N_16500,N_17409);
nor U20045 (N_20045,N_17246,N_10616);
nand U20046 (N_20046,N_17987,N_10938);
nand U20047 (N_20047,N_12268,N_19052);
and U20048 (N_20048,N_19789,N_18619);
xor U20049 (N_20049,N_14407,N_16576);
or U20050 (N_20050,N_18899,N_12134);
nand U20051 (N_20051,N_17034,N_13116);
nor U20052 (N_20052,N_14661,N_12186);
or U20053 (N_20053,N_12886,N_16694);
xnor U20054 (N_20054,N_12218,N_14993);
or U20055 (N_20055,N_13157,N_16687);
nor U20056 (N_20056,N_13769,N_16454);
nor U20057 (N_20057,N_10170,N_12794);
and U20058 (N_20058,N_16855,N_15605);
nand U20059 (N_20059,N_13276,N_10733);
and U20060 (N_20060,N_13306,N_11207);
xor U20061 (N_20061,N_19199,N_12893);
or U20062 (N_20062,N_13004,N_17882);
and U20063 (N_20063,N_17210,N_12876);
nor U20064 (N_20064,N_13470,N_15321);
or U20065 (N_20065,N_15026,N_10104);
xor U20066 (N_20066,N_14353,N_15543);
and U20067 (N_20067,N_13387,N_13831);
nand U20068 (N_20068,N_16691,N_15510);
nor U20069 (N_20069,N_19917,N_18135);
or U20070 (N_20070,N_15646,N_13482);
nor U20071 (N_20071,N_13007,N_10627);
nand U20072 (N_20072,N_18971,N_16131);
or U20073 (N_20073,N_15182,N_14380);
or U20074 (N_20074,N_14793,N_17138);
xnor U20075 (N_20075,N_19349,N_13922);
nor U20076 (N_20076,N_12639,N_19222);
or U20077 (N_20077,N_16307,N_12852);
xor U20078 (N_20078,N_12091,N_14972);
xor U20079 (N_20079,N_16693,N_15558);
and U20080 (N_20080,N_16752,N_16996);
and U20081 (N_20081,N_12427,N_12467);
and U20082 (N_20082,N_11766,N_13466);
or U20083 (N_20083,N_15502,N_17725);
nand U20084 (N_20084,N_12031,N_12707);
nand U20085 (N_20085,N_10156,N_16856);
or U20086 (N_20086,N_12778,N_15181);
or U20087 (N_20087,N_11687,N_13258);
or U20088 (N_20088,N_19755,N_14391);
nor U20089 (N_20089,N_11850,N_17068);
or U20090 (N_20090,N_18656,N_18141);
or U20091 (N_20091,N_14147,N_17405);
nor U20092 (N_20092,N_17368,N_18629);
nand U20093 (N_20093,N_13183,N_13485);
nand U20094 (N_20094,N_19028,N_11107);
nand U20095 (N_20095,N_16795,N_18192);
nand U20096 (N_20096,N_12292,N_17392);
nand U20097 (N_20097,N_13612,N_14221);
and U20098 (N_20098,N_16053,N_14425);
or U20099 (N_20099,N_17627,N_17247);
nor U20100 (N_20100,N_11635,N_18461);
nand U20101 (N_20101,N_18071,N_10353);
and U20102 (N_20102,N_17915,N_19497);
and U20103 (N_20103,N_14317,N_10710);
or U20104 (N_20104,N_16496,N_10331);
or U20105 (N_20105,N_17080,N_16132);
nor U20106 (N_20106,N_14710,N_14582);
or U20107 (N_20107,N_14479,N_17266);
nand U20108 (N_20108,N_13580,N_17006);
nor U20109 (N_20109,N_18621,N_13483);
and U20110 (N_20110,N_13223,N_17182);
nor U20111 (N_20111,N_11867,N_19491);
nor U20112 (N_20112,N_10597,N_19360);
and U20113 (N_20113,N_12949,N_16703);
nand U20114 (N_20114,N_14719,N_13884);
and U20115 (N_20115,N_16945,N_19729);
nor U20116 (N_20116,N_17402,N_14512);
nand U20117 (N_20117,N_16524,N_15107);
and U20118 (N_20118,N_17188,N_10185);
nand U20119 (N_20119,N_12073,N_11785);
nand U20120 (N_20120,N_14509,N_17863);
nor U20121 (N_20121,N_16139,N_12050);
or U20122 (N_20122,N_19692,N_18824);
nand U20123 (N_20123,N_18917,N_15263);
nor U20124 (N_20124,N_15127,N_18394);
nand U20125 (N_20125,N_13731,N_10501);
nand U20126 (N_20126,N_15405,N_12108);
nor U20127 (N_20127,N_16381,N_12258);
or U20128 (N_20128,N_10498,N_12354);
and U20129 (N_20129,N_11809,N_13239);
and U20130 (N_20130,N_14003,N_17346);
nand U20131 (N_20131,N_11771,N_17791);
or U20132 (N_20132,N_18988,N_12747);
and U20133 (N_20133,N_18561,N_14025);
and U20134 (N_20134,N_17901,N_19981);
or U20135 (N_20135,N_19424,N_19730);
nand U20136 (N_20136,N_13591,N_18252);
and U20137 (N_20137,N_16372,N_15239);
and U20138 (N_20138,N_16651,N_13304);
or U20139 (N_20139,N_16584,N_11847);
and U20140 (N_20140,N_14751,N_12016);
or U20141 (N_20141,N_13989,N_15986);
nor U20142 (N_20142,N_16827,N_10187);
or U20143 (N_20143,N_10297,N_16543);
or U20144 (N_20144,N_10916,N_15707);
nor U20145 (N_20145,N_10626,N_10666);
and U20146 (N_20146,N_15449,N_11001);
xnor U20147 (N_20147,N_14297,N_16376);
nand U20148 (N_20148,N_19943,N_18378);
nor U20149 (N_20149,N_16509,N_14144);
nor U20150 (N_20150,N_11853,N_14953);
nand U20151 (N_20151,N_17698,N_18504);
nand U20152 (N_20152,N_15630,N_18827);
xnor U20153 (N_20153,N_17554,N_16879);
nand U20154 (N_20154,N_15472,N_17448);
nand U20155 (N_20155,N_14838,N_17197);
nand U20156 (N_20156,N_17353,N_10067);
nand U20157 (N_20157,N_12514,N_16602);
nor U20158 (N_20158,N_19207,N_12421);
nand U20159 (N_20159,N_10912,N_18983);
and U20160 (N_20160,N_18502,N_10814);
and U20161 (N_20161,N_12320,N_10399);
or U20162 (N_20162,N_19370,N_14129);
or U20163 (N_20163,N_19811,N_15092);
nand U20164 (N_20164,N_18466,N_12360);
nand U20165 (N_20165,N_12978,N_16830);
nor U20166 (N_20166,N_15160,N_13904);
or U20167 (N_20167,N_14554,N_10869);
or U20168 (N_20168,N_16325,N_16130);
nand U20169 (N_20169,N_15208,N_19608);
xor U20170 (N_20170,N_12349,N_13853);
and U20171 (N_20171,N_16750,N_10580);
nor U20172 (N_20172,N_17002,N_19812);
nor U20173 (N_20173,N_12128,N_18133);
nand U20174 (N_20174,N_18435,N_17831);
xor U20175 (N_20175,N_12741,N_11415);
or U20176 (N_20176,N_16142,N_17676);
nor U20177 (N_20177,N_19393,N_10727);
nand U20178 (N_20178,N_19131,N_18352);
nand U20179 (N_20179,N_12845,N_17672);
xnor U20180 (N_20180,N_10781,N_15491);
nor U20181 (N_20181,N_16464,N_14911);
and U20182 (N_20182,N_19467,N_10782);
nand U20183 (N_20183,N_11544,N_11138);
and U20184 (N_20184,N_17503,N_17768);
nor U20185 (N_20185,N_14056,N_19470);
nand U20186 (N_20186,N_16705,N_15667);
nor U20187 (N_20187,N_16812,N_15083);
nor U20188 (N_20188,N_19797,N_10208);
nand U20189 (N_20189,N_17680,N_11061);
nor U20190 (N_20190,N_13189,N_11627);
nand U20191 (N_20191,N_19447,N_14529);
and U20192 (N_20192,N_17261,N_14522);
nand U20193 (N_20193,N_12358,N_17692);
nand U20194 (N_20194,N_15523,N_13906);
or U20195 (N_20195,N_11350,N_10771);
nand U20196 (N_20196,N_13866,N_12938);
nor U20197 (N_20197,N_17171,N_12951);
nand U20198 (N_20198,N_12720,N_11045);
or U20199 (N_20199,N_18398,N_14173);
xor U20200 (N_20200,N_11671,N_12677);
and U20201 (N_20201,N_17185,N_18861);
nor U20202 (N_20202,N_18332,N_13133);
nor U20203 (N_20203,N_12924,N_18677);
nor U20204 (N_20204,N_15933,N_18322);
nand U20205 (N_20205,N_11799,N_15873);
nor U20206 (N_20206,N_14603,N_18553);
nor U20207 (N_20207,N_13272,N_14285);
nor U20208 (N_20208,N_12615,N_17723);
xnor U20209 (N_20209,N_17015,N_13015);
nor U20210 (N_20210,N_19206,N_15290);
nor U20211 (N_20211,N_14322,N_15637);
and U20212 (N_20212,N_17875,N_15411);
nor U20213 (N_20213,N_12155,N_15671);
nand U20214 (N_20214,N_14002,N_15685);
and U20215 (N_20215,N_18754,N_10473);
and U20216 (N_20216,N_15328,N_19637);
nor U20217 (N_20217,N_11842,N_14271);
nand U20218 (N_20218,N_18505,N_12718);
nor U20219 (N_20219,N_15017,N_19466);
xnor U20220 (N_20220,N_17218,N_10550);
and U20221 (N_20221,N_15512,N_14106);
nor U20222 (N_20222,N_11127,N_14517);
or U20223 (N_20223,N_15769,N_11583);
nand U20224 (N_20224,N_17881,N_10116);
nand U20225 (N_20225,N_10920,N_11199);
or U20226 (N_20226,N_16732,N_14920);
nand U20227 (N_20227,N_17076,N_18701);
nor U20228 (N_20228,N_10345,N_12275);
nand U20229 (N_20229,N_13102,N_19213);
nand U20230 (N_20230,N_18651,N_18779);
and U20231 (N_20231,N_19615,N_10101);
nor U20232 (N_20232,N_16551,N_12167);
or U20233 (N_20233,N_14471,N_12995);
nor U20234 (N_20234,N_18512,N_10654);
nand U20235 (N_20235,N_14216,N_16063);
and U20236 (N_20236,N_15498,N_15675);
xnor U20237 (N_20237,N_16066,N_18529);
and U20238 (N_20238,N_13799,N_14747);
and U20239 (N_20239,N_12971,N_11593);
nand U20240 (N_20240,N_19579,N_14762);
and U20241 (N_20241,N_13548,N_19119);
or U20242 (N_20242,N_15420,N_14931);
or U20243 (N_20243,N_11776,N_11651);
or U20244 (N_20244,N_19104,N_19862);
nor U20245 (N_20245,N_13518,N_16967);
nor U20246 (N_20246,N_19455,N_13281);
and U20247 (N_20247,N_13105,N_19378);
or U20248 (N_20248,N_11320,N_12248);
and U20249 (N_20249,N_19779,N_10184);
or U20250 (N_20250,N_11324,N_10567);
xnor U20251 (N_20251,N_13733,N_14359);
nand U20252 (N_20252,N_14589,N_11835);
nand U20253 (N_20253,N_12868,N_13581);
and U20254 (N_20254,N_19149,N_12664);
nand U20255 (N_20255,N_17230,N_16483);
or U20256 (N_20256,N_10930,N_14867);
nand U20257 (N_20257,N_15978,N_10466);
nand U20258 (N_20258,N_15979,N_11598);
and U20259 (N_20259,N_18851,N_17564);
and U20260 (N_20260,N_18932,N_18823);
nand U20261 (N_20261,N_16156,N_18054);
and U20262 (N_20262,N_10739,N_19567);
and U20263 (N_20263,N_10203,N_11726);
xnor U20264 (N_20264,N_12244,N_19271);
and U20265 (N_20265,N_17484,N_16636);
or U20266 (N_20266,N_14375,N_15976);
and U20267 (N_20267,N_11128,N_19815);
nand U20268 (N_20268,N_16530,N_18216);
or U20269 (N_20269,N_10443,N_19158);
nor U20270 (N_20270,N_12979,N_11910);
xor U20271 (N_20271,N_14796,N_14694);
or U20272 (N_20272,N_11570,N_12694);
nand U20273 (N_20273,N_19536,N_14184);
and U20274 (N_20274,N_14503,N_12007);
nor U20275 (N_20275,N_17844,N_15090);
and U20276 (N_20276,N_13727,N_17505);
xnor U20277 (N_20277,N_13386,N_14677);
nor U20278 (N_20278,N_16112,N_10014);
and U20279 (N_20279,N_10846,N_16616);
and U20280 (N_20280,N_14215,N_11304);
nand U20281 (N_20281,N_13136,N_14905);
and U20282 (N_20282,N_11861,N_11969);
and U20283 (N_20283,N_14430,N_15853);
and U20284 (N_20284,N_14121,N_19887);
nor U20285 (N_20285,N_14089,N_13093);
nor U20286 (N_20286,N_12039,N_18246);
or U20287 (N_20287,N_10629,N_16428);
and U20288 (N_20288,N_12630,N_18140);
and U20289 (N_20289,N_14846,N_14812);
and U20290 (N_20290,N_18060,N_15117);
nor U20291 (N_20291,N_17551,N_12879);
and U20292 (N_20292,N_17852,N_16587);
nand U20293 (N_20293,N_13011,N_11984);
nor U20294 (N_20294,N_17119,N_12026);
or U20295 (N_20295,N_14681,N_19550);
or U20296 (N_20296,N_17956,N_16012);
and U20297 (N_20297,N_15442,N_11574);
and U20298 (N_20298,N_15206,N_19046);
nand U20299 (N_20299,N_10157,N_16900);
or U20300 (N_20300,N_19510,N_13441);
nand U20301 (N_20301,N_19184,N_19949);
and U20302 (N_20302,N_14961,N_18969);
xnor U20303 (N_20303,N_19234,N_15705);
nor U20304 (N_20304,N_10385,N_13729);
and U20305 (N_20305,N_18439,N_16233);
or U20306 (N_20306,N_17038,N_11442);
nand U20307 (N_20307,N_12503,N_16612);
and U20308 (N_20308,N_17673,N_15219);
nor U20309 (N_20309,N_10624,N_18552);
or U20310 (N_20310,N_10973,N_13583);
or U20311 (N_20311,N_18263,N_18535);
xnor U20312 (N_20312,N_13089,N_18238);
nor U20313 (N_20313,N_14605,N_18325);
nor U20314 (N_20314,N_18503,N_13090);
nand U20315 (N_20315,N_10420,N_19521);
nor U20316 (N_20316,N_14732,N_19761);
nor U20317 (N_20317,N_19896,N_10432);
nand U20318 (N_20318,N_13233,N_16221);
or U20319 (N_20319,N_17345,N_19471);
nand U20320 (N_20320,N_13422,N_13500);
or U20321 (N_20321,N_14679,N_17947);
nand U20322 (N_20322,N_13000,N_14564);
or U20323 (N_20323,N_13888,N_15551);
and U20324 (N_20324,N_19636,N_12806);
or U20325 (N_20325,N_11961,N_13859);
and U20326 (N_20326,N_10484,N_18302);
and U20327 (N_20327,N_11351,N_12369);
and U20328 (N_20328,N_14822,N_13926);
nor U20329 (N_20329,N_17737,N_13900);
and U20330 (N_20330,N_14767,N_19894);
xnor U20331 (N_20331,N_15141,N_17308);
or U20332 (N_20332,N_15254,N_13746);
nand U20333 (N_20333,N_14177,N_10133);
nand U20334 (N_20334,N_10741,N_10428);
and U20335 (N_20335,N_13380,N_18058);
and U20336 (N_20336,N_17443,N_17634);
nor U20337 (N_20337,N_19354,N_16627);
nand U20338 (N_20338,N_16475,N_19633);
nand U20339 (N_20339,N_13508,N_13653);
nor U20340 (N_20340,N_10859,N_19531);
or U20341 (N_20341,N_17647,N_18806);
nand U20342 (N_20342,N_13098,N_11747);
nand U20343 (N_20343,N_10748,N_12609);
nand U20344 (N_20344,N_15082,N_17380);
and U20345 (N_20345,N_12093,N_16242);
nor U20346 (N_20346,N_18579,N_10034);
nand U20347 (N_20347,N_14361,N_14636);
nand U20348 (N_20348,N_10499,N_11550);
or U20349 (N_20349,N_17435,N_10472);
nor U20350 (N_20350,N_11988,N_17733);
nor U20351 (N_20351,N_16238,N_12245);
xnor U20352 (N_20352,N_17646,N_18608);
and U20353 (N_20353,N_16251,N_11801);
and U20354 (N_20354,N_13827,N_12149);
nor U20355 (N_20355,N_12575,N_10437);
and U20356 (N_20356,N_10056,N_16976);
and U20357 (N_20357,N_18496,N_13851);
nor U20358 (N_20358,N_15526,N_15474);
and U20359 (N_20359,N_17532,N_16745);
and U20360 (N_20360,N_18515,N_16357);
and U20361 (N_20361,N_19082,N_11689);
nand U20362 (N_20362,N_13046,N_14206);
nand U20363 (N_20363,N_19100,N_12424);
or U20364 (N_20364,N_12836,N_10984);
and U20365 (N_20365,N_16973,N_18180);
nor U20366 (N_20366,N_10915,N_10253);
and U20367 (N_20367,N_12184,N_19547);
nand U20368 (N_20368,N_16441,N_12351);
nand U20369 (N_20369,N_13114,N_10848);
and U20370 (N_20370,N_11158,N_15844);
nand U20371 (N_20371,N_13975,N_18097);
nand U20372 (N_20372,N_18412,N_19033);
and U20373 (N_20373,N_15692,N_10078);
and U20374 (N_20374,N_19012,N_18888);
nor U20375 (N_20375,N_11298,N_18789);
or U20376 (N_20376,N_11954,N_15482);
xnor U20377 (N_20377,N_12085,N_18421);
nor U20378 (N_20378,N_15199,N_15106);
and U20379 (N_20379,N_11178,N_10564);
and U20380 (N_20380,N_19589,N_16974);
and U20381 (N_20381,N_12107,N_12635);
xor U20382 (N_20382,N_19495,N_11393);
nand U20383 (N_20383,N_13848,N_14853);
and U20384 (N_20384,N_11716,N_19468);
or U20385 (N_20385,N_14921,N_16890);
xor U20386 (N_20386,N_18032,N_17041);
and U20387 (N_20387,N_16948,N_16726);
nand U20388 (N_20388,N_17565,N_17284);
or U20389 (N_20389,N_15195,N_12197);
and U20390 (N_20390,N_18819,N_14898);
xor U20391 (N_20391,N_13571,N_14585);
xor U20392 (N_20392,N_14854,N_19445);
nand U20393 (N_20393,N_18499,N_15387);
nand U20394 (N_20394,N_17450,N_17026);
or U20395 (N_20395,N_11560,N_13228);
and U20396 (N_20396,N_17487,N_11422);
nand U20397 (N_20397,N_14658,N_18541);
or U20398 (N_20398,N_18782,N_18012);
nand U20399 (N_20399,N_16677,N_15170);
nand U20400 (N_20400,N_12823,N_12614);
nor U20401 (N_20401,N_19923,N_15694);
and U20402 (N_20402,N_15786,N_18778);
or U20403 (N_20403,N_19386,N_18755);
and U20404 (N_20404,N_19725,N_14883);
nor U20405 (N_20405,N_12054,N_18893);
nor U20406 (N_20406,N_10444,N_14524);
nor U20407 (N_20407,N_15114,N_17625);
nand U20408 (N_20408,N_11763,N_11959);
or U20409 (N_20409,N_13495,N_16596);
or U20410 (N_20410,N_11077,N_10937);
xor U20411 (N_20411,N_18614,N_16350);
and U20412 (N_20412,N_14871,N_10887);
nor U20413 (N_20413,N_15492,N_10663);
nand U20414 (N_20414,N_10182,N_17282);
nor U20415 (N_20415,N_14030,N_18189);
or U20416 (N_20416,N_14332,N_10097);
and U20417 (N_20417,N_18057,N_10296);
and U20418 (N_20418,N_10488,N_10482);
nor U20419 (N_20419,N_13073,N_13957);
and U20420 (N_20420,N_16158,N_17475);
and U20421 (N_20421,N_16570,N_12544);
nor U20422 (N_20422,N_15884,N_13174);
or U20423 (N_20423,N_19118,N_11056);
nor U20424 (N_20424,N_13311,N_15426);
or U20425 (N_20425,N_18127,N_11235);
nor U20426 (N_20426,N_17681,N_17050);
or U20427 (N_20427,N_19898,N_17577);
nand U20428 (N_20428,N_11846,N_11586);
or U20429 (N_20429,N_13165,N_17980);
xor U20430 (N_20430,N_13303,N_16582);
xor U20431 (N_20431,N_10284,N_10803);
or U20432 (N_20432,N_15467,N_18316);
and U20433 (N_20433,N_10142,N_14486);
or U20434 (N_20434,N_10953,N_11386);
and U20435 (N_20435,N_12885,N_18815);
xor U20436 (N_20436,N_16457,N_13976);
nand U20437 (N_20437,N_13080,N_18210);
or U20438 (N_20438,N_17787,N_12873);
and U20439 (N_20439,N_18202,N_13118);
nor U20440 (N_20440,N_18069,N_18284);
nand U20441 (N_20441,N_14559,N_14368);
nand U20442 (N_20442,N_18123,N_10502);
or U20443 (N_20443,N_18793,N_15923);
or U20444 (N_20444,N_10998,N_19243);
nand U20445 (N_20445,N_12533,N_13456);
or U20446 (N_20446,N_18879,N_16824);
and U20447 (N_20447,N_14253,N_12185);
and U20448 (N_20448,N_18718,N_15522);
or U20449 (N_20449,N_16215,N_15257);
and U20450 (N_20450,N_19128,N_13014);
nor U20451 (N_20451,N_11622,N_18315);
or U20452 (N_20452,N_19317,N_19478);
and U20453 (N_20453,N_17399,N_13864);
and U20454 (N_20454,N_19630,N_16067);
xor U20455 (N_20455,N_12444,N_10907);
and U20456 (N_20456,N_18338,N_11302);
nor U20457 (N_20457,N_19599,N_10398);
nand U20458 (N_20458,N_17338,N_19150);
xor U20459 (N_20459,N_19942,N_15759);
xnor U20460 (N_20460,N_13211,N_18685);
or U20461 (N_20461,N_15528,N_17113);
or U20462 (N_20462,N_13562,N_18237);
nor U20463 (N_20463,N_17310,N_16924);
or U20464 (N_20464,N_14408,N_13787);
nor U20465 (N_20465,N_16971,N_13603);
nor U20466 (N_20466,N_13496,N_11339);
xor U20467 (N_20467,N_18543,N_16147);
and U20468 (N_20468,N_15155,N_11182);
nor U20469 (N_20469,N_16828,N_15470);
or U20470 (N_20470,N_14260,N_18478);
nor U20471 (N_20471,N_14474,N_18389);
and U20472 (N_20472,N_13546,N_14499);
or U20473 (N_20473,N_17880,N_12018);
nand U20474 (N_20474,N_14434,N_18273);
and U20475 (N_20475,N_15299,N_14688);
or U20476 (N_20476,N_16462,N_15863);
or U20477 (N_20477,N_12835,N_13987);
nor U20478 (N_20478,N_17196,N_19764);
and U20479 (N_20479,N_14096,N_17229);
or U20480 (N_20480,N_16127,N_16774);
or U20481 (N_20481,N_12669,N_11945);
nand U20482 (N_20482,N_16575,N_17952);
and U20483 (N_20483,N_11909,N_14876);
and U20484 (N_20484,N_17615,N_12584);
nor U20485 (N_20485,N_13151,N_14240);
nor U20486 (N_20486,N_14996,N_12223);
nor U20487 (N_20487,N_11623,N_12997);
nand U20488 (N_20488,N_18716,N_16787);
nand U20489 (N_20489,N_16079,N_10225);
nand U20490 (N_20490,N_17144,N_12772);
or U20491 (N_20491,N_12912,N_19098);
nor U20492 (N_20492,N_17355,N_19530);
and U20493 (N_20493,N_12483,N_16170);
xor U20494 (N_20494,N_17391,N_11002);
nor U20495 (N_20495,N_18171,N_10053);
nor U20496 (N_20496,N_18021,N_12058);
or U20497 (N_20497,N_18312,N_11624);
nor U20498 (N_20498,N_12527,N_11818);
nor U20499 (N_20499,N_11484,N_14712);
and U20500 (N_20500,N_16721,N_16057);
and U20501 (N_20501,N_17430,N_11461);
nor U20502 (N_20502,N_19888,N_15267);
nand U20503 (N_20503,N_12222,N_18562);
and U20504 (N_20504,N_14709,N_13036);
nand U20505 (N_20505,N_18230,N_16392);
or U20506 (N_20506,N_11337,N_10659);
and U20507 (N_20507,N_19622,N_16807);
nand U20508 (N_20508,N_19808,N_10596);
and U20509 (N_20509,N_14182,N_19605);
or U20510 (N_20510,N_14141,N_15274);
and U20511 (N_20511,N_14477,N_12083);
nor U20512 (N_20512,N_19836,N_15910);
or U20513 (N_20513,N_15806,N_12974);
or U20514 (N_20514,N_12629,N_19787);
xnor U20515 (N_20515,N_19237,N_10177);
nor U20516 (N_20516,N_10683,N_16114);
nor U20517 (N_20517,N_16507,N_11232);
nor U20518 (N_20518,N_13213,N_14954);
and U20519 (N_20519,N_12468,N_11340);
or U20520 (N_20520,N_14084,N_10205);
and U20521 (N_20521,N_14922,N_13516);
nand U20522 (N_20522,N_14252,N_18558);
nor U20523 (N_20523,N_15917,N_17526);
or U20524 (N_20524,N_15653,N_14689);
nand U20525 (N_20525,N_16135,N_14330);
and U20526 (N_20526,N_16652,N_19810);
nor U20527 (N_20527,N_19733,N_11252);
nor U20528 (N_20528,N_12964,N_17317);
nand U20529 (N_20529,N_15345,N_10464);
nor U20530 (N_20530,N_17258,N_17059);
nand U20531 (N_20531,N_19160,N_11829);
nor U20532 (N_20532,N_16369,N_12840);
nor U20533 (N_20533,N_19773,N_15276);
nand U20534 (N_20534,N_10414,N_11514);
or U20535 (N_20535,N_17764,N_18872);
and U20536 (N_20536,N_18700,N_16660);
nor U20537 (N_20537,N_13682,N_17242);
xor U20538 (N_20538,N_17751,N_18086);
and U20539 (N_20539,N_17250,N_12751);
or U20540 (N_20540,N_11911,N_15376);
and U20541 (N_20541,N_12326,N_14530);
or U20542 (N_20542,N_17711,N_14641);
xor U20543 (N_20543,N_11675,N_14535);
nor U20544 (N_20544,N_10510,N_10013);
nand U20545 (N_20545,N_11804,N_12290);
and U20546 (N_20546,N_12570,N_17794);
or U20547 (N_20547,N_19783,N_13395);
nand U20548 (N_20548,N_13614,N_17360);
nand U20549 (N_20549,N_17704,N_12592);
and U20550 (N_20550,N_14286,N_12286);
or U20551 (N_20551,N_17807,N_11349);
nand U20552 (N_20552,N_12561,N_14713);
nor U20553 (N_20553,N_12067,N_12591);
or U20554 (N_20554,N_15793,N_16738);
and U20555 (N_20555,N_16234,N_13047);
and U20556 (N_20556,N_15521,N_16150);
or U20557 (N_20557,N_15792,N_15304);
or U20558 (N_20558,N_10295,N_15047);
or U20559 (N_20559,N_11871,N_10540);
or U20560 (N_20560,N_15158,N_11558);
or U20561 (N_20561,N_19054,N_18379);
and U20562 (N_20562,N_19249,N_10827);
nor U20563 (N_20563,N_13028,N_16223);
nor U20564 (N_20564,N_16175,N_14784);
or U20565 (N_20565,N_15353,N_19274);
and U20566 (N_20566,N_10988,N_19353);
or U20567 (N_20567,N_16848,N_13567);
xnor U20568 (N_20568,N_12111,N_11405);
nand U20569 (N_20569,N_15623,N_10820);
and U20570 (N_20570,N_11403,N_15691);
or U20571 (N_20571,N_12750,N_19347);
nor U20572 (N_20572,N_17056,N_18834);
nand U20573 (N_20573,N_12628,N_17480);
and U20574 (N_20574,N_11900,N_16762);
nand U20575 (N_20575,N_19763,N_16571);
nand U20576 (N_20576,N_14450,N_15845);
nand U20577 (N_20577,N_16418,N_19934);
nor U20578 (N_20578,N_19745,N_11366);
and U20579 (N_20579,N_10857,N_14031);
or U20580 (N_20580,N_18646,N_17005);
nand U20581 (N_20581,N_18774,N_16345);
and U20582 (N_20582,N_13231,N_18798);
xnor U20583 (N_20583,N_17879,N_18550);
nor U20584 (N_20584,N_17624,N_11389);
nand U20585 (N_20585,N_11990,N_12471);
nand U20586 (N_20586,N_10119,N_13366);
nand U20587 (N_20587,N_19690,N_17699);
and U20588 (N_20588,N_15303,N_18592);
nor U20589 (N_20589,N_18241,N_18990);
and U20590 (N_20590,N_14825,N_13930);
or U20591 (N_20591,N_17608,N_19268);
nand U20592 (N_20592,N_15144,N_13458);
and U20593 (N_20593,N_18481,N_16933);
and U20594 (N_20594,N_13792,N_10128);
or U20595 (N_20595,N_17683,N_17500);
or U20596 (N_20596,N_19405,N_18723);
xnor U20597 (N_20597,N_18741,N_10963);
and U20598 (N_20598,N_17581,N_17281);
nand U20599 (N_20599,N_17651,N_17083);
nor U20600 (N_20600,N_13867,N_14550);
and U20601 (N_20601,N_14316,N_15739);
nor U20602 (N_20602,N_11779,N_10434);
nor U20603 (N_20603,N_18878,N_16099);
and U20604 (N_20604,N_14849,N_14109);
nor U20605 (N_20605,N_11115,N_12168);
nor U20606 (N_20606,N_11048,N_16818);
xor U20607 (N_20607,N_10747,N_16487);
and U20608 (N_20608,N_12428,N_16167);
xnor U20609 (N_20609,N_13167,N_11342);
or U20610 (N_20610,N_10129,N_11015);
and U20611 (N_20611,N_14721,N_11976);
or U20612 (N_20612,N_12379,N_12910);
nor U20613 (N_20613,N_10453,N_15587);
nand U20614 (N_20614,N_16436,N_18912);
nand U20615 (N_20615,N_17716,N_14179);
and U20616 (N_20616,N_10003,N_18612);
nand U20617 (N_20617,N_19844,N_14655);
and U20618 (N_20618,N_16629,N_10162);
nand U20619 (N_20619,N_14454,N_19067);
nor U20620 (N_20620,N_19074,N_15357);
and U20621 (N_20621,N_18007,N_10516);
or U20622 (N_20622,N_19649,N_18908);
nand U20623 (N_20623,N_11834,N_16166);
or U20624 (N_20624,N_19083,N_15837);
nand U20625 (N_20625,N_15875,N_12182);
or U20626 (N_20626,N_19640,N_18050);
xnor U20627 (N_20627,N_15668,N_15688);
and U20628 (N_20628,N_15732,N_19952);
and U20629 (N_20629,N_10012,N_10409);
nand U20630 (N_20630,N_10695,N_14125);
or U20631 (N_20631,N_10892,N_17873);
or U20632 (N_20632,N_19905,N_11155);
and U20633 (N_20633,N_10390,N_14313);
or U20634 (N_20634,N_10775,N_18172);
xor U20635 (N_20635,N_14153,N_10214);
nor U20636 (N_20636,N_16380,N_17722);
and U20637 (N_20637,N_12216,N_17935);
xnor U20638 (N_20638,N_15483,N_18687);
and U20639 (N_20639,N_12625,N_18124);
and U20640 (N_20640,N_18967,N_17201);
nand U20641 (N_20641,N_19968,N_11259);
xor U20642 (N_20642,N_15055,N_18549);
nor U20643 (N_20643,N_10036,N_10850);
nand U20644 (N_20644,N_15159,N_17654);
and U20645 (N_20645,N_19573,N_14470);
nand U20646 (N_20646,N_19085,N_11067);
nor U20647 (N_20647,N_12140,N_14302);
or U20648 (N_20648,N_19088,N_17136);
and U20649 (N_20649,N_10393,N_10720);
nor U20650 (N_20650,N_14250,N_12156);
nand U20651 (N_20651,N_13432,N_14360);
nand U20652 (N_20652,N_11402,N_17192);
xor U20653 (N_20653,N_16288,N_14717);
xor U20654 (N_20654,N_15989,N_16021);
nor U20655 (N_20655,N_15690,N_13389);
or U20656 (N_20656,N_15589,N_19865);
xnor U20657 (N_20657,N_11156,N_16113);
and U20658 (N_20658,N_14738,N_10634);
and U20659 (N_20659,N_19039,N_17412);
and U20660 (N_20660,N_19841,N_16348);
and U20661 (N_20661,N_11788,N_16661);
nand U20662 (N_20662,N_19072,N_11543);
nand U20663 (N_20663,N_11258,N_19216);
nand U20664 (N_20664,N_13550,N_13627);
xor U20665 (N_20665,N_19646,N_12565);
nor U20666 (N_20666,N_17327,N_19303);
nand U20667 (N_20667,N_12773,N_19697);
and U20668 (N_20668,N_10969,N_17320);
or U20669 (N_20669,N_12923,N_14242);
nor U20670 (N_20670,N_11164,N_12464);
nor U20671 (N_20671,N_18492,N_10590);
or U20672 (N_20672,N_12578,N_15150);
nand U20673 (N_20673,N_16306,N_12151);
and U20674 (N_20674,N_14553,N_18295);
and U20675 (N_20675,N_14639,N_11761);
and U20676 (N_20676,N_16712,N_17087);
nor U20677 (N_20677,N_16561,N_14749);
nor U20678 (N_20678,N_11962,N_19154);
and U20679 (N_20679,N_16329,N_14647);
or U20680 (N_20680,N_12636,N_10019);
and U20681 (N_20681,N_19232,N_17396);
or U20682 (N_20682,N_16999,N_15109);
nor U20683 (N_20683,N_11595,N_15225);
or U20684 (N_20684,N_16126,N_12501);
nor U20685 (N_20685,N_11264,N_14785);
nand U20686 (N_20686,N_17053,N_15650);
nor U20687 (N_20687,N_12809,N_12036);
nand U20688 (N_20688,N_10363,N_18797);
nor U20689 (N_20689,N_14574,N_16379);
or U20690 (N_20690,N_19047,N_10858);
or U20691 (N_20691,N_14860,N_16591);
or U20692 (N_20692,N_16568,N_14243);
xnor U20693 (N_20693,N_19439,N_11986);
nor U20694 (N_20694,N_11932,N_15687);
nand U20695 (N_20695,N_13712,N_15217);
nand U20696 (N_20696,N_10840,N_10377);
nand U20697 (N_20697,N_12675,N_15693);
and U20698 (N_20698,N_17775,N_18763);
or U20699 (N_20699,N_11043,N_14932);
nor U20700 (N_20700,N_11755,N_19765);
and U20701 (N_20701,N_13002,N_16926);
nand U20702 (N_20702,N_14850,N_16360);
and U20703 (N_20703,N_19791,N_19832);
and U20704 (N_20704,N_18817,N_18130);
or U20705 (N_20705,N_18094,N_14923);
or U20706 (N_20706,N_11243,N_13807);
nor U20707 (N_20707,N_15358,N_11548);
and U20708 (N_20708,N_17571,N_14298);
nand U20709 (N_20709,N_16015,N_18093);
xor U20710 (N_20710,N_16521,N_19744);
nor U20711 (N_20711,N_18875,N_19638);
nand U20712 (N_20712,N_12289,N_17377);
and U20713 (N_20713,N_13103,N_10982);
nand U20714 (N_20714,N_16672,N_19087);
nand U20715 (N_20715,N_16314,N_17085);
or U20716 (N_20716,N_19659,N_12362);
nand U20717 (N_20717,N_19916,N_10424);
and U20718 (N_20718,N_14718,N_12703);
xnor U20719 (N_20719,N_10090,N_17965);
nor U20720 (N_20720,N_16946,N_10762);
and U20721 (N_20721,N_15956,N_19867);
or U20722 (N_20722,N_15015,N_18884);
nor U20723 (N_20723,N_17040,N_16962);
nand U20724 (N_20724,N_18837,N_15504);
nand U20725 (N_20725,N_14806,N_11108);
nand U20726 (N_20726,N_19781,N_14590);
nor U20727 (N_20727,N_17322,N_18787);
nor U20728 (N_20728,N_14929,N_15061);
nand U20729 (N_20729,N_11101,N_11830);
or U20730 (N_20730,N_15703,N_16859);
nand U20731 (N_20731,N_13615,N_14768);
nor U20732 (N_20732,N_11661,N_17370);
xnor U20733 (N_20733,N_19404,N_16748);
nand U20734 (N_20734,N_18092,N_12192);
nand U20735 (N_20735,N_16310,N_10594);
and U20736 (N_20736,N_10378,N_10589);
xor U20737 (N_20737,N_17552,N_18683);
and U20738 (N_20738,N_10586,N_14342);
nand U20739 (N_20739,N_19966,N_10439);
and U20740 (N_20740,N_12960,N_14384);
or U20741 (N_20741,N_10721,N_13812);
and U20742 (N_20742,N_10001,N_11881);
xor U20743 (N_20743,N_19448,N_15962);
nor U20744 (N_20744,N_10000,N_10171);
and U20745 (N_20745,N_18791,N_18276);
xnor U20746 (N_20746,N_16188,N_12262);
or U20747 (N_20747,N_14017,N_14799);
or U20748 (N_20748,N_16182,N_18215);
nand U20749 (N_20749,N_11775,N_19507);
nand U20750 (N_20750,N_15036,N_16465);
or U20751 (N_20751,N_19132,N_12211);
and U20752 (N_20752,N_10864,N_14114);
nand U20753 (N_20753,N_19854,N_10059);
nand U20754 (N_20754,N_15670,N_15591);
and U20755 (N_20755,N_10343,N_13915);
and U20756 (N_20756,N_18968,N_19103);
nand U20757 (N_20757,N_16904,N_17344);
and U20758 (N_20758,N_18702,N_19537);
and U20759 (N_20759,N_16912,N_15716);
nand U20760 (N_20760,N_19875,N_10671);
or U20761 (N_20761,N_15184,N_18672);
and U20762 (N_20762,N_10048,N_11475);
or U20763 (N_20763,N_12368,N_17172);
xor U20764 (N_20764,N_10583,N_19983);
xor U20765 (N_20765,N_14861,N_15389);
nor U20766 (N_20766,N_19450,N_15260);
xnor U20767 (N_20767,N_11907,N_16343);
xnor U20768 (N_20768,N_19494,N_14703);
nor U20769 (N_20769,N_14792,N_13065);
xnor U20770 (N_20770,N_17576,N_11166);
and U20771 (N_20771,N_13707,N_15342);
and U20772 (N_20772,N_17106,N_12859);
xor U20773 (N_20773,N_16645,N_16797);
nand U20774 (N_20774,N_15011,N_12829);
and U20775 (N_20775,N_14736,N_18907);
xor U20776 (N_20776,N_19414,N_16821);
and U20777 (N_20777,N_12177,N_10194);
nand U20778 (N_20778,N_19965,N_15718);
nor U20779 (N_20779,N_10362,N_13874);
nand U20780 (N_20780,N_14064,N_14219);
nand U20781 (N_20781,N_12433,N_13986);
nand U20782 (N_20782,N_17203,N_18674);
nor U20783 (N_20783,N_12704,N_15810);
and U20784 (N_20784,N_17924,N_13086);
nor U20785 (N_20785,N_12564,N_14068);
xor U20786 (N_20786,N_14420,N_16276);
and U20787 (N_20787,N_13179,N_16852);
nand U20788 (N_20788,N_11044,N_17870);
and U20789 (N_20789,N_13984,N_18191);
or U20790 (N_20790,N_10729,N_16857);
nor U20791 (N_20791,N_15750,N_11681);
nor U20792 (N_20792,N_18373,N_17243);
nor U20793 (N_20793,N_11789,N_18134);
or U20794 (N_20794,N_19933,N_18809);
and U20795 (N_20795,N_14674,N_10628);
nand U20796 (N_20796,N_18536,N_12608);
nand U20797 (N_20797,N_16209,N_17102);
xnor U20798 (N_20798,N_12415,N_17697);
or U20799 (N_20799,N_19549,N_10492);
nor U20800 (N_20800,N_10070,N_10467);
or U20801 (N_20801,N_11144,N_12497);
nand U20802 (N_20802,N_16052,N_10430);
nor U20803 (N_20803,N_18594,N_13125);
or U20804 (N_20804,N_16143,N_13880);
nand U20805 (N_20805,N_12315,N_10480);
and U20806 (N_20806,N_11017,N_14981);
nand U20807 (N_20807,N_13461,N_17100);
or U20808 (N_20808,N_15065,N_13206);
xnor U20809 (N_20809,N_10648,N_18707);
nand U20810 (N_20810,N_17156,N_16706);
or U20811 (N_20811,N_16684,N_11210);
nor U20812 (N_20812,N_11920,N_16628);
nand U20813 (N_20813,N_16410,N_10330);
or U20814 (N_20814,N_13772,N_16196);
and U20815 (N_20815,N_19911,N_12963);
and U20816 (N_20816,N_16301,N_15385);
or U20817 (N_20817,N_10576,N_11359);
and U20818 (N_20818,N_17275,N_17506);
or U20819 (N_20819,N_11737,N_18278);
nand U20820 (N_20820,N_10224,N_11578);
xnor U20821 (N_20821,N_14874,N_18448);
nor U20822 (N_20822,N_11950,N_16178);
nand U20823 (N_20823,N_10446,N_13703);
or U20824 (N_20824,N_13824,N_11826);
or U20825 (N_20825,N_10717,N_13315);
nand U20826 (N_20826,N_17350,N_11365);
and U20827 (N_20827,N_14551,N_19873);
nor U20828 (N_20828,N_17007,N_13601);
or U20829 (N_20829,N_18361,N_13798);
nor U20830 (N_20830,N_14282,N_18041);
and U20831 (N_20831,N_17065,N_17361);
or U20832 (N_20832,N_15635,N_19462);
and U20833 (N_20833,N_12512,N_19824);
and U20834 (N_20834,N_11698,N_16986);
or U20835 (N_20835,N_16897,N_10160);
nand U20836 (N_20836,N_16461,N_19291);
and U20837 (N_20837,N_12319,N_15927);
and U20838 (N_20838,N_19816,N_18131);
and U20839 (N_20839,N_12983,N_11515);
nand U20840 (N_20840,N_12602,N_12402);
or U20841 (N_20841,N_14615,N_17490);
and U20842 (N_20842,N_10731,N_19108);
and U20843 (N_20843,N_17213,N_17761);
nor U20844 (N_20844,N_12807,N_19379);
nand U20845 (N_20845,N_13322,N_17496);
and U20846 (N_20846,N_15816,N_13832);
or U20847 (N_20847,N_18142,N_16760);
and U20848 (N_20848,N_19111,N_16548);
nor U20849 (N_20849,N_10608,N_17069);
xnor U20850 (N_20850,N_14009,N_17516);
nand U20851 (N_20851,N_11883,N_15937);
and U20852 (N_20852,N_19284,N_13646);
and U20853 (N_20853,N_11616,N_18662);
nor U20854 (N_20854,N_16367,N_19346);
or U20855 (N_20855,N_14120,N_19015);
nor U20856 (N_20856,N_18049,N_18300);
nand U20857 (N_20857,N_18661,N_11756);
nand U20858 (N_20858,N_18829,N_15790);
xnor U20859 (N_20859,N_11851,N_14586);
nand U20860 (N_20860,N_11283,N_17289);
nor U20861 (N_20861,N_11572,N_15463);
or U20862 (N_20862,N_13417,N_17348);
nand U20863 (N_20863,N_11944,N_17479);
or U20864 (N_20864,N_11410,N_12242);
nor U20865 (N_20865,N_12370,N_15074);
or U20866 (N_20866,N_11700,N_12339);
and U20867 (N_20867,N_12484,N_18089);
nand U20868 (N_20868,N_17063,N_19356);
nand U20869 (N_20869,N_13362,N_10314);
nor U20870 (N_20870,N_11518,N_14163);
nor U20871 (N_20871,N_19662,N_19180);
and U20872 (N_20872,N_15365,N_17849);
and U20873 (N_20873,N_14890,N_13202);
nand U20874 (N_20874,N_12702,N_12015);
and U20875 (N_20875,N_12463,N_12002);
and U20876 (N_20876,N_18477,N_10532);
xnor U20877 (N_20877,N_13554,N_16960);
nand U20878 (N_20878,N_13540,N_18105);
and U20879 (N_20879,N_15297,N_15547);
nand U20880 (N_20880,N_10706,N_16635);
nor U20881 (N_20881,N_14656,N_16386);
nand U20882 (N_20882,N_14315,N_13743);
nor U20883 (N_20883,N_15919,N_19591);
nor U20884 (N_20884,N_15573,N_11225);
nand U20885 (N_20885,N_16756,N_14916);
nand U20886 (N_20886,N_13094,N_17972);
nand U20887 (N_20887,N_13563,N_14797);
or U20888 (N_20888,N_10603,N_19784);
nor U20889 (N_20889,N_12695,N_14402);
and U20890 (N_20890,N_17114,N_18268);
nand U20891 (N_20891,N_19262,N_16202);
nand U20892 (N_20892,N_12895,N_19264);
xnor U20893 (N_20893,N_10697,N_14651);
or U20894 (N_20894,N_14082,N_14006);
nand U20895 (N_20895,N_18765,N_11073);
or U20896 (N_20896,N_19011,N_16577);
or U20897 (N_20897,N_19434,N_19505);
and U20898 (N_20898,N_15081,N_19701);
nand U20899 (N_20899,N_12145,N_11517);
or U20900 (N_20900,N_19800,N_18523);
and U20901 (N_20901,N_15110,N_15295);
and U20902 (N_20902,N_17948,N_18953);
xnor U20903 (N_20903,N_19629,N_12040);
nand U20904 (N_20904,N_15748,N_19133);
and U20905 (N_20905,N_18365,N_12928);
nand U20906 (N_20906,N_17279,N_19019);
nor U20907 (N_20907,N_10043,N_17337);
or U20908 (N_20908,N_10599,N_12408);
nand U20909 (N_20909,N_13043,N_19563);
and U20910 (N_20910,N_10367,N_13071);
xnor U20911 (N_20911,N_11975,N_12361);
and U20912 (N_20912,N_17942,N_12399);
nor U20913 (N_20913,N_14595,N_17135);
nor U20914 (N_20914,N_13709,N_10358);
or U20915 (N_20915,N_13256,N_10272);
nor U20916 (N_20916,N_17719,N_18331);
or U20917 (N_20917,N_15248,N_11936);
or U20918 (N_20918,N_11236,N_15256);
or U20919 (N_20919,N_18630,N_10561);
nand U20920 (N_20920,N_10904,N_11628);
or U20921 (N_20921,N_11308,N_19539);
and U20922 (N_20922,N_17176,N_12172);
nor U20923 (N_20923,N_10962,N_12678);
nand U20924 (N_20924,N_16755,N_13368);
or U20925 (N_20925,N_12384,N_18464);
and U20926 (N_20926,N_15789,N_19163);
and U20927 (N_20927,N_11648,N_13935);
nor U20928 (N_20928,N_16610,N_14511);
or U20929 (N_20929,N_13131,N_15763);
nor U20930 (N_20930,N_19312,N_18209);
nor U20931 (N_20931,N_10932,N_13943);
and U20932 (N_20932,N_16707,N_13009);
nand U20933 (N_20933,N_14731,N_12808);
nand U20934 (N_20934,N_16090,N_15665);
and U20935 (N_20935,N_13127,N_13048);
and U20936 (N_20936,N_12505,N_18108);
or U20937 (N_20937,N_13777,N_16294);
and U20938 (N_20938,N_19927,N_10828);
nand U20939 (N_20939,N_17161,N_13024);
xor U20940 (N_20940,N_15782,N_13793);
or U20941 (N_20941,N_13556,N_12753);
xnor U20942 (N_20942,N_15305,N_13051);
xnor U20943 (N_20943,N_11814,N_10553);
and U20944 (N_20944,N_11222,N_16115);
and U20945 (N_20945,N_12945,N_17311);
nand U20946 (N_20946,N_12118,N_18616);
or U20947 (N_20947,N_16330,N_16980);
and U20948 (N_20948,N_17189,N_17045);
nor U20949 (N_20949,N_18106,N_10989);
xnor U20950 (N_20950,N_15974,N_11545);
and U20951 (N_20951,N_16293,N_16850);
or U20952 (N_20952,N_11317,N_14005);
xor U20953 (N_20953,N_10077,N_14078);
nand U20954 (N_20954,N_17850,N_16515);
nand U20955 (N_20955,N_10812,N_14700);
and U20956 (N_20956,N_14016,N_12295);
xor U20957 (N_20957,N_13282,N_11172);
xor U20958 (N_20958,N_17765,N_12919);
and U20959 (N_20959,N_17703,N_19126);
and U20960 (N_20960,N_16423,N_19105);
nor U20961 (N_20961,N_14232,N_18970);
xnor U20962 (N_20962,N_12377,N_12423);
or U20963 (N_20963,N_10588,N_16228);
nand U20964 (N_20964,N_10197,N_15246);
and U20965 (N_20965,N_17186,N_19845);
or U20966 (N_20966,N_18285,N_12022);
xnor U20967 (N_20967,N_15583,N_12299);
nor U20968 (N_20968,N_10227,N_19696);
nor U20969 (N_20969,N_15495,N_13330);
or U20970 (N_20970,N_17910,N_14968);
or U20971 (N_20971,N_18517,N_14461);
xor U20972 (N_20972,N_12498,N_11508);
and U20973 (N_20973,N_12374,N_19871);
and U20974 (N_20974,N_17297,N_13850);
and U20975 (N_20975,N_18538,N_15647);
nand U20976 (N_20976,N_10256,N_10631);
nor U20977 (N_20977,N_13656,N_14947);
nand U20978 (N_20978,N_10623,N_17433);
and U20979 (N_20979,N_17398,N_16035);
and U20980 (N_20980,N_16567,N_19175);
nor U20981 (N_20981,N_11079,N_19377);
xnor U20982 (N_20982,N_16155,N_10082);
and U20983 (N_20983,N_14000,N_10948);
xor U20984 (N_20984,N_13665,N_17623);
and U20985 (N_20985,N_16136,N_17912);
nor U20986 (N_20986,N_18062,N_10708);
nand U20987 (N_20987,N_18321,N_19801);
nor U20988 (N_20988,N_12696,N_16217);
and U20989 (N_20989,N_12046,N_17418);
or U20990 (N_20990,N_10957,N_18955);
nor U20991 (N_20991,N_17951,N_15984);
and U20992 (N_20992,N_15585,N_11226);
nor U20993 (N_20993,N_19286,N_13290);
nor U20994 (N_20994,N_19322,N_13934);
xor U20995 (N_20995,N_16920,N_14101);
and U20996 (N_20996,N_13490,N_13755);
xor U20997 (N_20997,N_14132,N_17000);
nor U20998 (N_20998,N_16523,N_15284);
nand U20999 (N_20999,N_18583,N_18939);
and U21000 (N_21000,N_14443,N_14653);
or U21001 (N_21001,N_16029,N_11364);
nand U21002 (N_21002,N_14934,N_18075);
and U21003 (N_21003,N_12013,N_13954);
and U21004 (N_21004,N_14567,N_12553);
or U21005 (N_21005,N_10703,N_12573);
nand U21006 (N_21006,N_10972,N_16925);
nand U21007 (N_21007,N_17054,N_11000);
nor U21008 (N_21008,N_16634,N_17845);
or U21009 (N_21009,N_11499,N_19169);
and U21010 (N_21010,N_11822,N_15770);
and U21011 (N_21011,N_15214,N_16284);
nor U21012 (N_21012,N_13657,N_16539);
or U21013 (N_21013,N_14558,N_10630);
or U21014 (N_21014,N_15146,N_14197);
or U21015 (N_21015,N_12897,N_12671);
nand U21016 (N_21016,N_13331,N_18118);
or U21017 (N_21017,N_16885,N_13511);
nor U21018 (N_21018,N_14833,N_10158);
or U21019 (N_21019,N_15379,N_15001);
and U21020 (N_21020,N_16943,N_18266);
nand U21021 (N_21021,N_14705,N_13355);
nand U21022 (N_21022,N_17062,N_12606);
nor U21023 (N_21023,N_19454,N_10512);
and U21024 (N_21024,N_19244,N_11769);
nor U21025 (N_21025,N_17461,N_13129);
xnor U21026 (N_21026,N_12515,N_13359);
and U21027 (N_21027,N_14233,N_13471);
nor U21028 (N_21028,N_19259,N_12132);
and U21029 (N_21029,N_19897,N_11097);
and U21030 (N_21030,N_16124,N_14427);
or U21031 (N_21031,N_12357,N_19066);
nor U21032 (N_21032,N_15131,N_15998);
nor U21033 (N_21033,N_17696,N_19843);
and U21034 (N_21034,N_18363,N_19648);
and U21035 (N_21035,N_19757,N_16817);
and U21036 (N_21036,N_15259,N_10327);
xor U21037 (N_21037,N_17818,N_14982);
nor U21038 (N_21038,N_19515,N_17773);
and U21039 (N_21039,N_16199,N_17894);
or U21040 (N_21040,N_19551,N_12769);
xnor U21041 (N_21041,N_11702,N_13539);
and U21042 (N_21042,N_10423,N_11935);
nand U21043 (N_21043,N_16680,N_18353);
nand U21044 (N_21044,N_13414,N_12699);
or U21045 (N_21045,N_16785,N_12896);
or U21046 (N_21046,N_10143,N_19582);
or U21047 (N_21047,N_10945,N_15912);
nor U21048 (N_21048,N_14333,N_18045);
nand U21049 (N_21049,N_15243,N_12832);
and U21050 (N_21050,N_18233,N_10618);
nand U21051 (N_21051,N_19644,N_16692);
nor U21052 (N_21052,N_18156,N_10555);
nand U21053 (N_21053,N_13809,N_13621);
nor U21054 (N_21054,N_18752,N_13068);
and U21055 (N_21055,N_14741,N_19009);
or U21056 (N_21056,N_12510,N_19040);
nor U21057 (N_21057,N_13082,N_16168);
or U21058 (N_21058,N_16270,N_13181);
nand U21059 (N_21059,N_15066,N_13283);
or U21060 (N_21060,N_15957,N_11468);
and U21061 (N_21061,N_12651,N_14475);
and U21062 (N_21062,N_11399,N_14485);
and U21063 (N_21063,N_14432,N_18052);
nand U21064 (N_21064,N_16431,N_14608);
or U21065 (N_21065,N_16037,N_11112);
nor U21066 (N_21066,N_10872,N_16165);
and U21067 (N_21067,N_15384,N_19726);
nand U21068 (N_21068,N_17854,N_12041);
or U21069 (N_21069,N_14970,N_11787);
and U21070 (N_21070,N_19673,N_11116);
nand U21071 (N_21071,N_18996,N_13296);
nand U21072 (N_21072,N_12419,N_15890);
and U21073 (N_21073,N_13012,N_12030);
and U21074 (N_21074,N_15951,N_16466);
or U21075 (N_21075,N_12766,N_15731);
nor U21076 (N_21076,N_12929,N_14203);
or U21077 (N_21077,N_14403,N_14943);
and U21078 (N_21078,N_19383,N_11400);
and U21079 (N_21079,N_10838,N_12166);
nor U21080 (N_21080,N_11299,N_10572);
nor U21081 (N_21081,N_15287,N_15425);
nor U21082 (N_21082,N_16997,N_16622);
nor U21083 (N_21083,N_19932,N_18185);
nand U21084 (N_21084,N_18978,N_14410);
nand U21085 (N_21085,N_10766,N_11554);
nand U21086 (N_21086,N_15640,N_11939);
and U21087 (N_21087,N_15231,N_11511);
nor U21088 (N_21088,N_13940,N_12748);
nand U21089 (N_21089,N_12076,N_14676);
or U21090 (N_21090,N_14496,N_12793);
and U21091 (N_21091,N_12968,N_15701);
nor U21092 (N_21092,N_10517,N_17677);
nand U21093 (N_21093,N_11295,N_16681);
nor U21094 (N_21094,N_16390,N_12543);
or U21095 (N_21095,N_12712,N_18335);
nor U21096 (N_21096,N_10339,N_17848);
and U21097 (N_21097,N_11370,N_11063);
xor U21098 (N_21098,N_19806,N_18659);
or U21099 (N_21099,N_13437,N_19819);
xnor U21100 (N_21100,N_10568,N_14778);
or U21101 (N_21101,N_14451,N_12853);
or U21102 (N_21102,N_16563,N_14369);
nor U21103 (N_21103,N_13784,N_11479);
and U21104 (N_21104,N_10652,N_19529);
or U21105 (N_21105,N_14607,N_14967);
nor U21106 (N_21106,N_11401,N_11958);
nand U21107 (N_21107,N_19619,N_17300);
nand U21108 (N_21108,N_17891,N_19309);
nor U21109 (N_21109,N_13640,N_18769);
nor U21110 (N_21110,N_17825,N_18498);
nand U21111 (N_21111,N_15398,N_17215);
and U21112 (N_21112,N_11534,N_19627);
and U21113 (N_21113,N_14964,N_12519);
or U21114 (N_21114,N_10755,N_18166);
nor U21115 (N_21115,N_18340,N_14845);
and U21116 (N_21116,N_13289,N_13829);
nand U21117 (N_21117,N_11239,N_19924);
nor U21118 (N_21118,N_13216,N_16871);
or U21119 (N_21119,N_11654,N_13677);
or U21120 (N_21120,N_13234,N_19661);
and U21121 (N_21121,N_17713,N_14476);
or U21122 (N_21122,N_17543,N_17404);
nor U21123 (N_21123,N_11450,N_13529);
or U21124 (N_21124,N_18463,N_19129);
nand U21125 (N_21125,N_14347,N_19660);
or U21126 (N_21126,N_19449,N_19878);
nand U21127 (N_21127,N_16594,N_14226);
and U21128 (N_21128,N_10698,N_10315);
xor U21129 (N_21129,N_10391,N_15595);
xor U21130 (N_21130,N_17601,N_12077);
and U21131 (N_21131,N_12350,N_17556);
xnor U21132 (N_21132,N_12438,N_16264);
nor U21133 (N_21133,N_17889,N_18004);
xor U21134 (N_21134,N_16486,N_13585);
or U21135 (N_21135,N_19938,N_18919);
nand U21136 (N_21136,N_15593,N_10151);
xor U21137 (N_21137,N_14933,N_11591);
xnor U21138 (N_21138,N_17518,N_14835);
or U21139 (N_21139,N_17939,N_15115);
and U21140 (N_21140,N_11710,N_18460);
or U21141 (N_21141,N_14760,N_16144);
nor U21142 (N_21142,N_19420,N_15566);
or U21143 (N_21143,N_16213,N_18696);
nor U21144 (N_21144,N_17833,N_19564);
and U21145 (N_21145,N_12904,N_12958);
and U21146 (N_21146,N_16533,N_12927);
and U21147 (N_21147,N_14281,N_19910);
and U21148 (N_21148,N_15168,N_11923);
nand U21149 (N_21149,N_13574,N_15552);
and U21150 (N_21150,N_19705,N_16254);
nor U21151 (N_21151,N_18033,N_14334);
or U21152 (N_21152,N_19203,N_16529);
xnor U21153 (N_21153,N_10809,N_11735);
and U21154 (N_21154,N_13887,N_14312);
nand U21155 (N_21155,N_11838,N_16044);
nand U21156 (N_21156,N_10008,N_17789);
nor U21157 (N_21157,N_11396,N_18018);
or U21158 (N_21158,N_19101,N_10604);
or U21159 (N_21159,N_17665,N_12003);
and U21160 (N_21160,N_18356,N_16023);
nor U21161 (N_21161,N_14168,N_12768);
and U21162 (N_21162,N_12722,N_11524);
nor U21163 (N_21163,N_15814,N_13878);
and U21164 (N_21164,N_12092,N_18530);
nand U21165 (N_21165,N_18401,N_17049);
or U21166 (N_21166,N_18197,N_10757);
nand U21167 (N_21167,N_13358,N_14460);
nand U21168 (N_21168,N_14735,N_11579);
nand U21169 (N_21169,N_18984,N_18935);
nand U21170 (N_21170,N_15368,N_13629);
and U21171 (N_21171,N_14018,N_19857);
xor U21172 (N_21172,N_14699,N_11055);
nand U21173 (N_21173,N_16007,N_14208);
nand U21174 (N_21174,N_13825,N_13199);
and U21175 (N_21175,N_18883,N_17531);
and U21176 (N_21176,N_12153,N_15848);
and U21177 (N_21177,N_13527,N_13249);
and U21178 (N_21178,N_17778,N_19060);
or U21179 (N_21179,N_12229,N_10526);
nand U21180 (N_21180,N_13762,N_17913);
xor U21181 (N_21181,N_10665,N_15093);
nor U21182 (N_21182,N_12921,N_19006);
nand U21183 (N_21183,N_18928,N_11770);
and U21184 (N_21184,N_19273,N_11709);
or U21185 (N_21185,N_17527,N_10802);
nand U21186 (N_21186,N_17943,N_16318);
nor U21187 (N_21187,N_14378,N_18692);
nand U21188 (N_21188,N_11592,N_13191);
or U21189 (N_21189,N_14028,N_12693);
xnor U21190 (N_21190,N_19501,N_11249);
or U21191 (N_21191,N_14213,N_13662);
nand U21192 (N_21192,N_15166,N_13680);
xnor U21193 (N_21193,N_13153,N_13465);
nor U21194 (N_21194,N_12948,N_18048);
xor U21195 (N_21195,N_16716,N_16728);
and U21196 (N_21196,N_19853,N_11358);
and U21197 (N_21197,N_15281,N_14048);
nand U21198 (N_21198,N_16322,N_15586);
nand U21199 (N_21199,N_10269,N_14346);
and U21200 (N_21200,N_17969,N_13284);
nor U21201 (N_21201,N_12782,N_15437);
nor U21202 (N_21202,N_18051,N_16176);
or U21203 (N_21203,N_19919,N_18739);
and U21204 (N_21204,N_13372,N_16878);
or U21205 (N_21205,N_14382,N_15073);
and U21206 (N_21206,N_13947,N_11678);
nor U21207 (N_21207,N_10735,N_17900);
or U21208 (N_21208,N_13185,N_18442);
nand U21209 (N_21209,N_19925,N_16272);
or U21210 (N_21210,N_16440,N_16989);
and U21211 (N_21211,N_11856,N_17333);
nand U21212 (N_21212,N_13259,N_13770);
and U21213 (N_21213,N_19425,N_10952);
or U21214 (N_21214,N_11373,N_15067);
or U21215 (N_21215,N_11831,N_13740);
nor U21216 (N_21216,N_14602,N_17155);
xnor U21217 (N_21217,N_14844,N_14123);
or U21218 (N_21218,N_19336,N_17842);
or U21219 (N_21219,N_14908,N_10789);
nand U21220 (N_21220,N_18423,N_11163);
and U21221 (N_21221,N_16162,N_10460);
nor U21222 (N_21222,N_13982,N_10780);
nand U21223 (N_21223,N_19357,N_10961);
nor U21224 (N_21224,N_18319,N_11552);
nor U21225 (N_21225,N_19173,N_17207);
xnor U21226 (N_21226,N_14614,N_13560);
and U21227 (N_21227,N_17710,N_13724);
or U21228 (N_21228,N_18788,N_15285);
nor U21229 (N_21229,N_16562,N_17534);
and U21230 (N_21230,N_13463,N_17319);
nand U21231 (N_21231,N_10322,N_15592);
nor U21232 (N_21232,N_15832,N_12701);
nor U21233 (N_21233,N_19724,N_13720);
nand U21234 (N_21234,N_17033,N_13776);
nand U21235 (N_21235,N_19813,N_10232);
and U21236 (N_21236,N_15289,N_16699);
nand U21237 (N_21237,N_15596,N_19777);
and U21238 (N_21238,N_19775,N_18099);
nand U21239 (N_21239,N_14466,N_15903);
or U21240 (N_21240,N_19788,N_19953);
and U21241 (N_21241,N_11794,N_13031);
nand U21242 (N_21242,N_19670,N_16829);
and U21243 (N_21243,N_17511,N_15089);
and U21244 (N_21244,N_18333,N_17494);
or U21245 (N_21245,N_16799,N_14782);
xnor U21246 (N_21246,N_13439,N_15602);
nor U21247 (N_21247,N_16171,N_19506);
xnor U21248 (N_21248,N_13326,N_11004);
nand U21249 (N_21249,N_13008,N_12345);
nor U21250 (N_21250,N_16119,N_16928);
and U21251 (N_21251,N_16212,N_15471);
nand U21252 (N_21252,N_18487,N_11368);
and U21253 (N_21253,N_13019,N_11734);
or U21254 (N_21254,N_17025,N_15040);
xor U21255 (N_21255,N_14624,N_14244);
xor U21256 (N_21256,N_18973,N_19400);
and U21257 (N_21257,N_13100,N_13588);
nand U21258 (N_21258,N_18258,N_11849);
nor U21259 (N_21259,N_12196,N_19554);
and U21260 (N_21260,N_14525,N_14354);
xnor U21261 (N_21261,N_19251,N_12133);
or U21262 (N_21262,N_17941,N_18446);
xnor U21263 (N_21263,N_13124,N_14795);
or U21264 (N_21264,N_16711,N_14424);
or U21265 (N_21265,N_17356,N_19682);
xor U21266 (N_21266,N_14355,N_16664);
nor U21267 (N_21267,N_19200,N_13339);
nand U21268 (N_21268,N_10860,N_16082);
nor U21269 (N_21269,N_11145,N_16244);
or U21270 (N_21270,N_15314,N_16041);
nor U21271 (N_21271,N_17584,N_19948);
nor U21272 (N_21272,N_13802,N_14737);
nor U21273 (N_21273,N_17434,N_13017);
or U21274 (N_21274,N_17763,N_12878);
and U21275 (N_21275,N_17689,N_19544);
or U21276 (N_21276,N_15048,N_16275);
nor U21277 (N_21277,N_19823,N_15473);
xnor U21278 (N_21278,N_16769,N_19136);
and U21279 (N_21279,N_19899,N_13624);
and U21280 (N_21280,N_17286,N_10779);
nand U21281 (N_21281,N_11855,N_10738);
nand U21282 (N_21282,N_10258,N_10673);
nor U21283 (N_21283,N_12208,N_17920);
nand U21284 (N_21284,N_14327,N_12548);
nor U21285 (N_21285,N_10046,N_14744);
nor U21286 (N_21286,N_18509,N_11169);
nor U21287 (N_21287,N_15085,N_11690);
nor U21288 (N_21288,N_19613,N_11341);
and U21289 (N_21289,N_10066,N_18044);
xnor U21290 (N_21290,N_19369,N_10660);
or U21291 (N_21291,N_14519,N_14609);
nand U21292 (N_21292,N_13260,N_18582);
or U21293 (N_21293,N_10321,N_18892);
nor U21294 (N_21294,N_19433,N_17067);
nand U21295 (N_21295,N_16391,N_11894);
nand U21296 (N_21296,N_10981,N_16670);
xor U21297 (N_21297,N_14508,N_18116);
nand U21298 (N_21298,N_18730,N_19195);
or U21299 (N_21299,N_12406,N_13914);
nand U21300 (N_21300,N_11532,N_10139);
and U21301 (N_21301,N_17909,N_13785);
nor U21302 (N_21302,N_18084,N_16535);
xnor U21303 (N_21303,N_12101,N_15925);
xnor U21304 (N_21304,N_14247,N_13559);
xor U21305 (N_21305,N_16361,N_12754);
nor U21306 (N_21306,N_17633,N_15122);
or U21307 (N_21307,N_19327,N_10670);
and U21308 (N_21308,N_17321,N_10234);
nor U21309 (N_21309,N_15626,N_18545);
nor U21310 (N_21310,N_11020,N_18218);
and U21311 (N_21311,N_17668,N_16569);
or U21312 (N_21312,N_11275,N_12716);
and U21313 (N_21313,N_19711,N_16650);
and U21314 (N_21314,N_17524,N_17928);
nor U21315 (N_21315,N_11708,N_19316);
and U21316 (N_21316,N_11241,N_17349);
nor U21317 (N_21317,N_10329,N_16905);
or U21318 (N_21318,N_17152,N_14093);
and U21319 (N_21319,N_15215,N_19543);
xnor U21320 (N_21320,N_17904,N_19960);
and U21321 (N_21321,N_16003,N_16875);
nand U21322 (N_21322,N_12105,N_18111);
nand U21323 (N_21323,N_13318,N_13945);
nor U21324 (N_21324,N_14783,N_13186);
and U21325 (N_21325,N_19820,N_15604);
nand U21326 (N_21326,N_10344,N_18948);
and U21327 (N_21327,N_13894,N_11313);
or U21328 (N_21328,N_12935,N_13715);
and U21329 (N_21329,N_12648,N_16901);
nand U21330 (N_21330,N_14857,N_18786);
and U21331 (N_21331,N_15783,N_14887);
nand U21332 (N_21332,N_14704,N_19443);
nor U21333 (N_21333,N_18122,N_15945);
and U21334 (N_21334,N_13913,N_16062);
and U21335 (N_21335,N_17118,N_13147);
or U21336 (N_21336,N_14440,N_16197);
or U21337 (N_21337,N_14145,N_12014);
nand U21338 (N_21338,N_11501,N_11757);
and U21339 (N_21339,N_19698,N_17730);
nor U21340 (N_21340,N_18853,N_16245);
xor U21341 (N_21341,N_10966,N_10924);
nor U21342 (N_21342,N_10010,N_12837);
nand U21343 (N_21343,N_14764,N_19142);
nand U21344 (N_21344,N_15039,N_11784);
and U21345 (N_21345,N_15678,N_18925);
nor U21346 (N_21346,N_11274,N_14957);
nor U21347 (N_21347,N_12855,N_16511);
and U21348 (N_21348,N_13287,N_17269);
nor U21349 (N_21349,N_10009,N_14373);
nor U21350 (N_21350,N_16084,N_10396);
and U21351 (N_21351,N_18184,N_16630);
or U21352 (N_21352,N_11305,N_12536);
nor U21353 (N_21353,N_16277,N_16811);
and U21354 (N_21354,N_15883,N_11242);
and U21355 (N_21355,N_14075,N_10091);
nand U21356 (N_21356,N_11520,N_10023);
or U21357 (N_21357,N_10607,N_14321);
and U21358 (N_21358,N_10830,N_11347);
or U21359 (N_21359,N_12880,N_14335);
or U21360 (N_21360,N_11081,N_14740);
or U21361 (N_21361,N_14495,N_10361);
and U21362 (N_21362,N_18628,N_13566);
or U21363 (N_21363,N_17474,N_13870);
xnor U21364 (N_21364,N_10761,N_12324);
or U21365 (N_21365,N_12811,N_10855);
and U21366 (N_21366,N_18163,N_16780);
nor U21367 (N_21367,N_15336,N_10386);
xor U21368 (N_21368,N_11774,N_16894);
or U21369 (N_21369,N_16921,N_11934);
or U21370 (N_21370,N_10038,N_14351);
and U21371 (N_21371,N_15833,N_14885);
nand U21372 (N_21372,N_10882,N_13517);
nor U21373 (N_21373,N_16916,N_10123);
and U21374 (N_21374,N_15947,N_18091);
or U21375 (N_21375,N_19092,N_19431);
nor U21376 (N_21376,N_16526,N_17686);
nand U21377 (N_21377,N_17985,N_19635);
and U21378 (N_21378,N_14600,N_12035);
nand U21379 (N_21379,N_11903,N_19091);
nor U21380 (N_21380,N_15086,N_14306);
nand U21381 (N_21381,N_17178,N_11388);
nor U21382 (N_21382,N_11449,N_12281);
nor U21383 (N_21383,N_16813,N_13875);
or U21384 (N_21384,N_16918,N_19426);
nand U21385 (N_21385,N_11448,N_12973);
nor U21386 (N_21386,N_16565,N_16536);
xor U21387 (N_21387,N_14308,N_16030);
or U21388 (N_21388,N_13406,N_15955);
and U21389 (N_21389,N_18326,N_18434);
and U21390 (N_21390,N_15607,N_16554);
nand U21391 (N_21391,N_14819,N_14326);
xor U21392 (N_21392,N_18024,N_15611);
nand U21393 (N_21393,N_10287,N_13488);
nor U21394 (N_21394,N_12254,N_13959);
or U21395 (N_21395,N_15606,N_19732);
nand U21396 (N_21396,N_16100,N_17352);
nand U21397 (N_21397,N_18785,N_14318);
xnor U21398 (N_21398,N_13751,N_13219);
nand U21399 (N_21399,N_19463,N_16384);
nand U21400 (N_21400,N_11122,N_16203);
nor U21401 (N_21401,N_11824,N_14304);
nand U21402 (N_21402,N_11876,N_15035);
nor U21403 (N_21403,N_10593,N_16695);
nor U21404 (N_21404,N_12816,N_10725);
or U21405 (N_21405,N_16214,N_14510);
nand U21406 (N_21406,N_16405,N_15027);
and U21407 (N_21407,N_14826,N_11465);
xor U21408 (N_21408,N_13939,N_15101);
and U21409 (N_21409,N_19051,N_18602);
nor U21410 (N_21410,N_19374,N_14395);
nand U21411 (N_21411,N_18473,N_14300);
or U21412 (N_21412,N_19181,N_18096);
nand U21413 (N_21413,N_16078,N_11211);
and U21414 (N_21414,N_14482,N_10547);
nand U21415 (N_21415,N_10647,N_16490);
nand U21416 (N_21416,N_13600,N_10524);
nand U21417 (N_21417,N_19976,N_12367);
or U21418 (N_21418,N_12520,N_13159);
xnor U21419 (N_21419,N_12135,N_14178);
nor U21420 (N_21420,N_16560,N_12209);
nand U21421 (N_21421,N_11065,N_12518);
nor U21422 (N_21422,N_18068,N_13204);
nor U21423 (N_21423,N_11626,N_17838);
nor U21424 (N_21424,N_18768,N_15743);
and U21425 (N_21425,N_19581,N_14494);
and U21426 (N_21426,N_14851,N_16489);
or U21427 (N_21427,N_17607,N_12542);
and U21428 (N_21428,N_10994,N_10468);
nor U21429 (N_21429,N_12442,N_16323);
and U21430 (N_21430,N_18393,N_15419);
nor U21431 (N_21431,N_18387,N_18038);
and U21432 (N_21432,N_15537,N_18777);
xnor U21433 (N_21433,N_12781,N_16686);
xnor U21434 (N_21434,N_14552,N_14150);
or U21435 (N_21435,N_17239,N_16427);
nor U21436 (N_21436,N_17060,N_14727);
and U21437 (N_21437,N_18040,N_11764);
and U21438 (N_21438,N_11346,N_15570);
nand U21439 (N_21439,N_17238,N_13266);
nor U21440 (N_21440,N_11519,N_11599);
and U21441 (N_21441,N_18563,N_19172);
or U21442 (N_21442,N_11652,N_12232);
xnor U21443 (N_21443,N_14350,N_16474);
and U21444 (N_21444,N_14331,N_14730);
nand U21445 (N_21445,N_16479,N_12861);
and U21446 (N_21446,N_12170,N_18959);
nor U21447 (N_21447,N_10111,N_14061);
nand U21448 (N_21448,N_15916,N_10778);
nor U21449 (N_21449,N_19716,N_14416);
and U21450 (N_21450,N_17212,N_10083);
nand U21451 (N_21451,N_14807,N_11668);
xor U21452 (N_21452,N_12328,N_12645);
xor U21453 (N_21453,N_17868,N_16117);
and U21454 (N_21454,N_14013,N_14489);
nor U21455 (N_21455,N_11497,N_18359);
nor U21456 (N_21456,N_14862,N_10995);
nand U21457 (N_21457,N_10753,N_15313);
nand U21458 (N_21458,N_15755,N_14381);
nand U21459 (N_21459,N_13468,N_14255);
and U21460 (N_21460,N_11639,N_11781);
nor U21461 (N_21461,N_15964,N_10300);
and U21462 (N_21462,N_18547,N_17339);
and U21463 (N_21463,N_15663,N_11474);
nor U21464 (N_21464,N_13907,N_13379);
nand U21465 (N_21465,N_11408,N_18924);
xor U21466 (N_21466,N_13593,N_13401);
or U21467 (N_21467,N_18539,N_11813);
nor U21468 (N_21468,N_10169,N_15108);
or U21469 (N_21469,N_17472,N_16639);
or U21470 (N_21470,N_17802,N_11653);
nand U21471 (N_21471,N_10811,N_18507);
nand U21472 (N_21472,N_17257,N_11743);
nand U21473 (N_21473,N_19576,N_18267);
or U21474 (N_21474,N_19595,N_13291);
nor U21475 (N_21475,N_10294,N_10037);
or U21476 (N_21476,N_17649,N_17579);
and U21477 (N_21477,N_10061,N_19261);
nand U21478 (N_21478,N_17650,N_19995);
xnor U21479 (N_21479,N_13590,N_15247);
and U21480 (N_21480,N_11244,N_16723);
nand U21481 (N_21481,N_13789,N_12673);
or U21482 (N_21482,N_12190,N_19656);
xnor U21483 (N_21483,N_17072,N_11825);
or U21484 (N_21484,N_18986,N_11573);
nor U21485 (N_21485,N_12993,N_15464);
and U21486 (N_21486,N_18061,N_16463);
and U21487 (N_21487,N_17606,N_15865);
or U21488 (N_21488,N_11682,N_10419);
or U21489 (N_21489,N_15588,N_14119);
xnor U21490 (N_21490,N_10041,N_16258);
or U21491 (N_21491,N_10474,N_11303);
or U21492 (N_21492,N_16019,N_12764);
nor U21493 (N_21493,N_17994,N_17489);
or U21494 (N_21494,N_15987,N_10470);
nor U21495 (N_21495,N_18813,N_19157);
nand U21496 (N_21496,N_18158,N_11866);
and U21497 (N_21497,N_16932,N_16467);
or U21498 (N_21498,N_11741,N_12654);
or U21499 (N_21499,N_18534,N_15799);
nand U21500 (N_21500,N_19984,N_13267);
and U21501 (N_21501,N_14945,N_13717);
or U21502 (N_21502,N_11240,N_10335);
xnor U21503 (N_21503,N_17742,N_15139);
nand U21504 (N_21504,N_19931,N_12911);
xnor U21505 (N_21505,N_10006,N_17158);
and U21506 (N_21506,N_12045,N_10824);
xor U21507 (N_21507,N_18531,N_13083);
and U21508 (N_21508,N_12382,N_11760);
nor U21509 (N_21509,N_15896,N_14001);
or U21510 (N_21510,N_15493,N_11759);
and U21511 (N_21511,N_16257,N_12814);
or U21512 (N_21512,N_17664,N_17116);
and U21513 (N_21513,N_10183,N_14985);
or U21514 (N_21514,N_19846,N_11233);
or U21515 (N_21515,N_15230,N_17283);
and U21516 (N_21516,N_13066,N_12977);
and U21517 (N_21517,N_13628,N_18469);
and U21518 (N_21518,N_17630,N_12801);
nand U21519 (N_21519,N_13352,N_12019);
xnor U21520 (N_21520,N_17897,N_11718);
or U21521 (N_21521,N_16659,N_10832);
and U21522 (N_21522,N_19523,N_14128);
and U21523 (N_21523,N_11618,N_18745);
or U21524 (N_21524,N_10602,N_16074);
and U21525 (N_21525,N_13040,N_18916);
nor U21526 (N_21526,N_16295,N_15892);
xnor U21527 (N_21527,N_13925,N_17594);
and U21528 (N_21528,N_16606,N_11960);
nand U21529 (N_21529,N_14094,N_12117);
nor U21530 (N_21530,N_16740,N_15534);
or U21531 (N_21531,N_19196,N_13218);
nor U21532 (N_21532,N_16733,N_17240);
and U21533 (N_21533,N_19893,N_12940);
and U21534 (N_21534,N_19519,N_11877);
and U21535 (N_21535,N_11732,N_19500);
nor U21536 (N_21536,N_18115,N_17498);
nor U21537 (N_21537,N_17678,N_16534);
nand U21538 (N_21538,N_10354,N_13898);
and U21539 (N_21539,N_17429,N_12875);
nor U21540 (N_21540,N_14557,N_18043);
nor U21541 (N_21541,N_13744,N_18159);
and U21542 (N_21542,N_14560,N_16819);
xor U21543 (N_21543,N_16841,N_12667);
or U21544 (N_21544,N_18814,N_17927);
and U21545 (N_21545,N_10913,N_15209);
or U21546 (N_21546,N_16040,N_18047);
or U21547 (N_21547,N_17569,N_18839);
xnor U21548 (N_21548,N_15194,N_13711);
xor U21549 (N_21549,N_16332,N_10923);
nand U21550 (N_21550,N_17964,N_16619);
or U21551 (N_21551,N_10279,N_18013);
nor U21552 (N_21552,N_11957,N_14366);
nand U21553 (N_21553,N_10591,N_18749);
and U21554 (N_21554,N_12124,N_18449);
or U21555 (N_21555,N_11854,N_11502);
or U21556 (N_21556,N_19280,N_12659);
nand U21557 (N_21557,N_11151,N_14787);
nand U21558 (N_21558,N_10311,N_10292);
and U21559 (N_21559,N_11272,N_16382);
or U21560 (N_21560,N_15734,N_19250);
and U21561 (N_21561,N_19318,N_16761);
and U21562 (N_21562,N_10455,N_18506);
and U21563 (N_21563,N_12502,N_11815);
nor U21564 (N_21564,N_11898,N_12456);
nand U21565 (N_21565,N_19446,N_10164);
nand U21566 (N_21566,N_19735,N_18810);
or U21567 (N_21567,N_10987,N_19645);
nor U21568 (N_21568,N_12849,N_10275);
and U21569 (N_21569,N_12267,N_10861);
nand U21570 (N_21570,N_13039,N_14536);
nor U21571 (N_21571,N_13937,N_15444);
nor U21572 (N_21572,N_11208,N_14044);
and U21573 (N_21573,N_17949,N_18846);
and U21574 (N_21574,N_11455,N_19002);
or U21575 (N_21575,N_10688,N_13868);
and U21576 (N_21576,N_17903,N_16002);
or U21577 (N_21577,N_13594,N_14926);
and U21578 (N_21578,N_10956,N_13436);
nand U21579 (N_21579,N_19403,N_17470);
xnor U21580 (N_21580,N_11383,N_16138);
xnor U21581 (N_21581,N_15840,N_19388);
nor U21582 (N_21582,N_19684,N_11859);
nand U21583 (N_21583,N_18585,N_17456);
or U21584 (N_21584,N_13719,N_15200);
and U21585 (N_21585,N_17578,N_11140);
nor U21586 (N_21586,N_18425,N_14580);
and U21587 (N_21587,N_15056,N_15164);
or U21588 (N_21588,N_19479,N_11085);
nor U21589 (N_21589,N_17886,N_10507);
nand U21590 (N_21590,N_15879,N_16032);
or U21591 (N_21591,N_12042,N_16232);
nor U21592 (N_21592,N_14452,N_13879);
nand U21593 (N_21593,N_12725,N_11392);
and U21594 (N_21594,N_12265,N_15578);
xor U21595 (N_21595,N_12366,N_13530);
or U21596 (N_21596,N_19408,N_14079);
nand U21597 (N_21597,N_15273,N_12306);
nor U21598 (N_21598,N_16696,N_13795);
nand U21599 (N_21599,N_19568,N_15064);
and U21600 (N_21600,N_18364,N_14858);
xnor U21601 (N_21601,N_10569,N_12743);
xnor U21602 (N_21602,N_16844,N_11840);
nand U21603 (N_21603,N_17892,N_11367);
xor U21604 (N_21604,N_15715,N_19178);
or U21605 (N_21605,N_14696,N_18922);
nor U21606 (N_21606,N_10783,N_17612);
nor U21607 (N_21607,N_14015,N_10529);
or U21608 (N_21608,N_10058,N_10563);
or U21609 (N_21609,N_19453,N_14138);
nand U21610 (N_21610,N_13140,N_15179);
and U21611 (N_21611,N_14288,N_18720);
nand U21612 (N_21612,N_12779,N_19127);
or U21613 (N_21613,N_14999,N_18346);
or U21614 (N_21614,N_19939,N_10277);
nand U21615 (N_21615,N_17797,N_10841);
and U21616 (N_21616,N_12359,N_19731);
and U21617 (N_21617,N_14469,N_10405);
nor U21618 (N_21618,N_13018,N_10931);
nand U21619 (N_21619,N_15459,N_18711);
and U21620 (N_21620,N_19972,N_18993);
xnor U21621 (N_21621,N_18802,N_14671);
nor U21622 (N_21622,N_11325,N_13909);
nor U21623 (N_21623,N_19362,N_12783);
nand U21624 (N_21624,N_17750,N_15233);
nor U21625 (N_21625,N_19146,N_17220);
or U21626 (N_21626,N_14417,N_17720);
or U21627 (N_21627,N_11292,N_16274);
or U21628 (N_21628,N_18920,N_18028);
nand U21629 (N_21629,N_12436,N_11658);
nor U21630 (N_21630,N_14521,N_11011);
nand U21631 (N_21631,N_19986,N_10979);
and U21632 (N_21632,N_14891,N_14156);
nand U21633 (N_21633,N_18528,N_17463);
nand U21634 (N_21634,N_11816,N_10489);
nor U21635 (N_21635,N_17989,N_19977);
nand U21636 (N_21636,N_13783,N_19017);
nand U21637 (N_21637,N_12920,N_12860);
and U21638 (N_21638,N_10777,N_14756);
or U21639 (N_21639,N_18022,N_15154);
and U21640 (N_21640,N_16362,N_19306);
nor U21641 (N_21641,N_11819,N_12724);
and U21642 (N_21642,N_16580,N_13360);
nand U21643 (N_21643,N_19706,N_15468);
and U21644 (N_21644,N_13122,N_14032);
or U21645 (N_21645,N_16842,N_16601);
xor U21646 (N_21646,N_19719,N_16394);
nor U21647 (N_21647,N_11576,N_13419);
or U21648 (N_21648,N_13570,N_14545);
xor U21649 (N_21649,N_10506,N_18455);
nor U21650 (N_21650,N_19587,N_14561);
and U21651 (N_21651,N_17682,N_10433);
xor U21652 (N_21652,N_18416,N_17477);
xor U21653 (N_21653,N_18413,N_12340);
and U21654 (N_21654,N_15525,N_15070);
and U21655 (N_21655,N_10063,N_17585);
nor U21656 (N_21656,N_12327,N_13162);
nand U21657 (N_21657,N_13426,N_10210);
nor U21658 (N_21658,N_11982,N_10819);
nand U21659 (N_21659,N_17588,N_12871);
and U21660 (N_21660,N_15644,N_14225);
and U21661 (N_21661,N_15046,N_17874);
nor U21662 (N_21662,N_11862,N_10084);
or U21663 (N_21663,N_10518,N_17198);
or U21664 (N_21664,N_19971,N_18557);
nor U21665 (N_21665,N_13876,N_15548);
nand U21666 (N_21666,N_11526,N_16111);
nor U21667 (N_21667,N_15766,N_10881);
nor U21668 (N_21668,N_18126,N_13503);
or U21669 (N_21669,N_11507,N_13226);
or U21670 (N_21670,N_13063,N_11567);
or U21671 (N_21671,N_10469,N_11276);
and U21672 (N_21672,N_14579,N_13917);
nor U21673 (N_21673,N_12819,N_16118);
and U21674 (N_21674,N_18652,N_19256);
and U21675 (N_21675,N_10893,N_16011);
and U21676 (N_21676,N_13448,N_18420);
or U21677 (N_21677,N_17661,N_18129);
nor U21678 (N_21678,N_12256,N_17078);
or U21679 (N_21679,N_13222,N_11956);
nand U21680 (N_21680,N_12088,N_10804);
nor U21681 (N_21681,N_10088,N_15149);
nand U21682 (N_21682,N_16950,N_16839);
or U21683 (N_21683,N_17411,N_16374);
nand U21684 (N_21684,N_12500,N_13106);
or U21685 (N_21685,N_18161,N_17028);
nand U21686 (N_21686,N_18283,N_12434);
nand U21687 (N_21687,N_14377,N_14344);
nor U21688 (N_21688,N_12470,N_16746);
nor U21689 (N_21689,N_13025,N_12049);
and U21690 (N_21690,N_17657,N_10239);
and U21691 (N_21691,N_16344,N_15851);
nand U21692 (N_21692,N_19120,N_15780);
or U21693 (N_21693,N_16302,N_13236);
nor U21694 (N_21694,N_16017,N_17416);
and U21695 (N_21695,N_18565,N_12687);
and U21696 (N_21696,N_10382,N_19900);
or U21697 (N_21697,N_16578,N_10186);
nand U21698 (N_21698,N_18759,N_10073);
or U21699 (N_21699,N_18465,N_12385);
nor U21700 (N_21700,N_16383,N_18647);
or U21701 (N_21701,N_12535,N_10352);
xor U21702 (N_21702,N_15202,N_10173);
nand U21703 (N_21703,N_11667,N_15079);
or U21704 (N_21704,N_18840,N_16225);
nand U21705 (N_21705,N_10395,N_15943);
or U21706 (N_21706,N_19611,N_17946);
nor U21707 (N_21707,N_13433,N_17272);
or U21708 (N_21708,N_16055,N_19278);
nor U21709 (N_21709,N_14701,N_14060);
nand U21710 (N_21710,N_12813,N_13910);
xor U21711 (N_21711,N_16179,N_18279);
and U21712 (N_21712,N_15319,N_17030);
or U21713 (N_21713,N_13491,N_13060);
and U21714 (N_21714,N_19903,N_10388);
xnor U21715 (N_21715,N_14506,N_11254);
or U21716 (N_21716,N_19904,N_16387);
nand U21717 (N_21717,N_10018,N_11190);
nor U21718 (N_21718,N_14759,N_16697);
nor U21719 (N_21719,N_17139,N_10278);
nand U21720 (N_21720,N_18803,N_13721);
nand U21721 (N_21721,N_15400,N_19277);
xnor U21722 (N_21722,N_13928,N_16899);
nand U21723 (N_21723,N_17366,N_17256);
nor U21724 (N_21724,N_17559,N_17468);
or U21725 (N_21725,N_16292,N_19685);
nor U21726 (N_21726,N_18644,N_12933);
nand U21727 (N_21727,N_17860,N_14442);
xnor U21728 (N_21728,N_15432,N_12390);
or U21729 (N_21729,N_19148,N_13808);
or U21730 (N_21730,N_12159,N_18223);
and U21731 (N_21731,N_15714,N_19164);
and U21732 (N_21732,N_13698,N_18546);
and U21733 (N_21733,N_14218,N_11284);
nand U21734 (N_21734,N_19109,N_13912);
and U21735 (N_21735,N_12020,N_16425);
and U21736 (N_21736,N_13990,N_11973);
nand U21737 (N_21737,N_18575,N_12337);
nor U21738 (N_21738,N_13444,N_12828);
nor U21739 (N_21739,N_13152,N_16187);
xor U21740 (N_21740,N_17808,N_18395);
and U21741 (N_21741,N_10055,N_18836);
or U21742 (N_21742,N_19236,N_16354);
and U21743 (N_21743,N_16655,N_11090);
xor U21744 (N_21744,N_13184,N_19979);
nor U21745 (N_21745,N_12257,N_12247);
and U21746 (N_21746,N_14774,N_18877);
nor U21747 (N_21747,N_13669,N_15835);
or U21748 (N_21748,N_18974,N_14505);
nor U21749 (N_21749,N_19639,N_15930);
and U21750 (N_21750,N_19018,N_18511);
nor U21751 (N_21751,N_12249,N_11407);
or U21752 (N_21752,N_17095,N_17271);
or U21753 (N_21753,N_18445,N_14650);
or U21754 (N_21754,N_18600,N_14531);
nand U21755 (N_21755,N_19514,N_16151);
nor U21756 (N_21756,N_14183,N_13295);
nand U21757 (N_21757,N_11142,N_15639);
or U21758 (N_21758,N_14702,N_13460);
or U21759 (N_21759,N_19043,N_10285);
or U21760 (N_21760,N_19252,N_16237);
nor U21761 (N_21761,N_10600,N_11914);
nor U21762 (N_21762,N_10490,N_13528);
and U21763 (N_21763,N_12346,N_14363);
nand U21764 (N_21764,N_12728,N_16404);
or U21765 (N_21765,N_15513,N_17718);
nand U21766 (N_21766,N_11125,N_11677);
or U21767 (N_21767,N_14155,N_13344);
nor U21768 (N_21768,N_19325,N_11858);
and U21769 (N_21769,N_10217,N_13016);
nand U21770 (N_21770,N_15021,N_18117);
xnor U21771 (N_21771,N_12891,N_19401);
or U21772 (N_21772,N_11248,N_10312);
nor U21773 (N_21773,N_13697,N_18407);
xor U21774 (N_21774,N_19202,N_18663);
nand U21775 (N_21775,N_16315,N_14714);
or U21776 (N_21776,N_13428,N_18518);
nor U21777 (N_21777,N_10839,N_15292);
or U21778 (N_21778,N_14873,N_17988);
nor U21779 (N_21779,N_15929,N_11569);
nand U21780 (N_21780,N_17431,N_17747);
xor U21781 (N_21781,N_11808,N_18625);
nor U21782 (N_21782,N_10266,N_18452);
nand U21783 (N_21783,N_10704,N_17273);
or U21784 (N_21784,N_11420,N_13804);
xnor U21785 (N_21785,N_19130,N_15938);
nand U21786 (N_21786,N_18657,N_17805);
or U21787 (N_21787,N_18272,N_16480);
nand U21788 (N_21788,N_12762,N_14428);
nand U21789 (N_21789,N_18776,N_13839);
nor U21790 (N_21790,N_13846,N_15899);
nor U21791 (N_21791,N_15967,N_16038);
or U21792 (N_21792,N_16129,N_17400);
and U21793 (N_21793,N_16191,N_13950);
and U21794 (N_21794,N_12439,N_10120);
nor U21795 (N_21795,N_18500,N_18871);
nand U21796 (N_21796,N_16192,N_18444);
or U21797 (N_21797,N_13938,N_17525);
xnor U21798 (N_21798,N_18174,N_16122);
xnor U21799 (N_21799,N_14706,N_18078);
and U21800 (N_21800,N_11723,N_15538);
nor U21801 (N_21801,N_10758,N_16648);
xnor U21802 (N_21802,N_17774,N_11200);
or U21803 (N_21803,N_17793,N_18264);
or U21804 (N_21804,N_11742,N_11149);
xor U21805 (N_21805,N_12872,N_17132);
nand U21806 (N_21806,N_15348,N_14839);
or U21807 (N_21807,N_15699,N_11512);
nand U21808 (N_21808,N_13695,N_15784);
or U21809 (N_21809,N_10450,N_18229);
nand U21810 (N_21810,N_19770,N_15649);
or U21811 (N_21811,N_15991,N_15265);
nor U21812 (N_21812,N_17354,N_13427);
and U21813 (N_21813,N_11714,N_18438);
and U21814 (N_21814,N_10076,N_12335);
nand U21815 (N_21815,N_14855,N_19292);
and U21816 (N_21816,N_11629,N_15422);
xor U21817 (N_21817,N_11087,N_15296);
nand U21818 (N_21818,N_12060,N_17379);
and U21819 (N_21819,N_16451,N_13618);
xor U21820 (N_21820,N_17331,N_18399);
and U21821 (N_21821,N_12708,N_13497);
or U21822 (N_21822,N_19219,N_14770);
or U21823 (N_21823,N_10415,N_17590);
nand U21824 (N_21824,N_10380,N_18470);
nor U21825 (N_21825,N_11685,N_16290);
or U21826 (N_21826,N_13022,N_17732);
or U21827 (N_21827,N_13097,N_10328);
or U21828 (N_21828,N_18693,N_12767);
nand U21829 (N_21829,N_18102,N_15123);
xnor U21830 (N_21830,N_15133,N_15672);
and U21831 (N_21831,N_16366,N_10144);
and U21832 (N_21832,N_17439,N_10368);
nand U21833 (N_21833,N_19651,N_17758);
and U21834 (N_21834,N_10346,N_11695);
and U21835 (N_21835,N_13405,N_18101);
or U21836 (N_21836,N_11160,N_13353);
nor U21837 (N_21837,N_14900,N_18027);
and U21838 (N_21838,N_13449,N_17562);
or U21839 (N_21839,N_17039,N_19839);
nor U21840 (N_21840,N_11596,N_16439);
and U21841 (N_21841,N_16296,N_13737);
xor U21842 (N_21842,N_16940,N_10847);
nor U21843 (N_21843,N_18947,N_15125);
nand U21844 (N_21844,N_14587,N_15706);
and U21845 (N_21845,N_15221,N_12966);
and U21846 (N_21846,N_15479,N_10397);
nand U21847 (N_21847,N_11987,N_10657);
and U21848 (N_21848,N_17781,N_16611);
and U21849 (N_21849,N_17616,N_17495);
and U21850 (N_21850,N_18193,N_14116);
or U21851 (N_21851,N_14769,N_18243);
and U21852 (N_21852,N_13575,N_16892);
nor U21853 (N_21853,N_12079,N_10829);
or U21854 (N_21854,N_18519,N_12820);
and U21855 (N_21855,N_17835,N_18632);
nor U21856 (N_21856,N_18964,N_15774);
nand U21857 (N_21857,N_17539,N_15112);
and U21858 (N_21858,N_12937,N_13172);
nand U21859 (N_21859,N_17632,N_10650);
nand U21860 (N_21860,N_17193,N_14214);
and U21861 (N_21861,N_15948,N_13997);
and U21862 (N_21862,N_17962,N_11683);
nor U21863 (N_21863,N_10282,N_17483);
xnor U21864 (N_21864,N_11477,N_12932);
nor U21865 (N_21865,N_11369,N_18042);
nand U21866 (N_21866,N_13177,N_17316);
nor U21867 (N_21867,N_16068,N_18419);
and U21868 (N_21868,N_11631,N_11268);
and U21869 (N_21869,N_16579,N_13834);
and U21870 (N_21870,N_11100,N_10483);
xor U21871 (N_21871,N_16013,N_19073);
nor U21872 (N_21872,N_10767,N_12691);
nand U21873 (N_21873,N_12413,N_18781);
or U21874 (N_21874,N_15854,N_14198);
nand U21875 (N_21875,N_13391,N_16141);
or U21876 (N_21876,N_14052,N_18467);
nand U21877 (N_21877,N_18533,N_17803);
and U21878 (N_21878,N_15410,N_16482);
nand U21879 (N_21879,N_19320,N_14081);
and U21880 (N_21880,N_17259,N_18148);
nor U21881 (N_21881,N_19233,N_18577);
nor U21882 (N_21882,N_10252,N_12072);
and U21883 (N_21883,N_19350,N_16583);
nand U21884 (N_21884,N_13154,N_10712);
or U21885 (N_21885,N_12207,N_10447);
nor U21886 (N_21886,N_18551,N_17017);
or U21887 (N_21887,N_10316,N_10669);
nor U21888 (N_21888,N_18064,N_15397);
and U21889 (N_21889,N_14258,N_18617);
or U21890 (N_21890,N_16682,N_12276);
or U21891 (N_21891,N_16065,N_15173);
and U21892 (N_21892,N_12112,N_19215);
nor U21893 (N_21893,N_15002,N_18706);
or U21894 (N_21894,N_18029,N_14556);
nor U21895 (N_21895,N_13710,N_18889);
and U21896 (N_21896,N_11413,N_14907);
or U21897 (N_21897,N_18136,N_16792);
or U21898 (N_21898,N_13346,N_18943);
and U21899 (N_21899,N_17918,N_19214);
nand U21900 (N_21900,N_18909,N_13217);
xor U21901 (N_21901,N_13582,N_18762);
xnor U21902 (N_21902,N_11949,N_14668);
and U21903 (N_21903,N_10410,N_14765);
xnor U21904 (N_21904,N_17447,N_12652);
nor U21905 (N_21905,N_15097,N_12881);
nor U21906 (N_21906,N_15958,N_13149);
or U21907 (N_21907,N_13240,N_17993);
nor U21908 (N_21908,N_13995,N_10159);
nor U21909 (N_21909,N_17893,N_18368);
nand U21910 (N_21910,N_13764,N_15590);
or U21911 (N_21911,N_11912,N_16243);
nand U21912 (N_21912,N_17731,N_14745);
and U21913 (N_21913,N_14337,N_14245);
nor U21914 (N_21914,N_13313,N_17358);
or U21915 (N_21915,N_11664,N_13840);
nor U21916 (N_21916,N_18493,N_18615);
nand U21917 (N_21917,N_19742,N_18972);
nor U21918 (N_21918,N_11899,N_11948);
or U21919 (N_21919,N_16034,N_17406);
nand U21920 (N_21920,N_17223,N_18153);
nor U21921 (N_21921,N_10515,N_19535);
or U21922 (N_21922,N_12697,N_19328);
and U21923 (N_21923,N_11379,N_15033);
nand U21924 (N_21924,N_16250,N_16858);
and U21925 (N_21925,N_16195,N_11665);
nand U21926 (N_21926,N_10773,N_11273);
nor U21927 (N_21927,N_17252,N_11672);
or U21928 (N_21928,N_10130,N_12550);
nor U21929 (N_21929,N_12236,N_10863);
and U21930 (N_21930,N_15418,N_15852);
nor U21931 (N_21931,N_10910,N_15965);
or U21932 (N_21932,N_19665,N_15721);
nor U21933 (N_21933,N_14691,N_18887);
and U21934 (N_21934,N_13270,N_11811);
or U21935 (N_21935,N_13670,N_12640);
or U21936 (N_21936,N_17536,N_17415);
nor U21937 (N_21937,N_19817,N_18622);
or U21938 (N_21938,N_17890,N_17517);
and U21939 (N_21939,N_14283,N_14180);
nand U21940 (N_21940,N_19474,N_14447);
nand U21941 (N_21941,N_18334,N_12717);
xnor U21942 (N_21942,N_19238,N_17217);
and U21943 (N_21943,N_10674,N_19116);
nand U21944 (N_21944,N_15104,N_19592);
nor U21945 (N_21945,N_15264,N_18475);
nand U21946 (N_21946,N_10638,N_14604);
nand U21947 (N_21947,N_14071,N_12843);
and U21948 (N_21948,N_11064,N_10511);
nor U21949 (N_21949,N_19492,N_16134);
nor U21950 (N_21950,N_12761,N_11968);
nand U21951 (N_21951,N_18717,N_12440);
and U21952 (N_21952,N_13378,N_19081);
nand U21953 (N_21953,N_11187,N_10822);
and U21954 (N_21954,N_14241,N_17303);
or U21955 (N_21955,N_11647,N_14663);
nand U21956 (N_21956,N_14154,N_13803);
nand U21957 (N_21957,N_16321,N_15905);
or U21958 (N_21958,N_12081,N_16778);
nor U21959 (N_21959,N_13275,N_16309);
and U21960 (N_21960,N_17299,N_16246);
nand U21961 (N_21961,N_18721,N_11198);
xor U21962 (N_21962,N_13817,N_18747);
or U21963 (N_21963,N_12705,N_16872);
and U21964 (N_21964,N_14637,N_18689);
nand U21965 (N_21965,N_14879,N_12874);
nand U21966 (N_21966,N_14043,N_19486);
nand U21967 (N_21967,N_18727,N_17567);
or U21968 (N_21968,N_16981,N_15988);
nand U21969 (N_21969,N_11634,N_12954);
xor U21970 (N_21970,N_17851,N_10736);
and U21971 (N_21971,N_10571,N_14670);
xor U21972 (N_21972,N_18345,N_12304);
and U21973 (N_21973,N_18620,N_17968);
nand U21974 (N_21974,N_12395,N_14906);
or U21975 (N_21975,N_11192,N_16854);
or U21976 (N_21976,N_14418,N_15372);
xor U21977 (N_21977,N_19566,N_15452);
nor U21978 (N_21978,N_10943,N_18147);
and U21979 (N_21979,N_18910,N_14758);
nand U21980 (N_21980,N_13317,N_13010);
and U21981 (N_21981,N_11713,N_14174);
nand U21982 (N_21982,N_18286,N_15008);
nand U21983 (N_21983,N_14693,N_14555);
or U21984 (N_21984,N_14194,N_15708);
xor U21985 (N_21985,N_11720,N_17931);
nand U21986 (N_21986,N_19575,N_19068);
nor U21987 (N_21987,N_14794,N_18895);
xnor U21988 (N_21988,N_14299,N_14370);
or U21989 (N_21989,N_17364,N_15084);
xnor U21990 (N_21990,N_12263,N_12738);
nand U21991 (N_21991,N_18355,N_17679);
nand U21992 (N_21992,N_17541,N_18698);
nor U21993 (N_21993,N_10523,N_14399);
nand U21994 (N_21994,N_17685,N_16963);
nor U21995 (N_21995,N_12004,N_11336);
nand U21996 (N_21996,N_10022,N_11549);
and U21997 (N_21997,N_15245,N_15014);
nor U21998 (N_21998,N_11018,N_12297);
nand U21999 (N_21999,N_11991,N_16098);
or U22000 (N_22000,N_15315,N_12914);
and U22001 (N_22001,N_10435,N_12123);
or U22002 (N_22002,N_11269,N_14435);
xor U22003 (N_22003,N_10806,N_13602);
nor U22004 (N_22004,N_11267,N_12529);
xor U22005 (N_22005,N_16262,N_16116);
nand U22006 (N_22006,N_10889,N_17575);
or U22007 (N_22007,N_13683,N_16370);
or U22008 (N_22008,N_19786,N_15462);
nand U22009 (N_22009,N_14729,N_13902);
or U22010 (N_22010,N_10236,N_16352);
nor U22011 (N_22011,N_15388,N_13350);
or U22012 (N_22012,N_12882,N_13823);
and U22013 (N_22013,N_17023,N_19029);
nand U22014 (N_22014,N_13666,N_17896);
and U22015 (N_22015,N_12532,N_13182);
nor U22016 (N_22016,N_14966,N_19793);
nor U22017 (N_22017,N_11343,N_19013);
or U22018 (N_22018,N_17382,N_15527);
xor U22019 (N_22019,N_19802,N_16339);
nor U22020 (N_22020,N_17117,N_12169);
nor U22021 (N_22021,N_13908,N_14193);
or U22022 (N_22022,N_17175,N_14830);
and U22023 (N_22023,N_16393,N_17016);
and U22024 (N_22024,N_13790,N_18247);
nand U22025 (N_22025,N_11231,N_13980);
or U22026 (N_22026,N_18858,N_18304);
or U22027 (N_22027,N_10254,N_16224);
or U22028 (N_22028,N_11314,N_19534);
nor U22029 (N_22029,N_19242,N_12164);
nor U22030 (N_22030,N_18290,N_18751);
or U22031 (N_22031,N_16868,N_10970);
or U22032 (N_22032,N_15918,N_15094);
nor U22033 (N_22033,N_12668,N_15891);
nand U22034 (N_22034,N_10849,N_18655);
nor U22035 (N_22035,N_16261,N_10145);
or U22036 (N_22036,N_14091,N_13034);
xor U22037 (N_22037,N_18954,N_19435);
nand U22038 (N_22038,N_17195,N_18595);
or U22039 (N_22039,N_18601,N_19113);
xor U22040 (N_22040,N_15569,N_12986);
nand U22041 (N_22041,N_19423,N_14680);
and U22042 (N_22042,N_14014,N_19909);
nand U22043 (N_22043,N_13278,N_19883);
nand U22044 (N_22044,N_18146,N_15307);
and U22045 (N_22045,N_17485,N_16193);
or U22046 (N_22046,N_13235,N_15700);
or U22047 (N_22047,N_12027,N_12261);
xnor U22048 (N_22048,N_19978,N_11684);
and U22049 (N_22049,N_14918,N_17098);
and U22050 (N_22050,N_14946,N_12219);
nand U22051 (N_22051,N_15325,N_14881);
xnor U22052 (N_22052,N_15752,N_14935);
or U22053 (N_22053,N_11029,N_12900);
nor U22054 (N_22054,N_11423,N_14051);
or U22055 (N_22055,N_16249,N_12634);
or U22056 (N_22056,N_19512,N_16347);
nand U22057 (N_22057,N_14324,N_18371);
nor U22058 (N_22058,N_14401,N_18732);
or U22059 (N_22059,N_15013,N_12567);
xnor U22060 (N_22060,N_10801,N_13253);
or U22061 (N_22061,N_19484,N_15380);
and U22062 (N_22062,N_18868,N_19480);
and U22063 (N_22063,N_18865,N_13608);
nor U22064 (N_22064,N_15191,N_10456);
nand U22065 (N_22065,N_19680,N_10834);
nand U22066 (N_22066,N_14790,N_15080);
or U22067 (N_22067,N_11301,N_19556);
xnor U22068 (N_22068,N_14527,N_11216);
nand U22069 (N_22069,N_12850,N_15445);
nor U22070 (N_22070,N_16876,N_14397);
nor U22071 (N_22071,N_11895,N_19003);
nand U22072 (N_22072,N_15291,N_17658);
nand U22073 (N_22073,N_15098,N_18339);
nor U22074 (N_22074,N_16349,N_10146);
or U22075 (N_22075,N_16493,N_17533);
nor U22076 (N_22076,N_12460,N_11014);
nand U22077 (N_22077,N_13981,N_11332);
or U22078 (N_22078,N_12310,N_11636);
or U22079 (N_22079,N_18714,N_14383);
nand U22080 (N_22080,N_13660,N_15103);
nand U22081 (N_22081,N_18303,N_19681);
xor U22082 (N_22082,N_14951,N_13838);
and U22083 (N_22083,N_15095,N_19122);
and U22084 (N_22084,N_11165,N_14708);
or U22085 (N_22085,N_11841,N_10020);
nor U22086 (N_22086,N_17820,N_15323);
nand U22087 (N_22087,N_14374,N_19885);
nand U22088 (N_22088,N_18805,N_11008);
xor U22089 (N_22089,N_17938,N_16204);
nor U22090 (N_22090,N_14207,N_16010);
nor U22091 (N_22091,N_16365,N_19859);
xnor U22092 (N_22092,N_18946,N_17285);
nor U22093 (N_22093,N_15651,N_15658);
nor U22094 (N_22094,N_15240,N_17088);
nor U22095 (N_22095,N_15192,N_16669);
nand U22096 (N_22096,N_10941,N_12582);
or U22097 (N_22097,N_18490,N_10922);
nand U22098 (N_22098,N_12371,N_18025);
nor U22099 (N_22099,N_17253,N_18522);
or U22100 (N_22100,N_15354,N_16189);
or U22101 (N_22101,N_15129,N_19688);
nor U22102 (N_22102,N_18327,N_10371);
and U22103 (N_22103,N_13741,N_17815);
and U22104 (N_22104,N_18155,N_13385);
and U22105 (N_22105,N_11184,N_19842);
nand U22106 (N_22106,N_11994,N_10668);
and U22107 (N_22107,N_16683,N_19928);
or U22108 (N_22108,N_16613,N_15050);
and U22109 (N_22109,N_13176,N_13099);
nor U22110 (N_22110,N_17899,N_16356);
nand U22111 (N_22111,N_16208,N_14534);
nor U22112 (N_22112,N_10835,N_11471);
xor U22113 (N_22113,N_15333,N_16069);
and U22114 (N_22114,N_14834,N_19951);
xor U22115 (N_22115,N_11561,N_10263);
xor U22116 (N_22116,N_13109,N_16758);
and U22117 (N_22117,N_12763,N_14046);
nand U22118 (N_22118,N_13641,N_15901);
xnor U22119 (N_22119,N_13087,N_14175);
and U22120 (N_22120,N_11431,N_14962);
nor U22121 (N_22121,N_14236,N_13059);
nand U22122 (N_22122,N_12210,N_14588);
xnor U22123 (N_22123,N_13521,N_18167);
nor U22124 (N_22124,N_15134,N_17147);
nor U22125 (N_22125,N_18034,N_18607);
nor U22126 (N_22126,N_15224,N_11691);
or U22127 (N_22127,N_18598,N_11633);
and U22128 (N_22128,N_12489,N_17792);
nor U22129 (N_22129,N_19107,N_10662);
or U22130 (N_22130,N_14390,N_12410);
xnor U22131 (N_22131,N_15924,N_11296);
and U22132 (N_22132,N_12121,N_11452);
and U22133 (N_22133,N_13547,N_12446);
nand U22134 (N_22134,N_16432,N_15075);
nor U22135 (N_22135,N_15162,N_11655);
nand U22136 (N_22136,N_10454,N_12387);
or U22137 (N_22137,N_13229,N_12844);
or U22138 (N_22138,N_19247,N_13701);
xnor U22139 (N_22139,N_14269,N_19321);
or U22140 (N_22140,N_14571,N_17154);
nand U22141 (N_22141,N_18298,N_16403);
and U22142 (N_22142,N_19542,N_16572);
nand U22143 (N_22143,N_18666,N_11354);
or U22144 (N_22144,N_12098,N_14594);
or U22145 (N_22145,N_18330,N_16491);
and U22146 (N_22146,N_11315,N_10042);
nor U22147 (N_22147,N_13722,N_17999);
nand U22148 (N_22148,N_14266,N_13610);
and U22149 (N_22149,N_16618,N_12731);
nor U22150 (N_22150,N_19005,N_14365);
nor U22151 (N_22151,N_16922,N_14939);
and U22152 (N_22152,N_11905,N_19364);
or U22153 (N_22153,N_11049,N_19612);
nand U22154 (N_22154,N_12826,N_18800);
or U22155 (N_22155,N_13647,N_19260);
nor U22156 (N_22156,N_14823,N_12800);
or U22157 (N_22157,N_18437,N_15346);
nor U22158 (N_22158,N_13659,N_16873);
nand U22159 (N_22159,N_10108,N_16444);
nand U22160 (N_22160,N_10138,N_12250);
or U22161 (N_22161,N_17911,N_15250);
and U22162 (N_22162,N_19852,N_10401);
or U22163 (N_22163,N_17618,N_18235);
and U22164 (N_22164,N_14739,N_14055);
and U22165 (N_22165,N_10094,N_15461);
or U22166 (N_22166,N_10842,N_17570);
and U22167 (N_22167,N_13836,N_19217);
nand U22168 (N_22168,N_13143,N_15268);
xnor U22169 (N_22169,N_11382,N_14649);
nor U22170 (N_22170,N_15466,N_15751);
or U22171 (N_22171,N_17538,N_12341);
xnor U22172 (N_22172,N_14952,N_17992);
or U22173 (N_22173,N_18128,N_15698);
nand U22174 (N_22174,N_17687,N_18902);
nand U22175 (N_22175,N_18818,N_19593);
or U22176 (N_22176,N_19422,N_15894);
or U22177 (N_22177,N_13679,N_11608);
and U22178 (N_22178,N_13298,N_14618);
xnor U22179 (N_22179,N_16589,N_19352);
nor U22180 (N_22180,N_11506,N_14228);
or U22181 (N_22181,N_17887,N_12784);
nor U22182 (N_22182,N_16506,N_14610);
nor U22183 (N_22183,N_17855,N_18170);
nor U22184 (N_22184,N_13390,N_11398);
and U22185 (N_22185,N_16324,N_10646);
nor U22186 (N_22186,N_16499,N_11870);
nand U22187 (N_22187,N_16059,N_11659);
xor U22188 (N_22188,N_18734,N_14357);
nor U22189 (N_22189,N_12314,N_11600);
xor U22190 (N_22190,N_11605,N_14087);
or U22191 (N_22191,N_15788,N_10374);
nand U22192 (N_22192,N_12566,N_11201);
nand U22193 (N_22193,N_10281,N_11135);
nand U22194 (N_22194,N_18415,N_11848);
and U22195 (N_22195,N_16412,N_16205);
nand U22196 (N_22196,N_12526,N_11538);
nand U22197 (N_22197,N_15934,N_14393);
or U22198 (N_22198,N_14652,N_15953);
nand U22199 (N_22199,N_12043,N_11500);
nand U22200 (N_22200,N_19677,N_18635);
nor U22201 (N_22201,N_11280,N_19042);
and U22202 (N_22202,N_16226,N_13342);
nand U22203 (N_22203,N_15862,N_11725);
and U22204 (N_22204,N_17084,N_12985);
and U22205 (N_22205,N_16931,N_14083);
xor U22206 (N_22206,N_17869,N_14414);
nor U22207 (N_22207,N_12401,N_17395);
and U22208 (N_22208,N_10305,N_13280);
xor U22209 (N_22209,N_17596,N_13672);
nor U22210 (N_22210,N_13334,N_12394);
nor U22211 (N_22211,N_16229,N_17691);
nor U22212 (N_22212,N_18433,N_11940);
and U22213 (N_22213,N_16953,N_14436);
or U22214 (N_22214,N_17403,N_16775);
or U22215 (N_22215,N_17145,N_19330);
or U22216 (N_22216,N_15812,N_11891);
and U22217 (N_22217,N_15801,N_17885);
nand U22218 (N_22218,N_11030,N_17381);
and U22219 (N_22219,N_19829,N_19397);
and U22220 (N_22220,N_10598,N_17027);
or U22221 (N_22221,N_11409,N_16236);
nand U22222 (N_22222,N_16737,N_15367);
nor U22223 (N_22223,N_13156,N_18310);
nand U22224 (N_22224,N_16689,N_19860);
nand U22225 (N_22225,N_15719,N_13338);
xor U22226 (N_22226,N_13685,N_15364);
xnor U22227 (N_22227,N_16247,N_10024);
nor U22228 (N_22228,N_15761,N_15037);
or U22229 (N_22229,N_15369,N_19969);
nand U22230 (N_22230,N_17130,N_17214);
or U22231 (N_22231,N_11539,N_15395);
and U22232 (N_22232,N_14892,N_19351);
and U22233 (N_22233,N_17221,N_14453);
nor U22234 (N_22234,N_12956,N_13178);
xnor U22235 (N_22235,N_11712,N_11874);
nor U22236 (N_22236,N_18488,N_12102);
xnor U22237 (N_22237,N_14439,N_12803);
or U22238 (N_22238,N_19669,N_15116);
or U22239 (N_22239,N_12796,N_17232);
xnor U22240 (N_22240,N_17004,N_19945);
and U22241 (N_22241,N_17432,N_11234);
nand U22242 (N_22242,N_17620,N_14692);
nor U22243 (N_22243,N_14955,N_10007);
nand U22244 (N_22244,N_16287,N_13209);
nor U22245 (N_22245,N_14683,N_17978);
nor U22246 (N_22246,N_14648,N_18783);
or U22247 (N_22247,N_17120,N_14698);
and U22248 (N_22248,N_13800,N_18082);
nand U22249 (N_22249,N_16837,N_19475);
and U22250 (N_22250,N_17225,N_14810);
nor U22251 (N_22251,N_13373,N_14490);
or U22252 (N_22252,N_19269,N_17599);
and U22253 (N_22253,N_19922,N_14669);
or U22254 (N_22254,N_10768,N_14573);
nand U22255 (N_22255,N_13690,N_10031);
and U22256 (N_22256,N_15859,N_14584);
nor U22257 (N_22257,N_19590,N_10927);
or U22258 (N_22258,N_18862,N_15121);
nand U22259 (N_22259,N_12650,N_12323);
nor U22260 (N_22260,N_15458,N_14570);
and U22261 (N_22261,N_13365,N_10150);
nand U22262 (N_22262,N_13606,N_17819);
and U22263 (N_22263,N_16241,N_11322);
nand U22264 (N_22264,N_13113,N_11088);
or U22265 (N_22265,N_12864,N_13847);
nand U22266 (N_22266,N_13462,N_15681);
or U22267 (N_22267,N_18825,N_19165);
nor U22268 (N_22268,N_13431,N_19340);
and U22269 (N_22269,N_15996,N_11992);
or U22270 (N_22270,N_19021,N_17363);
or U22271 (N_22271,N_18890,N_15710);
and U22272 (N_22272,N_15679,N_12228);
xnor U22273 (N_22273,N_13622,N_15888);
nor U22274 (N_22274,N_17706,N_19297);
or U22275 (N_22275,N_17798,N_15038);
and U22276 (N_22276,N_13821,N_11478);
and U22277 (N_22277,N_14275,N_11762);
nor U22278 (N_22278,N_19208,N_13205);
and U22279 (N_22279,N_12506,N_14262);
or U22280 (N_22280,N_11844,N_17467);
or U22281 (N_22281,N_14726,N_13161);
or U22282 (N_22282,N_11309,N_10891);
xor U22283 (N_22283,N_12486,N_11466);
or U22284 (N_22284,N_18794,N_16983);
nand U22285 (N_22285,N_19258,N_11660);
nand U22286 (N_22286,N_16906,N_15007);
xnor U22287 (N_22287,N_19718,N_11328);
xnor U22288 (N_22288,N_19790,N_16869);
xnor U22289 (N_22289,N_17179,N_17960);
and U22290 (N_22290,N_17847,N_13321);
and U22291 (N_22291,N_14142,N_10074);
or U22292 (N_22292,N_12347,N_19441);
nand U22293 (N_22293,N_19825,N_14472);
and U22294 (N_22294,N_12665,N_19879);
and U22295 (N_22295,N_19477,N_18104);
and U22296 (N_22296,N_11845,N_18190);
or U22297 (N_22297,N_10971,N_15152);
nor U22298 (N_22298,N_14837,N_14780);
and U22299 (N_22299,N_18801,N_13408);
nor U22300 (N_22300,N_16516,N_19989);
and U22301 (N_22301,N_14067,N_12296);
nand U22302 (N_22302,N_11693,N_18476);
nand U22303 (N_22303,N_13891,N_11418);
and U22304 (N_22304,N_16853,N_19193);
or U22305 (N_22305,N_11528,N_18927);
and U22306 (N_22306,N_15882,N_18342);
and U22307 (N_22307,N_10291,N_10364);
and U22308 (N_22308,N_15077,N_18999);
nand U22309 (N_22309,N_17073,N_14502);
nand U22310 (N_22310,N_16653,N_17610);
and U22311 (N_22311,N_12982,N_10584);
and U22312 (N_22312,N_15950,N_13778);
or U22313 (N_22313,N_15850,N_10795);
and U22314 (N_22314,N_17481,N_14034);
nand U22315 (N_22315,N_13655,N_19869);
nor U22316 (N_22316,N_16520,N_14542);
xnor U22317 (N_22317,N_18985,N_13193);
or U22318 (N_22318,N_18009,N_13056);
or U22319 (N_22319,N_18441,N_15661);
or U22320 (N_22320,N_17954,N_12846);
and U22321 (N_22321,N_16668,N_16334);
nor U22322 (N_22322,N_16942,N_12205);
nand U22323 (N_22323,N_10218,N_10707);
or U22324 (N_22324,N_10372,N_13058);
nand U22325 (N_22325,N_13310,N_14773);
and U22326 (N_22326,N_16700,N_12331);
xor U22327 (N_22327,N_11374,N_13396);
nor U22328 (N_22328,N_11361,N_12944);
or U22329 (N_22329,N_11179,N_19987);
nor U22330 (N_22330,N_11220,N_13469);
nor U22331 (N_22331,N_11070,N_18344);
and U22332 (N_22332,N_15057,N_17884);
nor U22333 (N_22333,N_11697,N_12499);
nor U22334 (N_22334,N_10349,N_16470);
and U22335 (N_22335,N_10921,N_15204);
nor U22336 (N_22336,N_10201,N_16280);
or U22337 (N_22337,N_12642,N_18537);
xor U22338 (N_22338,N_15189,N_10107);
and U22339 (N_22339,N_19641,N_12201);
or U22340 (N_22340,N_18849,N_18260);
nor U22341 (N_22341,N_10862,N_13170);
nand U22342 (N_22342,N_10117,N_17944);
and U22343 (N_22343,N_11807,N_15779);
or U22344 (N_22344,N_15871,N_12825);
and U22345 (N_22345,N_14238,N_14446);
or U22346 (N_22346,N_10936,N_15020);
or U22347 (N_22347,N_15327,N_13381);
nor U22348 (N_22348,N_18705,N_14633);
nand U22349 (N_22349,N_10044,N_17659);
nor U22350 (N_22350,N_14386,N_15533);
nand U22351 (N_22351,N_12557,N_14989);
or U22352 (N_22352,N_14050,N_16657);
nor U22353 (N_22353,N_15415,N_10248);
nand U22354 (N_22354,N_14500,N_17573);
nor U22355 (N_22355,N_13992,N_18641);
xor U22356 (N_22356,N_15860,N_19365);
and U22357 (N_22357,N_17422,N_15802);
nor U22358 (N_22358,N_14268,N_15298);
and U22359 (N_22359,N_19020,N_17811);
nor U22360 (N_22360,N_10959,N_14724);
nor U22361 (N_22361,N_11974,N_10178);
nor U22362 (N_22362,N_14037,N_11188);
nand U22363 (N_22363,N_16644,N_19606);
or U22364 (N_22364,N_18217,N_10175);
nand U22365 (N_22365,N_14459,N_16783);
or U22366 (N_22366,N_19996,N_18016);
or U22367 (N_22367,N_14791,N_16566);
nand U22368 (N_22368,N_14789,N_14863);
nor U22369 (N_22369,N_15234,N_16446);
nand U22370 (N_22370,N_16734,N_15212);
and U22371 (N_22371,N_14623,N_17236);
or U22372 (N_22372,N_17149,N_14821);
and U22373 (N_22373,N_15235,N_15975);
and U22374 (N_22374,N_15440,N_13251);
and U22375 (N_22375,N_10347,N_17510);
or U22376 (N_22376,N_12981,N_16633);
nor U22377 (N_22377,N_17729,N_19794);
and U22378 (N_22378,N_13409,N_19699);
nor U22379 (N_22379,N_10383,N_15516);
or U22380 (N_22380,N_17359,N_11069);
and U22381 (N_22381,N_15829,N_12495);
nor U22382 (N_22382,N_15487,N_13941);
nor U22383 (N_22383,N_10220,N_11699);
or U22384 (N_22384,N_11129,N_10546);
or U22385 (N_22385,N_16709,N_17037);
nand U22386 (N_22386,N_14345,N_12698);
or U22387 (N_22387,N_14409,N_16426);
nor U22388 (N_22388,N_14753,N_15680);
nand U22389 (N_22389,N_18125,N_12925);
or U22390 (N_22390,N_11062,N_11162);
xor U22391 (N_22391,N_10215,N_18894);
nor U22392 (N_22392,N_11019,N_18811);
xor U22393 (N_22393,N_12322,N_14127);
nand U22394 (N_22394,N_12178,N_11371);
and U22395 (N_22395,N_11147,N_14063);
nand U22396 (N_22396,N_13750,N_15831);
and U22397 (N_22397,N_16538,N_10726);
nor U22398 (N_22398,N_12624,N_14949);
nand U22399 (N_22399,N_15830,N_10649);
and U22400 (N_22400,N_11951,N_15717);
and U22401 (N_22401,N_17013,N_11424);
or U22402 (N_22402,N_18559,N_19964);
nor U22403 (N_22403,N_18682,N_16285);
nand U22404 (N_22404,N_14229,N_16896);
or U22405 (N_22405,N_17164,N_19926);
xor U22406 (N_22406,N_14066,N_10095);
and U22407 (N_22407,N_16675,N_19197);
nand U22408 (N_22408,N_19227,N_11141);
and U22409 (N_22409,N_13145,N_14130);
nor U22410 (N_22410,N_18648,N_14188);
xor U22411 (N_22411,N_13609,N_15514);
nand U22412 (N_22412,N_10816,N_10026);
nand U22413 (N_22413,N_18570,N_15931);
and U22414 (N_22414,N_11227,N_10693);
and U22415 (N_22415,N_16615,N_15167);
and U22416 (N_22416,N_13732,N_16045);
nand U22417 (N_22417,N_15711,N_12775);
nor U22418 (N_22418,N_19890,N_17513);
or U22419 (N_22419,N_11767,N_12607);
and U22420 (N_22420,N_15754,N_18645);
nor U22421 (N_22421,N_13424,N_19618);
or U22422 (N_22422,N_16216,N_13148);
xnor U22423 (N_22423,N_18255,N_19585);
xor U22424 (N_22424,N_11031,N_10890);
nand U22425 (N_22425,N_13042,N_12907);
xor U22426 (N_22426,N_13773,N_16518);
nor U22427 (N_22427,N_12892,N_15961);
and U22428 (N_22428,N_14190,N_18758);
nor U22429 (N_22429,N_19913,N_15119);
nor U22430 (N_22430,N_17208,N_15781);
or U22431 (N_22431,N_19212,N_10914);
nand U22432 (N_22432,N_17828,N_15632);
nand U22433 (N_22433,N_17925,N_11421);
or U22434 (N_22434,N_17963,N_11864);
or U22435 (N_22435,N_15519,N_18634);
and U22436 (N_22436,N_10745,N_14969);
or U22437 (N_22437,N_15740,N_19460);
or U22438 (N_22438,N_13454,N_14501);
nor U22439 (N_22439,N_13979,N_17228);
and U22440 (N_22440,N_15695,N_12555);
nor U22441 (N_22441,N_13520,N_13141);
nor U22442 (N_22442,N_17991,N_12188);
nand U22443 (N_22443,N_12443,N_10029);
nand U22444 (N_22444,N_13486,N_15024);
or U22445 (N_22445,N_15712,N_14272);
and U22446 (N_22446,N_14750,N_15018);
or U22447 (N_22447,N_15034,N_19065);
nor U22448 (N_22448,N_15565,N_14779);
nor U22449 (N_22449,N_15612,N_15723);
or U22450 (N_22450,N_10788,N_17393);
nor U22451 (N_22451,N_17598,N_14274);
nand U22452 (N_22452,N_17177,N_16770);
nand U22453 (N_22453,N_12008,N_12239);
nand U22454 (N_22454,N_12269,N_14441);
and U22455 (N_22455,N_15561,N_17304);
xnor U22456 (N_22456,N_15156,N_18280);
nor U22457 (N_22457,N_18301,N_10845);
nor U22458 (N_22458,N_16698,N_10592);
nand U22459 (N_22459,N_10853,N_19037);
and U22460 (N_22460,N_14314,N_13132);
xor U22461 (N_22461,N_17667,N_16710);
or U22462 (N_22462,N_18305,N_12917);
and U22463 (N_22463,N_14808,N_10810);
and U22464 (N_22464,N_17173,N_17583);
and U22465 (N_22465,N_11355,N_16335);
and U22466 (N_22466,N_11051,N_14237);
and U22467 (N_22467,N_10976,N_14448);
xnor U22468 (N_22468,N_18882,N_15821);
nand U22469 (N_22469,N_10578,N_17572);
or U22470 (N_22470,N_19275,N_15485);
nor U22471 (N_22471,N_13865,N_11485);
nor U22472 (N_22472,N_16776,N_12103);
and U22473 (N_22473,N_10324,N_10875);
nand U22474 (N_22474,N_17876,N_18109);
and U22475 (N_22475,N_12593,N_10993);
or U22476 (N_22476,N_11291,N_13190);
nor U22477 (N_22477,N_13072,N_19410);
nand U22478 (N_22478,N_12173,N_13765);
and U22479 (N_22479,N_12065,N_13988);
nand U22480 (N_22480,N_12757,N_15169);
and U22481 (N_22481,N_18372,N_15499);
and U22482 (N_22482,N_12815,N_17211);
nand U22483 (N_22483,N_14284,N_19341);
nor U22484 (N_22484,N_15302,N_18866);
or U22485 (N_22485,N_19840,N_14158);
nor U22486 (N_22486,N_17637,N_19048);
nor U22487 (N_22487,N_17150,N_12352);
and U22488 (N_22488,N_19323,N_19031);
and U22489 (N_22489,N_10614,N_10200);
nor U22490 (N_22490,N_16420,N_13617);
nor U22491 (N_22491,N_12857,N_16704);
or U22492 (N_22492,N_15532,N_13806);
or U22493 (N_22493,N_16966,N_18982);
nand U22494 (N_22494,N_11970,N_11013);
nor U22495 (N_22495,N_16975,N_17800);
or U22496 (N_22496,N_16528,N_10644);
and U22497 (N_22497,N_11711,N_19294);
or U22498 (N_22498,N_13523,N_15553);
nor U22499 (N_22499,N_12308,N_16786);
or U22500 (N_22500,N_17707,N_17958);
xor U22501 (N_22501,N_10332,N_11203);
and U22502 (N_22502,N_17950,N_17440);
nor U22503 (N_22503,N_14685,N_10612);
xnor U22504 (N_22504,N_12138,N_10682);
nor U22505 (N_22505,N_18411,N_10509);
or U22506 (N_22506,N_14388,N_13794);
nor U22507 (N_22507,N_13579,N_11106);
and U22508 (N_22508,N_14492,N_19355);
nand U22509 (N_22509,N_14984,N_17859);
or U22510 (N_22510,N_16222,N_17521);
nand U22511 (N_22511,N_18686,N_10096);
and U22512 (N_22512,N_17809,N_18291);
or U22513 (N_22513,N_17502,N_18354);
or U22514 (N_22514,N_19007,N_12202);
and U22515 (N_22515,N_10011,N_15338);
nor U22516 (N_22516,N_15469,N_18074);
xor U22517 (N_22517,N_19738,N_18729);
xnor U22518 (N_22518,N_19668,N_14270);
xor U22519 (N_22519,N_19241,N_13702);
xnor U22520 (N_22520,N_12824,N_10556);
nand U22521 (N_22521,N_10815,N_16794);
or U22522 (N_22522,N_15645,N_11439);
nand U22523 (N_22523,N_14715,N_18145);
nand U22524 (N_22524,N_13126,N_16083);
nor U22525 (N_22525,N_17605,N_11878);
and U22526 (N_22526,N_13459,N_12459);
or U22527 (N_22527,N_16888,N_10636);
xnor U22528 (N_22528,N_16337,N_17744);
and U22529 (N_22529,N_13673,N_12011);
nor U22530 (N_22530,N_18753,N_14047);
and U22531 (N_22531,N_10235,N_19834);
nor U22532 (N_22532,N_15072,N_10622);
nand U22533 (N_22533,N_14976,N_16614);
nand U22534 (N_22534,N_10742,N_12863);
nor U22535 (N_22535,N_17035,N_15312);
nor U22536 (N_22536,N_12180,N_15370);
or U22537 (N_22537,N_18459,N_10274);
xnor U22538 (N_22538,N_11330,N_15433);
or U22539 (N_22539,N_16488,N_13752);
xor U22540 (N_22540,N_12788,N_14827);
nand U22541 (N_22541,N_12617,N_17553);
xor U22542 (N_22542,N_15475,N_15742);
or U22543 (N_22543,N_11103,N_13881);
or U22544 (N_22544,N_19381,N_10373);
and U22545 (N_22545,N_10867,N_11510);
nor U22546 (N_22546,N_13119,N_11580);
or U22547 (N_22547,N_17977,N_11947);
and U22548 (N_22548,N_14118,N_17301);
nand U22549 (N_22549,N_18080,N_15339);
xor U22550 (N_22550,N_14772,N_14008);
nand U22551 (N_22551,N_17919,N_14137);
or U22552 (N_22552,N_18447,N_13120);
or U22553 (N_22553,N_10167,N_10955);
nand U22554 (N_22554,N_19772,N_14310);
nand U22555 (N_22555,N_15666,N_12080);
and U22556 (N_22556,N_12448,N_13101);
xnor U22557 (N_22557,N_16049,N_10147);
nor U22558 (N_22558,N_10265,N_16452);
nand U22559 (N_22559,N_13775,N_17497);
xor U22560 (N_22560,N_12466,N_17318);
xor U22561 (N_22561,N_12252,N_17895);
nor U22562 (N_22562,N_17550,N_13479);
xor U22563 (N_22563,N_12730,N_11253);
and U22564 (N_22564,N_16304,N_17712);
and U22565 (N_22565,N_15349,N_14546);
nor U22566 (N_22566,N_11803,N_13572);
nor U22567 (N_22567,N_13736,N_15767);
nand U22568 (N_22568,N_11446,N_18376);
nor U22569 (N_22569,N_17684,N_19372);
or U22570 (N_22570,N_17777,N_18740);
nand U22571 (N_22571,N_14836,N_10728);
nor U22572 (N_22572,N_16865,N_16514);
nand U22573 (N_22573,N_19906,N_15087);
xnor U22574 (N_22574,N_13700,N_11139);
nand U22575 (N_22575,N_16806,N_17669);
and U22576 (N_22576,N_15330,N_11256);
nand U22577 (N_22577,N_16297,N_10052);
nand U22578 (N_22578,N_18995,N_10769);
nand U22579 (N_22579,N_10658,N_18639);
and U22580 (N_22580,N_11334,N_13411);
nor U22581 (N_22581,N_18650,N_11183);
nand U22582 (N_22582,N_10389,N_10734);
or U22583 (N_22583,N_19288,N_11282);
nand U22584 (N_22584,N_14404,N_13045);
nand U22585 (N_22585,N_17491,N_14990);
nand U22586 (N_22586,N_16190,N_18443);
and U22587 (N_22587,N_12417,N_11884);
nor U22588 (N_22588,N_14815,N_12631);
nor U22589 (N_22589,N_10213,N_17836);
and U22590 (N_22590,N_18213,N_17975);
or U22591 (N_22591,N_11927,N_17280);
nand U22592 (N_22592,N_10413,N_19359);
xor U22593 (N_22593,N_10581,N_11568);
xor U22594 (N_22594,N_14626,N_13115);
nand U22595 (N_22595,N_18288,N_10877);
nand U22596 (N_22596,N_17582,N_17862);
nor U22597 (N_22597,N_16415,N_15545);
nor U22598 (N_22598,N_18843,N_13779);
or U22599 (N_22599,N_17347,N_16662);
xor U22600 (N_22600,N_11701,N_17973);
or U22601 (N_22601,N_19090,N_11750);
nand U22602 (N_22602,N_13723,N_18831);
nand U22603 (N_22603,N_13972,N_18059);
or U22604 (N_22604,N_12810,N_13435);
or U22605 (N_22605,N_18402,N_16851);
nand U22606 (N_22606,N_16954,N_18179);
nor U22607 (N_22607,N_13965,N_11525);
nor U22608 (N_22608,N_19762,N_14195);
or U22609 (N_22609,N_11050,N_13549);
nand U22610 (N_22610,N_17051,N_12282);
nor U22611 (N_22611,N_11706,N_10537);
nand U22612 (N_22612,N_18548,N_11728);
nor U22613 (N_22613,N_18408,N_17840);
nand U22614 (N_22614,N_19451,N_10047);
xnor U22615 (N_22615,N_18113,N_15627);
nor U22616 (N_22616,N_14265,N_14533);
or U22617 (N_22617,N_19034,N_12240);
xnor U22618 (N_22618,N_11810,N_10940);
nand U22619 (N_22619,N_10528,N_19218);
nand U22620 (N_22620,N_11612,N_12271);
or U22621 (N_22621,N_15481,N_12383);
nor U22622 (N_22622,N_18199,N_16886);
and U22623 (N_22623,N_17981,N_14543);
nand U22624 (N_22624,N_18821,N_19305);
and U22625 (N_22625,N_19290,N_19967);
or U22626 (N_22626,N_10680,N_17383);
and U22627 (N_22627,N_11504,N_13849);
xnor U22628 (N_22628,N_17093,N_14613);
nand U22629 (N_22629,N_15536,N_19429);
or U22630 (N_22630,N_19963,N_14445);
or U22631 (N_22631,N_15249,N_10270);
nor U22632 (N_22632,N_14305,N_10230);
nor U22633 (N_22633,N_19115,N_11181);
nand U22634 (N_22634,N_14995,N_19756);
and U22635 (N_22635,N_14364,N_18728);
nand U22636 (N_22636,N_11288,N_18480);
and U22637 (N_22637,N_14323,N_10192);
nor U22638 (N_22638,N_14707,N_17428);
or U22639 (N_22639,N_10290,N_11996);
nor U22640 (N_22640,N_16621,N_12660);
xor U22641 (N_22641,N_19712,N_10021);
nand U22642 (N_22642,N_11024,N_10677);
or U22643 (N_22643,N_11730,N_11120);
xor U22644 (N_22644,N_15175,N_12095);
nand U22645 (N_22645,N_11441,N_10199);
nand U22646 (N_22646,N_19099,N_11214);
or U22647 (N_22647,N_19299,N_12161);
xor U22648 (N_22648,N_10950,N_16340);
and U22649 (N_22649,N_11611,N_19792);
or U22650 (N_22650,N_10543,N_17376);
and U22651 (N_22651,N_18886,N_16753);
and U22652 (N_22652,N_15508,N_16713);
nand U22653 (N_22653,N_10071,N_11644);
nor U22654 (N_22654,N_10152,N_18949);
and U22655 (N_22655,N_19112,N_17834);
nand U22656 (N_22656,N_13135,N_10620);
nand U22657 (N_22657,N_16443,N_17021);
or U22658 (N_22658,N_12203,N_13852);
nand U22659 (N_22659,N_16658,N_12524);
nor U22660 (N_22660,N_12688,N_14112);
and U22661 (N_22661,N_13869,N_14917);
and U22662 (N_22662,N_15542,N_17454);
nand U22663 (N_22663,N_18904,N_18593);
and U22664 (N_22664,N_12396,N_15006);
xnor U22665 (N_22665,N_12646,N_16009);
xnor U22666 (N_22666,N_19623,N_19776);
xor U22667 (N_22667,N_15579,N_10261);
and U22668 (N_22668,N_19740,N_12496);
or U22669 (N_22669,N_17806,N_16718);
nor U22670 (N_22670,N_12719,N_19314);
or U22671 (N_22671,N_15409,N_19704);
nor U22672 (N_22672,N_16430,N_15507);
nor U22673 (N_22673,N_18254,N_10942);
nand U22674 (N_22674,N_10908,N_11093);
nor U22675 (N_22675,N_16018,N_17019);
nor U22676 (N_22676,N_15867,N_12777);
nor U22677 (N_22677,N_13899,N_14979);
xnor U22678 (N_22678,N_17315,N_11221);
and U22679 (N_22679,N_11458,N_15196);
nand U22680 (N_22680,N_15363,N_10902);
nand U22681 (N_22681,N_10196,N_17047);
nand U22682 (N_22682,N_18063,N_16409);
nand U22683 (N_22683,N_10749,N_12613);
nor U22684 (N_22684,N_16177,N_13061);
and U22685 (N_22685,N_14149,N_19643);
and U22686 (N_22686,N_16417,N_12990);
nand U22687 (N_22687,N_11279,N_12888);
or U22688 (N_22688,N_13747,N_19076);
nor U22689 (N_22689,N_14592,N_14352);
or U22690 (N_22690,N_14516,N_17748);
xnor U22691 (N_22691,N_15335,N_13347);
nand U22692 (N_22692,N_13309,N_14875);
or U22693 (N_22693,N_16605,N_17444);
xor U22694 (N_22694,N_11559,N_18780);
and U22695 (N_22695,N_12749,N_13818);
or U22696 (N_22696,N_12069,N_11536);
and U22697 (N_22697,N_11092,N_19961);
and U22698 (N_22698,N_19419,N_15983);
xor U22699 (N_22699,N_19490,N_13292);
nand U22700 (N_22700,N_16883,N_15940);
nor U22701 (N_22701,N_11872,N_18497);
or U22702 (N_22702,N_11919,N_15005);
and U22703 (N_22703,N_16809,N_16140);
and U22704 (N_22704,N_19920,N_10040);
or U22705 (N_22705,N_16081,N_14148);
nand U22706 (N_22706,N_12348,N_19498);
nor U22707 (N_22707,N_13203,N_12032);
and U22708 (N_22708,N_13805,N_15952);
xnor U22709 (N_22709,N_11480,N_11469);
or U22710 (N_22710,N_11998,N_17568);
nor U22711 (N_22711,N_13077,N_16988);
or U22712 (N_22712,N_17839,N_12976);
and U22713 (N_22713,N_12412,N_17103);
nor U22714 (N_22714,N_10854,N_18977);
nand U22715 (N_22715,N_15990,N_15340);
xnor U22716 (N_22716,N_16020,N_14264);
or U22717 (N_22717,N_16800,N_13841);
or U22718 (N_22718,N_11071,N_17779);
and U22719 (N_22719,N_15942,N_10541);
nand U22720 (N_22720,N_17914,N_12303);
and U22721 (N_22721,N_18633,N_12044);
xnor U22722 (N_22722,N_10549,N_17137);
and U22723 (N_22723,N_10458,N_18690);
and U22724 (N_22724,N_19485,N_15071);
or U22725 (N_22725,N_19866,N_13037);
or U22726 (N_22726,N_17544,N_15641);
or U22727 (N_22727,N_10805,N_13526);
nand U22728 (N_22728,N_15443,N_10743);
and U22729 (N_22729,N_14398,N_15872);
nand U22730 (N_22730,N_15954,N_19625);
nor U22731 (N_22731,N_15453,N_11662);
xor U22732 (N_22732,N_15895,N_13893);
nor U22733 (N_22733,N_11131,N_11553);
nand U22734 (N_22734,N_17638,N_19946);
and U22735 (N_22735,N_13599,N_18257);
or U22736 (N_22736,N_18195,N_12786);
xor U22737 (N_22737,N_10740,N_11880);
xnor U22738 (N_22738,N_16838,N_15269);
and U22739 (N_22739,N_16014,N_13057);
or U22740 (N_22740,N_18030,N_19311);
xor U22741 (N_22741,N_18137,N_13964);
nand U22742 (N_22742,N_15827,N_18070);
xor U22743 (N_22743,N_18205,N_10500);
and U22744 (N_22744,N_12411,N_10878);
and U22745 (N_22745,N_14638,N_18196);
nor U22746 (N_22746,N_17473,N_18931);
xnor U22747 (N_22747,N_12877,N_18958);
and U22748 (N_22748,N_12033,N_11657);
nor U22749 (N_22749,N_15465,N_15689);
nor U22750 (N_22750,N_17934,N_14026);
or U22751 (N_22751,N_11157,N_13443);
nor U22752 (N_22752,N_10320,N_19342);
nor U22753 (N_22753,N_10319,N_11721);
xor U22754 (N_22754,N_14465,N_16972);
nor U22755 (N_22755,N_11993,N_16169);
nand U22756 (N_22756,N_11597,N_12291);
nor U22757 (N_22757,N_10575,N_15836);
nor U22758 (N_22758,N_15758,N_15124);
nand U22759 (N_22759,N_15412,N_18347);
and U22760 (N_22760,N_11832,N_11206);
or U22761 (N_22761,N_11727,N_16485);
nand U22762 (N_22762,N_15760,N_19522);
nand U22763 (N_22763,N_17305,N_12685);
nand U22764 (N_22764,N_14817,N_14092);
or U22765 (N_22765,N_19293,N_16072);
and U22766 (N_22766,N_17829,N_10732);
xnor U22767 (N_22767,N_11036,N_16763);
nor U22768 (N_22768,N_17446,N_11886);
nand U22769 (N_22769,N_17760,N_10667);
nor U22770 (N_22770,N_16768,N_16542);
and U22771 (N_22771,N_10206,N_15253);
or U22772 (N_22772,N_18737,N_13632);
xor U22773 (N_22773,N_14328,N_16874);
nor U22774 (N_22774,N_13748,N_14619);
nand U22775 (N_22775,N_18835,N_13412);
nand U22776 (N_22776,N_15825,N_13324);
and U22777 (N_22777,N_17560,N_16831);
nand U22778 (N_22778,N_15568,N_18095);
or U22779 (N_22779,N_12266,N_16788);
nor U22780 (N_22780,N_19343,N_14621);
and U22781 (N_22781,N_10992,N_12047);
and U22782 (N_22782,N_14062,N_15762);
nand U22783 (N_22783,N_17614,N_17827);
nand U22784 (N_22784,N_18422,N_14840);
or U22785 (N_22785,N_15099,N_19658);
nor U22786 (N_22786,N_19604,N_13706);
xor U22787 (N_22787,N_19767,N_13663);
xnor U22788 (N_22788,N_11989,N_11205);
xor U22789 (N_22789,N_15624,N_13364);
or U22790 (N_22790,N_19861,N_13452);
or U22791 (N_22791,N_12523,N_14843);
nand U22792 (N_22792,N_11357,N_11521);
nand U22793 (N_22793,N_19876,N_18770);
nand U22794 (N_22794,N_15857,N_17260);
xnor U22795 (N_22795,N_18757,N_13265);
or U22796 (N_22796,N_12633,N_14593);
xnor U22797 (N_22797,N_14192,N_14909);
xor U22798 (N_22798,N_16388,N_19580);
or U22799 (N_22799,N_19296,N_15546);
nand U22800 (N_22800,N_16814,N_11360);
and U22801 (N_22801,N_18750,N_16026);
nor U22802 (N_22802,N_14169,N_17244);
and U22803 (N_22803,N_18746,N_16545);
nand U22804 (N_22804,N_17459,N_17482);
nor U22805 (N_22805,N_19570,N_10965);
and U22806 (N_22806,N_15520,N_14597);
and U22807 (N_22807,N_19664,N_15042);
nand U22808 (N_22808,N_14146,N_17274);
or U22809 (N_22809,N_12554,N_10724);
nand U22810 (N_22810,N_12217,N_16559);
nand U22811 (N_22811,N_18679,N_13343);
and U22812 (N_22812,N_13519,N_10244);
nand U22813 (N_22813,N_17089,N_15143);
nand U22814 (N_22814,N_17604,N_17001);
nor U22815 (N_22815,N_13307,N_17394);
and U22816 (N_22816,N_11095,N_13942);
nand U22817 (N_22817,N_18850,N_17293);
nand U22818 (N_22818,N_16771,N_15028);
nor U22819 (N_22819,N_15044,N_17645);
or U22820 (N_22820,N_17734,N_13033);
and U22821 (N_22821,N_18090,N_18589);
nor U22822 (N_22822,N_11604,N_13220);
xnor U22823 (N_22823,N_10323,N_13857);
or U22824 (N_22824,N_15619,N_11540);
or U22825 (N_22825,N_14040,N_12805);
and U22826 (N_22826,N_14396,N_15843);
nand U22827 (N_22827,N_18722,N_12507);
nor U22828 (N_22828,N_10438,N_11026);
and U22829 (N_22829,N_13369,N_18613);
nor U22830 (N_22830,N_19345,N_12061);
nand U22831 (N_22831,N_13993,N_11908);
nand U22832 (N_22832,N_11023,N_13425);
or U22833 (N_22833,N_16836,N_12120);
nor U22834 (N_22834,N_13293,N_18712);
and U22835 (N_22835,N_15980,N_12902);
xnor U22836 (N_22836,N_19472,N_11758);
nand U22837 (N_22837,N_16722,N_11487);
and U22838 (N_22838,N_15749,N_17986);
nand U22839 (N_22839,N_17492,N_18397);
and U22840 (N_22840,N_13642,N_10131);
nor U22841 (N_22841,N_13718,N_10689);
xnor U22842 (N_22842,N_16153,N_16773);
nand U22843 (N_22843,N_10513,N_18930);
nor U22844 (N_22844,N_18311,N_14211);
nand U22845 (N_22845,N_16882,N_15629);
nand U22846 (N_22846,N_15995,N_19985);
nor U22847 (N_22847,N_13341,N_17413);
and U22848 (N_22848,N_16889,N_11297);
and U22849 (N_22849,N_16744,N_18860);
nand U22850 (N_22850,N_14387,N_12847);
nand U22851 (N_22851,N_16320,N_11971);
nand U22852 (N_22852,N_15999,N_13651);
nand U22853 (N_22853,N_12199,N_19502);
nand U22854 (N_22854,N_18002,N_16248);
and U22855 (N_22855,N_10118,N_18516);
nor U22856 (N_22856,N_12051,N_14894);
nand U22857 (N_22857,N_14800,N_19053);
nor U22858 (N_22858,N_18076,N_18881);
nand U22859 (N_22859,N_17922,N_16510);
nand U22860 (N_22860,N_14598,N_10060);
nor U22861 (N_22861,N_17245,N_17341);
or U22862 (N_22862,N_17776,N_12318);
xnor U22863 (N_22863,N_16959,N_11289);
nor U22864 (N_22864,N_17486,N_17265);
or U22865 (N_22865,N_14515,N_15866);
nand U22866 (N_22866,N_18906,N_10871);
and U22867 (N_22867,N_18313,N_18381);
and U22868 (N_22868,N_10796,N_17142);
or U22869 (N_22869,N_13788,N_16255);
xnor U22870 (N_22870,N_12525,N_16086);
nor U22871 (N_22871,N_10903,N_18526);
or U22872 (N_22872,N_11321,N_19517);
or U22873 (N_22873,N_18178,N_17020);
and U22874 (N_22874,N_11193,N_10870);
nor U22875 (N_22875,N_16316,N_10756);
nand U22876 (N_22876,N_12113,N_12157);
nor U22877 (N_22877,N_17111,N_11196);
nand U22878 (N_22878,N_11042,N_12038);
nor U22879 (N_22879,N_10392,N_16735);
or U22880 (N_22880,N_19713,N_13053);
xor U22881 (N_22881,N_16513,N_18453);
and U22882 (N_22882,N_19814,N_10301);
or U22883 (N_22883,N_11964,N_17426);
and U22884 (N_22884,N_19176,N_18822);
or U22885 (N_22885,N_16647,N_11204);
or U22886 (N_22886,N_19722,N_17595);
and U22887 (N_22887,N_18524,N_15659);
nor U22888 (N_22888,N_11262,N_19880);
nor U22889 (N_22889,N_12866,N_19061);
nand U22890 (N_22890,N_12721,N_11812);
nor U22891 (N_22891,N_13814,N_18744);
nand U22892 (N_22892,N_17180,N_17455);
nand U22893 (N_22893,N_11575,N_16326);
nor U22894 (N_22894,N_12472,N_10793);
nor U22895 (N_22895,N_11901,N_19552);
nand U22896 (N_22896,N_14202,N_16109);
nor U22897 (N_22897,N_15777,N_15977);
and U22898 (N_22898,N_16891,N_16160);
nand U22899 (N_22899,N_11266,N_14019);
and U22900 (N_22900,N_19671,N_16547);
nor U22901 (N_22901,N_16861,N_19830);
nor U22902 (N_22902,N_14171,N_19795);
nand U22903 (N_22903,N_13382,N_12686);
nor U22904 (N_22904,N_19493,N_11306);
nor U22905 (N_22905,N_11717,N_14257);
nor U22906 (N_22906,N_18169,N_17998);
xnor U22907 (N_22907,N_19499,N_13286);
nor U22908 (N_22908,N_14678,N_15741);
nand U22909 (N_22909,N_19598,N_14131);
nor U22910 (N_22910,N_12663,N_17401);
nor U22911 (N_22911,N_10436,N_19676);
or U22912 (N_22912,N_14977,N_15773);
xnor U22913 (N_22913,N_14757,N_14901);
nor U22914 (N_22914,N_12148,N_19642);
or U22915 (N_22915,N_19886,N_15203);
nand U22916 (N_22916,N_14852,N_19416);
nand U22917 (N_22917,N_14049,N_13946);
and U22918 (N_22918,N_17817,N_13243);
xor U22919 (N_22919,N_13686,N_13418);
nand U22920 (N_22920,N_19319,N_13573);
or U22921 (N_22921,N_15120,N_12726);
and U22922 (N_22922,N_10188,N_13254);
nand U22923 (N_22923,N_17743,N_12183);
or U22924 (N_22924,N_19106,N_12062);
nor U22925 (N_22925,N_13951,N_15279);
xnor U22926 (N_22926,N_16253,N_16968);
or U22927 (N_22927,N_15280,N_12915);
or U22928 (N_22928,N_11656,N_10027);
nand U22929 (N_22929,N_15163,N_11765);
nand U22930 (N_22930,N_18941,N_16123);
nor U22931 (N_22931,N_18349,N_19586);
nand U22932 (N_22932,N_16477,N_11261);
nor U22933 (N_22933,N_19044,N_13944);
and U22934 (N_22934,N_12052,N_17566);
nor U22935 (N_22935,N_10577,N_18713);
xnor U22936 (N_22936,N_19421,N_13107);
xor U22937 (N_22937,N_12126,N_13384);
or U22938 (N_22938,N_12416,N_10702);
nand U22939 (N_22939,N_10613,N_18150);
nor U22940 (N_22940,N_19168,N_15803);
nand U22941 (N_22941,N_10823,N_15654);
or U22942 (N_22942,N_10195,N_16553);
or U22943 (N_22943,N_11952,N_17810);
nand U22944 (N_22944,N_18508,N_19600);
nor U22945 (N_22945,N_11066,N_19210);
nor U22946 (N_22946,N_13027,N_18812);
xnor U22947 (N_22947,N_19533,N_13835);
nor U22948 (N_22948,N_10228,N_14562);
and U22949 (N_22949,N_11174,N_10268);
nand U22950 (N_22950,N_18510,N_15497);
and U22951 (N_22951,N_17837,N_12672);
or U22952 (N_22952,N_18586,N_10475);
nor U22953 (N_22953,N_12195,N_17767);
nor U22954 (N_22954,N_15251,N_10017);
xor U22955 (N_22955,N_18704,N_19891);
nor U22956 (N_22956,N_11130,N_13815);
and U22957 (N_22957,N_10451,N_17268);
nor U22958 (N_22958,N_17780,N_10422);
nand U22959 (N_22959,N_10625,N_10770);
nand U22960 (N_22960,N_12991,N_10141);
or U22961 (N_22961,N_19620,N_15928);
nor U22962 (N_22962,N_16808,N_18265);
nand U22963 (N_22963,N_11109,N_17324);
or U22964 (N_22964,N_19748,N_18175);
nor U22965 (N_22965,N_10911,N_16939);
nand U22966 (N_22966,N_13196,N_11033);
or U22967 (N_22967,N_14389,N_19907);
nor U22968 (N_22968,N_18514,N_10641);
nor U22969 (N_22969,N_19974,N_18694);
nand U22970 (N_22970,N_18926,N_15454);
nor U22971 (N_22971,N_15817,N_16070);
or U22972 (N_22972,N_18816,N_17233);
and U22973 (N_22973,N_19881,N_11523);
and U22974 (N_22974,N_15696,N_17465);
or U22975 (N_22975,N_11588,N_11416);
nor U22976 (N_22976,N_19380,N_18299);
and U22977 (N_22977,N_12556,N_18227);
nor U22978 (N_22978,N_14133,N_10246);
xor U22979 (N_22979,N_13584,N_11869);
xnor U22980 (N_22980,N_15185,N_11791);
nor U22981 (N_22981,N_10365,N_19167);
nor U22982 (N_22982,N_15855,N_16938);
or U22983 (N_22983,N_12336,N_13137);
and U22984 (N_22984,N_18715,N_14289);
nand U22985 (N_22985,N_11913,N_18631);
nor U22986 (N_22986,N_14057,N_19508);
nor U22987 (N_22987,N_10100,N_13429);
and U22988 (N_22988,N_13403,N_10494);
or U22989 (N_22989,N_14053,N_17445);
nor U22990 (N_22990,N_12580,N_19980);
nand U22991 (N_22991,N_13493,N_15053);
and U22992 (N_22992,N_16402,N_17867);
and U22993 (N_22993,N_19281,N_18606);
xor U22994 (N_22994,N_11943,N_15293);
or U22995 (N_22995,N_11084,N_15530);
nor U22996 (N_22996,N_12109,N_17165);
nor U22997 (N_22997,N_16626,N_11440);
nor U22998 (N_22998,N_13969,N_10245);
and U22999 (N_22999,N_16804,N_14581);
or U23000 (N_23000,N_13484,N_10813);
and U23001 (N_23001,N_18077,N_13555);
nor U23002 (N_23002,N_16784,N_11333);
nor U23003 (N_23003,N_15255,N_19707);
xor U23004 (N_23004,N_16717,N_16527);
nand U23005 (N_23005,N_15441,N_12174);
nand U23006 (N_23006,N_16497,N_19488);
nor U23007 (N_23007,N_18484,N_18143);
or U23008 (N_23008,N_16161,N_16363);
or U23009 (N_23009,N_16759,N_12142);
and U23010 (N_23010,N_10684,N_18653);
or U23011 (N_23011,N_17666,N_18256);
or U23012 (N_23012,N_17671,N_17746);
nand U23013 (N_23013,N_17204,N_15941);
and U23014 (N_23014,N_12780,N_13377);
xnor U23015 (N_23015,N_15580,N_14220);
nand U23016 (N_23016,N_19022,N_11555);
and U23017 (N_23017,N_19944,N_10818);
xor U23018 (N_23018,N_17745,N_13638);
and U23019 (N_23019,N_12700,N_17501);
xnor U23020 (N_23020,N_12474,N_13725);
and U23021 (N_23021,N_12137,N_19882);
xor U23022 (N_23022,N_12298,N_17292);
nor U23023 (N_23023,N_14514,N_13598);
and U23024 (N_23024,N_10181,N_12913);
nor U23025 (N_23025,N_12381,N_18544);
nor U23026 (N_23026,N_10615,N_13551);
nor U23027 (N_23027,N_18450,N_19230);
and U23028 (N_23028,N_15722,N_16097);
and U23029 (N_23029,N_10325,N_19626);
and U23030 (N_23030,N_10429,N_10681);
and U23031 (N_23031,N_11117,N_12540);
nor U23032 (N_23032,N_15322,N_19822);
nand U23033 (N_23033,N_14487,N_11427);
nand U23034 (N_23034,N_10306,N_12078);
nand U23035 (N_23035,N_16396,N_11098);
and U23036 (N_23036,N_18671,N_12152);
and U23037 (N_23037,N_17330,N_12760);
nand U23038 (N_23038,N_16194,N_15944);
and U23039 (N_23039,N_15435,N_18367);
or U23040 (N_23040,N_16736,N_15227);
or U23041 (N_23041,N_10355,N_12737);
nor U23042 (N_23042,N_11380,N_15213);
or U23043 (N_23043,N_17574,N_12146);
xnor U23044 (N_23044,N_15262,N_13681);
and U23045 (N_23045,N_11563,N_17688);
xnor U23046 (N_23046,N_12858,N_11082);
nor U23047 (N_23047,N_10798,N_15881);
nand U23048 (N_23048,N_18003,N_16798);
nor U23049 (N_23049,N_18605,N_19245);
xnor U23050 (N_23050,N_12420,N_12681);
or U23051 (N_23051,N_18165,N_17255);
and U23052 (N_23052,N_10406,N_15557);
or U23053 (N_23053,N_11589,N_14340);
nor U23054 (N_23054,N_14307,N_15096);
or U23055 (N_23055,N_11792,N_10479);
xor U23056 (N_23056,N_12253,N_15926);
or U23057 (N_23057,N_16469,N_13689);
or U23058 (N_23058,N_14877,N_14457);
or U23059 (N_23059,N_10113,N_17990);
nor U23060 (N_23060,N_14058,N_13388);
xnor U23061 (N_23061,N_13896,N_10752);
nand U23062 (N_23062,N_13694,N_14467);
nand U23063 (N_23063,N_15374,N_12139);
or U23064 (N_23064,N_18688,N_16095);
nor U23065 (N_23065,N_18251,N_17071);
nor U23066 (N_23066,N_16121,N_15383);
nand U23067 (N_23067,N_10610,N_11040);
nand U23068 (N_23068,N_19483,N_19663);
and U23069 (N_23069,N_16385,N_10457);
and U23070 (N_23070,N_10560,N_18114);
or U23071 (N_23071,N_15747,N_17641);
and U23072 (N_23072,N_14847,N_16433);
or U23073 (N_23073,N_17902,N_12887);
nand U23074 (N_23074,N_18366,N_11224);
xor U23075 (N_23075,N_15616,N_17923);
nand U23076 (N_23076,N_12279,N_18157);
and U23077 (N_23077,N_19283,N_16291);
nand U23078 (N_23078,N_10477,N_10716);
nor U23079 (N_23079,N_17199,N_13613);
and U23080 (N_23080,N_16351,N_17018);
and U23081 (N_23081,N_17795,N_14541);
and U23082 (N_23082,N_14405,N_12831);
nor U23083 (N_23083,N_14100,N_15052);
xor U23084 (N_23084,N_12053,N_12356);
or U23085 (N_23085,N_16186,N_12830);
or U23086 (N_23086,N_18208,N_18567);
nor U23087 (N_23087,N_18807,N_19289);
or U23088 (N_23088,N_15820,N_10843);
and U23089 (N_23089,N_14152,N_12006);
nand U23090 (N_23090,N_10356,N_17384);
or U23091 (N_23091,N_10350,N_14038);
nand U23092 (N_23092,N_11692,N_13774);
or U23093 (N_23093,N_13146,N_15874);
nand U23094 (N_23094,N_11057,N_14523);
or U23095 (N_23095,N_19524,N_18275);
nand U23096 (N_23096,N_19276,N_11663);
or U23097 (N_23097,N_11918,N_10260);
or U23098 (N_23098,N_16913,N_19902);
nor U23099 (N_23099,N_18571,N_17966);
or U23100 (N_23100,N_17631,N_18855);
nor U23101 (N_23101,N_13052,N_10656);
or U23102 (N_23102,N_16586,N_18790);
xor U23103 (N_23103,N_14752,N_12870);
nor U23104 (N_23104,N_10050,N_15344);
nand U23105 (N_23105,N_19363,N_18211);
xnor U23106 (N_23106,N_14544,N_11607);
or U23107 (N_23107,N_17593,N_10440);
nand U23108 (N_23108,N_11307,N_15795);
xnor U23109 (N_23109,N_15808,N_18957);
nor U23110 (N_23110,N_19084,N_15764);
nand U23111 (N_23111,N_14868,N_14992);
and U23112 (N_23112,N_10318,N_19170);
nor U23113 (N_23113,N_12833,N_16240);
and U23114 (N_23114,N_14520,N_15128);
nand U23115 (N_23115,N_11384,N_11372);
and U23116 (N_23116,N_14942,N_17663);
nand U23117 (N_23117,N_10445,N_16656);
nand U23118 (N_23118,N_19702,N_10212);
and U23119 (N_23119,N_14986,N_10960);
nand U23120 (N_23120,N_17766,N_18950);
nor U23121 (N_23121,N_15430,N_19947);
nand U23122 (N_23122,N_16259,N_12380);
or U23123 (N_23123,N_11926,N_10934);
or U23124 (N_23124,N_14673,N_11391);
nand U23125 (N_23125,N_14919,N_14222);
and U23126 (N_23126,N_12220,N_11797);
nand U23127 (N_23127,N_19407,N_14088);
nor U23128 (N_23128,N_17397,N_18337);
nand U23129 (N_23129,N_11566,N_15870);
xnor U23130 (N_23130,N_15921,N_17153);
nor U23131 (N_23131,N_17436,N_18005);
nor U23132 (N_23132,N_13687,N_14076);
or U23133 (N_23133,N_16266,N_19557);
and U23134 (N_23134,N_12647,N_10879);
and U23135 (N_23135,N_17278,N_16373);
xnor U23136 (N_23136,N_16676,N_18014);
xor U23137 (N_23137,N_14994,N_19657);
nor U23138 (N_23138,N_12393,N_14095);
or U23139 (N_23139,N_11493,N_16624);
and U23140 (N_23140,N_19520,N_13323);
xnor U23141 (N_23141,N_10418,N_13361);
or U23142 (N_23142,N_17757,N_18540);
or U23143 (N_23143,N_19138,N_15371);
or U23144 (N_23144,N_11483,N_19438);
xnor U23145 (N_23145,N_18573,N_11353);
nand U23146 (N_23146,N_13757,N_17287);
and U23147 (N_23147,N_18396,N_19411);
nand U23148 (N_23148,N_15960,N_10951);
and U23149 (N_23149,N_12931,N_11915);
nor U23150 (N_23150,N_13649,N_13413);
or U23151 (N_23151,N_13766,N_19999);
nand U23152 (N_23152,N_14329,N_17675);
nor U23153 (N_23153,N_16004,N_13445);
and U23154 (N_23154,N_17528,N_18414);
and U23155 (N_23155,N_15997,N_18323);
nor U23156 (N_23156,N_12867,N_18918);
nor U23157 (N_23157,N_13394,N_15448);
or U23158 (N_23158,N_16588,N_19889);
nor U23159 (N_23159,N_11212,N_18873);
and U23160 (N_23160,N_16815,N_13952);
nor U23161 (N_23161,N_11823,N_14684);
nand U23162 (N_23162,N_13949,N_18555);
and U23163 (N_23163,N_15393,N_12604);
and U23164 (N_23164,N_13675,N_15258);
nand U23165 (N_23165,N_16328,N_15177);
and U23166 (N_23166,N_10718,N_10054);
nor U23167 (N_23167,N_15396,N_19059);
xor U23168 (N_23168,N_16537,N_12546);
and U23169 (N_23169,N_17222,N_17163);
xnor U23170 (N_23170,N_12797,N_18432);
nand U23171 (N_23171,N_18019,N_15190);
and U23172 (N_23172,N_17112,N_11928);
nor U23173 (N_23173,N_11649,N_19538);
and U23174 (N_23174,N_14975,N_10463);
and U23175 (N_23175,N_14938,N_10190);
and U23176 (N_23176,N_16944,N_10002);
and U23177 (N_23177,N_14924,N_15970);
and U23178 (N_23178,N_13667,N_18358);
nand U23179 (N_23179,N_16164,N_18676);
nor U23180 (N_23180,N_17457,N_13791);
or U23181 (N_23181,N_13112,N_19114);
nand U23182 (N_23182,N_16642,N_17390);
nand U23183 (N_23183,N_12612,N_18680);
or U23184 (N_23184,N_16603,N_15051);
or U23185 (N_23185,N_16640,N_16289);
and U23186 (N_23186,N_10125,N_17546);
xnor U23187 (N_23187,N_13246,N_11703);
and U23188 (N_23188,N_10149,N_17312);
nor U23189 (N_23189,N_16823,N_13252);
xor U23190 (N_23190,N_19545,N_19187);
or U23191 (N_23191,N_19442,N_17226);
and U23192 (N_23192,N_13536,N_14108);
xor U23193 (N_23193,N_12537,N_11075);
nor U23194 (N_23194,N_12057,N_12558);
and U23195 (N_23195,N_10015,N_11729);
nand U23196 (N_23196,N_16714,N_15373);
nand U23197 (N_23197,N_10411,N_10404);
and U23198 (N_23198,N_16508,N_16549);
xnor U23199 (N_23199,N_13081,N_11503);
or U23200 (N_23200,N_13634,N_17507);
or U23201 (N_23201,N_12204,N_15911);
and U23202 (N_23202,N_12950,N_12452);
nand U23203 (N_23203,N_17295,N_10098);
or U23204 (N_23204,N_11917,N_14912);
nand U23205 (N_23205,N_18226,N_14841);
and U23206 (N_23206,N_18891,N_13481);
nor U23207 (N_23207,N_12689,N_16881);
nand U23208 (N_23208,N_18206,N_17369);
nand U23209 (N_23209,N_15744,N_19555);
or U23210 (N_23210,N_12926,N_15226);
and U23211 (N_23211,N_17721,N_17603);
nor U23212 (N_23212,N_17514,N_15392);
and U23213 (N_23213,N_16902,N_16359);
nor U23214 (N_23214,N_10179,N_19691);
nor U23215 (N_23215,N_19209,N_18046);
nand U23216 (N_23216,N_16557,N_14007);
nand U23217 (N_23217,N_15971,N_13963);
nor U23218 (N_23218,N_10025,N_10579);
nand U23219 (N_23219,N_13983,N_13166);
nor U23220 (N_23220,N_16371,N_13745);
and U23221 (N_23221,N_13349,N_13625);
or U23222 (N_23222,N_16742,N_13464);
or U23223 (N_23223,N_16088,N_19973);
nor U23224 (N_23224,N_12321,N_14176);
or U23225 (N_23225,N_16157,N_16747);
or U23226 (N_23226,N_14630,N_13308);
or U23227 (N_23227,N_12560,N_11406);
or U23228 (N_23228,N_19895,N_13221);
nand U23229 (N_23229,N_19695,N_14940);
xnor U23230 (N_23230,N_14205,N_17288);
nand U23231 (N_23231,N_14462,N_15753);
nor U23232 (N_23232,N_14565,N_12136);
and U23233 (N_23233,N_18269,N_16741);
nand U23234 (N_23234,N_19760,N_11513);
nand U23235 (N_23235,N_10140,N_16936);
nand U23236 (N_23236,N_18392,N_12752);
xnor U23237 (N_23237,N_10696,N_17052);
nor U23238 (N_23238,N_17930,N_13075);
and U23239 (N_23239,N_19398,N_10109);
and U23240 (N_23240,N_14963,N_19409);
and U23241 (N_23241,N_17984,N_10114);
and U23242 (N_23242,N_13895,N_13619);
xor U23243 (N_23243,N_12255,N_17066);
nand U23244 (N_23244,N_11053,N_19525);
or U23245 (N_23245,N_16042,N_14528);
nor U23246 (N_23246,N_19749,N_19577);
xor U23247 (N_23247,N_10917,N_11217);
or U23248 (N_23248,N_16910,N_11967);
xnor U23249 (N_23249,N_13862,N_17937);
xnor U23250 (N_23250,N_17157,N_18451);
nand U23251 (N_23251,N_18139,N_12590);
nand U23252 (N_23252,N_19818,N_12373);
xnor U23253 (N_23253,N_18719,N_11587);
xor U23254 (N_23254,N_12776,N_11977);
xnor U23255 (N_23255,N_14763,N_16595);
or U23256 (N_23256,N_16400,N_14449);
or U23257 (N_23257,N_10538,N_19809);
nand U23258 (N_23258,N_13734,N_16413);
or U23259 (N_23259,N_15684,N_10481);
nand U23260 (N_23260,N_19339,N_10675);
xor U23261 (N_23261,N_10062,N_16358);
nand U23262 (N_23262,N_14804,N_15505);
and U23263 (N_23263,N_13962,N_17662);
xnor U23264 (N_23264,N_17872,N_12785);
nand U23265 (N_23265,N_15634,N_16674);
and U23266 (N_23266,N_12494,N_18856);
nand U23267 (N_23267,N_19743,N_14103);
and U23268 (N_23268,N_19161,N_17636);
or U23269 (N_23269,N_11028,N_15010);
nor U23270 (N_23270,N_13506,N_13451);
nor U23271 (N_23271,N_19768,N_11293);
and U23272 (N_23272,N_10102,N_12130);
or U23273 (N_23273,N_13676,N_18660);
nand U23274 (N_23274,N_19959,N_14643);
nand U23275 (N_23275,N_12587,N_13392);
or U23276 (N_23276,N_12589,N_14160);
nand U23277 (N_23277,N_19368,N_17643);
nor U23278 (N_23278,N_19375,N_19614);
and U23279 (N_23279,N_18580,N_10525);
nand U23280 (N_23280,N_14742,N_13241);
nand U23281 (N_23281,N_12294,N_16597);
or U23282 (N_23282,N_11571,N_18699);
nand U23283 (N_23283,N_18841,N_16663);
xnor U23284 (N_23284,N_18055,N_15439);
nor U23285 (N_23285,N_10633,N_14259);
or U23286 (N_23286,N_18735,N_16089);
and U23287 (N_23287,N_15603,N_10137);
or U23288 (N_23288,N_15972,N_12270);
and U23289 (N_23289,N_16101,N_15914);
nor U23290 (N_23290,N_12706,N_19634);
nor U23291 (N_23291,N_12736,N_16484);
and U23292 (N_23292,N_13759,N_11143);
nor U23293 (N_23293,N_13288,N_17621);
and U23294 (N_23294,N_13611,N_18773);
or U23295 (N_23295,N_17908,N_19929);
nand U23296 (N_23296,N_12906,N_14181);
and U23297 (N_23297,N_12176,N_18079);
nand U23298 (N_23298,N_11009,N_18885);
nor U23299 (N_23299,N_13960,N_18568);
nor U23300 (N_23300,N_14599,N_14463);
nor U23301 (N_23301,N_19912,N_17542);
and U23302 (N_23302,N_13375,N_18308);
nor U23303 (N_23303,N_14104,N_16790);
or U23304 (N_23304,N_14438,N_16159);
xor U23305 (N_23305,N_19436,N_10112);
nand U23306 (N_23306,N_19035,N_12213);
and U23307 (N_23307,N_15709,N_17695);
or U23308 (N_23308,N_13180,N_14458);
nand U23309 (N_23309,N_13861,N_12017);
nor U23310 (N_23310,N_10336,N_17967);
or U23311 (N_23311,N_17010,N_11786);
nand U23312 (N_23312,N_11463,N_19395);
nor U23313 (N_23313,N_17101,N_18277);
or U23314 (N_23314,N_16937,N_15118);
nand U23315 (N_23315,N_18897,N_10028);
and U23316 (N_23316,N_19503,N_15386);
nand U23317 (N_23317,N_11154,N_14230);
and U23318 (N_23318,N_18281,N_19458);
nor U23319 (N_23319,N_17611,N_19248);
xor U23320 (N_23320,N_13415,N_18870);
nor U23321 (N_23321,N_12068,N_11363);
nand U23322 (N_23322,N_14628,N_18527);
and U23323 (N_23323,N_19958,N_16146);
or U23324 (N_23324,N_13901,N_16495);
and U23325 (N_23325,N_10651,N_10545);
nor U23326 (N_23326,N_19754,N_12233);
nor U23327 (N_23327,N_12163,N_13696);
or U23328 (N_23328,N_10204,N_18742);
nor U23329 (N_23329,N_14023,N_17421);
and U23330 (N_23330,N_16096,N_10558);
or U23331 (N_23331,N_19304,N_18733);
xor U23332 (N_23332,N_18236,N_12154);
xnor U23333 (N_23333,N_14065,N_18020);
nand U23334 (N_23334,N_18624,N_18784);
nand U23335 (N_23335,N_19674,N_13320);
nor U23336 (N_23336,N_12234,N_10337);
nand U23337 (N_23337,N_17629,N_17342);
nand U23338 (N_23338,N_18603,N_15597);
xnor U23339 (N_23339,N_14415,N_15188);
or U23340 (N_23340,N_15423,N_15509);
or U23341 (N_23341,N_14227,N_10898);
or U23342 (N_23342,N_18336,N_10264);
nand U23343 (N_23343,N_17234,N_12226);
nand U23344 (N_23344,N_19848,N_13892);
or U23345 (N_23345,N_10709,N_13537);
nand U23346 (N_23346,N_11843,N_18994);
nor U23347 (N_23347,N_12947,N_15029);
xor U23348 (N_23348,N_12012,N_15486);
xor U23349 (N_23349,N_17031,N_13164);
nor U23350 (N_23350,N_13076,N_13446);
nor U23351 (N_23351,N_16056,N_15847);
nand U23352 (N_23352,N_15176,N_19452);
xor U23353 (N_23353,N_11430,N_15137);
or U23354 (N_23354,N_11238,N_10632);
and U23355 (N_23355,N_11546,N_16207);
and U23356 (N_23356,N_13819,N_11016);
and U23357 (N_23357,N_11195,N_13197);
and U23358 (N_23358,N_18225,N_10557);
nor U23359 (N_23359,N_17202,N_10873);
nor U23360 (N_23360,N_14722,N_14903);
and U23361 (N_23361,N_15211,N_14069);
and U23362 (N_23362,N_15220,N_16375);
nor U23363 (N_23363,N_19647,N_17997);
and U23364 (N_23364,N_12490,N_14831);
and U23365 (N_23365,N_18710,N_17656);
nor U23366 (N_23366,N_12165,N_17187);
or U23367 (N_23367,N_19162,N_16949);
nand U23368 (N_23368,N_12798,N_19666);
and U23369 (N_23369,N_18198,N_15288);
and U23370 (N_23370,N_10705,N_14720);
or U23371 (N_23371,N_17466,N_13604);
nand U23372 (N_23372,N_19338,N_15683);
and U23373 (N_23373,N_17522,N_10968);
nor U23374 (N_23374,N_14612,N_16947);
nand U23375 (N_23375,N_14102,N_11281);
and U23376 (N_23376,N_12770,N_15210);
nor U23377 (N_23377,N_14734,N_16992);
and U23378 (N_23378,N_14011,N_11806);
nand U23379 (N_23379,N_16604,N_12469);
xor U23380 (N_23380,N_15518,N_18221);
xor U23381 (N_23381,N_10617,N_12407);
or U23382 (N_23382,N_16378,N_18626);
xnor U23383 (N_23383,N_15054,N_13524);
and U23384 (N_23384,N_16725,N_18748);
nand U23385 (N_23385,N_13049,N_14606);
nand U23386 (N_23386,N_14566,N_18590);
xor U23387 (N_23387,N_13279,N_17194);
nand U23388 (N_23388,N_17058,N_17670);
nand U23389 (N_23389,N_19198,N_16006);
nor U23390 (N_23390,N_11795,N_19221);
and U23391 (N_23391,N_15720,N_14276);
nand U23392 (N_23392,N_13074,N_11180);
nor U23393 (N_23393,N_11827,N_12476);
or U23394 (N_23394,N_11798,N_18775);
nand U23395 (N_23395,N_13589,N_13383);
and U23396 (N_23396,N_16181,N_15822);
or U23397 (N_23397,N_14301,N_18001);
nand U23398 (N_23398,N_12641,N_12375);
nor U23399 (N_23399,N_13872,N_18328);
or U23400 (N_23400,N_19758,N_17547);
and U23401 (N_23401,N_15356,N_12970);
nand U23402 (N_23402,N_18385,N_11437);
and U23403 (N_23403,N_16956,N_11821);
nor U23404 (N_23404,N_13929,N_19753);
and U23405 (N_23405,N_15880,N_10619);
nor U23406 (N_23406,N_11828,N_10714);
nor U23407 (N_23407,N_11176,N_18898);
and U23408 (N_23408,N_12179,N_14675);
nand U23409 (N_23409,N_19628,N_13871);
or U23410 (N_23410,N_10536,N_12955);
nand U23411 (N_23411,N_18863,N_15669);
or U23412 (N_23412,N_19708,N_11885);
nand U23413 (N_23413,N_12398,N_11486);
or U23414 (N_23414,N_11707,N_12450);
and U23415 (N_23415,N_18031,N_13410);
nor U23416 (N_23416,N_15598,N_13948);
and U23417 (N_23417,N_11035,N_16305);
nand U23418 (N_23418,N_14122,N_14291);
or U23419 (N_23419,N_17291,N_18743);
nor U23420 (N_23420,N_17635,N_12994);
or U23421 (N_23421,N_19063,N_11676);
or U23422 (N_23422,N_17365,N_14151);
and U23423 (N_23423,N_17216,N_19855);
nor U23424 (N_23424,N_10471,N_18611);
or U23425 (N_23425,N_10302,N_16448);
or U23426 (N_23426,N_10527,N_14400);
and U23427 (N_23427,N_17866,N_18681);
or U23428 (N_23428,N_12627,N_18486);
and U23429 (N_23429,N_13933,N_13416);
or U23430 (N_23430,N_18271,N_18261);
or U23431 (N_23431,N_17325,N_11852);
nor U23432 (N_23432,N_11601,N_13300);
nor U23433 (N_23433,N_16969,N_11529);
xor U23434 (N_23434,N_15939,N_19078);
xor U23435 (N_23435,N_16453,N_18292);
nand U23436 (N_23436,N_14497,N_15727);
and U23437 (N_23437,N_16994,N_15301);
and U23438 (N_23438,N_16107,N_16822);
and U23439 (N_23439,N_17335,N_17249);
or U23440 (N_23440,N_11603,N_19041);
or U23441 (N_23441,N_12787,N_15457);
or U23442 (N_23442,N_18842,N_14904);
nand U23443 (N_23443,N_17979,N_13477);
or U23444 (N_23444,N_10967,N_14187);
and U23445 (N_23445,N_12657,N_10791);
nor U23446 (N_23446,N_11696,N_15864);
and U23447 (N_23447,N_11820,N_17864);
and U23448 (N_23448,N_12541,N_19616);
nand U23449 (N_23449,N_16887,N_11738);
nor U23450 (N_23450,N_15151,N_19376);
and U23451 (N_23451,N_17022,N_17277);
nand U23452 (N_23452,N_18458,N_19678);
nor U23453 (N_23453,N_19461,N_13297);
and U23454 (N_23454,N_18936,N_14886);
and U23455 (N_23455,N_10894,N_11890);
nor U23456 (N_23456,N_18454,N_17075);
nor U23457 (N_23457,N_14766,N_11547);
nand U23458 (N_23458,N_16211,N_12834);
xor U23459 (N_23459,N_19141,N_11110);
xor U23460 (N_23460,N_11557,N_10421);
and U23461 (N_23461,N_19016,N_15252);
and U23462 (N_23462,N_13117,N_19300);
xnor U23463 (N_23463,N_13450,N_16825);
nand U23464 (N_23464,N_11310,N_11072);
and U23465 (N_23465,N_13498,N_17241);
and U23466 (N_23466,N_18039,N_19513);
and U23467 (N_23467,N_18418,N_16459);
nor U23468 (N_23468,N_11285,N_13592);
nand U23469 (N_23469,N_18494,N_11637);
and U23470 (N_23470,N_14971,N_15403);
or U23471 (N_23471,N_16447,N_11096);
nand U23472 (N_23472,N_12889,N_14813);
nand U23473 (N_23473,N_13542,N_12812);
nand U23474 (N_23474,N_16094,N_18643);
or U23475 (N_23475,N_11783,N_14666);
and U23476 (N_23476,N_13605,N_11751);
or U23477 (N_23477,N_11537,N_11613);
xor U23478 (N_23478,N_15324,N_17959);
nor U23479 (N_23479,N_16564,N_13903);
nand U23480 (N_23480,N_13363,N_12461);
nor U23481 (N_23481,N_10640,N_10387);
nor U23482 (N_23482,N_13474,N_14803);
nor U23483 (N_23483,N_14303,N_15807);
and U23484 (N_23484,N_17602,N_16273);
nand U23485 (N_23485,N_16585,N_13163);
or U23486 (N_23486,N_11173,N_10304);
or U23487 (N_23487,N_15564,N_16678);
or U23488 (N_23488,N_10868,N_15375);
or U23489 (N_23489,N_10193,N_16492);
and U23490 (N_23490,N_10986,N_16331);
nand U23491 (N_23491,N_11074,N_17906);
and U23492 (N_23492,N_16401,N_12023);
xnor U23493 (N_23493,N_19182,N_19851);
and U23494 (N_23494,N_19998,N_10222);
or U23495 (N_23495,N_15981,N_15238);
nand U23496 (N_23496,N_19962,N_12432);
nor U23497 (N_23497,N_16279,N_17357);
and U23498 (N_23498,N_11460,N_12082);
xnor U23499 (N_23499,N_10690,N_13781);
or U23500 (N_23500,N_11104,N_14431);
or U23501 (N_23501,N_19440,N_16471);
or U23502 (N_23502,N_12715,N_13558);
nor U23503 (N_23503,N_18513,N_16064);
nand U23504 (N_23504,N_15140,N_11086);
nand U23505 (N_23505,N_10533,N_13225);
nor U23506 (N_23506,N_14657,N_14296);
xnor U23507 (N_23507,N_10876,N_16552);
or U23508 (N_23508,N_17451,N_12386);
or U23509 (N_23509,N_19226,N_19588);
nor U23510 (N_23510,N_18324,N_10247);
nand U23511 (N_23511,N_10655,N_19532);
nor U23512 (N_23512,N_17057,N_19955);
nor U23513 (N_23513,N_14622,N_14437);
xor U23514 (N_23514,N_15060,N_15031);
or U23515 (N_23515,N_17125,N_17109);
or U23516 (N_23516,N_14124,N_17929);
and U23517 (N_23517,N_19134,N_10985);
nor U23518 (N_23518,N_12147,N_16914);
nor U23519 (N_23519,N_15186,N_12989);
and U23520 (N_23520,N_10465,N_13956);
xor U23521 (N_23521,N_18578,N_19856);
or U23522 (N_23522,N_10601,N_11171);
and U23523 (N_23523,N_10163,N_14956);
and U23524 (N_23524,N_15756,N_19191);
nor U23525 (N_23525,N_11323,N_19185);
or U23526 (N_23526,N_18188,N_10991);
and U23527 (N_23527,N_18766,N_15625);
nor U23528 (N_23528,N_17096,N_12378);
or U23529 (N_23529,N_16183,N_12437);
nor U23530 (N_23530,N_19799,N_12009);
and U23531 (N_23531,N_18220,N_16128);
xor U23532 (N_23532,N_14077,N_15908);
nand U23533 (N_23533,N_16919,N_15878);
nand U23534 (N_23534,N_11704,N_15638);
nand U23535 (N_23535,N_14848,N_12455);
nor U23536 (N_23536,N_17323,N_11300);
or U23537 (N_23537,N_16071,N_19110);
nor U23538 (N_23538,N_12300,N_15136);
nor U23539 (N_23539,N_13325,N_18542);
xnor U23540 (N_23540,N_10664,N_15728);
nand U23541 (N_23541,N_16688,N_15877);
xnor U23542 (N_23542,N_16862,N_14029);
and U23543 (N_23543,N_11263,N_10110);
nor U23544 (N_23544,N_15889,N_10521);
and U23545 (N_23545,N_15360,N_13402);
and U23546 (N_23546,N_15922,N_18121);
or U23547 (N_23547,N_17708,N_19267);
nand U23548 (N_23548,N_15796,N_13274);
and U23549 (N_23549,N_16411,N_12125);
or U23550 (N_23550,N_11590,N_12392);
or U23551 (N_23551,N_19821,N_18587);
or U23552 (N_23552,N_19055,N_14983);
and U23553 (N_23553,N_11213,N_17771);
nor U23554 (N_23554,N_16043,N_16820);
or U23555 (N_23555,N_19070,N_16608);
nand U23556 (N_23556,N_18296,N_14937);
and U23557 (N_23557,N_19970,N_12070);
and U23558 (N_23558,N_12599,N_16556);
nand U23559 (N_23559,N_13522,N_13480);
or U23560 (N_23560,N_16298,N_18207);
nor U23561 (N_23561,N_12571,N_11790);
and U23562 (N_23562,N_15222,N_12941);
or U23563 (N_23563,N_19000,N_13195);
xor U23564 (N_23564,N_17419,N_19225);
nor U23565 (N_23565,N_12854,N_15045);
or U23566 (N_23566,N_13294,N_12684);
nand U23567 (N_23567,N_16638,N_19653);
nor U23568 (N_23568,N_15406,N_11983);
or U23569 (N_23569,N_18520,N_17932);
nor U23570 (N_23570,N_12946,N_10503);
and U23571 (N_23571,N_11091,N_15993);
or U23572 (N_23572,N_11584,N_19391);
nor U23573 (N_23573,N_16498,N_13577);
nand U23574 (N_23574,N_11375,N_14634);
nor U23575 (N_23575,N_18820,N_19847);
nand U23576 (N_23576,N_14899,N_12274);
nor U23577 (N_23577,N_15402,N_15282);
and U23578 (N_23578,N_19139,N_14036);
and U23579 (N_23579,N_18471,N_18799);
and U23580 (N_23580,N_14455,N_13780);
or U23581 (N_23581,N_15088,N_17709);
nand U23582 (N_23582,N_16929,N_13543);
xor U23583 (N_23583,N_11223,N_13918);
nand U23584 (N_23584,N_18360,N_14801);
and U23585 (N_23585,N_18979,N_16764);
or U23586 (N_23586,N_13455,N_14775);
or U23587 (N_23587,N_19693,N_13525);
or U23588 (N_23588,N_11237,N_10068);
or U23589 (N_23589,N_11111,N_13538);
nor U23590 (N_23590,N_12099,N_14022);
or U23591 (N_23591,N_15622,N_18259);
or U23592 (N_23592,N_18253,N_17437);
or U23593 (N_23593,N_13877,N_10574);
and U23594 (N_23594,N_18428,N_10286);
nand U23595 (N_23595,N_18026,N_13067);
or U23596 (N_23596,N_15132,N_17523);
or U23597 (N_23597,N_16864,N_12241);
and U23598 (N_23598,N_17375,N_15907);
and U23599 (N_23599,N_18796,N_18100);
xor U23600 (N_23600,N_17814,N_13092);
nand U23601 (N_23601,N_11646,N_17784);
nor U23602 (N_23602,N_17128,N_14422);
and U23603 (N_23603,N_17974,N_15025);
or U23604 (N_23604,N_17127,N_15030);
and U23605 (N_23605,N_10539,N_19988);
or U23606 (N_23606,N_12302,N_17753);
and U23607 (N_23607,N_11387,N_19930);
and U23608 (N_23608,N_19415,N_19089);
nor U23609 (N_23609,N_10700,N_17014);
or U23610 (N_23610,N_12674,N_16898);
or U23611 (N_23611,N_13920,N_15628);
xnor U23612 (N_23612,N_11754,N_12309);
nand U23613 (N_23613,N_12965,N_10165);
or U23614 (N_23614,N_11916,N_19596);
nand U23615 (N_23615,N_16137,N_19430);
nand U23616 (N_23616,N_14811,N_18228);
nand U23617 (N_23617,N_10049,N_13200);
and U23618 (N_23618,N_10400,N_13069);
nand U23619 (N_23619,N_15535,N_16001);
nand U23620 (N_23620,N_14616,N_16105);
and U23621 (N_23621,N_16679,N_11451);
and U23622 (N_23622,N_11311,N_19739);
nand U23623 (N_23623,N_17091,N_10999);
and U23624 (N_23624,N_12594,N_17520);
and U23625 (N_23625,N_15294,N_10309);
nor U23626 (N_23626,N_12939,N_11344);
or U23627 (N_23627,N_19444,N_16407);
or U23628 (N_23628,N_18200,N_12451);
nand U23629 (N_23629,N_19574,N_18177);
or U23630 (N_23630,N_17488,N_13345);
nor U23631 (N_23631,N_12962,N_10366);
nand U23632 (N_23632,N_10661,N_14888);
or U23633 (N_23633,N_13771,N_10449);
and U23634 (N_23634,N_14537,N_15959);
or U23635 (N_23635,N_18485,N_12278);
xnor U23636 (N_23636,N_17877,N_13822);
and U23637 (N_23637,N_16504,N_12280);
nor U23638 (N_23638,N_11679,N_13911);
or U23639 (N_23639,N_12330,N_13150);
xnor U23640 (N_23640,N_16777,N_13504);
nor U23641 (N_23641,N_10136,N_12934);
xnor U23642 (N_23642,N_17613,N_17752);
or U23643 (N_23643,N_10293,N_10135);
or U23644 (N_23644,N_18965,N_16219);
and U23645 (N_23645,N_14280,N_18289);
nor U23646 (N_23646,N_19246,N_14856);
nand U23647 (N_23647,N_17499,N_18880);
and U23648 (N_23648,N_15906,N_16895);
nor U23649 (N_23649,N_14654,N_13314);
nor U23650 (N_23650,N_12759,N_13248);
and U23651 (N_23651,N_15270,N_10746);
or U23652 (N_23652,N_17782,N_12264);
and U23653 (N_23653,N_10153,N_13201);
and U23654 (N_23654,N_17205,N_15138);
nor U23655 (N_23655,N_12445,N_16540);
nand U23656 (N_23656,N_16282,N_11153);
nand U23657 (N_23657,N_18669,N_17453);
nand U23658 (N_23658,N_12485,N_19667);
nand U23659 (N_23659,N_15674,N_17107);
or U23660 (N_23660,N_11119,N_11897);
and U23661 (N_23661,N_17622,N_16031);
nand U23662 (N_23662,N_19578,N_10722);
and U23663 (N_23663,N_13932,N_13393);
or U23664 (N_23664,N_12894,N_16133);
nor U23665 (N_23665,N_18981,N_19603);
and U23666 (N_23666,N_14927,N_13238);
and U23667 (N_23667,N_11609,N_12301);
nor U23668 (N_23668,N_12610,N_18035);
and U23669 (N_23669,N_10267,N_13035);
and U23670 (N_23670,N_10605,N_11312);
or U23671 (N_23671,N_19632,N_17362);
nand U23672 (N_23672,N_10787,N_18903);
nor U23673 (N_23673,N_15571,N_14771);
and U23674 (N_23674,N_10338,N_11978);
xor U23675 (N_23675,N_19287,N_17557);
and U23676 (N_23676,N_12332,N_12597);
or U23677 (N_23677,N_13860,N_16047);
and U23678 (N_23678,N_14498,N_17129);
nor U23679 (N_23679,N_15308,N_16077);
nor U23680 (N_23680,N_19778,N_12539);
xnor U23681 (N_23681,N_13175,N_17237);
nor U23682 (N_23682,N_16152,N_10209);
nand U23683 (N_23683,N_17756,N_15100);
and U23684 (N_23684,N_13210,N_13568);
nor U23685 (N_23685,N_13257,N_14072);
nand U23686 (N_23686,N_10417,N_13597);
nor U23687 (N_23687,N_14884,N_10221);
nor U23688 (N_23688,N_13232,N_18975);
or U23689 (N_23689,N_10611,N_14210);
and U23690 (N_23690,N_12563,N_11121);
and U23691 (N_23691,N_10534,N_14139);
nor U23692 (N_23692,N_17442,N_19504);
or U23693 (N_23693,N_15216,N_10792);
or U23694 (N_23694,N_16442,N_19270);
and U23695 (N_23695,N_15352,N_16327);
nor U23696 (N_23696,N_12513,N_11046);
or U23697 (N_23697,N_16481,N_19752);
or U23698 (N_23698,N_13552,N_19004);
and U23699 (N_23699,N_16108,N_12818);
or U23700 (N_23700,N_12237,N_14882);
nand U23701 (N_23701,N_18738,N_17600);
xor U23702 (N_23702,N_15609,N_19609);
and U23703 (N_23703,N_11265,N_17452);
nand U23704 (N_23704,N_19335,N_15885);
nand U23705 (N_23705,N_18832,N_15584);
nand U23706 (N_23706,N_14292,N_10856);
and U23707 (N_23707,N_19030,N_15900);
nand U23708 (N_23708,N_16546,N_15427);
nand U23709 (N_23709,N_17476,N_19679);
nand U23710 (N_23710,N_12221,N_17878);
or U23711 (N_23711,N_17099,N_19427);
and U23712 (N_23712,N_10379,N_13192);
nand U23713 (N_23713,N_16421,N_15205);
and U23714 (N_23714,N_16163,N_19489);
nor U23715 (N_23715,N_18431,N_13845);
xnor U23716 (N_23716,N_10086,N_12795);
nor U23717 (N_23717,N_16231,N_15549);
nand U23718 (N_23718,N_16252,N_16145);
or U23719 (N_23719,N_12918,N_17174);
or U23720 (N_23720,N_17865,N_16765);
nand U23721 (N_23721,N_19266,N_11953);
nand U23722 (N_23722,N_15725,N_14572);
or U23723 (N_23723,N_13664,N_11327);
nand U23724 (N_23724,N_12936,N_17036);
nand U23725 (N_23725,N_16843,N_10570);
xor U23726 (N_23726,N_11516,N_16308);
and U23727 (N_23727,N_13811,N_18474);
nor U23728 (N_23728,N_17388,N_19036);
nand U23729 (N_23729,N_18564,N_18201);
nand U23730 (N_23730,N_19892,N_12528);
xnor U23731 (N_23731,N_13041,N_16893);
nor U23732 (N_23732,N_18489,N_18826);
and U23733 (N_23733,N_19121,N_10764);
and U23734 (N_23734,N_10587,N_13173);
xnor U23735 (N_23735,N_15113,N_14820);
nand U23736 (N_23736,N_13050,N_15778);
nor U23737 (N_23737,N_12372,N_17597);
and U23738 (N_23738,N_19392,N_14456);
nor U23739 (N_23739,N_10425,N_15105);
nand U23740 (N_23740,N_11041,N_17740);
and U23741 (N_23741,N_15456,N_18584);
nor U23742 (N_23742,N_16846,N_15091);
or U23743 (N_23743,N_19511,N_13921);
or U23744 (N_23744,N_11436,N_15617);
and U23745 (N_23745,N_18375,N_18736);
nor U23746 (N_23746,N_17077,N_15135);
or U23747 (N_23747,N_18417,N_15686);
or U23748 (N_23748,N_15362,N_17378);
or U23749 (N_23749,N_10808,N_19253);
and U23750 (N_23750,N_14098,N_16033);
nand U23751 (N_23751,N_10189,N_18410);
and U23752 (N_23752,N_17843,N_18183);
and U23753 (N_23753,N_10064,N_11257);
nand U23754 (N_23754,N_12171,N_18708);
nor U23755 (N_23755,N_11052,N_14974);
nor U23756 (N_23756,N_12952,N_13557);
nor U23757 (N_23757,N_11941,N_15477);
or U23758 (N_23758,N_18756,N_14507);
and U23759 (N_23759,N_12198,N_10080);
and U23760 (N_23760,N_17254,N_12005);
xnor U23761 (N_23761,N_13510,N_19631);
xor U23762 (N_23762,N_17159,N_12957);
or U23763 (N_23763,N_17970,N_19741);
and U23764 (N_23764,N_15414,N_18406);
xnor U23765 (N_23765,N_15223,N_15183);
or U23766 (N_23766,N_10964,N_15642);
xor U23767 (N_23767,N_12478,N_11457);
nand U23768 (N_23768,N_10765,N_17115);
nor U23769 (N_23769,N_11643,N_17167);
and U23770 (N_23770,N_19406,N_12110);
xor U23771 (N_23771,N_14115,N_13966);
nand U23772 (N_23772,N_12581,N_19572);
nor U23773 (N_23773,N_13635,N_19990);
and U23774 (N_23774,N_16801,N_12899);
or U23775 (N_23775,N_11625,N_12338);
or U23776 (N_23776,N_10691,N_14814);
xor U23777 (N_23777,N_16609,N_10348);
nor U23778 (N_23778,N_16991,N_10918);
and U23779 (N_23779,N_15575,N_12545);
or U23780 (N_23780,N_11428,N_18405);
nand U23781 (N_23781,N_16230,N_14889);
nor U23782 (N_23782,N_12075,N_14761);
nor U23783 (N_23783,N_17983,N_13854);
nor U23784 (N_23784,N_12802,N_19456);
xnor U23785 (N_23785,N_13763,N_17933);
xor U23786 (N_23786,N_14483,N_17408);
xor U23787 (N_23787,N_13078,N_13357);
or U23788 (N_23788,N_10223,N_11247);
nand U23789 (N_23789,N_11136,N_13208);
nor U23790 (N_23790,N_10360,N_12792);
xor U23791 (N_23791,N_16200,N_19402);
xor U23792 (N_23792,N_16849,N_10880);
and U23793 (N_23793,N_13399,N_19750);
nand U23794 (N_23794,N_12601,N_18581);
nor U23795 (N_23795,N_15043,N_18618);
nand U23796 (N_23796,N_16460,N_13738);
and U23797 (N_23797,N_13578,N_11395);
and U23798 (N_23798,N_10486,N_14659);
or U23799 (N_23799,N_14086,N_11531);
nor U23800 (N_23800,N_16269,N_17143);
or U23801 (N_23801,N_19366,N_16990);
or U23802 (N_23802,N_11326,N_15676);
nand U23803 (N_23803,N_14267,N_14099);
and U23804 (N_23804,N_10672,N_17644);
nand U23805 (N_23805,N_10198,N_17469);
nand U23806 (N_23806,N_13973,N_17871);
nor U23807 (N_23807,N_11930,N_12739);
nor U23808 (N_23808,N_13513,N_18609);
nand U23809 (N_23809,N_19159,N_12656);
or U23810 (N_23810,N_13768,N_12116);
or U23811 (N_23811,N_16473,N_19094);
nand U23812 (N_23812,N_17785,N_15041);
nand U23813 (N_23813,N_10497,N_12569);
or U23814 (N_23814,N_10431,N_10997);
nor U23815 (N_23815,N_12972,N_15316);
or U23816 (N_23816,N_18317,N_19655);
nor U23817 (N_23817,N_19553,N_14987);
nor U23818 (N_23818,N_18962,N_19179);
nor U23819 (N_23819,N_16927,N_12733);
or U23820 (N_23820,N_13977,N_18638);
nand U23821 (N_23821,N_19751,N_12620);
nor U23822 (N_23822,N_18869,N_14776);
xnor U23823 (N_23823,N_11012,N_10694);
nand U23824 (N_23824,N_14073,N_12619);
nor U23825 (N_23825,N_13708,N_18574);
nor U23826 (N_23826,N_16271,N_18085);
and U23827 (N_23827,N_10504,N_13023);
nand U23828 (N_23828,N_13271,N_13434);
nor U23829 (N_23829,N_15682,N_19941);
nand U23830 (N_23830,N_11836,N_13692);
nand U23831 (N_23831,N_10774,N_19171);
and U23832 (N_23832,N_15431,N_18664);
nand U23833 (N_23833,N_16877,N_16503);
nand U23834 (N_23834,N_17741,N_10800);
or U23835 (N_23835,N_11817,N_19272);
nor U23836 (N_23836,N_17905,N_15915);
nand U23837 (N_23837,N_17617,N_15447);
nand U23838 (N_23838,N_10621,N_13961);
or U23839 (N_23839,N_12670,N_14433);
and U23840 (N_23840,N_16505,N_15148);
and U23841 (N_23841,N_13643,N_19561);
nand U23842 (N_23842,N_14777,N_16286);
nor U23843 (N_23843,N_12585,N_16435);
and U23844 (N_23844,N_10944,N_18495);
nor U23845 (N_23845,N_16419,N_13423);
or U23846 (N_23846,N_13688,N_13749);
nand U23847 (N_23847,N_17351,N_14547);
and U23848 (N_23848,N_16227,N_11316);
xnor U23849 (N_23849,N_12572,N_13936);
or U23850 (N_23850,N_13214,N_16599);
and U23851 (N_23851,N_19798,N_17754);
xor U23852 (N_23852,N_18937,N_15887);
xnor U23853 (N_23853,N_15982,N_16957);
nand U23854 (N_23854,N_19125,N_16437);
or U23855 (N_23855,N_11175,N_16702);
xnor U23856 (N_23856,N_11039,N_14278);
nand U23857 (N_23857,N_16076,N_10065);
and U23858 (N_23858,N_12119,N_16620);
nand U23859 (N_23859,N_15016,N_13897);
nor U23860 (N_23860,N_17586,N_13535);
or U23861 (N_23861,N_16103,N_16445);
and U23862 (N_23862,N_16581,N_13735);
or U23863 (N_23863,N_10376,N_12127);
nor U23864 (N_23864,N_10954,N_14235);
or U23865 (N_23865,N_15757,N_13595);
or U23866 (N_23866,N_19602,N_11168);
xor U23867 (N_23867,N_19282,N_12084);
nor U23868 (N_23868,N_12817,N_15735);
or U23869 (N_23869,N_10947,N_12547);
or U23870 (N_23870,N_18847,N_12449);
and U23871 (N_23871,N_18262,N_14191);
nor U23872 (N_23872,N_12838,N_17783);
nor U23873 (N_23873,N_15968,N_12559);
or U23874 (N_23874,N_10035,N_10288);
nor U23875 (N_23875,N_15765,N_13756);
nor U23876 (N_23876,N_19687,N_12001);
xor U23877 (N_23877,N_10357,N_16880);
nand U23878 (N_23878,N_10906,N_18951);
or U23879 (N_23879,N_16641,N_15823);
or U23880 (N_23880,N_18913,N_19805);
xnor U23881 (N_23881,N_12122,N_11632);
nand U23882 (N_23882,N_19371,N_19045);
nor U23883 (N_23883,N_12071,N_13003);
and U23884 (N_23884,N_12277,N_13623);
xor U23885 (N_23885,N_18604,N_12284);
and U23886 (N_23886,N_16050,N_14224);
and U23887 (N_23887,N_14309,N_17816);
nand U23888 (N_23888,N_17591,N_15662);
and U23889 (N_23889,N_10520,N_13828);
and U23890 (N_23890,N_13354,N_15556);
nor U23891 (N_23891,N_11209,N_16979);
nand U23892 (N_23892,N_11564,N_17738);
nand U23893 (N_23893,N_17982,N_16046);
or U23894 (N_23894,N_18006,N_17248);
and U23895 (N_23895,N_11123,N_13953);
or U23896 (N_23896,N_12441,N_19683);
or U23897 (N_23897,N_19540,N_10127);
nor U23898 (N_23898,N_15489,N_14033);
or U23899 (N_23899,N_14249,N_14162);
or U23900 (N_23900,N_14576,N_19850);
xnor U23901 (N_23901,N_11542,N_13531);
nor U23902 (N_23902,N_10895,N_11694);
nand U23903 (N_23903,N_15909,N_19123);
nand U23904 (N_23904,N_12600,N_17328);
and U23905 (N_23905,N_10844,N_14991);
or U23906 (N_23906,N_11922,N_17823);
nor U23907 (N_23907,N_17727,N_10653);
and U23908 (N_23908,N_19621,N_11453);
or U23909 (N_23909,N_19077,N_18072);
and U23910 (N_23910,N_17302,N_18684);
and U23911 (N_23911,N_17580,N_16456);
nor U23912 (N_23912,N_11481,N_18390);
xnor U23913 (N_23913,N_12344,N_18597);
or U23914 (N_23914,N_11444,N_14161);
nor U23915 (N_23915,N_12643,N_10105);
xor U23916 (N_23916,N_19050,N_14234);
and U23917 (N_23917,N_16210,N_17609);
and U23918 (N_23918,N_13499,N_11445);
or U23919 (N_23919,N_14295,N_13398);
and U23920 (N_23920,N_13400,N_18231);
nand U23921 (N_23921,N_16406,N_15655);
nor U23922 (N_23922,N_19032,N_16590);
or U23923 (N_23923,N_12425,N_15704);
nand U23924 (N_23924,N_11134,N_15413);
nor U23925 (N_23925,N_19102,N_14895);
or U23926 (N_23926,N_18610,N_14200);
nand U23927 (N_23927,N_13919,N_19025);
or U23928 (N_23928,N_15615,N_18329);
nor U23929 (N_23929,N_10562,N_10359);
or U23930 (N_23930,N_15355,N_10154);
nor U23931 (N_23931,N_19255,N_14532);
xnor U23932 (N_23932,N_11492,N_10257);
and U23933 (N_23933,N_11617,N_11556);
nand U23934 (N_23934,N_11673,N_12493);
nor U23935 (N_23935,N_15172,N_17184);
nand U23936 (N_23936,N_14645,N_11034);
nor U23937 (N_23937,N_18320,N_14423);
nor U23938 (N_23938,N_19279,N_14818);
nor U23939 (N_23939,N_10317,N_13207);
or U23940 (N_23940,N_16048,N_12409);
nand U23941 (N_23941,N_15241,N_15936);
and U23942 (N_23942,N_15652,N_16701);
and U23943 (N_23943,N_13644,N_15501);
nor U23944 (N_23944,N_12621,N_17423);
or U23945 (N_23945,N_19709,N_13108);
nand U23946 (N_23946,N_16867,N_16720);
nand U23947 (N_23947,N_11397,N_11997);
and U23948 (N_23948,N_16816,N_10817);
and U23949 (N_23949,N_19717,N_14167);
nor U23950 (N_23950,N_17162,N_17976);
or U23951 (N_23951,N_12901,N_10744);
and U23952 (N_23952,N_14468,N_17032);
and U23953 (N_23953,N_17846,N_16952);
nand U23954 (N_23954,N_16027,N_13971);
xor U23955 (N_23955,N_12638,N_11186);
nand U23956 (N_23956,N_11748,N_12530);
nand U23957 (N_23957,N_19373,N_17821);
nand U23958 (N_23958,N_13335,N_16312);
or U23959 (N_23959,N_18944,N_10115);
and U23960 (N_23960,N_11793,N_13544);
or U23961 (N_23961,N_13155,N_12742);
nor U23962 (N_23962,N_15846,N_17788);
and U23963 (N_23963,N_11906,N_11955);
nor U23964 (N_23964,N_11669,N_19069);
or U23965 (N_23965,N_16715,N_13268);
or U23966 (N_23966,N_17504,N_11021);
or U23967 (N_23967,N_16449,N_14816);
or U23968 (N_23968,N_18934,N_11963);
nand U23969 (N_23969,N_18914,N_12710);
and U23970 (N_23970,N_11185,N_19487);
nor U23971 (N_23971,N_12025,N_12376);
or U23972 (N_23972,N_17628,N_10886);
nor U23973 (N_23973,N_10606,N_16154);
or U23974 (N_23974,N_12404,N_10678);
or U23975 (N_23975,N_18348,N_15394);
xnor U23976 (N_23976,N_10241,N_11404);
or U23977 (N_23977,N_10790,N_10885);
and U23978 (N_23978,N_14251,N_16574);
nand U23979 (N_23979,N_11752,N_10033);
or U23980 (N_23980,N_10925,N_13978);
or U23981 (N_23981,N_17012,N_19145);
nor U23982 (N_23982,N_16218,N_10901);
nand U23983 (N_23983,N_11150,N_14010);
nor U23984 (N_23984,N_10642,N_17407);
and U23985 (N_23985,N_15320,N_14419);
nor U23986 (N_23986,N_19727,N_14859);
nand U23987 (N_23987,N_11965,N_12158);
and U23988 (N_23988,N_19601,N_15572);
xnor U23989 (N_23989,N_12273,N_16649);
nor U23990 (N_23990,N_12596,N_15738);
nor U23991 (N_23991,N_16174,N_12312);
or U23992 (N_23992,N_18987,N_17024);
and U23993 (N_23993,N_15187,N_15729);
and U23994 (N_23994,N_16623,N_12568);
or U23995 (N_23995,N_12435,N_13564);
nor U23996 (N_23996,N_12959,N_14074);
and U23997 (N_23997,N_15310,N_12883);
nand U23998 (N_23998,N_19220,N_12998);
nor U23999 (N_23999,N_11170,N_15515);
or U24000 (N_24000,N_19835,N_11059);
and U24001 (N_24001,N_11893,N_11942);
and U24002 (N_24002,N_11290,N_15198);
and U24003 (N_24003,N_17090,N_16256);
nand U24004 (N_24004,N_17086,N_19774);
and U24005 (N_24005,N_16995,N_11715);
xnor U24006 (N_24006,N_17589,N_12595);
and U24007 (N_24007,N_14620,N_18429);
or U24008 (N_24008,N_19239,N_17916);
xor U24009 (N_24009,N_15601,N_14959);
nand U24010 (N_24010,N_12583,N_14338);
nor U24011 (N_24011,N_11938,N_13367);
nand U24012 (N_24012,N_10416,N_14695);
and U24013 (N_24013,N_11736,N_17389);
nand U24014 (N_24014,N_19689,N_10759);
and U24015 (N_24015,N_13187,N_14958);
nor U24016 (N_24016,N_18852,N_15815);
nand U24017 (N_24017,N_17509,N_16080);
xnor U24018 (N_24018,N_17313,N_12106);
nand U24019 (N_24019,N_17853,N_18828);
or U24020 (N_24020,N_15920,N_13329);
and U24021 (N_24021,N_17655,N_12662);
or U24022 (N_24022,N_19560,N_17824);
and U24023 (N_24023,N_18144,N_10030);
nand U24024 (N_24024,N_14376,N_10106);
or U24025 (N_24025,N_15826,N_14212);
nand U24026 (N_24026,N_12549,N_14385);
nor U24027 (N_24027,N_14672,N_15772);
nor U24028 (N_24028,N_19265,N_16398);
nand U24029 (N_24029,N_10180,N_13489);
nand U24030 (N_24030,N_17046,N_14513);
and U24031 (N_24031,N_13596,N_12682);
or U24032 (N_24032,N_19804,N_15237);
or U24033 (N_24033,N_18037,N_14413);
and U24034 (N_24034,N_14140,N_19331);
and U24035 (N_24035,N_18245,N_14660);
nor U24036 (N_24036,N_17558,N_11447);
nor U24037 (N_24037,N_13250,N_13299);
nor U24038 (N_24038,N_11686,N_17151);
or U24039 (N_24039,N_10461,N_15381);
or U24040 (N_24040,N_19334,N_10202);
xnor U24041 (N_24041,N_16278,N_18036);
and U24042 (N_24042,N_18440,N_19056);
and U24043 (N_24043,N_11530,N_13467);
nor U24044 (N_24044,N_13916,N_17857);
nor U24045 (N_24045,N_17131,N_17642);
or U24046 (N_24046,N_19144,N_14640);
or U24047 (N_24047,N_15631,N_18151);
or U24048 (N_24048,N_16025,N_10639);
nor U24049 (N_24049,N_16075,N_18287);
nand U24050 (N_24050,N_12212,N_14687);
nor U24051 (N_24051,N_12144,N_16961);
or U24052 (N_24052,N_10103,N_12729);
nand U24053 (N_24053,N_19117,N_16779);
or U24054 (N_24054,N_10081,N_14172);
or U24055 (N_24055,N_18966,N_17971);
and U24056 (N_24056,N_15424,N_18098);
nor U24057 (N_24057,N_19915,N_18162);
and U24058 (N_24058,N_12658,N_15897);
xor U24059 (N_24059,N_13305,N_14185);
and U24060 (N_24060,N_16729,N_18248);
xor U24061 (N_24061,N_14872,N_18250);
xnor U24062 (N_24062,N_15271,N_15377);
or U24063 (N_24063,N_14336,N_10595);
nor U24064 (N_24064,N_10865,N_13356);
and U24065 (N_24065,N_15488,N_18952);
xor U24066 (N_24066,N_18623,N_18940);
and U24067 (N_24067,N_15529,N_16845);
nand U24068 (N_24068,N_17530,N_13079);
nand U24069 (N_24069,N_15000,N_10760);
nor U24070 (N_24070,N_10750,N_17619);
nand U24071 (N_24071,N_16399,N_16607);
and U24072 (N_24072,N_19361,N_12074);
nor U24073 (N_24073,N_18232,N_12576);
or U24074 (N_24074,N_17094,N_14411);
or U24075 (N_24075,N_17830,N_10271);
nor U24076 (N_24076,N_19308,N_18187);
or U24077 (N_24077,N_10737,N_14239);
nor U24078 (N_24078,N_10949,N_13569);
nand U24079 (N_24079,N_17883,N_14915);
nand U24080 (N_24080,N_13269,N_18436);
or U24081 (N_24081,N_19188,N_10958);
nor U24082 (N_24082,N_13714,N_13786);
nand U24083 (N_24083,N_16333,N_14578);
nor U24084 (N_24084,N_19975,N_18306);
nor U24085 (N_24085,N_11425,N_17796);
nand U24086 (N_24086,N_18357,N_16148);
or U24087 (N_24087,N_15003,N_13138);
and U24088 (N_24088,N_17755,N_14591);
nand U24089 (N_24089,N_15434,N_16757);
or U24090 (N_24090,N_19650,N_15286);
nand U24091 (N_24091,N_16671,N_11390);
or U24092 (N_24092,N_12114,N_17826);
nand U24093 (N_24093,N_18859,N_14723);
xor U24094 (N_24094,N_12129,N_18525);
and U24095 (N_24095,N_15563,N_10946);
or U24096 (N_24096,N_13586,N_16766);
or U24097 (N_24097,N_11228,N_16826);
and U24098 (N_24098,N_17181,N_14864);
or U24099 (N_24099,N_11385,N_11433);
nand U24100 (N_24100,N_13533,N_16730);
or U24101 (N_24101,N_18560,N_19394);
nor U24102 (N_24102,N_15171,N_14568);
nand U24103 (N_24103,N_19597,N_18403);
or U24104 (N_24104,N_19982,N_10508);
nand U24105 (N_24105,N_19624,N_16311);
xnor U24106 (N_24106,N_14504,N_17183);
nor U24107 (N_24107,N_10216,N_11581);
or U24108 (N_24108,N_14941,N_13348);
or U24109 (N_24109,N_16377,N_18658);
nand U24110 (N_24110,N_11527,N_11674);
nor U24111 (N_24111,N_12709,N_19329);
and U24112 (N_24112,N_17438,N_19147);
nand U24113 (N_24113,N_15745,N_17048);
xor U24114 (N_24114,N_12842,N_11197);
and U24115 (N_24115,N_11782,N_13654);
or U24116 (N_24116,N_18244,N_18923);
and U24117 (N_24117,N_14743,N_16727);
or U24118 (N_24118,N_10687,N_13699);
nand U24119 (N_24119,N_11394,N_18065);
and U24120 (N_24120,N_18000,N_10219);
xnor U24121 (N_24121,N_17907,N_19826);
nor U24122 (N_24122,N_16260,N_15613);
xnor U24123 (N_24123,N_15102,N_14896);
nor U24124 (N_24124,N_19326,N_12666);
or U24125 (N_24125,N_10032,N_19064);
nand U24126 (N_24126,N_18764,N_19558);
and U24127 (N_24127,N_17070,N_13830);
or U24128 (N_24128,N_14629,N_12422);
xor U24129 (N_24129,N_11724,N_13730);
or U24130 (N_24130,N_11873,N_11286);
nor U24131 (N_24131,N_14319,N_17262);
or U24132 (N_24132,N_13553,N_13160);
or U24133 (N_24133,N_13130,N_13316);
nand U24134 (N_24134,N_19177,N_17110);
nand U24135 (N_24135,N_18678,N_17736);
or U24136 (N_24136,N_19518,N_11642);
xnor U24137 (N_24137,N_18017,N_17373);
nand U24138 (N_24138,N_17535,N_11882);
and U24139 (N_24139,N_14664,N_13302);
nand U24140 (N_24140,N_19389,N_14412);
nor U24141 (N_24141,N_16870,N_10679);
or U24142 (N_24142,N_16964,N_13754);
nor U24143 (N_24143,N_11377,N_14348);
nand U24144 (N_24144,N_17519,N_11159);
nand U24145 (N_24145,N_10251,N_10375);
or U24146 (N_24146,N_19201,N_18173);
nand U24147 (N_24147,N_13758,N_14728);
nand U24148 (N_24148,N_12225,N_11467);
or U24149 (N_24149,N_12577,N_12355);
nor U24150 (N_24150,N_15804,N_12181);
nor U24151 (N_24151,N_10079,N_15805);
and U24152 (N_24152,N_14980,N_19516);
or U24153 (N_24153,N_16833,N_17626);
xor U24154 (N_24154,N_10303,N_15408);
and U24155 (N_24155,N_17372,N_18767);
and U24156 (N_24156,N_19562,N_15332);
nand U24157 (N_24157,N_13438,N_14928);
or U24158 (N_24158,N_16985,N_16789);
and U24159 (N_24159,N_14893,N_12329);
and U24160 (N_24160,N_12325,N_18808);
and U24161 (N_24161,N_17104,N_19174);
or U24162 (N_24162,N_11902,N_14936);
nand U24163 (N_24163,N_12492,N_15946);
nand U24164 (N_24164,N_11146,N_14392);
nand U24165 (N_24165,N_18482,N_17592);
or U24166 (N_24166,N_11865,N_12305);
nor U24167 (N_24167,N_14343,N_16024);
and U24168 (N_24168,N_15450,N_10485);
xor U24169 (N_24169,N_17329,N_19014);
nor U24170 (N_24170,N_18107,N_17227);
or U24171 (N_24171,N_16265,N_16935);
and U24172 (N_24172,N_17029,N_18015);
or U24173 (N_24173,N_11551,N_10554);
or U24174 (N_24174,N_15992,N_14166);
xor U24175 (N_24175,N_18149,N_11946);
and U24176 (N_24176,N_15531,N_11638);
or U24177 (N_24177,N_15932,N_17417);
nor U24178 (N_24178,N_19459,N_12160);
or U24179 (N_24179,N_17009,N_10459);
or U24180 (N_24180,N_16909,N_11562);
xnor U24181 (N_24181,N_14134,N_17387);
nor U24182 (N_24182,N_19991,N_13837);
and U24183 (N_24183,N_15329,N_17011);
or U24184 (N_24184,N_14493,N_15838);
nand U24185 (N_24185,N_18724,N_13931);
nor U24186 (N_24186,N_11378,N_15973);
nor U24187 (N_24187,N_16494,N_18804);
or U24188 (N_24188,N_18341,N_17926);
nor U24189 (N_24189,N_10996,N_11980);
or U24190 (N_24190,N_11489,N_14356);
nand U24191 (N_24191,N_13797,N_15111);
and U24192 (N_24192,N_10530,N_10713);
nand U24193 (N_24193,N_19285,N_17640);
or U24194 (N_24194,N_14263,N_12508);
or U24195 (N_24195,N_15849,N_12848);
nand U24196 (N_24196,N_12454,N_12562);
and U24197 (N_24197,N_13312,N_10926);
or U24198 (N_24198,N_17749,N_18760);
or U24199 (N_24199,N_17921,N_16982);
nand U24200 (N_24200,N_15004,N_10069);
xor U24201 (N_24201,N_15550,N_19720);
and U24202 (N_24202,N_15232,N_10176);
nor U24203 (N_24203,N_19093,N_15599);
or U24204 (N_24204,N_19921,N_13704);
or U24205 (N_24205,N_15278,N_19997);
or U24206 (N_24206,N_19190,N_12930);
and U24207 (N_24207,N_16338,N_11476);
or U24208 (N_24208,N_11005,N_16555);
and U24209 (N_24209,N_11260,N_11746);
and U24210 (N_24210,N_18382,N_13985);
nor U24211 (N_24211,N_12632,N_19465);
or U24212 (N_24212,N_13111,N_14686);
and U24213 (N_24213,N_19496,N_10794);
or U24214 (N_24214,N_16478,N_16724);
or U24215 (N_24215,N_19095,N_15876);
nor U24216 (N_24216,N_10072,N_11602);
nor U24217 (N_24217,N_12141,N_18242);
or U24218 (N_24218,N_12477,N_15913);
and U24219 (N_24219,N_16267,N_16840);
and U24220 (N_24220,N_15063,N_18282);
nor U24221 (N_24221,N_15713,N_14261);
nor U24222 (N_24222,N_19137,N_11868);
nor U24223 (N_24223,N_12791,N_14045);
and U24224 (N_24224,N_19992,N_13301);
and U24225 (N_24225,N_13336,N_12745);
or U24226 (N_24226,N_12230,N_18008);
nor U24227 (N_24227,N_14209,N_14136);
nor U24228 (N_24228,N_15277,N_11615);
or U24229 (N_24229,N_17508,N_18521);
nor U24230 (N_24230,N_16028,N_13813);
or U24231 (N_24231,N_16283,N_19096);
nor U24232 (N_24232,N_11929,N_19584);
or U24233 (N_24233,N_17209,N_12365);
nor U24234 (N_24234,N_15417,N_19864);
nand U24235 (N_24235,N_12056,N_14473);
or U24236 (N_24236,N_17079,N_18667);
or U24237 (N_24237,N_13194,N_16036);
xnor U24238 (N_24238,N_13816,N_16667);
or U24239 (N_24239,N_16834,N_13873);
and U24240 (N_24240,N_17122,N_17441);
xnor U24241 (N_24241,N_10821,N_12626);
or U24242 (N_24242,N_16172,N_13030);
nor U24243 (N_24243,N_15197,N_13337);
nand U24244 (N_24244,N_13327,N_10751);
nand U24245 (N_24245,N_10699,N_15174);
nor U24246 (N_24246,N_14617,N_17832);
xor U24247 (N_24247,N_11585,N_15359);
and U24248 (N_24248,N_15541,N_11888);
xor U24249 (N_24249,N_17386,N_17263);
nand U24250 (N_24250,N_14828,N_14478);
nor U24251 (N_24251,N_14625,N_14273);
xor U24252 (N_24252,N_13123,N_17856);
xor U24253 (N_24253,N_12087,N_13652);
nor U24254 (N_24254,N_19872,N_11533);
nand U24255 (N_24255,N_10237,N_17996);
nor U24256 (N_24256,N_10825,N_15677);
nor U24257 (N_24257,N_13842,N_15576);
or U24258 (N_24258,N_11879,N_13668);
xnor U24259 (N_24259,N_14746,N_13224);
xor U24260 (N_24260,N_12251,N_11137);
or U24261 (N_24261,N_10505,N_12431);
and U24262 (N_24262,N_17003,N_18929);
nor U24263 (N_24263,N_18703,N_14805);
and U24264 (N_24264,N_18792,N_15218);
and U24265 (N_24265,N_13782,N_19240);
xnor U24266 (N_24266,N_16860,N_11494);
nand U24267 (N_24267,N_16847,N_16346);
nor U24268 (N_24268,N_15019,N_16598);
nand U24269 (N_24269,N_12214,N_12175);
xnor U24270 (N_24270,N_19796,N_16450);
nand U24271 (N_24271,N_16977,N_15785);
nor U24272 (N_24272,N_12097,N_10211);
nand U24273 (N_24273,N_10155,N_19396);
and U24274 (N_24274,N_19310,N_11863);
and U24275 (N_24275,N_15311,N_11105);
or U24276 (N_24276,N_13021,N_16353);
nor U24277 (N_24277,N_14878,N_12479);
xor U24278 (N_24278,N_13494,N_17148);
xor U24279 (N_24279,N_14426,N_11456);
nand U24280 (N_24280,N_12100,N_19528);
nor U24281 (N_24281,N_18224,N_18864);
or U24282 (N_24282,N_13658,N_17458);
nor U24283 (N_24283,N_13263,N_11113);
and U24284 (N_24284,N_14042,N_18404);
and U24285 (N_24285,N_15656,N_11981);
nor U24286 (N_24286,N_19746,N_18351);
or U24287 (N_24287,N_14223,N_15049);
nand U24288 (N_24288,N_12488,N_18214);
or U24289 (N_24289,N_14824,N_18073);
and U24290 (N_24290,N_15382,N_10542);
nand U24291 (N_24291,N_13198,N_14965);
or U24292 (N_24292,N_13991,N_17160);
or U24293 (N_24293,N_15813,N_16201);
and U24294 (N_24294,N_19344,N_18532);
nand U24295 (N_24295,N_15023,N_19901);
or U24296 (N_24296,N_19737,N_12342);
nand U24297 (N_24297,N_18154,N_12574);
nor U24298 (N_24298,N_18874,N_15147);
nor U24299 (N_24299,N_14159,N_17917);
or U24300 (N_24300,N_10763,N_16592);
nand U24301 (N_24301,N_14631,N_12622);
or U24302 (N_24302,N_15660,N_12063);
and U24303 (N_24303,N_14569,N_12821);
nand U24304 (N_24304,N_11535,N_16512);
nand U24305 (N_24305,N_13168,N_14538);
nor U24306 (N_24306,N_17940,N_13661);
xnor U24307 (N_24307,N_10831,N_13967);
nand U24308 (N_24308,N_13351,N_11443);
nor U24309 (N_24309,N_16051,N_17343);
nor U24310 (N_24310,N_10412,N_11126);
or U24311 (N_24311,N_18726,N_12992);
or U24312 (N_24312,N_16281,N_11294);
or U24313 (N_24313,N_11417,N_10582);
xnor U24314 (N_24314,N_15985,N_16092);
and U24315 (N_24315,N_17772,N_13753);
and U24316 (N_24316,N_12653,N_12735);
nor U24317 (N_24317,N_15436,N_18479);
nor U24318 (N_24318,N_14914,N_15341);
or U24319 (N_24319,N_10645,N_15621);
xor U24320 (N_24320,N_11124,N_11318);
nor U24321 (N_24321,N_19428,N_15207);
nor U24322 (N_24322,N_15618,N_12388);
and U24323 (N_24323,N_19384,N_10273);
and U24324 (N_24324,N_12285,N_15994);
or U24325 (N_24325,N_14930,N_10807);
nand U24326 (N_24326,N_13509,N_18384);
nand U24327 (N_24327,N_15511,N_12307);
and U24328 (N_24328,N_12465,N_18222);
nor U24329 (N_24329,N_11271,N_12804);
nand U24330 (N_24330,N_14748,N_13085);
nor U24331 (N_24331,N_17449,N_10776);
and U24332 (N_24332,N_12414,N_11381);
xor U24333 (N_24333,N_18343,N_11857);
or U24334 (N_24334,N_16541,N_14111);
nor U24335 (N_24335,N_16173,N_15326);
xor U24336 (N_24336,N_19211,N_10307);
and U24337 (N_24337,N_13515,N_16884);
or U24338 (N_24338,N_13856,N_17813);
and U24339 (N_24339,N_14199,N_18900);
or U24340 (N_24340,N_17425,N_19993);
or U24341 (N_24341,N_12131,N_13110);
and U24342 (N_24342,N_18915,N_11459);
and U24343 (N_24343,N_13029,N_15559);
and U24344 (N_24344,N_10975,N_17191);
nor U24345 (N_24345,N_18691,N_12676);
or U24346 (N_24346,N_12516,N_16198);
and U24347 (N_24347,N_18830,N_13084);
nor U24348 (N_24348,N_17995,N_10250);
nand U24349 (N_24349,N_15776,N_17804);
and U24350 (N_24350,N_16930,N_17371);
and U24351 (N_24351,N_15614,N_15811);
xnor U24352 (N_24352,N_13885,N_16429);
or U24353 (N_24353,N_16087,N_19884);
or U24354 (N_24354,N_17064,N_19097);
or U24355 (N_24355,N_13013,N_15478);
nor U24356 (N_24356,N_14135,N_11219);
nand U24357 (N_24357,N_15078,N_12287);
nor U24358 (N_24358,N_11892,N_18274);
and U24359 (N_24359,N_19509,N_10243);
or U24360 (N_24360,N_18181,N_16832);
or U24361 (N_24361,N_19155,N_18709);
or U24362 (N_24362,N_19559,N_12391);
and U24363 (N_24363,N_13882,N_11645);
nand U24364 (N_24364,N_13505,N_13607);
nand U24365 (N_24365,N_17841,N_11719);
xor U24366 (N_24366,N_14635,N_16550);
and U24367 (N_24367,N_16907,N_18293);
and U24368 (N_24368,N_11229,N_10797);
or U24369 (N_24369,N_14733,N_11426);
and U24370 (N_24370,N_12059,N_18675);
xnor U24371 (N_24371,N_17700,N_17936);
and U24372 (N_24372,N_15966,N_15347);
nor U24373 (N_24373,N_18857,N_14020);
xnor U24374 (N_24374,N_16022,N_12162);
and U24375 (N_24375,N_12711,N_14682);
nand U24376 (N_24376,N_10522,N_12458);
nand U24377 (N_24377,N_17141,N_10174);
and U24378 (N_24378,N_10723,N_15737);
xnor U24379 (N_24379,N_19652,N_10289);
xnor U24380 (N_24380,N_12732,N_13826);
nor U24381 (N_24381,N_15724,N_13630);
or U24382 (N_24382,N_19863,N_17298);
or U24383 (N_24383,N_17515,N_12771);
nand U24384 (N_24384,N_17276,N_13844);
and U24385 (N_24385,N_19473,N_12094);
nor U24386 (N_24386,N_17953,N_10551);
or U24387 (N_24387,N_18119,N_14563);
and U24388 (N_24388,N_19728,N_17548);
nor U24389 (N_24389,N_13001,N_16263);
nand U24390 (N_24390,N_12096,N_11454);
nor U24391 (N_24391,N_11032,N_10310);
or U24392 (N_24392,N_19333,N_18219);
nor U24393 (N_24393,N_15460,N_18695);
or U24394 (N_24394,N_10427,N_18212);
nor U24395 (N_24395,N_15904,N_13674);
nor U24396 (N_24396,N_18456,N_16455);
nor U24397 (N_24397,N_10980,N_13843);
and U24398 (N_24398,N_16782,N_13512);
or U24399 (N_24399,N_15318,N_10585);
and U24400 (N_24400,N_11037,N_15361);
and U24401 (N_24401,N_10676,N_16235);
xnor U24402 (N_24402,N_15643,N_13371);
and U24403 (N_24403,N_11270,N_13476);
nor U24404 (N_24404,N_11966,N_15800);
nor U24405 (N_24405,N_16781,N_13121);
nor U24406 (N_24406,N_15664,N_19301);
nor U24407 (N_24407,N_12579,N_19337);
nor U24408 (N_24408,N_11773,N_11251);
or U24409 (N_24409,N_17121,N_15902);
nor U24410 (N_24410,N_10799,N_18588);
nand U24411 (N_24411,N_16239,N_17190);
nor U24412 (N_24412,N_18011,N_17471);
nand U24413 (N_24413,N_12243,N_19914);
nand U24414 (N_24414,N_11745,N_13620);
and U24415 (N_24415,N_15317,N_12534);
nand U24416 (N_24416,N_11995,N_19166);
or U24417 (N_24417,N_15404,N_13889);
or U24418 (N_24418,N_19747,N_12723);
or U24419 (N_24419,N_17092,N_10692);
xnor U24420 (N_24420,N_10730,N_17097);
xnor U24421 (N_24421,N_16673,N_16908);
nand U24422 (N_24422,N_13924,N_13890);
nand U24423 (N_24423,N_12028,N_16923);
xnor U24424 (N_24424,N_15438,N_12623);
nor U24425 (N_24425,N_15272,N_10226);
or U24426 (N_24426,N_11250,N_10276);
xnor U24427 (N_24427,N_19785,N_14367);
and U24428 (N_24428,N_16731,N_12909);
and U24429 (N_24429,N_15428,N_15809);
or U24430 (N_24430,N_10711,N_11833);
nor U24431 (N_24431,N_12048,N_14406);
or U24432 (N_24432,N_19390,N_16525);
xnor U24433 (N_24433,N_14518,N_13453);
xor U24434 (N_24434,N_10566,N_18992);
nor U24435 (N_24435,N_19143,N_15620);
or U24436 (N_24436,N_18066,N_12333);
and U24437 (N_24437,N_12839,N_14662);
or U24438 (N_24438,N_11007,N_17652);
or U24439 (N_24439,N_15366,N_12758);
nand U24440 (N_24440,N_11411,N_15446);
or U24441 (N_24441,N_10496,N_18501);
nor U24442 (N_24442,N_18204,N_12789);
and U24443 (N_24443,N_13171,N_11047);
xor U24444 (N_24444,N_15062,N_10231);
nand U24445 (N_24445,N_14105,N_12191);
nand U24446 (N_24446,N_11837,N_17555);
or U24447 (N_24447,N_14549,N_14973);
nor U24448 (N_24448,N_19833,N_18901);
and U24449 (N_24449,N_15337,N_18854);
and U24450 (N_24450,N_19315,N_15407);
nor U24451 (N_24451,N_12865,N_16965);
or U24452 (N_24452,N_19057,N_18386);
xor U24453 (N_24453,N_10977,N_15455);
nor U24454 (N_24454,N_13442,N_12311);
nand U24455 (N_24455,N_16125,N_12405);
nand U24456 (N_24456,N_16313,N_14809);
nand U24457 (N_24457,N_16754,N_12224);
nand U24458 (N_24458,N_11038,N_14910);
and U24459 (N_24459,N_11089,N_11161);
and U24460 (N_24460,N_13820,N_14339);
and U24461 (N_24461,N_12206,N_13996);
nor U24462 (N_24462,N_14254,N_18572);
nor U24463 (N_24463,N_17133,N_17786);
or U24464 (N_24464,N_19874,N_15733);
or U24465 (N_24465,N_10928,N_13005);
nor U24466 (N_24466,N_18370,N_14480);
and U24467 (N_24467,N_18998,N_10495);
nand U24468 (N_24468,N_19526,N_13514);
nor U24469 (N_24469,N_11705,N_14170);
or U24470 (N_24470,N_14526,N_14754);
nand U24471 (N_24471,N_12538,N_18152);
nand U24472 (N_24472,N_13142,N_13333);
or U24473 (N_24473,N_16395,N_19382);
or U24474 (N_24474,N_16000,N_12746);
or U24475 (N_24475,N_19263,N_18053);
and U24476 (N_24476,N_14464,N_13637);
and U24477 (N_24477,N_17648,N_17770);
xor U24478 (N_24478,N_15768,N_19192);
or U24479 (N_24479,N_19766,N_11348);
xor U24480 (N_24480,N_10051,N_11777);
nand U24481 (N_24481,N_18963,N_11025);
and U24482 (N_24482,N_16998,N_13104);
and U24483 (N_24483,N_19224,N_19086);
nor U24484 (N_24484,N_16085,N_11641);
xor U24485 (N_24485,N_16951,N_15421);
xnor U24486 (N_24486,N_17858,N_13863);
nor U24487 (N_24487,N_15506,N_11904);
nor U24488 (N_24488,N_18942,N_10493);
and U24489 (N_24489,N_12487,N_13319);
nand U24490 (N_24490,N_19849,N_11780);
and U24491 (N_24491,N_10308,N_19140);
and U24492 (N_24492,N_10408,N_10299);
or U24493 (N_24493,N_11749,N_13332);
and U24494 (N_24494,N_11022,N_19152);
and U24495 (N_24495,N_12430,N_15058);
xor U24496 (N_24496,N_17206,N_10442);
nand U24497 (N_24497,N_19418,N_12238);
nand U24498 (N_24498,N_11739,N_14059);
nor U24499 (N_24499,N_16903,N_18023);
nand U24500 (N_24500,N_10686,N_18388);
xor U24501 (N_24501,N_17888,N_13420);
or U24502 (N_24502,N_12187,N_17705);
nand U24503 (N_24503,N_14248,N_17267);
or U24504 (N_24504,N_12511,N_15022);
nor U24505 (N_24505,N_10519,N_19837);
or U24506 (N_24506,N_15610,N_12429);
xor U24507 (N_24507,N_13974,N_11619);
or U24508 (N_24508,N_13561,N_19432);
nand U24509 (N_24509,N_14988,N_13264);
and U24510 (N_24510,N_14627,N_18239);
xnor U24511 (N_24511,N_16501,N_11772);
nor U24512 (N_24512,N_14866,N_15390);
or U24513 (N_24513,N_18867,N_13245);
nor U24514 (N_24514,N_11287,N_11094);
nand U24515 (N_24515,N_10548,N_17561);
xor U24516 (N_24516,N_16008,N_19870);
or U24517 (N_24517,N_14832,N_18186);
xor U24518 (N_24518,N_16984,N_12364);
nor U24519 (N_24519,N_17200,N_15949);
xor U24520 (N_24520,N_12605,N_17307);
and U24521 (N_24521,N_12260,N_12400);
or U24522 (N_24522,N_12916,N_10899);
nand U24523 (N_24523,N_19156,N_11054);
and U24524 (N_24524,N_19332,N_18010);
and U24525 (N_24525,N_14143,N_11338);
nand U24526 (N_24526,N_11805,N_13091);
or U24527 (N_24527,N_14944,N_12531);
nand U24528 (N_24528,N_16835,N_11432);
nand U24529 (N_24529,N_11582,N_18554);
and U24530 (N_24530,N_18961,N_19313);
nand U24531 (N_24531,N_17822,N_10784);
nor U24532 (N_24532,N_16502,N_12288);
and U24533 (N_24533,N_10426,N_12334);
and U24534 (N_24534,N_12680,N_18637);
and U24535 (N_24535,N_17294,N_17314);
or U24536 (N_24536,N_14041,N_12740);
nand U24537 (N_24537,N_18654,N_13691);
xor U24538 (N_24538,N_10085,N_18844);
or U24539 (N_24539,N_19527,N_15193);
or U24540 (N_24540,N_18569,N_11218);
or U24541 (N_24541,N_10836,N_10016);
or U24542 (N_24542,N_13693,N_12481);
or U24543 (N_24543,N_10326,N_10089);
or U24544 (N_24544,N_17108,N_15861);
or U24545 (N_24545,N_14107,N_19607);
or U24546 (N_24546,N_13096,N_15229);
nor U24547 (N_24547,N_11722,N_13244);
and U24548 (N_24548,N_13261,N_15673);
xor U24549 (N_24549,N_12235,N_19694);
or U24550 (N_24550,N_10719,N_16863);
nand U24551 (N_24551,N_19994,N_12999);
nor U24552 (N_24552,N_17460,N_15726);
or U24553 (N_24553,N_19771,N_14755);
nand U24554 (N_24554,N_17082,N_11132);
nand U24555 (N_24555,N_17728,N_16665);
or U24556 (N_24556,N_10161,N_11650);
nand U24557 (N_24557,N_11731,N_18636);
and U24558 (N_24558,N_10207,N_13285);
or U24559 (N_24559,N_16911,N_19071);
and U24560 (N_24560,N_17042,N_12522);
and U24561 (N_24561,N_19229,N_18294);
nand U24562 (N_24562,N_15594,N_12316);
or U24563 (N_24563,N_19135,N_11230);
or U24564 (N_24564,N_15893,N_17529);
nand U24565 (N_24565,N_19464,N_13144);
and U24566 (N_24566,N_11412,N_15898);
or U24567 (N_24567,N_15886,N_10874);
or U24568 (N_24568,N_15600,N_17545);
nor U24569 (N_24569,N_19075,N_11753);
nor U24570 (N_24570,N_11889,N_16058);
and U24571 (N_24571,N_12841,N_14279);
or U24572 (N_24572,N_15608,N_13026);
nor U24573 (N_24573,N_13576,N_18240);
nor U24574 (N_24574,N_19807,N_11414);
or U24575 (N_24575,N_10262,N_11472);
or U24576 (N_24576,N_18668,N_12727);
and U24577 (N_24577,N_16631,N_10883);
or U24578 (N_24578,N_13237,N_12898);
and U24579 (N_24579,N_16005,N_16184);
and U24580 (N_24580,N_18067,N_16073);
nand U24581 (N_24581,N_12453,N_19412);
nand U24582 (N_24582,N_13501,N_11189);
and U24583 (N_24583,N_14646,N_10351);
or U24584 (N_24584,N_16472,N_13810);
and U24585 (N_24585,N_16810,N_10754);
nand U24586 (N_24586,N_19008,N_18164);
xor U24587 (N_24587,N_17715,N_19183);
nor U24588 (N_24588,N_12884,N_13636);
or U24589 (N_24589,N_17549,N_14186);
and U24590 (N_24590,N_19358,N_18772);
and U24591 (N_24591,N_12215,N_15798);
nand U24592 (N_24592,N_18640,N_12283);
nor U24593 (N_24593,N_10573,N_19936);
nor U24594 (N_24594,N_12637,N_14311);
xnor U24595 (N_24595,N_17146,N_16060);
or U24596 (N_24596,N_13545,N_15142);
nor U24597 (N_24597,N_16414,N_13532);
xnor U24598 (N_24598,N_19298,N_13188);
nand U24599 (N_24599,N_15554,N_11999);
nand U24600 (N_24600,N_15636,N_10148);
nor U24601 (N_24601,N_11496,N_13128);
or U24602 (N_24602,N_12090,N_19831);
or U24603 (N_24603,N_12194,N_17540);
or U24604 (N_24604,N_12755,N_11003);
or U24605 (N_24605,N_14786,N_14601);
nand U24606 (N_24606,N_12010,N_15351);
nor U24607 (N_24607,N_18203,N_17169);
nor U24608 (N_24608,N_15574,N_16039);
and U24609 (N_24609,N_17334,N_14539);
or U24610 (N_24610,N_13728,N_12200);
xor U24611 (N_24611,N_11670,N_17374);
or U24612 (N_24612,N_15819,N_11167);
nor U24613 (N_24613,N_12827,N_19617);
or U24614 (N_24614,N_10491,N_13994);
nand U24615 (N_24615,N_19780,N_15261);
or U24616 (N_24616,N_14429,N_11522);
nand U24617 (N_24617,N_19469,N_16749);
xnor U24618 (N_24618,N_16336,N_17385);
or U24619 (N_24619,N_10826,N_13886);
or U24620 (N_24620,N_15401,N_16093);
and U24621 (N_24621,N_18725,N_10866);
or U24622 (N_24622,N_17799,N_12504);
and U24623 (N_24623,N_15242,N_11152);
and U24624 (N_24624,N_18377,N_18491);
or U24625 (N_24625,N_11352,N_13883);
and U24626 (N_24626,N_14021,N_14204);
or U24627 (N_24627,N_14842,N_17735);
and U24628 (N_24628,N_17462,N_19023);
nor U24629 (N_24629,N_11245,N_14024);
nand U24630 (N_24630,N_12679,N_19569);
nor U24631 (N_24631,N_13421,N_11060);
or U24632 (N_24632,N_18848,N_16941);
and U24633 (N_24633,N_12683,N_13487);
nand U24634 (N_24634,N_10233,N_11278);
and U24635 (N_24635,N_14379,N_18833);
or U24636 (N_24636,N_19058,N_12418);
and U24637 (N_24637,N_15300,N_13648);
or U24638 (N_24638,N_16805,N_19546);
nand U24639 (N_24639,N_16772,N_10514);
or U24640 (N_24640,N_19302,N_10933);
xnor U24641 (N_24641,N_15178,N_15775);
and U24642 (N_24642,N_19049,N_18176);
nand U24643 (N_24643,N_15236,N_12890);
or U24644 (N_24644,N_14256,N_11080);
and U24645 (N_24645,N_18182,N_17306);
and U24646 (N_24646,N_10462,N_17694);
and U24647 (N_24647,N_17264,N_15126);
or U24648 (N_24648,N_19827,N_16802);
nor U24649 (N_24649,N_15391,N_13705);
and U24650 (N_24650,N_18599,N_12104);
nand U24651 (N_24651,N_13430,N_14349);
nor U24652 (N_24652,N_19482,N_14540);
and U24653 (N_24653,N_13633,N_15153);
and U24654 (N_24654,N_15842,N_11099);
and U24655 (N_24655,N_12586,N_16091);
xor U24656 (N_24656,N_12000,N_14548);
xor U24657 (N_24657,N_12475,N_17170);
nand U24658 (N_24658,N_12029,N_17336);
or U24659 (N_24659,N_14611,N_19908);
and U24660 (N_24660,N_12143,N_10045);
and U24661 (N_24661,N_11778,N_16389);
nand U24662 (N_24662,N_15935,N_16416);
or U24663 (N_24663,N_17714,N_13541);
nand U24664 (N_24664,N_16993,N_17702);
and U24665 (N_24665,N_18088,N_12905);
and U24666 (N_24666,N_14583,N_16593);
nor U24667 (N_24667,N_16796,N_12353);
nand U24668 (N_24668,N_12482,N_14126);
nand U24669 (N_24669,N_11345,N_12024);
nor U24670 (N_24670,N_15309,N_13277);
nand U24671 (N_24671,N_14711,N_10544);
and U24672 (N_24672,N_14421,N_15012);
nand U24673 (N_24673,N_16104,N_18960);
nand U24674 (N_24674,N_16341,N_17724);
and U24675 (N_24675,N_13158,N_18673);
or U24676 (N_24676,N_10785,N_11462);
or U24677 (N_24677,N_14788,N_14362);
nor U24678 (N_24678,N_12984,N_11802);
or U24679 (N_24679,N_15582,N_14277);
nand U24680 (N_24680,N_14484,N_10990);
and U24681 (N_24681,N_17762,N_18297);
and U24682 (N_24682,N_16803,N_10342);
nand U24683 (N_24683,N_11621,N_18427);
nor U24684 (N_24684,N_17224,N_19736);
and U24685 (N_24685,N_11006,N_16519);
xor U24686 (N_24686,N_13139,N_12690);
nor U24687 (N_24687,N_14575,N_11666);
or U24688 (N_24688,N_18576,N_10407);
xnor U24689 (N_24689,N_18087,N_11438);
nor U24690 (N_24690,N_13447,N_14097);
or U24691 (N_24691,N_19940,N_10900);
or U24692 (N_24692,N_14950,N_10093);
nand U24693 (N_24693,N_12363,N_16458);
and U24694 (N_24694,N_10635,N_19956);
or U24695 (N_24695,N_16342,N_19307);
or U24696 (N_24696,N_19918,N_13397);
nor U24697 (N_24697,N_14632,N_10004);
or U24698 (N_24698,N_15283,N_15244);
nor U24699 (N_24699,N_15180,N_12661);
and U24700 (N_24700,N_16303,N_18309);
or U24701 (N_24701,N_15841,N_11102);
or U24702 (N_24702,N_13070,N_17898);
and U24703 (N_24703,N_11191,N_10559);
nand U24704 (N_24704,N_17537,N_18424);
nor U24705 (N_24705,N_19324,N_14798);
xnor U24706 (N_24706,N_13242,N_14117);
or U24707 (N_24707,N_12943,N_18697);
nand U24708 (N_24708,N_13616,N_19476);
and U24709 (N_24709,N_15797,N_10685);
and U24710 (N_24710,N_17410,N_16102);
nand U24711 (N_24711,N_18249,N_18566);
nor U24712 (N_24712,N_17653,N_19675);
nor U24713 (N_24713,N_16364,N_12227);
nor U24714 (N_24714,N_11925,N_15503);
xor U24715 (N_24715,N_19001,N_18234);
nor U24716 (N_24716,N_13713,N_15824);
or U24717 (N_24717,N_16468,N_18194);
nand U24718 (N_24718,N_13055,N_15494);
or U24719 (N_24719,N_19769,N_18976);
and U24720 (N_24720,N_10240,N_16934);
or U24721 (N_24721,N_15839,N_15648);
nor U24722 (N_24722,N_11620,N_17055);
or U24723 (N_24723,N_18400,N_11329);
nand U24724 (N_24724,N_16793,N_15032);
and U24725 (N_24725,N_13905,N_10255);
xnor U24726 (N_24726,N_10122,N_16434);
xor U24727 (N_24727,N_12343,N_12611);
nor U24728 (N_24728,N_13134,N_10786);
nand U24729 (N_24729,N_19457,N_10381);
and U24730 (N_24730,N_10121,N_18627);
nor U24731 (N_24731,N_17231,N_14358);
xor U24732 (N_24732,N_15577,N_10166);
xnor U24733 (N_24733,N_13678,N_11688);
nand U24734 (N_24734,N_19413,N_18362);
xnor U24735 (N_24735,N_16654,N_12862);
and U24736 (N_24736,N_19223,N_12967);
nor U24737 (N_24737,N_18731,N_14293);
nor U24738 (N_24738,N_13478,N_10313);
nand U24739 (N_24739,N_11488,N_13227);
or U24740 (N_24740,N_11800,N_18120);
and U24741 (N_24741,N_19417,N_14491);
and U24742 (N_24742,N_13095,N_13858);
or U24743 (N_24743,N_19348,N_14644);
nand U24744 (N_24744,N_12618,N_18056);
xnor U24745 (N_24745,N_14913,N_11319);
and U24746 (N_24746,N_16743,N_19235);
xor U24747 (N_24747,N_16708,N_14164);
nor U24748 (N_24748,N_19957,N_15416);
or U24749 (N_24749,N_17861,N_17367);
nand U24750 (N_24750,N_16866,N_15794);
and U24751 (N_24751,N_13761,N_18997);
nor U24752 (N_24752,N_18110,N_16299);
xor U24753 (N_24753,N_11640,N_15856);
or U24754 (N_24754,N_11246,N_10478);
nor U24755 (N_24755,N_14196,N_18472);
nand U24756 (N_24756,N_12509,N_16719);
nand U24757 (N_24757,N_17126,N_15963);
and U24758 (N_24758,N_11896,N_12517);
or U24759 (N_24759,N_10168,N_18318);
xnor U24760 (N_24760,N_10334,N_15480);
xor U24761 (N_24761,N_11594,N_15306);
and U24762 (N_24762,N_13407,N_14157);
and U24763 (N_24763,N_19189,N_14246);
nor U24764 (N_24764,N_15076,N_14869);
nand U24765 (N_24765,N_10191,N_10238);
or U24766 (N_24766,N_11068,N_12552);
nor U24767 (N_24767,N_17739,N_12996);
xor U24768 (N_24768,N_17290,N_18138);
or U24769 (N_24769,N_10075,N_16317);
xnor U24770 (N_24770,N_18112,N_11335);
or U24771 (N_24771,N_16643,N_12987);
and U24772 (N_24772,N_14110,N_15490);
or U24773 (N_24773,N_13440,N_11118);
and U24774 (N_24774,N_13923,N_13273);
nor U24775 (N_24775,N_15378,N_14294);
xor U24776 (N_24776,N_13739,N_12480);
and U24777 (N_24777,N_19803,N_10283);
and U24778 (N_24778,N_14725,N_18168);
nor U24779 (N_24779,N_17008,N_13457);
nor U24780 (N_24780,N_11860,N_12037);
and U24781 (N_24781,N_12655,N_13340);
nor U24782 (N_24782,N_16751,N_14290);
or U24783 (N_24783,N_15484,N_18160);
and U24784 (N_24784,N_19877,N_12756);
and U24785 (N_24785,N_16532,N_19937);
or U24786 (N_24786,N_13631,N_16422);
nand U24787 (N_24787,N_14165,N_13212);
and U24788 (N_24788,N_18989,N_11194);
nor U24789 (N_24789,N_11362,N_10837);
or U24790 (N_24790,N_16690,N_13507);
or U24791 (N_24791,N_18642,N_17219);
xnor U24792 (N_24792,N_15736,N_10039);
nand U24793 (N_24793,N_17769,N_17424);
and U24794 (N_24794,N_12064,N_12491);
and U24795 (N_24795,N_18771,N_14978);
nand U24796 (N_24796,N_12975,N_11010);
nand U24797 (N_24797,N_17140,N_15633);
or U24798 (N_24798,N_13044,N_12150);
or U24799 (N_24799,N_14997,N_14948);
nor U24800 (N_24800,N_13855,N_12603);
and U24801 (N_24801,N_12189,N_10565);
nand U24802 (N_24802,N_14070,N_18911);
and U24803 (N_24803,N_16268,N_12462);
nand U24804 (N_24804,N_18556,N_17332);
and U24805 (N_24805,N_17043,N_16544);
and U24806 (N_24806,N_10637,N_17044);
nor U24807 (N_24807,N_13262,N_15828);
and U24808 (N_24808,N_13998,N_16397);
nand U24809 (N_24809,N_14201,N_16531);
nor U24810 (N_24810,N_13032,N_15555);
nor U24811 (N_24811,N_17235,N_18905);
nor U24812 (N_24812,N_12115,N_15331);
or U24813 (N_24813,N_18132,N_11083);
or U24814 (N_24814,N_13565,N_13054);
nor U24815 (N_24815,N_11215,N_10124);
nand U24816 (N_24816,N_15130,N_11733);
and U24817 (N_24817,N_19080,N_10298);
nor U24818 (N_24818,N_14642,N_13716);
nor U24819 (N_24819,N_17759,N_17340);
and U24820 (N_24820,N_15228,N_12744);
nand U24821 (N_24821,N_14667,N_15524);
nor U24822 (N_24822,N_10280,N_17061);
nor U24823 (N_24823,N_14287,N_12734);
and U24824 (N_24824,N_18383,N_16915);
and U24825 (N_24825,N_14880,N_18083);
nor U24826 (N_24826,N_11331,N_11202);
nand U24827 (N_24827,N_14870,N_19295);
nor U24828 (N_24828,N_14665,N_14371);
nor U24829 (N_24829,N_11680,N_12598);
or U24830 (N_24830,N_12790,N_11255);
nor U24831 (N_24831,N_15818,N_13958);
and U24832 (N_24832,N_15834,N_10896);
nand U24833 (N_24833,N_11985,N_11356);
nor U24834 (N_24834,N_10888,N_19571);
and U24835 (N_24835,N_12856,N_11933);
nand U24836 (N_24836,N_12272,N_13088);
and U24837 (N_24837,N_15702,N_15540);
and U24838 (N_24838,N_15068,N_11740);
nand U24839 (N_24839,N_14054,N_12851);
xnor U24840 (N_24840,N_13587,N_19228);
and U24841 (N_24841,N_11979,N_18896);
or U24842 (N_24842,N_10643,N_10242);
nor U24843 (N_24843,N_19010,N_13230);
or U24844 (N_24844,N_11464,N_12903);
nand U24845 (N_24845,N_13671,N_15562);
nor U24846 (N_24846,N_14039,N_18426);
or U24847 (N_24847,N_12988,N_17134);
and U24848 (N_24848,N_15791,N_10905);
nand U24849 (N_24849,N_18991,N_13215);
nor U24850 (N_24850,N_18081,N_12426);
or U24851 (N_24851,N_15657,N_10057);
and U24852 (N_24852,N_19715,N_16016);
xnor U24853 (N_24853,N_14325,N_13370);
nor U24854 (N_24854,N_12822,N_11277);
and U24855 (N_24855,N_13970,N_10394);
nor U24856 (N_24856,N_19858,N_10935);
xor U24857 (N_24857,N_19594,N_14697);
or U24858 (N_24858,N_18103,N_15266);
nor U24859 (N_24859,N_15069,N_16149);
nand U24860 (N_24860,N_14231,N_15161);
nand U24861 (N_24861,N_15201,N_15697);
nand U24862 (N_24862,N_14372,N_15350);
nor U24863 (N_24863,N_11768,N_13534);
or U24864 (N_24864,N_11177,N_18350);
or U24865 (N_24865,N_12473,N_19935);
or U24866 (N_24866,N_13767,N_16476);
nor U24867 (N_24867,N_13742,N_15476);
or U24868 (N_24868,N_11875,N_16958);
nor U24869 (N_24869,N_16180,N_12953);
nand U24870 (N_24870,N_10452,N_18369);
nor U24871 (N_24871,N_13247,N_17464);
or U24872 (N_24872,N_19782,N_19686);
and U24873 (N_24873,N_16206,N_13833);
and U24874 (N_24874,N_18483,N_17961);
xnor U24875 (N_24875,N_11435,N_19714);
nand U24876 (N_24876,N_15581,N_10134);
nand U24877 (N_24877,N_12055,N_17955);
nor U24878 (N_24878,N_19700,N_18596);
or U24879 (N_24879,N_15969,N_15496);
and U24880 (N_24880,N_14444,N_16368);
and U24881 (N_24881,N_15165,N_10552);
nand U24882 (N_24882,N_16517,N_16220);
or U24883 (N_24883,N_15343,N_11473);
xor U24884 (N_24884,N_19654,N_16185);
or U24885 (N_24885,N_19024,N_10369);
and U24886 (N_24886,N_12922,N_13968);
and U24887 (N_24887,N_10126,N_19828);
and U24888 (N_24888,N_12649,N_13376);
nor U24889 (N_24889,N_15451,N_17726);
and U24890 (N_24890,N_16061,N_13684);
or U24891 (N_24891,N_19703,N_13645);
or U24892 (N_24892,N_18876,N_10939);
nor U24893 (N_24893,N_17945,N_16767);
xor U24894 (N_24894,N_12193,N_16987);
or U24895 (N_24895,N_14481,N_16110);
nand U24896 (N_24896,N_14004,N_18462);
nor U24897 (N_24897,N_10909,N_10851);
nand U24898 (N_24898,N_17124,N_12021);
or U24899 (N_24899,N_16522,N_10531);
nand U24900 (N_24900,N_16625,N_17251);
nand U24901 (N_24901,N_11076,N_17074);
nor U24902 (N_24902,N_17801,N_18761);
nand U24903 (N_24903,N_10370,N_16978);
xnor U24904 (N_24904,N_11630,N_11606);
nor U24905 (N_24905,N_10441,N_14716);
nor U24906 (N_24906,N_12714,N_18430);
xor U24907 (N_24907,N_11027,N_10715);
and U24908 (N_24908,N_17478,N_14085);
or U24909 (N_24909,N_13639,N_17563);
and U24910 (N_24910,N_10172,N_19723);
and U24911 (N_24911,N_11921,N_12616);
nand U24912 (N_24912,N_19437,N_10884);
and U24913 (N_24913,N_18380,N_16438);
and U24914 (N_24914,N_15009,N_18838);
or U24915 (N_24915,N_14577,N_13020);
nand U24916 (N_24916,N_11577,N_10897);
nand U24917 (N_24917,N_19868,N_13374);
or U24918 (N_24918,N_17512,N_11482);
or U24919 (N_24919,N_10833,N_19194);
nor U24920 (N_24920,N_16666,N_12908);
nand U24921 (N_24921,N_14897,N_16917);
and U24922 (N_24922,N_12980,N_17105);
nand U24923 (N_24923,N_10092,N_14090);
and U24924 (N_24924,N_16424,N_19583);
or U24925 (N_24925,N_19079,N_10772);
or U24926 (N_24926,N_14781,N_17790);
and U24927 (N_24927,N_13064,N_11614);
nand U24928 (N_24928,N_18938,N_19759);
nand U24929 (N_24929,N_11505,N_16685);
nand U24930 (N_24930,N_12066,N_16319);
nor U24931 (N_24931,N_12961,N_11972);
nand U24932 (N_24932,N_10983,N_15539);
or U24933 (N_24933,N_18307,N_11565);
and U24934 (N_24934,N_14027,N_12403);
and U24935 (N_24935,N_13169,N_17081);
or U24936 (N_24936,N_14865,N_19399);
nand U24937 (N_24937,N_10340,N_15730);
nand U24938 (N_24938,N_11924,N_18670);
and U24939 (N_24939,N_12313,N_10099);
nand U24940 (N_24940,N_19541,N_10384);
nand U24941 (N_24941,N_16791,N_16408);
nor U24942 (N_24942,N_16600,N_12447);
and U24943 (N_24943,N_19124,N_12034);
nor U24944 (N_24944,N_13927,N_10978);
and U24945 (N_24945,N_13472,N_18391);
and U24946 (N_24946,N_18591,N_10005);
nand U24947 (N_24947,N_11058,N_16106);
and U24948 (N_24948,N_15145,N_18468);
nor U24949 (N_24949,N_14802,N_11490);
nand U24950 (N_24950,N_19026,N_10333);
or U24951 (N_24951,N_11931,N_10701);
nor U24952 (N_24952,N_16739,N_14341);
or U24953 (N_24953,N_11495,N_19610);
nor U24954 (N_24954,N_15500,N_15567);
nand U24955 (N_24955,N_13796,N_19062);
and U24956 (N_24956,N_11839,N_18314);
xnor U24957 (N_24957,N_13650,N_18374);
nor U24958 (N_24958,N_19734,N_17427);
and U24959 (N_24959,N_19385,N_17166);
xor U24960 (N_24960,N_10402,N_19153);
or U24961 (N_24961,N_14998,N_12086);
or U24962 (N_24962,N_11887,N_11148);
and U24963 (N_24963,N_10132,N_19387);
nor U24964 (N_24964,N_17309,N_13473);
or U24965 (N_24965,N_14189,N_17690);
or U24966 (N_24966,N_14829,N_16617);
nor U24967 (N_24967,N_16355,N_18933);
or U24968 (N_24968,N_11429,N_16300);
xor U24969 (N_24969,N_15399,N_14080);
nor U24970 (N_24970,N_17587,N_17660);
or U24971 (N_24971,N_10448,N_10341);
and U24972 (N_24972,N_19710,N_12259);
xnor U24973 (N_24973,N_11498,N_17717);
xnor U24974 (N_24974,N_12942,N_18270);
nand U24975 (N_24975,N_10929,N_19027);
and U24976 (N_24976,N_10249,N_12521);
and U24977 (N_24977,N_13038,N_19672);
nand U24978 (N_24978,N_19231,N_19481);
or U24979 (N_24979,N_10852,N_15858);
or U24980 (N_24980,N_15544,N_14217);
or U24981 (N_24981,N_19254,N_15517);
nor U24982 (N_24982,N_18845,N_10974);
and U24983 (N_24983,N_16054,N_12551);
xor U24984 (N_24984,N_13328,N_18956);
nor U24985 (N_24985,N_11078,N_12588);
nand U24986 (N_24986,N_15157,N_17420);
or U24987 (N_24987,N_18980,N_11541);
and U24988 (N_24988,N_12293,N_16970);
nand U24989 (N_24989,N_19838,N_11114);
nor U24990 (N_24990,N_12317,N_17123);
and U24991 (N_24991,N_11491,N_10229);
xor U24992 (N_24992,N_14925,N_17674);
xor U24993 (N_24993,N_11744,N_11610);
nand U24994 (N_24994,N_13475,N_12246);
nor U24995 (N_24995,N_11796,N_19151);
or U24996 (N_24996,N_12799,N_10476);
nand U24997 (N_24997,N_18457,N_12869);
nor U24998 (N_24998,N_10403,N_19038);
or U24999 (N_24999,N_18945,N_13999);
and U25000 (N_25000,N_19888,N_10208);
nand U25001 (N_25001,N_14235,N_10594);
nand U25002 (N_25002,N_16361,N_16546);
nand U25003 (N_25003,N_10850,N_12139);
and U25004 (N_25004,N_16537,N_15390);
and U25005 (N_25005,N_16312,N_11339);
nor U25006 (N_25006,N_14886,N_11794);
nand U25007 (N_25007,N_10825,N_14141);
nor U25008 (N_25008,N_18241,N_16781);
nor U25009 (N_25009,N_11241,N_19629);
and U25010 (N_25010,N_14277,N_17377);
or U25011 (N_25011,N_16835,N_14101);
nand U25012 (N_25012,N_15173,N_14825);
nor U25013 (N_25013,N_16178,N_15144);
or U25014 (N_25014,N_19475,N_10697);
and U25015 (N_25015,N_15298,N_11981);
nor U25016 (N_25016,N_19373,N_13318);
or U25017 (N_25017,N_11145,N_17756);
nor U25018 (N_25018,N_12058,N_18009);
nand U25019 (N_25019,N_14955,N_18045);
and U25020 (N_25020,N_10429,N_18682);
xnor U25021 (N_25021,N_15954,N_17974);
and U25022 (N_25022,N_14748,N_11334);
nand U25023 (N_25023,N_13493,N_17472);
nor U25024 (N_25024,N_14136,N_13401);
nor U25025 (N_25025,N_15146,N_13984);
nor U25026 (N_25026,N_13014,N_18072);
or U25027 (N_25027,N_18421,N_14567);
or U25028 (N_25028,N_18023,N_16737);
nand U25029 (N_25029,N_19394,N_13875);
xnor U25030 (N_25030,N_19862,N_12299);
and U25031 (N_25031,N_14708,N_19002);
and U25032 (N_25032,N_11343,N_11369);
and U25033 (N_25033,N_13107,N_13267);
or U25034 (N_25034,N_13991,N_10246);
xnor U25035 (N_25035,N_13891,N_19136);
nor U25036 (N_25036,N_12145,N_18074);
or U25037 (N_25037,N_16063,N_13702);
nor U25038 (N_25038,N_18144,N_16275);
or U25039 (N_25039,N_18775,N_11344);
nand U25040 (N_25040,N_15652,N_13287);
xor U25041 (N_25041,N_14881,N_11866);
and U25042 (N_25042,N_11410,N_19347);
or U25043 (N_25043,N_18653,N_11064);
or U25044 (N_25044,N_17495,N_13076);
and U25045 (N_25045,N_13240,N_15337);
nand U25046 (N_25046,N_11743,N_16844);
and U25047 (N_25047,N_14644,N_18106);
nand U25048 (N_25048,N_17454,N_16809);
nand U25049 (N_25049,N_13484,N_12314);
nand U25050 (N_25050,N_13984,N_15245);
nand U25051 (N_25051,N_18806,N_12193);
nand U25052 (N_25052,N_17713,N_14970);
nor U25053 (N_25053,N_12448,N_17076);
and U25054 (N_25054,N_10271,N_18648);
nand U25055 (N_25055,N_11560,N_17140);
nand U25056 (N_25056,N_18502,N_19145);
or U25057 (N_25057,N_17579,N_10511);
nor U25058 (N_25058,N_17705,N_19229);
nand U25059 (N_25059,N_18181,N_13246);
or U25060 (N_25060,N_14527,N_18427);
and U25061 (N_25061,N_14945,N_10689);
nand U25062 (N_25062,N_14412,N_13792);
nor U25063 (N_25063,N_12253,N_13006);
nand U25064 (N_25064,N_14911,N_11972);
nor U25065 (N_25065,N_12655,N_13826);
or U25066 (N_25066,N_13371,N_11128);
and U25067 (N_25067,N_14050,N_15692);
or U25068 (N_25068,N_15561,N_16278);
xnor U25069 (N_25069,N_16233,N_10925);
nor U25070 (N_25070,N_12994,N_14088);
or U25071 (N_25071,N_12235,N_16924);
xor U25072 (N_25072,N_10398,N_14750);
and U25073 (N_25073,N_16675,N_18132);
or U25074 (N_25074,N_11361,N_13514);
nor U25075 (N_25075,N_11637,N_15412);
xnor U25076 (N_25076,N_18298,N_12038);
or U25077 (N_25077,N_12253,N_17990);
and U25078 (N_25078,N_17306,N_17677);
and U25079 (N_25079,N_11374,N_17588);
nor U25080 (N_25080,N_14341,N_13432);
or U25081 (N_25081,N_18357,N_19252);
nand U25082 (N_25082,N_14027,N_16468);
or U25083 (N_25083,N_13457,N_19159);
or U25084 (N_25084,N_19381,N_16618);
and U25085 (N_25085,N_14950,N_15590);
nor U25086 (N_25086,N_17069,N_17411);
xor U25087 (N_25087,N_12031,N_13756);
nand U25088 (N_25088,N_17436,N_13835);
or U25089 (N_25089,N_16892,N_15046);
nand U25090 (N_25090,N_12006,N_18594);
nand U25091 (N_25091,N_13323,N_11285);
or U25092 (N_25092,N_18459,N_11537);
nand U25093 (N_25093,N_12566,N_14718);
nor U25094 (N_25094,N_16776,N_16409);
nor U25095 (N_25095,N_11491,N_11226);
or U25096 (N_25096,N_16789,N_10450);
nor U25097 (N_25097,N_11660,N_14718);
nand U25098 (N_25098,N_15584,N_19662);
nor U25099 (N_25099,N_13528,N_16432);
and U25100 (N_25100,N_13013,N_16042);
nor U25101 (N_25101,N_19821,N_11681);
nor U25102 (N_25102,N_19473,N_10302);
and U25103 (N_25103,N_17138,N_19244);
nor U25104 (N_25104,N_18553,N_11628);
or U25105 (N_25105,N_11976,N_13909);
or U25106 (N_25106,N_17043,N_14471);
and U25107 (N_25107,N_11588,N_17533);
nor U25108 (N_25108,N_18332,N_13396);
nor U25109 (N_25109,N_18902,N_10405);
nor U25110 (N_25110,N_12265,N_13336);
xnor U25111 (N_25111,N_15512,N_12927);
or U25112 (N_25112,N_16003,N_10802);
nand U25113 (N_25113,N_11356,N_11542);
nand U25114 (N_25114,N_16756,N_13026);
nand U25115 (N_25115,N_10812,N_11984);
nor U25116 (N_25116,N_19222,N_16271);
nand U25117 (N_25117,N_10916,N_13233);
or U25118 (N_25118,N_11139,N_19786);
and U25119 (N_25119,N_12385,N_18668);
and U25120 (N_25120,N_17369,N_16438);
or U25121 (N_25121,N_10635,N_12466);
or U25122 (N_25122,N_13020,N_11210);
nand U25123 (N_25123,N_18490,N_15198);
nand U25124 (N_25124,N_10775,N_13478);
or U25125 (N_25125,N_11213,N_11817);
and U25126 (N_25126,N_12454,N_13716);
nor U25127 (N_25127,N_18350,N_14482);
or U25128 (N_25128,N_15152,N_16443);
nor U25129 (N_25129,N_12163,N_17267);
nand U25130 (N_25130,N_14974,N_15988);
nor U25131 (N_25131,N_16070,N_15599);
or U25132 (N_25132,N_19526,N_17615);
nand U25133 (N_25133,N_11746,N_13847);
and U25134 (N_25134,N_16486,N_10256);
nand U25135 (N_25135,N_10119,N_13357);
xor U25136 (N_25136,N_17352,N_17703);
nor U25137 (N_25137,N_19119,N_15808);
nand U25138 (N_25138,N_10797,N_10061);
nor U25139 (N_25139,N_14568,N_14582);
or U25140 (N_25140,N_15454,N_12740);
nand U25141 (N_25141,N_11893,N_17892);
nand U25142 (N_25142,N_10362,N_13335);
xnor U25143 (N_25143,N_17735,N_11604);
nand U25144 (N_25144,N_19270,N_15379);
or U25145 (N_25145,N_15314,N_15846);
nand U25146 (N_25146,N_12717,N_18749);
and U25147 (N_25147,N_17751,N_13938);
or U25148 (N_25148,N_10398,N_15958);
or U25149 (N_25149,N_18399,N_14304);
and U25150 (N_25150,N_11356,N_17420);
or U25151 (N_25151,N_13380,N_19181);
or U25152 (N_25152,N_17431,N_16724);
or U25153 (N_25153,N_10816,N_15696);
nor U25154 (N_25154,N_18834,N_10960);
or U25155 (N_25155,N_13618,N_16580);
or U25156 (N_25156,N_14979,N_14754);
and U25157 (N_25157,N_17166,N_16660);
and U25158 (N_25158,N_11580,N_17986);
nand U25159 (N_25159,N_16252,N_12378);
and U25160 (N_25160,N_16304,N_17383);
xnor U25161 (N_25161,N_15894,N_11441);
nor U25162 (N_25162,N_12972,N_19132);
and U25163 (N_25163,N_17716,N_10417);
and U25164 (N_25164,N_15728,N_19548);
or U25165 (N_25165,N_14761,N_11542);
and U25166 (N_25166,N_10036,N_14983);
nor U25167 (N_25167,N_17543,N_15178);
nand U25168 (N_25168,N_15602,N_18514);
nor U25169 (N_25169,N_19899,N_17555);
or U25170 (N_25170,N_12026,N_19447);
nand U25171 (N_25171,N_19217,N_19228);
or U25172 (N_25172,N_11327,N_18749);
or U25173 (N_25173,N_10211,N_13501);
xnor U25174 (N_25174,N_17560,N_14402);
and U25175 (N_25175,N_17127,N_13010);
nand U25176 (N_25176,N_18570,N_14300);
and U25177 (N_25177,N_17274,N_16519);
nand U25178 (N_25178,N_16658,N_10728);
nand U25179 (N_25179,N_14156,N_10748);
and U25180 (N_25180,N_18418,N_14860);
and U25181 (N_25181,N_13461,N_11839);
or U25182 (N_25182,N_12742,N_18641);
nand U25183 (N_25183,N_12934,N_17806);
nand U25184 (N_25184,N_16182,N_10460);
and U25185 (N_25185,N_19815,N_10222);
xnor U25186 (N_25186,N_15968,N_10252);
and U25187 (N_25187,N_18963,N_17039);
or U25188 (N_25188,N_12140,N_16207);
xnor U25189 (N_25189,N_17413,N_12928);
and U25190 (N_25190,N_11171,N_11119);
and U25191 (N_25191,N_19905,N_13245);
nand U25192 (N_25192,N_12560,N_11991);
or U25193 (N_25193,N_19259,N_10455);
or U25194 (N_25194,N_15029,N_13119);
nand U25195 (N_25195,N_11031,N_12405);
and U25196 (N_25196,N_16557,N_15569);
nor U25197 (N_25197,N_10963,N_19605);
or U25198 (N_25198,N_10278,N_13869);
and U25199 (N_25199,N_18707,N_17100);
or U25200 (N_25200,N_19207,N_17250);
nand U25201 (N_25201,N_17139,N_16450);
and U25202 (N_25202,N_17540,N_10821);
nand U25203 (N_25203,N_13788,N_18043);
xor U25204 (N_25204,N_12885,N_12292);
and U25205 (N_25205,N_15551,N_14170);
xor U25206 (N_25206,N_10476,N_12951);
or U25207 (N_25207,N_17764,N_16866);
nand U25208 (N_25208,N_16662,N_15768);
nand U25209 (N_25209,N_15791,N_15241);
or U25210 (N_25210,N_12022,N_19158);
nand U25211 (N_25211,N_18571,N_12419);
nor U25212 (N_25212,N_19861,N_18734);
or U25213 (N_25213,N_13776,N_17390);
nor U25214 (N_25214,N_19515,N_18241);
xor U25215 (N_25215,N_18770,N_15162);
xnor U25216 (N_25216,N_16048,N_10226);
and U25217 (N_25217,N_17986,N_14095);
nand U25218 (N_25218,N_17316,N_12445);
or U25219 (N_25219,N_19125,N_18911);
xor U25220 (N_25220,N_15194,N_14521);
nor U25221 (N_25221,N_11377,N_11374);
xnor U25222 (N_25222,N_15040,N_11388);
nand U25223 (N_25223,N_19892,N_19194);
or U25224 (N_25224,N_18342,N_13109);
and U25225 (N_25225,N_14293,N_14132);
and U25226 (N_25226,N_11799,N_15577);
nor U25227 (N_25227,N_16993,N_19322);
or U25228 (N_25228,N_15800,N_19108);
nor U25229 (N_25229,N_14626,N_19058);
nand U25230 (N_25230,N_18653,N_10056);
and U25231 (N_25231,N_19552,N_14596);
xor U25232 (N_25232,N_12187,N_13353);
nor U25233 (N_25233,N_15813,N_12629);
nor U25234 (N_25234,N_10692,N_13438);
nor U25235 (N_25235,N_14934,N_12327);
or U25236 (N_25236,N_15870,N_10613);
nand U25237 (N_25237,N_16954,N_15037);
or U25238 (N_25238,N_18404,N_18608);
nand U25239 (N_25239,N_18162,N_15977);
and U25240 (N_25240,N_17157,N_18197);
nand U25241 (N_25241,N_14020,N_17670);
nand U25242 (N_25242,N_17917,N_13132);
xor U25243 (N_25243,N_15946,N_19130);
or U25244 (N_25244,N_18913,N_14618);
or U25245 (N_25245,N_15875,N_12936);
nand U25246 (N_25246,N_17826,N_10391);
and U25247 (N_25247,N_10656,N_12085);
or U25248 (N_25248,N_13035,N_18395);
nand U25249 (N_25249,N_18727,N_17525);
nand U25250 (N_25250,N_19366,N_18536);
or U25251 (N_25251,N_19473,N_14929);
xnor U25252 (N_25252,N_10076,N_17714);
nor U25253 (N_25253,N_10042,N_11858);
nand U25254 (N_25254,N_10475,N_17378);
xnor U25255 (N_25255,N_12634,N_11882);
and U25256 (N_25256,N_11335,N_11391);
nand U25257 (N_25257,N_11524,N_18557);
and U25258 (N_25258,N_16637,N_13943);
and U25259 (N_25259,N_15582,N_13704);
or U25260 (N_25260,N_14972,N_13803);
or U25261 (N_25261,N_12105,N_13109);
and U25262 (N_25262,N_10666,N_19218);
nand U25263 (N_25263,N_12190,N_18497);
and U25264 (N_25264,N_18182,N_10516);
and U25265 (N_25265,N_19616,N_15190);
or U25266 (N_25266,N_11315,N_14165);
nand U25267 (N_25267,N_10571,N_16503);
or U25268 (N_25268,N_11855,N_19883);
and U25269 (N_25269,N_19152,N_19499);
or U25270 (N_25270,N_10556,N_12908);
xnor U25271 (N_25271,N_19954,N_16750);
nand U25272 (N_25272,N_16264,N_10719);
or U25273 (N_25273,N_18013,N_16031);
xnor U25274 (N_25274,N_11036,N_10176);
and U25275 (N_25275,N_17939,N_17733);
nor U25276 (N_25276,N_17552,N_17459);
nor U25277 (N_25277,N_12517,N_15057);
nor U25278 (N_25278,N_12784,N_14502);
and U25279 (N_25279,N_11003,N_13727);
nand U25280 (N_25280,N_14771,N_16167);
nand U25281 (N_25281,N_15776,N_17911);
nand U25282 (N_25282,N_19092,N_12153);
or U25283 (N_25283,N_16180,N_15101);
or U25284 (N_25284,N_14051,N_11861);
or U25285 (N_25285,N_12899,N_17369);
and U25286 (N_25286,N_12982,N_16064);
nand U25287 (N_25287,N_19741,N_17778);
nand U25288 (N_25288,N_18548,N_16308);
and U25289 (N_25289,N_19614,N_12644);
and U25290 (N_25290,N_12537,N_15412);
nand U25291 (N_25291,N_16551,N_16577);
nor U25292 (N_25292,N_16780,N_10322);
and U25293 (N_25293,N_18039,N_16649);
or U25294 (N_25294,N_15083,N_18369);
or U25295 (N_25295,N_12314,N_14955);
and U25296 (N_25296,N_10747,N_16215);
xnor U25297 (N_25297,N_16299,N_17514);
and U25298 (N_25298,N_19699,N_16233);
and U25299 (N_25299,N_10905,N_11693);
and U25300 (N_25300,N_11917,N_15112);
and U25301 (N_25301,N_13518,N_18579);
nand U25302 (N_25302,N_12167,N_19812);
and U25303 (N_25303,N_12088,N_10228);
nand U25304 (N_25304,N_13476,N_18615);
and U25305 (N_25305,N_12920,N_19264);
or U25306 (N_25306,N_18807,N_15089);
nand U25307 (N_25307,N_11161,N_13672);
nor U25308 (N_25308,N_10821,N_14570);
and U25309 (N_25309,N_10757,N_13010);
nor U25310 (N_25310,N_15847,N_15878);
nand U25311 (N_25311,N_16786,N_19070);
and U25312 (N_25312,N_11694,N_11224);
and U25313 (N_25313,N_17280,N_14742);
or U25314 (N_25314,N_18807,N_15693);
or U25315 (N_25315,N_19547,N_19564);
or U25316 (N_25316,N_19965,N_18647);
nand U25317 (N_25317,N_10830,N_14176);
or U25318 (N_25318,N_14919,N_15792);
nand U25319 (N_25319,N_15874,N_10055);
and U25320 (N_25320,N_17390,N_17038);
and U25321 (N_25321,N_17918,N_15097);
and U25322 (N_25322,N_11173,N_15337);
or U25323 (N_25323,N_11168,N_14350);
nor U25324 (N_25324,N_18473,N_16504);
or U25325 (N_25325,N_13387,N_10764);
nand U25326 (N_25326,N_10360,N_16411);
or U25327 (N_25327,N_15746,N_18041);
or U25328 (N_25328,N_11798,N_13513);
nor U25329 (N_25329,N_16732,N_16193);
and U25330 (N_25330,N_11224,N_14064);
and U25331 (N_25331,N_18761,N_17930);
and U25332 (N_25332,N_13484,N_19929);
and U25333 (N_25333,N_15317,N_15143);
or U25334 (N_25334,N_18759,N_14401);
nor U25335 (N_25335,N_14234,N_14973);
nor U25336 (N_25336,N_19338,N_15029);
nor U25337 (N_25337,N_12242,N_19958);
and U25338 (N_25338,N_11854,N_18192);
or U25339 (N_25339,N_11418,N_18738);
or U25340 (N_25340,N_15447,N_18614);
nand U25341 (N_25341,N_13100,N_10706);
nor U25342 (N_25342,N_13469,N_17752);
or U25343 (N_25343,N_14544,N_15689);
nand U25344 (N_25344,N_15270,N_17932);
or U25345 (N_25345,N_17294,N_18243);
nor U25346 (N_25346,N_10696,N_13204);
nor U25347 (N_25347,N_17552,N_18884);
or U25348 (N_25348,N_10149,N_11152);
nor U25349 (N_25349,N_14329,N_10884);
nand U25350 (N_25350,N_17995,N_17162);
nand U25351 (N_25351,N_17470,N_19075);
nand U25352 (N_25352,N_10341,N_15989);
and U25353 (N_25353,N_14634,N_14414);
xnor U25354 (N_25354,N_11110,N_19242);
or U25355 (N_25355,N_10983,N_16931);
nand U25356 (N_25356,N_13001,N_10413);
nand U25357 (N_25357,N_16996,N_14766);
or U25358 (N_25358,N_16436,N_18512);
xnor U25359 (N_25359,N_14311,N_14428);
and U25360 (N_25360,N_14410,N_17241);
nand U25361 (N_25361,N_17713,N_18933);
nand U25362 (N_25362,N_11525,N_17253);
nor U25363 (N_25363,N_10067,N_14951);
nor U25364 (N_25364,N_13786,N_15648);
and U25365 (N_25365,N_19384,N_14593);
or U25366 (N_25366,N_11735,N_16741);
nand U25367 (N_25367,N_17678,N_11870);
xnor U25368 (N_25368,N_10186,N_13284);
xnor U25369 (N_25369,N_16784,N_12799);
xnor U25370 (N_25370,N_10166,N_19964);
xnor U25371 (N_25371,N_15995,N_19673);
nand U25372 (N_25372,N_10071,N_12750);
xnor U25373 (N_25373,N_10580,N_11078);
and U25374 (N_25374,N_15605,N_12640);
xor U25375 (N_25375,N_13921,N_15724);
or U25376 (N_25376,N_12032,N_17268);
and U25377 (N_25377,N_10623,N_17839);
or U25378 (N_25378,N_15955,N_11252);
and U25379 (N_25379,N_10339,N_11270);
nand U25380 (N_25380,N_14673,N_14245);
nand U25381 (N_25381,N_15027,N_13027);
nand U25382 (N_25382,N_11392,N_12381);
and U25383 (N_25383,N_14726,N_16290);
and U25384 (N_25384,N_14612,N_15720);
nor U25385 (N_25385,N_19942,N_13304);
and U25386 (N_25386,N_15270,N_15688);
nand U25387 (N_25387,N_15532,N_14318);
nand U25388 (N_25388,N_11472,N_17862);
nor U25389 (N_25389,N_13911,N_16289);
xor U25390 (N_25390,N_18660,N_19444);
nand U25391 (N_25391,N_10596,N_10978);
nor U25392 (N_25392,N_17536,N_19136);
xnor U25393 (N_25393,N_11289,N_15097);
and U25394 (N_25394,N_15816,N_18369);
xor U25395 (N_25395,N_18985,N_14057);
nand U25396 (N_25396,N_16926,N_13615);
xor U25397 (N_25397,N_14787,N_16494);
nand U25398 (N_25398,N_14223,N_18478);
nand U25399 (N_25399,N_18859,N_16926);
xnor U25400 (N_25400,N_16502,N_11142);
nor U25401 (N_25401,N_11392,N_19816);
or U25402 (N_25402,N_15826,N_11738);
or U25403 (N_25403,N_17231,N_10352);
and U25404 (N_25404,N_19979,N_12296);
or U25405 (N_25405,N_17278,N_16022);
nand U25406 (N_25406,N_13104,N_16566);
and U25407 (N_25407,N_19134,N_16631);
nand U25408 (N_25408,N_11549,N_10873);
nor U25409 (N_25409,N_16879,N_12421);
or U25410 (N_25410,N_18128,N_10133);
and U25411 (N_25411,N_10825,N_18590);
or U25412 (N_25412,N_13385,N_19995);
and U25413 (N_25413,N_14529,N_10527);
nand U25414 (N_25414,N_12845,N_16134);
or U25415 (N_25415,N_14222,N_10363);
nand U25416 (N_25416,N_14336,N_12190);
or U25417 (N_25417,N_19721,N_15046);
and U25418 (N_25418,N_19335,N_14706);
nand U25419 (N_25419,N_16100,N_18463);
xnor U25420 (N_25420,N_16367,N_11878);
xnor U25421 (N_25421,N_13831,N_14189);
xnor U25422 (N_25422,N_13825,N_16639);
and U25423 (N_25423,N_16252,N_18008);
nor U25424 (N_25424,N_19283,N_18777);
and U25425 (N_25425,N_10312,N_14376);
nor U25426 (N_25426,N_18408,N_18490);
nand U25427 (N_25427,N_15035,N_13175);
xor U25428 (N_25428,N_17068,N_14975);
or U25429 (N_25429,N_18038,N_16653);
nand U25430 (N_25430,N_14332,N_14288);
xnor U25431 (N_25431,N_11462,N_11559);
nor U25432 (N_25432,N_16725,N_11019);
nand U25433 (N_25433,N_10347,N_17638);
and U25434 (N_25434,N_11886,N_16706);
nand U25435 (N_25435,N_19642,N_16390);
and U25436 (N_25436,N_11327,N_17297);
and U25437 (N_25437,N_15799,N_18456);
or U25438 (N_25438,N_19673,N_15332);
nor U25439 (N_25439,N_10298,N_19638);
and U25440 (N_25440,N_17795,N_10681);
nand U25441 (N_25441,N_18526,N_10608);
nor U25442 (N_25442,N_17119,N_10670);
nor U25443 (N_25443,N_12950,N_13730);
and U25444 (N_25444,N_14446,N_15671);
or U25445 (N_25445,N_13423,N_14703);
nor U25446 (N_25446,N_17129,N_16530);
or U25447 (N_25447,N_17890,N_16627);
nand U25448 (N_25448,N_11279,N_18952);
nor U25449 (N_25449,N_12861,N_19058);
nor U25450 (N_25450,N_18130,N_16960);
nand U25451 (N_25451,N_17626,N_11623);
xnor U25452 (N_25452,N_15100,N_15819);
xor U25453 (N_25453,N_13078,N_14533);
or U25454 (N_25454,N_18861,N_10866);
or U25455 (N_25455,N_17657,N_15499);
nor U25456 (N_25456,N_18138,N_12335);
nand U25457 (N_25457,N_10870,N_16131);
nand U25458 (N_25458,N_13254,N_13017);
nor U25459 (N_25459,N_16608,N_13934);
and U25460 (N_25460,N_12628,N_17407);
and U25461 (N_25461,N_16203,N_14315);
and U25462 (N_25462,N_12573,N_14799);
nor U25463 (N_25463,N_11336,N_18301);
nor U25464 (N_25464,N_14081,N_11643);
xor U25465 (N_25465,N_13833,N_19429);
and U25466 (N_25466,N_18103,N_14349);
or U25467 (N_25467,N_10638,N_15322);
and U25468 (N_25468,N_11908,N_17303);
xor U25469 (N_25469,N_17385,N_18716);
and U25470 (N_25470,N_19610,N_17425);
nor U25471 (N_25471,N_18921,N_19775);
and U25472 (N_25472,N_15884,N_10997);
nor U25473 (N_25473,N_18465,N_13271);
or U25474 (N_25474,N_12119,N_15628);
or U25475 (N_25475,N_10547,N_17367);
nor U25476 (N_25476,N_17886,N_15526);
and U25477 (N_25477,N_14724,N_15437);
xnor U25478 (N_25478,N_11864,N_16633);
and U25479 (N_25479,N_13116,N_10391);
xor U25480 (N_25480,N_17130,N_13537);
nand U25481 (N_25481,N_18406,N_19013);
nor U25482 (N_25482,N_13528,N_15821);
or U25483 (N_25483,N_11296,N_15891);
or U25484 (N_25484,N_11887,N_10104);
nand U25485 (N_25485,N_10501,N_17286);
xor U25486 (N_25486,N_12368,N_10047);
or U25487 (N_25487,N_17815,N_19509);
and U25488 (N_25488,N_11294,N_10051);
or U25489 (N_25489,N_17783,N_12575);
or U25490 (N_25490,N_12101,N_19088);
or U25491 (N_25491,N_11440,N_19983);
or U25492 (N_25492,N_11510,N_15695);
nor U25493 (N_25493,N_17165,N_13025);
nor U25494 (N_25494,N_12161,N_18512);
and U25495 (N_25495,N_17993,N_10515);
nand U25496 (N_25496,N_11727,N_15367);
or U25497 (N_25497,N_16330,N_18836);
or U25498 (N_25498,N_14072,N_11839);
nor U25499 (N_25499,N_10995,N_18363);
nand U25500 (N_25500,N_19059,N_13481);
xor U25501 (N_25501,N_12020,N_17261);
and U25502 (N_25502,N_10927,N_18356);
or U25503 (N_25503,N_16176,N_19615);
xor U25504 (N_25504,N_19878,N_12884);
or U25505 (N_25505,N_13176,N_16174);
nand U25506 (N_25506,N_14012,N_16978);
nor U25507 (N_25507,N_13826,N_19389);
and U25508 (N_25508,N_15133,N_19769);
or U25509 (N_25509,N_14370,N_13673);
nor U25510 (N_25510,N_19592,N_14653);
xnor U25511 (N_25511,N_10042,N_15368);
nand U25512 (N_25512,N_19682,N_13293);
nand U25513 (N_25513,N_16972,N_11656);
xnor U25514 (N_25514,N_13211,N_18841);
or U25515 (N_25515,N_18133,N_13310);
or U25516 (N_25516,N_10810,N_12480);
and U25517 (N_25517,N_16863,N_18046);
or U25518 (N_25518,N_13407,N_16204);
or U25519 (N_25519,N_15820,N_12620);
and U25520 (N_25520,N_19396,N_16261);
xnor U25521 (N_25521,N_11763,N_12552);
and U25522 (N_25522,N_14692,N_19250);
nand U25523 (N_25523,N_19307,N_16117);
or U25524 (N_25524,N_11746,N_19995);
xnor U25525 (N_25525,N_17363,N_12345);
xnor U25526 (N_25526,N_18152,N_10708);
nand U25527 (N_25527,N_17555,N_11077);
or U25528 (N_25528,N_12557,N_12859);
nand U25529 (N_25529,N_15649,N_18744);
nor U25530 (N_25530,N_17776,N_12262);
nand U25531 (N_25531,N_13066,N_13967);
nand U25532 (N_25532,N_14840,N_18776);
nand U25533 (N_25533,N_14804,N_17458);
or U25534 (N_25534,N_10138,N_11756);
and U25535 (N_25535,N_12298,N_10893);
nand U25536 (N_25536,N_11072,N_12847);
xnor U25537 (N_25537,N_15811,N_11794);
nand U25538 (N_25538,N_12548,N_15113);
and U25539 (N_25539,N_16002,N_15007);
nor U25540 (N_25540,N_18344,N_15120);
and U25541 (N_25541,N_19303,N_16912);
and U25542 (N_25542,N_13218,N_11722);
or U25543 (N_25543,N_19922,N_19119);
nand U25544 (N_25544,N_10639,N_10997);
or U25545 (N_25545,N_16801,N_11133);
nor U25546 (N_25546,N_14188,N_12840);
and U25547 (N_25547,N_12146,N_13602);
xnor U25548 (N_25548,N_12903,N_15197);
nor U25549 (N_25549,N_14176,N_16253);
and U25550 (N_25550,N_17266,N_12729);
nor U25551 (N_25551,N_11474,N_15547);
nor U25552 (N_25552,N_17226,N_19873);
nor U25553 (N_25553,N_19106,N_14751);
or U25554 (N_25554,N_15704,N_19189);
nand U25555 (N_25555,N_11748,N_14928);
or U25556 (N_25556,N_10484,N_10405);
nand U25557 (N_25557,N_17011,N_17083);
and U25558 (N_25558,N_19887,N_11402);
nand U25559 (N_25559,N_11736,N_13720);
nor U25560 (N_25560,N_15477,N_14469);
or U25561 (N_25561,N_16612,N_15295);
or U25562 (N_25562,N_13583,N_17716);
and U25563 (N_25563,N_12482,N_16457);
nand U25564 (N_25564,N_13613,N_11937);
xor U25565 (N_25565,N_13396,N_18101);
and U25566 (N_25566,N_17894,N_17278);
or U25567 (N_25567,N_18600,N_17012);
nor U25568 (N_25568,N_11870,N_14936);
nor U25569 (N_25569,N_10348,N_19374);
xnor U25570 (N_25570,N_17367,N_18045);
nor U25571 (N_25571,N_13020,N_14379);
nor U25572 (N_25572,N_14313,N_12219);
and U25573 (N_25573,N_15982,N_11261);
nand U25574 (N_25574,N_14391,N_17859);
nor U25575 (N_25575,N_13291,N_12530);
and U25576 (N_25576,N_12391,N_16801);
or U25577 (N_25577,N_13119,N_18127);
and U25578 (N_25578,N_18605,N_14599);
and U25579 (N_25579,N_17965,N_11462);
nor U25580 (N_25580,N_15431,N_11736);
or U25581 (N_25581,N_17106,N_14814);
and U25582 (N_25582,N_11299,N_16022);
and U25583 (N_25583,N_15384,N_11487);
and U25584 (N_25584,N_17209,N_13432);
or U25585 (N_25585,N_10017,N_17264);
nor U25586 (N_25586,N_13381,N_18414);
or U25587 (N_25587,N_12404,N_12208);
xnor U25588 (N_25588,N_14644,N_13584);
or U25589 (N_25589,N_17634,N_13279);
or U25590 (N_25590,N_17757,N_19033);
or U25591 (N_25591,N_10458,N_17665);
nor U25592 (N_25592,N_10043,N_19912);
or U25593 (N_25593,N_13264,N_10810);
nor U25594 (N_25594,N_16360,N_12654);
nand U25595 (N_25595,N_17383,N_14069);
nor U25596 (N_25596,N_13294,N_19142);
nand U25597 (N_25597,N_19429,N_15269);
and U25598 (N_25598,N_16590,N_19777);
or U25599 (N_25599,N_12767,N_16414);
or U25600 (N_25600,N_10334,N_13962);
nor U25601 (N_25601,N_10884,N_15315);
or U25602 (N_25602,N_15149,N_17484);
and U25603 (N_25603,N_15724,N_13827);
nand U25604 (N_25604,N_11937,N_15257);
xor U25605 (N_25605,N_17823,N_19134);
or U25606 (N_25606,N_17320,N_12090);
and U25607 (N_25607,N_17926,N_17611);
nand U25608 (N_25608,N_12024,N_14448);
nand U25609 (N_25609,N_11881,N_11254);
nor U25610 (N_25610,N_12203,N_19604);
nor U25611 (N_25611,N_15119,N_17690);
or U25612 (N_25612,N_16736,N_11343);
nor U25613 (N_25613,N_11734,N_19672);
or U25614 (N_25614,N_13949,N_15659);
nand U25615 (N_25615,N_17301,N_12518);
nand U25616 (N_25616,N_17076,N_12803);
and U25617 (N_25617,N_12596,N_17153);
nand U25618 (N_25618,N_17677,N_11444);
nand U25619 (N_25619,N_10152,N_12761);
and U25620 (N_25620,N_10460,N_15343);
or U25621 (N_25621,N_14766,N_15590);
nand U25622 (N_25622,N_17627,N_17543);
nand U25623 (N_25623,N_16757,N_15381);
nand U25624 (N_25624,N_13688,N_17372);
xnor U25625 (N_25625,N_12632,N_10527);
nor U25626 (N_25626,N_18220,N_17877);
nor U25627 (N_25627,N_14842,N_10762);
nand U25628 (N_25628,N_13034,N_13677);
or U25629 (N_25629,N_17576,N_12274);
or U25630 (N_25630,N_11455,N_16285);
nor U25631 (N_25631,N_16276,N_18498);
and U25632 (N_25632,N_14490,N_10073);
or U25633 (N_25633,N_19216,N_10284);
and U25634 (N_25634,N_10614,N_14342);
or U25635 (N_25635,N_11225,N_14665);
nor U25636 (N_25636,N_17499,N_17384);
nor U25637 (N_25637,N_16559,N_17036);
nor U25638 (N_25638,N_11072,N_11289);
or U25639 (N_25639,N_18037,N_15147);
nor U25640 (N_25640,N_12184,N_15056);
and U25641 (N_25641,N_18618,N_11291);
nor U25642 (N_25642,N_13014,N_16798);
or U25643 (N_25643,N_14644,N_15052);
nand U25644 (N_25644,N_17238,N_19233);
nor U25645 (N_25645,N_19498,N_13109);
xnor U25646 (N_25646,N_15475,N_14064);
xnor U25647 (N_25647,N_11695,N_17507);
or U25648 (N_25648,N_19793,N_18152);
or U25649 (N_25649,N_16740,N_10262);
nand U25650 (N_25650,N_12552,N_18864);
or U25651 (N_25651,N_11379,N_17213);
nand U25652 (N_25652,N_17549,N_19966);
nand U25653 (N_25653,N_10714,N_19160);
nand U25654 (N_25654,N_10912,N_16160);
nor U25655 (N_25655,N_16366,N_13859);
nor U25656 (N_25656,N_15402,N_14635);
or U25657 (N_25657,N_12794,N_18841);
and U25658 (N_25658,N_13722,N_12042);
nor U25659 (N_25659,N_11127,N_19280);
xor U25660 (N_25660,N_16388,N_18518);
nor U25661 (N_25661,N_15361,N_15714);
nand U25662 (N_25662,N_13811,N_16620);
and U25663 (N_25663,N_13941,N_17872);
xnor U25664 (N_25664,N_16626,N_15712);
xor U25665 (N_25665,N_13504,N_10306);
and U25666 (N_25666,N_10680,N_15153);
nand U25667 (N_25667,N_10320,N_15285);
nand U25668 (N_25668,N_14008,N_16575);
xnor U25669 (N_25669,N_17032,N_10246);
xnor U25670 (N_25670,N_14614,N_11520);
nand U25671 (N_25671,N_18815,N_17809);
nor U25672 (N_25672,N_16995,N_14250);
or U25673 (N_25673,N_16773,N_17153);
and U25674 (N_25674,N_19889,N_18457);
nor U25675 (N_25675,N_19086,N_19560);
and U25676 (N_25676,N_12831,N_19600);
and U25677 (N_25677,N_12231,N_17940);
and U25678 (N_25678,N_17788,N_17866);
xnor U25679 (N_25679,N_15603,N_11677);
and U25680 (N_25680,N_17564,N_19425);
nand U25681 (N_25681,N_19930,N_10711);
nand U25682 (N_25682,N_13576,N_18033);
or U25683 (N_25683,N_17812,N_17839);
and U25684 (N_25684,N_11781,N_19744);
nand U25685 (N_25685,N_16680,N_15062);
and U25686 (N_25686,N_13676,N_18730);
and U25687 (N_25687,N_13709,N_12171);
or U25688 (N_25688,N_15028,N_12337);
nand U25689 (N_25689,N_14794,N_15517);
nand U25690 (N_25690,N_18388,N_18656);
and U25691 (N_25691,N_17449,N_13420);
nor U25692 (N_25692,N_12776,N_11952);
and U25693 (N_25693,N_15411,N_12249);
nor U25694 (N_25694,N_16508,N_15509);
or U25695 (N_25695,N_15772,N_11221);
nor U25696 (N_25696,N_10823,N_10435);
xor U25697 (N_25697,N_15839,N_17395);
and U25698 (N_25698,N_17443,N_19991);
and U25699 (N_25699,N_11852,N_11441);
nand U25700 (N_25700,N_19585,N_13220);
or U25701 (N_25701,N_16504,N_19430);
xor U25702 (N_25702,N_13947,N_13557);
and U25703 (N_25703,N_15120,N_10751);
or U25704 (N_25704,N_16061,N_19485);
and U25705 (N_25705,N_12523,N_10751);
nor U25706 (N_25706,N_10721,N_11590);
or U25707 (N_25707,N_10448,N_18204);
nor U25708 (N_25708,N_14996,N_10966);
and U25709 (N_25709,N_19546,N_17489);
nand U25710 (N_25710,N_11002,N_11483);
or U25711 (N_25711,N_11730,N_14220);
or U25712 (N_25712,N_17471,N_15294);
and U25713 (N_25713,N_10622,N_19596);
xnor U25714 (N_25714,N_13055,N_12873);
and U25715 (N_25715,N_17135,N_17401);
nand U25716 (N_25716,N_18167,N_19152);
and U25717 (N_25717,N_12785,N_12533);
nand U25718 (N_25718,N_15087,N_17549);
or U25719 (N_25719,N_15097,N_15433);
or U25720 (N_25720,N_13244,N_15356);
or U25721 (N_25721,N_19458,N_18624);
and U25722 (N_25722,N_15782,N_17331);
or U25723 (N_25723,N_12930,N_14382);
or U25724 (N_25724,N_12265,N_10071);
or U25725 (N_25725,N_11274,N_15632);
and U25726 (N_25726,N_18853,N_17746);
nor U25727 (N_25727,N_12213,N_13610);
and U25728 (N_25728,N_13076,N_10670);
nand U25729 (N_25729,N_18889,N_15081);
xor U25730 (N_25730,N_13417,N_18076);
or U25731 (N_25731,N_14140,N_13832);
and U25732 (N_25732,N_18164,N_19558);
nand U25733 (N_25733,N_12031,N_16509);
nand U25734 (N_25734,N_14508,N_18573);
nand U25735 (N_25735,N_13384,N_18672);
nand U25736 (N_25736,N_11002,N_12816);
nand U25737 (N_25737,N_11384,N_10587);
and U25738 (N_25738,N_19827,N_14363);
nor U25739 (N_25739,N_12265,N_12967);
and U25740 (N_25740,N_16929,N_19591);
nor U25741 (N_25741,N_12335,N_16505);
nand U25742 (N_25742,N_14059,N_10360);
or U25743 (N_25743,N_17223,N_13198);
nor U25744 (N_25744,N_10249,N_14438);
and U25745 (N_25745,N_14784,N_10463);
or U25746 (N_25746,N_13811,N_15703);
nor U25747 (N_25747,N_17912,N_10085);
and U25748 (N_25748,N_13322,N_17763);
nand U25749 (N_25749,N_14252,N_12546);
nand U25750 (N_25750,N_18762,N_11748);
nor U25751 (N_25751,N_10766,N_18637);
xor U25752 (N_25752,N_10119,N_15253);
nor U25753 (N_25753,N_13385,N_17011);
nor U25754 (N_25754,N_12916,N_15990);
nor U25755 (N_25755,N_19051,N_15753);
nor U25756 (N_25756,N_13442,N_17274);
nand U25757 (N_25757,N_19739,N_19879);
and U25758 (N_25758,N_11324,N_16136);
nor U25759 (N_25759,N_14786,N_18229);
and U25760 (N_25760,N_18466,N_13910);
or U25761 (N_25761,N_10864,N_12668);
or U25762 (N_25762,N_14831,N_18547);
nor U25763 (N_25763,N_14794,N_15450);
and U25764 (N_25764,N_12714,N_16479);
nand U25765 (N_25765,N_17154,N_17863);
xnor U25766 (N_25766,N_14758,N_13729);
nand U25767 (N_25767,N_11215,N_10993);
and U25768 (N_25768,N_14675,N_17832);
nand U25769 (N_25769,N_12736,N_13404);
nand U25770 (N_25770,N_13805,N_11995);
or U25771 (N_25771,N_14420,N_13856);
xnor U25772 (N_25772,N_14653,N_14946);
nor U25773 (N_25773,N_10344,N_11845);
or U25774 (N_25774,N_16666,N_13363);
or U25775 (N_25775,N_16038,N_19251);
or U25776 (N_25776,N_13309,N_11583);
and U25777 (N_25777,N_16644,N_19494);
xor U25778 (N_25778,N_17016,N_11295);
and U25779 (N_25779,N_11467,N_16419);
nand U25780 (N_25780,N_17858,N_10139);
nand U25781 (N_25781,N_11184,N_14237);
and U25782 (N_25782,N_10179,N_14545);
and U25783 (N_25783,N_17960,N_13193);
or U25784 (N_25784,N_10089,N_13399);
or U25785 (N_25785,N_11310,N_14650);
and U25786 (N_25786,N_19284,N_18894);
nand U25787 (N_25787,N_18537,N_11748);
nor U25788 (N_25788,N_17321,N_11011);
or U25789 (N_25789,N_18730,N_14704);
and U25790 (N_25790,N_16947,N_10368);
nand U25791 (N_25791,N_11599,N_15117);
nor U25792 (N_25792,N_16799,N_10815);
and U25793 (N_25793,N_14804,N_16194);
nor U25794 (N_25794,N_14125,N_12819);
nand U25795 (N_25795,N_17108,N_13386);
nor U25796 (N_25796,N_14646,N_17320);
nand U25797 (N_25797,N_18329,N_19377);
or U25798 (N_25798,N_15918,N_10925);
and U25799 (N_25799,N_16711,N_19361);
nor U25800 (N_25800,N_18884,N_16249);
or U25801 (N_25801,N_16837,N_13760);
or U25802 (N_25802,N_10828,N_15746);
or U25803 (N_25803,N_13486,N_18069);
and U25804 (N_25804,N_15845,N_15556);
xor U25805 (N_25805,N_10640,N_18189);
and U25806 (N_25806,N_13924,N_11980);
nand U25807 (N_25807,N_18553,N_18862);
nor U25808 (N_25808,N_11379,N_19519);
and U25809 (N_25809,N_19001,N_12259);
nor U25810 (N_25810,N_19714,N_11327);
nand U25811 (N_25811,N_13031,N_18972);
nor U25812 (N_25812,N_19094,N_11785);
nand U25813 (N_25813,N_15203,N_10089);
or U25814 (N_25814,N_16287,N_11579);
nand U25815 (N_25815,N_15095,N_13487);
or U25816 (N_25816,N_13030,N_10721);
or U25817 (N_25817,N_15930,N_19095);
and U25818 (N_25818,N_14968,N_17243);
xnor U25819 (N_25819,N_13325,N_19204);
nor U25820 (N_25820,N_12644,N_15755);
nor U25821 (N_25821,N_11074,N_13917);
and U25822 (N_25822,N_14951,N_17169);
nand U25823 (N_25823,N_12104,N_16249);
and U25824 (N_25824,N_13909,N_11024);
or U25825 (N_25825,N_11785,N_10543);
nor U25826 (N_25826,N_18896,N_17677);
or U25827 (N_25827,N_19949,N_12375);
and U25828 (N_25828,N_12798,N_16364);
nand U25829 (N_25829,N_12377,N_14777);
or U25830 (N_25830,N_18586,N_11535);
nor U25831 (N_25831,N_19413,N_14031);
nand U25832 (N_25832,N_15789,N_12986);
and U25833 (N_25833,N_15690,N_17281);
nor U25834 (N_25834,N_12596,N_18072);
nand U25835 (N_25835,N_12408,N_11822);
nand U25836 (N_25836,N_14574,N_13587);
nor U25837 (N_25837,N_17158,N_13944);
or U25838 (N_25838,N_15943,N_12067);
and U25839 (N_25839,N_19731,N_14329);
or U25840 (N_25840,N_19251,N_15532);
and U25841 (N_25841,N_13825,N_10789);
and U25842 (N_25842,N_14487,N_15509);
nor U25843 (N_25843,N_15269,N_11323);
nand U25844 (N_25844,N_14382,N_18861);
or U25845 (N_25845,N_18307,N_13174);
or U25846 (N_25846,N_13253,N_13836);
nand U25847 (N_25847,N_18725,N_15752);
xor U25848 (N_25848,N_17183,N_18485);
and U25849 (N_25849,N_19187,N_13540);
nor U25850 (N_25850,N_12973,N_17809);
nand U25851 (N_25851,N_10154,N_13159);
nand U25852 (N_25852,N_10956,N_13559);
or U25853 (N_25853,N_10849,N_16721);
nand U25854 (N_25854,N_17886,N_13513);
nor U25855 (N_25855,N_13703,N_16353);
xnor U25856 (N_25856,N_18144,N_14400);
and U25857 (N_25857,N_18391,N_18905);
nand U25858 (N_25858,N_16033,N_10957);
and U25859 (N_25859,N_12702,N_12290);
or U25860 (N_25860,N_16716,N_10635);
nand U25861 (N_25861,N_13228,N_19751);
nand U25862 (N_25862,N_16352,N_15066);
nand U25863 (N_25863,N_19267,N_19724);
nor U25864 (N_25864,N_13211,N_16387);
and U25865 (N_25865,N_11279,N_12366);
nand U25866 (N_25866,N_13046,N_15707);
nor U25867 (N_25867,N_10009,N_16772);
nor U25868 (N_25868,N_18336,N_10619);
nor U25869 (N_25869,N_17597,N_10806);
nor U25870 (N_25870,N_12979,N_11211);
or U25871 (N_25871,N_15617,N_16835);
and U25872 (N_25872,N_15023,N_12183);
and U25873 (N_25873,N_15089,N_15564);
nand U25874 (N_25874,N_16273,N_14505);
and U25875 (N_25875,N_18250,N_10723);
xor U25876 (N_25876,N_13227,N_18794);
nor U25877 (N_25877,N_11772,N_10004);
xnor U25878 (N_25878,N_15381,N_11601);
nor U25879 (N_25879,N_18975,N_16280);
and U25880 (N_25880,N_12737,N_15947);
xor U25881 (N_25881,N_10522,N_10825);
or U25882 (N_25882,N_12766,N_17464);
xnor U25883 (N_25883,N_13230,N_12984);
xnor U25884 (N_25884,N_13911,N_19846);
nor U25885 (N_25885,N_19586,N_14319);
nand U25886 (N_25886,N_12730,N_14328);
nand U25887 (N_25887,N_18725,N_12844);
nor U25888 (N_25888,N_15270,N_14755);
nand U25889 (N_25889,N_17555,N_14746);
nand U25890 (N_25890,N_17371,N_10501);
and U25891 (N_25891,N_11082,N_12637);
nor U25892 (N_25892,N_17708,N_16853);
or U25893 (N_25893,N_16977,N_15651);
or U25894 (N_25894,N_16168,N_18671);
or U25895 (N_25895,N_13487,N_19192);
nand U25896 (N_25896,N_14001,N_11593);
or U25897 (N_25897,N_18450,N_11113);
xnor U25898 (N_25898,N_10316,N_12015);
nor U25899 (N_25899,N_12906,N_18831);
and U25900 (N_25900,N_14616,N_11620);
and U25901 (N_25901,N_15667,N_11253);
nand U25902 (N_25902,N_11605,N_14026);
nand U25903 (N_25903,N_14661,N_10819);
or U25904 (N_25904,N_15979,N_18196);
and U25905 (N_25905,N_17354,N_10570);
nand U25906 (N_25906,N_13705,N_14305);
nand U25907 (N_25907,N_16362,N_14649);
nand U25908 (N_25908,N_14044,N_13136);
nor U25909 (N_25909,N_19723,N_18664);
or U25910 (N_25910,N_11304,N_18797);
nand U25911 (N_25911,N_10975,N_14375);
nand U25912 (N_25912,N_13395,N_19434);
nand U25913 (N_25913,N_11577,N_14319);
nor U25914 (N_25914,N_11380,N_14077);
or U25915 (N_25915,N_12919,N_13050);
nand U25916 (N_25916,N_14746,N_13426);
or U25917 (N_25917,N_18220,N_16424);
nor U25918 (N_25918,N_10816,N_14901);
nand U25919 (N_25919,N_18103,N_18070);
or U25920 (N_25920,N_19011,N_12176);
nand U25921 (N_25921,N_15533,N_15870);
xor U25922 (N_25922,N_19804,N_16611);
nor U25923 (N_25923,N_13410,N_10214);
xnor U25924 (N_25924,N_13809,N_19810);
and U25925 (N_25925,N_11291,N_15482);
nor U25926 (N_25926,N_15350,N_19960);
and U25927 (N_25927,N_19877,N_11863);
nor U25928 (N_25928,N_18254,N_13735);
and U25929 (N_25929,N_10845,N_10720);
and U25930 (N_25930,N_12444,N_18138);
or U25931 (N_25931,N_16692,N_16880);
and U25932 (N_25932,N_12972,N_18299);
nor U25933 (N_25933,N_12265,N_16390);
and U25934 (N_25934,N_17688,N_15022);
nand U25935 (N_25935,N_19934,N_18758);
nor U25936 (N_25936,N_16603,N_18160);
xor U25937 (N_25937,N_15536,N_15366);
or U25938 (N_25938,N_16436,N_16773);
nor U25939 (N_25939,N_10667,N_10258);
and U25940 (N_25940,N_16250,N_11451);
nand U25941 (N_25941,N_12383,N_10119);
xnor U25942 (N_25942,N_14521,N_16711);
or U25943 (N_25943,N_11326,N_15063);
and U25944 (N_25944,N_14849,N_10005);
nand U25945 (N_25945,N_17985,N_11686);
and U25946 (N_25946,N_16503,N_12275);
nand U25947 (N_25947,N_11983,N_12981);
xor U25948 (N_25948,N_14434,N_12159);
or U25949 (N_25949,N_12746,N_17448);
and U25950 (N_25950,N_14172,N_11800);
nand U25951 (N_25951,N_16675,N_14691);
nand U25952 (N_25952,N_13249,N_19779);
and U25953 (N_25953,N_14398,N_12191);
nand U25954 (N_25954,N_16179,N_18634);
xor U25955 (N_25955,N_16046,N_10791);
nor U25956 (N_25956,N_17676,N_16633);
nor U25957 (N_25957,N_14473,N_10797);
and U25958 (N_25958,N_15895,N_11725);
and U25959 (N_25959,N_15143,N_16148);
nor U25960 (N_25960,N_15222,N_18884);
or U25961 (N_25961,N_14517,N_13065);
nor U25962 (N_25962,N_13153,N_10514);
nand U25963 (N_25963,N_10195,N_19158);
and U25964 (N_25964,N_11046,N_10277);
xnor U25965 (N_25965,N_14306,N_19160);
or U25966 (N_25966,N_19532,N_13399);
nand U25967 (N_25967,N_13716,N_10726);
nand U25968 (N_25968,N_12867,N_19052);
nand U25969 (N_25969,N_13482,N_16701);
nor U25970 (N_25970,N_16030,N_16390);
and U25971 (N_25971,N_11156,N_14113);
and U25972 (N_25972,N_19728,N_12018);
xnor U25973 (N_25973,N_12364,N_15615);
nor U25974 (N_25974,N_14524,N_12557);
nor U25975 (N_25975,N_15591,N_11579);
or U25976 (N_25976,N_14383,N_16706);
or U25977 (N_25977,N_19409,N_11268);
and U25978 (N_25978,N_10777,N_14922);
nor U25979 (N_25979,N_16702,N_14859);
or U25980 (N_25980,N_13429,N_18057);
and U25981 (N_25981,N_11526,N_18128);
nor U25982 (N_25982,N_12218,N_18912);
xnor U25983 (N_25983,N_15173,N_12745);
xnor U25984 (N_25984,N_17579,N_19576);
and U25985 (N_25985,N_13717,N_11374);
or U25986 (N_25986,N_14848,N_18629);
or U25987 (N_25987,N_11001,N_11970);
and U25988 (N_25988,N_18190,N_13965);
and U25989 (N_25989,N_12440,N_18785);
nand U25990 (N_25990,N_17178,N_10406);
nand U25991 (N_25991,N_19955,N_17222);
nor U25992 (N_25992,N_13488,N_13939);
nor U25993 (N_25993,N_15506,N_13657);
nand U25994 (N_25994,N_11661,N_10909);
nand U25995 (N_25995,N_11795,N_16140);
xor U25996 (N_25996,N_10134,N_10866);
or U25997 (N_25997,N_17102,N_15631);
nand U25998 (N_25998,N_11035,N_16845);
nand U25999 (N_25999,N_11231,N_16319);
xor U26000 (N_26000,N_14846,N_18857);
and U26001 (N_26001,N_14545,N_13801);
and U26002 (N_26002,N_16353,N_11283);
nor U26003 (N_26003,N_19229,N_13980);
xnor U26004 (N_26004,N_19602,N_17473);
and U26005 (N_26005,N_10957,N_16054);
nor U26006 (N_26006,N_12226,N_13500);
and U26007 (N_26007,N_13276,N_15446);
and U26008 (N_26008,N_11349,N_13158);
nand U26009 (N_26009,N_11641,N_11126);
or U26010 (N_26010,N_13253,N_14282);
nand U26011 (N_26011,N_16666,N_10067);
and U26012 (N_26012,N_16621,N_11388);
nor U26013 (N_26013,N_19416,N_16929);
or U26014 (N_26014,N_13994,N_14045);
nand U26015 (N_26015,N_16572,N_13156);
xnor U26016 (N_26016,N_17961,N_12330);
nor U26017 (N_26017,N_14497,N_12125);
and U26018 (N_26018,N_15777,N_12621);
nand U26019 (N_26019,N_15324,N_16867);
nand U26020 (N_26020,N_12216,N_11844);
or U26021 (N_26021,N_19688,N_10956);
nor U26022 (N_26022,N_14702,N_14959);
nor U26023 (N_26023,N_13763,N_16103);
or U26024 (N_26024,N_18676,N_19203);
and U26025 (N_26025,N_18279,N_12923);
nor U26026 (N_26026,N_11736,N_16737);
nor U26027 (N_26027,N_10217,N_19598);
nor U26028 (N_26028,N_18130,N_12626);
nor U26029 (N_26029,N_11515,N_14017);
or U26030 (N_26030,N_14431,N_15688);
or U26031 (N_26031,N_10368,N_15084);
xor U26032 (N_26032,N_13315,N_13377);
nand U26033 (N_26033,N_11664,N_10060);
and U26034 (N_26034,N_14753,N_13595);
or U26035 (N_26035,N_12979,N_15004);
xnor U26036 (N_26036,N_15394,N_15711);
or U26037 (N_26037,N_12094,N_16056);
and U26038 (N_26038,N_14816,N_15688);
xnor U26039 (N_26039,N_17685,N_13288);
nor U26040 (N_26040,N_15255,N_15319);
nand U26041 (N_26041,N_12957,N_16412);
nor U26042 (N_26042,N_18496,N_12983);
and U26043 (N_26043,N_12998,N_19915);
or U26044 (N_26044,N_15472,N_11493);
nor U26045 (N_26045,N_13964,N_19953);
and U26046 (N_26046,N_16428,N_12109);
nand U26047 (N_26047,N_11493,N_13462);
nor U26048 (N_26048,N_15532,N_17723);
nand U26049 (N_26049,N_10287,N_14286);
or U26050 (N_26050,N_13972,N_15731);
nor U26051 (N_26051,N_11696,N_16055);
nor U26052 (N_26052,N_15147,N_13090);
and U26053 (N_26053,N_19980,N_11283);
or U26054 (N_26054,N_10065,N_17485);
or U26055 (N_26055,N_10829,N_11059);
and U26056 (N_26056,N_16436,N_13170);
nor U26057 (N_26057,N_15517,N_14395);
and U26058 (N_26058,N_18535,N_12581);
nor U26059 (N_26059,N_12518,N_18813);
or U26060 (N_26060,N_11672,N_10047);
or U26061 (N_26061,N_16081,N_13691);
nand U26062 (N_26062,N_14146,N_11848);
and U26063 (N_26063,N_19201,N_13008);
xor U26064 (N_26064,N_11910,N_13096);
nor U26065 (N_26065,N_10799,N_18703);
or U26066 (N_26066,N_13090,N_13119);
xor U26067 (N_26067,N_19130,N_17411);
nand U26068 (N_26068,N_19842,N_11135);
and U26069 (N_26069,N_12518,N_12340);
nand U26070 (N_26070,N_16040,N_18146);
and U26071 (N_26071,N_17192,N_10303);
or U26072 (N_26072,N_15924,N_11668);
nand U26073 (N_26073,N_11406,N_13868);
nor U26074 (N_26074,N_14057,N_18501);
or U26075 (N_26075,N_17642,N_13682);
and U26076 (N_26076,N_11417,N_19829);
xor U26077 (N_26077,N_12392,N_15895);
nand U26078 (N_26078,N_18167,N_19824);
or U26079 (N_26079,N_10250,N_11913);
nand U26080 (N_26080,N_13921,N_10808);
nand U26081 (N_26081,N_13866,N_10221);
or U26082 (N_26082,N_11029,N_19528);
and U26083 (N_26083,N_11836,N_13394);
or U26084 (N_26084,N_17550,N_14580);
xnor U26085 (N_26085,N_18184,N_19838);
nand U26086 (N_26086,N_11323,N_11578);
or U26087 (N_26087,N_13489,N_18096);
xnor U26088 (N_26088,N_19374,N_17874);
or U26089 (N_26089,N_19464,N_16711);
nand U26090 (N_26090,N_13534,N_14341);
or U26091 (N_26091,N_10525,N_11215);
nor U26092 (N_26092,N_10257,N_19474);
or U26093 (N_26093,N_10753,N_11210);
and U26094 (N_26094,N_18347,N_11400);
nand U26095 (N_26095,N_16528,N_17223);
nor U26096 (N_26096,N_18161,N_15503);
nand U26097 (N_26097,N_12606,N_12751);
nand U26098 (N_26098,N_17718,N_13816);
nor U26099 (N_26099,N_14677,N_14062);
xor U26100 (N_26100,N_10809,N_12902);
nand U26101 (N_26101,N_14369,N_16586);
and U26102 (N_26102,N_10127,N_12782);
nand U26103 (N_26103,N_12450,N_11375);
or U26104 (N_26104,N_15018,N_10146);
and U26105 (N_26105,N_16961,N_17490);
or U26106 (N_26106,N_10617,N_13172);
or U26107 (N_26107,N_15080,N_13680);
nand U26108 (N_26108,N_14360,N_12220);
nor U26109 (N_26109,N_18589,N_12265);
xnor U26110 (N_26110,N_15034,N_19483);
or U26111 (N_26111,N_11173,N_13043);
nand U26112 (N_26112,N_10825,N_10894);
nand U26113 (N_26113,N_16066,N_11645);
or U26114 (N_26114,N_19604,N_12628);
nor U26115 (N_26115,N_13660,N_15497);
and U26116 (N_26116,N_16274,N_15736);
nor U26117 (N_26117,N_11620,N_18469);
or U26118 (N_26118,N_15953,N_19101);
nor U26119 (N_26119,N_13318,N_16379);
xnor U26120 (N_26120,N_18637,N_19681);
or U26121 (N_26121,N_14266,N_10677);
and U26122 (N_26122,N_19227,N_19278);
nand U26123 (N_26123,N_11292,N_19351);
and U26124 (N_26124,N_10895,N_13225);
and U26125 (N_26125,N_11652,N_17289);
nor U26126 (N_26126,N_16020,N_14330);
and U26127 (N_26127,N_16928,N_18617);
nand U26128 (N_26128,N_14492,N_14883);
nand U26129 (N_26129,N_10642,N_14166);
and U26130 (N_26130,N_12779,N_16951);
xor U26131 (N_26131,N_17438,N_18779);
or U26132 (N_26132,N_13107,N_15178);
and U26133 (N_26133,N_12592,N_12873);
nand U26134 (N_26134,N_12901,N_15492);
or U26135 (N_26135,N_14493,N_18099);
nor U26136 (N_26136,N_10340,N_18282);
nand U26137 (N_26137,N_12567,N_12865);
and U26138 (N_26138,N_15492,N_13350);
or U26139 (N_26139,N_18250,N_17972);
or U26140 (N_26140,N_10343,N_10354);
and U26141 (N_26141,N_12347,N_11504);
nor U26142 (N_26142,N_18232,N_19786);
and U26143 (N_26143,N_13588,N_13647);
nor U26144 (N_26144,N_18162,N_13294);
xor U26145 (N_26145,N_10863,N_11067);
xnor U26146 (N_26146,N_19297,N_11216);
or U26147 (N_26147,N_12350,N_14481);
or U26148 (N_26148,N_12409,N_12255);
nor U26149 (N_26149,N_17414,N_14764);
nand U26150 (N_26150,N_12642,N_15603);
or U26151 (N_26151,N_16171,N_12465);
or U26152 (N_26152,N_12571,N_13585);
nand U26153 (N_26153,N_15461,N_12867);
or U26154 (N_26154,N_14452,N_13272);
or U26155 (N_26155,N_10386,N_15211);
and U26156 (N_26156,N_11265,N_11115);
xor U26157 (N_26157,N_13504,N_13149);
or U26158 (N_26158,N_13980,N_10170);
and U26159 (N_26159,N_11502,N_10869);
xnor U26160 (N_26160,N_14693,N_17410);
xor U26161 (N_26161,N_11680,N_19583);
nor U26162 (N_26162,N_17466,N_17737);
nor U26163 (N_26163,N_12436,N_15562);
or U26164 (N_26164,N_16196,N_17858);
or U26165 (N_26165,N_19695,N_11083);
and U26166 (N_26166,N_14280,N_13385);
and U26167 (N_26167,N_10457,N_13743);
nand U26168 (N_26168,N_10334,N_19893);
nor U26169 (N_26169,N_16672,N_12662);
nor U26170 (N_26170,N_12914,N_16276);
xnor U26171 (N_26171,N_19037,N_17088);
and U26172 (N_26172,N_17050,N_10785);
nand U26173 (N_26173,N_17520,N_10479);
nor U26174 (N_26174,N_18516,N_13279);
nand U26175 (N_26175,N_13839,N_18711);
nor U26176 (N_26176,N_17404,N_17624);
and U26177 (N_26177,N_18591,N_19074);
xnor U26178 (N_26178,N_19254,N_17187);
or U26179 (N_26179,N_19136,N_14414);
nand U26180 (N_26180,N_12191,N_12565);
nand U26181 (N_26181,N_19876,N_10245);
xor U26182 (N_26182,N_19059,N_14078);
xnor U26183 (N_26183,N_14994,N_17311);
nand U26184 (N_26184,N_11698,N_16786);
or U26185 (N_26185,N_10811,N_19258);
or U26186 (N_26186,N_12197,N_18187);
nor U26187 (N_26187,N_19935,N_10853);
and U26188 (N_26188,N_15324,N_11832);
or U26189 (N_26189,N_19321,N_18029);
nor U26190 (N_26190,N_18464,N_13448);
or U26191 (N_26191,N_19646,N_17422);
and U26192 (N_26192,N_17964,N_14935);
nor U26193 (N_26193,N_16546,N_16629);
and U26194 (N_26194,N_14655,N_19038);
and U26195 (N_26195,N_15831,N_13498);
and U26196 (N_26196,N_10439,N_19882);
nor U26197 (N_26197,N_13221,N_12411);
nor U26198 (N_26198,N_17187,N_18796);
nand U26199 (N_26199,N_18828,N_16538);
nand U26200 (N_26200,N_12080,N_12391);
or U26201 (N_26201,N_13276,N_11684);
and U26202 (N_26202,N_10355,N_15551);
nor U26203 (N_26203,N_14934,N_13828);
and U26204 (N_26204,N_11461,N_18566);
nand U26205 (N_26205,N_10588,N_15725);
nor U26206 (N_26206,N_19506,N_11767);
nand U26207 (N_26207,N_11094,N_18511);
and U26208 (N_26208,N_11519,N_14136);
xnor U26209 (N_26209,N_16772,N_16830);
and U26210 (N_26210,N_18696,N_18530);
nand U26211 (N_26211,N_11325,N_16251);
or U26212 (N_26212,N_17657,N_16254);
and U26213 (N_26213,N_19188,N_14993);
nand U26214 (N_26214,N_12215,N_18487);
nor U26215 (N_26215,N_11399,N_18761);
or U26216 (N_26216,N_12533,N_16370);
or U26217 (N_26217,N_14013,N_19804);
or U26218 (N_26218,N_13754,N_15551);
and U26219 (N_26219,N_13334,N_12746);
or U26220 (N_26220,N_15169,N_12740);
nor U26221 (N_26221,N_15360,N_15374);
nand U26222 (N_26222,N_13604,N_17902);
nand U26223 (N_26223,N_19115,N_11295);
nand U26224 (N_26224,N_13132,N_13563);
and U26225 (N_26225,N_14527,N_10902);
and U26226 (N_26226,N_15633,N_17551);
and U26227 (N_26227,N_10483,N_13156);
or U26228 (N_26228,N_18199,N_16644);
and U26229 (N_26229,N_15548,N_18672);
nand U26230 (N_26230,N_14707,N_10598);
and U26231 (N_26231,N_12560,N_16844);
and U26232 (N_26232,N_13242,N_11840);
nor U26233 (N_26233,N_13193,N_18292);
xnor U26234 (N_26234,N_12031,N_11431);
nand U26235 (N_26235,N_10397,N_11035);
and U26236 (N_26236,N_14705,N_12395);
and U26237 (N_26237,N_19936,N_14370);
xnor U26238 (N_26238,N_14272,N_11571);
or U26239 (N_26239,N_11149,N_12103);
nand U26240 (N_26240,N_12120,N_15826);
nand U26241 (N_26241,N_11276,N_11140);
or U26242 (N_26242,N_16831,N_16615);
nand U26243 (N_26243,N_16239,N_16919);
nand U26244 (N_26244,N_10725,N_12346);
nor U26245 (N_26245,N_15651,N_19602);
or U26246 (N_26246,N_14592,N_17197);
nor U26247 (N_26247,N_14444,N_16416);
xor U26248 (N_26248,N_10939,N_13664);
nand U26249 (N_26249,N_10550,N_11458);
or U26250 (N_26250,N_10343,N_14953);
or U26251 (N_26251,N_19900,N_15692);
nand U26252 (N_26252,N_16445,N_13064);
and U26253 (N_26253,N_19721,N_19459);
nor U26254 (N_26254,N_16522,N_12223);
and U26255 (N_26255,N_10714,N_13468);
nor U26256 (N_26256,N_10948,N_12835);
and U26257 (N_26257,N_12613,N_12840);
nor U26258 (N_26258,N_15946,N_13126);
nand U26259 (N_26259,N_16926,N_18325);
nand U26260 (N_26260,N_13642,N_13644);
nand U26261 (N_26261,N_14344,N_19949);
xnor U26262 (N_26262,N_12905,N_16898);
nor U26263 (N_26263,N_13545,N_12774);
nand U26264 (N_26264,N_10907,N_18493);
xnor U26265 (N_26265,N_10731,N_17093);
nor U26266 (N_26266,N_10337,N_13365);
nand U26267 (N_26267,N_19937,N_11375);
and U26268 (N_26268,N_12481,N_16707);
nand U26269 (N_26269,N_16348,N_17755);
and U26270 (N_26270,N_15970,N_19871);
or U26271 (N_26271,N_18447,N_19493);
or U26272 (N_26272,N_14279,N_17298);
nand U26273 (N_26273,N_18761,N_12680);
nor U26274 (N_26274,N_13766,N_17084);
and U26275 (N_26275,N_13425,N_16332);
xnor U26276 (N_26276,N_18886,N_18102);
xnor U26277 (N_26277,N_17604,N_16296);
or U26278 (N_26278,N_12310,N_17351);
and U26279 (N_26279,N_13578,N_12391);
or U26280 (N_26280,N_18086,N_18650);
nand U26281 (N_26281,N_17661,N_14987);
or U26282 (N_26282,N_15713,N_14961);
nand U26283 (N_26283,N_17934,N_15571);
nor U26284 (N_26284,N_19839,N_19252);
or U26285 (N_26285,N_19426,N_17697);
and U26286 (N_26286,N_19022,N_15694);
and U26287 (N_26287,N_18168,N_14919);
nor U26288 (N_26288,N_12952,N_14554);
and U26289 (N_26289,N_17987,N_11040);
xnor U26290 (N_26290,N_15892,N_18875);
and U26291 (N_26291,N_16957,N_16923);
and U26292 (N_26292,N_13437,N_12270);
nor U26293 (N_26293,N_13543,N_13003);
and U26294 (N_26294,N_16287,N_11150);
and U26295 (N_26295,N_11600,N_18223);
or U26296 (N_26296,N_19386,N_14149);
and U26297 (N_26297,N_10035,N_13570);
or U26298 (N_26298,N_19276,N_19133);
xnor U26299 (N_26299,N_14518,N_18315);
or U26300 (N_26300,N_16455,N_13288);
nor U26301 (N_26301,N_11437,N_14599);
or U26302 (N_26302,N_16231,N_12622);
or U26303 (N_26303,N_19471,N_10762);
or U26304 (N_26304,N_11489,N_15606);
nand U26305 (N_26305,N_16213,N_14577);
and U26306 (N_26306,N_12042,N_11358);
or U26307 (N_26307,N_12652,N_17701);
nor U26308 (N_26308,N_12181,N_18891);
xor U26309 (N_26309,N_11302,N_18339);
nand U26310 (N_26310,N_15629,N_10213);
or U26311 (N_26311,N_11908,N_16890);
nor U26312 (N_26312,N_12267,N_11783);
and U26313 (N_26313,N_14074,N_17651);
or U26314 (N_26314,N_15292,N_16232);
and U26315 (N_26315,N_11904,N_16679);
nor U26316 (N_26316,N_14677,N_13174);
and U26317 (N_26317,N_17338,N_15426);
nor U26318 (N_26318,N_12453,N_17420);
and U26319 (N_26319,N_16429,N_17296);
nor U26320 (N_26320,N_12095,N_16136);
nand U26321 (N_26321,N_19475,N_14575);
xor U26322 (N_26322,N_14683,N_11249);
or U26323 (N_26323,N_17514,N_19288);
nor U26324 (N_26324,N_15442,N_19928);
nand U26325 (N_26325,N_14389,N_12011);
nand U26326 (N_26326,N_13276,N_17379);
nand U26327 (N_26327,N_14695,N_14315);
or U26328 (N_26328,N_15181,N_18887);
or U26329 (N_26329,N_14865,N_17151);
or U26330 (N_26330,N_11992,N_18537);
nand U26331 (N_26331,N_18198,N_10007);
or U26332 (N_26332,N_18058,N_16570);
or U26333 (N_26333,N_10895,N_16126);
and U26334 (N_26334,N_11341,N_11143);
and U26335 (N_26335,N_18083,N_10514);
or U26336 (N_26336,N_16787,N_17888);
or U26337 (N_26337,N_12381,N_11629);
or U26338 (N_26338,N_15936,N_11610);
nor U26339 (N_26339,N_18394,N_19704);
nand U26340 (N_26340,N_18964,N_10581);
and U26341 (N_26341,N_19790,N_12616);
and U26342 (N_26342,N_18393,N_15754);
nand U26343 (N_26343,N_11893,N_13690);
nand U26344 (N_26344,N_14040,N_16560);
nor U26345 (N_26345,N_18946,N_16985);
xor U26346 (N_26346,N_10184,N_18076);
nor U26347 (N_26347,N_10190,N_15226);
and U26348 (N_26348,N_15719,N_18757);
nand U26349 (N_26349,N_17194,N_14612);
nand U26350 (N_26350,N_15961,N_15441);
nor U26351 (N_26351,N_11993,N_13262);
nand U26352 (N_26352,N_17160,N_15876);
nand U26353 (N_26353,N_15651,N_19251);
and U26354 (N_26354,N_10895,N_12759);
nor U26355 (N_26355,N_18598,N_19426);
or U26356 (N_26356,N_11178,N_16573);
or U26357 (N_26357,N_18477,N_15035);
and U26358 (N_26358,N_16167,N_15732);
or U26359 (N_26359,N_13929,N_16595);
and U26360 (N_26360,N_13294,N_18146);
and U26361 (N_26361,N_17610,N_14209);
nand U26362 (N_26362,N_14763,N_14839);
and U26363 (N_26363,N_18279,N_15427);
or U26364 (N_26364,N_17320,N_11941);
nand U26365 (N_26365,N_15575,N_12801);
or U26366 (N_26366,N_17664,N_16437);
nand U26367 (N_26367,N_13626,N_14679);
nor U26368 (N_26368,N_10601,N_17196);
nor U26369 (N_26369,N_18118,N_14303);
nor U26370 (N_26370,N_16058,N_12976);
nand U26371 (N_26371,N_12685,N_13019);
or U26372 (N_26372,N_14237,N_10909);
nor U26373 (N_26373,N_11078,N_13366);
and U26374 (N_26374,N_19484,N_16721);
or U26375 (N_26375,N_18469,N_19424);
nor U26376 (N_26376,N_19457,N_19432);
nor U26377 (N_26377,N_16645,N_10730);
or U26378 (N_26378,N_13915,N_19596);
xor U26379 (N_26379,N_10344,N_14509);
nand U26380 (N_26380,N_16086,N_17625);
nand U26381 (N_26381,N_10080,N_10843);
nor U26382 (N_26382,N_16335,N_12868);
or U26383 (N_26383,N_15665,N_18680);
and U26384 (N_26384,N_14593,N_18584);
nor U26385 (N_26385,N_14708,N_11542);
nor U26386 (N_26386,N_14187,N_19517);
nor U26387 (N_26387,N_14283,N_10893);
nand U26388 (N_26388,N_18770,N_16434);
or U26389 (N_26389,N_17480,N_19423);
nor U26390 (N_26390,N_13537,N_12254);
nor U26391 (N_26391,N_17812,N_12844);
or U26392 (N_26392,N_11369,N_19106);
or U26393 (N_26393,N_18485,N_10774);
nor U26394 (N_26394,N_14229,N_13921);
and U26395 (N_26395,N_15469,N_11225);
and U26396 (N_26396,N_18769,N_14126);
or U26397 (N_26397,N_14508,N_17052);
xnor U26398 (N_26398,N_17340,N_10081);
nor U26399 (N_26399,N_14929,N_12264);
nand U26400 (N_26400,N_16145,N_18876);
and U26401 (N_26401,N_11262,N_14280);
or U26402 (N_26402,N_15511,N_17007);
or U26403 (N_26403,N_14840,N_11147);
and U26404 (N_26404,N_11305,N_19413);
or U26405 (N_26405,N_10053,N_17121);
xnor U26406 (N_26406,N_17227,N_12719);
and U26407 (N_26407,N_12758,N_19204);
or U26408 (N_26408,N_10941,N_11570);
nand U26409 (N_26409,N_14376,N_12505);
xor U26410 (N_26410,N_11459,N_12358);
nor U26411 (N_26411,N_17725,N_13931);
or U26412 (N_26412,N_12701,N_18930);
and U26413 (N_26413,N_19797,N_11019);
nand U26414 (N_26414,N_15770,N_11032);
and U26415 (N_26415,N_10890,N_13526);
xnor U26416 (N_26416,N_17899,N_18126);
nor U26417 (N_26417,N_17147,N_13942);
and U26418 (N_26418,N_10150,N_16367);
or U26419 (N_26419,N_15428,N_14140);
and U26420 (N_26420,N_14372,N_19222);
nor U26421 (N_26421,N_11457,N_11851);
nor U26422 (N_26422,N_15398,N_15973);
or U26423 (N_26423,N_18009,N_10633);
or U26424 (N_26424,N_16980,N_12529);
and U26425 (N_26425,N_11346,N_11717);
or U26426 (N_26426,N_13648,N_14936);
xor U26427 (N_26427,N_13876,N_13771);
nor U26428 (N_26428,N_10498,N_19767);
and U26429 (N_26429,N_15878,N_19346);
nor U26430 (N_26430,N_17773,N_11265);
nor U26431 (N_26431,N_12205,N_18256);
nand U26432 (N_26432,N_11498,N_13485);
or U26433 (N_26433,N_11699,N_15730);
xnor U26434 (N_26434,N_16704,N_17653);
or U26435 (N_26435,N_18711,N_13568);
or U26436 (N_26436,N_14779,N_12565);
or U26437 (N_26437,N_11795,N_14659);
nor U26438 (N_26438,N_10074,N_15221);
or U26439 (N_26439,N_15983,N_12944);
nor U26440 (N_26440,N_18612,N_12361);
and U26441 (N_26441,N_16158,N_12627);
nand U26442 (N_26442,N_18371,N_17793);
xor U26443 (N_26443,N_10561,N_11330);
nand U26444 (N_26444,N_10277,N_10129);
xor U26445 (N_26445,N_15431,N_15292);
and U26446 (N_26446,N_16590,N_15721);
and U26447 (N_26447,N_16377,N_11522);
nor U26448 (N_26448,N_10963,N_10880);
nand U26449 (N_26449,N_11226,N_15428);
nand U26450 (N_26450,N_19611,N_12424);
xnor U26451 (N_26451,N_16426,N_12166);
xor U26452 (N_26452,N_11306,N_19666);
xor U26453 (N_26453,N_19925,N_16564);
or U26454 (N_26454,N_15467,N_15722);
xor U26455 (N_26455,N_14268,N_14926);
or U26456 (N_26456,N_11192,N_19244);
nor U26457 (N_26457,N_17643,N_17630);
or U26458 (N_26458,N_13968,N_12414);
nor U26459 (N_26459,N_13611,N_14498);
nand U26460 (N_26460,N_16839,N_15217);
nand U26461 (N_26461,N_13106,N_11344);
or U26462 (N_26462,N_18336,N_19723);
nand U26463 (N_26463,N_16170,N_17535);
nor U26464 (N_26464,N_11517,N_16499);
and U26465 (N_26465,N_17220,N_15671);
nand U26466 (N_26466,N_19402,N_14262);
and U26467 (N_26467,N_11097,N_12787);
nand U26468 (N_26468,N_10235,N_13402);
and U26469 (N_26469,N_16685,N_19424);
nor U26470 (N_26470,N_10440,N_16539);
nor U26471 (N_26471,N_12816,N_17826);
or U26472 (N_26472,N_19273,N_19231);
or U26473 (N_26473,N_14672,N_16467);
or U26474 (N_26474,N_15234,N_19590);
or U26475 (N_26475,N_19298,N_11712);
nor U26476 (N_26476,N_17620,N_10359);
nand U26477 (N_26477,N_18993,N_11003);
and U26478 (N_26478,N_15750,N_14974);
or U26479 (N_26479,N_15634,N_11486);
and U26480 (N_26480,N_12961,N_10892);
or U26481 (N_26481,N_11126,N_13736);
or U26482 (N_26482,N_16527,N_13215);
and U26483 (N_26483,N_16020,N_12151);
or U26484 (N_26484,N_16228,N_13717);
and U26485 (N_26485,N_14574,N_13040);
nand U26486 (N_26486,N_18199,N_12742);
or U26487 (N_26487,N_13129,N_17772);
nand U26488 (N_26488,N_16241,N_11003);
nor U26489 (N_26489,N_12625,N_18843);
nor U26490 (N_26490,N_13729,N_17242);
or U26491 (N_26491,N_16510,N_13170);
or U26492 (N_26492,N_19831,N_14243);
nand U26493 (N_26493,N_16596,N_14239);
xor U26494 (N_26494,N_12115,N_14501);
nor U26495 (N_26495,N_14755,N_11376);
nor U26496 (N_26496,N_12318,N_17395);
or U26497 (N_26497,N_14699,N_10002);
nor U26498 (N_26498,N_12669,N_13081);
nand U26499 (N_26499,N_16903,N_18932);
nand U26500 (N_26500,N_10199,N_17692);
or U26501 (N_26501,N_10779,N_13178);
nor U26502 (N_26502,N_16187,N_11126);
nor U26503 (N_26503,N_13559,N_13095);
or U26504 (N_26504,N_12620,N_15753);
and U26505 (N_26505,N_19693,N_18938);
or U26506 (N_26506,N_11344,N_13233);
nand U26507 (N_26507,N_19829,N_13998);
and U26508 (N_26508,N_10898,N_11689);
or U26509 (N_26509,N_12887,N_15038);
and U26510 (N_26510,N_15405,N_16632);
or U26511 (N_26511,N_12442,N_15856);
nor U26512 (N_26512,N_13945,N_14644);
and U26513 (N_26513,N_11903,N_19363);
or U26514 (N_26514,N_12743,N_17914);
or U26515 (N_26515,N_19731,N_12068);
and U26516 (N_26516,N_14744,N_13522);
nand U26517 (N_26517,N_18324,N_10163);
or U26518 (N_26518,N_15640,N_10070);
xnor U26519 (N_26519,N_10701,N_15753);
nor U26520 (N_26520,N_13515,N_19708);
or U26521 (N_26521,N_15860,N_18862);
xnor U26522 (N_26522,N_11570,N_11762);
or U26523 (N_26523,N_14880,N_11050);
nor U26524 (N_26524,N_17790,N_12153);
and U26525 (N_26525,N_13759,N_11521);
and U26526 (N_26526,N_12974,N_11010);
nor U26527 (N_26527,N_10658,N_10959);
and U26528 (N_26528,N_13660,N_15449);
nand U26529 (N_26529,N_11850,N_13022);
or U26530 (N_26530,N_16520,N_17675);
nor U26531 (N_26531,N_18035,N_16061);
or U26532 (N_26532,N_19917,N_17468);
or U26533 (N_26533,N_12441,N_17189);
nand U26534 (N_26534,N_14245,N_15241);
or U26535 (N_26535,N_12333,N_10456);
or U26536 (N_26536,N_13677,N_12333);
nor U26537 (N_26537,N_17999,N_17507);
and U26538 (N_26538,N_12044,N_17186);
xnor U26539 (N_26539,N_12725,N_18172);
and U26540 (N_26540,N_14216,N_12922);
nor U26541 (N_26541,N_19682,N_16635);
or U26542 (N_26542,N_14352,N_19347);
nor U26543 (N_26543,N_19265,N_11808);
nor U26544 (N_26544,N_15799,N_19470);
and U26545 (N_26545,N_10903,N_17839);
and U26546 (N_26546,N_16312,N_13048);
nor U26547 (N_26547,N_10297,N_17470);
and U26548 (N_26548,N_10813,N_18815);
and U26549 (N_26549,N_10208,N_18284);
and U26550 (N_26550,N_12183,N_15370);
or U26551 (N_26551,N_11174,N_14880);
nor U26552 (N_26552,N_15109,N_10365);
or U26553 (N_26553,N_11070,N_13013);
nor U26554 (N_26554,N_15312,N_18988);
nand U26555 (N_26555,N_12931,N_11376);
nor U26556 (N_26556,N_16551,N_13612);
nor U26557 (N_26557,N_18592,N_11873);
and U26558 (N_26558,N_12403,N_14052);
or U26559 (N_26559,N_16958,N_11494);
or U26560 (N_26560,N_18246,N_19634);
or U26561 (N_26561,N_11717,N_12848);
nor U26562 (N_26562,N_11832,N_13538);
nor U26563 (N_26563,N_11369,N_10116);
and U26564 (N_26564,N_17178,N_15707);
or U26565 (N_26565,N_18175,N_10548);
and U26566 (N_26566,N_19120,N_18209);
and U26567 (N_26567,N_19392,N_14034);
xor U26568 (N_26568,N_18377,N_17567);
and U26569 (N_26569,N_18637,N_13373);
nor U26570 (N_26570,N_18516,N_19992);
nand U26571 (N_26571,N_19746,N_15616);
nand U26572 (N_26572,N_19499,N_11846);
nand U26573 (N_26573,N_19903,N_17884);
nand U26574 (N_26574,N_16524,N_17641);
nand U26575 (N_26575,N_19640,N_19590);
nor U26576 (N_26576,N_19946,N_14177);
and U26577 (N_26577,N_18259,N_11779);
nor U26578 (N_26578,N_12038,N_13237);
nand U26579 (N_26579,N_16421,N_14364);
nand U26580 (N_26580,N_16700,N_13788);
or U26581 (N_26581,N_14234,N_12164);
nand U26582 (N_26582,N_13131,N_15957);
nand U26583 (N_26583,N_15498,N_18305);
and U26584 (N_26584,N_19230,N_18261);
and U26585 (N_26585,N_15172,N_15526);
xnor U26586 (N_26586,N_13894,N_18753);
nor U26587 (N_26587,N_10838,N_19694);
nand U26588 (N_26588,N_11834,N_15271);
nand U26589 (N_26589,N_19864,N_16943);
nand U26590 (N_26590,N_10008,N_17383);
and U26591 (N_26591,N_11913,N_14868);
nor U26592 (N_26592,N_18011,N_14555);
xor U26593 (N_26593,N_13403,N_15047);
or U26594 (N_26594,N_15153,N_15999);
and U26595 (N_26595,N_14253,N_15278);
nor U26596 (N_26596,N_15884,N_10616);
xnor U26597 (N_26597,N_16360,N_19360);
or U26598 (N_26598,N_12079,N_19017);
and U26599 (N_26599,N_19515,N_10656);
nor U26600 (N_26600,N_17376,N_11773);
nand U26601 (N_26601,N_16883,N_12084);
nor U26602 (N_26602,N_19613,N_17293);
nor U26603 (N_26603,N_19228,N_15182);
and U26604 (N_26604,N_12749,N_16682);
and U26605 (N_26605,N_16155,N_11119);
or U26606 (N_26606,N_10648,N_14718);
nor U26607 (N_26607,N_17762,N_13633);
nor U26608 (N_26608,N_14596,N_14498);
and U26609 (N_26609,N_17324,N_17189);
nor U26610 (N_26610,N_18982,N_17391);
xnor U26611 (N_26611,N_14198,N_18606);
and U26612 (N_26612,N_16737,N_18766);
or U26613 (N_26613,N_19510,N_18997);
nor U26614 (N_26614,N_14915,N_14106);
and U26615 (N_26615,N_12179,N_13849);
and U26616 (N_26616,N_15065,N_15336);
nor U26617 (N_26617,N_16733,N_12778);
and U26618 (N_26618,N_11458,N_17978);
nand U26619 (N_26619,N_14264,N_16380);
nor U26620 (N_26620,N_11980,N_16108);
nor U26621 (N_26621,N_17208,N_16138);
nor U26622 (N_26622,N_10168,N_12253);
and U26623 (N_26623,N_13715,N_13792);
nor U26624 (N_26624,N_17885,N_18119);
nor U26625 (N_26625,N_12489,N_14735);
xnor U26626 (N_26626,N_14799,N_10278);
and U26627 (N_26627,N_11178,N_18752);
nand U26628 (N_26628,N_11313,N_19370);
nor U26629 (N_26629,N_12136,N_15814);
nor U26630 (N_26630,N_13646,N_18297);
and U26631 (N_26631,N_18723,N_12601);
nand U26632 (N_26632,N_13225,N_16873);
or U26633 (N_26633,N_19976,N_13876);
and U26634 (N_26634,N_17936,N_15162);
or U26635 (N_26635,N_12527,N_18021);
or U26636 (N_26636,N_14649,N_10403);
nor U26637 (N_26637,N_11447,N_10176);
nor U26638 (N_26638,N_13883,N_19110);
and U26639 (N_26639,N_11873,N_18673);
nor U26640 (N_26640,N_11407,N_16352);
nand U26641 (N_26641,N_14487,N_19703);
or U26642 (N_26642,N_14264,N_12749);
nand U26643 (N_26643,N_15420,N_16692);
or U26644 (N_26644,N_18669,N_10618);
nand U26645 (N_26645,N_19766,N_18464);
nand U26646 (N_26646,N_16775,N_15697);
nand U26647 (N_26647,N_18736,N_13426);
nand U26648 (N_26648,N_18883,N_12156);
nand U26649 (N_26649,N_13570,N_19200);
and U26650 (N_26650,N_17428,N_10175);
or U26651 (N_26651,N_17604,N_13475);
nor U26652 (N_26652,N_12015,N_14293);
nor U26653 (N_26653,N_12872,N_11402);
nand U26654 (N_26654,N_11622,N_19244);
nand U26655 (N_26655,N_15569,N_18853);
nand U26656 (N_26656,N_17196,N_12475);
nor U26657 (N_26657,N_12746,N_17152);
nand U26658 (N_26658,N_17391,N_16477);
and U26659 (N_26659,N_17342,N_16098);
nand U26660 (N_26660,N_12454,N_11270);
and U26661 (N_26661,N_16744,N_17063);
nor U26662 (N_26662,N_19497,N_10044);
nor U26663 (N_26663,N_19184,N_16569);
nand U26664 (N_26664,N_10952,N_11454);
nor U26665 (N_26665,N_11018,N_14374);
nor U26666 (N_26666,N_18558,N_16016);
or U26667 (N_26667,N_10753,N_15601);
or U26668 (N_26668,N_15713,N_19703);
or U26669 (N_26669,N_15653,N_19243);
nand U26670 (N_26670,N_17419,N_13662);
or U26671 (N_26671,N_17251,N_18202);
nand U26672 (N_26672,N_11175,N_11854);
and U26673 (N_26673,N_16862,N_17120);
and U26674 (N_26674,N_18840,N_17730);
or U26675 (N_26675,N_18437,N_19704);
nand U26676 (N_26676,N_11628,N_15895);
or U26677 (N_26677,N_15464,N_15075);
nand U26678 (N_26678,N_17043,N_16954);
nor U26679 (N_26679,N_12368,N_14183);
and U26680 (N_26680,N_16798,N_17427);
nor U26681 (N_26681,N_17998,N_11941);
xnor U26682 (N_26682,N_10096,N_10345);
nand U26683 (N_26683,N_17757,N_13298);
nand U26684 (N_26684,N_17480,N_19216);
xnor U26685 (N_26685,N_17649,N_11950);
nor U26686 (N_26686,N_13800,N_17246);
xnor U26687 (N_26687,N_12523,N_18962);
and U26688 (N_26688,N_12594,N_17326);
nor U26689 (N_26689,N_17550,N_11955);
or U26690 (N_26690,N_15590,N_10952);
nor U26691 (N_26691,N_13050,N_11240);
nand U26692 (N_26692,N_10920,N_12109);
nor U26693 (N_26693,N_11037,N_10758);
nand U26694 (N_26694,N_11952,N_19278);
nor U26695 (N_26695,N_11525,N_15459);
or U26696 (N_26696,N_10896,N_14071);
nor U26697 (N_26697,N_14356,N_12196);
nand U26698 (N_26698,N_16994,N_15023);
or U26699 (N_26699,N_16581,N_16154);
and U26700 (N_26700,N_15380,N_12144);
or U26701 (N_26701,N_17506,N_10840);
nor U26702 (N_26702,N_15439,N_19751);
or U26703 (N_26703,N_16271,N_19492);
xnor U26704 (N_26704,N_11379,N_19810);
nand U26705 (N_26705,N_12329,N_14338);
and U26706 (N_26706,N_18336,N_18724);
and U26707 (N_26707,N_17823,N_14244);
and U26708 (N_26708,N_17472,N_18234);
nand U26709 (N_26709,N_18953,N_11148);
nand U26710 (N_26710,N_11134,N_16088);
or U26711 (N_26711,N_16338,N_16144);
nand U26712 (N_26712,N_16455,N_17874);
and U26713 (N_26713,N_15455,N_19625);
and U26714 (N_26714,N_14740,N_17061);
nand U26715 (N_26715,N_16483,N_11761);
nor U26716 (N_26716,N_12242,N_10916);
xnor U26717 (N_26717,N_13929,N_12920);
nand U26718 (N_26718,N_14038,N_18351);
and U26719 (N_26719,N_17592,N_12883);
xnor U26720 (N_26720,N_13203,N_19310);
nand U26721 (N_26721,N_12185,N_17098);
nor U26722 (N_26722,N_17466,N_11807);
nor U26723 (N_26723,N_19660,N_13889);
nand U26724 (N_26724,N_13078,N_17226);
nor U26725 (N_26725,N_11892,N_18098);
nand U26726 (N_26726,N_11515,N_17325);
nand U26727 (N_26727,N_19023,N_11963);
or U26728 (N_26728,N_15817,N_19776);
or U26729 (N_26729,N_13555,N_17215);
and U26730 (N_26730,N_12006,N_14933);
or U26731 (N_26731,N_13561,N_14489);
nor U26732 (N_26732,N_15226,N_11999);
nor U26733 (N_26733,N_17445,N_12852);
or U26734 (N_26734,N_15851,N_12397);
and U26735 (N_26735,N_11536,N_14877);
nand U26736 (N_26736,N_16363,N_18997);
nor U26737 (N_26737,N_14015,N_10079);
nor U26738 (N_26738,N_15615,N_12832);
nor U26739 (N_26739,N_18294,N_15335);
and U26740 (N_26740,N_17172,N_15620);
nand U26741 (N_26741,N_10902,N_17465);
or U26742 (N_26742,N_11816,N_19401);
nor U26743 (N_26743,N_18791,N_15217);
nor U26744 (N_26744,N_17483,N_17989);
and U26745 (N_26745,N_18576,N_18263);
nand U26746 (N_26746,N_19684,N_16454);
nand U26747 (N_26747,N_17402,N_10379);
nor U26748 (N_26748,N_15688,N_12539);
and U26749 (N_26749,N_11586,N_16402);
nor U26750 (N_26750,N_13946,N_15772);
and U26751 (N_26751,N_10841,N_16717);
or U26752 (N_26752,N_15473,N_19711);
nor U26753 (N_26753,N_12552,N_11904);
nand U26754 (N_26754,N_19699,N_13002);
nand U26755 (N_26755,N_19911,N_17204);
and U26756 (N_26756,N_12478,N_13831);
nor U26757 (N_26757,N_18498,N_11887);
xor U26758 (N_26758,N_17617,N_17520);
and U26759 (N_26759,N_17094,N_19905);
nor U26760 (N_26760,N_18467,N_10725);
or U26761 (N_26761,N_14103,N_11661);
and U26762 (N_26762,N_11005,N_19184);
and U26763 (N_26763,N_13582,N_15888);
xnor U26764 (N_26764,N_17356,N_17030);
and U26765 (N_26765,N_14728,N_11903);
nand U26766 (N_26766,N_15445,N_11746);
and U26767 (N_26767,N_18405,N_11759);
or U26768 (N_26768,N_10870,N_17942);
nor U26769 (N_26769,N_18749,N_10611);
nand U26770 (N_26770,N_19059,N_18514);
nor U26771 (N_26771,N_14799,N_15784);
nor U26772 (N_26772,N_19647,N_15757);
nand U26773 (N_26773,N_18945,N_16925);
and U26774 (N_26774,N_12300,N_12782);
and U26775 (N_26775,N_10277,N_12461);
xor U26776 (N_26776,N_18183,N_19838);
xnor U26777 (N_26777,N_12394,N_11372);
or U26778 (N_26778,N_18859,N_19921);
nand U26779 (N_26779,N_19355,N_11504);
xnor U26780 (N_26780,N_14665,N_11701);
xor U26781 (N_26781,N_10432,N_16791);
and U26782 (N_26782,N_19857,N_12985);
xnor U26783 (N_26783,N_15100,N_19366);
xnor U26784 (N_26784,N_19310,N_18365);
or U26785 (N_26785,N_11998,N_14439);
or U26786 (N_26786,N_16055,N_15831);
nor U26787 (N_26787,N_10524,N_11961);
nand U26788 (N_26788,N_13442,N_16333);
or U26789 (N_26789,N_19930,N_10159);
nor U26790 (N_26790,N_15110,N_11065);
or U26791 (N_26791,N_18536,N_14125);
nand U26792 (N_26792,N_10365,N_15279);
xnor U26793 (N_26793,N_12623,N_12501);
nor U26794 (N_26794,N_12922,N_10927);
nor U26795 (N_26795,N_11329,N_18841);
or U26796 (N_26796,N_15923,N_10099);
nand U26797 (N_26797,N_10550,N_13865);
or U26798 (N_26798,N_19210,N_11311);
nand U26799 (N_26799,N_16950,N_13188);
xor U26800 (N_26800,N_16502,N_19863);
or U26801 (N_26801,N_15796,N_14625);
nand U26802 (N_26802,N_16295,N_10927);
nor U26803 (N_26803,N_17490,N_18356);
and U26804 (N_26804,N_13587,N_11871);
and U26805 (N_26805,N_19727,N_14803);
or U26806 (N_26806,N_14191,N_10634);
nand U26807 (N_26807,N_14156,N_16062);
nor U26808 (N_26808,N_18833,N_10629);
and U26809 (N_26809,N_19352,N_17728);
or U26810 (N_26810,N_18903,N_12332);
and U26811 (N_26811,N_19540,N_17880);
or U26812 (N_26812,N_17685,N_10449);
nand U26813 (N_26813,N_14428,N_18475);
and U26814 (N_26814,N_18193,N_14823);
or U26815 (N_26815,N_16635,N_13214);
nand U26816 (N_26816,N_11902,N_17112);
nor U26817 (N_26817,N_12959,N_10468);
nand U26818 (N_26818,N_16400,N_12075);
and U26819 (N_26819,N_16844,N_18263);
nand U26820 (N_26820,N_16531,N_18782);
nand U26821 (N_26821,N_11281,N_18783);
and U26822 (N_26822,N_15948,N_11933);
or U26823 (N_26823,N_10312,N_13898);
nor U26824 (N_26824,N_13727,N_18682);
nor U26825 (N_26825,N_18971,N_11103);
nor U26826 (N_26826,N_17178,N_16672);
or U26827 (N_26827,N_18821,N_13697);
or U26828 (N_26828,N_14349,N_15445);
xnor U26829 (N_26829,N_13785,N_10859);
and U26830 (N_26830,N_18998,N_10653);
nand U26831 (N_26831,N_14445,N_17298);
nand U26832 (N_26832,N_15942,N_18911);
and U26833 (N_26833,N_15856,N_19156);
nand U26834 (N_26834,N_10224,N_14577);
xor U26835 (N_26835,N_11962,N_15572);
nor U26836 (N_26836,N_11500,N_19717);
and U26837 (N_26837,N_19685,N_14809);
or U26838 (N_26838,N_18934,N_11432);
and U26839 (N_26839,N_12530,N_13525);
or U26840 (N_26840,N_13270,N_15566);
nor U26841 (N_26841,N_13257,N_11704);
and U26842 (N_26842,N_19806,N_12724);
nand U26843 (N_26843,N_11993,N_18582);
xor U26844 (N_26844,N_12405,N_16880);
or U26845 (N_26845,N_18347,N_14584);
nor U26846 (N_26846,N_16707,N_12801);
or U26847 (N_26847,N_12961,N_19075);
or U26848 (N_26848,N_13838,N_17350);
nor U26849 (N_26849,N_12164,N_17011);
nand U26850 (N_26850,N_18752,N_12239);
and U26851 (N_26851,N_16762,N_14251);
xnor U26852 (N_26852,N_13210,N_15482);
or U26853 (N_26853,N_19651,N_10433);
and U26854 (N_26854,N_17535,N_13921);
or U26855 (N_26855,N_18837,N_17901);
and U26856 (N_26856,N_11616,N_15179);
and U26857 (N_26857,N_15028,N_18027);
and U26858 (N_26858,N_16153,N_10963);
or U26859 (N_26859,N_16518,N_19925);
and U26860 (N_26860,N_13272,N_15387);
nand U26861 (N_26861,N_12686,N_16567);
nand U26862 (N_26862,N_19128,N_13027);
and U26863 (N_26863,N_14655,N_11377);
or U26864 (N_26864,N_14049,N_17957);
and U26865 (N_26865,N_15820,N_12838);
nor U26866 (N_26866,N_13266,N_10732);
or U26867 (N_26867,N_11104,N_12477);
and U26868 (N_26868,N_18429,N_11389);
and U26869 (N_26869,N_16757,N_18634);
and U26870 (N_26870,N_19851,N_15027);
or U26871 (N_26871,N_14619,N_14086);
or U26872 (N_26872,N_11971,N_19375);
nand U26873 (N_26873,N_10141,N_17658);
xnor U26874 (N_26874,N_18061,N_10654);
or U26875 (N_26875,N_18870,N_17218);
and U26876 (N_26876,N_17534,N_11698);
nand U26877 (N_26877,N_14325,N_17974);
nand U26878 (N_26878,N_15533,N_10880);
nand U26879 (N_26879,N_18350,N_11168);
and U26880 (N_26880,N_14459,N_14742);
nand U26881 (N_26881,N_13250,N_14464);
nor U26882 (N_26882,N_12664,N_15041);
and U26883 (N_26883,N_19485,N_18128);
nor U26884 (N_26884,N_19800,N_19859);
or U26885 (N_26885,N_10057,N_15556);
nor U26886 (N_26886,N_18303,N_15287);
nand U26887 (N_26887,N_11773,N_19692);
nand U26888 (N_26888,N_15260,N_13000);
nand U26889 (N_26889,N_14939,N_13935);
or U26890 (N_26890,N_17259,N_17700);
or U26891 (N_26891,N_18429,N_10087);
xor U26892 (N_26892,N_12252,N_11332);
or U26893 (N_26893,N_12302,N_14023);
nor U26894 (N_26894,N_15538,N_16357);
xor U26895 (N_26895,N_14998,N_10135);
and U26896 (N_26896,N_11182,N_11582);
nor U26897 (N_26897,N_19313,N_16627);
nor U26898 (N_26898,N_17717,N_16218);
nor U26899 (N_26899,N_19838,N_13350);
xnor U26900 (N_26900,N_18022,N_11447);
nor U26901 (N_26901,N_14739,N_17405);
nor U26902 (N_26902,N_15483,N_13116);
and U26903 (N_26903,N_11653,N_13865);
or U26904 (N_26904,N_15166,N_14008);
and U26905 (N_26905,N_10693,N_10108);
xnor U26906 (N_26906,N_15985,N_17507);
xnor U26907 (N_26907,N_17923,N_19456);
nor U26908 (N_26908,N_19111,N_17678);
and U26909 (N_26909,N_10235,N_11085);
and U26910 (N_26910,N_17782,N_13491);
or U26911 (N_26911,N_19452,N_15564);
or U26912 (N_26912,N_12303,N_14272);
and U26913 (N_26913,N_17040,N_11271);
nor U26914 (N_26914,N_12730,N_17915);
or U26915 (N_26915,N_18957,N_17131);
and U26916 (N_26916,N_11528,N_19128);
nand U26917 (N_26917,N_18824,N_16875);
nor U26918 (N_26918,N_11280,N_15028);
and U26919 (N_26919,N_17051,N_13927);
xor U26920 (N_26920,N_14419,N_15680);
nand U26921 (N_26921,N_10445,N_14666);
nor U26922 (N_26922,N_18176,N_19236);
and U26923 (N_26923,N_15793,N_14238);
nor U26924 (N_26924,N_17132,N_19803);
xnor U26925 (N_26925,N_15261,N_17899);
xnor U26926 (N_26926,N_17349,N_10111);
xnor U26927 (N_26927,N_19848,N_16223);
and U26928 (N_26928,N_14668,N_11793);
and U26929 (N_26929,N_19416,N_16934);
and U26930 (N_26930,N_18628,N_10438);
and U26931 (N_26931,N_15924,N_19198);
or U26932 (N_26932,N_11215,N_14693);
nor U26933 (N_26933,N_18364,N_11328);
nand U26934 (N_26934,N_11064,N_12935);
nor U26935 (N_26935,N_10965,N_17181);
xor U26936 (N_26936,N_16575,N_12249);
or U26937 (N_26937,N_16316,N_16745);
xnor U26938 (N_26938,N_14446,N_13446);
nor U26939 (N_26939,N_16226,N_15381);
or U26940 (N_26940,N_14772,N_17474);
nor U26941 (N_26941,N_15935,N_10710);
nand U26942 (N_26942,N_15678,N_11255);
and U26943 (N_26943,N_15677,N_18777);
xnor U26944 (N_26944,N_13583,N_18456);
or U26945 (N_26945,N_19460,N_18997);
nor U26946 (N_26946,N_12032,N_16430);
nor U26947 (N_26947,N_17053,N_14429);
nor U26948 (N_26948,N_13908,N_19881);
nor U26949 (N_26949,N_15597,N_15968);
nand U26950 (N_26950,N_18159,N_10371);
nor U26951 (N_26951,N_10460,N_16535);
or U26952 (N_26952,N_12320,N_12221);
nand U26953 (N_26953,N_13512,N_16673);
nand U26954 (N_26954,N_15447,N_18779);
nor U26955 (N_26955,N_14715,N_10338);
nand U26956 (N_26956,N_12389,N_16759);
or U26957 (N_26957,N_11210,N_12133);
nor U26958 (N_26958,N_14699,N_19352);
or U26959 (N_26959,N_14549,N_12189);
nor U26960 (N_26960,N_17360,N_17011);
nand U26961 (N_26961,N_15164,N_11317);
nand U26962 (N_26962,N_12417,N_10990);
nand U26963 (N_26963,N_19141,N_19879);
nand U26964 (N_26964,N_12886,N_17353);
and U26965 (N_26965,N_11743,N_17377);
or U26966 (N_26966,N_17699,N_14753);
nor U26967 (N_26967,N_16391,N_10701);
nand U26968 (N_26968,N_15173,N_17848);
and U26969 (N_26969,N_16630,N_14625);
or U26970 (N_26970,N_19045,N_17982);
or U26971 (N_26971,N_14553,N_18100);
nor U26972 (N_26972,N_19197,N_18369);
nor U26973 (N_26973,N_11207,N_10105);
nand U26974 (N_26974,N_12300,N_13347);
nand U26975 (N_26975,N_19697,N_18612);
or U26976 (N_26976,N_14369,N_11667);
nor U26977 (N_26977,N_17334,N_12144);
nand U26978 (N_26978,N_17850,N_18277);
nand U26979 (N_26979,N_15125,N_15402);
nor U26980 (N_26980,N_11930,N_18667);
and U26981 (N_26981,N_17060,N_19682);
nand U26982 (N_26982,N_10044,N_18726);
nand U26983 (N_26983,N_15745,N_18059);
and U26984 (N_26984,N_13277,N_10750);
nor U26985 (N_26985,N_17383,N_12352);
or U26986 (N_26986,N_13445,N_12594);
or U26987 (N_26987,N_18763,N_14744);
xnor U26988 (N_26988,N_14710,N_12654);
or U26989 (N_26989,N_17223,N_14356);
nand U26990 (N_26990,N_16154,N_18939);
nand U26991 (N_26991,N_16402,N_10588);
nand U26992 (N_26992,N_18505,N_18857);
nand U26993 (N_26993,N_16889,N_17406);
or U26994 (N_26994,N_16355,N_15314);
nand U26995 (N_26995,N_16271,N_16731);
nor U26996 (N_26996,N_17145,N_14501);
nand U26997 (N_26997,N_14777,N_12362);
nand U26998 (N_26998,N_18384,N_10488);
nor U26999 (N_26999,N_16231,N_10613);
nand U27000 (N_27000,N_18083,N_12639);
nor U27001 (N_27001,N_11163,N_13869);
or U27002 (N_27002,N_11119,N_18015);
xor U27003 (N_27003,N_15995,N_19954);
and U27004 (N_27004,N_12581,N_11608);
and U27005 (N_27005,N_14810,N_19489);
nand U27006 (N_27006,N_12358,N_19919);
and U27007 (N_27007,N_12732,N_16287);
or U27008 (N_27008,N_14035,N_11442);
nor U27009 (N_27009,N_14663,N_11830);
or U27010 (N_27010,N_19107,N_16224);
and U27011 (N_27011,N_18264,N_13522);
nor U27012 (N_27012,N_11025,N_14431);
nand U27013 (N_27013,N_14321,N_11352);
and U27014 (N_27014,N_17237,N_11613);
nor U27015 (N_27015,N_11258,N_16558);
nand U27016 (N_27016,N_13419,N_10203);
nand U27017 (N_27017,N_13848,N_17831);
or U27018 (N_27018,N_19681,N_14818);
xor U27019 (N_27019,N_16818,N_13535);
nand U27020 (N_27020,N_13679,N_16429);
or U27021 (N_27021,N_11578,N_10500);
and U27022 (N_27022,N_14234,N_14599);
nor U27023 (N_27023,N_16182,N_15599);
nor U27024 (N_27024,N_14186,N_16065);
nor U27025 (N_27025,N_19830,N_12475);
xnor U27026 (N_27026,N_18593,N_15176);
nand U27027 (N_27027,N_13444,N_16665);
nor U27028 (N_27028,N_14976,N_11467);
and U27029 (N_27029,N_19265,N_17232);
and U27030 (N_27030,N_11722,N_10683);
nor U27031 (N_27031,N_19405,N_16422);
and U27032 (N_27032,N_14260,N_16851);
or U27033 (N_27033,N_13186,N_18250);
nor U27034 (N_27034,N_14731,N_18547);
nor U27035 (N_27035,N_19833,N_14075);
and U27036 (N_27036,N_18443,N_11028);
or U27037 (N_27037,N_12983,N_17672);
and U27038 (N_27038,N_13053,N_12299);
and U27039 (N_27039,N_18221,N_14642);
nor U27040 (N_27040,N_14473,N_17098);
nor U27041 (N_27041,N_11286,N_19460);
or U27042 (N_27042,N_11348,N_18035);
and U27043 (N_27043,N_10410,N_12019);
nor U27044 (N_27044,N_18230,N_17921);
or U27045 (N_27045,N_19572,N_17280);
or U27046 (N_27046,N_14861,N_18037);
xor U27047 (N_27047,N_13020,N_12900);
and U27048 (N_27048,N_18312,N_11231);
or U27049 (N_27049,N_16832,N_10157);
nand U27050 (N_27050,N_19639,N_11852);
nor U27051 (N_27051,N_12917,N_11247);
nand U27052 (N_27052,N_19386,N_15638);
and U27053 (N_27053,N_11545,N_17214);
and U27054 (N_27054,N_15937,N_19330);
and U27055 (N_27055,N_10226,N_17878);
nand U27056 (N_27056,N_15246,N_11162);
nand U27057 (N_27057,N_17596,N_12233);
or U27058 (N_27058,N_19196,N_16982);
or U27059 (N_27059,N_17931,N_14193);
and U27060 (N_27060,N_17197,N_15535);
or U27061 (N_27061,N_17325,N_14743);
and U27062 (N_27062,N_10466,N_19046);
nand U27063 (N_27063,N_15289,N_12913);
or U27064 (N_27064,N_19193,N_17587);
nor U27065 (N_27065,N_12797,N_19130);
nand U27066 (N_27066,N_13885,N_13361);
nand U27067 (N_27067,N_10957,N_10731);
nor U27068 (N_27068,N_15156,N_14245);
nor U27069 (N_27069,N_16476,N_11198);
nor U27070 (N_27070,N_15824,N_17330);
nand U27071 (N_27071,N_11125,N_16224);
and U27072 (N_27072,N_14923,N_19110);
and U27073 (N_27073,N_11549,N_14309);
nor U27074 (N_27074,N_13985,N_11360);
nor U27075 (N_27075,N_16531,N_13820);
or U27076 (N_27076,N_18240,N_14110);
nor U27077 (N_27077,N_13099,N_16665);
xor U27078 (N_27078,N_12668,N_15844);
nand U27079 (N_27079,N_16817,N_15770);
nor U27080 (N_27080,N_11887,N_17668);
and U27081 (N_27081,N_13662,N_13340);
or U27082 (N_27082,N_10601,N_13769);
xor U27083 (N_27083,N_13941,N_14060);
nand U27084 (N_27084,N_12623,N_13765);
xnor U27085 (N_27085,N_12457,N_19731);
or U27086 (N_27086,N_17697,N_18639);
or U27087 (N_27087,N_16455,N_10853);
and U27088 (N_27088,N_12401,N_18332);
or U27089 (N_27089,N_14796,N_14355);
nand U27090 (N_27090,N_14174,N_15299);
nand U27091 (N_27091,N_17772,N_10189);
or U27092 (N_27092,N_11563,N_12863);
or U27093 (N_27093,N_17948,N_16961);
or U27094 (N_27094,N_14636,N_19552);
nand U27095 (N_27095,N_19812,N_15464);
and U27096 (N_27096,N_18910,N_11117);
and U27097 (N_27097,N_13207,N_12923);
nand U27098 (N_27098,N_18053,N_10978);
nor U27099 (N_27099,N_17290,N_14169);
nand U27100 (N_27100,N_17309,N_13513);
nand U27101 (N_27101,N_10698,N_12531);
and U27102 (N_27102,N_16410,N_10460);
nor U27103 (N_27103,N_14551,N_16081);
and U27104 (N_27104,N_12587,N_16456);
and U27105 (N_27105,N_11633,N_15586);
and U27106 (N_27106,N_10893,N_11246);
xnor U27107 (N_27107,N_15115,N_10131);
nand U27108 (N_27108,N_18537,N_14139);
nand U27109 (N_27109,N_15446,N_14389);
nand U27110 (N_27110,N_18499,N_10253);
or U27111 (N_27111,N_19759,N_14694);
or U27112 (N_27112,N_17564,N_17172);
nand U27113 (N_27113,N_11782,N_10401);
nor U27114 (N_27114,N_14371,N_10595);
nand U27115 (N_27115,N_19950,N_13992);
nor U27116 (N_27116,N_13890,N_12374);
or U27117 (N_27117,N_12098,N_16727);
nor U27118 (N_27118,N_12405,N_10590);
or U27119 (N_27119,N_15880,N_14170);
or U27120 (N_27120,N_12827,N_10457);
and U27121 (N_27121,N_18073,N_18224);
and U27122 (N_27122,N_16770,N_11986);
and U27123 (N_27123,N_15506,N_17349);
nand U27124 (N_27124,N_18936,N_12798);
nand U27125 (N_27125,N_17242,N_15566);
xnor U27126 (N_27126,N_14648,N_13619);
nand U27127 (N_27127,N_13504,N_13738);
or U27128 (N_27128,N_13051,N_15314);
nand U27129 (N_27129,N_19240,N_16608);
nand U27130 (N_27130,N_10443,N_16802);
nand U27131 (N_27131,N_15680,N_19386);
nor U27132 (N_27132,N_18411,N_19399);
and U27133 (N_27133,N_18755,N_13091);
nand U27134 (N_27134,N_15108,N_17408);
nand U27135 (N_27135,N_11654,N_18625);
nor U27136 (N_27136,N_15838,N_10488);
nand U27137 (N_27137,N_10429,N_11243);
nand U27138 (N_27138,N_17458,N_12933);
nand U27139 (N_27139,N_17907,N_13546);
and U27140 (N_27140,N_12332,N_19445);
and U27141 (N_27141,N_14456,N_14900);
or U27142 (N_27142,N_10987,N_16400);
or U27143 (N_27143,N_18355,N_19125);
nand U27144 (N_27144,N_19113,N_17298);
nor U27145 (N_27145,N_11493,N_19334);
or U27146 (N_27146,N_13287,N_19877);
nor U27147 (N_27147,N_16662,N_13267);
nor U27148 (N_27148,N_15523,N_19597);
nor U27149 (N_27149,N_18513,N_17711);
or U27150 (N_27150,N_17340,N_16026);
nor U27151 (N_27151,N_11097,N_16793);
or U27152 (N_27152,N_18872,N_16197);
xor U27153 (N_27153,N_10035,N_15549);
and U27154 (N_27154,N_18043,N_14634);
and U27155 (N_27155,N_19540,N_17428);
and U27156 (N_27156,N_10485,N_15101);
nor U27157 (N_27157,N_10719,N_13679);
or U27158 (N_27158,N_13929,N_16059);
and U27159 (N_27159,N_10736,N_16516);
nand U27160 (N_27160,N_12416,N_11428);
or U27161 (N_27161,N_10860,N_18391);
xor U27162 (N_27162,N_15713,N_15840);
nand U27163 (N_27163,N_11715,N_10604);
and U27164 (N_27164,N_19378,N_10003);
and U27165 (N_27165,N_19203,N_13936);
nor U27166 (N_27166,N_13709,N_17451);
nor U27167 (N_27167,N_13351,N_12804);
or U27168 (N_27168,N_13671,N_13434);
nor U27169 (N_27169,N_14695,N_18956);
nand U27170 (N_27170,N_13964,N_17318);
or U27171 (N_27171,N_13976,N_11079);
nand U27172 (N_27172,N_11839,N_15043);
nor U27173 (N_27173,N_10158,N_17324);
and U27174 (N_27174,N_18852,N_18041);
or U27175 (N_27175,N_16171,N_17562);
or U27176 (N_27176,N_14347,N_12942);
nor U27177 (N_27177,N_15564,N_14299);
and U27178 (N_27178,N_13076,N_15033);
or U27179 (N_27179,N_10347,N_14092);
or U27180 (N_27180,N_12571,N_11218);
nor U27181 (N_27181,N_12355,N_11063);
or U27182 (N_27182,N_17619,N_15305);
or U27183 (N_27183,N_14059,N_18582);
nand U27184 (N_27184,N_11544,N_10098);
nand U27185 (N_27185,N_14984,N_19002);
nand U27186 (N_27186,N_16801,N_14766);
and U27187 (N_27187,N_12467,N_19050);
nor U27188 (N_27188,N_14645,N_13099);
nor U27189 (N_27189,N_16698,N_18176);
nand U27190 (N_27190,N_10132,N_12681);
or U27191 (N_27191,N_17180,N_12211);
and U27192 (N_27192,N_12746,N_15838);
or U27193 (N_27193,N_19004,N_16124);
nand U27194 (N_27194,N_19313,N_14276);
xor U27195 (N_27195,N_14719,N_14135);
nand U27196 (N_27196,N_12695,N_17559);
or U27197 (N_27197,N_18722,N_13286);
and U27198 (N_27198,N_15107,N_11982);
nor U27199 (N_27199,N_15418,N_19934);
nand U27200 (N_27200,N_18550,N_13591);
nor U27201 (N_27201,N_18942,N_12015);
nor U27202 (N_27202,N_16376,N_19260);
and U27203 (N_27203,N_16168,N_12615);
nand U27204 (N_27204,N_15219,N_19807);
and U27205 (N_27205,N_16840,N_17791);
nand U27206 (N_27206,N_15463,N_11601);
nor U27207 (N_27207,N_16852,N_17074);
and U27208 (N_27208,N_13212,N_16743);
nor U27209 (N_27209,N_18700,N_16601);
xnor U27210 (N_27210,N_14433,N_10123);
or U27211 (N_27211,N_19683,N_15833);
and U27212 (N_27212,N_10295,N_18113);
xnor U27213 (N_27213,N_14392,N_19205);
nor U27214 (N_27214,N_16275,N_15291);
nor U27215 (N_27215,N_17285,N_14362);
nor U27216 (N_27216,N_18859,N_13606);
and U27217 (N_27217,N_19829,N_13545);
nand U27218 (N_27218,N_10820,N_11965);
nand U27219 (N_27219,N_12932,N_15493);
nand U27220 (N_27220,N_19607,N_12857);
nor U27221 (N_27221,N_11511,N_13716);
nand U27222 (N_27222,N_19552,N_13679);
or U27223 (N_27223,N_10214,N_11064);
or U27224 (N_27224,N_10016,N_12723);
or U27225 (N_27225,N_12501,N_15674);
nand U27226 (N_27226,N_18497,N_13355);
nor U27227 (N_27227,N_11882,N_12326);
nand U27228 (N_27228,N_13206,N_10852);
or U27229 (N_27229,N_18080,N_12144);
and U27230 (N_27230,N_14938,N_16825);
or U27231 (N_27231,N_18712,N_14356);
nor U27232 (N_27232,N_13234,N_16447);
or U27233 (N_27233,N_10044,N_10806);
or U27234 (N_27234,N_19407,N_10190);
and U27235 (N_27235,N_16837,N_19264);
nand U27236 (N_27236,N_13080,N_11062);
nand U27237 (N_27237,N_17243,N_14094);
nand U27238 (N_27238,N_14065,N_18956);
and U27239 (N_27239,N_15459,N_18191);
and U27240 (N_27240,N_16451,N_19328);
nand U27241 (N_27241,N_14521,N_12395);
nor U27242 (N_27242,N_12900,N_14070);
and U27243 (N_27243,N_15216,N_16930);
nand U27244 (N_27244,N_19650,N_13646);
nor U27245 (N_27245,N_15052,N_16879);
nor U27246 (N_27246,N_18952,N_12143);
nor U27247 (N_27247,N_13474,N_14122);
or U27248 (N_27248,N_17835,N_12684);
or U27249 (N_27249,N_18908,N_13553);
nor U27250 (N_27250,N_16150,N_16549);
xor U27251 (N_27251,N_17260,N_15234);
or U27252 (N_27252,N_15146,N_10673);
nor U27253 (N_27253,N_13105,N_19034);
and U27254 (N_27254,N_10607,N_18817);
and U27255 (N_27255,N_15485,N_16173);
or U27256 (N_27256,N_19540,N_10257);
nand U27257 (N_27257,N_10136,N_19759);
nand U27258 (N_27258,N_13967,N_19885);
nand U27259 (N_27259,N_15018,N_14501);
and U27260 (N_27260,N_13579,N_19598);
nor U27261 (N_27261,N_12607,N_17762);
and U27262 (N_27262,N_11418,N_12697);
nor U27263 (N_27263,N_18928,N_12289);
and U27264 (N_27264,N_11422,N_17919);
nand U27265 (N_27265,N_19779,N_10510);
and U27266 (N_27266,N_16073,N_15372);
and U27267 (N_27267,N_19467,N_19635);
nor U27268 (N_27268,N_13129,N_17883);
xnor U27269 (N_27269,N_19973,N_10399);
and U27270 (N_27270,N_19543,N_17147);
or U27271 (N_27271,N_12087,N_16780);
or U27272 (N_27272,N_15721,N_12771);
and U27273 (N_27273,N_11554,N_15080);
or U27274 (N_27274,N_12416,N_16512);
or U27275 (N_27275,N_16555,N_13616);
or U27276 (N_27276,N_18630,N_17326);
or U27277 (N_27277,N_12635,N_15602);
or U27278 (N_27278,N_13056,N_14738);
and U27279 (N_27279,N_19581,N_15840);
nor U27280 (N_27280,N_16084,N_18933);
and U27281 (N_27281,N_14409,N_18067);
nor U27282 (N_27282,N_11963,N_18217);
xnor U27283 (N_27283,N_12201,N_12003);
xor U27284 (N_27284,N_17711,N_15221);
xor U27285 (N_27285,N_13569,N_16254);
xor U27286 (N_27286,N_13503,N_10604);
or U27287 (N_27287,N_12680,N_15925);
or U27288 (N_27288,N_10705,N_12005);
nand U27289 (N_27289,N_18420,N_16071);
and U27290 (N_27290,N_12460,N_11466);
nor U27291 (N_27291,N_14695,N_17164);
or U27292 (N_27292,N_13920,N_16496);
and U27293 (N_27293,N_12226,N_19810);
or U27294 (N_27294,N_13630,N_13889);
nor U27295 (N_27295,N_11519,N_18620);
nor U27296 (N_27296,N_17063,N_17394);
and U27297 (N_27297,N_12132,N_17986);
nand U27298 (N_27298,N_12584,N_11483);
nand U27299 (N_27299,N_19178,N_17616);
nand U27300 (N_27300,N_14874,N_19110);
or U27301 (N_27301,N_11341,N_10472);
or U27302 (N_27302,N_11764,N_12503);
nor U27303 (N_27303,N_16787,N_12473);
or U27304 (N_27304,N_15967,N_14414);
or U27305 (N_27305,N_18486,N_15721);
or U27306 (N_27306,N_18604,N_11213);
nor U27307 (N_27307,N_10467,N_10375);
and U27308 (N_27308,N_17673,N_16042);
and U27309 (N_27309,N_19088,N_12677);
xnor U27310 (N_27310,N_18253,N_13181);
and U27311 (N_27311,N_17512,N_15492);
or U27312 (N_27312,N_15752,N_14934);
nor U27313 (N_27313,N_12842,N_13186);
or U27314 (N_27314,N_15223,N_13911);
nor U27315 (N_27315,N_18345,N_16942);
nand U27316 (N_27316,N_10675,N_10689);
nand U27317 (N_27317,N_14621,N_17539);
nand U27318 (N_27318,N_15883,N_16150);
or U27319 (N_27319,N_18400,N_13536);
and U27320 (N_27320,N_13796,N_17235);
xnor U27321 (N_27321,N_17799,N_18833);
or U27322 (N_27322,N_11415,N_17250);
nand U27323 (N_27323,N_15581,N_13932);
or U27324 (N_27324,N_15857,N_11739);
xnor U27325 (N_27325,N_13400,N_13731);
and U27326 (N_27326,N_19636,N_16411);
nand U27327 (N_27327,N_16352,N_14100);
nor U27328 (N_27328,N_11404,N_12225);
nand U27329 (N_27329,N_17679,N_19160);
or U27330 (N_27330,N_19224,N_18563);
nand U27331 (N_27331,N_17994,N_18239);
nor U27332 (N_27332,N_12551,N_11272);
nor U27333 (N_27333,N_12744,N_16534);
nor U27334 (N_27334,N_17749,N_10907);
nand U27335 (N_27335,N_19807,N_18891);
nor U27336 (N_27336,N_13989,N_18646);
or U27337 (N_27337,N_14974,N_16223);
nand U27338 (N_27338,N_12286,N_10609);
and U27339 (N_27339,N_11487,N_16490);
nor U27340 (N_27340,N_13860,N_15601);
nand U27341 (N_27341,N_15988,N_12598);
nor U27342 (N_27342,N_13628,N_10120);
nand U27343 (N_27343,N_19485,N_11106);
and U27344 (N_27344,N_12296,N_12137);
or U27345 (N_27345,N_13649,N_17048);
nand U27346 (N_27346,N_15363,N_19686);
and U27347 (N_27347,N_18861,N_13609);
nand U27348 (N_27348,N_13608,N_17508);
nand U27349 (N_27349,N_19762,N_15345);
and U27350 (N_27350,N_17695,N_11971);
and U27351 (N_27351,N_18287,N_17576);
and U27352 (N_27352,N_12722,N_12956);
and U27353 (N_27353,N_19479,N_16197);
nor U27354 (N_27354,N_14514,N_15834);
nand U27355 (N_27355,N_16851,N_13187);
and U27356 (N_27356,N_10851,N_13998);
nand U27357 (N_27357,N_12467,N_13687);
nor U27358 (N_27358,N_10486,N_15824);
or U27359 (N_27359,N_16017,N_10176);
and U27360 (N_27360,N_15718,N_12693);
nor U27361 (N_27361,N_19117,N_14422);
and U27362 (N_27362,N_12164,N_18558);
nand U27363 (N_27363,N_13380,N_17472);
xor U27364 (N_27364,N_19238,N_12810);
or U27365 (N_27365,N_19124,N_10959);
nor U27366 (N_27366,N_15986,N_10897);
nor U27367 (N_27367,N_18923,N_17394);
xnor U27368 (N_27368,N_16862,N_15872);
nor U27369 (N_27369,N_10330,N_13272);
and U27370 (N_27370,N_11018,N_19592);
nand U27371 (N_27371,N_13643,N_17095);
nand U27372 (N_27372,N_14965,N_15012);
xor U27373 (N_27373,N_18779,N_15197);
and U27374 (N_27374,N_18597,N_19188);
and U27375 (N_27375,N_19060,N_17973);
xnor U27376 (N_27376,N_12951,N_15470);
nor U27377 (N_27377,N_11701,N_18407);
nor U27378 (N_27378,N_10674,N_10999);
or U27379 (N_27379,N_11048,N_16147);
nor U27380 (N_27380,N_17385,N_17749);
and U27381 (N_27381,N_17569,N_15771);
and U27382 (N_27382,N_19528,N_13980);
xnor U27383 (N_27383,N_18728,N_12592);
or U27384 (N_27384,N_19149,N_14450);
nand U27385 (N_27385,N_16656,N_12839);
and U27386 (N_27386,N_12336,N_13452);
xnor U27387 (N_27387,N_19231,N_10062);
nand U27388 (N_27388,N_16984,N_12841);
nand U27389 (N_27389,N_14963,N_15784);
nor U27390 (N_27390,N_15903,N_15055);
and U27391 (N_27391,N_13551,N_14031);
nor U27392 (N_27392,N_19766,N_11747);
nand U27393 (N_27393,N_12580,N_16438);
and U27394 (N_27394,N_15278,N_17578);
and U27395 (N_27395,N_12736,N_16962);
and U27396 (N_27396,N_12424,N_18707);
and U27397 (N_27397,N_14411,N_13941);
xor U27398 (N_27398,N_18409,N_17967);
nand U27399 (N_27399,N_17703,N_14295);
and U27400 (N_27400,N_15171,N_15593);
nor U27401 (N_27401,N_15393,N_12469);
and U27402 (N_27402,N_16307,N_10674);
nor U27403 (N_27403,N_17737,N_12118);
nand U27404 (N_27404,N_15029,N_18742);
nor U27405 (N_27405,N_15494,N_19414);
xor U27406 (N_27406,N_10852,N_14216);
and U27407 (N_27407,N_11188,N_17025);
and U27408 (N_27408,N_19829,N_12105);
nor U27409 (N_27409,N_18690,N_14317);
and U27410 (N_27410,N_12251,N_12416);
nand U27411 (N_27411,N_10076,N_19888);
nor U27412 (N_27412,N_18817,N_13351);
or U27413 (N_27413,N_14078,N_16712);
nor U27414 (N_27414,N_17275,N_14639);
nor U27415 (N_27415,N_14053,N_11438);
or U27416 (N_27416,N_19861,N_12790);
or U27417 (N_27417,N_10507,N_17838);
or U27418 (N_27418,N_10249,N_11758);
and U27419 (N_27419,N_11061,N_19060);
or U27420 (N_27420,N_18012,N_18247);
or U27421 (N_27421,N_17727,N_10862);
nand U27422 (N_27422,N_19050,N_13041);
nor U27423 (N_27423,N_18128,N_17793);
and U27424 (N_27424,N_16853,N_18052);
and U27425 (N_27425,N_18282,N_18382);
nor U27426 (N_27426,N_14566,N_18084);
nor U27427 (N_27427,N_18184,N_13036);
xor U27428 (N_27428,N_14535,N_12447);
xnor U27429 (N_27429,N_16425,N_10921);
nand U27430 (N_27430,N_13751,N_19566);
xor U27431 (N_27431,N_13116,N_14555);
or U27432 (N_27432,N_11756,N_13843);
xnor U27433 (N_27433,N_14126,N_19476);
or U27434 (N_27434,N_12187,N_15752);
or U27435 (N_27435,N_12934,N_11043);
nand U27436 (N_27436,N_17500,N_11013);
and U27437 (N_27437,N_10517,N_19242);
or U27438 (N_27438,N_17561,N_17850);
and U27439 (N_27439,N_10154,N_10877);
nand U27440 (N_27440,N_15761,N_19569);
nor U27441 (N_27441,N_16099,N_10004);
or U27442 (N_27442,N_13402,N_12847);
or U27443 (N_27443,N_11538,N_12606);
and U27444 (N_27444,N_17177,N_10452);
and U27445 (N_27445,N_13374,N_10735);
and U27446 (N_27446,N_14256,N_10635);
or U27447 (N_27447,N_14778,N_15269);
nor U27448 (N_27448,N_10421,N_16113);
and U27449 (N_27449,N_10183,N_10677);
nand U27450 (N_27450,N_14024,N_12219);
or U27451 (N_27451,N_17802,N_16442);
nand U27452 (N_27452,N_16406,N_17240);
nand U27453 (N_27453,N_11671,N_16172);
nand U27454 (N_27454,N_15443,N_11440);
xor U27455 (N_27455,N_11652,N_12785);
or U27456 (N_27456,N_17578,N_12235);
nor U27457 (N_27457,N_14873,N_15190);
nand U27458 (N_27458,N_12524,N_13775);
nand U27459 (N_27459,N_11487,N_13040);
and U27460 (N_27460,N_11323,N_10741);
nor U27461 (N_27461,N_16356,N_12676);
and U27462 (N_27462,N_18347,N_19796);
nor U27463 (N_27463,N_11530,N_17429);
and U27464 (N_27464,N_14540,N_17414);
and U27465 (N_27465,N_17077,N_11774);
nor U27466 (N_27466,N_17384,N_13673);
nor U27467 (N_27467,N_10974,N_14352);
nor U27468 (N_27468,N_10687,N_12413);
xor U27469 (N_27469,N_19567,N_13220);
nand U27470 (N_27470,N_17591,N_11725);
and U27471 (N_27471,N_19902,N_16331);
and U27472 (N_27472,N_18611,N_10115);
and U27473 (N_27473,N_17455,N_19968);
and U27474 (N_27474,N_10272,N_13936);
nand U27475 (N_27475,N_13730,N_14579);
nand U27476 (N_27476,N_11373,N_10774);
nand U27477 (N_27477,N_19631,N_12821);
nand U27478 (N_27478,N_15515,N_19887);
nand U27479 (N_27479,N_12203,N_15118);
nor U27480 (N_27480,N_16006,N_11662);
nor U27481 (N_27481,N_18317,N_12623);
and U27482 (N_27482,N_16194,N_14240);
nor U27483 (N_27483,N_14831,N_13003);
nand U27484 (N_27484,N_16287,N_18186);
nor U27485 (N_27485,N_13117,N_10842);
nor U27486 (N_27486,N_15432,N_16886);
nand U27487 (N_27487,N_19912,N_10992);
or U27488 (N_27488,N_18713,N_12732);
nor U27489 (N_27489,N_15828,N_16221);
nand U27490 (N_27490,N_12487,N_11390);
and U27491 (N_27491,N_16891,N_16460);
and U27492 (N_27492,N_18169,N_11139);
or U27493 (N_27493,N_17249,N_11500);
and U27494 (N_27494,N_19425,N_18023);
xor U27495 (N_27495,N_18847,N_10223);
xor U27496 (N_27496,N_14345,N_11396);
nor U27497 (N_27497,N_14860,N_18630);
and U27498 (N_27498,N_11404,N_19400);
nand U27499 (N_27499,N_19151,N_16335);
nand U27500 (N_27500,N_11541,N_18029);
and U27501 (N_27501,N_11263,N_17996);
nor U27502 (N_27502,N_15158,N_15627);
nand U27503 (N_27503,N_15418,N_12348);
and U27504 (N_27504,N_12588,N_15345);
and U27505 (N_27505,N_10926,N_10950);
and U27506 (N_27506,N_10986,N_16753);
and U27507 (N_27507,N_15990,N_10535);
or U27508 (N_27508,N_17440,N_17293);
nand U27509 (N_27509,N_15915,N_16378);
or U27510 (N_27510,N_15394,N_15503);
and U27511 (N_27511,N_16193,N_16639);
or U27512 (N_27512,N_19601,N_17101);
and U27513 (N_27513,N_12050,N_14840);
or U27514 (N_27514,N_19787,N_16294);
and U27515 (N_27515,N_10285,N_17029);
nor U27516 (N_27516,N_14287,N_14639);
or U27517 (N_27517,N_15052,N_11044);
and U27518 (N_27518,N_11370,N_16765);
or U27519 (N_27519,N_11517,N_12801);
or U27520 (N_27520,N_18016,N_16488);
nand U27521 (N_27521,N_10703,N_12551);
nor U27522 (N_27522,N_15317,N_15188);
xor U27523 (N_27523,N_13812,N_13473);
nor U27524 (N_27524,N_12051,N_13621);
and U27525 (N_27525,N_17144,N_18464);
nor U27526 (N_27526,N_13907,N_13858);
nor U27527 (N_27527,N_12999,N_18106);
nor U27528 (N_27528,N_12028,N_14141);
nor U27529 (N_27529,N_17833,N_10225);
xor U27530 (N_27530,N_11002,N_15010);
nor U27531 (N_27531,N_15819,N_11847);
or U27532 (N_27532,N_11263,N_13127);
nand U27533 (N_27533,N_17315,N_15397);
nand U27534 (N_27534,N_13660,N_13658);
or U27535 (N_27535,N_11120,N_12147);
nor U27536 (N_27536,N_10743,N_16650);
nor U27537 (N_27537,N_15041,N_16939);
or U27538 (N_27538,N_18654,N_16502);
and U27539 (N_27539,N_16255,N_11053);
nand U27540 (N_27540,N_12420,N_12755);
xnor U27541 (N_27541,N_14791,N_18686);
nor U27542 (N_27542,N_13276,N_18219);
and U27543 (N_27543,N_17938,N_14035);
nor U27544 (N_27544,N_16389,N_16846);
nand U27545 (N_27545,N_18481,N_13187);
or U27546 (N_27546,N_11115,N_13651);
nor U27547 (N_27547,N_15757,N_18639);
or U27548 (N_27548,N_18907,N_16372);
nand U27549 (N_27549,N_12369,N_10510);
and U27550 (N_27550,N_10628,N_17612);
or U27551 (N_27551,N_12425,N_13204);
or U27552 (N_27552,N_14228,N_17756);
and U27553 (N_27553,N_12327,N_13907);
and U27554 (N_27554,N_19343,N_18270);
nor U27555 (N_27555,N_10113,N_14311);
nor U27556 (N_27556,N_18632,N_17426);
and U27557 (N_27557,N_15540,N_17226);
nor U27558 (N_27558,N_10178,N_11204);
nor U27559 (N_27559,N_15919,N_10898);
and U27560 (N_27560,N_11747,N_16177);
nand U27561 (N_27561,N_19038,N_16745);
nand U27562 (N_27562,N_17195,N_15517);
and U27563 (N_27563,N_19321,N_13218);
or U27564 (N_27564,N_18771,N_18484);
nor U27565 (N_27565,N_10100,N_19417);
nor U27566 (N_27566,N_10070,N_10983);
or U27567 (N_27567,N_15916,N_14746);
and U27568 (N_27568,N_15873,N_12020);
nor U27569 (N_27569,N_18967,N_17330);
nor U27570 (N_27570,N_11323,N_15611);
or U27571 (N_27571,N_19380,N_19919);
or U27572 (N_27572,N_19201,N_17751);
or U27573 (N_27573,N_17259,N_18037);
nor U27574 (N_27574,N_14521,N_19507);
xnor U27575 (N_27575,N_15736,N_15264);
nand U27576 (N_27576,N_17528,N_17672);
nor U27577 (N_27577,N_13985,N_12348);
and U27578 (N_27578,N_17661,N_11591);
and U27579 (N_27579,N_10511,N_10633);
nand U27580 (N_27580,N_18649,N_18727);
nor U27581 (N_27581,N_12566,N_17288);
and U27582 (N_27582,N_12488,N_14934);
or U27583 (N_27583,N_14262,N_14707);
or U27584 (N_27584,N_17137,N_11114);
and U27585 (N_27585,N_10312,N_12341);
nor U27586 (N_27586,N_18641,N_10042);
nor U27587 (N_27587,N_18616,N_15629);
and U27588 (N_27588,N_11497,N_11955);
and U27589 (N_27589,N_18027,N_18035);
nor U27590 (N_27590,N_14335,N_15888);
or U27591 (N_27591,N_16130,N_11388);
nor U27592 (N_27592,N_18447,N_19076);
nand U27593 (N_27593,N_18336,N_12488);
nor U27594 (N_27594,N_12872,N_19142);
or U27595 (N_27595,N_18042,N_18210);
nand U27596 (N_27596,N_19041,N_19890);
nor U27597 (N_27597,N_11580,N_19579);
and U27598 (N_27598,N_17282,N_15454);
or U27599 (N_27599,N_17828,N_17784);
xnor U27600 (N_27600,N_15468,N_16749);
nor U27601 (N_27601,N_10571,N_13033);
nor U27602 (N_27602,N_19886,N_18451);
nor U27603 (N_27603,N_13283,N_11230);
nand U27604 (N_27604,N_19546,N_17777);
nand U27605 (N_27605,N_19092,N_18675);
nor U27606 (N_27606,N_14886,N_15711);
or U27607 (N_27607,N_17094,N_19491);
or U27608 (N_27608,N_18970,N_19460);
nor U27609 (N_27609,N_19598,N_11963);
and U27610 (N_27610,N_17520,N_13531);
nor U27611 (N_27611,N_15287,N_16474);
xor U27612 (N_27612,N_15422,N_13108);
or U27613 (N_27613,N_14413,N_12234);
nand U27614 (N_27614,N_12137,N_13728);
nor U27615 (N_27615,N_13787,N_10836);
nand U27616 (N_27616,N_15047,N_12329);
nor U27617 (N_27617,N_16713,N_14075);
nand U27618 (N_27618,N_19316,N_15799);
nor U27619 (N_27619,N_19038,N_13255);
and U27620 (N_27620,N_19433,N_18503);
and U27621 (N_27621,N_15378,N_13266);
and U27622 (N_27622,N_12336,N_14153);
nor U27623 (N_27623,N_13640,N_16835);
or U27624 (N_27624,N_13632,N_17828);
or U27625 (N_27625,N_18132,N_18001);
nor U27626 (N_27626,N_17282,N_15735);
or U27627 (N_27627,N_11053,N_19587);
nor U27628 (N_27628,N_18956,N_17964);
or U27629 (N_27629,N_18372,N_13871);
nor U27630 (N_27630,N_16943,N_10244);
nand U27631 (N_27631,N_14675,N_10608);
or U27632 (N_27632,N_16695,N_16091);
nand U27633 (N_27633,N_14344,N_18890);
nand U27634 (N_27634,N_13026,N_10934);
nor U27635 (N_27635,N_19191,N_14843);
nand U27636 (N_27636,N_16229,N_19046);
nand U27637 (N_27637,N_16406,N_16061);
nor U27638 (N_27638,N_14351,N_12040);
and U27639 (N_27639,N_14854,N_10311);
nand U27640 (N_27640,N_19026,N_18585);
nand U27641 (N_27641,N_15703,N_12102);
nor U27642 (N_27642,N_16428,N_16990);
nor U27643 (N_27643,N_12075,N_14003);
nor U27644 (N_27644,N_19491,N_11448);
and U27645 (N_27645,N_16255,N_18793);
and U27646 (N_27646,N_16523,N_12357);
or U27647 (N_27647,N_10914,N_15066);
nor U27648 (N_27648,N_13603,N_19528);
nor U27649 (N_27649,N_18560,N_18581);
nor U27650 (N_27650,N_15031,N_17934);
nand U27651 (N_27651,N_16366,N_18724);
or U27652 (N_27652,N_12650,N_16152);
or U27653 (N_27653,N_11446,N_10316);
xnor U27654 (N_27654,N_19030,N_19222);
or U27655 (N_27655,N_16864,N_14259);
and U27656 (N_27656,N_15066,N_11127);
nor U27657 (N_27657,N_11017,N_19878);
nor U27658 (N_27658,N_10428,N_16445);
nand U27659 (N_27659,N_12537,N_17583);
nand U27660 (N_27660,N_14531,N_12143);
and U27661 (N_27661,N_12679,N_14497);
or U27662 (N_27662,N_18664,N_13436);
nor U27663 (N_27663,N_17192,N_10352);
or U27664 (N_27664,N_19169,N_16977);
xnor U27665 (N_27665,N_10398,N_13208);
and U27666 (N_27666,N_12795,N_10711);
nand U27667 (N_27667,N_10339,N_13050);
nand U27668 (N_27668,N_14768,N_15464);
xor U27669 (N_27669,N_15650,N_19078);
or U27670 (N_27670,N_12637,N_19794);
or U27671 (N_27671,N_16320,N_18334);
nor U27672 (N_27672,N_13321,N_14638);
nand U27673 (N_27673,N_16723,N_11263);
or U27674 (N_27674,N_17669,N_10026);
nand U27675 (N_27675,N_11958,N_14792);
nand U27676 (N_27676,N_12317,N_14169);
and U27677 (N_27677,N_12898,N_15428);
xor U27678 (N_27678,N_15118,N_10959);
nor U27679 (N_27679,N_18986,N_12765);
or U27680 (N_27680,N_10480,N_10301);
and U27681 (N_27681,N_18472,N_13772);
nor U27682 (N_27682,N_18612,N_12802);
nand U27683 (N_27683,N_16692,N_13572);
xor U27684 (N_27684,N_18463,N_11720);
nor U27685 (N_27685,N_18242,N_17266);
nor U27686 (N_27686,N_14978,N_15124);
nor U27687 (N_27687,N_14809,N_19814);
xnor U27688 (N_27688,N_16825,N_11174);
or U27689 (N_27689,N_19052,N_14377);
or U27690 (N_27690,N_17341,N_11649);
or U27691 (N_27691,N_13172,N_11322);
and U27692 (N_27692,N_19999,N_15575);
nand U27693 (N_27693,N_16449,N_18094);
nand U27694 (N_27694,N_17210,N_18207);
nor U27695 (N_27695,N_10793,N_10243);
or U27696 (N_27696,N_11623,N_10101);
nand U27697 (N_27697,N_11587,N_19201);
nor U27698 (N_27698,N_18708,N_12516);
or U27699 (N_27699,N_10494,N_10228);
nor U27700 (N_27700,N_10978,N_15896);
or U27701 (N_27701,N_13997,N_13014);
and U27702 (N_27702,N_16720,N_16115);
or U27703 (N_27703,N_10272,N_12369);
nor U27704 (N_27704,N_10424,N_15864);
nand U27705 (N_27705,N_17527,N_16908);
or U27706 (N_27706,N_13655,N_14148);
or U27707 (N_27707,N_16787,N_16440);
xnor U27708 (N_27708,N_17694,N_18984);
or U27709 (N_27709,N_13570,N_10789);
and U27710 (N_27710,N_13345,N_18995);
nor U27711 (N_27711,N_19473,N_19092);
xnor U27712 (N_27712,N_13254,N_19577);
or U27713 (N_27713,N_17562,N_15802);
nor U27714 (N_27714,N_18038,N_19146);
and U27715 (N_27715,N_14789,N_12618);
nand U27716 (N_27716,N_19390,N_13936);
nand U27717 (N_27717,N_16070,N_15656);
and U27718 (N_27718,N_18395,N_19913);
nand U27719 (N_27719,N_18443,N_10927);
nor U27720 (N_27720,N_11372,N_13400);
nand U27721 (N_27721,N_19257,N_10962);
or U27722 (N_27722,N_11379,N_15893);
nor U27723 (N_27723,N_16065,N_11597);
or U27724 (N_27724,N_13177,N_17420);
nand U27725 (N_27725,N_14728,N_18379);
nand U27726 (N_27726,N_11862,N_17521);
nor U27727 (N_27727,N_12615,N_17972);
or U27728 (N_27728,N_16529,N_14549);
and U27729 (N_27729,N_14390,N_14288);
and U27730 (N_27730,N_14870,N_11529);
nand U27731 (N_27731,N_17131,N_10456);
and U27732 (N_27732,N_10813,N_17076);
nor U27733 (N_27733,N_11384,N_19247);
nand U27734 (N_27734,N_19061,N_19675);
nand U27735 (N_27735,N_12730,N_10140);
and U27736 (N_27736,N_12808,N_13400);
nand U27737 (N_27737,N_10979,N_16842);
or U27738 (N_27738,N_10977,N_11417);
or U27739 (N_27739,N_10354,N_18760);
or U27740 (N_27740,N_13650,N_13542);
xnor U27741 (N_27741,N_16713,N_12616);
nand U27742 (N_27742,N_14133,N_17181);
nor U27743 (N_27743,N_11653,N_18747);
nor U27744 (N_27744,N_18926,N_11488);
nand U27745 (N_27745,N_10678,N_12775);
and U27746 (N_27746,N_10596,N_12391);
and U27747 (N_27747,N_19117,N_11392);
or U27748 (N_27748,N_13739,N_19302);
nor U27749 (N_27749,N_19761,N_19798);
nand U27750 (N_27750,N_18934,N_13285);
nand U27751 (N_27751,N_12965,N_17112);
and U27752 (N_27752,N_16540,N_19519);
nand U27753 (N_27753,N_15532,N_14152);
and U27754 (N_27754,N_13261,N_15499);
and U27755 (N_27755,N_12684,N_11359);
and U27756 (N_27756,N_17964,N_18553);
nor U27757 (N_27757,N_15151,N_15600);
nor U27758 (N_27758,N_19495,N_14753);
or U27759 (N_27759,N_19342,N_13699);
and U27760 (N_27760,N_16413,N_15255);
nor U27761 (N_27761,N_12946,N_19865);
or U27762 (N_27762,N_13010,N_17481);
nor U27763 (N_27763,N_11900,N_18208);
and U27764 (N_27764,N_14348,N_13461);
and U27765 (N_27765,N_11229,N_19343);
nor U27766 (N_27766,N_15925,N_10902);
and U27767 (N_27767,N_11382,N_14862);
xor U27768 (N_27768,N_12039,N_10597);
nor U27769 (N_27769,N_17393,N_18871);
and U27770 (N_27770,N_11054,N_11145);
nand U27771 (N_27771,N_13488,N_19389);
nand U27772 (N_27772,N_18553,N_10909);
xnor U27773 (N_27773,N_14944,N_19609);
or U27774 (N_27774,N_15477,N_10640);
and U27775 (N_27775,N_15415,N_19518);
xor U27776 (N_27776,N_17725,N_10981);
nand U27777 (N_27777,N_13108,N_15067);
xnor U27778 (N_27778,N_10764,N_18665);
and U27779 (N_27779,N_10543,N_15773);
or U27780 (N_27780,N_11286,N_13716);
nand U27781 (N_27781,N_10651,N_14104);
nor U27782 (N_27782,N_14911,N_16769);
nand U27783 (N_27783,N_19419,N_17376);
or U27784 (N_27784,N_10166,N_10891);
or U27785 (N_27785,N_15989,N_14000);
nand U27786 (N_27786,N_18742,N_18987);
nor U27787 (N_27787,N_14020,N_16373);
nor U27788 (N_27788,N_11000,N_10637);
xor U27789 (N_27789,N_16182,N_13656);
nand U27790 (N_27790,N_12639,N_17039);
or U27791 (N_27791,N_16520,N_10344);
nor U27792 (N_27792,N_17871,N_16692);
nor U27793 (N_27793,N_12609,N_18812);
or U27794 (N_27794,N_10123,N_10462);
and U27795 (N_27795,N_14323,N_16807);
or U27796 (N_27796,N_19738,N_12190);
nand U27797 (N_27797,N_13218,N_17940);
nor U27798 (N_27798,N_15379,N_17065);
nand U27799 (N_27799,N_14492,N_18283);
or U27800 (N_27800,N_13957,N_19490);
and U27801 (N_27801,N_11911,N_10959);
nor U27802 (N_27802,N_19621,N_19361);
nand U27803 (N_27803,N_10270,N_18486);
nor U27804 (N_27804,N_11082,N_16716);
and U27805 (N_27805,N_10929,N_17181);
or U27806 (N_27806,N_12167,N_17987);
or U27807 (N_27807,N_10861,N_17867);
nor U27808 (N_27808,N_17341,N_18618);
nand U27809 (N_27809,N_14064,N_17116);
nor U27810 (N_27810,N_13495,N_16422);
and U27811 (N_27811,N_17292,N_10413);
nor U27812 (N_27812,N_13388,N_13398);
nor U27813 (N_27813,N_15322,N_17590);
or U27814 (N_27814,N_18313,N_18925);
nand U27815 (N_27815,N_12125,N_19394);
nand U27816 (N_27816,N_11355,N_12771);
nand U27817 (N_27817,N_14255,N_18046);
nor U27818 (N_27818,N_16828,N_11774);
nor U27819 (N_27819,N_12685,N_14612);
or U27820 (N_27820,N_12384,N_11645);
nand U27821 (N_27821,N_11903,N_13973);
nor U27822 (N_27822,N_13921,N_18216);
or U27823 (N_27823,N_13210,N_19259);
nor U27824 (N_27824,N_10552,N_17141);
nand U27825 (N_27825,N_16539,N_15461);
nand U27826 (N_27826,N_14434,N_10253);
nor U27827 (N_27827,N_15715,N_11982);
or U27828 (N_27828,N_14015,N_17284);
nand U27829 (N_27829,N_14915,N_18735);
and U27830 (N_27830,N_16552,N_18272);
nor U27831 (N_27831,N_12367,N_19359);
nor U27832 (N_27832,N_16421,N_13619);
or U27833 (N_27833,N_17427,N_18238);
and U27834 (N_27834,N_16930,N_16147);
nand U27835 (N_27835,N_12946,N_11891);
xnor U27836 (N_27836,N_19770,N_17573);
and U27837 (N_27837,N_10953,N_13341);
or U27838 (N_27838,N_15008,N_19510);
xnor U27839 (N_27839,N_11072,N_18980);
nor U27840 (N_27840,N_19230,N_14057);
and U27841 (N_27841,N_10083,N_13262);
nand U27842 (N_27842,N_18698,N_19400);
xnor U27843 (N_27843,N_18361,N_11643);
nand U27844 (N_27844,N_18423,N_15742);
xnor U27845 (N_27845,N_11614,N_10657);
nand U27846 (N_27846,N_19592,N_11098);
or U27847 (N_27847,N_19728,N_14084);
xnor U27848 (N_27848,N_10493,N_10786);
nand U27849 (N_27849,N_12666,N_19105);
nand U27850 (N_27850,N_19307,N_14924);
or U27851 (N_27851,N_14402,N_17478);
nand U27852 (N_27852,N_13428,N_10363);
and U27853 (N_27853,N_14343,N_17545);
and U27854 (N_27854,N_14870,N_16479);
or U27855 (N_27855,N_19745,N_10014);
nor U27856 (N_27856,N_14725,N_10270);
nand U27857 (N_27857,N_14708,N_19721);
nand U27858 (N_27858,N_13173,N_10038);
nor U27859 (N_27859,N_12478,N_13132);
and U27860 (N_27860,N_13721,N_10569);
nor U27861 (N_27861,N_14149,N_16703);
xor U27862 (N_27862,N_18859,N_19251);
or U27863 (N_27863,N_11745,N_17043);
or U27864 (N_27864,N_11356,N_17243);
or U27865 (N_27865,N_12488,N_18415);
nand U27866 (N_27866,N_11883,N_17590);
and U27867 (N_27867,N_16645,N_11268);
nor U27868 (N_27868,N_14368,N_19141);
xnor U27869 (N_27869,N_14356,N_16502);
or U27870 (N_27870,N_11819,N_10420);
xnor U27871 (N_27871,N_14075,N_17312);
nor U27872 (N_27872,N_19796,N_11018);
or U27873 (N_27873,N_19259,N_14801);
nand U27874 (N_27874,N_14609,N_16243);
xnor U27875 (N_27875,N_17526,N_16717);
nand U27876 (N_27876,N_13576,N_10955);
xnor U27877 (N_27877,N_12650,N_11958);
nor U27878 (N_27878,N_14973,N_10040);
or U27879 (N_27879,N_10822,N_16264);
and U27880 (N_27880,N_15928,N_14628);
xor U27881 (N_27881,N_15397,N_18603);
nand U27882 (N_27882,N_11376,N_16886);
and U27883 (N_27883,N_17494,N_19334);
nor U27884 (N_27884,N_15850,N_18818);
or U27885 (N_27885,N_18745,N_19383);
and U27886 (N_27886,N_13547,N_12008);
and U27887 (N_27887,N_19715,N_19250);
or U27888 (N_27888,N_17868,N_14794);
and U27889 (N_27889,N_18856,N_10177);
nor U27890 (N_27890,N_14239,N_12550);
xnor U27891 (N_27891,N_16518,N_18063);
xnor U27892 (N_27892,N_15593,N_18793);
xor U27893 (N_27893,N_17161,N_11360);
nor U27894 (N_27894,N_11209,N_14728);
or U27895 (N_27895,N_18938,N_13801);
or U27896 (N_27896,N_17364,N_19924);
nand U27897 (N_27897,N_11902,N_13428);
nor U27898 (N_27898,N_14656,N_17148);
and U27899 (N_27899,N_18079,N_17954);
nand U27900 (N_27900,N_11117,N_16669);
nor U27901 (N_27901,N_17510,N_11245);
nand U27902 (N_27902,N_19603,N_15882);
nand U27903 (N_27903,N_18983,N_13845);
nand U27904 (N_27904,N_16795,N_11219);
or U27905 (N_27905,N_12733,N_14476);
nor U27906 (N_27906,N_14550,N_13252);
or U27907 (N_27907,N_15725,N_18929);
nand U27908 (N_27908,N_12665,N_16024);
or U27909 (N_27909,N_13957,N_12469);
and U27910 (N_27910,N_14749,N_15539);
nand U27911 (N_27911,N_10377,N_15441);
nor U27912 (N_27912,N_13510,N_18731);
nand U27913 (N_27913,N_16194,N_13937);
nand U27914 (N_27914,N_16429,N_11100);
nand U27915 (N_27915,N_19250,N_11334);
and U27916 (N_27916,N_18901,N_14647);
and U27917 (N_27917,N_10187,N_17223);
or U27918 (N_27918,N_19207,N_17197);
and U27919 (N_27919,N_14601,N_16923);
nor U27920 (N_27920,N_14667,N_15937);
nand U27921 (N_27921,N_17710,N_19429);
nand U27922 (N_27922,N_16918,N_18540);
and U27923 (N_27923,N_13295,N_15985);
or U27924 (N_27924,N_18316,N_14415);
or U27925 (N_27925,N_11772,N_12256);
xor U27926 (N_27926,N_16688,N_17046);
and U27927 (N_27927,N_19608,N_15106);
or U27928 (N_27928,N_17365,N_10938);
xor U27929 (N_27929,N_12894,N_18946);
nand U27930 (N_27930,N_18550,N_18849);
nand U27931 (N_27931,N_18479,N_16745);
and U27932 (N_27932,N_13027,N_12005);
nand U27933 (N_27933,N_12314,N_18662);
and U27934 (N_27934,N_12927,N_18762);
nand U27935 (N_27935,N_16726,N_16412);
and U27936 (N_27936,N_10611,N_15551);
nor U27937 (N_27937,N_15357,N_16398);
or U27938 (N_27938,N_16335,N_10664);
or U27939 (N_27939,N_16059,N_14327);
and U27940 (N_27940,N_18918,N_14067);
nand U27941 (N_27941,N_12679,N_16951);
xnor U27942 (N_27942,N_11548,N_19165);
or U27943 (N_27943,N_15145,N_11000);
nand U27944 (N_27944,N_16436,N_18492);
nor U27945 (N_27945,N_13736,N_12695);
nor U27946 (N_27946,N_10066,N_12922);
or U27947 (N_27947,N_18840,N_16377);
or U27948 (N_27948,N_10810,N_14998);
nor U27949 (N_27949,N_16412,N_15114);
or U27950 (N_27950,N_16878,N_15699);
or U27951 (N_27951,N_14978,N_18427);
nand U27952 (N_27952,N_13018,N_19236);
or U27953 (N_27953,N_11928,N_14596);
and U27954 (N_27954,N_17110,N_15716);
or U27955 (N_27955,N_18309,N_11309);
nand U27956 (N_27956,N_17512,N_10019);
nor U27957 (N_27957,N_11627,N_18493);
nor U27958 (N_27958,N_18653,N_15186);
nor U27959 (N_27959,N_19472,N_17381);
nor U27960 (N_27960,N_10733,N_14282);
or U27961 (N_27961,N_16492,N_18860);
and U27962 (N_27962,N_15501,N_19816);
nor U27963 (N_27963,N_18791,N_18788);
xor U27964 (N_27964,N_10992,N_14143);
and U27965 (N_27965,N_10589,N_18275);
or U27966 (N_27966,N_17298,N_16493);
nand U27967 (N_27967,N_18600,N_18895);
xnor U27968 (N_27968,N_13293,N_16180);
and U27969 (N_27969,N_18159,N_18429);
and U27970 (N_27970,N_18386,N_18615);
and U27971 (N_27971,N_18867,N_12716);
or U27972 (N_27972,N_14305,N_17715);
nor U27973 (N_27973,N_13405,N_11192);
and U27974 (N_27974,N_13243,N_12087);
nand U27975 (N_27975,N_12997,N_12026);
nand U27976 (N_27976,N_12901,N_19085);
nand U27977 (N_27977,N_19547,N_14902);
and U27978 (N_27978,N_13838,N_16313);
nor U27979 (N_27979,N_10902,N_12149);
nor U27980 (N_27980,N_16734,N_14445);
nor U27981 (N_27981,N_15995,N_15461);
nor U27982 (N_27982,N_17272,N_15923);
nand U27983 (N_27983,N_16941,N_19609);
nor U27984 (N_27984,N_10812,N_10519);
nand U27985 (N_27985,N_12547,N_12301);
nor U27986 (N_27986,N_13771,N_13869);
nor U27987 (N_27987,N_17249,N_16715);
nor U27988 (N_27988,N_17587,N_19081);
xnor U27989 (N_27989,N_17395,N_12334);
nand U27990 (N_27990,N_13770,N_16382);
and U27991 (N_27991,N_11529,N_13645);
nor U27992 (N_27992,N_15215,N_16260);
and U27993 (N_27993,N_15796,N_19053);
nor U27994 (N_27994,N_17713,N_19522);
nor U27995 (N_27995,N_14735,N_16178);
nand U27996 (N_27996,N_10657,N_17578);
xor U27997 (N_27997,N_12146,N_10667);
nor U27998 (N_27998,N_13199,N_17602);
and U27999 (N_27999,N_11339,N_19115);
and U28000 (N_28000,N_12656,N_10378);
nor U28001 (N_28001,N_10978,N_19371);
nor U28002 (N_28002,N_15628,N_17219);
and U28003 (N_28003,N_14190,N_19202);
nor U28004 (N_28004,N_16875,N_13607);
nor U28005 (N_28005,N_17160,N_15241);
nor U28006 (N_28006,N_18732,N_13913);
or U28007 (N_28007,N_10891,N_18797);
nand U28008 (N_28008,N_19243,N_10535);
xor U28009 (N_28009,N_13917,N_15150);
and U28010 (N_28010,N_13926,N_10170);
or U28011 (N_28011,N_10714,N_19248);
xnor U28012 (N_28012,N_16082,N_18196);
or U28013 (N_28013,N_12365,N_16037);
xnor U28014 (N_28014,N_17407,N_13625);
nand U28015 (N_28015,N_14213,N_14465);
nand U28016 (N_28016,N_13647,N_18713);
xor U28017 (N_28017,N_19895,N_19499);
nand U28018 (N_28018,N_18870,N_10001);
or U28019 (N_28019,N_16141,N_12955);
and U28020 (N_28020,N_11321,N_16064);
nor U28021 (N_28021,N_12186,N_11225);
or U28022 (N_28022,N_18747,N_15509);
xor U28023 (N_28023,N_14960,N_17220);
nand U28024 (N_28024,N_19525,N_19333);
and U28025 (N_28025,N_16708,N_17803);
nand U28026 (N_28026,N_15625,N_17030);
and U28027 (N_28027,N_16320,N_11059);
nor U28028 (N_28028,N_14184,N_10061);
or U28029 (N_28029,N_15036,N_10347);
nand U28030 (N_28030,N_19217,N_12690);
nand U28031 (N_28031,N_14544,N_14922);
or U28032 (N_28032,N_17576,N_15382);
nand U28033 (N_28033,N_16671,N_18867);
and U28034 (N_28034,N_10159,N_18892);
and U28035 (N_28035,N_19622,N_13430);
xnor U28036 (N_28036,N_16397,N_12204);
xnor U28037 (N_28037,N_17690,N_19156);
nand U28038 (N_28038,N_11609,N_12247);
xnor U28039 (N_28039,N_15366,N_16129);
nor U28040 (N_28040,N_11301,N_16673);
nand U28041 (N_28041,N_17430,N_13452);
nand U28042 (N_28042,N_15010,N_16513);
nor U28043 (N_28043,N_19743,N_10183);
xnor U28044 (N_28044,N_18387,N_15489);
nor U28045 (N_28045,N_19088,N_11422);
nor U28046 (N_28046,N_12401,N_14859);
and U28047 (N_28047,N_17075,N_16654);
or U28048 (N_28048,N_15937,N_19754);
nand U28049 (N_28049,N_18962,N_17645);
xor U28050 (N_28050,N_12753,N_14041);
or U28051 (N_28051,N_12925,N_17385);
nor U28052 (N_28052,N_15886,N_15709);
nor U28053 (N_28053,N_14742,N_12008);
or U28054 (N_28054,N_15767,N_12844);
xor U28055 (N_28055,N_12581,N_15628);
nor U28056 (N_28056,N_11618,N_12670);
nand U28057 (N_28057,N_14960,N_14679);
nand U28058 (N_28058,N_17293,N_12326);
and U28059 (N_28059,N_13522,N_11690);
or U28060 (N_28060,N_15597,N_10142);
and U28061 (N_28061,N_12531,N_19086);
nand U28062 (N_28062,N_13892,N_19911);
nor U28063 (N_28063,N_18014,N_11697);
or U28064 (N_28064,N_19346,N_17206);
xnor U28065 (N_28065,N_14599,N_16395);
and U28066 (N_28066,N_18213,N_19845);
or U28067 (N_28067,N_11081,N_12065);
and U28068 (N_28068,N_14628,N_16871);
and U28069 (N_28069,N_17790,N_11152);
nor U28070 (N_28070,N_15762,N_17750);
and U28071 (N_28071,N_16245,N_10019);
or U28072 (N_28072,N_12324,N_12723);
or U28073 (N_28073,N_15566,N_11886);
and U28074 (N_28074,N_13118,N_11240);
xnor U28075 (N_28075,N_15576,N_16323);
or U28076 (N_28076,N_10819,N_15874);
nand U28077 (N_28077,N_17909,N_14407);
xnor U28078 (N_28078,N_15080,N_10405);
nand U28079 (N_28079,N_18529,N_14854);
nand U28080 (N_28080,N_13516,N_15385);
and U28081 (N_28081,N_18394,N_13352);
and U28082 (N_28082,N_16397,N_15225);
nand U28083 (N_28083,N_15373,N_14657);
nor U28084 (N_28084,N_10199,N_16444);
xnor U28085 (N_28085,N_15582,N_17115);
and U28086 (N_28086,N_11305,N_18196);
nor U28087 (N_28087,N_16989,N_12258);
and U28088 (N_28088,N_15416,N_11142);
and U28089 (N_28089,N_10217,N_16154);
and U28090 (N_28090,N_11349,N_11604);
and U28091 (N_28091,N_10858,N_15581);
and U28092 (N_28092,N_11654,N_16647);
nand U28093 (N_28093,N_18047,N_10771);
or U28094 (N_28094,N_15676,N_16856);
nor U28095 (N_28095,N_17126,N_13169);
and U28096 (N_28096,N_18310,N_11366);
or U28097 (N_28097,N_17650,N_16290);
or U28098 (N_28098,N_16736,N_11504);
nor U28099 (N_28099,N_12860,N_10026);
nor U28100 (N_28100,N_10995,N_14765);
or U28101 (N_28101,N_10126,N_10441);
nand U28102 (N_28102,N_12930,N_16380);
xor U28103 (N_28103,N_15095,N_12668);
nand U28104 (N_28104,N_17213,N_18665);
and U28105 (N_28105,N_18280,N_18932);
or U28106 (N_28106,N_17973,N_12557);
xnor U28107 (N_28107,N_13962,N_11225);
or U28108 (N_28108,N_15144,N_16471);
nor U28109 (N_28109,N_11186,N_19545);
and U28110 (N_28110,N_15750,N_19338);
and U28111 (N_28111,N_17266,N_17329);
nand U28112 (N_28112,N_10576,N_10347);
and U28113 (N_28113,N_15861,N_17089);
nor U28114 (N_28114,N_12464,N_11793);
nor U28115 (N_28115,N_15697,N_12394);
or U28116 (N_28116,N_10614,N_11650);
or U28117 (N_28117,N_15120,N_17014);
and U28118 (N_28118,N_12402,N_14785);
and U28119 (N_28119,N_19554,N_11790);
nor U28120 (N_28120,N_14181,N_19740);
or U28121 (N_28121,N_17279,N_16241);
xor U28122 (N_28122,N_16070,N_17717);
xor U28123 (N_28123,N_15445,N_12544);
or U28124 (N_28124,N_16827,N_15680);
nand U28125 (N_28125,N_10378,N_17809);
xor U28126 (N_28126,N_16247,N_19277);
and U28127 (N_28127,N_11716,N_16719);
xor U28128 (N_28128,N_19800,N_14833);
nand U28129 (N_28129,N_10187,N_17706);
xnor U28130 (N_28130,N_13540,N_11417);
and U28131 (N_28131,N_13259,N_16129);
or U28132 (N_28132,N_14453,N_16565);
or U28133 (N_28133,N_14597,N_19850);
and U28134 (N_28134,N_16672,N_19116);
nor U28135 (N_28135,N_10176,N_17608);
and U28136 (N_28136,N_17274,N_18209);
nor U28137 (N_28137,N_17970,N_18312);
nor U28138 (N_28138,N_19951,N_11311);
or U28139 (N_28139,N_15187,N_13633);
or U28140 (N_28140,N_17353,N_17314);
nand U28141 (N_28141,N_16326,N_10907);
or U28142 (N_28142,N_13321,N_14844);
or U28143 (N_28143,N_11067,N_19139);
and U28144 (N_28144,N_13885,N_18606);
or U28145 (N_28145,N_16787,N_11425);
or U28146 (N_28146,N_17409,N_18795);
or U28147 (N_28147,N_16368,N_17093);
nand U28148 (N_28148,N_10528,N_17657);
and U28149 (N_28149,N_15149,N_17278);
nor U28150 (N_28150,N_12563,N_17025);
nor U28151 (N_28151,N_16579,N_15243);
xnor U28152 (N_28152,N_19079,N_17148);
or U28153 (N_28153,N_17746,N_19950);
xnor U28154 (N_28154,N_15255,N_19635);
and U28155 (N_28155,N_10582,N_14573);
nand U28156 (N_28156,N_17340,N_13108);
or U28157 (N_28157,N_18642,N_18627);
or U28158 (N_28158,N_14539,N_12101);
and U28159 (N_28159,N_10475,N_10683);
or U28160 (N_28160,N_14116,N_11829);
nand U28161 (N_28161,N_18352,N_18848);
and U28162 (N_28162,N_12032,N_12714);
or U28163 (N_28163,N_10036,N_19934);
nand U28164 (N_28164,N_11128,N_13298);
and U28165 (N_28165,N_13241,N_10738);
xor U28166 (N_28166,N_19668,N_13919);
nor U28167 (N_28167,N_16701,N_10190);
and U28168 (N_28168,N_15020,N_10085);
or U28169 (N_28169,N_12390,N_10973);
and U28170 (N_28170,N_16767,N_13156);
or U28171 (N_28171,N_11884,N_13113);
and U28172 (N_28172,N_13180,N_12825);
nand U28173 (N_28173,N_13173,N_13986);
xnor U28174 (N_28174,N_18951,N_18807);
xnor U28175 (N_28175,N_13935,N_17346);
nand U28176 (N_28176,N_19885,N_14920);
nand U28177 (N_28177,N_12991,N_15768);
xor U28178 (N_28178,N_13744,N_18037);
nor U28179 (N_28179,N_16432,N_19640);
nor U28180 (N_28180,N_11481,N_15869);
nand U28181 (N_28181,N_12960,N_18731);
or U28182 (N_28182,N_18033,N_19996);
nand U28183 (N_28183,N_12022,N_16930);
nor U28184 (N_28184,N_12753,N_19032);
and U28185 (N_28185,N_11333,N_14064);
or U28186 (N_28186,N_10203,N_18548);
nand U28187 (N_28187,N_18078,N_19946);
or U28188 (N_28188,N_12536,N_14425);
or U28189 (N_28189,N_16466,N_11713);
or U28190 (N_28190,N_10345,N_16475);
xnor U28191 (N_28191,N_18423,N_16518);
or U28192 (N_28192,N_19447,N_11543);
or U28193 (N_28193,N_14180,N_17823);
xor U28194 (N_28194,N_11648,N_10684);
or U28195 (N_28195,N_15878,N_16149);
nor U28196 (N_28196,N_10589,N_16843);
nand U28197 (N_28197,N_16640,N_13312);
nor U28198 (N_28198,N_14971,N_17609);
xor U28199 (N_28199,N_14348,N_11104);
or U28200 (N_28200,N_18257,N_15568);
or U28201 (N_28201,N_19028,N_18516);
or U28202 (N_28202,N_18062,N_13000);
or U28203 (N_28203,N_13702,N_12868);
and U28204 (N_28204,N_11504,N_19023);
nor U28205 (N_28205,N_10255,N_14183);
xor U28206 (N_28206,N_13869,N_17135);
and U28207 (N_28207,N_15894,N_19792);
or U28208 (N_28208,N_10084,N_13865);
or U28209 (N_28209,N_19488,N_17228);
or U28210 (N_28210,N_13790,N_18770);
and U28211 (N_28211,N_16626,N_17919);
xor U28212 (N_28212,N_15346,N_19116);
nand U28213 (N_28213,N_19596,N_10860);
and U28214 (N_28214,N_15580,N_19550);
xnor U28215 (N_28215,N_17009,N_14898);
and U28216 (N_28216,N_15513,N_11830);
nand U28217 (N_28217,N_19182,N_19322);
nor U28218 (N_28218,N_13101,N_11456);
xnor U28219 (N_28219,N_10863,N_12038);
or U28220 (N_28220,N_18732,N_15408);
or U28221 (N_28221,N_15005,N_18172);
nand U28222 (N_28222,N_15424,N_19922);
or U28223 (N_28223,N_14385,N_16482);
or U28224 (N_28224,N_11799,N_11819);
nand U28225 (N_28225,N_19569,N_15406);
nand U28226 (N_28226,N_19095,N_10106);
nand U28227 (N_28227,N_18316,N_10033);
and U28228 (N_28228,N_18760,N_19627);
and U28229 (N_28229,N_10605,N_12874);
and U28230 (N_28230,N_12952,N_11482);
nand U28231 (N_28231,N_10611,N_15843);
nor U28232 (N_28232,N_19622,N_19310);
or U28233 (N_28233,N_18714,N_13418);
and U28234 (N_28234,N_12828,N_16567);
nor U28235 (N_28235,N_15816,N_18868);
nand U28236 (N_28236,N_15681,N_17173);
xor U28237 (N_28237,N_19249,N_15069);
nor U28238 (N_28238,N_14179,N_10047);
and U28239 (N_28239,N_13451,N_14335);
nor U28240 (N_28240,N_12013,N_14779);
and U28241 (N_28241,N_11867,N_18062);
and U28242 (N_28242,N_17586,N_11289);
or U28243 (N_28243,N_12243,N_19362);
and U28244 (N_28244,N_14959,N_16483);
nand U28245 (N_28245,N_19503,N_10155);
nand U28246 (N_28246,N_17771,N_11719);
or U28247 (N_28247,N_13934,N_15137);
xor U28248 (N_28248,N_15574,N_17591);
and U28249 (N_28249,N_14439,N_18479);
and U28250 (N_28250,N_14180,N_17947);
nand U28251 (N_28251,N_19982,N_10285);
or U28252 (N_28252,N_10909,N_11574);
and U28253 (N_28253,N_14989,N_19807);
or U28254 (N_28254,N_11665,N_16819);
and U28255 (N_28255,N_10696,N_17701);
or U28256 (N_28256,N_10263,N_12184);
xnor U28257 (N_28257,N_10694,N_15812);
nand U28258 (N_28258,N_16592,N_19378);
nand U28259 (N_28259,N_11239,N_13193);
nor U28260 (N_28260,N_16233,N_18752);
and U28261 (N_28261,N_14520,N_16418);
and U28262 (N_28262,N_11984,N_18406);
nor U28263 (N_28263,N_16016,N_16739);
and U28264 (N_28264,N_19339,N_11119);
and U28265 (N_28265,N_19732,N_18492);
and U28266 (N_28266,N_15995,N_16901);
nand U28267 (N_28267,N_15753,N_10755);
or U28268 (N_28268,N_19547,N_10628);
and U28269 (N_28269,N_12828,N_17419);
nand U28270 (N_28270,N_16462,N_14211);
nand U28271 (N_28271,N_10046,N_17826);
and U28272 (N_28272,N_10781,N_14209);
nor U28273 (N_28273,N_13222,N_15723);
nor U28274 (N_28274,N_17271,N_15622);
and U28275 (N_28275,N_10022,N_10039);
and U28276 (N_28276,N_18720,N_14444);
or U28277 (N_28277,N_18792,N_18377);
and U28278 (N_28278,N_19734,N_18182);
or U28279 (N_28279,N_16761,N_11929);
nor U28280 (N_28280,N_13235,N_14616);
and U28281 (N_28281,N_13247,N_19651);
nand U28282 (N_28282,N_12096,N_10945);
nor U28283 (N_28283,N_14844,N_19355);
or U28284 (N_28284,N_18622,N_11960);
nor U28285 (N_28285,N_15958,N_14001);
nor U28286 (N_28286,N_14845,N_14166);
nor U28287 (N_28287,N_19931,N_16882);
nand U28288 (N_28288,N_19860,N_11481);
nor U28289 (N_28289,N_18672,N_13750);
or U28290 (N_28290,N_10616,N_14772);
or U28291 (N_28291,N_15062,N_13481);
and U28292 (N_28292,N_16835,N_19472);
nor U28293 (N_28293,N_15326,N_19585);
nor U28294 (N_28294,N_12383,N_12762);
xnor U28295 (N_28295,N_16916,N_17931);
or U28296 (N_28296,N_17568,N_18792);
or U28297 (N_28297,N_16748,N_10021);
nand U28298 (N_28298,N_12163,N_17597);
xor U28299 (N_28299,N_18524,N_16447);
nand U28300 (N_28300,N_10117,N_12175);
and U28301 (N_28301,N_18223,N_15857);
nand U28302 (N_28302,N_16616,N_13036);
and U28303 (N_28303,N_15139,N_18936);
or U28304 (N_28304,N_19801,N_13524);
and U28305 (N_28305,N_11855,N_15448);
xnor U28306 (N_28306,N_16790,N_15760);
and U28307 (N_28307,N_12873,N_12365);
nand U28308 (N_28308,N_12036,N_10893);
nor U28309 (N_28309,N_19577,N_14661);
nand U28310 (N_28310,N_10694,N_14429);
nor U28311 (N_28311,N_19919,N_19917);
and U28312 (N_28312,N_19186,N_16494);
nor U28313 (N_28313,N_11623,N_14032);
nand U28314 (N_28314,N_15247,N_17462);
or U28315 (N_28315,N_11695,N_13022);
and U28316 (N_28316,N_13100,N_14088);
nor U28317 (N_28317,N_10697,N_18423);
and U28318 (N_28318,N_10057,N_19292);
or U28319 (N_28319,N_12657,N_12240);
nor U28320 (N_28320,N_18025,N_18683);
nor U28321 (N_28321,N_12205,N_17637);
and U28322 (N_28322,N_18119,N_12710);
xor U28323 (N_28323,N_14088,N_11487);
nand U28324 (N_28324,N_15187,N_15254);
nand U28325 (N_28325,N_15788,N_12458);
or U28326 (N_28326,N_16194,N_12879);
nand U28327 (N_28327,N_13238,N_17251);
nand U28328 (N_28328,N_13396,N_15181);
or U28329 (N_28329,N_19622,N_10405);
nand U28330 (N_28330,N_17119,N_18889);
and U28331 (N_28331,N_11096,N_15143);
or U28332 (N_28332,N_10753,N_17102);
nand U28333 (N_28333,N_17736,N_15393);
nand U28334 (N_28334,N_19643,N_19702);
and U28335 (N_28335,N_12531,N_11931);
and U28336 (N_28336,N_14539,N_11886);
nand U28337 (N_28337,N_16544,N_10022);
or U28338 (N_28338,N_12101,N_18670);
nand U28339 (N_28339,N_13226,N_14420);
nor U28340 (N_28340,N_12028,N_16212);
nand U28341 (N_28341,N_14258,N_17044);
nor U28342 (N_28342,N_18380,N_19826);
and U28343 (N_28343,N_15846,N_13166);
or U28344 (N_28344,N_14223,N_17113);
nor U28345 (N_28345,N_15729,N_16320);
or U28346 (N_28346,N_10444,N_10823);
nand U28347 (N_28347,N_19558,N_13727);
nor U28348 (N_28348,N_12209,N_17811);
nor U28349 (N_28349,N_15337,N_10222);
xnor U28350 (N_28350,N_12802,N_11605);
or U28351 (N_28351,N_17625,N_14795);
nand U28352 (N_28352,N_18387,N_15437);
nor U28353 (N_28353,N_16021,N_18173);
nand U28354 (N_28354,N_13291,N_17844);
nand U28355 (N_28355,N_15966,N_10928);
or U28356 (N_28356,N_12271,N_13665);
nand U28357 (N_28357,N_13037,N_17490);
or U28358 (N_28358,N_15924,N_19580);
nand U28359 (N_28359,N_16379,N_10447);
or U28360 (N_28360,N_17281,N_16552);
nor U28361 (N_28361,N_12315,N_15438);
or U28362 (N_28362,N_19421,N_10625);
or U28363 (N_28363,N_13242,N_16614);
xor U28364 (N_28364,N_11458,N_11419);
xnor U28365 (N_28365,N_13082,N_14090);
and U28366 (N_28366,N_12131,N_12629);
nand U28367 (N_28367,N_11728,N_18273);
and U28368 (N_28368,N_10277,N_10172);
nor U28369 (N_28369,N_15962,N_14741);
xnor U28370 (N_28370,N_15272,N_15850);
nand U28371 (N_28371,N_18170,N_10600);
or U28372 (N_28372,N_15364,N_14360);
xnor U28373 (N_28373,N_17890,N_10422);
nand U28374 (N_28374,N_13893,N_15980);
nor U28375 (N_28375,N_12905,N_18555);
nand U28376 (N_28376,N_12740,N_18732);
nand U28377 (N_28377,N_11834,N_15256);
nor U28378 (N_28378,N_15900,N_13762);
nor U28379 (N_28379,N_14983,N_14837);
nand U28380 (N_28380,N_11037,N_14914);
nand U28381 (N_28381,N_10459,N_17095);
nand U28382 (N_28382,N_13706,N_13627);
nand U28383 (N_28383,N_16998,N_16021);
nor U28384 (N_28384,N_10192,N_16832);
and U28385 (N_28385,N_18607,N_18299);
or U28386 (N_28386,N_13360,N_12503);
nand U28387 (N_28387,N_11609,N_19699);
or U28388 (N_28388,N_14604,N_18889);
nor U28389 (N_28389,N_16765,N_12743);
nand U28390 (N_28390,N_11669,N_10306);
and U28391 (N_28391,N_11646,N_18602);
nand U28392 (N_28392,N_10967,N_14446);
or U28393 (N_28393,N_15064,N_16715);
nor U28394 (N_28394,N_12315,N_13713);
nand U28395 (N_28395,N_16052,N_13830);
and U28396 (N_28396,N_11680,N_19386);
or U28397 (N_28397,N_18489,N_16477);
or U28398 (N_28398,N_11592,N_16434);
or U28399 (N_28399,N_13215,N_18144);
nor U28400 (N_28400,N_11211,N_12711);
or U28401 (N_28401,N_10278,N_11909);
and U28402 (N_28402,N_18278,N_17525);
nor U28403 (N_28403,N_12063,N_19550);
nand U28404 (N_28404,N_11970,N_12000);
nor U28405 (N_28405,N_14205,N_17041);
and U28406 (N_28406,N_19941,N_15351);
nor U28407 (N_28407,N_11375,N_18801);
and U28408 (N_28408,N_12013,N_19301);
and U28409 (N_28409,N_11811,N_17657);
or U28410 (N_28410,N_15499,N_17664);
xor U28411 (N_28411,N_10717,N_12967);
and U28412 (N_28412,N_17822,N_18095);
and U28413 (N_28413,N_11331,N_13788);
nor U28414 (N_28414,N_18482,N_18486);
nor U28415 (N_28415,N_10057,N_12085);
xnor U28416 (N_28416,N_15386,N_13334);
or U28417 (N_28417,N_13414,N_18835);
or U28418 (N_28418,N_19880,N_11391);
or U28419 (N_28419,N_18594,N_16529);
or U28420 (N_28420,N_15575,N_11060);
nor U28421 (N_28421,N_16204,N_14510);
or U28422 (N_28422,N_13710,N_19253);
xnor U28423 (N_28423,N_11557,N_19050);
and U28424 (N_28424,N_14718,N_16867);
and U28425 (N_28425,N_19876,N_12882);
or U28426 (N_28426,N_11621,N_16490);
nand U28427 (N_28427,N_10359,N_11327);
nor U28428 (N_28428,N_18223,N_11010);
or U28429 (N_28429,N_17127,N_10744);
and U28430 (N_28430,N_15279,N_15595);
nand U28431 (N_28431,N_17670,N_18389);
nor U28432 (N_28432,N_13716,N_17303);
or U28433 (N_28433,N_17328,N_10670);
nand U28434 (N_28434,N_12605,N_17465);
nand U28435 (N_28435,N_12155,N_15833);
or U28436 (N_28436,N_18429,N_16888);
xnor U28437 (N_28437,N_19598,N_19395);
or U28438 (N_28438,N_16583,N_18284);
nand U28439 (N_28439,N_15564,N_11457);
xnor U28440 (N_28440,N_19834,N_17356);
nand U28441 (N_28441,N_14578,N_17351);
nor U28442 (N_28442,N_10140,N_15779);
or U28443 (N_28443,N_13332,N_13432);
and U28444 (N_28444,N_17101,N_17075);
nand U28445 (N_28445,N_18402,N_12944);
or U28446 (N_28446,N_12297,N_13414);
nand U28447 (N_28447,N_11087,N_14359);
nand U28448 (N_28448,N_15043,N_11412);
nor U28449 (N_28449,N_11549,N_13489);
nand U28450 (N_28450,N_13830,N_19415);
and U28451 (N_28451,N_13432,N_14466);
and U28452 (N_28452,N_12132,N_14458);
nor U28453 (N_28453,N_14905,N_17241);
nand U28454 (N_28454,N_15512,N_12456);
nand U28455 (N_28455,N_18445,N_10992);
nor U28456 (N_28456,N_10476,N_17222);
nor U28457 (N_28457,N_18021,N_11216);
xnor U28458 (N_28458,N_18006,N_17679);
or U28459 (N_28459,N_15686,N_18123);
nand U28460 (N_28460,N_18416,N_15583);
nor U28461 (N_28461,N_16950,N_15354);
nor U28462 (N_28462,N_19187,N_12191);
and U28463 (N_28463,N_12344,N_15648);
nor U28464 (N_28464,N_18860,N_10139);
nand U28465 (N_28465,N_10039,N_11724);
nor U28466 (N_28466,N_17984,N_10784);
xnor U28467 (N_28467,N_12337,N_14175);
and U28468 (N_28468,N_11731,N_12176);
and U28469 (N_28469,N_12314,N_15588);
or U28470 (N_28470,N_16841,N_12436);
nor U28471 (N_28471,N_11748,N_18177);
nand U28472 (N_28472,N_16212,N_17996);
nand U28473 (N_28473,N_18313,N_11466);
nor U28474 (N_28474,N_13856,N_11288);
or U28475 (N_28475,N_12728,N_19994);
or U28476 (N_28476,N_11525,N_13980);
nand U28477 (N_28477,N_13587,N_10798);
and U28478 (N_28478,N_17554,N_16156);
nor U28479 (N_28479,N_12205,N_12397);
nor U28480 (N_28480,N_19356,N_18792);
nand U28481 (N_28481,N_12565,N_12609);
xor U28482 (N_28482,N_18049,N_14043);
and U28483 (N_28483,N_16675,N_19549);
and U28484 (N_28484,N_13616,N_13414);
xor U28485 (N_28485,N_11121,N_16253);
nand U28486 (N_28486,N_17982,N_10521);
xor U28487 (N_28487,N_11626,N_18566);
and U28488 (N_28488,N_12339,N_10701);
nand U28489 (N_28489,N_16507,N_15196);
or U28490 (N_28490,N_13706,N_15873);
and U28491 (N_28491,N_17513,N_14723);
xor U28492 (N_28492,N_12052,N_15551);
nand U28493 (N_28493,N_11899,N_17266);
and U28494 (N_28494,N_11192,N_10679);
nand U28495 (N_28495,N_11055,N_10470);
xnor U28496 (N_28496,N_12059,N_17390);
nor U28497 (N_28497,N_15739,N_14419);
nor U28498 (N_28498,N_18807,N_17707);
nor U28499 (N_28499,N_14004,N_13179);
and U28500 (N_28500,N_16213,N_17921);
xor U28501 (N_28501,N_16499,N_17671);
nor U28502 (N_28502,N_16869,N_11015);
and U28503 (N_28503,N_17328,N_11135);
nand U28504 (N_28504,N_14841,N_19373);
and U28505 (N_28505,N_10841,N_15132);
and U28506 (N_28506,N_13914,N_18341);
nor U28507 (N_28507,N_16632,N_12546);
nand U28508 (N_28508,N_19776,N_19475);
nor U28509 (N_28509,N_12958,N_13293);
or U28510 (N_28510,N_11775,N_18682);
nor U28511 (N_28511,N_13398,N_11951);
and U28512 (N_28512,N_14377,N_16594);
xor U28513 (N_28513,N_16582,N_14559);
nand U28514 (N_28514,N_11935,N_18509);
xor U28515 (N_28515,N_11068,N_12616);
or U28516 (N_28516,N_15843,N_14299);
and U28517 (N_28517,N_12507,N_11280);
and U28518 (N_28518,N_16595,N_19273);
or U28519 (N_28519,N_19268,N_16603);
xnor U28520 (N_28520,N_15061,N_16367);
nand U28521 (N_28521,N_17410,N_14428);
nand U28522 (N_28522,N_19035,N_11562);
or U28523 (N_28523,N_14368,N_13717);
nand U28524 (N_28524,N_17515,N_13742);
and U28525 (N_28525,N_15540,N_13930);
xor U28526 (N_28526,N_17553,N_12106);
nor U28527 (N_28527,N_17949,N_11213);
and U28528 (N_28528,N_16960,N_18243);
or U28529 (N_28529,N_16884,N_10740);
nor U28530 (N_28530,N_13321,N_13066);
and U28531 (N_28531,N_13654,N_18898);
nand U28532 (N_28532,N_17025,N_18540);
nand U28533 (N_28533,N_15526,N_17841);
or U28534 (N_28534,N_10294,N_18875);
nor U28535 (N_28535,N_10408,N_19026);
and U28536 (N_28536,N_15840,N_10452);
and U28537 (N_28537,N_15531,N_12273);
nand U28538 (N_28538,N_10503,N_17501);
and U28539 (N_28539,N_12935,N_16136);
or U28540 (N_28540,N_17319,N_18074);
nand U28541 (N_28541,N_15583,N_11251);
or U28542 (N_28542,N_13565,N_15750);
xnor U28543 (N_28543,N_11313,N_19379);
and U28544 (N_28544,N_14229,N_19941);
nand U28545 (N_28545,N_14763,N_13900);
and U28546 (N_28546,N_15519,N_13122);
and U28547 (N_28547,N_12689,N_12743);
and U28548 (N_28548,N_10996,N_14887);
or U28549 (N_28549,N_10931,N_12188);
and U28550 (N_28550,N_15663,N_14167);
or U28551 (N_28551,N_18397,N_16457);
or U28552 (N_28552,N_16543,N_10232);
nor U28553 (N_28553,N_11907,N_13560);
or U28554 (N_28554,N_11970,N_15146);
nand U28555 (N_28555,N_18312,N_19038);
nand U28556 (N_28556,N_18747,N_13144);
and U28557 (N_28557,N_12606,N_11417);
nand U28558 (N_28558,N_13530,N_12264);
or U28559 (N_28559,N_16311,N_14226);
nand U28560 (N_28560,N_11072,N_16263);
and U28561 (N_28561,N_12614,N_12436);
nand U28562 (N_28562,N_17614,N_17586);
nand U28563 (N_28563,N_16456,N_11450);
nand U28564 (N_28564,N_12019,N_18509);
nor U28565 (N_28565,N_15359,N_19955);
nor U28566 (N_28566,N_11307,N_15608);
nor U28567 (N_28567,N_18171,N_11997);
xnor U28568 (N_28568,N_16418,N_16741);
and U28569 (N_28569,N_16714,N_18132);
xnor U28570 (N_28570,N_17366,N_16093);
nand U28571 (N_28571,N_14790,N_10265);
or U28572 (N_28572,N_11078,N_16972);
and U28573 (N_28573,N_15361,N_16915);
or U28574 (N_28574,N_14135,N_12516);
and U28575 (N_28575,N_12862,N_19133);
nand U28576 (N_28576,N_12499,N_17631);
and U28577 (N_28577,N_16970,N_16748);
nor U28578 (N_28578,N_17165,N_16093);
or U28579 (N_28579,N_12748,N_12692);
nor U28580 (N_28580,N_19073,N_19774);
nor U28581 (N_28581,N_17871,N_14612);
and U28582 (N_28582,N_11234,N_16921);
or U28583 (N_28583,N_19852,N_19220);
nand U28584 (N_28584,N_12634,N_10794);
xnor U28585 (N_28585,N_11262,N_15212);
nor U28586 (N_28586,N_16552,N_18162);
or U28587 (N_28587,N_14048,N_15971);
nor U28588 (N_28588,N_18676,N_13425);
or U28589 (N_28589,N_10447,N_10194);
nor U28590 (N_28590,N_12755,N_10998);
or U28591 (N_28591,N_10922,N_19575);
nor U28592 (N_28592,N_18063,N_11141);
or U28593 (N_28593,N_15808,N_15970);
nand U28594 (N_28594,N_14971,N_12181);
nor U28595 (N_28595,N_19476,N_11440);
and U28596 (N_28596,N_10780,N_11051);
or U28597 (N_28597,N_12390,N_18497);
and U28598 (N_28598,N_16100,N_15076);
nor U28599 (N_28599,N_17731,N_14530);
nor U28600 (N_28600,N_18571,N_14250);
nand U28601 (N_28601,N_10812,N_19733);
xnor U28602 (N_28602,N_16111,N_15332);
and U28603 (N_28603,N_11097,N_11421);
nand U28604 (N_28604,N_17580,N_10189);
nand U28605 (N_28605,N_17411,N_12659);
nor U28606 (N_28606,N_18215,N_15460);
or U28607 (N_28607,N_13757,N_12998);
or U28608 (N_28608,N_10844,N_14148);
and U28609 (N_28609,N_18246,N_11829);
nor U28610 (N_28610,N_19544,N_12765);
nor U28611 (N_28611,N_15170,N_13502);
xor U28612 (N_28612,N_11365,N_11116);
nand U28613 (N_28613,N_10842,N_17212);
and U28614 (N_28614,N_14699,N_13725);
or U28615 (N_28615,N_19361,N_11753);
or U28616 (N_28616,N_10225,N_18919);
and U28617 (N_28617,N_16596,N_17512);
xnor U28618 (N_28618,N_12928,N_11775);
nor U28619 (N_28619,N_16564,N_11411);
and U28620 (N_28620,N_15589,N_10083);
nand U28621 (N_28621,N_10619,N_18188);
nand U28622 (N_28622,N_12493,N_16104);
or U28623 (N_28623,N_16253,N_14540);
nor U28624 (N_28624,N_16824,N_13293);
nand U28625 (N_28625,N_12095,N_16182);
and U28626 (N_28626,N_14148,N_15497);
nor U28627 (N_28627,N_17665,N_15904);
nor U28628 (N_28628,N_14297,N_16885);
and U28629 (N_28629,N_15789,N_12407);
nor U28630 (N_28630,N_17425,N_12716);
nand U28631 (N_28631,N_12417,N_19401);
nor U28632 (N_28632,N_19412,N_17885);
and U28633 (N_28633,N_10263,N_17630);
or U28634 (N_28634,N_10035,N_17930);
nor U28635 (N_28635,N_12158,N_19687);
and U28636 (N_28636,N_12172,N_17948);
and U28637 (N_28637,N_11053,N_12845);
xor U28638 (N_28638,N_12878,N_15495);
nand U28639 (N_28639,N_14373,N_12398);
or U28640 (N_28640,N_12794,N_11263);
and U28641 (N_28641,N_16536,N_10504);
nor U28642 (N_28642,N_18698,N_11650);
and U28643 (N_28643,N_16169,N_11855);
and U28644 (N_28644,N_16598,N_12954);
and U28645 (N_28645,N_13796,N_18085);
nor U28646 (N_28646,N_13311,N_10999);
xor U28647 (N_28647,N_12839,N_18842);
nand U28648 (N_28648,N_14523,N_12786);
xor U28649 (N_28649,N_16641,N_18186);
or U28650 (N_28650,N_14595,N_10695);
and U28651 (N_28651,N_12290,N_13859);
nand U28652 (N_28652,N_13017,N_17573);
or U28653 (N_28653,N_13731,N_10922);
nand U28654 (N_28654,N_13983,N_14189);
or U28655 (N_28655,N_11489,N_15924);
and U28656 (N_28656,N_12590,N_18225);
nand U28657 (N_28657,N_19973,N_13416);
xor U28658 (N_28658,N_18431,N_12431);
xnor U28659 (N_28659,N_13653,N_13518);
and U28660 (N_28660,N_16920,N_14728);
nor U28661 (N_28661,N_19884,N_15028);
or U28662 (N_28662,N_19589,N_11286);
and U28663 (N_28663,N_19880,N_18894);
nor U28664 (N_28664,N_15537,N_16607);
xor U28665 (N_28665,N_11810,N_18351);
nand U28666 (N_28666,N_18127,N_16831);
and U28667 (N_28667,N_18386,N_12201);
and U28668 (N_28668,N_19463,N_16786);
nor U28669 (N_28669,N_13139,N_11854);
nor U28670 (N_28670,N_11831,N_10201);
or U28671 (N_28671,N_18776,N_15163);
nand U28672 (N_28672,N_13303,N_19630);
nor U28673 (N_28673,N_18742,N_12452);
nand U28674 (N_28674,N_14235,N_14866);
or U28675 (N_28675,N_15938,N_10647);
and U28676 (N_28676,N_11451,N_18621);
nor U28677 (N_28677,N_13902,N_17798);
or U28678 (N_28678,N_13562,N_16990);
nor U28679 (N_28679,N_16707,N_12142);
and U28680 (N_28680,N_19861,N_16246);
nand U28681 (N_28681,N_12620,N_17302);
and U28682 (N_28682,N_19050,N_11826);
and U28683 (N_28683,N_12126,N_19832);
nand U28684 (N_28684,N_13821,N_12068);
and U28685 (N_28685,N_12530,N_18943);
nor U28686 (N_28686,N_19338,N_13663);
nand U28687 (N_28687,N_14187,N_10637);
or U28688 (N_28688,N_12783,N_12898);
nor U28689 (N_28689,N_16381,N_11247);
and U28690 (N_28690,N_13678,N_14005);
or U28691 (N_28691,N_12633,N_10831);
and U28692 (N_28692,N_14131,N_19017);
or U28693 (N_28693,N_10168,N_10944);
or U28694 (N_28694,N_18646,N_18644);
nand U28695 (N_28695,N_16206,N_15502);
nand U28696 (N_28696,N_15017,N_10388);
and U28697 (N_28697,N_15922,N_10331);
nand U28698 (N_28698,N_14204,N_16742);
and U28699 (N_28699,N_11123,N_18608);
nor U28700 (N_28700,N_16614,N_18137);
or U28701 (N_28701,N_10522,N_13551);
nor U28702 (N_28702,N_19514,N_14273);
nand U28703 (N_28703,N_17309,N_16368);
and U28704 (N_28704,N_10599,N_12050);
or U28705 (N_28705,N_10596,N_17214);
and U28706 (N_28706,N_16828,N_19250);
nand U28707 (N_28707,N_16985,N_11106);
or U28708 (N_28708,N_17831,N_12887);
and U28709 (N_28709,N_16588,N_13005);
nor U28710 (N_28710,N_18156,N_10645);
or U28711 (N_28711,N_13992,N_10887);
nor U28712 (N_28712,N_13812,N_19547);
nor U28713 (N_28713,N_13994,N_10573);
nand U28714 (N_28714,N_19123,N_14218);
nor U28715 (N_28715,N_11585,N_18240);
nor U28716 (N_28716,N_14488,N_14387);
nand U28717 (N_28717,N_15805,N_10868);
and U28718 (N_28718,N_14680,N_11578);
or U28719 (N_28719,N_17331,N_10959);
nand U28720 (N_28720,N_15249,N_18268);
and U28721 (N_28721,N_19835,N_15795);
xnor U28722 (N_28722,N_19416,N_11827);
nor U28723 (N_28723,N_14047,N_15258);
nor U28724 (N_28724,N_13031,N_13374);
or U28725 (N_28725,N_13907,N_15390);
nor U28726 (N_28726,N_12178,N_11290);
nand U28727 (N_28727,N_11396,N_17058);
nand U28728 (N_28728,N_14906,N_14952);
xor U28729 (N_28729,N_16314,N_18672);
nor U28730 (N_28730,N_12351,N_12656);
nor U28731 (N_28731,N_15236,N_11712);
nand U28732 (N_28732,N_10039,N_16721);
nand U28733 (N_28733,N_19618,N_14586);
xnor U28734 (N_28734,N_14175,N_17738);
nand U28735 (N_28735,N_12210,N_15339);
or U28736 (N_28736,N_19601,N_16014);
nand U28737 (N_28737,N_16488,N_11602);
and U28738 (N_28738,N_15727,N_14620);
or U28739 (N_28739,N_15787,N_15187);
or U28740 (N_28740,N_16309,N_17297);
nor U28741 (N_28741,N_16549,N_11850);
nand U28742 (N_28742,N_12343,N_13536);
and U28743 (N_28743,N_14127,N_13070);
or U28744 (N_28744,N_18274,N_14517);
and U28745 (N_28745,N_18558,N_18082);
nor U28746 (N_28746,N_18310,N_15654);
and U28747 (N_28747,N_12461,N_11697);
nor U28748 (N_28748,N_10428,N_10736);
or U28749 (N_28749,N_12544,N_18027);
or U28750 (N_28750,N_16896,N_19576);
nand U28751 (N_28751,N_17487,N_19175);
or U28752 (N_28752,N_14064,N_18820);
nor U28753 (N_28753,N_13079,N_11655);
and U28754 (N_28754,N_12414,N_16404);
xnor U28755 (N_28755,N_11561,N_19886);
or U28756 (N_28756,N_16275,N_11739);
nor U28757 (N_28757,N_11116,N_15461);
and U28758 (N_28758,N_10897,N_14721);
or U28759 (N_28759,N_12901,N_15385);
nor U28760 (N_28760,N_19844,N_13505);
nand U28761 (N_28761,N_11608,N_13584);
or U28762 (N_28762,N_14409,N_15204);
nand U28763 (N_28763,N_11067,N_13535);
or U28764 (N_28764,N_19971,N_17774);
nand U28765 (N_28765,N_15307,N_10855);
nand U28766 (N_28766,N_18842,N_15903);
or U28767 (N_28767,N_19382,N_12732);
or U28768 (N_28768,N_16318,N_17666);
nor U28769 (N_28769,N_15709,N_17740);
xnor U28770 (N_28770,N_17290,N_18413);
nor U28771 (N_28771,N_13207,N_13120);
xor U28772 (N_28772,N_19297,N_19217);
or U28773 (N_28773,N_18547,N_10499);
xor U28774 (N_28774,N_13705,N_11165);
and U28775 (N_28775,N_19438,N_10913);
nor U28776 (N_28776,N_13457,N_10029);
xor U28777 (N_28777,N_15225,N_18044);
nor U28778 (N_28778,N_16512,N_16220);
or U28779 (N_28779,N_14093,N_16471);
or U28780 (N_28780,N_10918,N_12825);
nor U28781 (N_28781,N_12661,N_11842);
xnor U28782 (N_28782,N_15563,N_18823);
and U28783 (N_28783,N_13957,N_19003);
or U28784 (N_28784,N_18277,N_18480);
nor U28785 (N_28785,N_10808,N_18046);
nor U28786 (N_28786,N_16148,N_16702);
and U28787 (N_28787,N_17273,N_12056);
nor U28788 (N_28788,N_13928,N_14693);
nor U28789 (N_28789,N_15848,N_17996);
nand U28790 (N_28790,N_17520,N_14505);
or U28791 (N_28791,N_17409,N_16308);
nand U28792 (N_28792,N_18325,N_15325);
nor U28793 (N_28793,N_15732,N_12924);
or U28794 (N_28794,N_17087,N_18360);
nand U28795 (N_28795,N_15305,N_11655);
or U28796 (N_28796,N_13014,N_11797);
nand U28797 (N_28797,N_19782,N_13662);
nand U28798 (N_28798,N_11807,N_16527);
nand U28799 (N_28799,N_14494,N_12959);
and U28800 (N_28800,N_17368,N_10517);
nand U28801 (N_28801,N_12862,N_13404);
and U28802 (N_28802,N_12324,N_14816);
xor U28803 (N_28803,N_17403,N_16372);
or U28804 (N_28804,N_14139,N_10314);
or U28805 (N_28805,N_16318,N_19170);
and U28806 (N_28806,N_13102,N_10067);
nand U28807 (N_28807,N_11574,N_14057);
nand U28808 (N_28808,N_11155,N_11410);
or U28809 (N_28809,N_12857,N_17135);
nor U28810 (N_28810,N_14572,N_16240);
or U28811 (N_28811,N_13302,N_14899);
and U28812 (N_28812,N_19028,N_13146);
nand U28813 (N_28813,N_11400,N_10252);
nand U28814 (N_28814,N_17704,N_12007);
or U28815 (N_28815,N_11691,N_13000);
and U28816 (N_28816,N_12835,N_14873);
and U28817 (N_28817,N_12963,N_15672);
and U28818 (N_28818,N_10097,N_13104);
and U28819 (N_28819,N_15589,N_17911);
xor U28820 (N_28820,N_19814,N_13162);
or U28821 (N_28821,N_11323,N_10862);
xor U28822 (N_28822,N_15707,N_16273);
nor U28823 (N_28823,N_11055,N_13741);
or U28824 (N_28824,N_10818,N_13385);
and U28825 (N_28825,N_15674,N_18146);
or U28826 (N_28826,N_10236,N_12986);
and U28827 (N_28827,N_14427,N_18086);
or U28828 (N_28828,N_17478,N_11063);
or U28829 (N_28829,N_11137,N_14751);
and U28830 (N_28830,N_18495,N_16751);
nand U28831 (N_28831,N_13113,N_13057);
nor U28832 (N_28832,N_15796,N_17767);
and U28833 (N_28833,N_14567,N_12223);
and U28834 (N_28834,N_17517,N_15802);
or U28835 (N_28835,N_15518,N_12255);
nor U28836 (N_28836,N_19432,N_12061);
and U28837 (N_28837,N_15137,N_16295);
or U28838 (N_28838,N_10043,N_14794);
nand U28839 (N_28839,N_19888,N_12082);
nor U28840 (N_28840,N_12942,N_14903);
nand U28841 (N_28841,N_19012,N_17183);
nand U28842 (N_28842,N_17063,N_15075);
or U28843 (N_28843,N_16786,N_10115);
and U28844 (N_28844,N_13249,N_16886);
nand U28845 (N_28845,N_11126,N_17125);
or U28846 (N_28846,N_16208,N_17310);
nor U28847 (N_28847,N_14741,N_13478);
nand U28848 (N_28848,N_14603,N_18800);
and U28849 (N_28849,N_18398,N_13424);
nand U28850 (N_28850,N_12489,N_11710);
nor U28851 (N_28851,N_18503,N_18441);
and U28852 (N_28852,N_14380,N_12700);
and U28853 (N_28853,N_12571,N_14891);
or U28854 (N_28854,N_18282,N_19997);
or U28855 (N_28855,N_18893,N_10672);
or U28856 (N_28856,N_15080,N_11585);
and U28857 (N_28857,N_19786,N_10208);
and U28858 (N_28858,N_10970,N_13413);
or U28859 (N_28859,N_19412,N_10126);
and U28860 (N_28860,N_18245,N_19250);
or U28861 (N_28861,N_11608,N_15961);
nor U28862 (N_28862,N_18498,N_10525);
or U28863 (N_28863,N_14728,N_17452);
and U28864 (N_28864,N_12834,N_14025);
nand U28865 (N_28865,N_14184,N_15751);
and U28866 (N_28866,N_15042,N_15383);
and U28867 (N_28867,N_18929,N_17998);
or U28868 (N_28868,N_18412,N_10023);
nor U28869 (N_28869,N_11794,N_10275);
xnor U28870 (N_28870,N_14416,N_16966);
nand U28871 (N_28871,N_17828,N_19411);
nand U28872 (N_28872,N_12247,N_19845);
or U28873 (N_28873,N_18260,N_11578);
xnor U28874 (N_28874,N_17421,N_15020);
xnor U28875 (N_28875,N_19189,N_13368);
nor U28876 (N_28876,N_16551,N_17370);
and U28877 (N_28877,N_14119,N_11486);
nor U28878 (N_28878,N_13125,N_19742);
or U28879 (N_28879,N_18391,N_12677);
nand U28880 (N_28880,N_19232,N_18376);
nand U28881 (N_28881,N_17660,N_15242);
nor U28882 (N_28882,N_10215,N_10663);
or U28883 (N_28883,N_13075,N_12660);
and U28884 (N_28884,N_18431,N_16267);
and U28885 (N_28885,N_18960,N_12987);
nor U28886 (N_28886,N_10442,N_14498);
nor U28887 (N_28887,N_17912,N_15751);
or U28888 (N_28888,N_11755,N_11078);
and U28889 (N_28889,N_13279,N_17536);
or U28890 (N_28890,N_11614,N_16416);
or U28891 (N_28891,N_16932,N_15714);
and U28892 (N_28892,N_13615,N_19008);
or U28893 (N_28893,N_12295,N_16256);
or U28894 (N_28894,N_15189,N_18275);
nor U28895 (N_28895,N_10045,N_14490);
and U28896 (N_28896,N_16795,N_11861);
and U28897 (N_28897,N_10754,N_10090);
or U28898 (N_28898,N_18918,N_14876);
nor U28899 (N_28899,N_18369,N_18102);
nor U28900 (N_28900,N_17598,N_13326);
nand U28901 (N_28901,N_17821,N_19447);
and U28902 (N_28902,N_18107,N_17189);
nand U28903 (N_28903,N_16866,N_18456);
nor U28904 (N_28904,N_15227,N_16069);
nand U28905 (N_28905,N_17994,N_10323);
or U28906 (N_28906,N_15706,N_13389);
or U28907 (N_28907,N_16728,N_12411);
nand U28908 (N_28908,N_17671,N_17614);
nor U28909 (N_28909,N_13820,N_11458);
nand U28910 (N_28910,N_19752,N_10290);
nand U28911 (N_28911,N_17371,N_19672);
nor U28912 (N_28912,N_14276,N_13309);
nand U28913 (N_28913,N_19891,N_12762);
and U28914 (N_28914,N_13187,N_12910);
nor U28915 (N_28915,N_15455,N_16062);
and U28916 (N_28916,N_11720,N_18208);
nand U28917 (N_28917,N_17139,N_16073);
nand U28918 (N_28918,N_11477,N_15102);
or U28919 (N_28919,N_14791,N_10371);
or U28920 (N_28920,N_17105,N_18148);
or U28921 (N_28921,N_13104,N_17059);
nor U28922 (N_28922,N_19646,N_18038);
xor U28923 (N_28923,N_12061,N_16488);
nand U28924 (N_28924,N_11906,N_17072);
and U28925 (N_28925,N_13566,N_11892);
xor U28926 (N_28926,N_15148,N_10132);
nor U28927 (N_28927,N_16565,N_11109);
or U28928 (N_28928,N_15502,N_11969);
or U28929 (N_28929,N_14426,N_18795);
nor U28930 (N_28930,N_17844,N_11911);
nand U28931 (N_28931,N_10359,N_19790);
nor U28932 (N_28932,N_19183,N_18049);
or U28933 (N_28933,N_11526,N_18557);
nor U28934 (N_28934,N_18837,N_12476);
and U28935 (N_28935,N_15651,N_17661);
nor U28936 (N_28936,N_17049,N_18332);
or U28937 (N_28937,N_12818,N_12158);
xor U28938 (N_28938,N_14792,N_19570);
nor U28939 (N_28939,N_18903,N_19470);
nand U28940 (N_28940,N_19475,N_11408);
or U28941 (N_28941,N_15947,N_12693);
nor U28942 (N_28942,N_14231,N_18600);
or U28943 (N_28943,N_11978,N_14289);
and U28944 (N_28944,N_11495,N_11658);
and U28945 (N_28945,N_12103,N_13686);
or U28946 (N_28946,N_14692,N_11527);
xor U28947 (N_28947,N_18356,N_12087);
or U28948 (N_28948,N_16249,N_17049);
nand U28949 (N_28949,N_19145,N_15470);
and U28950 (N_28950,N_12139,N_17920);
nor U28951 (N_28951,N_18265,N_18182);
and U28952 (N_28952,N_18938,N_17624);
nor U28953 (N_28953,N_15017,N_10477);
nor U28954 (N_28954,N_14030,N_15906);
and U28955 (N_28955,N_15701,N_19252);
nand U28956 (N_28956,N_10758,N_10781);
or U28957 (N_28957,N_19409,N_14084);
nand U28958 (N_28958,N_10325,N_11639);
or U28959 (N_28959,N_12882,N_10673);
nand U28960 (N_28960,N_17394,N_19454);
nor U28961 (N_28961,N_17704,N_13228);
nor U28962 (N_28962,N_14270,N_12403);
or U28963 (N_28963,N_19282,N_12226);
and U28964 (N_28964,N_13338,N_12756);
nand U28965 (N_28965,N_17942,N_14559);
nor U28966 (N_28966,N_10136,N_13990);
and U28967 (N_28967,N_17933,N_12835);
nand U28968 (N_28968,N_16312,N_13276);
xor U28969 (N_28969,N_12810,N_15744);
nor U28970 (N_28970,N_16172,N_15906);
xor U28971 (N_28971,N_17384,N_15961);
and U28972 (N_28972,N_15799,N_11456);
nor U28973 (N_28973,N_17698,N_10305);
nor U28974 (N_28974,N_16815,N_12342);
nor U28975 (N_28975,N_19156,N_12342);
and U28976 (N_28976,N_16587,N_11983);
nor U28977 (N_28977,N_10341,N_10786);
nand U28978 (N_28978,N_14210,N_18836);
nor U28979 (N_28979,N_13697,N_14188);
nand U28980 (N_28980,N_17099,N_19617);
and U28981 (N_28981,N_19059,N_14086);
or U28982 (N_28982,N_19617,N_15816);
and U28983 (N_28983,N_10890,N_10550);
and U28984 (N_28984,N_18370,N_10027);
nand U28985 (N_28985,N_17100,N_18505);
and U28986 (N_28986,N_12144,N_18073);
nand U28987 (N_28987,N_19074,N_15110);
and U28988 (N_28988,N_16161,N_10056);
xnor U28989 (N_28989,N_12951,N_17576);
nor U28990 (N_28990,N_16777,N_17921);
or U28991 (N_28991,N_13693,N_17476);
nor U28992 (N_28992,N_17806,N_17310);
nor U28993 (N_28993,N_17658,N_17398);
or U28994 (N_28994,N_12675,N_17201);
or U28995 (N_28995,N_16767,N_14337);
and U28996 (N_28996,N_14024,N_15759);
nand U28997 (N_28997,N_17131,N_19086);
or U28998 (N_28998,N_16468,N_10548);
nand U28999 (N_28999,N_11570,N_12947);
nand U29000 (N_29000,N_17328,N_15779);
xnor U29001 (N_29001,N_17414,N_15064);
and U29002 (N_29002,N_19471,N_10852);
or U29003 (N_29003,N_17836,N_13649);
xnor U29004 (N_29004,N_15343,N_18061);
or U29005 (N_29005,N_18739,N_17705);
nand U29006 (N_29006,N_17170,N_12009);
nand U29007 (N_29007,N_13494,N_10755);
xor U29008 (N_29008,N_14864,N_13456);
nor U29009 (N_29009,N_10362,N_15435);
nand U29010 (N_29010,N_17410,N_12442);
nor U29011 (N_29011,N_16089,N_16125);
and U29012 (N_29012,N_10934,N_12274);
nand U29013 (N_29013,N_18600,N_13162);
or U29014 (N_29014,N_12369,N_15602);
and U29015 (N_29015,N_19673,N_14007);
or U29016 (N_29016,N_10754,N_11119);
or U29017 (N_29017,N_15301,N_16504);
or U29018 (N_29018,N_16707,N_10966);
or U29019 (N_29019,N_15347,N_15839);
or U29020 (N_29020,N_16053,N_19410);
nor U29021 (N_29021,N_12671,N_12609);
and U29022 (N_29022,N_16552,N_12664);
nand U29023 (N_29023,N_17301,N_12450);
nor U29024 (N_29024,N_15540,N_19098);
or U29025 (N_29025,N_13857,N_15136);
nor U29026 (N_29026,N_19950,N_10543);
nor U29027 (N_29027,N_15445,N_16005);
and U29028 (N_29028,N_15429,N_14342);
xnor U29029 (N_29029,N_19025,N_14507);
nand U29030 (N_29030,N_10854,N_11042);
or U29031 (N_29031,N_10275,N_12268);
and U29032 (N_29032,N_14570,N_13912);
or U29033 (N_29033,N_12738,N_10272);
or U29034 (N_29034,N_17769,N_18831);
nor U29035 (N_29035,N_13586,N_17252);
nor U29036 (N_29036,N_12664,N_17507);
nand U29037 (N_29037,N_15228,N_13197);
nand U29038 (N_29038,N_13696,N_19897);
and U29039 (N_29039,N_12255,N_16806);
and U29040 (N_29040,N_10256,N_18935);
nand U29041 (N_29041,N_13969,N_13597);
or U29042 (N_29042,N_12623,N_10639);
or U29043 (N_29043,N_11088,N_13098);
nor U29044 (N_29044,N_11176,N_11332);
nor U29045 (N_29045,N_12568,N_10051);
nand U29046 (N_29046,N_17686,N_15185);
nand U29047 (N_29047,N_15215,N_11634);
nand U29048 (N_29048,N_12016,N_17127);
and U29049 (N_29049,N_12906,N_17418);
or U29050 (N_29050,N_16487,N_11283);
xnor U29051 (N_29051,N_13737,N_17142);
and U29052 (N_29052,N_11603,N_14623);
nor U29053 (N_29053,N_18025,N_13796);
xor U29054 (N_29054,N_10372,N_13042);
nor U29055 (N_29055,N_19347,N_13291);
and U29056 (N_29056,N_18847,N_14305);
nand U29057 (N_29057,N_13884,N_11605);
and U29058 (N_29058,N_10595,N_14896);
and U29059 (N_29059,N_13256,N_11647);
nor U29060 (N_29060,N_19825,N_10830);
or U29061 (N_29061,N_16697,N_19652);
nand U29062 (N_29062,N_17725,N_11069);
and U29063 (N_29063,N_19931,N_15542);
nor U29064 (N_29064,N_19959,N_10638);
nor U29065 (N_29065,N_13932,N_10752);
nor U29066 (N_29066,N_18275,N_14289);
nor U29067 (N_29067,N_17448,N_13762);
nand U29068 (N_29068,N_15084,N_17782);
nand U29069 (N_29069,N_10269,N_17475);
nand U29070 (N_29070,N_19329,N_12915);
or U29071 (N_29071,N_16596,N_17280);
and U29072 (N_29072,N_16295,N_14611);
nand U29073 (N_29073,N_18473,N_19364);
or U29074 (N_29074,N_11628,N_10653);
and U29075 (N_29075,N_15585,N_15431);
nor U29076 (N_29076,N_14627,N_10558);
and U29077 (N_29077,N_12932,N_15951);
or U29078 (N_29078,N_17858,N_10649);
or U29079 (N_29079,N_14504,N_10172);
or U29080 (N_29080,N_10685,N_12037);
nand U29081 (N_29081,N_16159,N_16170);
or U29082 (N_29082,N_11597,N_16133);
nand U29083 (N_29083,N_19587,N_13419);
xnor U29084 (N_29084,N_19309,N_18328);
and U29085 (N_29085,N_10667,N_12481);
and U29086 (N_29086,N_18015,N_17804);
nor U29087 (N_29087,N_11923,N_10559);
xor U29088 (N_29088,N_10112,N_13840);
xor U29089 (N_29089,N_13738,N_17948);
nand U29090 (N_29090,N_13554,N_19381);
nor U29091 (N_29091,N_18269,N_15146);
nor U29092 (N_29092,N_15868,N_10693);
xor U29093 (N_29093,N_19575,N_18678);
and U29094 (N_29094,N_15861,N_17441);
nor U29095 (N_29095,N_16883,N_10858);
nand U29096 (N_29096,N_16717,N_11910);
nor U29097 (N_29097,N_18321,N_13476);
or U29098 (N_29098,N_19463,N_15376);
and U29099 (N_29099,N_15353,N_14230);
and U29100 (N_29100,N_16566,N_10834);
nand U29101 (N_29101,N_12791,N_11358);
and U29102 (N_29102,N_14049,N_10550);
and U29103 (N_29103,N_18843,N_12960);
or U29104 (N_29104,N_15179,N_12829);
and U29105 (N_29105,N_11941,N_18761);
nor U29106 (N_29106,N_16772,N_13232);
xnor U29107 (N_29107,N_13066,N_13703);
nor U29108 (N_29108,N_16725,N_12527);
and U29109 (N_29109,N_17651,N_19515);
or U29110 (N_29110,N_13328,N_13688);
nand U29111 (N_29111,N_13470,N_14611);
nor U29112 (N_29112,N_18250,N_18310);
or U29113 (N_29113,N_14576,N_10396);
or U29114 (N_29114,N_14143,N_17240);
nand U29115 (N_29115,N_18076,N_17202);
nand U29116 (N_29116,N_14850,N_16091);
xor U29117 (N_29117,N_19768,N_18177);
and U29118 (N_29118,N_13387,N_14327);
nand U29119 (N_29119,N_11870,N_18615);
nand U29120 (N_29120,N_11256,N_16446);
and U29121 (N_29121,N_15297,N_17343);
or U29122 (N_29122,N_15250,N_17468);
or U29123 (N_29123,N_13149,N_17039);
and U29124 (N_29124,N_11361,N_11251);
xnor U29125 (N_29125,N_12320,N_12309);
nor U29126 (N_29126,N_12242,N_17578);
xnor U29127 (N_29127,N_16207,N_19083);
and U29128 (N_29128,N_10119,N_10605);
nor U29129 (N_29129,N_17131,N_14769);
nand U29130 (N_29130,N_19365,N_12291);
nor U29131 (N_29131,N_16441,N_14253);
nand U29132 (N_29132,N_10201,N_17169);
nor U29133 (N_29133,N_10212,N_11310);
xnor U29134 (N_29134,N_11464,N_16406);
xor U29135 (N_29135,N_11737,N_15738);
or U29136 (N_29136,N_11521,N_18112);
nor U29137 (N_29137,N_17234,N_13301);
nand U29138 (N_29138,N_12181,N_16713);
or U29139 (N_29139,N_16691,N_10047);
or U29140 (N_29140,N_11164,N_18786);
nand U29141 (N_29141,N_16947,N_12372);
and U29142 (N_29142,N_11915,N_11614);
xor U29143 (N_29143,N_18744,N_11671);
and U29144 (N_29144,N_17055,N_14660);
nand U29145 (N_29145,N_18267,N_16591);
nor U29146 (N_29146,N_10812,N_11699);
or U29147 (N_29147,N_13243,N_10500);
nand U29148 (N_29148,N_18626,N_19142);
and U29149 (N_29149,N_14420,N_17009);
nand U29150 (N_29150,N_19763,N_11436);
nor U29151 (N_29151,N_15350,N_14975);
and U29152 (N_29152,N_19275,N_12111);
or U29153 (N_29153,N_16151,N_14907);
nor U29154 (N_29154,N_11081,N_17617);
and U29155 (N_29155,N_12062,N_11648);
or U29156 (N_29156,N_11159,N_18821);
nor U29157 (N_29157,N_10033,N_18586);
or U29158 (N_29158,N_15245,N_14047);
nor U29159 (N_29159,N_15856,N_18777);
nand U29160 (N_29160,N_19056,N_11164);
nand U29161 (N_29161,N_16028,N_14719);
or U29162 (N_29162,N_15024,N_11560);
xor U29163 (N_29163,N_10450,N_14730);
nor U29164 (N_29164,N_17568,N_17526);
nand U29165 (N_29165,N_15727,N_19731);
nand U29166 (N_29166,N_14753,N_15239);
nor U29167 (N_29167,N_19449,N_14501);
or U29168 (N_29168,N_15660,N_15210);
nand U29169 (N_29169,N_18050,N_14744);
nand U29170 (N_29170,N_18271,N_11910);
nand U29171 (N_29171,N_14866,N_17421);
nor U29172 (N_29172,N_13187,N_19783);
or U29173 (N_29173,N_12146,N_11206);
or U29174 (N_29174,N_16042,N_19403);
nand U29175 (N_29175,N_16974,N_14818);
nor U29176 (N_29176,N_10942,N_11341);
nor U29177 (N_29177,N_14264,N_10010);
nand U29178 (N_29178,N_14952,N_18633);
or U29179 (N_29179,N_15758,N_19171);
nor U29180 (N_29180,N_16654,N_12599);
or U29181 (N_29181,N_11680,N_18674);
nand U29182 (N_29182,N_18074,N_17445);
and U29183 (N_29183,N_18353,N_15706);
or U29184 (N_29184,N_11863,N_17612);
or U29185 (N_29185,N_17948,N_15952);
nor U29186 (N_29186,N_13321,N_18689);
nand U29187 (N_29187,N_10456,N_14505);
nand U29188 (N_29188,N_17642,N_15052);
nand U29189 (N_29189,N_11009,N_18752);
xnor U29190 (N_29190,N_15303,N_13369);
nor U29191 (N_29191,N_10249,N_10403);
or U29192 (N_29192,N_11193,N_12295);
and U29193 (N_29193,N_17438,N_17056);
nor U29194 (N_29194,N_14321,N_10060);
or U29195 (N_29195,N_11243,N_17462);
nor U29196 (N_29196,N_10919,N_12412);
nor U29197 (N_29197,N_17711,N_12036);
nor U29198 (N_29198,N_16830,N_12797);
nand U29199 (N_29199,N_19953,N_12161);
and U29200 (N_29200,N_12200,N_10419);
and U29201 (N_29201,N_18026,N_15256);
and U29202 (N_29202,N_11890,N_13944);
and U29203 (N_29203,N_17634,N_13267);
and U29204 (N_29204,N_11903,N_18144);
and U29205 (N_29205,N_14158,N_16115);
and U29206 (N_29206,N_17857,N_12680);
and U29207 (N_29207,N_14570,N_12084);
nor U29208 (N_29208,N_19020,N_11084);
and U29209 (N_29209,N_15160,N_15996);
and U29210 (N_29210,N_18522,N_12099);
or U29211 (N_29211,N_15826,N_12700);
nor U29212 (N_29212,N_16735,N_15229);
and U29213 (N_29213,N_13114,N_12919);
nand U29214 (N_29214,N_17179,N_12145);
nand U29215 (N_29215,N_12434,N_10316);
nor U29216 (N_29216,N_10796,N_11811);
xnor U29217 (N_29217,N_12547,N_13163);
and U29218 (N_29218,N_13725,N_17356);
or U29219 (N_29219,N_19907,N_14662);
nor U29220 (N_29220,N_14371,N_12641);
nor U29221 (N_29221,N_18665,N_15161);
xor U29222 (N_29222,N_12045,N_19320);
or U29223 (N_29223,N_18169,N_17885);
and U29224 (N_29224,N_18066,N_11573);
or U29225 (N_29225,N_13854,N_12024);
xnor U29226 (N_29226,N_17569,N_18379);
or U29227 (N_29227,N_14437,N_13289);
nor U29228 (N_29228,N_14841,N_17584);
nor U29229 (N_29229,N_10152,N_16644);
nand U29230 (N_29230,N_14146,N_12451);
or U29231 (N_29231,N_18609,N_18975);
nor U29232 (N_29232,N_11860,N_18574);
and U29233 (N_29233,N_12018,N_16317);
or U29234 (N_29234,N_18180,N_15741);
nor U29235 (N_29235,N_18206,N_10029);
nor U29236 (N_29236,N_18317,N_19428);
nand U29237 (N_29237,N_17869,N_10927);
or U29238 (N_29238,N_17214,N_15472);
nand U29239 (N_29239,N_16215,N_13574);
nor U29240 (N_29240,N_17378,N_17820);
nor U29241 (N_29241,N_16203,N_10307);
xor U29242 (N_29242,N_17465,N_13706);
and U29243 (N_29243,N_18846,N_12682);
or U29244 (N_29244,N_12329,N_18662);
or U29245 (N_29245,N_10730,N_10736);
or U29246 (N_29246,N_17223,N_10518);
nand U29247 (N_29247,N_19247,N_17856);
nand U29248 (N_29248,N_12414,N_14106);
nor U29249 (N_29249,N_19698,N_10826);
and U29250 (N_29250,N_15589,N_17517);
nand U29251 (N_29251,N_17036,N_15679);
xor U29252 (N_29252,N_12029,N_13463);
nand U29253 (N_29253,N_14238,N_10812);
nand U29254 (N_29254,N_18532,N_18456);
nand U29255 (N_29255,N_18845,N_13745);
and U29256 (N_29256,N_18782,N_14273);
nand U29257 (N_29257,N_12285,N_10505);
nor U29258 (N_29258,N_18210,N_17318);
or U29259 (N_29259,N_13295,N_18542);
nand U29260 (N_29260,N_19081,N_10586);
nand U29261 (N_29261,N_10111,N_17866);
and U29262 (N_29262,N_16316,N_16914);
xnor U29263 (N_29263,N_12601,N_16836);
and U29264 (N_29264,N_16934,N_11460);
nor U29265 (N_29265,N_11212,N_17819);
nor U29266 (N_29266,N_19272,N_17976);
xnor U29267 (N_29267,N_13672,N_12995);
nor U29268 (N_29268,N_17612,N_11931);
nand U29269 (N_29269,N_19666,N_10215);
and U29270 (N_29270,N_15132,N_16666);
and U29271 (N_29271,N_11009,N_14820);
xnor U29272 (N_29272,N_17539,N_12886);
nor U29273 (N_29273,N_12934,N_18253);
or U29274 (N_29274,N_12641,N_11027);
xor U29275 (N_29275,N_13682,N_15380);
or U29276 (N_29276,N_11321,N_13939);
nor U29277 (N_29277,N_14210,N_13139);
nand U29278 (N_29278,N_17959,N_19533);
nor U29279 (N_29279,N_10139,N_14604);
nand U29280 (N_29280,N_12495,N_18460);
or U29281 (N_29281,N_18260,N_11559);
nand U29282 (N_29282,N_13588,N_15271);
nand U29283 (N_29283,N_17677,N_17784);
xor U29284 (N_29284,N_14221,N_17585);
nand U29285 (N_29285,N_19410,N_15859);
nor U29286 (N_29286,N_16297,N_10433);
nor U29287 (N_29287,N_13050,N_12621);
nor U29288 (N_29288,N_11505,N_12859);
and U29289 (N_29289,N_16509,N_13115);
nand U29290 (N_29290,N_15050,N_10401);
nor U29291 (N_29291,N_13997,N_13325);
and U29292 (N_29292,N_17908,N_13668);
and U29293 (N_29293,N_17506,N_14879);
or U29294 (N_29294,N_18423,N_14834);
nor U29295 (N_29295,N_17698,N_12590);
xnor U29296 (N_29296,N_10502,N_15206);
and U29297 (N_29297,N_19294,N_19157);
nor U29298 (N_29298,N_10026,N_17320);
nor U29299 (N_29299,N_16257,N_10068);
xor U29300 (N_29300,N_17182,N_16467);
or U29301 (N_29301,N_14996,N_10931);
and U29302 (N_29302,N_15902,N_10980);
nand U29303 (N_29303,N_19138,N_10556);
and U29304 (N_29304,N_16675,N_13819);
nand U29305 (N_29305,N_17353,N_16675);
nand U29306 (N_29306,N_15609,N_14442);
or U29307 (N_29307,N_17296,N_18313);
nor U29308 (N_29308,N_14065,N_13741);
nor U29309 (N_29309,N_13124,N_15819);
and U29310 (N_29310,N_12199,N_18886);
nor U29311 (N_29311,N_14596,N_17945);
and U29312 (N_29312,N_16743,N_16184);
nand U29313 (N_29313,N_10963,N_16506);
and U29314 (N_29314,N_14517,N_17216);
or U29315 (N_29315,N_16655,N_11993);
nand U29316 (N_29316,N_11246,N_11994);
and U29317 (N_29317,N_12219,N_19104);
nand U29318 (N_29318,N_11917,N_18475);
and U29319 (N_29319,N_11326,N_13518);
nor U29320 (N_29320,N_16945,N_15388);
nand U29321 (N_29321,N_18783,N_16163);
nand U29322 (N_29322,N_12415,N_16738);
nor U29323 (N_29323,N_11331,N_13900);
xnor U29324 (N_29324,N_17946,N_19381);
nand U29325 (N_29325,N_13286,N_17248);
nor U29326 (N_29326,N_16672,N_11884);
or U29327 (N_29327,N_16352,N_15881);
or U29328 (N_29328,N_19124,N_19164);
or U29329 (N_29329,N_18972,N_10415);
or U29330 (N_29330,N_10738,N_15223);
or U29331 (N_29331,N_12065,N_15596);
nor U29332 (N_29332,N_19941,N_12054);
or U29333 (N_29333,N_10121,N_19871);
or U29334 (N_29334,N_15837,N_17866);
or U29335 (N_29335,N_19524,N_13212);
or U29336 (N_29336,N_12417,N_18865);
xor U29337 (N_29337,N_14043,N_17726);
or U29338 (N_29338,N_13964,N_12106);
and U29339 (N_29339,N_16647,N_11600);
xor U29340 (N_29340,N_17188,N_12096);
or U29341 (N_29341,N_11600,N_11624);
and U29342 (N_29342,N_17205,N_10640);
and U29343 (N_29343,N_16759,N_14058);
xnor U29344 (N_29344,N_13922,N_18554);
nor U29345 (N_29345,N_16305,N_17781);
and U29346 (N_29346,N_14296,N_16476);
or U29347 (N_29347,N_18549,N_13640);
nand U29348 (N_29348,N_11546,N_14220);
and U29349 (N_29349,N_15893,N_15773);
nand U29350 (N_29350,N_17635,N_15397);
nand U29351 (N_29351,N_11850,N_15079);
nand U29352 (N_29352,N_14403,N_12054);
nand U29353 (N_29353,N_18052,N_15605);
or U29354 (N_29354,N_11425,N_10796);
nor U29355 (N_29355,N_12808,N_19403);
nor U29356 (N_29356,N_17150,N_10149);
nand U29357 (N_29357,N_16329,N_18649);
or U29358 (N_29358,N_10444,N_15019);
or U29359 (N_29359,N_12589,N_17750);
or U29360 (N_29360,N_18795,N_13084);
nand U29361 (N_29361,N_13442,N_13458);
or U29362 (N_29362,N_11405,N_14342);
and U29363 (N_29363,N_10106,N_19631);
and U29364 (N_29364,N_16767,N_19238);
and U29365 (N_29365,N_14863,N_11917);
nand U29366 (N_29366,N_13391,N_16102);
or U29367 (N_29367,N_10826,N_18598);
and U29368 (N_29368,N_15775,N_15970);
and U29369 (N_29369,N_15625,N_17177);
or U29370 (N_29370,N_18524,N_17578);
xnor U29371 (N_29371,N_10509,N_10435);
and U29372 (N_29372,N_15462,N_17052);
nor U29373 (N_29373,N_19229,N_17382);
nor U29374 (N_29374,N_16182,N_12637);
xor U29375 (N_29375,N_13107,N_10986);
and U29376 (N_29376,N_13578,N_18780);
and U29377 (N_29377,N_11990,N_11834);
nand U29378 (N_29378,N_15425,N_15399);
or U29379 (N_29379,N_14344,N_19351);
nor U29380 (N_29380,N_19861,N_13895);
or U29381 (N_29381,N_17096,N_11438);
xor U29382 (N_29382,N_14074,N_17991);
nand U29383 (N_29383,N_14937,N_17058);
or U29384 (N_29384,N_10865,N_12710);
and U29385 (N_29385,N_14104,N_16744);
or U29386 (N_29386,N_15459,N_12403);
nand U29387 (N_29387,N_18819,N_18824);
and U29388 (N_29388,N_10072,N_18930);
and U29389 (N_29389,N_10505,N_16568);
nand U29390 (N_29390,N_14387,N_13370);
nand U29391 (N_29391,N_19686,N_12033);
and U29392 (N_29392,N_13920,N_16366);
nor U29393 (N_29393,N_11975,N_18430);
nand U29394 (N_29394,N_17253,N_12450);
nand U29395 (N_29395,N_13359,N_15553);
or U29396 (N_29396,N_18802,N_16776);
nand U29397 (N_29397,N_19919,N_11089);
nand U29398 (N_29398,N_11752,N_11346);
nand U29399 (N_29399,N_12657,N_16750);
and U29400 (N_29400,N_12128,N_15457);
nand U29401 (N_29401,N_10591,N_16747);
and U29402 (N_29402,N_10976,N_13364);
and U29403 (N_29403,N_13574,N_14144);
or U29404 (N_29404,N_13416,N_12148);
xnor U29405 (N_29405,N_14276,N_14364);
xnor U29406 (N_29406,N_15772,N_15544);
or U29407 (N_29407,N_11380,N_18078);
nand U29408 (N_29408,N_14856,N_17737);
or U29409 (N_29409,N_15069,N_12462);
nor U29410 (N_29410,N_16674,N_10386);
and U29411 (N_29411,N_10060,N_18454);
nor U29412 (N_29412,N_12458,N_16491);
xnor U29413 (N_29413,N_15978,N_13378);
nand U29414 (N_29414,N_11384,N_15889);
nor U29415 (N_29415,N_13923,N_14962);
xnor U29416 (N_29416,N_12380,N_13880);
nor U29417 (N_29417,N_13057,N_11501);
and U29418 (N_29418,N_16093,N_11532);
xnor U29419 (N_29419,N_15111,N_13813);
nand U29420 (N_29420,N_16084,N_13176);
or U29421 (N_29421,N_17690,N_12943);
and U29422 (N_29422,N_14092,N_18922);
and U29423 (N_29423,N_14610,N_11247);
nand U29424 (N_29424,N_14912,N_14753);
and U29425 (N_29425,N_13906,N_19343);
nor U29426 (N_29426,N_18132,N_10232);
nor U29427 (N_29427,N_17331,N_15243);
and U29428 (N_29428,N_10880,N_18223);
nand U29429 (N_29429,N_14648,N_10900);
xnor U29430 (N_29430,N_10701,N_10189);
and U29431 (N_29431,N_15618,N_15497);
or U29432 (N_29432,N_10474,N_14413);
or U29433 (N_29433,N_12960,N_13910);
or U29434 (N_29434,N_10519,N_11439);
or U29435 (N_29435,N_11112,N_19387);
and U29436 (N_29436,N_18039,N_18576);
nand U29437 (N_29437,N_16988,N_16699);
nand U29438 (N_29438,N_17883,N_13471);
nor U29439 (N_29439,N_13807,N_13117);
or U29440 (N_29440,N_15390,N_11352);
xnor U29441 (N_29441,N_10164,N_11523);
or U29442 (N_29442,N_11192,N_18204);
xnor U29443 (N_29443,N_10827,N_17144);
and U29444 (N_29444,N_14758,N_19151);
and U29445 (N_29445,N_11973,N_18800);
or U29446 (N_29446,N_13867,N_13923);
nand U29447 (N_29447,N_18867,N_14675);
or U29448 (N_29448,N_11822,N_17444);
nand U29449 (N_29449,N_15972,N_11103);
nor U29450 (N_29450,N_13283,N_13352);
xor U29451 (N_29451,N_13084,N_17054);
and U29452 (N_29452,N_15149,N_17105);
or U29453 (N_29453,N_10135,N_15763);
xor U29454 (N_29454,N_15158,N_16499);
or U29455 (N_29455,N_14480,N_13778);
or U29456 (N_29456,N_18493,N_12786);
nand U29457 (N_29457,N_16562,N_19188);
and U29458 (N_29458,N_14048,N_16131);
xor U29459 (N_29459,N_18576,N_10975);
nor U29460 (N_29460,N_12043,N_14443);
or U29461 (N_29461,N_14268,N_14851);
xor U29462 (N_29462,N_10345,N_15412);
or U29463 (N_29463,N_12536,N_18627);
nand U29464 (N_29464,N_19808,N_13533);
and U29465 (N_29465,N_17495,N_13013);
nand U29466 (N_29466,N_16354,N_12765);
or U29467 (N_29467,N_15050,N_10820);
nor U29468 (N_29468,N_14849,N_15959);
and U29469 (N_29469,N_10803,N_14155);
nand U29470 (N_29470,N_18093,N_15298);
and U29471 (N_29471,N_10186,N_11209);
or U29472 (N_29472,N_12507,N_16867);
xnor U29473 (N_29473,N_18290,N_13835);
and U29474 (N_29474,N_19588,N_14604);
nand U29475 (N_29475,N_19100,N_17994);
nand U29476 (N_29476,N_12364,N_15381);
nor U29477 (N_29477,N_19189,N_15775);
nand U29478 (N_29478,N_14171,N_18440);
nand U29479 (N_29479,N_10569,N_17226);
nor U29480 (N_29480,N_11225,N_11058);
nand U29481 (N_29481,N_10352,N_14707);
or U29482 (N_29482,N_19923,N_18083);
or U29483 (N_29483,N_14517,N_12987);
or U29484 (N_29484,N_18699,N_18144);
nand U29485 (N_29485,N_11047,N_17120);
nand U29486 (N_29486,N_11282,N_12658);
nand U29487 (N_29487,N_10116,N_12207);
nor U29488 (N_29488,N_14951,N_18341);
nor U29489 (N_29489,N_13293,N_16621);
nor U29490 (N_29490,N_13960,N_11908);
nor U29491 (N_29491,N_13959,N_10575);
nor U29492 (N_29492,N_16052,N_17609);
nand U29493 (N_29493,N_12078,N_14057);
nand U29494 (N_29494,N_16174,N_15182);
nand U29495 (N_29495,N_11037,N_17008);
nand U29496 (N_29496,N_18489,N_10702);
or U29497 (N_29497,N_10106,N_11387);
and U29498 (N_29498,N_14891,N_14306);
xor U29499 (N_29499,N_12052,N_14579);
xor U29500 (N_29500,N_16473,N_18814);
and U29501 (N_29501,N_18703,N_13933);
and U29502 (N_29502,N_19938,N_17734);
nand U29503 (N_29503,N_19165,N_18777);
or U29504 (N_29504,N_12595,N_19226);
and U29505 (N_29505,N_19124,N_15841);
or U29506 (N_29506,N_12911,N_12238);
or U29507 (N_29507,N_14097,N_15078);
and U29508 (N_29508,N_11627,N_15157);
and U29509 (N_29509,N_19836,N_17057);
and U29510 (N_29510,N_11683,N_10940);
nand U29511 (N_29511,N_12829,N_19568);
or U29512 (N_29512,N_11907,N_15950);
and U29513 (N_29513,N_11235,N_15244);
or U29514 (N_29514,N_16845,N_10347);
or U29515 (N_29515,N_13862,N_17226);
nor U29516 (N_29516,N_16771,N_18981);
and U29517 (N_29517,N_15182,N_15977);
nor U29518 (N_29518,N_18198,N_12949);
nor U29519 (N_29519,N_17959,N_15756);
and U29520 (N_29520,N_14904,N_12389);
nor U29521 (N_29521,N_17523,N_12390);
nand U29522 (N_29522,N_16150,N_13248);
or U29523 (N_29523,N_10174,N_10313);
nand U29524 (N_29524,N_15944,N_15966);
or U29525 (N_29525,N_17878,N_15074);
nor U29526 (N_29526,N_12195,N_17456);
nor U29527 (N_29527,N_18540,N_11974);
nor U29528 (N_29528,N_11216,N_17832);
or U29529 (N_29529,N_12222,N_16776);
xor U29530 (N_29530,N_17933,N_13114);
and U29531 (N_29531,N_14731,N_11933);
or U29532 (N_29532,N_17456,N_13869);
nor U29533 (N_29533,N_19665,N_14677);
or U29534 (N_29534,N_15167,N_11025);
nor U29535 (N_29535,N_11485,N_12562);
and U29536 (N_29536,N_12806,N_11932);
nand U29537 (N_29537,N_11471,N_10426);
and U29538 (N_29538,N_16483,N_15462);
nor U29539 (N_29539,N_15016,N_15361);
nand U29540 (N_29540,N_17791,N_16299);
and U29541 (N_29541,N_11820,N_14636);
or U29542 (N_29542,N_11015,N_19324);
and U29543 (N_29543,N_12568,N_10461);
or U29544 (N_29544,N_19103,N_17592);
and U29545 (N_29545,N_17092,N_11322);
and U29546 (N_29546,N_11341,N_13953);
xor U29547 (N_29547,N_17103,N_15537);
nor U29548 (N_29548,N_13730,N_10885);
nand U29549 (N_29549,N_10881,N_10313);
nand U29550 (N_29550,N_15575,N_19178);
or U29551 (N_29551,N_12046,N_13527);
xnor U29552 (N_29552,N_18884,N_13363);
and U29553 (N_29553,N_10202,N_12308);
nand U29554 (N_29554,N_10060,N_11538);
or U29555 (N_29555,N_15090,N_18489);
nor U29556 (N_29556,N_15511,N_11398);
xnor U29557 (N_29557,N_10815,N_14568);
and U29558 (N_29558,N_12404,N_10828);
nand U29559 (N_29559,N_11101,N_19898);
nand U29560 (N_29560,N_10455,N_19627);
xnor U29561 (N_29561,N_17816,N_10022);
nor U29562 (N_29562,N_19989,N_13636);
or U29563 (N_29563,N_19149,N_10756);
or U29564 (N_29564,N_16826,N_10292);
xor U29565 (N_29565,N_10832,N_16081);
nor U29566 (N_29566,N_17859,N_18098);
nand U29567 (N_29567,N_14144,N_14984);
xnor U29568 (N_29568,N_10155,N_10822);
xnor U29569 (N_29569,N_14224,N_16837);
xor U29570 (N_29570,N_11422,N_15775);
and U29571 (N_29571,N_13341,N_13879);
or U29572 (N_29572,N_12100,N_13866);
nand U29573 (N_29573,N_10840,N_14182);
and U29574 (N_29574,N_12715,N_15241);
nand U29575 (N_29575,N_10963,N_16832);
nand U29576 (N_29576,N_12421,N_11080);
or U29577 (N_29577,N_13728,N_17828);
and U29578 (N_29578,N_18956,N_18087);
or U29579 (N_29579,N_12296,N_14736);
nor U29580 (N_29580,N_18803,N_13732);
and U29581 (N_29581,N_16252,N_10558);
nand U29582 (N_29582,N_17631,N_16430);
or U29583 (N_29583,N_15634,N_18252);
or U29584 (N_29584,N_17201,N_16944);
and U29585 (N_29585,N_11402,N_14051);
xnor U29586 (N_29586,N_12380,N_18822);
nor U29587 (N_29587,N_17288,N_10394);
nand U29588 (N_29588,N_10990,N_19113);
and U29589 (N_29589,N_17689,N_14756);
nand U29590 (N_29590,N_15026,N_12570);
nor U29591 (N_29591,N_16111,N_12230);
nand U29592 (N_29592,N_17775,N_16653);
nand U29593 (N_29593,N_18760,N_16933);
nor U29594 (N_29594,N_10733,N_14156);
nand U29595 (N_29595,N_10169,N_10019);
and U29596 (N_29596,N_14331,N_18796);
xor U29597 (N_29597,N_15585,N_13771);
and U29598 (N_29598,N_14236,N_14598);
and U29599 (N_29599,N_11757,N_19590);
xor U29600 (N_29600,N_18350,N_14546);
nand U29601 (N_29601,N_12456,N_17970);
xor U29602 (N_29602,N_11849,N_16384);
xnor U29603 (N_29603,N_16332,N_18825);
and U29604 (N_29604,N_14366,N_17970);
xor U29605 (N_29605,N_12360,N_16510);
or U29606 (N_29606,N_19221,N_13406);
nand U29607 (N_29607,N_11136,N_11554);
nand U29608 (N_29608,N_11113,N_15520);
and U29609 (N_29609,N_11278,N_11364);
nor U29610 (N_29610,N_11118,N_15700);
nand U29611 (N_29611,N_13705,N_13448);
or U29612 (N_29612,N_17761,N_11990);
or U29613 (N_29613,N_11303,N_15179);
nand U29614 (N_29614,N_19753,N_10268);
nand U29615 (N_29615,N_15644,N_18450);
xnor U29616 (N_29616,N_13972,N_18937);
or U29617 (N_29617,N_16805,N_11186);
xnor U29618 (N_29618,N_10779,N_19980);
nor U29619 (N_29619,N_15370,N_16382);
and U29620 (N_29620,N_10305,N_14180);
or U29621 (N_29621,N_17318,N_17387);
or U29622 (N_29622,N_17514,N_16942);
or U29623 (N_29623,N_19591,N_10988);
and U29624 (N_29624,N_15832,N_11726);
nand U29625 (N_29625,N_13271,N_13951);
xnor U29626 (N_29626,N_18333,N_11723);
or U29627 (N_29627,N_15681,N_18407);
and U29628 (N_29628,N_18878,N_15047);
xor U29629 (N_29629,N_17969,N_14721);
and U29630 (N_29630,N_15999,N_14805);
or U29631 (N_29631,N_10286,N_14662);
nor U29632 (N_29632,N_14752,N_13185);
or U29633 (N_29633,N_14692,N_14212);
or U29634 (N_29634,N_18364,N_19675);
or U29635 (N_29635,N_15706,N_12682);
nor U29636 (N_29636,N_12858,N_16375);
and U29637 (N_29637,N_13399,N_12913);
nand U29638 (N_29638,N_14093,N_12511);
nand U29639 (N_29639,N_17498,N_12837);
and U29640 (N_29640,N_15566,N_11062);
xnor U29641 (N_29641,N_10610,N_10627);
and U29642 (N_29642,N_10121,N_12751);
nand U29643 (N_29643,N_14435,N_10592);
or U29644 (N_29644,N_19947,N_10366);
nor U29645 (N_29645,N_12632,N_12369);
nor U29646 (N_29646,N_11027,N_15796);
and U29647 (N_29647,N_19455,N_14293);
nand U29648 (N_29648,N_17462,N_14046);
or U29649 (N_29649,N_16735,N_12067);
and U29650 (N_29650,N_16606,N_13841);
nand U29651 (N_29651,N_13669,N_11924);
or U29652 (N_29652,N_17946,N_17743);
nor U29653 (N_29653,N_12054,N_12381);
and U29654 (N_29654,N_18823,N_10720);
nand U29655 (N_29655,N_11112,N_11558);
and U29656 (N_29656,N_19929,N_10922);
and U29657 (N_29657,N_14740,N_10579);
nand U29658 (N_29658,N_14386,N_11022);
nor U29659 (N_29659,N_14505,N_10409);
nand U29660 (N_29660,N_15763,N_11216);
nor U29661 (N_29661,N_16651,N_12037);
nor U29662 (N_29662,N_17973,N_12445);
or U29663 (N_29663,N_16684,N_11647);
or U29664 (N_29664,N_13261,N_10355);
and U29665 (N_29665,N_13688,N_16970);
nor U29666 (N_29666,N_13659,N_19972);
and U29667 (N_29667,N_11408,N_14667);
or U29668 (N_29668,N_13611,N_11914);
and U29669 (N_29669,N_19344,N_17129);
and U29670 (N_29670,N_19095,N_14368);
and U29671 (N_29671,N_17906,N_18136);
nand U29672 (N_29672,N_19943,N_14094);
and U29673 (N_29673,N_13691,N_11543);
or U29674 (N_29674,N_10075,N_11599);
nor U29675 (N_29675,N_12618,N_13561);
xor U29676 (N_29676,N_12868,N_19913);
or U29677 (N_29677,N_18169,N_19303);
xnor U29678 (N_29678,N_13313,N_14698);
nand U29679 (N_29679,N_12517,N_19531);
or U29680 (N_29680,N_16839,N_10918);
and U29681 (N_29681,N_17612,N_14568);
or U29682 (N_29682,N_10399,N_13251);
nor U29683 (N_29683,N_18512,N_16973);
nor U29684 (N_29684,N_15128,N_12664);
and U29685 (N_29685,N_14286,N_14182);
xor U29686 (N_29686,N_13827,N_18248);
and U29687 (N_29687,N_17560,N_18247);
and U29688 (N_29688,N_14921,N_16843);
xnor U29689 (N_29689,N_13283,N_19872);
xor U29690 (N_29690,N_13056,N_11168);
and U29691 (N_29691,N_11630,N_19982);
and U29692 (N_29692,N_19856,N_15069);
nand U29693 (N_29693,N_14212,N_13756);
and U29694 (N_29694,N_19485,N_16946);
and U29695 (N_29695,N_16849,N_12634);
and U29696 (N_29696,N_10661,N_12473);
nor U29697 (N_29697,N_11710,N_13694);
or U29698 (N_29698,N_19031,N_11681);
or U29699 (N_29699,N_16131,N_12011);
nor U29700 (N_29700,N_14974,N_14207);
and U29701 (N_29701,N_13913,N_16317);
nor U29702 (N_29702,N_15212,N_15609);
nand U29703 (N_29703,N_14877,N_19549);
xor U29704 (N_29704,N_14550,N_15949);
nor U29705 (N_29705,N_12754,N_13183);
or U29706 (N_29706,N_10071,N_15928);
nor U29707 (N_29707,N_12633,N_18003);
nand U29708 (N_29708,N_10506,N_12607);
and U29709 (N_29709,N_12608,N_14296);
or U29710 (N_29710,N_14149,N_11490);
nand U29711 (N_29711,N_19138,N_10581);
or U29712 (N_29712,N_18885,N_10341);
or U29713 (N_29713,N_19253,N_10801);
nor U29714 (N_29714,N_13312,N_14602);
nand U29715 (N_29715,N_16974,N_13733);
nand U29716 (N_29716,N_18651,N_10331);
or U29717 (N_29717,N_16027,N_15987);
xor U29718 (N_29718,N_14462,N_11848);
or U29719 (N_29719,N_18399,N_16999);
nor U29720 (N_29720,N_12116,N_17346);
and U29721 (N_29721,N_14239,N_17157);
nor U29722 (N_29722,N_18154,N_13042);
and U29723 (N_29723,N_16062,N_16405);
xor U29724 (N_29724,N_11798,N_17086);
xnor U29725 (N_29725,N_16052,N_13126);
nor U29726 (N_29726,N_14293,N_13844);
or U29727 (N_29727,N_17890,N_15958);
or U29728 (N_29728,N_19297,N_15638);
and U29729 (N_29729,N_13453,N_11572);
or U29730 (N_29730,N_11729,N_15487);
nand U29731 (N_29731,N_10771,N_15451);
nand U29732 (N_29732,N_16375,N_16387);
or U29733 (N_29733,N_19770,N_11915);
or U29734 (N_29734,N_14129,N_11108);
and U29735 (N_29735,N_13713,N_12638);
xnor U29736 (N_29736,N_12710,N_17542);
nor U29737 (N_29737,N_17716,N_16470);
nor U29738 (N_29738,N_18635,N_19633);
and U29739 (N_29739,N_18655,N_11602);
nand U29740 (N_29740,N_15766,N_17968);
nand U29741 (N_29741,N_18944,N_19353);
nor U29742 (N_29742,N_17292,N_16026);
nand U29743 (N_29743,N_19834,N_12875);
nand U29744 (N_29744,N_17328,N_13110);
and U29745 (N_29745,N_10102,N_18137);
and U29746 (N_29746,N_16462,N_14548);
nor U29747 (N_29747,N_11439,N_17372);
nor U29748 (N_29748,N_19429,N_15133);
or U29749 (N_29749,N_13487,N_15637);
nand U29750 (N_29750,N_12805,N_11729);
nor U29751 (N_29751,N_16462,N_14647);
or U29752 (N_29752,N_18515,N_19605);
nor U29753 (N_29753,N_17455,N_14092);
nand U29754 (N_29754,N_18451,N_15713);
xor U29755 (N_29755,N_14733,N_17967);
and U29756 (N_29756,N_19098,N_19141);
xnor U29757 (N_29757,N_10758,N_14375);
or U29758 (N_29758,N_13126,N_16133);
nand U29759 (N_29759,N_14207,N_17544);
nand U29760 (N_29760,N_17513,N_19570);
or U29761 (N_29761,N_13172,N_15672);
and U29762 (N_29762,N_19942,N_11410);
nand U29763 (N_29763,N_12538,N_19049);
and U29764 (N_29764,N_14871,N_12588);
nor U29765 (N_29765,N_15669,N_13363);
or U29766 (N_29766,N_14231,N_13844);
nand U29767 (N_29767,N_17547,N_12764);
and U29768 (N_29768,N_15842,N_18885);
and U29769 (N_29769,N_11060,N_17045);
nand U29770 (N_29770,N_10435,N_11973);
and U29771 (N_29771,N_13602,N_16413);
and U29772 (N_29772,N_10981,N_10108);
and U29773 (N_29773,N_12838,N_11200);
or U29774 (N_29774,N_10198,N_11257);
nand U29775 (N_29775,N_13750,N_19573);
or U29776 (N_29776,N_17769,N_11552);
nand U29777 (N_29777,N_13266,N_13975);
nor U29778 (N_29778,N_10635,N_19986);
and U29779 (N_29779,N_15818,N_15718);
or U29780 (N_29780,N_13571,N_15972);
nand U29781 (N_29781,N_12985,N_12672);
nor U29782 (N_29782,N_16669,N_18217);
xnor U29783 (N_29783,N_11834,N_12918);
or U29784 (N_29784,N_10592,N_15765);
or U29785 (N_29785,N_10311,N_18582);
nor U29786 (N_29786,N_18425,N_19128);
nor U29787 (N_29787,N_12279,N_16772);
nand U29788 (N_29788,N_19754,N_11016);
or U29789 (N_29789,N_16584,N_14349);
and U29790 (N_29790,N_14520,N_19070);
nor U29791 (N_29791,N_14969,N_13473);
nor U29792 (N_29792,N_11582,N_14709);
nor U29793 (N_29793,N_11952,N_16376);
nor U29794 (N_29794,N_12255,N_17464);
and U29795 (N_29795,N_18758,N_17165);
xnor U29796 (N_29796,N_19510,N_12223);
nand U29797 (N_29797,N_19067,N_19667);
nand U29798 (N_29798,N_10780,N_16891);
or U29799 (N_29799,N_12186,N_17135);
nand U29800 (N_29800,N_14674,N_19546);
nand U29801 (N_29801,N_14248,N_14970);
or U29802 (N_29802,N_17212,N_18367);
and U29803 (N_29803,N_12205,N_15726);
xnor U29804 (N_29804,N_13463,N_17708);
nor U29805 (N_29805,N_12134,N_19980);
xor U29806 (N_29806,N_16112,N_15869);
nor U29807 (N_29807,N_13313,N_10455);
or U29808 (N_29808,N_17665,N_10325);
xor U29809 (N_29809,N_17435,N_17579);
and U29810 (N_29810,N_18334,N_16174);
and U29811 (N_29811,N_10648,N_14053);
nand U29812 (N_29812,N_11934,N_17426);
nand U29813 (N_29813,N_12237,N_16593);
nand U29814 (N_29814,N_14872,N_17676);
nand U29815 (N_29815,N_15955,N_18732);
nor U29816 (N_29816,N_10281,N_12482);
nor U29817 (N_29817,N_18416,N_18230);
xnor U29818 (N_29818,N_11873,N_16730);
or U29819 (N_29819,N_17863,N_17879);
and U29820 (N_29820,N_10694,N_11841);
nand U29821 (N_29821,N_14522,N_19428);
or U29822 (N_29822,N_17903,N_11669);
or U29823 (N_29823,N_17358,N_13753);
xor U29824 (N_29824,N_18356,N_13156);
or U29825 (N_29825,N_10047,N_18195);
and U29826 (N_29826,N_17769,N_17958);
nor U29827 (N_29827,N_16745,N_10271);
nand U29828 (N_29828,N_12214,N_16605);
xnor U29829 (N_29829,N_13399,N_13425);
nand U29830 (N_29830,N_17420,N_13259);
and U29831 (N_29831,N_17306,N_10742);
or U29832 (N_29832,N_13368,N_19048);
and U29833 (N_29833,N_19216,N_17123);
and U29834 (N_29834,N_12652,N_15407);
nand U29835 (N_29835,N_10402,N_14750);
and U29836 (N_29836,N_18133,N_18104);
nand U29837 (N_29837,N_18638,N_19690);
or U29838 (N_29838,N_17915,N_12694);
or U29839 (N_29839,N_12429,N_16123);
or U29840 (N_29840,N_10747,N_15828);
or U29841 (N_29841,N_14023,N_19482);
nand U29842 (N_29842,N_17441,N_18089);
nand U29843 (N_29843,N_16639,N_15889);
nand U29844 (N_29844,N_10707,N_13864);
nand U29845 (N_29845,N_16789,N_14953);
or U29846 (N_29846,N_15661,N_11531);
or U29847 (N_29847,N_17164,N_14749);
and U29848 (N_29848,N_10147,N_15938);
nand U29849 (N_29849,N_12627,N_16400);
nand U29850 (N_29850,N_14836,N_12149);
nand U29851 (N_29851,N_19653,N_14838);
nand U29852 (N_29852,N_13254,N_19738);
nor U29853 (N_29853,N_10326,N_17385);
nor U29854 (N_29854,N_13792,N_15258);
and U29855 (N_29855,N_19679,N_16107);
nand U29856 (N_29856,N_16657,N_10609);
or U29857 (N_29857,N_14042,N_10523);
nor U29858 (N_29858,N_12675,N_19200);
xor U29859 (N_29859,N_14383,N_14791);
nor U29860 (N_29860,N_16241,N_11176);
and U29861 (N_29861,N_18105,N_18059);
nand U29862 (N_29862,N_18911,N_16451);
and U29863 (N_29863,N_10842,N_14399);
and U29864 (N_29864,N_18763,N_14034);
xnor U29865 (N_29865,N_17196,N_10829);
nor U29866 (N_29866,N_13343,N_13311);
and U29867 (N_29867,N_15135,N_13771);
nand U29868 (N_29868,N_12063,N_16658);
nand U29869 (N_29869,N_16435,N_14877);
nor U29870 (N_29870,N_11449,N_14125);
or U29871 (N_29871,N_11832,N_18099);
nand U29872 (N_29872,N_14428,N_10895);
and U29873 (N_29873,N_18776,N_15293);
nand U29874 (N_29874,N_19159,N_19926);
xor U29875 (N_29875,N_19316,N_18931);
nand U29876 (N_29876,N_19681,N_13473);
nor U29877 (N_29877,N_10737,N_12273);
xnor U29878 (N_29878,N_13810,N_19656);
and U29879 (N_29879,N_10471,N_17535);
nand U29880 (N_29880,N_10448,N_18755);
nor U29881 (N_29881,N_16031,N_16252);
or U29882 (N_29882,N_15790,N_19746);
xor U29883 (N_29883,N_17889,N_11558);
and U29884 (N_29884,N_16792,N_13283);
nand U29885 (N_29885,N_12958,N_18752);
nand U29886 (N_29886,N_18296,N_19195);
nor U29887 (N_29887,N_15888,N_11077);
nor U29888 (N_29888,N_13564,N_15304);
and U29889 (N_29889,N_14516,N_16936);
nand U29890 (N_29890,N_18489,N_12458);
nand U29891 (N_29891,N_10263,N_12956);
nand U29892 (N_29892,N_18625,N_19237);
nand U29893 (N_29893,N_13276,N_17846);
xnor U29894 (N_29894,N_12043,N_17070);
and U29895 (N_29895,N_15686,N_12109);
or U29896 (N_29896,N_11084,N_12092);
nand U29897 (N_29897,N_11489,N_14567);
and U29898 (N_29898,N_10954,N_14251);
or U29899 (N_29899,N_10207,N_15237);
and U29900 (N_29900,N_19274,N_19824);
or U29901 (N_29901,N_10221,N_15294);
nand U29902 (N_29902,N_13930,N_11036);
and U29903 (N_29903,N_11163,N_19432);
nor U29904 (N_29904,N_14142,N_13186);
nand U29905 (N_29905,N_13060,N_14599);
nor U29906 (N_29906,N_12825,N_16596);
xor U29907 (N_29907,N_18727,N_10911);
or U29908 (N_29908,N_18391,N_11650);
or U29909 (N_29909,N_11428,N_15283);
xor U29910 (N_29910,N_17820,N_14270);
nor U29911 (N_29911,N_15554,N_19253);
nor U29912 (N_29912,N_10706,N_14882);
xor U29913 (N_29913,N_14445,N_14878);
nand U29914 (N_29914,N_11247,N_12516);
nand U29915 (N_29915,N_14085,N_14059);
xor U29916 (N_29916,N_18632,N_11588);
xnor U29917 (N_29917,N_14498,N_19384);
and U29918 (N_29918,N_13062,N_16875);
or U29919 (N_29919,N_12030,N_10870);
nand U29920 (N_29920,N_10723,N_14015);
and U29921 (N_29921,N_19813,N_17612);
xnor U29922 (N_29922,N_13496,N_14648);
and U29923 (N_29923,N_16009,N_18023);
and U29924 (N_29924,N_16177,N_17216);
and U29925 (N_29925,N_19546,N_19360);
xor U29926 (N_29926,N_15807,N_13846);
and U29927 (N_29927,N_18133,N_19795);
nor U29928 (N_29928,N_12461,N_17257);
and U29929 (N_29929,N_10347,N_13659);
nand U29930 (N_29930,N_12770,N_11556);
nand U29931 (N_29931,N_16044,N_13724);
or U29932 (N_29932,N_16894,N_11481);
or U29933 (N_29933,N_12932,N_11093);
nand U29934 (N_29934,N_14824,N_11922);
nand U29935 (N_29935,N_13107,N_11553);
xnor U29936 (N_29936,N_14661,N_17237);
nand U29937 (N_29937,N_15006,N_13666);
or U29938 (N_29938,N_15498,N_17236);
nand U29939 (N_29939,N_19711,N_19992);
and U29940 (N_29940,N_16704,N_16468);
or U29941 (N_29941,N_12697,N_12220);
nor U29942 (N_29942,N_19860,N_14812);
and U29943 (N_29943,N_18644,N_10921);
nor U29944 (N_29944,N_12246,N_18891);
xor U29945 (N_29945,N_13478,N_18900);
or U29946 (N_29946,N_10073,N_11423);
nor U29947 (N_29947,N_18381,N_18459);
or U29948 (N_29948,N_14271,N_16832);
and U29949 (N_29949,N_16634,N_12484);
xor U29950 (N_29950,N_19409,N_13268);
nand U29951 (N_29951,N_17420,N_13207);
or U29952 (N_29952,N_13496,N_14441);
and U29953 (N_29953,N_14322,N_13582);
nand U29954 (N_29954,N_13386,N_16227);
xor U29955 (N_29955,N_11085,N_18586);
or U29956 (N_29956,N_18490,N_13912);
nor U29957 (N_29957,N_14821,N_13127);
xnor U29958 (N_29958,N_19161,N_18437);
or U29959 (N_29959,N_19434,N_19423);
nor U29960 (N_29960,N_19896,N_11665);
or U29961 (N_29961,N_11866,N_11788);
nor U29962 (N_29962,N_11659,N_11614);
nand U29963 (N_29963,N_11343,N_10537);
and U29964 (N_29964,N_13499,N_18757);
nand U29965 (N_29965,N_10939,N_18244);
and U29966 (N_29966,N_18057,N_15665);
nor U29967 (N_29967,N_15037,N_15541);
or U29968 (N_29968,N_13352,N_17743);
or U29969 (N_29969,N_15975,N_13200);
and U29970 (N_29970,N_13800,N_16151);
or U29971 (N_29971,N_19535,N_17824);
xnor U29972 (N_29972,N_15371,N_14065);
nor U29973 (N_29973,N_16558,N_17353);
nor U29974 (N_29974,N_15516,N_15833);
and U29975 (N_29975,N_17187,N_17729);
nor U29976 (N_29976,N_11860,N_16871);
and U29977 (N_29977,N_18580,N_10435);
nand U29978 (N_29978,N_19052,N_15672);
and U29979 (N_29979,N_14867,N_14681);
and U29980 (N_29980,N_17030,N_10965);
and U29981 (N_29981,N_13586,N_15133);
nor U29982 (N_29982,N_17856,N_16313);
nor U29983 (N_29983,N_15679,N_14385);
and U29984 (N_29984,N_19631,N_10381);
nor U29985 (N_29985,N_17813,N_11475);
and U29986 (N_29986,N_10686,N_10651);
or U29987 (N_29987,N_18984,N_12570);
and U29988 (N_29988,N_12728,N_17551);
nor U29989 (N_29989,N_17993,N_16926);
nor U29990 (N_29990,N_14980,N_12144);
nor U29991 (N_29991,N_19465,N_10552);
nor U29992 (N_29992,N_15498,N_18160);
nand U29993 (N_29993,N_16991,N_15570);
xnor U29994 (N_29994,N_18784,N_12180);
or U29995 (N_29995,N_11801,N_10145);
and U29996 (N_29996,N_16517,N_12113);
nand U29997 (N_29997,N_16016,N_11500);
and U29998 (N_29998,N_10241,N_16533);
or U29999 (N_29999,N_14275,N_12383);
or U30000 (N_30000,N_21298,N_23732);
nor U30001 (N_30001,N_24130,N_23281);
and U30002 (N_30002,N_28161,N_22747);
nand U30003 (N_30003,N_28878,N_21339);
or U30004 (N_30004,N_20923,N_28099);
nor U30005 (N_30005,N_20132,N_29836);
and U30006 (N_30006,N_25004,N_26256);
nor U30007 (N_30007,N_25084,N_27628);
or U30008 (N_30008,N_25674,N_24869);
and U30009 (N_30009,N_27255,N_25147);
and U30010 (N_30010,N_28281,N_29268);
nand U30011 (N_30011,N_22742,N_29657);
nand U30012 (N_30012,N_23078,N_21698);
nor U30013 (N_30013,N_27268,N_22302);
xor U30014 (N_30014,N_27245,N_25047);
nor U30015 (N_30015,N_22314,N_24925);
or U30016 (N_30016,N_20528,N_25847);
or U30017 (N_30017,N_23497,N_20362);
and U30018 (N_30018,N_20385,N_28179);
nor U30019 (N_30019,N_24849,N_23693);
xnor U30020 (N_30020,N_20148,N_21693);
nor U30021 (N_30021,N_21842,N_28298);
and U30022 (N_30022,N_28305,N_20598);
xor U30023 (N_30023,N_29603,N_28160);
nand U30024 (N_30024,N_29900,N_28303);
nand U30025 (N_30025,N_21552,N_29259);
nand U30026 (N_30026,N_28159,N_29373);
nand U30027 (N_30027,N_26655,N_21178);
nand U30028 (N_30028,N_28747,N_28682);
nand U30029 (N_30029,N_25610,N_25080);
or U30030 (N_30030,N_29665,N_28611);
nor U30031 (N_30031,N_26956,N_22117);
or U30032 (N_30032,N_27722,N_29950);
or U30033 (N_30033,N_20881,N_26483);
nand U30034 (N_30034,N_25714,N_24218);
nand U30035 (N_30035,N_20036,N_22008);
nand U30036 (N_30036,N_22956,N_20878);
nor U30037 (N_30037,N_21566,N_23509);
or U30038 (N_30038,N_20802,N_20630);
nand U30039 (N_30039,N_29348,N_22692);
and U30040 (N_30040,N_22086,N_26239);
and U30041 (N_30041,N_21471,N_23050);
nand U30042 (N_30042,N_27307,N_22865);
nand U30043 (N_30043,N_27822,N_21223);
nor U30044 (N_30044,N_23066,N_25780);
and U30045 (N_30045,N_28331,N_20302);
xnor U30046 (N_30046,N_29250,N_27981);
xor U30047 (N_30047,N_21765,N_22024);
or U30048 (N_30048,N_21961,N_23978);
nor U30049 (N_30049,N_27163,N_29894);
or U30050 (N_30050,N_21214,N_21717);
nor U30051 (N_30051,N_20759,N_23756);
nand U30052 (N_30052,N_29620,N_23857);
and U30053 (N_30053,N_28104,N_24492);
nand U30054 (N_30054,N_25155,N_24173);
nand U30055 (N_30055,N_22010,N_21240);
xnor U30056 (N_30056,N_22179,N_21506);
and U30057 (N_30057,N_29756,N_29690);
and U30058 (N_30058,N_25994,N_21222);
and U30059 (N_30059,N_21117,N_20344);
and U30060 (N_30060,N_20080,N_23774);
nand U30061 (N_30061,N_22062,N_21541);
and U30062 (N_30062,N_28545,N_22777);
or U30063 (N_30063,N_23881,N_22690);
or U30064 (N_30064,N_23533,N_26487);
or U30065 (N_30065,N_29421,N_26167);
or U30066 (N_30066,N_26079,N_20777);
and U30067 (N_30067,N_22477,N_25591);
nor U30068 (N_30068,N_26430,N_26441);
and U30069 (N_30069,N_22574,N_25419);
nor U30070 (N_30070,N_21664,N_25222);
nand U30071 (N_30071,N_23241,N_28195);
or U30072 (N_30072,N_29863,N_25765);
nand U30073 (N_30073,N_28356,N_24561);
and U30074 (N_30074,N_20869,N_21073);
xor U30075 (N_30075,N_25217,N_20276);
nor U30076 (N_30076,N_29452,N_20667);
or U30077 (N_30077,N_26446,N_22945);
nand U30078 (N_30078,N_26205,N_21301);
nor U30079 (N_30079,N_28977,N_21375);
and U30080 (N_30080,N_28049,N_21767);
or U30081 (N_30081,N_27638,N_23257);
and U30082 (N_30082,N_26259,N_23571);
or U30083 (N_30083,N_20313,N_26092);
and U30084 (N_30084,N_28144,N_22389);
xor U30085 (N_30085,N_21040,N_29360);
nand U30086 (N_30086,N_27217,N_23741);
nand U30087 (N_30087,N_28771,N_27005);
or U30088 (N_30088,N_26922,N_23474);
and U30089 (N_30089,N_29551,N_26068);
or U30090 (N_30090,N_24495,N_24363);
or U30091 (N_30091,N_21898,N_28639);
nor U30092 (N_30092,N_27546,N_27224);
xor U30093 (N_30093,N_29957,N_24224);
and U30094 (N_30094,N_20394,N_28288);
nand U30095 (N_30095,N_26209,N_24529);
or U30096 (N_30096,N_25926,N_26346);
xnor U30097 (N_30097,N_25881,N_20697);
xnor U30098 (N_30098,N_25191,N_26244);
nor U30099 (N_30099,N_25411,N_22514);
and U30100 (N_30100,N_23747,N_28572);
nand U30101 (N_30101,N_25381,N_26003);
nand U30102 (N_30102,N_20990,N_24271);
or U30103 (N_30103,N_29928,N_27838);
nand U30104 (N_30104,N_26577,N_26095);
or U30105 (N_30105,N_27079,N_21169);
nand U30106 (N_30106,N_22143,N_29285);
nor U30107 (N_30107,N_21447,N_22898);
nand U30108 (N_30108,N_22186,N_24190);
nand U30109 (N_30109,N_24933,N_29264);
and U30110 (N_30110,N_26666,N_24053);
nand U30111 (N_30111,N_22071,N_26046);
nor U30112 (N_30112,N_29135,N_20412);
nor U30113 (N_30113,N_23075,N_24096);
nand U30114 (N_30114,N_23195,N_20430);
or U30115 (N_30115,N_24023,N_21643);
or U30116 (N_30116,N_27292,N_29037);
xor U30117 (N_30117,N_28508,N_25198);
or U30118 (N_30118,N_23005,N_20659);
nand U30119 (N_30119,N_25484,N_23567);
nor U30120 (N_30120,N_28362,N_28558);
or U30121 (N_30121,N_20684,N_26644);
nor U30122 (N_30122,N_28686,N_29987);
and U30123 (N_30123,N_28974,N_29578);
xnor U30124 (N_30124,N_24668,N_25200);
and U30125 (N_30125,N_29240,N_22700);
or U30126 (N_30126,N_22111,N_24140);
and U30127 (N_30127,N_26066,N_27837);
and U30128 (N_30128,N_25285,N_21590);
and U30129 (N_30129,N_27149,N_21423);
or U30130 (N_30130,N_26713,N_29010);
nor U30131 (N_30131,N_23702,N_23468);
nor U30132 (N_30132,N_23271,N_29464);
nor U30133 (N_30133,N_29016,N_24221);
nand U30134 (N_30134,N_27387,N_22000);
and U30135 (N_30135,N_28412,N_25406);
or U30136 (N_30136,N_27897,N_25039);
nor U30137 (N_30137,N_24533,N_29461);
xor U30138 (N_30138,N_20242,N_27426);
and U30139 (N_30139,N_22834,N_27481);
nor U30140 (N_30140,N_21244,N_26833);
or U30141 (N_30141,N_26583,N_28888);
and U30142 (N_30142,N_26082,N_22684);
and U30143 (N_30143,N_24845,N_22942);
nand U30144 (N_30144,N_26820,N_22182);
and U30145 (N_30145,N_26747,N_24108);
nand U30146 (N_30146,N_27443,N_27688);
and U30147 (N_30147,N_23392,N_29524);
nor U30148 (N_30148,N_21793,N_22555);
or U30149 (N_30149,N_25002,N_24797);
nand U30150 (N_30150,N_24894,N_25949);
and U30151 (N_30151,N_25159,N_24362);
or U30152 (N_30152,N_29675,N_29732);
xnor U30153 (N_30153,N_25624,N_21659);
or U30154 (N_30154,N_20357,N_24214);
and U30155 (N_30155,N_22586,N_26172);
nand U30156 (N_30156,N_20559,N_25982);
and U30157 (N_30157,N_25062,N_25688);
nand U30158 (N_30158,N_27081,N_20826);
xor U30159 (N_30159,N_29721,N_25941);
and U30160 (N_30160,N_20382,N_23088);
and U30161 (N_30161,N_26452,N_27357);
and U30162 (N_30162,N_20520,N_25126);
nand U30163 (N_30163,N_25954,N_27640);
xor U30164 (N_30164,N_25997,N_28538);
nand U30165 (N_30165,N_22646,N_28677);
or U30166 (N_30166,N_23561,N_28014);
or U30167 (N_30167,N_25832,N_23234);
and U30168 (N_30168,N_28957,N_28086);
xnor U30169 (N_30169,N_22910,N_20600);
nor U30170 (N_30170,N_24227,N_29586);
nor U30171 (N_30171,N_21030,N_21412);
nor U30172 (N_30172,N_27869,N_22827);
nor U30173 (N_30173,N_25265,N_24259);
and U30174 (N_30174,N_28285,N_20710);
and U30175 (N_30175,N_26214,N_22900);
nor U30176 (N_30176,N_27083,N_27596);
nand U30177 (N_30177,N_20805,N_23775);
nand U30178 (N_30178,N_22936,N_23937);
and U30179 (N_30179,N_26969,N_24826);
xor U30180 (N_30180,N_25189,N_24673);
nand U30181 (N_30181,N_21808,N_25594);
nand U30182 (N_30182,N_27177,N_22264);
and U30183 (N_30183,N_25247,N_23018);
or U30184 (N_30184,N_28634,N_28627);
nand U30185 (N_30185,N_24297,N_24088);
xor U30186 (N_30186,N_26516,N_26165);
nor U30187 (N_30187,N_28689,N_23546);
nand U30188 (N_30188,N_21848,N_20367);
nand U30189 (N_30189,N_27369,N_29147);
and U30190 (N_30190,N_24855,N_21327);
nor U30191 (N_30191,N_26805,N_22554);
or U30192 (N_30192,N_28829,N_28643);
nand U30193 (N_30193,N_26254,N_23489);
or U30194 (N_30194,N_29402,N_24906);
xnor U30195 (N_30195,N_26825,N_28128);
nor U30196 (N_30196,N_25322,N_28896);
nand U30197 (N_30197,N_24528,N_21668);
or U30198 (N_30198,N_21788,N_26898);
and U30199 (N_30199,N_25344,N_29580);
or U30200 (N_30200,N_28234,N_28991);
xor U30201 (N_30201,N_28515,N_28588);
or U30202 (N_30202,N_29216,N_21391);
or U30203 (N_30203,N_24991,N_28058);
or U30204 (N_30204,N_21311,N_25606);
nor U30205 (N_30205,N_20363,N_26579);
nor U30206 (N_30206,N_27290,N_24509);
nand U30207 (N_30207,N_26984,N_21657);
or U30208 (N_30208,N_21238,N_27138);
xnor U30209 (N_30209,N_21367,N_24784);
and U30210 (N_30210,N_22868,N_24829);
nor U30211 (N_30211,N_25793,N_29293);
and U30212 (N_30212,N_23655,N_24386);
nor U30213 (N_30213,N_20319,N_21175);
and U30214 (N_30214,N_26679,N_29230);
and U30215 (N_30215,N_26901,N_21746);
or U30216 (N_30216,N_24724,N_27371);
or U30217 (N_30217,N_20162,N_20198);
or U30218 (N_30218,N_23428,N_25990);
or U30219 (N_30219,N_21398,N_29362);
nor U30220 (N_30220,N_28735,N_25557);
xnor U30221 (N_30221,N_22539,N_25014);
and U30222 (N_30222,N_20271,N_20890);
or U30223 (N_30223,N_26566,N_29084);
nand U30224 (N_30224,N_21686,N_25609);
or U30225 (N_30225,N_24425,N_26316);
xnor U30226 (N_30226,N_24475,N_23033);
and U30227 (N_30227,N_22896,N_25474);
or U30228 (N_30228,N_22361,N_27750);
nor U30229 (N_30229,N_25188,N_24084);
and U30230 (N_30230,N_29335,N_22097);
or U30231 (N_30231,N_29270,N_24637);
or U30232 (N_30232,N_21797,N_29177);
or U30233 (N_30233,N_27557,N_22031);
nor U30234 (N_30234,N_24620,N_20937);
xor U30235 (N_30235,N_22153,N_26301);
nand U30236 (N_30236,N_27437,N_29496);
or U30237 (N_30237,N_20793,N_26948);
xor U30238 (N_30238,N_20556,N_22369);
and U30239 (N_30239,N_20120,N_27478);
nor U30240 (N_30240,N_21957,N_27210);
and U30241 (N_30241,N_28369,N_27273);
and U30242 (N_30242,N_28494,N_21160);
or U30243 (N_30243,N_24120,N_26424);
and U30244 (N_30244,N_22850,N_24195);
and U30245 (N_30245,N_26628,N_26626);
or U30246 (N_30246,N_27696,N_21906);
or U30247 (N_30247,N_24154,N_23983);
nor U30248 (N_30248,N_22205,N_26699);
or U30249 (N_30249,N_23904,N_25644);
nor U30250 (N_30250,N_24632,N_20568);
nand U30251 (N_30251,N_28139,N_26366);
nand U30252 (N_30252,N_28419,N_28425);
nor U30253 (N_30253,N_20491,N_27040);
nand U30254 (N_30254,N_27013,N_21394);
nor U30255 (N_30255,N_29890,N_21294);
xnor U30256 (N_30256,N_21069,N_24257);
and U30257 (N_30257,N_23849,N_23322);
nor U30258 (N_30258,N_27260,N_26704);
and U30259 (N_30259,N_28310,N_26284);
nand U30260 (N_30260,N_23815,N_20643);
nand U30261 (N_30261,N_23593,N_27413);
or U30262 (N_30262,N_24278,N_20701);
or U30263 (N_30263,N_23758,N_29035);
nand U30264 (N_30264,N_21673,N_27657);
nor U30265 (N_30265,N_28764,N_29613);
nor U30266 (N_30266,N_26940,N_27489);
and U30267 (N_30267,N_29069,N_24794);
and U30268 (N_30268,N_22036,N_20790);
or U30269 (N_30269,N_26022,N_20455);
or U30270 (N_30270,N_27700,N_21665);
nand U30271 (N_30271,N_25685,N_25494);
and U30272 (N_30272,N_20415,N_29549);
nand U30273 (N_30273,N_29482,N_26450);
and U30274 (N_30274,N_20870,N_29581);
or U30275 (N_30275,N_24114,N_25544);
and U30276 (N_30276,N_26861,N_21909);
and U30277 (N_30277,N_20993,N_23047);
and U30278 (N_30278,N_29503,N_27731);
and U30279 (N_30279,N_24150,N_21652);
or U30280 (N_30280,N_23357,N_27488);
nor U30281 (N_30281,N_28085,N_29101);
or U30282 (N_30282,N_22531,N_24378);
or U30283 (N_30283,N_23012,N_22126);
nand U30284 (N_30284,N_23114,N_29656);
xor U30285 (N_30285,N_22052,N_21736);
xnor U30286 (N_30286,N_29639,N_26162);
and U30287 (N_30287,N_27353,N_28266);
nand U30288 (N_30288,N_21393,N_26943);
nand U30289 (N_30289,N_24578,N_26983);
nand U30290 (N_30290,N_28065,N_22164);
nor U30291 (N_30291,N_23805,N_25110);
xnor U30292 (N_30292,N_28672,N_25236);
and U30293 (N_30293,N_20166,N_20096);
and U30294 (N_30294,N_20517,N_21733);
or U30295 (N_30295,N_25719,N_25028);
or U30296 (N_30296,N_24564,N_29880);
or U30297 (N_30297,N_25393,N_28067);
and U30298 (N_30298,N_22216,N_29847);
or U30299 (N_30299,N_24743,N_28683);
or U30300 (N_30300,N_20816,N_24872);
and U30301 (N_30301,N_25827,N_21714);
nand U30302 (N_30302,N_29772,N_28370);
and U30303 (N_30303,N_20263,N_22760);
and U30304 (N_30304,N_24865,N_27970);
or U30305 (N_30305,N_25262,N_22025);
xnor U30306 (N_30306,N_24061,N_26409);
or U30307 (N_30307,N_26767,N_23198);
xor U30308 (N_30308,N_21533,N_22523);
or U30309 (N_30309,N_27356,N_29915);
nand U30310 (N_30310,N_21565,N_26740);
nand U30311 (N_30311,N_22858,N_28509);
nor U30312 (N_30312,N_20590,N_27439);
nand U30313 (N_30313,N_28716,N_27418);
nor U30314 (N_30314,N_22547,N_24634);
or U30315 (N_30315,N_21575,N_21563);
or U30316 (N_30316,N_28311,N_28731);
and U30317 (N_30317,N_28059,N_29363);
and U30318 (N_30318,N_26934,N_22388);
and U30319 (N_30319,N_21726,N_21264);
or U30320 (N_30320,N_21364,N_29097);
nand U30321 (N_30321,N_28187,N_26090);
nor U30322 (N_30322,N_29056,N_24508);
nand U30323 (N_30323,N_28913,N_24220);
or U30324 (N_30324,N_23364,N_23036);
nand U30325 (N_30325,N_28006,N_27687);
nand U30326 (N_30326,N_23801,N_25331);
nor U30327 (N_30327,N_28981,N_28021);
nand U30328 (N_30328,N_25248,N_28920);
nor U30329 (N_30329,N_25261,N_24299);
and U30330 (N_30330,N_26818,N_26911);
nand U30331 (N_30331,N_25421,N_26122);
nand U30332 (N_30332,N_27367,N_20899);
or U30333 (N_30333,N_23220,N_29741);
or U30334 (N_30334,N_26721,N_20406);
and U30335 (N_30335,N_29131,N_26139);
and U30336 (N_30336,N_21308,N_22217);
and U30337 (N_30337,N_27678,N_29782);
xnor U30338 (N_30338,N_21607,N_22570);
and U30339 (N_30339,N_23710,N_28025);
or U30340 (N_30340,N_26846,N_24357);
nand U30341 (N_30341,N_29686,N_20593);
and U30342 (N_30342,N_21997,N_22620);
or U30343 (N_30343,N_22508,N_27860);
and U30344 (N_30344,N_29419,N_28431);
xor U30345 (N_30345,N_28376,N_29407);
or U30346 (N_30346,N_20980,N_27251);
nand U30347 (N_30347,N_23784,N_20786);
or U30348 (N_30348,N_22141,N_27244);
nand U30349 (N_30349,N_27794,N_21556);
and U30350 (N_30350,N_25479,N_23288);
nor U30351 (N_30351,N_24851,N_25659);
nand U30352 (N_30352,N_28610,N_22593);
and U30353 (N_30353,N_25882,N_26023);
nand U30354 (N_30354,N_29939,N_23549);
or U30355 (N_30355,N_21690,N_23676);
nor U30356 (N_30356,N_27036,N_20836);
nand U30357 (N_30357,N_21782,N_28983);
nand U30358 (N_30358,N_28740,N_20461);
or U30359 (N_30359,N_20072,N_23961);
nand U30360 (N_30360,N_29051,N_29630);
and U30361 (N_30361,N_26445,N_23164);
nor U30362 (N_30362,N_25276,N_22444);
nand U30363 (N_30363,N_29884,N_23006);
xnor U30364 (N_30364,N_24432,N_26754);
nor U30365 (N_30365,N_29239,N_21372);
nand U30366 (N_30366,N_24370,N_22676);
and U30367 (N_30367,N_27520,N_24955);
and U30368 (N_30368,N_26141,N_20865);
nor U30369 (N_30369,N_29027,N_23771);
or U30370 (N_30370,N_20007,N_25566);
and U30371 (N_30371,N_26104,N_25304);
nand U30372 (N_30372,N_29989,N_23440);
nand U30373 (N_30373,N_24079,N_25316);
or U30374 (N_30374,N_22710,N_22298);
or U30375 (N_30375,N_24908,N_20687);
and U30376 (N_30376,N_21897,N_20585);
nor U30377 (N_30377,N_29930,N_27004);
or U30378 (N_30378,N_24556,N_24042);
nor U30379 (N_30379,N_29601,N_26174);
and U30380 (N_30380,N_20090,N_28522);
and U30381 (N_30381,N_20025,N_20750);
or U30382 (N_30382,N_24428,N_27770);
nor U30383 (N_30383,N_28391,N_23292);
nand U30384 (N_30384,N_26942,N_26258);
nand U30385 (N_30385,N_29684,N_29903);
nor U30386 (N_30386,N_28833,N_28265);
and U30387 (N_30387,N_24775,N_23753);
nor U30388 (N_30388,N_24523,N_22017);
nand U30389 (N_30389,N_23600,N_23082);
nor U30390 (N_30390,N_28937,N_23995);
nor U30391 (N_30391,N_21635,N_27117);
nand U30392 (N_30392,N_26431,N_29314);
or U30393 (N_30393,N_26006,N_28063);
nand U30394 (N_30394,N_27153,N_25090);
or U30395 (N_30395,N_26604,N_29610);
xor U30396 (N_30396,N_28927,N_21642);
or U30397 (N_30397,N_20438,N_21731);
and U30398 (N_30398,N_20566,N_27764);
nand U30399 (N_30399,N_28566,N_29937);
nor U30400 (N_30400,N_21812,N_24587);
or U30401 (N_30401,N_20800,N_25924);
and U30402 (N_30402,N_20938,N_20292);
or U30403 (N_30403,N_27852,N_29800);
and U30404 (N_30404,N_23466,N_24263);
nor U30405 (N_30405,N_29463,N_24585);
xor U30406 (N_30406,N_29605,N_27175);
or U30407 (N_30407,N_26933,N_22300);
or U30408 (N_30408,N_24124,N_22659);
nor U30409 (N_30409,N_28151,N_20743);
and U30410 (N_30410,N_26788,N_27704);
nand U30411 (N_30411,N_23478,N_22500);
nand U30412 (N_30412,N_29976,N_26500);
nand U30413 (N_30413,N_28788,N_29985);
or U30414 (N_30414,N_28599,N_20646);
or U30415 (N_30415,N_21151,N_25942);
and U30416 (N_30416,N_22725,N_28465);
or U30417 (N_30417,N_29597,N_29660);
and U30418 (N_30418,N_20698,N_27589);
and U30419 (N_30419,N_27570,N_25687);
or U30420 (N_30420,N_22633,N_29735);
xor U30421 (N_30421,N_26429,N_21768);
nand U30422 (N_30422,N_27730,N_21576);
nand U30423 (N_30423,N_23273,N_27509);
or U30424 (N_30424,N_20337,N_28393);
nand U30425 (N_30425,N_25617,N_25181);
and U30426 (N_30426,N_26935,N_24020);
nand U30427 (N_30427,N_27326,N_26183);
nor U30428 (N_30428,N_27476,N_27455);
nand U30429 (N_30429,N_22044,N_23465);
or U30430 (N_30430,N_28345,N_28277);
or U30431 (N_30431,N_26063,N_22230);
nand U30432 (N_30432,N_23347,N_25391);
xnor U30433 (N_30433,N_20004,N_24940);
and U30434 (N_30434,N_21280,N_27646);
xor U30435 (N_30435,N_29401,N_29801);
and U30436 (N_30436,N_21687,N_29679);
nor U30437 (N_30437,N_26683,N_27874);
nor U30438 (N_30438,N_29541,N_28307);
or U30439 (N_30439,N_25409,N_20506);
or U30440 (N_30440,N_23620,N_29980);
or U30441 (N_30441,N_27862,N_22140);
xnor U30442 (N_30442,N_25660,N_27465);
and U30443 (N_30443,N_27352,N_20466);
and U30444 (N_30444,N_21709,N_28280);
and U30445 (N_30445,N_26702,N_28073);
nand U30446 (N_30446,N_22457,N_23487);
or U30447 (N_30447,N_29831,N_23882);
and U30448 (N_30448,N_27077,N_22004);
nand U30449 (N_30449,N_26652,N_28999);
and U30450 (N_30450,N_22675,N_28846);
nor U30451 (N_30451,N_20981,N_24537);
and U30452 (N_30452,N_25721,N_21177);
and U30453 (N_30453,N_28678,N_26708);
and U30454 (N_30454,N_29638,N_21161);
nand U30455 (N_30455,N_21544,N_27950);
or U30456 (N_30456,N_28680,N_25343);
and U30457 (N_30457,N_21928,N_22014);
or U30458 (N_30458,N_29307,N_28842);
and U30459 (N_30459,N_22360,N_25356);
nand U30460 (N_30460,N_25910,N_29116);
and U30461 (N_30461,N_27365,N_29918);
nand U30462 (N_30462,N_26012,N_21963);
nor U30463 (N_30463,N_28479,N_26601);
nor U30464 (N_30464,N_27567,N_27714);
nand U30465 (N_30465,N_29310,N_24880);
nor U30466 (N_30466,N_28226,N_20859);
nor U30467 (N_30467,N_24978,N_27533);
xnor U30468 (N_30468,N_24435,N_22304);
nor U30469 (N_30469,N_28687,N_29150);
nor U30470 (N_30470,N_20119,N_20613);
or U30471 (N_30471,N_20549,N_24462);
xnor U30472 (N_30472,N_26472,N_23932);
xnor U30473 (N_30473,N_29413,N_25530);
and U30474 (N_30474,N_22482,N_21958);
nand U30475 (N_30475,N_22480,N_25903);
and U30476 (N_30476,N_24867,N_25462);
or U30477 (N_30477,N_23851,N_20943);
or U30478 (N_30478,N_22697,N_21065);
or U30479 (N_30479,N_22866,N_28252);
nand U30480 (N_30480,N_25715,N_21070);
nor U30481 (N_30481,N_29914,N_28493);
nor U30482 (N_30482,N_25923,N_29462);
or U30483 (N_30483,N_24466,N_24708);
nand U30484 (N_30484,N_26438,N_25224);
nand U30485 (N_30485,N_28803,N_21883);
and U30486 (N_30486,N_22963,N_22999);
nand U30487 (N_30487,N_20038,N_29932);
nand U30488 (N_30488,N_29953,N_20485);
or U30489 (N_30489,N_28595,N_27161);
nand U30490 (N_30490,N_29817,N_21139);
and U30491 (N_30491,N_29923,N_24814);
nor U30492 (N_30492,N_29171,N_23768);
nand U30493 (N_30493,N_24074,N_23626);
nor U30494 (N_30494,N_23134,N_20015);
nor U30495 (N_30495,N_29893,N_25974);
and U30496 (N_30496,N_20041,N_20904);
nor U30497 (N_30497,N_20592,N_26649);
nor U30498 (N_30498,N_21388,N_25420);
or U30499 (N_30499,N_25952,N_20222);
nand U30500 (N_30500,N_20835,N_22410);
or U30501 (N_30501,N_20423,N_27065);
nor U30502 (N_30502,N_25182,N_29655);
nor U30503 (N_30503,N_21526,N_23944);
or U30504 (N_30504,N_27111,N_23960);
and U30505 (N_30505,N_20425,N_29938);
xnor U30506 (N_30506,N_21921,N_28759);
xor U30507 (N_30507,N_29559,N_22378);
nor U30508 (N_30508,N_20744,N_24029);
nor U30509 (N_30509,N_25490,N_21209);
nor U30510 (N_30510,N_26444,N_27767);
xnor U30511 (N_30511,N_24963,N_21130);
or U30512 (N_30512,N_27444,N_24179);
nand U30513 (N_30513,N_27491,N_28782);
and U30514 (N_30514,N_28971,N_20308);
xor U30515 (N_30515,N_26945,N_27994);
or U30516 (N_30516,N_27716,N_24476);
nand U30517 (N_30517,N_24075,N_29678);
and U30518 (N_30518,N_28886,N_25428);
and U30519 (N_30519,N_26608,N_24417);
and U30520 (N_30520,N_25519,N_29378);
nor U30521 (N_30521,N_27402,N_25938);
and U30522 (N_30522,N_29723,N_24718);
nand U30523 (N_30523,N_28631,N_29438);
or U30524 (N_30524,N_24004,N_25446);
or U30525 (N_30525,N_24300,N_25332);
nor U30526 (N_30526,N_20087,N_20747);
or U30527 (N_30527,N_24958,N_27474);
nand U30528 (N_30528,N_29044,N_28273);
nor U30529 (N_30529,N_26010,N_26199);
nor U30530 (N_30530,N_22561,N_24011);
nand U30531 (N_30531,N_20247,N_24209);
nor U30532 (N_30532,N_28567,N_23651);
and U30533 (N_30533,N_29192,N_21107);
and U30534 (N_30534,N_24071,N_27254);
nand U30535 (N_30535,N_27243,N_20186);
or U30536 (N_30536,N_24474,N_24590);
and U30537 (N_30537,N_25588,N_28109);
nor U30538 (N_30538,N_25444,N_28730);
and U30539 (N_30539,N_20028,N_28456);
or U30540 (N_30540,N_23624,N_23720);
or U30541 (N_30541,N_21404,N_29102);
nand U30542 (N_30542,N_26799,N_21524);
or U30543 (N_30543,N_22098,N_21080);
nand U30544 (N_30544,N_28923,N_28662);
nand U30545 (N_30545,N_27929,N_29468);
and U30546 (N_30546,N_24460,N_26734);
nand U30547 (N_30547,N_27425,N_25346);
or U30548 (N_30548,N_21985,N_21578);
nand U30549 (N_30549,N_22305,N_21111);
nand U30550 (N_30550,N_23760,N_22654);
and U30551 (N_30551,N_22094,N_22825);
nor U30552 (N_30552,N_21165,N_21405);
or U30553 (N_30553,N_29138,N_24823);
and U30554 (N_30554,N_25257,N_21125);
xor U30555 (N_30555,N_20712,N_29561);
nor U30556 (N_30556,N_26851,N_25587);
nor U30557 (N_30557,N_21622,N_27689);
nand U30558 (N_30558,N_22994,N_24810);
and U30559 (N_30559,N_29005,N_24285);
and U30560 (N_30560,N_24352,N_25007);
and U30561 (N_30561,N_28818,N_28755);
xnor U30562 (N_30562,N_29471,N_21328);
nor U30563 (N_30563,N_20088,N_26944);
or U30564 (N_30564,N_21152,N_26133);
or U30565 (N_30565,N_23356,N_29243);
xor U30566 (N_30566,N_28414,N_20019);
nand U30567 (N_30567,N_26808,N_20654);
nand U30568 (N_30568,N_24083,N_20874);
nand U30569 (N_30569,N_29296,N_25339);
and U30570 (N_30570,N_26558,N_26345);
and U30571 (N_30571,N_28898,N_21778);
nor U30572 (N_30572,N_26522,N_26766);
or U30573 (N_30573,N_21675,N_21755);
or U30574 (N_30574,N_24579,N_29784);
nand U30575 (N_30575,N_26508,N_29526);
nor U30576 (N_30576,N_24703,N_22463);
or U30577 (N_30577,N_23388,N_24660);
nand U30578 (N_30578,N_23106,N_29276);
nand U30579 (N_30579,N_25472,N_20778);
or U30580 (N_30580,N_25541,N_22609);
nor U30581 (N_30581,N_28719,N_22954);
nor U30582 (N_30582,N_29076,N_26333);
or U30583 (N_30583,N_21206,N_27158);
nor U30584 (N_30584,N_28229,N_24534);
and U30585 (N_30585,N_27612,N_26996);
and U30586 (N_30586,N_23024,N_23381);
or U30587 (N_30587,N_22683,N_28455);
nor U30588 (N_30588,N_27811,N_24532);
nand U30589 (N_30589,N_29442,N_23612);
nor U30590 (N_30590,N_24323,N_21012);
nand U30591 (N_30591,N_24487,N_29637);
xnor U30592 (N_30592,N_20649,N_25743);
or U30593 (N_30593,N_21470,N_21783);
and U30594 (N_30594,N_28103,N_29090);
nor U30595 (N_30595,N_29540,N_28758);
or U30596 (N_30596,N_22419,N_29345);
nor U30597 (N_30597,N_21996,N_21067);
nand U30598 (N_30598,N_21128,N_22672);
or U30599 (N_30599,N_26681,N_21155);
nor U30600 (N_30600,N_22198,N_22163);
nand U30601 (N_30601,N_22712,N_20725);
and U30602 (N_30602,N_29619,N_22969);
and U30603 (N_30603,N_20154,N_24177);
and U30604 (N_30604,N_21403,N_24593);
nand U30605 (N_30605,N_21530,N_21754);
nand U30606 (N_30606,N_27129,N_22413);
xor U30607 (N_30607,N_29019,N_22124);
or U30608 (N_30608,N_27076,N_24344);
nor U30609 (N_30609,N_26462,N_22716);
or U30610 (N_30610,N_29874,N_24719);
or U30611 (N_30611,N_27216,N_26017);
and U30612 (N_30612,N_24031,N_26947);
or U30613 (N_30613,N_25518,N_25324);
nor U30614 (N_30614,N_20400,N_28606);
and U30615 (N_30615,N_27228,N_27599);
nand U30616 (N_30616,N_27400,N_24948);
and U30617 (N_30617,N_25488,N_20705);
nor U30618 (N_30618,N_29904,N_23382);
nand U30619 (N_30619,N_26866,N_28125);
or U30620 (N_30620,N_29380,N_23298);
nand U30621 (N_30621,N_21959,N_25577);
or U30622 (N_30622,N_26596,N_27671);
nand U30623 (N_30623,N_28986,N_20822);
or U30624 (N_30624,N_21250,N_24419);
or U30625 (N_30625,N_22821,N_22813);
nand U30626 (N_30626,N_21638,N_22829);
or U30627 (N_30627,N_27055,N_28210);
or U30628 (N_30628,N_24793,N_22063);
nand U30629 (N_30629,N_28022,N_23216);
or U30630 (N_30630,N_22665,N_25957);
or U30631 (N_30631,N_25639,N_25169);
nand U30632 (N_30632,N_27033,N_22248);
nor U30633 (N_30633,N_25897,N_25750);
and U30634 (N_30634,N_21730,N_22422);
nand U30635 (N_30635,N_29822,N_25469);
nor U30636 (N_30636,N_21931,N_29271);
and U30637 (N_30637,N_20969,N_27440);
nor U30638 (N_30638,N_25445,N_21216);
or U30639 (N_30639,N_29257,N_25218);
nor U30640 (N_30640,N_29261,N_24237);
nor U30641 (N_30641,N_27692,N_23121);
or U30642 (N_30642,N_21572,N_27791);
or U30643 (N_30643,N_26988,N_23245);
and U30644 (N_30644,N_28030,N_25079);
and U30645 (N_30645,N_21305,N_29127);
nor U30646 (N_30646,N_28612,N_27459);
xnor U30647 (N_30647,N_26386,N_20254);
and U30648 (N_30648,N_22830,N_25766);
and U30649 (N_30649,N_21794,N_28840);
nand U30650 (N_30650,N_23200,N_22734);
nand U30651 (N_30651,N_26067,N_23723);
and U30652 (N_30652,N_27293,N_29798);
nor U30653 (N_30653,N_26829,N_22493);
nand U30654 (N_30654,N_25289,N_22433);
and U30655 (N_30655,N_25986,N_20801);
and U30656 (N_30656,N_28300,N_29592);
nand U30657 (N_30657,N_25120,N_23543);
nand U30658 (N_30658,N_24366,N_20525);
nor U30659 (N_30659,N_28048,N_26850);
and U30660 (N_30660,N_25884,N_24858);
nor U30661 (N_30661,N_21993,N_25310);
nand U30662 (N_30662,N_26817,N_28212);
nor U30663 (N_30663,N_26226,N_20497);
nor U30664 (N_30664,N_23658,N_27749);
and U30665 (N_30665,N_20315,N_22214);
nand U30666 (N_30666,N_28597,N_27257);
nor U30667 (N_30667,N_20273,N_20233);
and U30668 (N_30668,N_22925,N_21331);
nor U30669 (N_30669,N_23031,N_23646);
and U30670 (N_30670,N_20930,N_24510);
and U30671 (N_30671,N_29397,N_20365);
nand U30672 (N_30672,N_24542,N_26932);
nand U30673 (N_30673,N_26555,N_26100);
xnor U30674 (N_30674,N_23371,N_21967);
nand U30675 (N_30675,N_26189,N_25368);
and U30676 (N_30676,N_24575,N_21817);
or U30677 (N_30677,N_26647,N_21953);
xnor U30678 (N_30678,N_23412,N_23685);
or U30679 (N_30679,N_28355,N_21670);
or U30680 (N_30680,N_22235,N_27484);
or U30681 (N_30681,N_28660,N_23080);
xor U30682 (N_30682,N_29773,N_24565);
or U30683 (N_30683,N_24560,N_25290);
or U30684 (N_30684,N_29579,N_24044);
or U30685 (N_30685,N_24843,N_28365);
nor U30686 (N_30686,N_20806,N_24208);
nand U30687 (N_30687,N_23287,N_22985);
nor U30688 (N_30688,N_20396,N_28736);
nor U30689 (N_30689,N_23502,N_29693);
xor U30690 (N_30690,N_20726,N_28931);
nor U30691 (N_30691,N_26044,N_26282);
nand U30692 (N_30692,N_26298,N_23186);
nor U30693 (N_30693,N_27346,N_21129);
nand U30694 (N_30694,N_25128,N_25716);
nand U30695 (N_30695,N_28570,N_21983);
nand U30696 (N_30696,N_20979,N_23380);
or U30697 (N_30697,N_28428,N_29183);
or U30698 (N_30698,N_20526,N_29746);
and U30699 (N_30699,N_24841,N_29720);
nand U30700 (N_30700,N_21377,N_22628);
nand U30701 (N_30701,N_22458,N_29248);
nand U30702 (N_30702,N_21505,N_29372);
nor U30703 (N_30703,N_26222,N_24687);
or U30704 (N_30704,N_20887,N_21469);
nand U30705 (N_30705,N_24412,N_23258);
nand U30706 (N_30706,N_26490,N_29159);
nor U30707 (N_30707,N_25657,N_21738);
nor U30708 (N_30708,N_27234,N_24439);
nor U30709 (N_30709,N_22515,N_29403);
or U30710 (N_30710,N_29262,N_25953);
xnor U30711 (N_30711,N_23687,N_25782);
nand U30712 (N_30712,N_27751,N_21987);
nor U30713 (N_30713,N_20460,N_25975);
and U30714 (N_30714,N_24382,N_21234);
xor U30715 (N_30715,N_21531,N_23856);
and U30716 (N_30716,N_25347,N_22918);
xor U30717 (N_30717,N_25048,N_24456);
or U30718 (N_30718,N_21704,N_22642);
xnor U30719 (N_30719,N_27900,N_25187);
and U30720 (N_30720,N_23898,N_26928);
nor U30721 (N_30721,N_27310,N_24392);
nor U30722 (N_30722,N_23860,N_25729);
or U30723 (N_30723,N_26640,N_22540);
or U30724 (N_30724,N_29323,N_22801);
xor U30725 (N_30725,N_25811,N_22793);
and U30726 (N_30726,N_26469,N_25710);
or U30727 (N_30727,N_23934,N_29614);
or U30728 (N_30728,N_25589,N_25727);
nand U30729 (N_30729,N_22992,N_20228);
xnor U30730 (N_30730,N_21561,N_25861);
nor U30731 (N_30731,N_25655,N_25638);
or U30732 (N_30732,N_21202,N_26630);
or U30733 (N_30733,N_24822,N_28954);
nor U30734 (N_30734,N_21499,N_28912);
nor U30735 (N_30735,N_25452,N_22588);
nor U30736 (N_30736,N_29696,N_28628);
nor U30737 (N_30737,N_28379,N_27626);
and U30738 (N_30738,N_26529,N_27313);
or U30739 (N_30739,N_21086,N_29572);
or U30740 (N_30740,N_21924,N_24969);
nor U30741 (N_30741,N_21351,N_22766);
and U30742 (N_30742,N_26470,N_29908);
xor U30743 (N_30743,N_26563,N_29398);
and U30744 (N_30744,N_27768,N_22694);
nor U30745 (N_30745,N_20736,N_29085);
nor U30746 (N_30746,N_28395,N_26521);
nor U30747 (N_30747,N_21137,N_25050);
nor U30748 (N_30748,N_27911,N_21232);
nand U30749 (N_30749,N_24167,N_24287);
xor U30750 (N_30750,N_25195,N_29713);
or U30751 (N_30751,N_20212,N_27102);
or U30752 (N_30752,N_28869,N_22113);
nor U30753 (N_30753,N_20541,N_21038);
nor U30754 (N_30754,N_26049,N_25451);
nor U30755 (N_30755,N_21041,N_23192);
nor U30756 (N_30756,N_28045,N_26008);
nand U30757 (N_30757,N_20748,N_26363);
nand U30758 (N_30758,N_22079,N_23376);
nor U30759 (N_30759,N_21281,N_23202);
xor U30760 (N_30760,N_29783,N_23935);
nor U30761 (N_30761,N_22181,N_21615);
or U30762 (N_30762,N_28155,N_29180);
nand U30763 (N_30763,N_23517,N_21358);
xor U30764 (N_30764,N_23349,N_23452);
or U30765 (N_30765,N_23902,N_24946);
and U30766 (N_30766,N_22091,N_21094);
xnor U30767 (N_30767,N_24280,N_27584);
or U30768 (N_30768,N_26706,N_25575);
or U30769 (N_30769,N_26636,N_25641);
nor U30770 (N_30770,N_21057,N_27054);
and U30771 (N_30771,N_28404,N_25175);
nor U30772 (N_30772,N_27789,N_23605);
nor U30773 (N_30773,N_29095,N_28505);
or U30774 (N_30774,N_25790,N_20815);
nor U30775 (N_30775,N_27632,N_26709);
or U30776 (N_30776,N_27442,N_23333);
or U30777 (N_30777,N_26168,N_20419);
nor U30778 (N_30778,N_28062,N_25122);
or U30779 (N_30779,N_26210,N_26705);
and U30780 (N_30780,N_25177,N_26761);
or U30781 (N_30781,N_27798,N_24063);
nand U30782 (N_30782,N_20515,N_24191);
and U30783 (N_30783,N_29266,N_25355);
nand U30784 (N_30784,N_28517,N_26349);
or U30785 (N_30785,N_25692,N_20264);
nand U30786 (N_30786,N_21774,N_20947);
or U30787 (N_30787,N_21215,N_23049);
nand U30788 (N_30788,N_29507,N_25022);
or U30789 (N_30789,N_20692,N_24712);
or U30790 (N_30790,N_21103,N_26553);
nor U30791 (N_30791,N_23188,N_28241);
nor U30792 (N_30792,N_23848,N_23171);
and U30793 (N_30793,N_29269,N_27378);
nor U30794 (N_30794,N_20901,N_27139);
and U30795 (N_30795,N_22407,N_25935);
nand U30796 (N_30796,N_29064,N_21660);
and U30797 (N_30797,N_23947,N_29554);
nor U30798 (N_30798,N_21131,N_23738);
and U30799 (N_30799,N_29855,N_21120);
or U30800 (N_30800,N_28038,N_21661);
and U30801 (N_30801,N_23048,N_20807);
and U30802 (N_30802,N_23500,N_20789);
and U30803 (N_30803,N_25708,N_21399);
or U30804 (N_30804,N_29877,N_26877);
or U30805 (N_30805,N_27912,N_29539);
or U30806 (N_30806,N_28361,N_23203);
nor U30807 (N_30807,N_24754,N_29867);
nand U30808 (N_30808,N_21624,N_21150);
nor U30809 (N_30809,N_29733,N_26473);
nor U30810 (N_30810,N_25510,N_23148);
or U30811 (N_30811,N_29821,N_28651);
nor U30812 (N_30812,N_26714,N_24945);
and U30813 (N_30813,N_21247,N_25814);
xnor U30814 (N_30814,N_25493,N_20230);
or U30815 (N_30815,N_21899,N_20459);
nand U30816 (N_30816,N_28259,N_23352);
and U30817 (N_30817,N_20427,N_24710);
xor U30818 (N_30818,N_25670,N_21691);
nor U30819 (N_30819,N_26703,N_26399);
and U30820 (N_30820,N_20324,N_23175);
nor U30821 (N_30821,N_25826,N_27002);
or U30822 (N_30822,N_20959,N_28711);
nand U30823 (N_30823,N_22686,N_25009);
nand U30824 (N_30824,N_26893,N_24757);
and U30825 (N_30825,N_28772,N_23230);
or U30826 (N_30826,N_20885,N_20075);
and U30827 (N_30827,N_23447,N_24998);
nand U30828 (N_30828,N_21000,N_27408);
or U30829 (N_30829,N_26160,N_25698);
xor U30830 (N_30830,N_24507,N_21426);
nand U30831 (N_30831,N_24711,N_25877);
nor U30832 (N_30832,N_28779,N_21310);
and U30833 (N_30833,N_22773,N_23637);
xnor U30834 (N_30834,N_20623,N_26595);
nand U30835 (N_30835,N_24269,N_29677);
nor U30836 (N_30836,N_26848,N_20368);
or U30837 (N_30837,N_25699,N_20799);
and U30838 (N_30838,N_25199,N_29254);
nand U30839 (N_30839,N_26633,N_21448);
and U30840 (N_30840,N_28386,N_26892);
or U30841 (N_30841,N_28261,N_27623);
nor U30842 (N_30842,N_22538,N_23389);
or U30843 (N_30843,N_28529,N_22730);
nand U30844 (N_30844,N_28530,N_23407);
or U30845 (N_30845,N_22888,N_22943);
nor U30846 (N_30846,N_26899,N_29544);
nor U30847 (N_30847,N_26930,N_23105);
nand U30848 (N_30848,N_24954,N_20996);
nor U30849 (N_30849,N_20282,N_24622);
or U30850 (N_30850,N_20309,N_20417);
and U30851 (N_30851,N_26195,N_20073);
xor U30852 (N_30852,N_28761,N_23967);
nor U30853 (N_30853,N_27999,N_20916);
nor U30854 (N_30854,N_28703,N_26632);
and U30855 (N_30855,N_27146,N_21342);
or U30856 (N_30856,N_23959,N_22729);
nand U30857 (N_30857,N_28542,N_27069);
or U30858 (N_30858,N_20443,N_21022);
nor U30859 (N_30859,N_24226,N_21024);
and U30860 (N_30860,N_22183,N_23086);
nand U30861 (N_30861,N_23766,N_21644);
and U30862 (N_30862,N_25680,N_24411);
and U30863 (N_30863,N_26304,N_23606);
nor U30864 (N_30864,N_29612,N_29122);
or U30865 (N_30865,N_26414,N_25948);
and U30866 (N_30866,N_27699,N_25314);
and U30867 (N_30867,N_26007,N_24681);
nor U30868 (N_30868,N_27593,N_26819);
nor U30869 (N_30869,N_22965,N_21752);
nor U30870 (N_30870,N_26142,N_28670);
nand U30871 (N_30871,N_23030,N_27782);
and U30872 (N_30872,N_29079,N_25676);
nand U30873 (N_30873,N_25731,N_21536);
nor U30874 (N_30874,N_20285,N_27571);
and U30875 (N_30875,N_20651,N_29487);
nor U30876 (N_30876,N_27532,N_21811);
xnor U30877 (N_30877,N_26164,N_20851);
nand U30878 (N_30878,N_27521,N_26085);
nor U30879 (N_30879,N_27775,N_24461);
or U30880 (N_30880,N_23840,N_20671);
and U30881 (N_30881,N_22617,N_20187);
and U30882 (N_30882,N_23614,N_22955);
and U30883 (N_30883,N_26330,N_23163);
nor U30884 (N_30884,N_24769,N_29699);
or U30885 (N_30885,N_23348,N_25424);
nand U30886 (N_30886,N_28079,N_23423);
or U30887 (N_30887,N_22191,N_26502);
and U30888 (N_30888,N_25538,N_29389);
and U30889 (N_30889,N_28069,N_20618);
nand U30890 (N_30890,N_27642,N_26786);
nand U30891 (N_30891,N_21074,N_23816);
nor U30892 (N_30892,N_20581,N_26515);
or U30893 (N_30893,N_23211,N_25377);
and U30894 (N_30894,N_23107,N_28858);
or U30895 (N_30895,N_22046,N_26274);
and U30896 (N_30896,N_26859,N_24844);
and U30897 (N_30897,N_27221,N_24599);
nand U30898 (N_30898,N_23536,N_28239);
nand U30899 (N_30899,N_27188,N_23762);
or U30900 (N_30900,N_23920,N_22223);
xor U30901 (N_30901,N_25037,N_27795);
nand U30902 (N_30902,N_22950,N_26671);
nor U30903 (N_30903,N_26087,N_23178);
or U30904 (N_30904,N_20732,N_29748);
and U30905 (N_30905,N_21023,N_27849);
nor U30906 (N_30906,N_24048,N_22818);
and U30907 (N_30907,N_21400,N_25299);
or U30908 (N_30908,N_27433,N_21413);
and U30909 (N_30909,N_27001,N_21267);
and U30910 (N_30910,N_23872,N_29356);
nor U30911 (N_30911,N_28247,N_29469);
and U30912 (N_30912,N_28600,N_26099);
nor U30913 (N_30913,N_25096,N_21791);
xor U30914 (N_30914,N_26405,N_27297);
xnor U30915 (N_30915,N_22750,N_25752);
nand U30916 (N_30916,N_21109,N_29692);
nor U30917 (N_30917,N_29476,N_26591);
and U30918 (N_30918,N_20450,N_21188);
or U30919 (N_30919,N_24694,N_29231);
or U30920 (N_30920,N_28691,N_24594);
nand U30921 (N_30921,N_29457,N_20912);
nand U30922 (N_30922,N_21770,N_22199);
xnor U30923 (N_30923,N_27583,N_22049);
nand U30924 (N_30924,N_24680,N_22543);
and U30925 (N_30925,N_25970,N_24773);
and U30926 (N_30926,N_21093,N_27736);
or U30927 (N_30927,N_28000,N_22651);
nand U30928 (N_30928,N_27043,N_28989);
nor U30929 (N_30929,N_21262,N_28092);
nand U30930 (N_30930,N_24170,N_23671);
nand U30931 (N_30931,N_20719,N_29891);
nor U30932 (N_30932,N_23845,N_27894);
and U30933 (N_30933,N_20633,N_24818);
and U30934 (N_30934,N_23940,N_20142);
nor U30935 (N_30935,N_21751,N_26777);
nor U30936 (N_30936,N_29514,N_24765);
nor U30937 (N_30937,N_25250,N_27560);
or U30938 (N_30938,N_25992,N_22940);
nand U30939 (N_30939,N_23025,N_24957);
nor U30940 (N_30940,N_29780,N_21346);
nor U30941 (N_30941,N_26966,N_27885);
nor U30942 (N_30942,N_29789,N_29922);
nand U30943 (N_30943,N_22544,N_23424);
nor U30944 (N_30944,N_25480,N_27516);
nor U30945 (N_30945,N_24887,N_24633);
nand U30946 (N_30946,N_20206,N_24207);
nand U30947 (N_30947,N_25255,N_23063);
nor U30948 (N_30948,N_21558,N_21970);
and U30949 (N_30949,N_28679,N_26311);
or U30950 (N_30950,N_25907,N_21500);
xor U30951 (N_30951,N_20421,N_27142);
nor U30952 (N_30952,N_29654,N_24790);
or U30953 (N_30953,N_24835,N_24974);
nor U30954 (N_30954,N_27645,N_23808);
or U30955 (N_30955,N_25442,N_27741);
nand U30956 (N_30956,N_23956,N_22204);
and U30957 (N_30957,N_29816,N_22273);
or U30958 (N_30958,N_27710,N_29473);
nand U30959 (N_30959,N_24142,N_26520);
or U30960 (N_30960,N_29099,N_25036);
nor U30961 (N_30961,N_24804,N_29343);
nor U30962 (N_30962,N_25945,N_25776);
nor U30963 (N_30963,N_27644,N_24943);
or U30964 (N_30964,N_25071,N_28617);
or U30965 (N_30965,N_22938,N_29344);
and U30966 (N_30966,N_26736,N_25691);
or U30967 (N_30967,N_26069,N_25388);
or U30968 (N_30968,N_21460,N_26976);
xnor U30969 (N_30969,N_28156,N_23141);
xnor U30970 (N_30970,N_22081,N_26519);
or U30971 (N_30971,N_26912,N_27604);
xnor U30972 (N_30972,N_23270,N_27157);
nor U30973 (N_30973,N_29244,N_23948);
or U30974 (N_30974,N_21297,N_28996);
and U30975 (N_30975,N_24553,N_28965);
or U30976 (N_30976,N_28463,N_25740);
xor U30977 (N_30977,N_28825,N_22059);
or U30978 (N_30978,N_23664,N_25139);
nand U30979 (N_30979,N_23174,N_23425);
nand U30980 (N_30980,N_20641,N_25001);
nor U30981 (N_30981,N_26925,N_26009);
nor U30982 (N_30982,N_25929,N_26075);
or U30983 (N_30983,N_24640,N_27724);
and U30984 (N_30984,N_27718,N_27391);
nand U30985 (N_30985,N_29878,N_29764);
and U30986 (N_30986,N_29924,N_20632);
or U30987 (N_30987,N_25764,N_23070);
nand U30988 (N_30988,N_27682,N_23302);
and U30989 (N_30989,N_23821,N_23340);
or U30990 (N_30990,N_27824,N_20194);
and U30991 (N_30991,N_21678,N_20487);
xnor U30992 (N_30992,N_29448,N_20017);
or U30993 (N_30993,N_25675,N_25160);
nor U30994 (N_30994,N_21149,N_26803);
nand U30995 (N_30995,N_21674,N_21205);
or U30996 (N_30996,N_22631,N_26919);
nand U30997 (N_30997,N_23733,N_24258);
and U30998 (N_30998,N_26689,N_28106);
and U30999 (N_30999,N_27333,N_22737);
nor U31000 (N_31000,N_29224,N_27891);
or U31001 (N_31001,N_22048,N_27527);
nor U31002 (N_31002,N_28131,N_29394);
nor U31003 (N_31003,N_21349,N_27713);
and U31004 (N_31004,N_22721,N_26262);
nand U31005 (N_31005,N_25554,N_21942);
and U31006 (N_31006,N_20567,N_20444);
nor U31007 (N_31007,N_20657,N_26690);
nor U31008 (N_31008,N_25958,N_29232);
xnor U31009 (N_31009,N_29447,N_25225);
or U31010 (N_31010,N_20408,N_29775);
and U31011 (N_31011,N_29523,N_23866);
nand U31012 (N_31012,N_29907,N_24162);
nor U31013 (N_31013,N_25098,N_27152);
and U31014 (N_31014,N_20334,N_20796);
nand U31015 (N_31015,N_22296,N_24666);
nor U31016 (N_31016,N_27349,N_26026);
nor U31017 (N_31017,N_20418,N_24816);
xnor U31018 (N_31018,N_20299,N_20426);
nor U31019 (N_31019,N_20537,N_23089);
or U31020 (N_31020,N_22090,N_23527);
and U31021 (N_31021,N_24194,N_22979);
nor U31022 (N_31022,N_28725,N_26824);
nand U31023 (N_31023,N_22848,N_23575);
or U31024 (N_31024,N_22393,N_23009);
or U31025 (N_31025,N_28838,N_27384);
and U31026 (N_31026,N_27321,N_25622);
or U31027 (N_31027,N_20863,N_23032);
nor U31028 (N_31028,N_24700,N_20986);
or U31029 (N_31029,N_28743,N_26796);
nand U31030 (N_31030,N_27441,N_27253);
or U31031 (N_31031,N_24264,N_22812);
nand U31032 (N_31032,N_24484,N_28801);
xnor U31033 (N_31033,N_22161,N_23386);
nor U31034 (N_31034,N_25099,N_28642);
nand U31035 (N_31035,N_22804,N_26959);
nand U31036 (N_31036,N_28077,N_26564);
nand U31037 (N_31037,N_26643,N_24043);
nand U31038 (N_31038,N_23451,N_23659);
nand U31039 (N_31039,N_21920,N_22698);
nor U31040 (N_31040,N_20488,N_24035);
nand U31041 (N_31041,N_29041,N_23643);
nand U31042 (N_31042,N_28536,N_22967);
nand U31043 (N_31043,N_27434,N_20615);
and U31044 (N_31044,N_28720,N_26290);
nor U31045 (N_31045,N_22887,N_20243);
and U31046 (N_31046,N_25856,N_20984);
and U31047 (N_31047,N_28620,N_28396);
or U31048 (N_31048,N_24821,N_27427);
nor U31049 (N_31049,N_29711,N_28120);
or U31050 (N_31050,N_26823,N_22029);
nor U31051 (N_31051,N_27219,N_28222);
and U31052 (N_31052,N_28745,N_29589);
nor U31053 (N_31053,N_24452,N_27181);
nand U31054 (N_31054,N_23485,N_27424);
and U31055 (N_31055,N_21816,N_26211);
nor U31056 (N_31056,N_20647,N_22611);
and U31057 (N_31057,N_23187,N_24605);
xnor U31058 (N_31058,N_28648,N_20280);
nand U31059 (N_31059,N_26722,N_26200);
nand U31060 (N_31060,N_25559,N_26781);
and U31061 (N_31061,N_24592,N_23071);
and U31062 (N_31062,N_29458,N_29320);
nor U31063 (N_31063,N_25156,N_23430);
nor U31064 (N_31064,N_21503,N_28944);
or U31065 (N_31065,N_21629,N_24355);
xnor U31066 (N_31066,N_23445,N_22265);
or U31067 (N_31067,N_24658,N_23043);
or U31068 (N_31068,N_21941,N_27487);
and U31069 (N_31069,N_27832,N_25792);
and U31070 (N_31070,N_28990,N_24239);
and U31071 (N_31071,N_27565,N_29865);
nor U31072 (N_31072,N_27979,N_21633);
nor U31073 (N_31073,N_22893,N_27558);
or U31074 (N_31074,N_25946,N_28193);
nor U31075 (N_31075,N_26348,N_25802);
nand U31076 (N_31076,N_21599,N_22241);
and U31077 (N_31077,N_27968,N_25450);
nand U31078 (N_31078,N_21560,N_22512);
nor U31079 (N_31079,N_24589,N_29054);
nor U31080 (N_31080,N_24010,N_22285);
or U31081 (N_31081,N_25466,N_27492);
and U31082 (N_31082,N_23928,N_24895);
nand U31083 (N_31083,N_20255,N_23145);
and U31084 (N_31084,N_25410,N_23826);
xor U31085 (N_31085,N_21326,N_22038);
or U31086 (N_31086,N_24055,N_22343);
or U31087 (N_31087,N_29222,N_20795);
or U31088 (N_31088,N_21621,N_24961);
and U31089 (N_31089,N_26687,N_21265);
or U31090 (N_31090,N_26691,N_24430);
nand U31091 (N_31091,N_22338,N_23183);
xor U31092 (N_31092,N_21606,N_20475);
and U31093 (N_31093,N_28763,N_25143);
or U31094 (N_31094,N_21374,N_24763);
nor U31095 (N_31095,N_29607,N_27906);
and U31096 (N_31096,N_25586,N_28078);
and U31097 (N_31097,N_22897,N_26741);
or U31098 (N_31098,N_23633,N_20290);
nor U31099 (N_31099,N_26377,N_28956);
xnor U31100 (N_31100,N_26241,N_23833);
xnor U31101 (N_31101,N_27569,N_25060);
nand U31102 (N_31102,N_22536,N_29165);
nor U31103 (N_31103,N_27339,N_24905);
nand U31104 (N_31104,N_28717,N_21835);
nand U31105 (N_31105,N_21380,N_25024);
nor U31106 (N_31106,N_23966,N_25183);
and U31107 (N_31107,N_22261,N_22375);
nor U31108 (N_31108,N_27238,N_27507);
nor U31109 (N_31109,N_24197,N_24279);
or U31110 (N_31110,N_29573,N_24881);
or U31111 (N_31111,N_20857,N_21148);
or U31112 (N_31112,N_24072,N_25461);
nand U31113 (N_31113,N_22479,N_23321);
or U31114 (N_31114,N_20597,N_28778);
nand U31115 (N_31115,N_24902,N_29548);
or U31116 (N_31116,N_26518,N_29528);
or U31117 (N_31117,N_28091,N_20554);
nor U31118 (N_31118,N_28117,N_22162);
nand U31119 (N_31119,N_23476,N_23662);
and U31120 (N_31120,N_23102,N_20405);
xor U31121 (N_31121,N_28945,N_22772);
nor U31122 (N_31122,N_25744,N_28844);
nand U31123 (N_31123,N_23223,N_23154);
nand U31124 (N_31124,N_29491,N_22249);
or U31125 (N_31125,N_29154,N_20079);
xor U31126 (N_31126,N_27878,N_21352);
or U31127 (N_31127,N_29556,N_28841);
or U31128 (N_31128,N_26960,N_21005);
nand U31129 (N_31129,N_27263,N_28126);
nand U31130 (N_31130,N_20298,N_29502);
and U31131 (N_31131,N_20794,N_27477);
nor U31132 (N_31132,N_29022,N_24988);
nor U31133 (N_31133,N_20398,N_22202);
nand U31134 (N_31134,N_23246,N_24796);
nor U31135 (N_31135,N_22392,N_29162);
and U31136 (N_31136,N_25798,N_25647);
and U31137 (N_31137,N_28359,N_26598);
nor U31138 (N_31138,N_28287,N_23590);
and U31139 (N_31139,N_28897,N_23244);
and U31140 (N_31140,N_20023,N_23690);
nand U31141 (N_31141,N_20495,N_22279);
nor U31142 (N_31142,N_24465,N_26804);
nand U31143 (N_31143,N_22233,N_22920);
and U31144 (N_31144,N_29636,N_22661);
or U31145 (N_31145,N_27937,N_25652);
or U31146 (N_31146,N_26479,N_26394);
and U31147 (N_31147,N_20757,N_27250);
nor U31148 (N_31148,N_27658,N_26735);
or U31149 (N_31149,N_21248,N_26419);
and U31150 (N_31150,N_25073,N_22774);
nand U31151 (N_31151,N_29088,N_20650);
or U31152 (N_31152,N_21058,N_23558);
nor U31153 (N_31153,N_23120,N_28650);
xor U31154 (N_31154,N_28649,N_25841);
and U31155 (N_31155,N_23158,N_21667);
nor U31156 (N_31156,N_29596,N_23666);
xnor U31157 (N_31157,N_22318,N_26957);
nand U31158 (N_31158,N_23044,N_24698);
or U31159 (N_31159,N_26225,N_25735);
and U31160 (N_31160,N_25663,N_26020);
or U31161 (N_31161,N_22852,N_28851);
or U31162 (N_31162,N_27345,N_24085);
or U31163 (N_31163,N_23514,N_28978);
nor U31164 (N_31164,N_26865,N_28541);
or U31165 (N_31165,N_23746,N_20077);
or U31166 (N_31166,N_28003,N_24759);
and U31167 (N_31167,N_21379,N_21594);
nand U31168 (N_31168,N_21366,N_28980);
nand U31169 (N_31169,N_26550,N_29701);
nor U31170 (N_31170,N_24714,N_22608);
nor U31171 (N_31171,N_20903,N_21208);
xor U31172 (N_31172,N_20449,N_23609);
nand U31173 (N_31173,N_21325,N_20306);
and U31174 (N_31174,N_28527,N_26789);
nand U31175 (N_31175,N_25601,N_20699);
xnor U31176 (N_31176,N_24722,N_25112);
or U31177 (N_31177,N_22974,N_28712);
or U31178 (N_31178,N_25202,N_21976);
or U31179 (N_31179,N_27172,N_27998);
and U31180 (N_31180,N_20374,N_29742);
and U31181 (N_31181,N_25679,N_26461);
nor U31182 (N_31182,N_23253,N_26822);
or U31183 (N_31183,N_27525,N_27888);
nor U31184 (N_31184,N_22489,N_24524);
nand U31185 (N_31185,N_26181,N_29687);
xnor U31186 (N_31186,N_26359,N_29410);
and U31187 (N_31187,N_20213,N_27104);
xnor U31188 (N_31188,N_25234,N_23681);
nand U31189 (N_31189,N_28799,N_27506);
nor U31190 (N_31190,N_27758,N_20676);
nand U31191 (N_31191,N_23061,N_27029);
or U31192 (N_31192,N_27022,N_29411);
or U31193 (N_31193,N_25810,N_24650);
nor U31194 (N_31194,N_21535,N_24627);
nand U31195 (N_31195,N_24500,N_24748);
or U31196 (N_31196,N_20326,N_23692);
nor U31197 (N_31197,N_26064,N_26309);
and U31198 (N_31198,N_28008,N_27866);
nand U31199 (N_31199,N_28258,N_21189);
or U31200 (N_31200,N_29897,N_22043);
xor U31201 (N_31201,N_27531,N_21443);
and U31202 (N_31202,N_26464,N_22101);
nor U31203 (N_31203,N_21397,N_28462);
nand U31204 (N_31204,N_27256,N_27744);
and U31205 (N_31205,N_29121,N_26816);
and U31206 (N_31206,N_25784,N_23418);
or U31207 (N_31207,N_23448,N_24669);
or U31208 (N_31208,N_29854,N_21588);
or U31209 (N_31209,N_21888,N_25645);
nor U31210 (N_31210,N_28847,N_29347);
and U31211 (N_31211,N_27996,N_27624);
nand U31212 (N_31212,N_20519,N_21540);
and U31213 (N_31213,N_25819,N_24408);
xnor U31214 (N_31214,N_25352,N_28794);
xnor U31215 (N_31215,N_29201,N_26731);
and U31216 (N_31216,N_23854,N_22767);
nor U31217 (N_31217,N_23136,N_26654);
nand U31218 (N_31218,N_29542,N_26674);
nand U31219 (N_31219,N_29641,N_21945);
nand U31220 (N_31220,N_28580,N_24696);
or U31221 (N_31221,N_26616,N_26831);
nor U31222 (N_31222,N_24678,N_21999);
or U31223 (N_31223,N_22937,N_23906);
or U31224 (N_31224,N_26109,N_22465);
nand U31225 (N_31225,N_22833,N_25010);
nor U31226 (N_31226,N_24158,N_20456);
nor U31227 (N_31227,N_21097,N_23743);
and U31228 (N_31228,N_27207,N_20691);
and U31229 (N_31229,N_25718,N_23432);
and U31230 (N_31230,N_22281,N_24045);
xnor U31231 (N_31231,N_21361,N_26979);
and U31232 (N_31232,N_28426,N_29706);
xnor U31233 (N_31233,N_20416,N_20086);
nand U31234 (N_31234,N_23852,N_20071);
nand U31235 (N_31235,N_25011,N_20891);
xor U31236 (N_31236,N_20124,N_28441);
or U31237 (N_31237,N_21172,N_27611);
nor U31238 (N_31238,N_20231,N_26697);
nor U31239 (N_31239,N_28817,N_20403);
nor U31240 (N_31240,N_20156,N_25570);
nand U31241 (N_31241,N_29451,N_24888);
nand U31242 (N_31242,N_22427,N_26371);
nand U31243 (N_31243,N_24999,N_23110);
nand U31244 (N_31244,N_29255,N_20902);
xnor U31245 (N_31245,N_26688,N_24809);
and U31246 (N_31246,N_24917,N_26275);
nor U31247 (N_31247,N_28632,N_29003);
nand U31248 (N_31248,N_23411,N_25298);
nand U31249 (N_31249,N_22299,N_28262);
nand U31250 (N_31250,N_27050,N_29148);
and U31251 (N_31251,N_29132,N_25626);
nand U31252 (N_31252,N_26054,N_27582);
nor U31253 (N_31253,N_28552,N_28154);
or U31254 (N_31254,N_21602,N_29001);
and U31255 (N_31255,N_20779,N_25390);
or U31256 (N_31256,N_27992,N_21849);
or U31257 (N_31257,N_26083,N_22123);
or U31258 (N_31258,N_25761,N_29642);
nand U31259 (N_31259,N_23711,N_27222);
nand U31260 (N_31260,N_26501,N_23559);
and U31261 (N_31261,N_24535,N_28921);
nor U31262 (N_31262,N_23504,N_26182);
or U31263 (N_31263,N_27728,N_22418);
nand U31264 (N_31264,N_25523,N_29490);
nor U31265 (N_31265,N_28206,N_28654);
nor U31266 (N_31266,N_26765,N_25017);
nor U31267 (N_31267,N_22412,N_23788);
nand U31268 (N_31268,N_28684,N_22147);
and U31269 (N_31269,N_29718,N_25860);
or U31270 (N_31270,N_20066,N_25375);
xor U31271 (N_31271,N_21968,N_24322);
or U31272 (N_31272,N_26574,N_26242);
nor U31273 (N_31273,N_21047,N_29595);
and U31274 (N_31274,N_22165,N_28953);
and U31275 (N_31275,N_20341,N_25286);
nand U31276 (N_31276,N_26058,N_29492);
or U31277 (N_31277,N_26232,N_21185);
nand U31278 (N_31278,N_25888,N_27925);
nor U31279 (N_31279,N_20521,N_21591);
or U31280 (N_31280,N_28057,N_29428);
nand U31281 (N_31281,N_24645,N_20608);
nor U31282 (N_31282,N_23354,N_22935);
xnor U31283 (N_31283,N_27779,N_20220);
nor U31284 (N_31284,N_26406,N_26081);
or U31285 (N_31285,N_20876,N_21981);
nand U31286 (N_31286,N_24097,N_22677);
or U31287 (N_31287,N_23034,N_25432);
or U31288 (N_31288,N_22128,N_26523);
nor U31289 (N_31289,N_22624,N_23237);
and U31290 (N_31290,N_27180,N_21960);
and U31291 (N_31291,N_22175,N_22220);
nand U31292 (N_31292,N_26169,N_27733);
and U31293 (N_31293,N_24240,N_27887);
nor U31294 (N_31294,N_29273,N_28785);
and U31295 (N_31295,N_25397,N_21049);
nor U31296 (N_31296,N_27872,N_24336);
or U31297 (N_31297,N_22626,N_29112);
nand U31298 (N_31298,N_22751,N_27904);
nand U31299 (N_31299,N_29946,N_23568);
or U31300 (N_31300,N_20988,N_24041);
and U31301 (N_31301,N_24171,N_27813);
nand U31302 (N_31302,N_25012,N_23433);
or U31303 (N_31303,N_20706,N_22291);
or U31304 (N_31304,N_23717,N_27124);
and U31305 (N_31305,N_29067,N_22549);
nor U31306 (N_31306,N_21431,N_24981);
nand U31307 (N_31307,N_21759,N_21786);
nand U31308 (N_31308,N_22268,N_22277);
nor U31309 (N_31309,N_24569,N_22409);
nand U31310 (N_31310,N_26606,N_26720);
xor U31311 (N_31311,N_20168,N_24375);
xnor U31312 (N_31312,N_26179,N_29313);
or U31313 (N_31313,N_22495,N_23058);
xnor U31314 (N_31314,N_26283,N_26440);
nand U31315 (N_31315,N_25906,N_22883);
nand U31316 (N_31316,N_28357,N_26382);
nand U31317 (N_31317,N_23718,N_23081);
nand U31318 (N_31318,N_21237,N_25831);
nand U31319 (N_31319,N_27643,N_24749);
or U31320 (N_31320,N_27771,N_22911);
nand U31321 (N_31321,N_24586,N_29670);
or U31322 (N_31322,N_29472,N_22599);
or U31323 (N_31323,N_28253,N_20960);
nand U31324 (N_31324,N_20888,N_20482);
nand U31325 (N_31325,N_26364,N_20065);
or U31326 (N_31326,N_22506,N_23941);
nand U31327 (N_31327,N_24022,N_28271);
and U31328 (N_31328,N_28750,N_27627);
nand U31329 (N_31329,N_24402,N_24693);
nand U31330 (N_31330,N_24836,N_28899);
nor U31331 (N_31331,N_28015,N_25820);
nand U31332 (N_31332,N_26651,N_27281);
or U31333 (N_31333,N_28440,N_23007);
xnor U31334 (N_31334,N_20703,N_28973);
nor U31335 (N_31335,N_25673,N_24467);
and U31336 (N_31336,N_29253,N_20958);
nand U31337 (N_31337,N_26124,N_24418);
nor U31338 (N_31338,N_25027,N_24482);
nand U31339 (N_31339,N_27513,N_23400);
or U31340 (N_31340,N_25088,N_23598);
or U31341 (N_31341,N_23143,N_24312);
and U31342 (N_31342,N_20602,N_29365);
xnor U31343 (N_31343,N_28321,N_29861);
nor U31344 (N_31344,N_29316,N_23919);
and U31345 (N_31345,N_25141,N_26138);
nand U31346 (N_31346,N_26622,N_22461);
nand U31347 (N_31347,N_20906,N_26562);
and U31348 (N_31348,N_26481,N_23101);
nor U31349 (N_31349,N_21497,N_21676);
nand U31350 (N_31350,N_29060,N_25534);
and U31351 (N_31351,N_20561,N_29206);
and U31352 (N_31352,N_24741,N_25434);
and U31353 (N_31353,N_28168,N_24774);
and U31354 (N_31354,N_27421,N_23785);
or U31355 (N_31355,N_27030,N_29998);
nor U31356 (N_31356,N_26845,N_29866);
or U31357 (N_31357,N_26663,N_25506);
nand U31358 (N_31358,N_29286,N_27276);
and U31359 (N_31359,N_24690,N_22861);
or U31360 (N_31360,N_24598,N_28766);
nor U31361 (N_31361,N_20201,N_22385);
nor U31362 (N_31362,N_20376,N_26999);
nand U31363 (N_31363,N_29256,N_25093);
nor U31364 (N_31364,N_23972,N_29103);
and U31365 (N_31365,N_26427,N_23952);
or U31366 (N_31366,N_21982,N_29799);
nand U31367 (N_31367,N_26980,N_21872);
nand U31368 (N_31368,N_26061,N_23538);
and U31369 (N_31369,N_22988,N_20005);
and U31370 (N_31370,N_21807,N_23254);
xnor U31371 (N_31371,N_28700,N_29207);
nor U31372 (N_31372,N_27026,N_23938);
or U31373 (N_31373,N_21283,N_21557);
nand U31374 (N_31374,N_28448,N_21159);
and U31375 (N_31375,N_24017,N_28352);
or U31376 (N_31376,N_26476,N_24246);
and U31377 (N_31377,N_22847,N_24670);
nand U31378 (N_31378,N_22971,N_24728);
or U31379 (N_31379,N_27415,N_27360);
nand U31380 (N_31380,N_28337,N_23283);
or U31381 (N_31381,N_24661,N_29766);
nand U31382 (N_31382,N_23293,N_29114);
and U31383 (N_31383,N_25890,N_21697);
nor U31384 (N_31384,N_25706,N_21449);
and U31385 (N_31385,N_27910,N_20672);
and U31386 (N_31386,N_28843,N_21634);
or U31387 (N_31387,N_27317,N_21954);
or U31388 (N_31388,N_20717,N_22188);
or U31389 (N_31389,N_23780,N_26638);
and U31390 (N_31390,N_24721,N_24117);
and U31391 (N_31391,N_20811,N_25111);
and U31392 (N_31392,N_22042,N_26227);
nor U31393 (N_31393,N_28633,N_29193);
and U31394 (N_31394,N_21515,N_23663);
nand U31395 (N_31395,N_20843,N_27618);
or U31396 (N_31396,N_21282,N_25464);
or U31397 (N_31397,N_26879,N_24252);
or U31398 (N_31398,N_25618,N_29226);
and U31399 (N_31399,N_23397,N_23510);
and U31400 (N_31400,N_24308,N_24924);
or U31401 (N_31401,N_22382,N_24276);
and U31402 (N_31402,N_24512,N_24436);
nand U31403 (N_31403,N_25274,N_29141);
or U31404 (N_31404,N_23697,N_29515);
xnor U31405 (N_31405,N_21879,N_28009);
or U31406 (N_31406,N_23767,N_26177);
or U31407 (N_31407,N_29034,N_20366);
xnor U31408 (N_31408,N_28554,N_27539);
and U31409 (N_31409,N_29512,N_20393);
or U31410 (N_31410,N_21173,N_20193);
nor U31411 (N_31411,N_24288,N_27137);
or U31412 (N_31412,N_22740,N_29305);
and U31413 (N_31413,N_27056,N_24009);
nor U31414 (N_31414,N_21803,N_20229);
and U31415 (N_31415,N_27000,N_22610);
xnor U31416 (N_31416,N_23874,N_22478);
or U31417 (N_31417,N_21304,N_25943);
xor U31418 (N_31418,N_24146,N_21118);
or U31419 (N_31419,N_26759,N_24313);
or U31420 (N_31420,N_28952,N_23677);
nand U31421 (N_31421,N_25777,N_24196);
nand U31422 (N_31422,N_27672,N_20677);
nand U31423 (N_31423,N_26230,N_21777);
and U31424 (N_31424,N_20172,N_23507);
or U31425 (N_31425,N_27202,N_23222);
and U31426 (N_31426,N_25807,N_27457);
and U31427 (N_31427,N_24238,N_23776);
xor U31428 (N_31428,N_22648,N_26034);
and U31429 (N_31429,N_26872,N_29322);
and U31430 (N_31430,N_27958,N_25648);
xor U31431 (N_31431,N_26048,N_21126);
nand U31432 (N_31432,N_22085,N_25869);
nand U31433 (N_31433,N_27381,N_27126);
or U31434 (N_31434,N_29238,N_21457);
or U31435 (N_31435,N_27098,N_29486);
or U31436 (N_31436,N_27542,N_29981);
xor U31437 (N_31437,N_27483,N_25788);
nand U31438 (N_31438,N_23572,N_20603);
nor U31439 (N_31439,N_27665,N_27261);
nor U31440 (N_31440,N_21900,N_29470);
or U31441 (N_31441,N_25630,N_24976);
and U31442 (N_31442,N_28467,N_25854);
nand U31443 (N_31443,N_29814,N_20508);
or U31444 (N_31444,N_29560,N_22315);
and U31445 (N_31445,N_26793,N_24689);
nor U31446 (N_31446,N_21392,N_24713);
nor U31447 (N_31447,N_29252,N_24538);
and U31448 (N_31448,N_27252,N_23975);
xor U31449 (N_31449,N_27812,N_28868);
or U31450 (N_31450,N_23577,N_29386);
or U31451 (N_31451,N_25690,N_28304);
nand U31452 (N_31452,N_21227,N_26723);
and U31453 (N_31453,N_23375,N_29883);
or U31454 (N_31454,N_24215,N_21513);
and U31455 (N_31455,N_27545,N_26711);
and U31456 (N_31456,N_25387,N_22439);
nor U31457 (N_31457,N_23554,N_22530);
nor U31458 (N_31458,N_28934,N_21804);
or U31459 (N_31459,N_28225,N_22408);
nand U31460 (N_31460,N_24868,N_20810);
nand U31461 (N_31461,N_20694,N_27880);
xor U31462 (N_31462,N_21554,N_24514);
nand U31463 (N_31463,N_22831,N_27587);
or U31464 (N_31464,N_29249,N_25876);
nand U31465 (N_31465,N_28503,N_26014);
or U31466 (N_31466,N_24772,N_24198);
or U31467 (N_31467,N_27099,N_27068);
nand U31468 (N_31468,N_22026,N_28969);
nand U31469 (N_31469,N_29172,N_28421);
nor U31470 (N_31470,N_20246,N_28608);
and U31471 (N_31471,N_23638,N_27893);
and U31472 (N_31472,N_29385,N_24399);
nand U31473 (N_31473,N_22144,N_22192);
or U31474 (N_31474,N_28754,N_28951);
or U31475 (N_31475,N_22351,N_25067);
nand U31476 (N_31476,N_26101,N_24388);
nand U31477 (N_31477,N_22324,N_23683);
and U31478 (N_31478,N_27523,N_21245);
nand U31479 (N_31479,N_23971,N_24318);
nor U31480 (N_31480,N_26391,N_25220);
nor U31481 (N_31481,N_28113,N_24119);
nand U31482 (N_31482,N_27264,N_20039);
nand U31483 (N_31483,N_20138,N_28458);
nand U31484 (N_31484,N_21766,N_27915);
nand U31485 (N_31485,N_25762,N_23142);
or U31486 (N_31486,N_22064,N_23661);
nor U31487 (N_31487,N_20284,N_28874);
or U31488 (N_31488,N_26196,N_20879);
or U31489 (N_31489,N_25614,N_22678);
nand U31490 (N_31490,N_20044,N_20791);
nor U31491 (N_31491,N_25287,N_23535);
nor U31492 (N_31492,N_28016,N_27786);
nor U31493 (N_31493,N_27480,N_26415);
nor U31494 (N_31494,N_27277,N_24189);
or U31495 (N_31495,N_29966,N_27568);
nor U31496 (N_31496,N_27695,N_21295);
xnor U31497 (N_31497,N_27190,N_20587);
or U31498 (N_31498,N_20913,N_25360);
nand U31499 (N_31499,N_26132,N_24573);
or U31500 (N_31500,N_26991,N_29283);
or U31501 (N_31501,N_23858,N_25215);
nand U31502 (N_31502,N_28774,N_22695);
nor U31503 (N_31503,N_22504,N_27882);
or U31504 (N_31504,N_26594,N_29011);
or U31505 (N_31505,N_28384,N_23039);
and U31506 (N_31506,N_27969,N_22527);
and U31507 (N_31507,N_27902,N_21157);
xor U31508 (N_31508,N_24473,N_24975);
or U31509 (N_31509,N_27092,N_25203);
or U31510 (N_31510,N_28324,N_29842);
nand U31511 (N_31511,N_22011,N_23266);
or U31512 (N_31512,N_22404,N_22118);
or U31513 (N_31513,N_26474,N_25422);
nor U31514 (N_31514,N_28007,N_28932);
xor U31515 (N_31515,N_23770,N_24109);
and U31516 (N_31516,N_20511,N_26155);
nor U31517 (N_31517,N_21800,N_21539);
nor U31518 (N_31518,N_23064,N_22687);
or U31519 (N_31519,N_26434,N_29736);
xor U31520 (N_31520,N_29049,N_22980);
or U31521 (N_31521,N_22598,N_29885);
and U31522 (N_31522,N_29737,N_24614);
nand U31523 (N_31523,N_27399,N_29004);
and U31524 (N_31524,N_22380,N_22340);
nor U31525 (N_31525,N_24600,N_29621);
and U31526 (N_31526,N_27340,N_20839);
nand U31527 (N_31527,N_21776,N_29896);
and U31528 (N_31528,N_24113,N_28174);
nor U31529 (N_31529,N_24760,N_29300);
nand U31530 (N_31530,N_20762,N_29214);
or U31531 (N_31531,N_23829,N_24874);
and U31532 (N_31532,N_23149,N_29768);
or U31533 (N_31533,N_23170,N_22790);
nand U31534 (N_31534,N_24139,N_24813);
and U31535 (N_31535,N_28399,N_20838);
nand U31536 (N_31536,N_24582,N_28336);
and U31537 (N_31537,N_28255,N_23524);
nor U31538 (N_31538,N_26572,N_26908);
or U31539 (N_31539,N_24186,N_23168);
or U31540 (N_31540,N_26978,N_24739);
and U31541 (N_31541,N_23750,N_20543);
nand U31542 (N_31542,N_28149,N_25374);
or U31543 (N_31543,N_20821,N_27726);
nor U31544 (N_31544,N_21102,N_24199);
xnor U31545 (N_31545,N_27614,N_23038);
nand U31546 (N_31546,N_25431,N_28322);
nand U31547 (N_31547,N_23629,N_28012);
nor U31548 (N_31548,N_23495,N_23842);
nand U31549 (N_31549,N_27526,N_24707);
or U31550 (N_31550,N_27299,N_20992);
and U31551 (N_31551,N_22649,N_24409);
xor U31552 (N_31552,N_22019,N_26125);
and U31553 (N_31553,N_20565,N_25686);
nand U31554 (N_31554,N_25325,N_28918);
and U31555 (N_31555,N_22061,N_20707);
xnor U31556 (N_31556,N_24986,N_21171);
and U31557 (N_31557,N_29277,N_21919);
nand U31558 (N_31558,N_25653,N_25219);
nor U31559 (N_31559,N_21350,N_20209);
and U31560 (N_31560,N_28857,N_22484);
nand U31561 (N_31561,N_24697,N_28484);
nor U31562 (N_31562,N_24860,N_26305);
nand U31563 (N_31563,N_20846,N_25795);
and U31564 (N_31564,N_27540,N_28575);
xnor U31565 (N_31565,N_20462,N_25833);
nand U31566 (N_31566,N_28111,N_25911);
or U31567 (N_31567,N_23908,N_29858);
nand U31568 (N_31568,N_27128,N_29187);
nor U31569 (N_31569,N_29169,N_24455);
and U31570 (N_31570,N_22415,N_26448);
nand U31571 (N_31571,N_21076,N_22337);
xor U31572 (N_31572,N_27301,N_20975);
or U31573 (N_31573,N_20045,N_24468);
nand U31574 (N_31574,N_23265,N_22680);
nand U31575 (N_31575,N_26247,N_21272);
nor U31576 (N_31576,N_28275,N_20303);
nand U31577 (N_31577,N_20895,N_23636);
or U31578 (N_31578,N_25927,N_22764);
and U31579 (N_31579,N_29023,N_21156);
and U31580 (N_31580,N_29000,N_24959);
xnor U31581 (N_31581,N_23057,N_26004);
nand U31582 (N_31582,N_23290,N_23267);
and U31583 (N_31583,N_22158,N_22987);
nor U31584 (N_31584,N_26123,N_27773);
nand U31585 (N_31585,N_20208,N_21482);
nor U31586 (N_31586,N_23473,N_25046);
nand U31587 (N_31587,N_26190,N_22227);
nand U31588 (N_31588,N_28915,N_29845);
nor U31589 (N_31589,N_24440,N_22084);
or U31590 (N_31590,N_20639,N_25180);
nor U31591 (N_31591,N_27064,N_21532);
and U31592 (N_31592,N_27808,N_22219);
and U31593 (N_31593,N_26416,N_28349);
and U31594 (N_31594,N_27169,N_22964);
or U31595 (N_31595,N_20931,N_27471);
or U31596 (N_31596,N_21992,N_21881);
nor U31597 (N_31597,N_27676,N_26153);
or U31598 (N_31598,N_23668,N_21604);
nor U31599 (N_31599,N_23859,N_28656);
nand U31600 (N_31600,N_27809,N_29530);
nor U31601 (N_31601,N_22169,N_27034);
and U31602 (N_31602,N_22293,N_22377);
nand U31603 (N_31603,N_27524,N_25755);
or U31604 (N_31604,N_21014,N_22150);
xor U31605 (N_31605,N_26051,N_27919);
or U31606 (N_31606,N_21386,N_22130);
and U31607 (N_31607,N_28392,N_23903);
and U31608 (N_31608,N_22703,N_25400);
or U31609 (N_31609,N_22707,N_27435);
nand U31610 (N_31610,N_26782,N_28722);
xor U31611 (N_31611,N_29495,N_24153);
nor U31612 (N_31612,N_21596,N_27209);
nand U31613 (N_31613,N_21229,N_29519);
or U31614 (N_31614,N_20827,N_22706);
xnor U31615 (N_31615,N_23460,N_24558);
and U31616 (N_31616,N_29909,N_23761);
and U31617 (N_31617,N_28150,N_26270);
nand U31618 (N_31618,N_23393,N_23004);
nand U31619 (N_31619,N_24268,N_20783);
nor U31620 (N_31620,N_25123,N_20591);
nor U31621 (N_31621,N_22856,N_26967);
nor U31622 (N_31622,N_29483,N_27075);
nor U31623 (N_31623,N_25899,N_20447);
or U31624 (N_31624,N_24385,N_29604);
nor U31625 (N_31625,N_28098,N_25486);
or U31626 (N_31626,N_22781,N_28583);
xor U31627 (N_31627,N_23021,N_25983);
xnor U31628 (N_31628,N_25689,N_20125);
or U31629 (N_31629,N_24302,N_23515);
xnor U31630 (N_31630,N_29815,N_28192);
nor U31631 (N_31631,N_24886,N_21357);
and U31632 (N_31632,N_23403,N_23420);
nand U31633 (N_31633,N_24997,N_27534);
xnor U31634 (N_31634,N_21692,N_25000);
or U31635 (N_31635,N_29500,N_23931);
and U31636 (N_31636,N_28449,N_22070);
nand U31637 (N_31637,N_29882,N_22780);
nand U31638 (N_31638,N_29336,N_23167);
nor U31639 (N_31639,N_28815,N_26982);
xor U31640 (N_31640,N_26176,N_25369);
or U31641 (N_31641,N_24726,N_22232);
nor U31642 (N_31642,N_20318,N_25176);
or U31643 (N_31643,N_26395,N_24138);
nand U31644 (N_31644,N_25678,N_26094);
nor U31645 (N_31645,N_24144,N_21829);
or U31646 (N_31646,N_27350,N_25013);
nor U31647 (N_31647,N_26147,N_26677);
and U31648 (N_31648,N_26202,N_24889);
or U31649 (N_31649,N_23867,N_22441);
or U31650 (N_31650,N_21371,N_27541);
nand U31651 (N_31651,N_25770,N_27417);
nand U31652 (N_31652,N_23694,N_29971);
xnor U31653 (N_31653,N_23013,N_20735);
and U31654 (N_31654,N_27518,N_22016);
nand U31655 (N_31655,N_20940,N_22923);
and U31656 (N_31656,N_27155,N_24251);
or U31657 (N_31657,N_24852,N_22982);
and U31658 (N_31658,N_20116,N_21852);
nand U31659 (N_31659,N_27062,N_24241);
or U31660 (N_31660,N_28415,N_20844);
and U31661 (N_31661,N_25382,N_28498);
nand U31662 (N_31662,N_22221,N_24516);
nor U31663 (N_31663,N_25632,N_29967);
and U31664 (N_31664,N_29752,N_25967);
or U31665 (N_31665,N_22745,N_24606);
and U31666 (N_31666,N_24546,N_23625);
nor U31667 (N_31667,N_26302,N_21220);
nand U31668 (N_31668,N_20414,N_24919);
nor U31669 (N_31669,N_21758,N_25207);
nand U31670 (N_31670,N_25971,N_21454);
nand U31671 (N_31671,N_20656,N_26120);
nand U31672 (N_31672,N_20774,N_22681);
nor U31673 (N_31673,N_26992,N_28993);
xnor U31674 (N_31674,N_27021,N_28017);
or U31675 (N_31675,N_25223,N_24541);
xor U31676 (N_31676,N_25604,N_21333);
or U31677 (N_31677,N_21823,N_23974);
and U31678 (N_31678,N_25608,N_24768);
or U31679 (N_31679,N_28473,N_23921);
or U31680 (N_31680,N_29390,N_27997);
or U31681 (N_31681,N_27512,N_26806);
nor U31682 (N_31682,N_23307,N_27337);
nand U31683 (N_31683,N_28439,N_28429);
nor U31684 (N_31684,N_28539,N_21940);
xor U31685 (N_31685,N_22800,N_27859);
and U31686 (N_31686,N_24298,N_21850);
nor U31687 (N_31687,N_21628,N_24936);
xnor U31688 (N_31688,N_26624,N_29424);
nor U31689 (N_31689,N_29574,N_22131);
and U31690 (N_31690,N_26748,N_28143);
and U31691 (N_31691,N_24290,N_29312);
xor U31692 (N_31692,N_29509,N_23126);
nand U31693 (N_31693,N_26535,N_27482);
nor U31694 (N_31694,N_24335,N_29785);
and U31695 (N_31695,N_26997,N_23224);
and U31696 (N_31696,N_24636,N_25791);
or U31697 (N_31697,N_22630,N_26465);
or U31698 (N_31698,N_29263,N_27184);
nor U31699 (N_31699,N_26920,N_25395);
nand U31700 (N_31700,N_26993,N_23160);
nand U31701 (N_31701,N_29557,N_22251);
or U31702 (N_31702,N_22702,N_22234);
nand U31703 (N_31703,N_28593,N_23706);
and U31704 (N_31704,N_21884,N_26053);
or U31705 (N_31705,N_23885,N_25756);
nand U31706 (N_31706,N_24618,N_24262);
xnor U31707 (N_31707,N_27530,N_27431);
nand U31708 (N_31708,N_29427,N_22685);
nand U31709 (N_31709,N_28061,N_21060);
xor U31710 (N_31710,N_25668,N_24459);
nor U31711 (N_31711,N_23159,N_27564);
and U31712 (N_31712,N_21434,N_27649);
nor U31713 (N_31713,N_23015,N_22584);
xor U31714 (N_31714,N_22995,N_20532);
nand U31715 (N_31715,N_28890,N_25433);
nand U31716 (N_31716,N_26329,N_20845);
nor U31717 (N_31717,N_28948,N_22786);
nand U31718 (N_31718,N_21343,N_25928);
or U31719 (N_31719,N_25104,N_24479);
or U31720 (N_31720,N_25739,N_27677);
nor U31721 (N_31721,N_21015,N_24890);
and U31722 (N_31722,N_28329,N_24018);
nor U31723 (N_31723,N_29113,N_20785);
or U31724 (N_31724,N_29972,N_22959);
nor U31725 (N_31725,N_21712,N_20224);
nor U31726 (N_31726,N_22423,N_20109);
xnor U31727 (N_31727,N_23765,N_24330);
or U31728 (N_31728,N_23865,N_21901);
nand U31729 (N_31729,N_29246,N_20262);
nor U31730 (N_31730,N_20361,N_29029);
xor U31731 (N_31731,N_23843,N_27121);
or U31732 (N_31732,N_21866,N_25295);
and U31733 (N_31733,N_27266,N_29128);
nand U31734 (N_31734,N_26257,N_28409);
nand U31735 (N_31735,N_24098,N_22284);
nor U31736 (N_31736,N_29712,N_23055);
or U31737 (N_31737,N_21468,N_29350);
or U31738 (N_31738,N_21123,N_22089);
nor U31739 (N_31739,N_20688,N_24780);
xnor U31740 (N_31740,N_22881,N_25467);
or U31741 (N_31741,N_25612,N_28491);
or U31742 (N_31742,N_23648,N_27361);
and U31743 (N_31743,N_27535,N_28430);
nand U31744 (N_31744,N_27792,N_28728);
nand U31745 (N_31745,N_24688,N_24116);
and U31746 (N_31746,N_24254,N_29617);
and U31747 (N_31747,N_22483,N_25378);
nand U31748 (N_31748,N_23803,N_27723);
nor U31749 (N_31749,N_22317,N_20238);
nand U31750 (N_31750,N_27084,N_28354);
nand U31751 (N_31751,N_27953,N_20594);
xor U31752 (N_31752,N_23190,N_28320);
nor U31753 (N_31753,N_20817,N_25448);
nor U31754 (N_31754,N_25794,N_26578);
nand U31755 (N_31755,N_29786,N_26617);
xor U31756 (N_31756,N_25696,N_20049);
nor U31757 (N_31757,N_22612,N_29702);
nand U31758 (N_31758,N_24212,N_27150);
nor U31759 (N_31759,N_23913,N_23660);
and U31760 (N_31760,N_22822,N_25069);
or U31761 (N_31761,N_24621,N_26770);
nor U31762 (N_31762,N_26159,N_22915);
or U31763 (N_31763,N_26554,N_22207);
or U31764 (N_31764,N_23642,N_22159);
or U31765 (N_31765,N_24995,N_27720);
nor U31766 (N_31766,N_26650,N_29337);
or U31767 (N_31767,N_23324,N_22670);
and U31768 (N_31768,N_26121,N_21081);
nor U31769 (N_31769,N_20093,N_26629);
nand U31770 (N_31770,N_29531,N_27563);
nand U31771 (N_31771,N_25625,N_20809);
xor U31772 (N_31772,N_25778,N_20512);
and U31773 (N_31773,N_28123,N_24024);
or U31774 (N_31774,N_28992,N_23422);
nor U31775 (N_31775,N_25695,N_22976);
or U31776 (N_31776,N_27309,N_28832);
or U31777 (N_31777,N_24210,N_27355);
xnor U31778 (N_31778,N_25969,N_23730);
and U31779 (N_31779,N_26949,N_26580);
or U31780 (N_31780,N_25597,N_28460);
nor U31781 (N_31781,N_20894,N_20617);
nand U31782 (N_31782,N_29408,N_28732);
xor U31783 (N_31783,N_24648,N_26867);
nand U31784 (N_31784,N_26540,N_23139);
and U31785 (N_31785,N_24840,N_29538);
nand U31786 (N_31786,N_29291,N_26958);
or U31787 (N_31787,N_25539,N_22312);
nand U31788 (N_31788,N_24699,N_25862);
nor U31789 (N_31789,N_25961,N_24332);
nand U31790 (N_31790,N_24562,N_21916);
and U31791 (N_31791,N_24026,N_24266);
nand U31792 (N_31792,N_27331,N_25590);
or U31793 (N_31793,N_24133,N_21571);
or U31794 (N_31794,N_23360,N_26680);
nand U31795 (N_31795,N_26480,N_25509);
or U31796 (N_31796,N_23810,N_21421);
and U31797 (N_31797,N_23305,N_29576);
nor U31798 (N_31798,N_28114,N_26293);
nor U31799 (N_31799,N_22498,N_25430);
or U31800 (N_31800,N_28621,N_22103);
nor U31801 (N_31801,N_23450,N_28565);
or U31802 (N_31802,N_27772,N_29341);
xor U31803 (N_31803,N_25809,N_24904);
nor U31804 (N_31804,N_26990,N_23249);
xnor U31805 (N_31805,N_29213,N_21249);
nor U31806 (N_31806,N_25867,N_20655);
nor U31807 (N_31807,N_29025,N_28312);
xor U31808 (N_31808,N_26489,N_24486);
and U31809 (N_31809,N_24414,N_25460);
nor U31810 (N_31810,N_27080,N_20560);
or U31811 (N_31811,N_20145,N_29434);
or U31812 (N_31812,N_27411,N_20458);
nor U31813 (N_31813,N_22912,N_26814);
and U31814 (N_31814,N_22301,N_20882);
nand U31815 (N_31815,N_20953,N_26145);
nand U31816 (N_31816,N_26567,N_22601);
nand U31817 (N_31817,N_27946,N_29805);
or U31818 (N_31818,N_23996,N_23275);
and U31819 (N_31819,N_26089,N_29133);
nor U31820 (N_31820,N_20503,N_23454);
nand U31821 (N_31821,N_27935,N_25077);
and U31822 (N_31822,N_21218,N_27147);
and U31823 (N_31823,N_23247,N_25384);
and U31824 (N_31824,N_21616,N_26973);
nor U31825 (N_31825,N_25741,N_28249);
and U31826 (N_31826,N_29376,N_24219);
and U31827 (N_31827,N_21910,N_20820);
or U31828 (N_31828,N_25873,N_28676);
xnor U31829 (N_31829,N_28594,N_24571);
xor U31830 (N_31830,N_26287,N_20610);
and U31831 (N_31831,N_29977,N_27165);
nand U31832 (N_31832,N_24446,N_23769);
and U31833 (N_31833,N_22327,N_23926);
nor U31834 (N_31834,N_20032,N_23909);
nor U31835 (N_31835,N_26313,N_29415);
nor U31836 (N_31836,N_21715,N_21780);
nor U31837 (N_31837,N_27712,N_26717);
nand U31838 (N_31838,N_28377,N_21911);
nor U31839 (N_31839,N_23980,N_26906);
or U31840 (N_31840,N_20967,N_27553);
nor U31841 (N_31841,N_28236,N_22559);
nand U31842 (N_31842,N_27229,N_22752);
or U31843 (N_31843,N_25089,N_21611);
and U31844 (N_31844,N_22618,N_23824);
or U31845 (N_31845,N_28084,N_28644);
nand U31846 (N_31846,N_26931,N_29153);
xor U31847 (N_31847,N_20501,N_23426);
xor U31848 (N_31848,N_25607,N_26510);
or U31849 (N_31849,N_26668,N_21312);
xor U31850 (N_31850,N_22605,N_27743);
nand U31851 (N_31851,N_23059,N_29917);
or U31852 (N_31852,N_25582,N_20498);
nor U31853 (N_31853,N_24485,N_25912);
or U31854 (N_31854,N_21509,N_20094);
and U31855 (N_31855,N_25279,N_27120);
or U31856 (N_31856,N_25555,N_22065);
nand U31857 (N_31857,N_22446,N_26367);
nand U31858 (N_31858,N_25281,N_21147);
nor U31859 (N_31859,N_24815,N_22099);
and U31860 (N_31860,N_23617,N_21006);
and U31861 (N_31861,N_22726,N_25823);
xor U31862 (N_31862,N_28433,N_25850);
nor U31863 (N_31863,N_26890,N_25879);
and U31864 (N_31864,N_27961,N_21512);
nor U31865 (N_31865,N_21143,N_22662);
or U31866 (N_31866,N_23068,N_28480);
xnor U31867 (N_31867,N_29658,N_21991);
and U31868 (N_31868,N_25376,N_26157);
or U31869 (N_31869,N_23413,N_25531);
nand U31870 (N_31870,N_28489,N_20768);
nor U31871 (N_31871,N_26985,N_24320);
nand U31872 (N_31872,N_22998,N_22194);
nor U31873 (N_31873,N_25213,N_20218);
or U31874 (N_31874,N_29368,N_23431);
nand U31875 (N_31875,N_25939,N_26568);
and U31876 (N_31876,N_20159,N_23965);
nor U31877 (N_31877,N_28578,N_27315);
and U31878 (N_31878,N_22266,N_26097);
nand U31879 (N_31879,N_23008,N_20547);
and U31880 (N_31880,N_24247,N_25730);
nor U31881 (N_31881,N_24876,N_26904);
xor U31882 (N_31882,N_28883,N_21984);
and U31883 (N_31883,N_28830,N_29835);
nor U31884 (N_31884,N_26340,N_28524);
nor U31885 (N_31885,N_28224,N_24702);
nor U31886 (N_31886,N_21484,N_22768);
nand U31887 (N_31887,N_27322,N_27024);
nand U31888 (N_31888,N_26485,N_27827);
and U31889 (N_31889,N_22170,N_24950);
xor U31890 (N_31890,N_23862,N_20686);
nand U31891 (N_31891,N_29926,N_29635);
and U31892 (N_31892,N_22824,N_23227);
and U31893 (N_31893,N_21528,N_27536);
nand U31894 (N_31894,N_25259,N_26096);
and U31895 (N_31895,N_22355,N_22114);
or U31896 (N_31896,N_21632,N_28966);
or U31897 (N_31897,N_26372,N_23943);
or U31898 (N_31898,N_21521,N_29681);
nor U31899 (N_31899,N_20808,N_28075);
and U31900 (N_31900,N_28976,N_26143);
nor U31901 (N_31901,N_28231,N_20291);
xor U31902 (N_31902,N_27136,N_25197);
or U31903 (N_31903,N_20572,N_25283);
nor U31904 (N_31904,N_28032,N_28279);
and U31905 (N_31905,N_22006,N_20129);
xor U31906 (N_31906,N_22641,N_29588);
or U31907 (N_31907,N_24684,N_25960);
xnor U31908 (N_31908,N_27922,N_23156);
xor U31909 (N_31909,N_23907,N_22321);
nor U31910 (N_31910,N_23657,N_22509);
or U31911 (N_31911,N_21951,N_25008);
nor U31912 (N_31912,N_25720,N_26937);
nor U31913 (N_31913,N_28910,N_26401);
nand U31914 (N_31914,N_21277,N_27059);
or U31915 (N_31915,N_29052,N_25038);
xnor U31916 (N_31916,N_27715,N_21637);
or U31917 (N_31917,N_20952,N_22105);
nor U31918 (N_31918,N_29210,N_26648);
nor U31919 (N_31919,N_20797,N_21990);
or U31920 (N_31920,N_20052,N_22660);
nand U31921 (N_31921,N_22869,N_27227);
and U31922 (N_31922,N_26033,N_26972);
or U31923 (N_31923,N_22826,N_26763);
and U31924 (N_31924,N_26836,N_22231);
and U31925 (N_31925,N_22120,N_27928);
nand U31926 (N_31926,N_24232,N_26635);
and U31927 (N_31927,N_27931,N_22003);
or U31928 (N_31928,N_22246,N_20150);
xnor U31929 (N_31929,N_24909,N_27130);
nor U31930 (N_31930,N_22732,N_22582);
or U31931 (N_31931,N_21446,N_24557);
xnor U31932 (N_31932,N_24360,N_29430);
and U31933 (N_31933,N_23505,N_24731);
nand U31934 (N_31934,N_29014,N_26864);
nor U31935 (N_31935,N_29024,N_22411);
or U31936 (N_31936,N_24129,N_27840);
nand U31937 (N_31937,N_24926,N_20420);
nor U31938 (N_31938,N_25722,N_26541);
and U31939 (N_31939,N_28564,N_22589);
nor U31940 (N_31940,N_20355,N_25522);
and U31941 (N_31941,N_28928,N_22556);
xor U31942 (N_31942,N_22425,N_22057);
or U31943 (N_31943,N_27515,N_25496);
xor U31944 (N_31944,N_20955,N_23523);
nor U31945 (N_31945,N_27861,N_27803);
nor U31946 (N_31946,N_29714,N_27947);
xnor U31947 (N_31947,N_29349,N_29666);
nor U31948 (N_31948,N_28901,N_28775);
or U31949 (N_31949,N_25329,N_25288);
and U31950 (N_31950,N_20546,N_25457);
xnor U31951 (N_31951,N_25965,N_20945);
nor U31952 (N_31952,N_25694,N_26884);
nor U31953 (N_31953,N_21939,N_21078);
or U31954 (N_31954,N_28338,N_29546);
nand U31955 (N_31955,N_28367,N_25914);
and U31956 (N_31956,N_25003,N_24663);
nand U31957 (N_31957,N_27982,N_22782);
nor U31958 (N_31958,N_22778,N_23988);
and U31959 (N_31959,N_20550,N_25988);
or U31960 (N_31960,N_27470,N_22040);
and U31961 (N_31961,N_20486,N_27964);
and U31962 (N_31962,N_27385,N_20850);
or U31963 (N_31963,N_25193,N_29302);
nand U31964 (N_31964,N_29338,N_23749);
or U31965 (N_31965,N_28856,N_24333);
nor U31966 (N_31966,N_23547,N_23739);
or U31967 (N_31967,N_23729,N_22148);
xnor U31968 (N_31968,N_28908,N_27330);
nor U31969 (N_31969,N_25704,N_23529);
xor U31970 (N_31970,N_27572,N_28837);
nor U31971 (N_31971,N_25768,N_27341);
nand U31972 (N_31972,N_29942,N_25478);
and U31973 (N_31973,N_21671,N_25767);
nor U31974 (N_31974,N_29719,N_22122);
nor U31975 (N_31975,N_23557,N_28807);
and U31976 (N_31976,N_21520,N_23052);
and U31977 (N_31977,N_27864,N_22689);
nand U31978 (N_31978,N_23455,N_29361);
and U31979 (N_31979,N_22240,N_28741);
and U31980 (N_31980,N_23544,N_21436);
nand U31981 (N_31981,N_24441,N_25055);
xnor U31982 (N_31982,N_28645,N_29552);
and U31983 (N_31983,N_27934,N_23695);
and U31984 (N_31984,N_27372,N_21851);
and U31985 (N_31985,N_21286,N_23131);
or U31986 (N_31986,N_25163,N_28485);
xor U31987 (N_31987,N_23530,N_28561);
nor U31988 (N_31988,N_24458,N_21732);
nand U31989 (N_31989,N_25848,N_28968);
xnor U31990 (N_31990,N_21775,N_26343);
or U31991 (N_31991,N_28939,N_24875);
nor U31992 (N_31992,N_28850,N_25133);
or U31993 (N_31993,N_28468,N_21747);
or U31994 (N_31994,N_21869,N_29906);
nand U31995 (N_31995,N_27220,N_24706);
nand U31996 (N_31996,N_22551,N_23623);
nor U31997 (N_31997,N_27697,N_25631);
or U31998 (N_31998,N_20106,N_24202);
nand U31999 (N_31999,N_27573,N_25064);
and U32000 (N_32000,N_21226,N_23513);
nor U32001 (N_32001,N_26265,N_21199);
or U32002 (N_32002,N_28373,N_27742);
xnor U32003 (N_32003,N_21964,N_22303);
or U32004 (N_32004,N_27494,N_23786);
nor U32005 (N_32005,N_21965,N_24234);
nand U32006 (N_32006,N_25818,N_27917);
nand U32007 (N_32007,N_29075,N_29391);
and U32008 (N_32008,N_26435,N_24205);
and U32009 (N_32009,N_20067,N_23566);
nand U32010 (N_32010,N_29708,N_21116);
nor U32011 (N_32011,N_24062,N_29743);
or U32012 (N_32012,N_21988,N_22055);
nand U32013 (N_32013,N_22308,N_29073);
nand U32014 (N_32014,N_20092,N_26778);
nand U32015 (N_32015,N_23883,N_25758);
and U32016 (N_32016,N_28074,N_27694);
nand U32017 (N_32017,N_21266,N_21485);
or U32018 (N_32018,N_26150,N_20434);
and U32019 (N_32019,N_22376,N_23589);
or U32020 (N_32020,N_29991,N_23272);
xor U32021 (N_32021,N_24242,N_24422);
nand U32022 (N_32022,N_24426,N_26970);
nand U32023 (N_32023,N_29730,N_21902);
nand U32024 (N_32024,N_25874,N_22704);
or U32025 (N_32025,N_24527,N_25918);
or U32026 (N_32026,N_23151,N_24672);
or U32027 (N_32027,N_21734,N_22603);
and U32028 (N_32028,N_24019,N_21864);
and U32029 (N_32029,N_22228,N_20738);
nand U32030 (N_32030,N_24792,N_24315);
nand U32031 (N_32031,N_22206,N_22843);
and U32032 (N_32032,N_23129,N_27113);
and U32033 (N_32033,N_24104,N_27600);
or U32034 (N_32034,N_21269,N_27351);
nand U32035 (N_32035,N_28385,N_25081);
nand U32036 (N_32036,N_24184,N_27833);
and U32037 (N_32037,N_29825,N_26255);
or U32038 (N_32038,N_26886,N_24824);
xor U32039 (N_32039,N_29143,N_25845);
or U32040 (N_32040,N_23449,N_25870);
or U32041 (N_32041,N_27848,N_21438);
nand U32042 (N_32042,N_23103,N_27995);
nor U32043 (N_32043,N_27555,N_23679);
nand U32044 (N_32044,N_24374,N_21517);
nor U32045 (N_32045,N_27898,N_29727);
nand U32046 (N_32046,N_29047,N_29040);
nor U32047 (N_32047,N_26547,N_20661);
nand U32048 (N_32048,N_20387,N_23649);
nor U32049 (N_32049,N_27965,N_21025);
nor U32050 (N_32050,N_26180,N_21948);
xnor U32051 (N_32051,N_22882,N_22503);
nand U32052 (N_32052,N_23686,N_29364);
nand U32053 (N_32053,N_23185,N_29158);
nand U32054 (N_32054,N_28118,N_29155);
nor U32055 (N_32055,N_25275,N_27927);
or U32056 (N_32056,N_21826,N_21187);
xnor U32057 (N_32057,N_23778,N_23490);
nor U32058 (N_32058,N_20780,N_27363);
nor U32059 (N_32059,N_26408,N_23077);
nor U32060 (N_32060,N_26267,N_25463);
or U32061 (N_32061,N_26102,N_20144);
nor U32062 (N_32062,N_20335,N_24038);
xor U32063 (N_32063,N_23976,N_23779);
xnor U32064 (N_32064,N_29152,N_25108);
nor U32065 (N_32065,N_20852,N_29747);
nand U32066 (N_32066,N_21779,N_25528);
nand U32067 (N_32067,N_20752,N_22953);
and U32068 (N_32068,N_27267,N_25370);
nor U32069 (N_32069,N_26374,N_29843);
nand U32070 (N_32070,N_23166,N_24365);
nor U32071 (N_32071,N_24611,N_23236);
nor U32072 (N_32072,N_26913,N_26451);
nor U32073 (N_32073,N_28459,N_25239);
and U32074 (N_32074,N_25086,N_26549);
xor U32075 (N_32075,N_28027,N_27166);
nor U32076 (N_32076,N_23259,N_20153);
or U32077 (N_32077,N_28116,N_21865);
nand U32078 (N_32078,N_26156,N_26312);
nand U32079 (N_32079,N_25700,N_29590);
nand U32080 (N_32080,N_26486,N_20626);
xnor U32081 (N_32081,N_29094,N_28291);
nand U32082 (N_32082,N_22282,N_24715);
nor U32083 (N_32083,N_28397,N_20245);
nand U32084 (N_32084,N_22015,N_26420);
nand U32085 (N_32085,N_25051,N_23435);
nor U32086 (N_32086,N_20974,N_27451);
nor U32087 (N_32087,N_27265,N_23673);
and U32088 (N_32088,N_24054,N_27107);
or U32089 (N_32089,N_23394,N_28760);
or U32090 (N_32090,N_23861,N_29852);
nand U32091 (N_32091,N_25171,N_20604);
nand U32092 (N_32092,N_20832,N_20307);
nand U32093 (N_32093,N_26251,N_23707);
nor U32094 (N_32094,N_28551,N_23855);
and U32095 (N_32095,N_21043,N_25501);
xnor U32096 (N_32096,N_29109,N_21119);
or U32097 (N_32097,N_28819,N_23644);
xor U32098 (N_32098,N_25835,N_22875);
nand U32099 (N_32099,N_26433,N_20217);
nand U32100 (N_32100,N_23863,N_29048);
nand U32101 (N_32101,N_23427,N_28060);
xor U32102 (N_32102,N_22166,N_29358);
nor U32103 (N_32103,N_20724,N_21414);
or U32104 (N_32104,N_27405,N_29017);
or U32105 (N_32105,N_20998,N_20678);
xor U32106 (N_32106,N_23992,N_22970);
xor U32107 (N_32107,N_29071,N_29920);
or U32108 (N_32108,N_20422,N_20761);
or U32109 (N_32109,N_25900,N_28658);
or U32110 (N_32110,N_25527,N_28071);
nor U32111 (N_32111,N_29382,N_28967);
xnor U32112 (N_32112,N_28525,N_22566);
nand U32113 (N_32113,N_23825,N_22809);
xnor U32114 (N_32114,N_21595,N_22899);
xor U32115 (N_32115,N_26737,N_26360);
nand U32116 (N_32116,N_25931,N_21389);
nor U32117 (N_32117,N_21707,N_20745);
xnor U32118 (N_32118,N_23215,N_22310);
nand U32119 (N_32119,N_24758,N_27754);
nor U32120 (N_32120,N_24776,N_21424);
nor U32121 (N_32121,N_29107,N_24427);
or U32122 (N_32122,N_20239,N_28804);
or U32123 (N_32123,N_26871,N_26895);
and U32124 (N_32124,N_29078,N_28940);
or U32125 (N_32125,N_22132,N_28876);
or U32126 (N_32126,N_26185,N_26050);
nand U32127 (N_32127,N_29734,N_20240);
and U32128 (N_32128,N_22476,N_23675);
nand U32129 (N_32129,N_21439,N_29229);
and U32130 (N_32130,N_24536,N_24920);
or U32131 (N_32131,N_24613,N_27851);
nor U32132 (N_32132,N_27344,N_26698);
or U32133 (N_32133,N_26858,N_22449);
or U32134 (N_32134,N_25053,N_26037);
nand U32135 (N_32135,N_28906,N_20454);
nor U32136 (N_32136,N_25769,N_24996);
nor U32137 (N_32137,N_21749,N_20082);
or U32138 (N_32138,N_29432,N_24597);
nand U32139 (N_32139,N_25091,N_22096);
or U32140 (N_32140,N_22841,N_28496);
or U32141 (N_32141,N_21994,N_28136);
or U32142 (N_32142,N_22185,N_23317);
and U32143 (N_32143,N_28872,N_22632);
or U32144 (N_32144,N_28780,N_26269);
or U32145 (N_32145,N_21549,N_23337);
and U32146 (N_32146,N_25307,N_24345);
or U32147 (N_32147,N_29668,N_21809);
nand U32148 (N_32148,N_27430,N_26667);
nor U32149 (N_32149,N_21839,N_27766);
or U32150 (N_32150,N_21729,N_21683);
nor U32151 (N_32151,N_27015,N_28709);
and U32152 (N_32152,N_20530,N_23130);
nor U32153 (N_32153,N_28824,N_23641);
and U32154 (N_32154,N_26148,N_28586);
or U32155 (N_32155,N_29279,N_20409);
and U32156 (N_32156,N_21529,N_23214);
or U32157 (N_32157,N_28635,N_27503);
and U32158 (N_32158,N_21061,N_21598);
and U32159 (N_32159,N_28220,N_20627);
and U32160 (N_32160,N_27936,N_28318);
xor U32161 (N_32161,N_27707,N_29716);
nand U32162 (N_32162,N_20126,N_23696);
and U32163 (N_32163,N_27547,N_23395);
nor U32164 (N_32164,N_22195,N_29369);
and U32165 (N_32165,N_29289,N_28861);
and U32166 (N_32166,N_27247,N_28814);
and U32167 (N_32167,N_29919,N_26511);
nand U32168 (N_32168,N_27605,N_27684);
nor U32169 (N_32169,N_26331,N_29295);
or U32170 (N_32170,N_20118,N_28102);
and U32171 (N_32171,N_27825,N_26115);
nor U32172 (N_32172,N_25453,N_22837);
and U32173 (N_32173,N_28765,N_23512);
nor U32174 (N_32174,N_20804,N_26175);
nor U32175 (N_32175,N_22155,N_28867);
and U32176 (N_32176,N_22238,N_29181);
nor U32177 (N_32177,N_25435,N_22636);
nor U32178 (N_32178,N_21815,N_27398);
and U32179 (N_32179,N_29077,N_29988);
nor U32180 (N_32180,N_28264,N_22909);
nand U32181 (N_32181,N_28158,N_27630);
or U32182 (N_32182,N_29824,N_27990);
and U32183 (N_32183,N_25922,N_28041);
and U32184 (N_32184,N_28826,N_25489);
nand U32185 (N_32185,N_27475,N_28521);
and U32186 (N_32186,N_25683,N_27389);
or U32187 (N_32187,N_29184,N_26233);
xor U32188 (N_32188,N_22402,N_22889);
and U32189 (N_32189,N_20723,N_20864);
xnor U32190 (N_32190,N_27348,N_25485);
nand U32191 (N_32191,N_24091,N_21384);
and U32192 (N_32192,N_21322,N_26047);
and U32193 (N_32193,N_20989,N_29104);
nand U32194 (N_32194,N_22032,N_22590);
nor U32195 (N_32195,N_24783,N_25863);
nor U32196 (N_32196,N_23193,N_23421);
nor U32197 (N_32197,N_26693,N_20897);
nor U32198 (N_32198,N_24544,N_23072);
and U32199 (N_32199,N_28854,N_20624);
nor U32200 (N_32200,N_27274,N_25909);
nor U32201 (N_32201,N_20234,N_24873);
and U32202 (N_32202,N_20311,N_26351);
and U32203 (N_32203,N_20500,N_23999);
or U32204 (N_32204,N_21889,N_22558);
nand U32205 (N_32205,N_26561,N_26111);
or U32206 (N_32206,N_23419,N_23791);
and U32207 (N_32207,N_20675,N_26910);
or U32208 (N_32208,N_23291,N_27106);
and U32209 (N_32209,N_29119,N_26074);
and U32210 (N_32210,N_29645,N_22880);
nand U32211 (N_32211,N_23069,N_25851);
or U32212 (N_32212,N_29889,N_29219);
nor U32213 (N_32213,N_20884,N_20991);
nand U32214 (N_32214,N_24635,N_27590);
or U32215 (N_32215,N_25125,N_24070);
and U32216 (N_32216,N_25291,N_27668);
and U32217 (N_32217,N_20814,N_29203);
and U32218 (N_32218,N_29792,N_25065);
or U32219 (N_32219,N_24178,N_21031);
nand U32220 (N_32220,N_26727,N_22335);
nor U32221 (N_32221,N_21975,N_28475);
nand U32222 (N_32222,N_25249,N_24200);
xnor U32223 (N_32223,N_20648,N_20130);
or U32224 (N_32224,N_29954,N_22473);
nand U32225 (N_32225,N_24078,N_26571);
or U32226 (N_32226,N_22154,N_25230);
nor U32227 (N_32227,N_25270,N_21472);
and U32228 (N_32228,N_27116,N_26308);
and U32229 (N_32229,N_26545,N_25371);
nor U32230 (N_32230,N_29460,N_23846);
or U32231 (N_32231,N_28813,N_25658);
and U32232 (N_32232,N_26915,N_20577);
nor U32233 (N_32233,N_22952,N_25925);
nand U32234 (N_32234,N_22045,N_27200);
nor U32235 (N_32235,N_23752,N_20051);
nand U32236 (N_32236,N_24652,N_21017);
or U32237 (N_32237,N_29117,N_26494);
nand U32238 (N_32238,N_26775,N_24812);
nor U32239 (N_32239,N_21085,N_21772);
or U32240 (N_32240,N_25107,N_29837);
nand U32241 (N_32241,N_25398,N_22908);
and U32242 (N_32242,N_28553,N_23650);
and U32243 (N_32243,N_24057,N_20776);
and U32244 (N_32244,N_29996,N_22947);
nor U32245 (N_32245,N_20192,N_21825);
nand U32246 (N_32246,N_23218,N_20314);
and U32247 (N_32247,N_29417,N_28727);
and U32248 (N_32248,N_25540,N_24832);
and U32249 (N_32249,N_24480,N_26425);
or U32250 (N_32250,N_27844,N_23201);
or U32251 (N_32251,N_26484,N_28512);
xnor U32252 (N_32252,N_21430,N_24503);
and U32253 (N_32253,N_28950,N_26961);
nand U32254 (N_32254,N_23511,N_22991);
and U32255 (N_32255,N_26238,N_22445);
and U32256 (N_32256,N_25379,N_27100);
and U32257 (N_32257,N_27460,N_21837);
nand U32258 (N_32258,N_24089,N_22776);
or U32259 (N_32259,N_29993,N_29425);
or U32260 (N_32260,N_22237,N_24128);
or U32261 (N_32261,N_22395,N_28268);
or U32262 (N_32262,N_20825,N_24077);
nor U32263 (N_32263,N_25302,N_29973);
nand U32264 (N_32264,N_27602,N_25843);
or U32265 (N_32265,N_23581,N_29803);
xnor U32266 (N_32266,N_26264,N_29820);
nand U32267 (N_32267,N_26889,N_25913);
xor U32268 (N_32268,N_29892,N_20504);
nand U32269 (N_32269,N_25294,N_22244);
or U32270 (N_32270,N_27295,N_29571);
or U32271 (N_32271,N_21004,N_24217);
xor U32272 (N_32272,N_23993,N_24076);
nor U32273 (N_32273,N_28366,N_29767);
and U32274 (N_32274,N_25865,N_24305);
nor U32275 (N_32275,N_24289,N_21442);
nor U32276 (N_32276,N_28768,N_29142);
nor U32277 (N_32277,N_24469,N_27101);
or U32278 (N_32278,N_25836,N_22455);
xor U32279 (N_32279,N_26055,N_28203);
nor U32280 (N_32280,N_28584,N_23248);
and U32281 (N_32281,N_20391,N_23229);
and U32282 (N_32282,N_20223,N_23108);
or U32283 (N_32283,N_20103,N_27871);
nor U32284 (N_32284,N_25405,N_23083);
and U32285 (N_32285,N_29533,N_26035);
nand U32286 (N_32286,N_24695,N_22828);
xnor U32287 (N_32287,N_22854,N_27191);
nor U32288 (N_32288,N_27097,N_24735);
and U32289 (N_32289,N_25627,N_26221);
nor U32290 (N_32290,N_20507,N_23703);
or U32291 (N_32291,N_21243,N_23387);
nand U32292 (N_32292,N_25726,N_22577);
nand U32293 (N_32293,N_23804,N_24530);
and U32294 (N_32294,N_28591,N_25905);
nand U32295 (N_32295,N_24464,N_23306);
or U32296 (N_32296,N_26801,N_22864);
and U32297 (N_32297,N_27458,N_27396);
nand U32298 (N_32298,N_24391,N_25078);
xor U32299 (N_32299,N_26223,N_25426);
xnor U32300 (N_32300,N_28053,N_20983);
nor U32301 (N_32301,N_28257,N_27242);
nor U32302 (N_32302,N_22184,N_20011);
xnor U32303 (N_32303,N_25201,N_27858);
nand U32304 (N_32304,N_27278,N_25492);
nand U32305 (N_32305,N_27393,N_27574);
nor U32306 (N_32306,N_28753,N_20274);
nand U32307 (N_32307,N_21158,N_23092);
xor U32308 (N_32308,N_22072,N_23630);
or U32309 (N_32309,N_22341,N_26201);
or U32310 (N_32310,N_27974,N_23280);
and U32311 (N_32311,N_23443,N_24903);
nor U32312 (N_32312,N_28573,N_24806);
nand U32313 (N_32313,N_21764,N_29275);
nand U32314 (N_32314,N_25705,N_26887);
nand U32315 (N_32315,N_27359,N_29788);
nor U32316 (N_32316,N_25620,N_25592);
or U32317 (N_32317,N_27262,N_21792);
and U32318 (N_32318,N_24549,N_26137);
or U32319 (N_32319,N_20061,N_25737);
xor U32320 (N_32320,N_21285,N_27122);
nor U32321 (N_32321,N_22696,N_29901);
nand U32322 (N_32322,N_23564,N_28798);
nand U32323 (N_32323,N_22657,N_26326);
nand U32324 (N_32324,N_28880,N_20428);
and U32325 (N_32325,N_22288,N_29475);
and U32326 (N_32326,N_24576,N_23176);
or U32327 (N_32327,N_29965,N_26570);
nor U32328 (N_32328,N_26432,N_27926);
xnor U32329 (N_32329,N_27143,N_24438);
or U32330 (N_32330,N_20429,N_29074);
nor U32331 (N_32331,N_24463,N_23924);
nor U32332 (N_32332,N_24953,N_28762);
nor U32333 (N_32333,N_24160,N_25886);
nand U32334 (N_32334,N_28877,N_21845);
xor U32335 (N_32335,N_24112,N_26410);
and U32336 (N_32336,N_21018,N_24073);
and U32337 (N_32337,N_22022,N_29818);
and U32338 (N_32338,N_24786,N_21314);
and U32339 (N_32339,N_20956,N_21170);
xor U32340 (N_32340,N_26573,N_25902);
and U32341 (N_32341,N_27403,N_27641);
or U32342 (N_32342,N_22417,N_24372);
nor U32343 (N_32343,N_20753,N_25312);
and U32344 (N_32344,N_24615,N_26499);
nand U32345 (N_32345,N_26353,N_26506);
and U32346 (N_32346,N_25917,N_22033);
or U32347 (N_32347,N_26862,N_26902);
nand U32348 (N_32348,N_25029,N_29879);
and U32349 (N_32349,N_25713,N_23338);
xnor U32350 (N_32350,N_29986,N_20287);
or U32351 (N_32351,N_21241,N_26791);
xnor U32352 (N_32352,N_20098,N_26750);
nand U32353 (N_32353,N_24554,N_20966);
nor U32354 (N_32354,N_29260,N_26610);
nand U32355 (N_32355,N_26768,N_26664);
xnor U32356 (N_32356,N_28590,N_25661);
or U32357 (N_32357,N_22534,N_26471);
nor U32358 (N_32358,N_23242,N_21784);
xnor U32359 (N_32359,N_20911,N_22492);
and U32360 (N_32360,N_29324,N_24270);
xnor U32361 (N_32361,N_24932,N_25049);
and U32362 (N_32362,N_26856,N_29284);
nor U32363 (N_32363,N_21141,N_24727);
xor U32364 (N_32364,N_25535,N_25829);
or U32365 (N_32365,N_22832,N_27748);
nor U32366 (N_32366,N_20915,N_26248);
or U32367 (N_32367,N_24067,N_23853);
or U32368 (N_32368,N_26272,N_25649);
xnor U32369 (N_32369,N_22436,N_22842);
or U32370 (N_32370,N_23342,N_26707);
nand U32371 (N_32371,N_20122,N_25455);
and U32372 (N_32372,N_20823,N_29532);
nor U32373 (N_32373,N_23569,N_23925);
nor U32374 (N_32374,N_23463,N_29332);
and U32375 (N_32375,N_22309,N_27548);
nor U32376 (N_32376,N_20818,N_22553);
nand U32377 (N_32377,N_27666,N_28382);
nor U32378 (N_32378,N_28718,N_20160);
nand U32379 (N_32379,N_27656,N_26963);
and U32380 (N_32380,N_22167,N_28661);
or U32381 (N_32381,N_22260,N_21651);
nor U32382 (N_32382,N_21465,N_29301);
nor U32383 (N_32383,N_24990,N_28466);
nor U32384 (N_32384,N_28949,N_24795);
and U32385 (N_32385,N_26552,N_25229);
nand U32386 (N_32386,N_21476,N_22986);
nor U32387 (N_32387,N_20161,N_20636);
nand U32388 (N_32388,N_22761,N_22996);
xor U32389 (N_32389,N_27703,N_28777);
nand U32390 (N_32390,N_27826,N_22973);
nand U32391 (N_32391,N_23878,N_26493);
and U32392 (N_32392,N_24907,N_25475);
and U32393 (N_32393,N_29161,N_26318);
nor U32394 (N_32394,N_27577,N_22125);
or U32395 (N_32395,N_29209,N_25399);
nand U32396 (N_32396,N_24261,N_27669);
and U32397 (N_32397,N_27072,N_28246);
and U32398 (N_32398,N_28497,N_22396);
nor U32399 (N_32399,N_26512,N_28403);
xor U32400 (N_32400,N_27719,N_25979);
nand U32401 (N_32401,N_25932,N_29466);
and U32402 (N_32402,N_28454,N_28319);
nor U32403 (N_32403,N_21106,N_27332);
or U32404 (N_32404,N_20178,N_26070);
nand U32405 (N_32405,N_29387,N_26170);
nand U32406 (N_32406,N_21072,N_26324);
or U32407 (N_32407,N_22051,N_25210);
and U32408 (N_32408,N_28013,N_27648);
and U32409 (N_32409,N_20999,N_22769);
or U32410 (N_32410,N_23310,N_22253);
and U32411 (N_32411,N_20555,N_24857);
xor U32412 (N_32412,N_23335,N_22387);
or U32413 (N_32413,N_20873,N_22722);
nand U32414 (N_32414,N_20267,N_24168);
or U32415 (N_32415,N_22621,N_21254);
nand U32416 (N_32416,N_28614,N_24762);
nor U32417 (N_32417,N_26581,N_20216);
nor U32418 (N_32418,N_21217,N_22481);
xor U32419 (N_32419,N_21108,N_26108);
or U32420 (N_32420,N_20682,N_26631);
nand U32421 (N_32421,N_22733,N_22009);
nor U32422 (N_32422,N_20062,N_25556);
nand U32423 (N_32423,N_23570,N_25437);
or U32424 (N_32424,N_26891,N_21502);
nand U32425 (N_32425,N_29087,N_28895);
nor U32426 (N_32426,N_27592,N_25383);
and U32427 (N_32427,N_29321,N_29395);
nand U32428 (N_32428,N_21410,N_21007);
or U32429 (N_32429,N_22791,N_21494);
or U32430 (N_32430,N_27436,N_22516);
xnor U32431 (N_32431,N_24767,N_28994);
xnor U32432 (N_32432,N_25115,N_25416);
or U32433 (N_32433,N_21306,N_24551);
or U32434 (N_32434,N_20742,N_23315);
nand U32435 (N_32435,N_27508,N_21066);
and U32436 (N_32436,N_20536,N_24803);
nand U32437 (N_32437,N_26280,N_20083);
nor U32438 (N_32438,N_26914,N_20001);
and U32439 (N_32439,N_25565,N_23157);
nor U32440 (N_32440,N_22669,N_29241);
or U32441 (N_32441,N_20316,N_20740);
nor U32442 (N_32442,N_20342,N_22401);
and U32443 (N_32443,N_28119,N_23045);
nand U32444 (N_32444,N_24753,N_28784);
nor U32445 (N_32445,N_28122,N_29043);
and U32446 (N_32446,N_28453,N_26418);
and U32447 (N_32447,N_22218,N_24657);
nand U32448 (N_32448,N_22613,N_27066);
nor U32449 (N_32449,N_25487,N_20463);
and U32450 (N_32450,N_25380,N_28088);
or U32451 (N_32451,N_20848,N_28514);
nand U32452 (N_32452,N_29233,N_27383);
nor U32453 (N_32453,N_21538,N_27855);
xnor U32454 (N_32454,N_29648,N_28739);
and U32455 (N_32455,N_26585,N_26615);
nand U32456 (N_32456,N_23773,N_24545);
nor U32457 (N_32457,N_21663,N_26855);
nand U32458 (N_32458,N_21493,N_23562);
nand U32459 (N_32459,N_25497,N_29968);
xor U32460 (N_32460,N_26347,N_24445);
nand U32461 (N_32461,N_24349,N_22656);
and U32462 (N_32462,N_21259,N_21203);
or U32463 (N_32463,N_28502,N_27164);
and U32464 (N_32464,N_23516,N_26213);
or U32465 (N_32465,N_26809,N_23525);
and U32466 (N_32466,N_28738,N_29070);
nor U32467 (N_32467,N_27651,N_28548);
or U32468 (N_32468,N_26422,N_26752);
nor U32469 (N_32469,N_22400,N_27615);
or U32470 (N_32470,N_27239,N_21021);
nand U32471 (N_32471,N_23182,N_20177);
or U32472 (N_32472,N_28051,N_26728);
or U32473 (N_32473,N_22879,N_25637);
or U32474 (N_32474,N_28618,N_21574);
xor U32475 (N_32475,N_24351,N_29745);
nor U32476 (N_32476,N_22397,N_29290);
or U32477 (N_32477,N_28055,N_26565);
nor U32478 (N_32478,N_20670,N_24359);
nand U32479 (N_32479,N_20666,N_29426);
or U32480 (N_32480,N_21204,N_25593);
or U32481 (N_32481,N_27225,N_24410);
and U32482 (N_32482,N_26428,N_27654);
xnor U32483 (N_32483,N_26716,N_29927);
or U32484 (N_32484,N_23233,N_27991);
nand U32485 (N_32485,N_26107,N_24420);
or U32486 (N_32486,N_20100,N_24094);
nand U32487 (N_32487,N_23807,N_27031);
xnor U32488 (N_32488,N_20297,N_28713);
or U32489 (N_32489,N_25883,N_27294);
nor U32490 (N_32490,N_20261,N_23997);
or U32491 (N_32491,N_24629,N_20535);
nor U32492 (N_32492,N_27125,N_22836);
nand U32493 (N_32493,N_24317,N_27259);
xnor U32494 (N_32494,N_27039,N_22486);
xor U32495 (N_32495,N_21875,N_21614);
xnor U32496 (N_32496,N_21381,N_23492);
nand U32497 (N_32497,N_28563,N_29565);
or U32498 (N_32498,N_26964,N_21335);
or U32499 (N_32499,N_22787,N_26813);
and U32500 (N_32500,N_28413,N_21051);
or U32501 (N_32501,N_25154,N_25338);
nand U32502 (N_32502,N_26834,N_28510);
and U32503 (N_32503,N_28669,N_21124);
nor U32504 (N_32504,N_20702,N_27637);
nand U32505 (N_32505,N_28438,N_20720);
or U32506 (N_32506,N_23125,N_22567);
nand U32507 (N_32507,N_26306,N_28596);
and U32508 (N_32508,N_24161,N_21268);
and U32509 (N_32509,N_22757,N_26989);
nand U32510 (N_32510,N_24235,N_20076);
or U32511 (N_32511,N_22594,N_22916);
and U32512 (N_32512,N_28469,N_23119);
nor U32513 (N_32513,N_28666,N_23416);
nand U32514 (N_32514,N_22428,N_25830);
and U32515 (N_32515,N_22679,N_28577);
and U32516 (N_32516,N_27850,N_26507);
or U32517 (N_32517,N_20665,N_25643);
nand U32518 (N_32518,N_29170,N_25547);
and U32519 (N_32519,N_28313,N_23372);
nand U32520 (N_32520,N_20737,N_28350);
and U32521 (N_32521,N_22723,N_21136);
nor U32522 (N_32522,N_27698,N_22855);
and U32523 (N_32523,N_21813,N_28424);
nand U32524 (N_32524,N_21406,N_24277);
xor U32525 (N_32525,N_28562,N_22939);
or U32526 (N_32526,N_28875,N_22391);
nand U32527 (N_32527,N_24127,N_20294);
nand U32528 (N_32528,N_20606,N_26924);
nand U32529 (N_32529,N_21501,N_26369);
nor U32530 (N_32530,N_22755,N_27052);
nor U32531 (N_32531,N_26383,N_21370);
nor U32532 (N_32532,N_29611,N_26018);
nand U32533 (N_32533,N_26762,N_27868);
or U32534 (N_32534,N_21140,N_22744);
nand U32535 (N_32535,N_27504,N_28663);
or U32536 (N_32536,N_23715,N_22807);
xnor U32537 (N_32537,N_29717,N_28808);
nand U32538 (N_32538,N_20855,N_20163);
or U32539 (N_32539,N_21720,N_20452);
nor U32540 (N_32540,N_20730,N_23213);
nand U32541 (N_32541,N_25070,N_27865);
and U32542 (N_32542,N_24856,N_29887);
and U32543 (N_32543,N_24387,N_28476);
nor U32544 (N_32544,N_21462,N_21492);
or U32545 (N_32545,N_24131,N_25578);
nand U32546 (N_32546,N_29118,N_25665);
nor U32547 (N_32547,N_27867,N_25512);
nand U32548 (N_32548,N_27159,N_22039);
or U32549 (N_32549,N_22406,N_25525);
nor U32550 (N_32550,N_22168,N_29212);
and U32551 (N_32551,N_27873,N_25984);
nor U32552 (N_32552,N_26126,N_20557);
nor U32553 (N_32553,N_25263,N_27316);
nor U32554 (N_32554,N_25319,N_25066);
nor U32555 (N_32555,N_27746,N_24040);
and U32556 (N_32556,N_20345,N_29436);
and U32557 (N_32557,N_26623,N_22701);
nor U32558 (N_32558,N_28284,N_20997);
or U32559 (N_32559,N_24922,N_20404);
and U32560 (N_32560,N_27701,N_20332);
xor U32561 (N_32561,N_29856,N_28054);
xnor U32562 (N_32562,N_28201,N_23370);
nor U32563 (N_32563,N_26041,N_25372);
and U32564 (N_32564,N_22857,N_28721);
and U32565 (N_32565,N_20900,N_26393);
or U32566 (N_32566,N_29860,N_22053);
or U32567 (N_32567,N_24342,N_22838);
xnor U32568 (N_32568,N_27042,N_23864);
and U32569 (N_32569,N_21514,N_23603);
nand U32570 (N_32570,N_23759,N_27270);
nand U32571 (N_32571,N_26384,N_28935);
or U32572 (N_32572,N_20199,N_24498);
nor U32573 (N_32573,N_23704,N_27140);
and U32574 (N_32574,N_23336,N_28490);
and U32575 (N_32575,N_22511,N_25264);
nor U32576 (N_32576,N_29640,N_23444);
nand U32577 (N_32577,N_29404,N_22667);
nand U32578 (N_32578,N_26794,N_26146);
nand U32579 (N_32579,N_20188,N_23712);
xnor U32580 (N_32580,N_21035,N_24324);
nor U32581 (N_32581,N_23205,N_27500);
and U32582 (N_32582,N_25500,N_22007);
or U32583 (N_32583,N_26774,N_21887);
nand U32584 (N_32584,N_27551,N_24834);
nand U32585 (N_32585,N_25889,N_28034);
or U32586 (N_32586,N_29329,N_29698);
nor U32587 (N_32587,N_23261,N_21194);
and U32588 (N_32588,N_22892,N_21190);
or U32589 (N_32589,N_26492,N_20136);
xor U32590 (N_32590,N_20696,N_22133);
nor U32591 (N_32591,N_24166,N_23152);
xnor U32592 (N_32592,N_22647,N_29450);
xnor U32593 (N_32593,N_21949,N_23274);
and U32594 (N_32594,N_22383,N_21934);
or U32595 (N_32595,N_20709,N_21198);
nand U32596 (N_32596,N_21838,N_21946);
and U32597 (N_32597,N_24899,N_26620);
xnor U32598 (N_32598,N_27945,N_28244);
nand U32599 (N_32599,N_21365,N_20259);
nor U32600 (N_32600,N_24572,N_22342);
or U32601 (N_32601,N_20616,N_27976);
nor U32602 (N_32602,N_28011,N_21201);
nand U32603 (N_32603,N_25977,N_23204);
and U32604 (N_32604,N_27319,N_29418);
and U32605 (N_32605,N_26575,N_28533);
nand U32606 (N_32606,N_29274,N_29646);
and U32607 (N_32607,N_25233,N_23553);
nand U32608 (N_32608,N_29494,N_20236);
or U32609 (N_32609,N_20638,N_26504);
and U32610 (N_32610,N_26072,N_24147);
nor U32611 (N_32611,N_23128,N_28622);
and U32612 (N_32612,N_26576,N_23225);
nor U32613 (N_32613,N_27683,N_20003);
nor U32614 (N_32614,N_28518,N_20283);
and U32615 (N_32615,N_22430,N_26036);
or U32616 (N_32616,N_25194,N_28624);
and U32617 (N_32617,N_21063,N_21649);
nor U32618 (N_32618,N_20596,N_23748);
nand U32619 (N_32619,N_29527,N_20210);
or U32620 (N_32620,N_25514,N_29974);
or U32621 (N_32621,N_28461,N_25443);
or U32622 (N_32622,N_20653,N_28315);
xor U32623 (N_32623,N_25697,N_27554);
and U32624 (N_32624,N_29039,N_29599);
and U32625 (N_32625,N_20339,N_25106);
or U32626 (N_32626,N_21133,N_25599);
or U32627 (N_32627,N_29994,N_23079);
nand U32628 (N_32628,N_20258,N_22728);
nand U32629 (N_32629,N_20771,N_28360);
nor U32630 (N_32630,N_25636,N_27382);
nor U32631 (N_32631,N_27984,N_26600);
or U32632 (N_32632,N_22560,N_27336);
xnor U32633 (N_32633,N_22851,N_25703);
xnor U32634 (N_32634,N_20445,N_22623);
nor U32635 (N_32635,N_25033,N_25855);
xnor U32636 (N_32636,N_20024,N_29065);
or U32637 (N_32637,N_20619,N_21653);
xor U32638 (N_32638,N_26411,N_26662);
and U32639 (N_32639,N_24364,N_21320);
nand U32640 (N_32640,N_27283,N_20031);
nor U32641 (N_32641,N_23789,N_24901);
nand U32642 (N_32642,N_24470,N_29984);
nand U32643 (N_32643,N_24574,N_28637);
and U32644 (N_32644,N_22496,N_29796);
nand U32645 (N_32645,N_25253,N_25803);
and U32646 (N_32646,N_26442,N_24766);
nand U32647 (N_32647,N_29292,N_20336);
or U32648 (N_32648,N_22270,N_23278);
nand U32649 (N_32649,N_23327,N_28218);
nor U32650 (N_32650,N_29725,N_28080);
nor U32651 (N_32651,N_22816,N_21896);
nor U32652 (N_32652,N_21258,N_29628);
nor U32653 (N_32653,N_21481,N_26712);
nor U32654 (N_32654,N_26764,N_21504);
xnor U32655 (N_32655,N_21321,N_27215);
nand U32656 (N_32656,N_24381,N_28929);
and U32657 (N_32657,N_26592,N_28146);
and U32658 (N_32658,N_24984,N_21037);
nor U32659 (N_32659,N_26463,N_29629);
nand U32660 (N_32660,N_20819,N_24293);
and U32661 (N_32661,N_23294,N_21867);
nand U32662 (N_32662,N_26953,N_25436);
and U32663 (N_32663,N_26897,N_29674);
nand U32664 (N_32664,N_26052,N_28500);
and U32665 (N_32665,N_26590,N_20579);
nand U32666 (N_32666,N_20134,N_21950);
and U32667 (N_32667,N_24027,N_25021);
nor U32668 (N_32668,N_20479,N_26665);
or U32669 (N_32669,N_26392,N_23607);
xnor U32670 (N_32670,N_24169,N_28297);
and U32671 (N_32671,N_23461,N_26362);
xor U32672 (N_32672,N_26045,N_22215);
nand U32673 (N_32673,N_28587,N_20448);
or U32674 (N_32674,N_26038,N_28900);
and U32675 (N_32675,N_23751,N_28537);
and U32676 (N_32676,N_22819,N_25529);
and U32677 (N_32677,N_21323,N_22517);
and U32678 (N_32678,N_25804,N_21219);
or U32679 (N_32679,N_20384,N_22028);
and U32680 (N_32680,N_20369,N_28630);
and U32681 (N_32681,N_26526,N_22058);
nand U32682 (N_32682,N_28574,N_23827);
xnor U32683 (N_32683,N_26505,N_24148);
and U32684 (N_32684,N_20968,N_22373);
and U32685 (N_32685,N_24122,N_21419);
nor U32686 (N_32686,N_26530,N_22872);
or U32687 (N_32687,N_20489,N_25799);
or U32688 (N_32688,N_29086,N_23212);
or U32689 (N_32689,N_20588,N_29534);
or U32690 (N_32690,N_20373,N_28961);
nor U32691 (N_32691,N_23796,N_26407);
and U32692 (N_32692,N_28859,N_28559);
xnor U32693 (N_32693,N_24653,N_29703);
and U32694 (N_32694,N_20020,N_26673);
and U32695 (N_32695,N_21274,N_27023);
nor U32696 (N_32696,N_24267,N_28924);
nor U32697 (N_32697,N_24282,N_26909);
nand U32698 (N_32698,N_22469,N_22583);
or U32699 (N_32699,N_29144,N_21613);
and U32700 (N_32700,N_28729,N_26951);
xor U32701 (N_32701,N_29705,N_22069);
nor U32702 (N_32702,N_21708,N_23916);
nor U32703 (N_32703,N_25297,N_23716);
nand U32704 (N_32704,N_23146,N_26149);
or U32705 (N_32705,N_24003,N_22420);
and U32706 (N_32706,N_29157,N_25581);
xor U32707 (N_32707,N_23016,N_26240);
nor U32708 (N_32708,N_28959,N_21456);
nand U32709 (N_32709,N_27966,N_20289);
nor U32710 (N_32710,N_21891,N_24596);
and U32711 (N_32711,N_28157,N_28852);
and U32712 (N_32712,N_26281,N_29306);
and U32713 (N_32713,N_24577,N_28866);
and U32714 (N_32714,N_25100,N_23453);
and U32715 (N_32715,N_21378,N_26219);
xnor U32716 (N_32716,N_26694,N_22691);
xnor U32717 (N_32717,N_28309,N_27342);
nor U32718 (N_32718,N_22839,N_25353);
or U32719 (N_32719,N_27519,N_28970);
and U32720 (N_32720,N_25196,N_21191);
or U32721 (N_32721,N_24568,N_23894);
nand U32722 (N_32722,N_26503,N_23672);
nor U32723 (N_32723,N_20249,N_26455);
or U32724 (N_32724,N_28450,N_26875);
or U32725 (N_32725,N_27212,N_22212);
nand U32726 (N_32726,N_28351,N_20772);
and U32727 (N_32727,N_27325,N_26300);
nand U32728 (N_32728,N_20985,N_29838);
and U32729 (N_32729,N_22280,N_24705);
and U32730 (N_32730,N_24893,N_29778);
nand U32731 (N_32731,N_25919,N_23285);
nor U32732 (N_32732,N_26676,N_20063);
or U32733 (N_32733,N_27145,N_29700);
xor U32734 (N_32734,N_28997,N_23117);
nor U32735 (N_32735,N_28153,N_26261);
nand U32736 (N_32736,N_26218,N_22635);
nand U32737 (N_32737,N_22592,N_20754);
xnor U32738 (N_32738,N_29567,N_23046);
nand U32739 (N_32739,N_21055,N_27132);
or U32740 (N_32740,N_24960,N_25394);
nor U32741 (N_32741,N_23209,N_27709);
nand U32742 (N_32742,N_23459,N_27784);
and U32743 (N_32743,N_27892,N_24400);
xnor U32744 (N_32744,N_25773,N_22708);
nor U32745 (N_32745,N_21587,N_27681);
nor U32746 (N_32746,N_20012,N_21742);
nand U32747 (N_32747,N_21589,N_20275);
nand U32748 (N_32748,N_24967,N_21427);
xor U32749 (N_32749,N_27061,N_24046);
or U32750 (N_32750,N_27108,N_24306);
and U32751 (N_32751,N_23434,N_27606);
nand U32752 (N_32752,N_21002,N_25348);
and U32753 (N_32753,N_24971,N_20069);
nor U32754 (N_32754,N_20513,N_26402);
xnor U32755 (N_32755,N_23763,N_26772);
xnor U32756 (N_32756,N_28068,N_28400);
or U32757 (N_32757,N_23927,N_21537);
and U32758 (N_32758,N_24647,N_20237);
nand U32759 (N_32759,N_22452,N_21703);
and U32760 (N_32760,N_20518,N_28724);
nand U32761 (N_32761,N_29493,N_21543);
xor U32762 (N_32762,N_26296,N_29057);
xnor U32763 (N_32763,N_29505,N_21480);
nand U32764 (N_32764,N_21252,N_24086);
or U32765 (N_32765,N_24013,N_23351);
or U32766 (N_32766,N_21559,N_26024);
nand U32767 (N_32767,N_26154,N_27598);
and U32768 (N_32768,N_25711,N_25800);
nand U32769 (N_32769,N_23320,N_29433);
nor U32770 (N_32770,N_22524,N_20014);
and U32771 (N_32771,N_23701,N_26136);
nor U32772 (N_32772,N_25786,N_20760);
nor U32773 (N_32773,N_25517,N_27810);
or U32774 (N_32774,N_24734,N_22919);
nor U32775 (N_32775,N_21211,N_26710);
nand U32776 (N_32776,N_29653,N_21847);
nand U32777 (N_32777,N_20123,N_23471);
or U32778 (N_32778,N_21753,N_28519);
nand U32779 (N_32779,N_21859,N_26113);
and U32780 (N_32780,N_29511,N_23277);
nor U32781 (N_32781,N_20544,N_24552);
or U32782 (N_32782,N_20932,N_27452);
xor U32783 (N_32783,N_23313,N_21508);
or U32784 (N_32784,N_23138,N_27298);
or U32785 (N_32785,N_21744,N_23930);
and U32786 (N_32786,N_29959,N_25401);
or U32787 (N_32787,N_22208,N_22116);
and U32788 (N_32788,N_28781,N_22922);
nor U32789 (N_32789,N_24898,N_21263);
nor U32790 (N_32790,N_29585,N_27801);
nor U32791 (N_32791,N_21796,N_26253);
and U32792 (N_32792,N_22467,N_29943);
nor U32793 (N_32793,N_21763,N_29429);
nand U32794 (N_32794,N_27788,N_28549);
nand U32795 (N_32795,N_21475,N_22933);
nor U32796 (N_32796,N_26084,N_20091);
and U32797 (N_32797,N_28516,N_25151);
nor U32798 (N_32798,N_23994,N_23250);
xor U32799 (N_32799,N_24339,N_25121);
or U32800 (N_32800,N_28443,N_26695);
and U32801 (N_32801,N_25023,N_28082);
xnor U32802 (N_32802,N_26589,N_25301);
nand U32803 (N_32803,N_27057,N_20356);
and U32804 (N_32804,N_27499,N_22859);
or U32805 (N_32805,N_29331,N_20102);
and U32806 (N_32806,N_27943,N_22785);
nor U32807 (N_32807,N_29130,N_24910);
or U32808 (N_32808,N_25595,N_20496);
and U32809 (N_32809,N_29790,N_24213);
nor U32810 (N_32810,N_20470,N_22548);
nand U32811 (N_32811,N_24016,N_22591);
or U32812 (N_32812,N_27096,N_29769);
nor U32813 (N_32813,N_29446,N_24884);
xnor U32814 (N_32814,N_27609,N_23969);
or U32815 (N_32815,N_28492,N_23194);
nand U32816 (N_32816,N_26513,N_23344);
nand U32817 (N_32817,N_25944,N_20171);
xor U32818 (N_32818,N_24539,N_26325);
nor U32819 (N_32819,N_26220,N_28550);
nor U32820 (N_32820,N_28914,N_24368);
and U32821 (N_32821,N_20510,N_24952);
nor U32822 (N_32822,N_29647,N_21121);
nor U32823 (N_32823,N_29634,N_27566);
or U32824 (N_32824,N_29190,N_27631);
or U32825 (N_32825,N_24610,N_21362);
nand U32826 (N_32826,N_22047,N_21806);
nand U32827 (N_32827,N_25584,N_24580);
nor U32828 (N_32828,N_28904,N_28863);
nand U32829 (N_32829,N_24405,N_26110);
nor U32830 (N_32830,N_26613,N_23318);
nand U32831 (N_32831,N_24416,N_23918);
and U32832 (N_32832,N_23580,N_27971);
or U32833 (N_32833,N_29680,N_21857);
nor U32834 (N_32834,N_23124,N_29615);
or U32835 (N_32835,N_28221,N_28371);
or U32836 (N_32836,N_26757,N_22668);
or U32837 (N_32837,N_22362,N_27463);
and U32838 (N_32838,N_28795,N_25386);
xnor U32839 (N_32839,N_27879,N_20200);
xor U32840 (N_32840,N_23311,N_23667);
or U32841 (N_32841,N_22035,N_27783);
xor U32842 (N_32842,N_20022,N_25402);
nand U32843 (N_32843,N_26030,N_26838);
nand U32844 (N_32844,N_28442,N_29709);
and U32845 (N_32845,N_28936,N_26883);
and U32846 (N_32846,N_26285,N_20457);
nand U32847 (N_32847,N_24520,N_24346);
and U32848 (N_32848,N_20935,N_25313);
and U32849 (N_32849,N_21291,N_27721);
nand U32850 (N_32850,N_21688,N_25962);
and U32851 (N_32851,N_29577,N_27502);
xor U32852 (N_32852,N_25145,N_21059);
nand U32853 (N_32853,N_26528,N_20658);
and U32854 (N_32854,N_20027,N_25521);
xnor U32855 (N_32855,N_26780,N_23982);
nand U32856 (N_32856,N_23950,N_23698);
and U32857 (N_32857,N_28248,N_28177);
or U32858 (N_32858,N_26466,N_29189);
or U32859 (N_32859,N_28200,N_28646);
nand U32860 (N_32860,N_28705,N_20286);
or U32861 (N_32861,N_26675,N_28138);
or U32862 (N_32862,N_23592,N_27777);
and U32863 (N_32863,N_29808,N_26758);
or U32864 (N_32864,N_23799,N_28282);
xor U32865 (N_32865,N_21092,N_24949);
xnor U32866 (N_32866,N_23023,N_21973);
xnor U32867 (N_32867,N_20907,N_20084);
and U32868 (N_32868,N_27366,N_27807);
or U32869 (N_32869,N_21432,N_23100);
xnor U32870 (N_32870,N_24729,N_26335);
nand U32871 (N_32871,N_20523,N_27379);
nor U32872 (N_32872,N_26844,N_23084);
or U32873 (N_32873,N_20893,N_21577);
nand U32874 (N_32874,N_26977,N_28960);
or U32875 (N_32875,N_21348,N_28520);
or U32876 (N_32876,N_23880,N_23207);
nor U32877 (N_32877,N_29830,N_23301);
or U32878 (N_32878,N_27450,N_22160);
nand U32879 (N_32879,N_25533,N_21395);
nor U32880 (N_32880,N_25978,N_25414);
or U32881 (N_32881,N_25574,N_21871);
nor U32882 (N_32882,N_21760,N_25309);
nor U32883 (N_32883,N_22262,N_21681);
nand U32884 (N_32884,N_26739,N_20173);
xor U32885 (N_32885,N_20301,N_29726);
nor U32886 (N_32886,N_27063,N_23299);
or U32887 (N_32887,N_26013,N_22100);
or U32888 (N_32888,N_22306,N_27347);
and U32889 (N_32889,N_23095,N_22135);
nand U32890 (N_32890,N_23811,N_24451);
and U32891 (N_32891,N_20883,N_28240);
nor U32892 (N_32892,N_25993,N_28963);
nand U32893 (N_32893,N_29151,N_22520);
and U32894 (N_32894,N_20256,N_23998);
nand U32895 (N_32895,N_23587,N_25118);
and U32896 (N_32896,N_21562,N_20278);
nor U32897 (N_32897,N_25231,N_22256);
nor U32898 (N_32898,N_22946,N_23054);
and U32899 (N_32899,N_27802,N_28314);
and U32900 (N_32900,N_27235,N_23206);
nand U32901 (N_32901,N_25269,N_29759);
or U32902 (N_32902,N_28301,N_26277);
nand U32903 (N_32903,N_25026,N_20211);
nand U32904 (N_32904,N_24156,N_25801);
xnor U32905 (N_32905,N_21082,N_25602);
nor U32906 (N_32906,N_26657,N_22177);
and U32907 (N_32907,N_29406,N_26532);
or U32908 (N_32908,N_26881,N_28695);
nor U32909 (N_32909,N_29108,N_24203);
and U32910 (N_32910,N_20564,N_24369);
and U32911 (N_32911,N_20359,N_25190);
or U32912 (N_32912,N_20853,N_21181);
or U32913 (N_32913,N_27105,N_20829);
or U32914 (N_32914,N_24989,N_28667);
nand U32915 (N_32915,N_25321,N_26536);
or U32916 (N_32916,N_28215,N_20483);
or U32917 (N_32917,N_27877,N_21437);
and U32918 (N_32918,N_29598,N_20013);
xor U32919 (N_32919,N_28604,N_28513);
xnor U32920 (N_32920,N_29355,N_21146);
nand U32921 (N_32921,N_21966,N_25895);
and U32922 (N_32922,N_29517,N_29371);
and U32923 (N_32923,N_26237,N_27881);
and U32924 (N_32924,N_24956,N_20866);
and U32925 (N_32925,N_23112,N_24802);
xnor U32926 (N_32926,N_24164,N_27468);
nor U32927 (N_32927,N_29807,N_25296);
nand U32928 (N_32928,N_20679,N_20741);
nand U32929 (N_32929,N_25709,N_20464);
nor U32930 (N_32930,N_29454,N_28987);
nand U32931 (N_32931,N_23542,N_21275);
nand U32932 (N_32932,N_22975,N_22329);
and U32933 (N_32933,N_27090,N_25403);
nor U32934 (N_32934,N_28452,N_26837);
nand U32935 (N_32935,N_23334,N_25772);
nor U32936 (N_32936,N_29420,N_26548);
nor U32937 (N_32937,N_27401,N_22093);
nand U32938 (N_32938,N_26161,N_26718);
nor U32939 (N_32939,N_22331,N_26797);
or U32940 (N_32940,N_27550,N_25373);
and U32941 (N_32941,N_25736,N_25438);
or U32942 (N_32942,N_29294,N_26338);
and U32943 (N_32943,N_26206,N_26002);
nand U32944 (N_32944,N_29006,N_25973);
nand U32945 (N_32945,N_25880,N_26198);
xnor U32946 (N_32946,N_21144,N_22311);
and U32947 (N_32947,N_29661,N_21034);
or U32948 (N_32948,N_27621,N_22352);
nand U32949 (N_32949,N_22082,N_20157);
nor U32950 (N_32950,N_28129,N_25723);
or U32951 (N_32951,N_22717,N_28328);
nor U32952 (N_32952,N_21020,N_21893);
and U32953 (N_32953,N_24006,N_27823);
nand U32954 (N_32954,N_23839,N_24515);
xor U32955 (N_32955,N_28178,N_28688);
or U32956 (N_32956,N_24755,N_26939);
nor U32957 (N_32957,N_26998,N_23800);
nand U32958 (N_32958,N_22981,N_20934);
and U32959 (N_32959,N_25771,N_21735);
or U32960 (N_32960,N_25751,N_23728);
and U32961 (N_32961,N_21235,N_28625);
and U32962 (N_32962,N_21242,N_20708);
nor U32963 (N_32963,N_28184,N_23496);
and U32964 (N_32964,N_24229,N_21255);
or U32965 (N_32965,N_25898,N_27226);
nand U32966 (N_32966,N_27078,N_25105);
and U32967 (N_32967,N_26417,N_25366);
nand U32968 (N_32968,N_21477,N_21003);
nor U32969 (N_32969,N_26288,N_28363);
nor U32970 (N_32970,N_29643,N_20372);
and U32971 (N_32971,N_27141,N_29516);
or U32972 (N_32972,N_25063,N_27805);
nand U32973 (N_32973,N_24692,N_28402);
nor U32974 (N_32974,N_26785,N_22190);
or U32975 (N_32975,N_25955,N_27197);
nor U32976 (N_32976,N_26586,N_22365);
xor U32977 (N_32977,N_21527,N_27168);
nand U32978 (N_32978,N_27118,N_21636);
and U32979 (N_32979,N_27941,N_21474);
nor U32980 (N_32980,N_20831,N_26028);
nand U32981 (N_32981,N_20599,N_25507);
and U32982 (N_32982,N_21601,N_23437);
or U32983 (N_32983,N_22110,N_20861);
or U32984 (N_32984,N_28930,N_26497);
or U32985 (N_32985,N_21233,N_23328);
or U32986 (N_32986,N_27422,N_29028);
and U32987 (N_32987,N_27899,N_27300);
nand U32988 (N_32988,N_28708,N_21260);
xnor U32989 (N_32989,N_20534,N_23284);
nor U32990 (N_32990,N_21425,N_28183);
and U32991 (N_32991,N_20279,N_20059);
and U32992 (N_32992,N_25985,N_21579);
nor U32993 (N_32993,N_29136,N_26077);
and U32994 (N_32994,N_26073,N_25968);
nand U32995 (N_32995,N_22779,N_24082);
nor U32996 (N_32996,N_29091,N_28238);
nor U32997 (N_32997,N_28710,N_21854);
xnor U32998 (N_32998,N_29055,N_24494);
nor U32999 (N_32999,N_25335,N_29910);
or U33000 (N_33000,N_28581,N_23705);
and U33001 (N_33001,N_29100,N_21042);
or U33002 (N_33002,N_25561,N_21573);
nor U33003 (N_33003,N_29625,N_22928);
xnor U33004 (N_33004,N_24331,N_29673);
and U33005 (N_33005,N_25357,N_23793);
nand U33006 (N_33006,N_28955,N_22977);
nor U33007 (N_33007,N_28110,N_28773);
nor U33008 (N_33008,N_20183,N_20493);
and U33009 (N_33009,N_24525,N_29707);
and U33010 (N_33010,N_22451,N_29497);
nand U33011 (N_33011,N_26776,N_24036);
or U33012 (N_33012,N_22557,N_23441);
or U33013 (N_33013,N_21757,N_22529);
and U33014 (N_33014,N_22034,N_25280);
xnor U33015 (N_33015,N_21345,N_27959);
or U33016 (N_33016,N_20175,N_28504);
nor U33017 (N_33017,N_23022,N_20573);
nor U33018 (N_33018,N_24334,N_23595);
and U33019 (N_33019,N_27213,N_23488);
xor U33020 (N_33020,N_23742,N_24944);
or U33021 (N_33021,N_23596,N_27956);
or U33022 (N_33022,N_29146,N_28474);
and U33023 (N_33023,N_25134,N_28746);
or U33024 (N_33024,N_22765,N_24316);
nand U33025 (N_33025,N_21923,N_27394);
xor U33026 (N_33026,N_23520,N_22075);
nand U33027 (N_33027,N_22550,N_27625);
and U33028 (N_33028,N_28925,N_25564);
xnor U33029 (N_33029,N_22471,N_26421);
xnor U33030 (N_33030,N_28213,N_21489);
nand U33031 (N_33031,N_25150,N_26771);
or U33032 (N_33032,N_22736,N_26341);
nand U33033 (N_33033,N_20957,N_24608);
or U33034 (N_33034,N_26354,N_22320);
nand U33035 (N_33035,N_22421,N_26266);
nand U33036 (N_33036,N_25603,N_20310);
and U33037 (N_33037,N_26870,N_26390);
nand U33038 (N_33038,N_22997,N_20442);
nand U33039 (N_33039,N_24730,N_22840);
nand U33040 (N_33040,N_29510,N_21907);
nor U33041 (N_33041,N_23876,N_25192);
nor U33042 (N_33042,N_24228,N_24488);
nand U33043 (N_33043,N_22332,N_27232);
xor U33044 (N_33044,N_26488,N_21600);
xor U33045 (N_33045,N_29963,N_21542);
xor U33046 (N_33046,N_22364,N_20781);
nand U33047 (N_33047,N_22056,N_20580);
nor U33048 (N_33048,N_21727,N_29453);
and U33049 (N_33049,N_25781,N_24176);
and U33050 (N_33050,N_27886,N_20933);
or U33051 (N_33051,N_29412,N_26091);
xnor U33052 (N_33052,N_28470,N_21569);
nor U33053 (N_33053,N_26246,N_24064);
or U33054 (N_33054,N_23745,N_25404);
and U33055 (N_33055,N_23573,N_26271);
nand U33056 (N_33056,N_25392,N_21270);
or U33057 (N_33057,N_27271,N_20964);
nand U33058 (N_33058,N_22027,N_28486);
nand U33059 (N_33059,N_24808,N_21978);
xor U33060 (N_33060,N_28375,N_21890);
and U33061 (N_33061,N_24720,N_22820);
or U33062 (N_33062,N_29208,N_22344);
nand U33063 (N_33063,N_24490,N_21841);
or U33064 (N_33064,N_20433,N_22092);
nand U33065 (N_33065,N_22271,N_26454);
or U33066 (N_33066,N_24882,N_29501);
nand U33067 (N_33067,N_25640,N_21455);
nand U33068 (N_33068,N_20551,N_26375);
or U33069 (N_33069,N_26186,N_29205);
or U33070 (N_33070,N_26936,N_26542);
and U33071 (N_33071,N_25018,N_21495);
nand U33072 (N_33072,N_29591,N_29393);
and U33073 (N_33073,N_20788,N_21368);
nor U33074 (N_33074,N_23721,N_27963);
nor U33075 (N_33075,N_28984,N_23264);
nand U33076 (N_33076,N_28834,N_23019);
and U33077 (N_33077,N_27328,N_29405);
xnor U33078 (N_33078,N_23537,N_22903);
xnor U33079 (N_33079,N_29649,N_20481);
nand U33080 (N_33080,N_23042,N_23289);
nor U33081 (N_33081,N_27610,N_23835);
nor U33082 (N_33082,N_29359,N_20226);
nor U33083 (N_33083,N_23090,N_22078);
or U33084 (N_33084,N_22435,N_29225);
nor U33085 (N_33085,N_28263,N_29441);
and U33086 (N_33086,N_28488,N_25763);
or U33087 (N_33087,N_25124,N_27957);
and U33088 (N_33088,N_23122,N_26986);
and U33089 (N_33089,N_26611,N_20392);
nand U33090 (N_33090,N_20167,N_29886);
nor U33091 (N_33091,N_23550,N_28809);
xnor U33092 (N_33092,N_20982,N_29009);
or U33093 (N_33093,N_23847,N_27842);
nor U33094 (N_33094,N_28175,N_24107);
and U33095 (N_33095,N_29145,N_26021);
nand U33096 (N_33096,N_28005,N_23464);
and U33097 (N_33097,N_26040,N_28325);
and U33098 (N_33098,N_24631,N_20576);
and U33099 (N_33099,N_20207,N_21246);
nand U33100 (N_33100,N_24192,N_28427);
nand U33101 (N_33101,N_27236,N_20749);
xor U33102 (N_33102,N_24380,N_26057);
nand U33103 (N_33103,N_22239,N_28451);
nand U33104 (N_33104,N_28176,N_25245);
and U33105 (N_33105,N_25396,N_20662);
or U33106 (N_33106,N_21810,N_24683);
and U33107 (N_33107,N_26593,N_25260);
and U33108 (N_33108,N_23656,N_25558);
nor U33109 (N_33109,N_25205,N_22867);
or U33110 (N_33110,N_29844,N_26453);
nand U33111 (N_33111,N_23844,N_24233);
or U33112 (N_33112,N_29999,N_21980);
nor U33113 (N_33113,N_26027,N_24987);
xnor U33114 (N_33114,N_23613,N_24033);
nor U33115 (N_33115,N_27875,N_25418);
and U33116 (N_33116,N_26678,N_22080);
and U33117 (N_33117,N_24965,N_24540);
nand U33118 (N_33118,N_27003,N_28726);
and U33119 (N_33119,N_29211,N_26456);
and U33120 (N_33120,N_27354,N_23096);
nor U33121 (N_33121,N_25211,N_20379);
nand U33122 (N_33122,N_24000,N_25320);
or U33123 (N_33123,N_25116,N_29449);
xor U33124 (N_33124,N_22106,N_24005);
nor U33125 (N_33125,N_29058,N_20492);
xnor U33126 (N_33126,N_22572,N_25114);
nor U33127 (N_33127,N_22578,N_29774);
nor U33128 (N_33128,N_25168,N_23619);
and U33129 (N_33129,N_22349,N_25074);
or U33130 (N_33130,N_21236,N_22587);
and U33131 (N_33131,N_23962,N_26863);
and U33132 (N_33132,N_29176,N_22358);
and U33133 (N_33133,N_25646,N_27467);
nand U33134 (N_33134,N_20139,N_23137);
or U33135 (N_33135,N_22983,N_21231);
or U33136 (N_33136,N_22272,N_21880);
or U33137 (N_33137,N_23532,N_20180);
nor U33138 (N_33138,N_21415,N_27178);
nor U33139 (N_33139,N_24137,N_20215);
nand U33140 (N_33140,N_23555,N_20645);
nand U33141 (N_33141,N_28681,N_26587);
nand U33142 (N_33142,N_25824,N_29072);
and U33143 (N_33143,N_23486,N_27284);
nor U33144 (N_33144,N_27528,N_21672);
nor U33145 (N_33145,N_28647,N_29030);
and U33146 (N_33146,N_23379,N_24056);
and U33147 (N_33147,N_21952,N_21585);
nor U33148 (N_33148,N_27420,N_28089);
and U33149 (N_33149,N_27633,N_27410);
nor U33150 (N_33150,N_29940,N_25916);
nor U33151 (N_33151,N_20628,N_25789);
nand U33152 (N_33152,N_24379,N_26273);
nand U33153 (N_33153,N_20108,N_20146);
xnor U33154 (N_33154,N_21340,N_22294);
xnor U33155 (N_33155,N_23494,N_26358);
nor U33156 (N_33156,N_27314,N_28870);
nor U33157 (N_33157,N_26962,N_22927);
nor U33158 (N_33158,N_25812,N_26955);
and U33159 (N_33159,N_22203,N_24423);
and U33160 (N_33160,N_26749,N_24493);
or U33161 (N_33161,N_27549,N_24491);
xnor U33162 (N_33162,N_26584,N_22474);
xnor U33163 (N_33163,N_29760,N_28406);
and U33164 (N_33164,N_20533,N_21113);
and U33165 (N_33165,N_27449,N_27967);
and U33166 (N_33166,N_23850,N_24513);
nor U33167 (N_33167,N_28081,N_23093);
nor U33168 (N_33168,N_29688,N_26080);
and U33169 (N_33169,N_23654,N_23744);
nand U33170 (N_33170,N_28481,N_21756);
and U33171 (N_33171,N_24477,N_22136);
nand U33172 (N_33172,N_28167,N_26544);
or U33173 (N_33173,N_24187,N_28701);
xor U33174 (N_33174,N_20660,N_28132);
and U33175 (N_33175,N_28652,N_22596);
nand U33176 (N_33176,N_29691,N_29663);
or U33177 (N_33177,N_25868,N_23133);
nand U33178 (N_33178,N_28242,N_22370);
nand U33179 (N_33179,N_25284,N_20030);
and U33180 (N_33180,N_26208,N_20971);
nand U33181 (N_33181,N_22784,N_28816);
nor U33182 (N_33182,N_26756,N_27613);
nor U33183 (N_33183,N_26742,N_27725);
nor U33184 (N_33184,N_25308,N_21905);
nand U33185 (N_33185,N_24877,N_22905);
nand U33186 (N_33186,N_29066,N_21363);
and U33187 (N_33187,N_25146,N_24973);
xor U33188 (N_33188,N_28690,N_25980);
or U33189 (N_33189,N_23963,N_24395);
nand U33190 (N_33190,N_26178,N_24934);
nor U33191 (N_33191,N_26127,N_20320);
nor U33192 (N_33192,N_26878,N_27016);
nor U33193 (N_33193,N_21210,N_22497);
and U33194 (N_33194,N_20644,N_23481);
or U33195 (N_33195,N_20828,N_22347);
xor U33196 (N_33196,N_25725,N_20950);
and U33197 (N_33197,N_27985,N_27303);
nor U33198 (N_33198,N_27690,N_29480);
or U33199 (N_33199,N_25717,N_20058);
nand U33200 (N_33200,N_24058,N_25278);
or U33201 (N_33201,N_24800,N_20078);
xor U33202 (N_33202,N_27230,N_28894);
nand U33203 (N_33203,N_29960,N_27058);
nor U33204 (N_33204,N_22535,N_20718);
and U33205 (N_33205,N_28540,N_22020);
or U33206 (N_33206,N_26981,N_23579);
or U33207 (N_33207,N_26882,N_21138);
nand U33208 (N_33208,N_29664,N_23123);
nor U33209 (N_33209,N_29765,N_27009);
xnor U33210 (N_33210,N_27755,N_20469);
and U33211 (N_33211,N_29160,N_24394);
nand U33212 (N_33212,N_24103,N_29008);
or U33213 (N_33213,N_28121,N_21761);
or U33214 (N_33214,N_26015,N_27060);
and U33215 (N_33215,N_24937,N_21441);
nor U33216 (N_33216,N_27799,N_24155);
and U33217 (N_33217,N_29839,N_26894);
xor U33218 (N_33218,N_20918,N_22741);
or U33219 (N_33219,N_29440,N_25349);
nor U33220 (N_33220,N_23140,N_22374);
nand U33221 (N_33221,N_29627,N_27324);
nand U33222 (N_33222,N_24704,N_25136);
nor U33223 (N_33223,N_25846,N_20867);
nand U33224 (N_33224,N_22653,N_21706);
xnor U33225 (N_33225,N_27373,N_20219);
nand U33226 (N_33226,N_28756,N_23879);
nand U33227 (N_33227,N_23391,N_27607);
xor U33228 (N_33228,N_20634,N_23819);
and U33229 (N_33229,N_27759,N_29319);
xnor U33230 (N_33230,N_26815,N_23584);
xor U33231 (N_33231,N_21937,N_25817);
nand U33232 (N_33232,N_20652,N_22917);
nor U33233 (N_33233,N_25634,N_29031);
nor U33234 (N_33234,N_20323,N_29445);
or U33235 (N_33235,N_26700,N_27940);
nand U33236 (N_33236,N_26224,N_23875);
nor U33237 (N_33237,N_26753,N_25277);
and U33238 (N_33238,N_28037,N_23708);
or U33239 (N_33239,N_28163,N_20631);
and U33240 (N_33240,N_22325,N_24296);
or U33241 (N_33241,N_25350,N_25351);
and U33242 (N_33242,N_29955,N_25358);
nand U33243 (N_33243,N_27035,N_27514);
and U33244 (N_33244,N_20695,N_20970);
and U33245 (N_33245,N_26276,N_21429);
nand U33246 (N_33246,N_23111,N_20195);
xor U33247 (N_33247,N_25816,N_29751);
and U33248 (N_33248,N_23631,N_21466);
nor U33249 (N_33249,N_22958,N_26467);
nand U33250 (N_33250,N_27601,N_27025);
nor U33251 (N_33251,N_21382,N_28848);
nand U33252 (N_33252,N_29600,N_24292);
nand U33253 (N_33253,N_21167,N_29583);
xor U33254 (N_33254,N_24248,N_24921);
or U33255 (N_33255,N_25087,N_29819);
or U33256 (N_33256,N_22705,N_28289);
nand U33257 (N_33257,N_28374,N_29545);
or U33258 (N_33258,N_29379,N_28216);
nand U33259 (N_33259,N_28148,N_20304);
or U33260 (N_33260,N_25238,N_28569);
and U33261 (N_33261,N_26514,N_25498);
nor U33262 (N_33262,N_27659,N_28534);
and U33263 (N_33263,N_24966,N_20927);
or U33264 (N_33264,N_23887,N_23286);
or U33265 (N_33265,N_21479,N_23150);
or U33266 (N_33266,N_20197,N_27591);
xnor U33267 (N_33267,N_27327,N_20140);
nand U33268 (N_33268,N_29979,N_27085);
xor U33269 (N_33269,N_21145,N_22724);
and U33270 (N_33270,N_25937,N_23446);
xnor U33271 (N_33271,N_23964,N_29945);
nand U33272 (N_33272,N_29357,N_25165);
or U33273 (N_33273,N_23232,N_23709);
xor U33274 (N_33274,N_24859,N_24329);
nor U33275 (N_33275,N_24896,N_27552);
nor U33276 (N_33276,N_22350,N_27854);
xor U33277 (N_33277,N_26207,N_27617);
or U33278 (N_33278,N_28800,N_22209);
or U33279 (N_33279,N_27127,N_27006);
nand U33280 (N_33280,N_28605,N_25103);
and U33281 (N_33281,N_20131,N_25153);
nor U33282 (N_33282,N_25204,N_25825);
nor U33283 (N_33283,N_26669,N_28626);
xnor U33284 (N_33284,N_28115,N_24619);
nor U33285 (N_33285,N_26524,N_24311);
and U33286 (N_33286,N_24938,N_24733);
nand U33287 (N_33287,N_23498,N_28941);
nand U33288 (N_33288,N_25317,N_23616);
nor U33289 (N_33289,N_27876,N_27288);
nor U33290 (N_33290,N_22313,N_21955);
or U33291 (N_33291,N_28845,N_25619);
nor U33292 (N_33292,N_20351,N_28207);
or U33293 (N_33293,N_22381,N_20397);
and U33294 (N_33294,N_24837,N_22604);
xor U33295 (N_33295,N_27774,N_20068);
or U33296 (N_33296,N_28797,N_26249);
and U33297 (N_33297,N_22013,N_29033);
nor U33298 (N_33298,N_26380,N_28820);
nand U33299 (N_33299,N_27921,N_22907);
nor U33300 (N_33300,N_28191,N_27924);
or U33301 (N_33301,N_24701,N_29722);
xnor U33302 (N_33302,N_28471,N_25760);
and U33303 (N_33303,N_26361,N_29431);
or U33304 (N_33304,N_29267,N_21619);
and U33305 (N_33305,N_26533,N_26339);
or U33306 (N_33306,N_22871,N_24750);
xor U33307 (N_33307,N_29194,N_22674);
and U33308 (N_33308,N_27051,N_23939);
and U33309 (N_33309,N_22187,N_25891);
or U33310 (N_33310,N_24651,N_22077);
and U33311 (N_33311,N_22625,N_27195);
nor U33312 (N_33312,N_23628,N_25681);
nor U33313 (N_33313,N_23945,N_22073);
nor U33314 (N_33314,N_21818,N_26719);
nor U33315 (N_33315,N_21933,N_24376);
nor U33316 (N_33316,N_25682,N_28946);
and U33317 (N_33317,N_25859,N_20057);
nand U33318 (N_33318,N_21831,N_26495);
or U33319 (N_33319,N_29731,N_25336);
nand U33320 (N_33320,N_26686,N_28378);
nand U33321 (N_33321,N_22112,N_28197);
and U33322 (N_33322,N_29367,N_20739);
and U33323 (N_33323,N_23153,N_22416);
nand U33324 (N_33324,N_21836,N_21737);
nand U33325 (N_33325,N_29399,N_21645);
and U33326 (N_33326,N_29857,N_23390);
nand U33327 (N_33327,N_26128,N_23118);
nor U33328 (N_33328,N_28004,N_28185);
nand U33329 (N_33329,N_29478,N_21416);
nand U33330 (N_33330,N_28673,N_22453);
nand U33331 (N_33331,N_22074,N_27479);
and U33332 (N_33332,N_27233,N_20922);
nand U33333 (N_33333,N_28306,N_26927);
or U33334 (N_33334,N_27841,N_28499);
or U33335 (N_33335,N_21009,N_24983);
xor U33336 (N_33336,N_26286,N_29622);
and U33337 (N_33337,N_28235,N_20880);
and U33338 (N_33338,N_24655,N_28802);
xnor U33339 (N_33339,N_23645,N_27983);
and U33340 (N_33340,N_28881,N_21276);
or U33341 (N_33341,N_25904,N_22394);
or U33342 (N_33342,N_21300,N_25185);
nor U33343 (N_33343,N_26787,N_27285);
xor U33344 (N_33344,N_27691,N_22873);
and U33345 (N_33345,N_21895,N_29757);
nand U33346 (N_33346,N_28988,N_22289);
or U33347 (N_33347,N_25417,N_26355);
or U33348 (N_33348,N_20642,N_20043);
nand U33349 (N_33349,N_27114,N_24444);
xnor U33350 (N_33350,N_22174,N_22447);
nand U33351 (N_33351,N_20381,N_27747);
nor U33352 (N_33352,N_26357,N_20439);
xor U33353 (N_33353,N_29202,N_21555);
or U33354 (N_33354,N_25246,N_21195);
and U33355 (N_33355,N_23724,N_27752);
and U33356 (N_33356,N_21853,N_28372);
or U33357 (N_33357,N_21344,N_29870);
and U33358 (N_33358,N_24397,N_29566);
nor U33359 (N_33359,N_29396,N_20364);
and U33360 (N_33360,N_24789,N_29710);
nor U33361 (N_33361,N_24126,N_25052);
nand U33362 (N_33362,N_27019,N_25209);
nor U33363 (N_33363,N_21682,N_24051);
nor U33364 (N_33364,N_22575,N_21618);
nand U33365 (N_33365,N_28340,N_27179);
and U33366 (N_33366,N_26685,N_26352);
nand U33367 (N_33367,N_28250,N_25757);
xnor U33368 (N_33368,N_27490,N_27989);
nand U33369 (N_33369,N_20152,N_24454);
and U33370 (N_33370,N_23794,N_23912);
or U33371 (N_33371,N_24204,N_24603);
nand U33372 (N_33372,N_24489,N_22510);
or U33373 (N_33373,N_20424,N_27374);
nor U33374 (N_33374,N_23062,N_25930);
nand U33375 (N_33375,N_21525,N_28389);
or U33376 (N_33376,N_25061,N_26212);
nor U33377 (N_33377,N_22475,N_26670);
xnor U33378 (N_33378,N_28100,N_29975);
and U33379 (N_33379,N_27608,N_27199);
nand U33380 (N_33380,N_25152,N_29770);
and U33381 (N_33381,N_20944,N_20327);
nand U33382 (N_33382,N_22957,N_29689);
xor U33383 (N_33383,N_25745,N_23792);
or U33384 (N_33384,N_21745,N_20729);
or U33385 (N_33385,N_26760,N_25842);
nand U33386 (N_33386,N_22229,N_25732);
or U33387 (N_33387,N_29370,N_27498);
nor U33388 (N_33388,N_23531,N_26457);
and U33389 (N_33389,N_25702,N_26350);
nand U33390 (N_33390,N_23378,N_20914);
and U33391 (N_33391,N_28436,N_27289);
nand U33392 (N_33392,N_22789,N_22798);
or U33393 (N_33393,N_24662,N_24230);
nand U33394 (N_33394,N_28342,N_20113);
nand U33395 (N_33395,N_23369,N_21943);
or U33396 (N_33396,N_27667,N_29609);
and U33397 (N_33397,N_22806,N_28335);
nand U33398 (N_33398,N_29929,N_22060);
and U33399 (N_33399,N_28166,N_29626);
xor U33400 (N_33400,N_21026,N_28791);
nand U33401 (N_33401,N_27038,N_20465);
xnor U33402 (N_33402,N_21724,N_24518);
or U33403 (N_33403,N_20860,N_23822);
and U33404 (N_33404,N_25635,N_21257);
nand U33405 (N_33405,N_22671,N_27800);
nor U33406 (N_33406,N_28326,N_29479);
and U33407 (N_33407,N_24172,N_24314);
nor U33408 (N_33408,N_27073,N_29186);
or U33409 (N_33409,N_29876,N_27510);
or U33410 (N_33410,N_24007,N_27890);
or U33411 (N_33411,N_20235,N_26062);
and U33412 (N_33412,N_22083,N_23332);
or U33413 (N_33413,N_25568,N_21303);
xnor U33414 (N_33414,N_21863,N_29853);
and U33415 (N_33415,N_28823,N_20792);
nand U33416 (N_33416,N_27087,N_22727);
or U33417 (N_33417,N_25385,N_21385);
nor U33418 (N_33418,N_25266,N_27160);
and U33419 (N_33419,N_28638,N_24825);
or U33420 (N_33420,N_20946,N_23611);
nand U33421 (N_33421,N_27511,N_23669);
nor U33422 (N_33422,N_21969,N_25006);
or U33423 (N_33423,N_20770,N_20963);
or U33424 (N_33424,N_28269,N_27790);
or U33425 (N_33425,N_27412,N_20872);
or U33426 (N_33426,N_23737,N_25044);
nand U33427 (N_33427,N_25684,N_24764);
nor U33428 (N_33428,N_28828,N_25972);
nor U33429 (N_33429,N_20225,N_20050);
or U33430 (N_33430,N_26755,N_23251);
nor U33431 (N_33431,N_20842,N_22050);
xor U33432 (N_33432,N_22334,N_27189);
nor U33433 (N_33433,N_28903,N_28180);
nor U33434 (N_33434,N_28182,N_24060);
nor U33435 (N_33435,N_22448,N_27944);
xor U33436 (N_33436,N_23180,N_26527);
nor U33437 (N_33437,N_22443,N_24994);
xor U33438 (N_33438,N_25258,N_21592);
and U33439 (N_33439,N_26291,N_24751);
xor U33440 (N_33440,N_27952,N_27047);
or U33441 (N_33441,N_25995,N_23503);
nand U33442 (N_33442,N_20766,N_25796);
or U33443 (N_33443,N_21401,N_25019);
and U33444 (N_33444,N_22356,N_29481);
nand U33445 (N_33445,N_20605,N_20751);
and U33446 (N_33446,N_21944,N_25148);
and U33447 (N_33447,N_24106,N_29631);
xor U33448 (N_33448,N_29311,N_29575);
xor U33449 (N_33449,N_23109,N_26368);
or U33450 (N_33450,N_28198,N_24866);
xnor U33451 (N_33451,N_20538,N_21609);
nor U33452 (N_33452,N_22966,N_23040);
and U33453 (N_33453,N_24502,N_29933);
or U33454 (N_33454,N_28145,N_22353);
nand U33455 (N_33455,N_27329,N_20383);
nor U33456 (N_33456,N_24581,N_22269);
nand U33457 (N_33457,N_21359,N_21284);
and U33458 (N_33458,N_24453,N_25864);
nor U33459 (N_33459,N_24801,N_26525);
and U33460 (N_33460,N_20637,N_21915);
nor U33461 (N_33461,N_23339,N_27975);
and U33462 (N_33462,N_24656,N_22431);
and U33463 (N_33463,N_24679,N_20669);
and U33464 (N_33464,N_23014,N_23085);
xnor U33465 (N_33465,N_28714,N_27027);
or U33466 (N_33466,N_21212,N_24231);
and U33467 (N_33467,N_28783,N_20115);
and U33468 (N_33468,N_29437,N_21039);
or U33469 (N_33469,N_25598,N_24223);
xnor U33470 (N_33470,N_20716,N_29898);
xnor U33471 (N_33471,N_24723,N_27496);
nor U33472 (N_33472,N_27889,N_26952);
nand U33473 (N_33473,N_26917,N_24012);
nor U33474 (N_33474,N_24431,N_29749);
or U33475 (N_33475,N_20293,N_20008);
nor U33476 (N_33476,N_28172,N_21882);
xnor U33477 (N_33477,N_26534,N_26496);
or U33478 (N_33478,N_27693,N_28916);
nor U33479 (N_33479,N_23518,N_23469);
or U33480 (N_33480,N_20620,N_27206);
nor U33481 (N_33481,N_28495,N_25600);
or U33482 (N_33482,N_21164,N_20478);
nor U33483 (N_33483,N_27816,N_27616);
nor U33484 (N_33484,N_25481,N_24854);
nor U33485 (N_33485,N_29841,N_23491);
and U33486 (N_33486,N_29916,N_22258);
or U33487 (N_33487,N_29317,N_22711);
or U33488 (N_33488,N_29272,N_21567);
nand U33489 (N_33489,N_22962,N_24878);
nand U33490 (N_33490,N_28254,N_25892);
nand U33491 (N_33491,N_20477,N_24037);
nor U33492 (N_33492,N_26941,N_24390);
and U33493 (N_33493,N_23922,N_20941);
nor U33494 (N_33494,N_20252,N_21834);
xnor U33495 (N_33495,N_23493,N_29810);
or U33496 (N_33496,N_27988,N_20269);
nor U33497 (N_33497,N_23837,N_20562);
nor U33498 (N_33498,N_27447,N_29771);
nor U33499 (N_33499,N_23915,N_27980);
or U33500 (N_33500,N_24505,N_23208);
or U33501 (N_33501,N_28188,N_24601);
and U33502 (N_33502,N_24805,N_21861);
or U33503 (N_33503,N_20179,N_22713);
or U33504 (N_33504,N_21876,N_22440);
nand U33505 (N_33505,N_25042,N_24183);
nor U33506 (N_33506,N_24811,N_26491);
nand U33507 (N_33507,N_29676,N_27296);
and U33508 (N_33508,N_29806,N_26134);
and U33509 (N_33509,N_28165,N_26802);
nand U33510 (N_33510,N_21174,N_23813);
or U33511 (N_33511,N_27119,N_29941);
xnor U33512 (N_33512,N_24671,N_25821);
and U33513 (N_33513,N_26682,N_25157);
nor U33514 (N_33514,N_20410,N_27185);
or U33515 (N_33515,N_21974,N_24885);
and U33516 (N_33516,N_27663,N_27705);
or U33517 (N_33517,N_23104,N_22068);
or U33518 (N_33518,N_20569,N_23343);
nor U33519 (N_33519,N_24337,N_24970);
or U33520 (N_33520,N_24972,N_26093);
and U33521 (N_33521,N_21273,N_26019);
nand U33522 (N_33522,N_23615,N_29899);
xnor U33523 (N_33523,N_22521,N_24736);
nand U33524 (N_33524,N_23297,N_22172);
xor U33525 (N_33525,N_24839,N_25775);
and U33526 (N_33526,N_24566,N_29667);
nor U33527 (N_33527,N_23832,N_20951);
nand U33528 (N_33528,N_27275,N_26319);
or U33529 (N_33529,N_28767,N_21833);
and U33530 (N_33530,N_29234,N_28405);
and U33531 (N_33531,N_28958,N_21354);
nor U33532 (N_33532,N_23226,N_21186);
or U33533 (N_33533,N_24931,N_21769);
and U33534 (N_33534,N_20693,N_20399);
nor U33535 (N_33535,N_20250,N_27196);
or U33536 (N_33536,N_28972,N_29330);
nand U33537 (N_33537,N_29895,N_23670);
or U33538 (N_33538,N_20505,N_25102);
nor U33539 (N_33539,N_27133,N_24833);
nor U33540 (N_33540,N_22142,N_29223);
nor U33541 (N_33541,N_26158,N_24015);
and U33542 (N_33542,N_26938,N_21914);
and U33543 (N_33543,N_23359,N_26197);
and U33544 (N_33544,N_26905,N_26365);
nand U33545 (N_33545,N_25553,N_23383);
nor U33546 (N_33546,N_25998,N_24401);
nand U33547 (N_33547,N_23981,N_23353);
nor U33548 (N_33548,N_25537,N_22606);
and U33549 (N_33549,N_27581,N_28330);
xnor U33550 (N_33550,N_27464,N_29992);
nand U33551 (N_33551,N_21356,N_28640);
nand U33552 (N_33552,N_22796,N_24499);
and U33553 (N_33553,N_27240,N_21110);
and U33554 (N_33554,N_28749,N_26812);
nor U33555 (N_33555,N_23196,N_25267);
nor U33556 (N_33556,N_21929,N_28317);
and U33557 (N_33557,N_25560,N_29185);
or U33558 (N_33558,N_23345,N_24848);
xor U33559 (N_33559,N_22384,N_23891);
nand U33560 (N_33560,N_26059,N_23787);
nor U33561 (N_33561,N_27280,N_24929);
or U33562 (N_33562,N_25849,N_29221);
nor U33563 (N_33563,N_22655,N_27685);
or U33564 (N_33564,N_21548,N_26619);
nor U33565 (N_33565,N_21253,N_23442);
and U33566 (N_33566,N_24050,N_27913);
nor U33567 (N_33567,N_25323,N_24326);
and U33568 (N_33568,N_27675,N_25166);
or U33569 (N_33569,N_21079,N_28108);
nand U33570 (N_33570,N_28776,N_28387);
and U33571 (N_33571,N_28097,N_29755);
or U33572 (N_33572,N_26517,N_24863);
nand U33573 (N_33573,N_22442,N_25878);
nand U33574 (N_33574,N_24548,N_24030);
or U33575 (N_33575,N_25097,N_21192);
nor U33576 (N_33576,N_24065,N_20331);
or U33577 (N_33577,N_29952,N_29779);
and U33578 (N_33578,N_21597,N_29840);
nor U33579 (N_33579,N_23539,N_23734);
nor U33580 (N_33580,N_24307,N_24328);
nor U33581 (N_33581,N_21196,N_24496);
nand U33582 (N_33582,N_22405,N_23556);
nand U33583 (N_33583,N_24583,N_22519);
or U33584 (N_33584,N_23781,N_25221);
and U33585 (N_33585,N_21716,N_21824);
nor U33586 (N_33586,N_22371,N_27485);
xor U33587 (N_33587,N_21721,N_20582);
nand U33588 (N_33588,N_21420,N_24087);
and U33589 (N_33589,N_29375,N_29110);
nor U33590 (N_33590,N_20494,N_28064);
and U33591 (N_33591,N_22250,N_21830);
nand U33592 (N_33592,N_20476,N_28589);
xor U33593 (N_33593,N_29123,N_21228);
xnor U33594 (N_33594,N_28283,N_28024);
nand U33595 (N_33595,N_23483,N_23764);
or U33596 (N_33596,N_27302,N_29593);
nand U33597 (N_33597,N_23011,N_28812);
nand U33598 (N_33598,N_26412,N_24201);
and U33599 (N_33599,N_23869,N_22738);
or U33600 (N_33600,N_25857,N_28787);
nand U33601 (N_33601,N_23147,N_23985);
nor U33602 (N_33602,N_24819,N_23684);
and U33603 (N_33603,N_24787,N_25057);
and U33604 (N_33604,N_21048,N_29227);
nor U33605 (N_33605,N_23901,N_28568);
or U33606 (N_33606,N_26642,N_24799);
or U33607 (N_33607,N_25746,N_20347);
and U33608 (N_33608,N_28228,N_24923);
xor U33609 (N_33609,N_22802,N_21230);
nor U33610 (N_33610,N_28020,N_21032);
and U33611 (N_33611,N_21433,N_20680);
nand U33612 (N_33612,N_22890,N_21646);
xor U33613 (N_33613,N_22693,N_22749);
or U33614 (N_33614,N_29134,N_26166);
or U33615 (N_33615,N_23946,N_23056);
or U33616 (N_33616,N_27948,N_29944);
nand U33617 (N_33617,N_22921,N_20040);
nand U33618 (N_33618,N_27466,N_21886);
xor U33619 (N_33619,N_27634,N_22664);
nand U33620 (N_33620,N_23838,N_24265);
nand U33621 (N_33621,N_29671,N_29050);
xnor U33622 (N_33622,N_27423,N_26327);
or U33623 (N_33623,N_28398,N_21666);
nor U33624 (N_33624,N_23065,N_29536);
nand U33625 (N_33625,N_23094,N_25138);
nand U33626 (N_33626,N_27071,N_27942);
and U33627 (N_33627,N_29569,N_25542);
and U33628 (N_33628,N_26229,N_20849);
or U33629 (N_33629,N_20305,N_29489);
nand U33630 (N_33630,N_28095,N_27597);
nor U33631 (N_33631,N_29913,N_21564);
xor U33632 (N_33632,N_29340,N_28737);
nand U33633 (N_33633,N_22354,N_26389);
and U33634 (N_33634,N_22152,N_29124);
and U33635 (N_33635,N_27151,N_20037);
nand U33636 (N_33636,N_20798,N_26900);
and U33637 (N_33637,N_21998,N_28096);
and U33638 (N_33638,N_21309,N_26144);
nor U33639 (N_33639,N_22874,N_28189);
nor U33640 (N_33640,N_29529,N_20509);
nor U33641 (N_33641,N_23053,N_26243);
and U33642 (N_33642,N_25186,N_29298);
and U33643 (N_33643,N_21922,N_28675);
xor U33644 (N_33644,N_25208,N_25340);
nor U33645 (N_33645,N_20714,N_23350);
nand U33646 (N_33646,N_29015,N_22438);
and U33647 (N_33647,N_23582,N_23255);
or U33648 (N_33648,N_25511,N_24159);
and U33649 (N_33649,N_26482,N_28278);
nand U33650 (N_33650,N_24093,N_25515);
or U33651 (N_33651,N_22569,N_23806);
nor U33652 (N_33652,N_27847,N_20575);
or U33653 (N_33653,N_29812,N_26874);
or U33654 (N_33654,N_23870,N_26118);
nor U33655 (N_33655,N_23312,N_22189);
and U33656 (N_33656,N_24879,N_22788);
nor U33657 (N_33657,N_26597,N_22581);
or U33658 (N_33658,N_26173,N_26191);
or U33659 (N_33659,N_25516,N_28535);
or U33660 (N_33660,N_28810,N_27711);
nor U33661 (N_33661,N_24281,N_28865);
xor U33662 (N_33662,N_28723,N_25747);
or U33663 (N_33663,N_24367,N_21045);
or U33664 (N_33664,N_25470,N_22629);
nand U33665 (N_33665,N_23172,N_22579);
and U33666 (N_33666,N_27918,N_25161);
and U33667 (N_33667,N_23599,N_22505);
and U33668 (N_33668,N_21507,N_20868);
xnor U33669 (N_33669,N_23002,N_25966);
nor U33670 (N_33670,N_27586,N_23323);
nor U33671 (N_33671,N_22292,N_24157);
xnor U33672 (N_33672,N_22037,N_22808);
and U33673 (N_33673,N_20174,N_27938);
nor U33674 (N_33674,N_27629,N_27406);
or U33675 (N_33675,N_25425,N_23583);
xnor U33676 (N_33676,N_29911,N_27046);
nand U33677 (N_33677,N_22906,N_26228);
nor U33678 (N_33678,N_21927,N_23097);
and U33679 (N_33679,N_28134,N_20046);
or U33680 (N_33680,N_23841,N_22803);
xnor U33681 (N_33681,N_20056,N_24828);
nand U33682 (N_33682,N_29106,N_23480);
nor U33683 (N_33683,N_26400,N_24225);
or U33684 (N_33684,N_20055,N_21814);
and U33685 (N_33685,N_21054,N_25045);
xor U33686 (N_33686,N_22518,N_21373);
nor U33687 (N_33687,N_20350,N_24985);
or U33688 (N_33688,N_29753,N_21337);
and U33689 (N_33689,N_27167,N_27883);
or U33690 (N_33690,N_21166,N_28323);
nand U33691 (N_33691,N_28613,N_23991);
nor U33692 (N_33692,N_25235,N_23552);
and U33693 (N_33693,N_20389,N_27461);
nand U33694 (N_33694,N_24616,N_24272);
and U33695 (N_33695,N_28256,N_24911);
nor U33696 (N_33696,N_25664,N_29568);
xor U33697 (N_33697,N_25085,N_27814);
nand U33698 (N_33698,N_27561,N_21088);
nor U33699 (N_33699,N_25871,N_21518);
xnor U33700 (N_33700,N_29318,N_27432);
or U33701 (N_33701,N_26043,N_23067);
or U33702 (N_33702,N_26321,N_26729);
xnor U33703 (N_33703,N_23868,N_26397);
xnor U33704 (N_33704,N_27407,N_27972);
and U33705 (N_33705,N_23990,N_22877);
and U33706 (N_33706,N_29982,N_26746);
nor U33707 (N_33707,N_29007,N_28133);
nand U33708 (N_33708,N_26459,N_28316);
nand U33709 (N_33709,N_24979,N_22913);
nor U33710 (N_33710,N_29459,N_25808);
nand U33711 (N_33711,N_25502,N_20042);
or U33712 (N_33712,N_28922,N_26557);
nand U33713 (N_33713,N_22699,N_21995);
nor U33714 (N_33714,N_25240,N_25341);
nand U33715 (N_33715,N_29594,N_22634);
nand U33716 (N_33716,N_25056,N_21892);
nand U33717 (N_33717,N_20340,N_20467);
or U33718 (N_33718,N_29948,N_28598);
or U33719 (N_33719,N_29823,N_20920);
nor U33720 (N_33720,N_27368,N_23462);
nor U33721 (N_33721,N_21821,N_21488);
or U33722 (N_33722,N_20924,N_22224);
or U33723 (N_33723,N_27279,N_27014);
nor U33724 (N_33724,N_29862,N_25054);
or U33725 (N_33725,N_29508,N_23308);
nor U33726 (N_33726,N_23722,N_24260);
or U33727 (N_33727,N_27409,N_27717);
and U33728 (N_33728,N_28002,N_29092);
nor U33729 (N_33729,N_20095,N_23326);
or U33730 (N_33730,N_28347,N_27362);
and U33731 (N_33731,N_23674,N_28181);
nand U33732 (N_33732,N_28105,N_28127);
or U33733 (N_33733,N_23355,N_23456);
xor U33734 (N_33734,N_20111,N_24449);
nor U33735 (N_33735,N_22541,N_20939);
and U33736 (N_33736,N_29139,N_20987);
or U33737 (N_33737,N_26907,N_28410);
nand U33738 (N_33738,N_21938,N_29105);
xor U33739 (N_33739,N_28211,N_29465);
and U33740 (N_33740,N_25779,N_20472);
nor U33741 (N_33741,N_25306,N_26437);
and U33742 (N_33742,N_24915,N_28333);
and U33743 (N_33743,N_26840,N_28334);
and U33744 (N_33744,N_29327,N_25940);
and U33745 (N_33745,N_25471,N_22336);
nand U33746 (N_33746,N_27835,N_27162);
nand U33747 (N_33747,N_27306,N_29485);
nand U33748 (N_33748,N_28831,N_28704);
or U33749 (N_33749,N_22688,N_25427);
nand U33750 (N_33750,N_20954,N_29195);
or U33751 (N_33751,N_21805,N_20165);
or U33752 (N_33752,N_25271,N_24511);
and U33753 (N_33753,N_27308,N_25834);
nor U33754 (N_33754,N_28792,N_20203);
xnor U33755 (N_33755,N_23754,N_25083);
or U33756 (N_33756,N_28555,N_21516);
and U33757 (N_33757,N_25354,N_25585);
or U33758 (N_33758,N_23020,N_27392);
nand U33759 (N_33759,N_25885,N_22197);
nor U33760 (N_33760,N_26551,N_23144);
or U33761 (N_33761,N_24102,N_28205);
and U33762 (N_33762,N_24761,N_21570);
nor U33763 (N_33763,N_28199,N_21947);
xor U33764 (N_33764,N_29758,N_24095);
and U33765 (N_33765,N_25334,N_21440);
nand U33766 (N_33766,N_22568,N_21387);
and U33767 (N_33767,N_20451,N_28557);
xor U33768 (N_33768,N_21699,N_21338);
and U33769 (N_33769,N_27192,N_29828);
xnor U33770 (N_33770,N_24180,N_20016);
nor U33771 (N_33771,N_24304,N_20270);
nor U33772 (N_33772,N_25361,N_24838);
or U33773 (N_33773,N_22173,N_22462);
nor U33774 (N_33774,N_24283,N_29499);
or U33775 (N_33775,N_22001,N_23548);
and U33776 (N_33776,N_29082,N_29616);
nand U33777 (N_33777,N_23914,N_28636);
nor U33778 (N_33778,N_20889,N_26317);
and U33779 (N_33779,N_24327,N_25532);
xor U33780 (N_33780,N_29750,N_24779);
or U33781 (N_33781,N_29281,N_29826);
nand U33782 (N_33782,N_23475,N_27395);
nor U33783 (N_33783,N_26011,N_23276);
xor U33784 (N_33784,N_22814,N_24716);
nor U33785 (N_33785,N_24273,N_29456);
nand U33786 (N_33786,N_20704,N_23417);
xor U33787 (N_33787,N_28507,N_21677);
or U33788 (N_33788,N_21773,N_29925);
and U33789 (N_33789,N_27920,N_21100);
or U33790 (N_33790,N_23895,N_29797);
nand U33791 (N_33791,N_24591,N_25082);
and U33792 (N_33792,N_23699,N_25901);
and U33793 (N_33793,N_23309,N_28619);
nor U33794 (N_33794,N_22771,N_21127);
or U33795 (N_33795,N_25184,N_28031);
nand U33796 (N_33796,N_21289,N_21176);
and U33797 (N_33797,N_26203,N_20176);
nand U33798 (N_33798,N_26659,N_27286);
nand U33799 (N_33799,N_21182,N_25367);
and U33800 (N_33800,N_25292,N_24752);
nand U33801 (N_33801,N_27495,N_27007);
nand U33802 (N_33802,N_24149,N_24847);
and U33803 (N_33803,N_20164,N_23621);
and U33804 (N_33804,N_21680,N_28975);
nor U33805 (N_33805,N_24135,N_20919);
or U33806 (N_33806,N_20830,N_28860);
or U33807 (N_33807,N_28243,N_27955);
nand U33808 (N_33808,N_21402,N_28685);
or U33809 (N_33809,N_27537,N_26289);
nand U33810 (N_33810,N_22295,N_20248);
nand U33811 (N_33811,N_24295,N_23243);
nor U33812 (N_33812,N_26215,N_22432);
nor U33813 (N_33813,N_27846,N_27173);
or U33814 (N_33814,N_29474,N_22176);
nor U33815 (N_33815,N_21411,N_25633);
nor U33816 (N_33816,N_21979,N_26204);
nand U33817 (N_33817,N_23954,N_29570);
xor U33818 (N_33818,N_20281,N_21743);
nand U33819 (N_33819,N_22501,N_28194);
nand U33820 (N_33820,N_27070,N_21586);
and U33821 (N_33821,N_24725,N_20021);
nor U33822 (N_33822,N_22709,N_20972);
nand U33823 (N_33823,N_26994,N_23802);
nor U33824 (N_33824,N_28276,N_21669);
and U33825 (N_33825,N_23470,N_27815);
nor U33826 (N_33826,N_23184,N_24404);
nor U33827 (N_33827,N_26876,N_22454);
xnor U33828 (N_33828,N_28186,N_29111);
nand U33829 (N_33829,N_22754,N_24424);
and U33830 (N_33830,N_28408,N_26065);
or U33831 (N_33831,N_25549,N_27650);
nand U33832 (N_33832,N_21062,N_27916);
or U33833 (N_33833,N_20755,N_25095);
or U33834 (N_33834,N_25562,N_27760);
nor U33835 (N_33835,N_28202,N_23942);
or U33836 (N_33836,N_25454,N_23341);
nand U33837 (N_33837,N_20862,N_22844);
nand U33838 (N_33838,N_29525,N_21789);
nor U33839 (N_33839,N_20402,N_25858);
and U33840 (N_33840,N_27845,N_23010);
nand U33841 (N_33841,N_21798,N_29951);
and U33842 (N_33842,N_25623,N_28744);
nor U33843 (N_33843,N_22739,N_22886);
nand U33844 (N_33844,N_26342,N_23727);
or U33845 (N_33845,N_27818,N_27636);
nand U33846 (N_33846,N_20265,N_21685);
or U33847 (N_33847,N_23429,N_26443);
nor U33848 (N_33848,N_23508,N_27674);
or U33849 (N_33849,N_29978,N_24643);
nand U33850 (N_33850,N_24211,N_24447);
or U33851 (N_33851,N_26873,N_27576);
nor U33852 (N_33852,N_24980,N_22799);
and U33853 (N_33853,N_22276,N_26916);
or U33854 (N_33854,N_23169,N_26810);
and U33855 (N_33855,N_29042,N_22600);
and U33856 (N_33856,N_26315,N_28571);
nor U33857 (N_33857,N_25131,N_21840);
and U33858 (N_33858,N_22491,N_27907);
xnor U33859 (N_33859,N_27857,N_27193);
nor U33860 (N_33860,N_21256,N_20009);
or U33861 (N_33861,N_27585,N_26625);
nand U33862 (N_33862,N_26849,N_29498);
xor U33863 (N_33863,N_29776,N_27735);
nor U33864 (N_33864,N_27853,N_28294);
nand U33865 (N_33865,N_28295,N_29020);
nand U33866 (N_33866,N_21122,N_21584);
and U33867 (N_33867,N_26790,N_26060);
or U33868 (N_33868,N_22437,N_27930);
or U33869 (N_33869,N_24188,N_21623);
and U33870 (N_33870,N_24626,N_24471);
or U33871 (N_33871,N_28233,N_29366);
nand U33872 (N_33872,N_29685,N_28272);
and U33873 (N_33873,N_28434,N_25543);
nor U33874 (N_33874,N_26098,N_22398);
nor U33875 (N_33875,N_25243,N_24039);
nand U33876 (N_33876,N_25149,N_28341);
nand U33877 (N_33877,N_23098,N_23482);
nand U33878 (N_33878,N_21418,N_22399);
or U33879 (N_33879,N_27376,N_25742);
nor U33880 (N_33880,N_22426,N_29962);
or U33881 (N_33881,N_25629,N_23534);
nor U33882 (N_33882,N_29564,N_22968);
nor U33883 (N_33883,N_28019,N_20948);
nor U33884 (N_33884,N_28546,N_23099);
or U33885 (N_33885,N_27017,N_28299);
nor U33886 (N_33886,N_24152,N_29834);
and U33887 (N_33887,N_21360,N_21912);
xnor U33888 (N_33888,N_23398,N_20155);
nor U33889 (N_33889,N_25232,N_21662);
or U33890 (N_33890,N_22563,N_22792);
nor U33891 (N_33891,N_27543,N_29477);
nor U33892 (N_33892,N_25576,N_27176);
and U33893 (N_33893,N_24174,N_21239);
nor U33894 (N_33894,N_20612,N_21332);
nand U33895 (N_33895,N_28358,N_27780);
xnor U33896 (N_33896,N_26278,N_29197);
xor U33897 (N_33897,N_22533,N_27737);
and U33898 (N_33898,N_24353,N_20746);
or U33899 (N_33899,N_29829,N_21741);
xor U33900 (N_33900,N_20542,N_20683);
nand U33901 (N_33901,N_20531,N_22758);
and U33902 (N_33902,N_27397,N_22622);
nand U33903 (N_33903,N_25666,N_28164);
nor U33904 (N_33904,N_29414,N_26807);
and U33905 (N_33905,N_20856,N_22139);
xor U33906 (N_33906,N_29012,N_25672);
or U33907 (N_33907,N_23777,N_20601);
and U33908 (N_33908,N_28655,N_22904);
nand U33909 (N_33909,N_22846,N_26645);
nor U33910 (N_33910,N_22894,N_23726);
nand U33911 (N_33911,N_27237,N_27438);
xnor U33912 (N_33912,N_23890,N_25505);
nor U33913 (N_33913,N_27088,N_25216);
nand U33914 (N_33914,N_22357,N_26078);
nand U33915 (N_33915,N_25520,N_23652);
and U33916 (N_33916,N_25893,N_20813);
nand U33917 (N_33917,N_21534,N_23029);
nor U33918 (N_33918,N_22614,N_25072);
nand U33919 (N_33919,N_29848,N_21271);
and U33920 (N_33920,N_27505,N_20622);
and U33921 (N_33921,N_25413,N_28487);
nor U33922 (N_33922,N_26965,N_21319);
and U33923 (N_33923,N_24373,N_21844);
or U33924 (N_33924,N_27781,N_20949);
and U33925 (N_33925,N_21334,N_20349);
and U33926 (N_33926,N_25837,N_21498);
and U33927 (N_33927,N_29697,N_25178);
nand U33928 (N_33928,N_23405,N_24827);
and U33929 (N_33929,N_24928,N_25337);
nor U33930 (N_33930,N_29096,N_28107);
nand U33931 (N_33931,N_23755,N_26732);
nor U33932 (N_33932,N_25468,N_24547);
nand U33933 (N_33933,N_27753,N_23893);
nand U33934 (N_33934,N_23917,N_24294);
nand U33935 (N_33935,N_25734,N_27575);
nand U33936 (N_33936,N_28223,N_28417);
nor U33937 (N_33937,N_28169,N_24136);
nor U33938 (N_33938,N_26458,N_24914);
or U33939 (N_33939,N_27821,N_20325);
or U33940 (N_33940,N_23181,N_22948);
nand U33941 (N_33941,N_22602,N_26130);
xor U33942 (N_33942,N_20584,N_29484);
nor U33943 (N_33943,N_29081,N_21860);
xor U33944 (N_33944,N_20589,N_28422);
nand U33945 (N_33945,N_29724,N_21801);
or U33946 (N_33946,N_20074,N_28917);
nor U33947 (N_33947,N_21046,N_22902);
or U33948 (N_33948,N_29062,N_26618);
and U33949 (N_33949,N_27497,N_20137);
nor U33950 (N_33950,N_25415,N_21376);
nand U33951 (N_33951,N_21718,N_26621);
nand U33952 (N_33952,N_21467,N_20973);
xnor U33953 (N_33953,N_23316,N_21696);
and U33954 (N_33954,N_26001,N_20196);
nand U33955 (N_33955,N_29935,N_26599);
xnor U33956 (N_33956,N_25701,N_28472);
nand U33957 (N_33957,N_22930,N_22863);
nor U33958 (N_33958,N_28526,N_27796);
nand U33959 (N_33959,N_22817,N_24110);
nor U33960 (N_33960,N_21224,N_26129);
nor U33961 (N_33961,N_22095,N_27375);
and U33962 (N_33962,N_23817,N_26827);
or U33963 (N_33963,N_28821,N_29729);
nand U33964 (N_33964,N_27660,N_27334);
nand U33965 (N_33965,N_29659,N_21077);
nor U33966 (N_33966,N_22715,N_28641);
nor U33967 (N_33967,N_21486,N_25040);
nand U33968 (N_33968,N_21511,N_28093);
and U33969 (N_33969,N_28141,N_27112);
xnor U33970 (N_33970,N_27819,N_26946);
or U33971 (N_33971,N_25251,N_20133);
nor U33972 (N_33972,N_29045,N_24644);
and U33973 (N_33973,N_27639,N_23073);
nor U33974 (N_33974,N_22720,N_23060);
and U33975 (N_33975,N_25167,N_24001);
or U33976 (N_33976,N_23506,N_25642);
and U33977 (N_33977,N_27580,N_22119);
nor U33978 (N_33978,N_23189,N_28142);
nand U33979 (N_33979,N_28292,N_24918);
xor U33980 (N_33980,N_29547,N_29217);
nand U33981 (N_33981,N_24641,N_25113);
or U33982 (N_33982,N_27241,N_28694);
and U33983 (N_33983,N_22088,N_25976);
xor U33984 (N_33984,N_22565,N_24132);
nor U33985 (N_33985,N_21296,N_22372);
nor U33986 (N_33986,N_21142,N_29353);
nand U33987 (N_33987,N_29811,N_25991);
nand U33988 (N_33988,N_23809,N_24685);
or U33989 (N_33989,N_25092,N_21608);
or U33990 (N_33990,N_23798,N_20767);
nor U33991 (N_33991,N_21827,N_28039);
nor U33992 (N_33992,N_23610,N_20006);
or U33993 (N_33993,N_21648,N_27453);
and U33994 (N_33994,N_28302,N_27187);
nand U33995 (N_33995,N_24531,N_24309);
and U33996 (N_33996,N_22470,N_28805);
or U33997 (N_33997,N_26639,N_21550);
and U33998 (N_33998,N_22884,N_24570);
or U33999 (N_33999,N_20833,N_23325);
nor U34000 (N_34000,N_29164,N_22941);
nor U34001 (N_34001,N_25996,N_22129);
nor U34002 (N_34002,N_23602,N_28657);
or U34003 (N_34003,N_25282,N_20097);
nand U34004 (N_34004,N_23979,N_25964);
xnor U34005 (N_34005,N_22333,N_27148);
and U34006 (N_34006,N_27603,N_21799);
and U34007 (N_34007,N_26336,N_27082);
and U34008 (N_34008,N_25254,N_20558);
and U34009 (N_34009,N_22961,N_28445);
or U34010 (N_34010,N_28715,N_21545);
nand U34011 (N_34011,N_28482,N_27462);
and U34012 (N_34012,N_23499,N_27884);
nor U34013 (N_34013,N_23541,N_23597);
nand U34014 (N_34014,N_20611,N_21640);
or U34015 (N_34015,N_21293,N_28152);
or U34016 (N_34016,N_20775,N_25408);
and U34017 (N_34017,N_27732,N_29871);
nor U34018 (N_34018,N_26792,N_23414);
nand U34019 (N_34019,N_23653,N_25887);
nand U34020 (N_34020,N_23521,N_24900);
nand U34021 (N_34021,N_21302,N_27544);
and U34022 (N_34022,N_28532,N_22236);
xor U34023 (N_34023,N_20976,N_22267);
nand U34024 (N_34024,N_21695,N_27269);
nand U34025 (N_34025,N_29351,N_23958);
nand U34026 (N_34026,N_20803,N_20892);
nor U34027 (N_34027,N_26614,N_24143);
and U34028 (N_34028,N_23028,N_25005);
nand U34029 (N_34029,N_23790,N_24732);
nand U34030 (N_34030,N_29297,N_24962);
nor U34031 (N_34031,N_21207,N_23519);
xnor U34032 (N_34032,N_28219,N_27186);
nor U34033 (N_34033,N_29558,N_26852);
and U34034 (N_34034,N_22972,N_29715);
and U34035 (N_34035,N_26449,N_24927);
and U34036 (N_34036,N_29258,N_24356);
nor U34037 (N_34037,N_23179,N_22845);
nor U34038 (N_34038,N_26076,N_24371);
nand U34039 (N_34039,N_25476,N_25244);
nor U34040 (N_34040,N_26263,N_23401);
nor U34041 (N_34041,N_28849,N_23719);
xor U34042 (N_34042,N_20586,N_21701);
xor U34043 (N_34043,N_25552,N_20516);
nand U34044 (N_34044,N_24350,N_27905);
nor U34045 (N_34045,N_27218,N_21603);
nand U34046 (N_34046,N_28659,N_20721);
xnor U34047 (N_34047,N_26303,N_24389);
nand U34048 (N_34048,N_25137,N_28938);
nand U34049 (N_34049,N_27032,N_22108);
nor U34050 (N_34050,N_20674,N_21977);
or U34051 (N_34051,N_24361,N_22363);
nand U34052 (N_34052,N_29002,N_21180);
and U34053 (N_34053,N_20288,N_22811);
nand U34054 (N_34054,N_21903,N_28383);
and U34055 (N_34055,N_29455,N_27903);
nand U34056 (N_34056,N_22464,N_26539);
nor U34057 (N_34057,N_25853,N_25132);
or U34058 (N_34058,N_21390,N_24604);
nor U34059 (N_34059,N_24588,N_23409);
nand U34060 (N_34060,N_23396,N_26888);
or U34061 (N_34061,N_27338,N_28245);
nor U34062 (N_34062,N_29809,N_24255);
xor U34063 (N_34063,N_25025,N_23691);
xnor U34064 (N_34064,N_23377,N_26841);
nor U34065 (N_34065,N_28998,N_26847);
nor U34066 (N_34066,N_27914,N_29182);
nand U34067 (N_34067,N_26715,N_21016);
nor U34068 (N_34068,N_27131,N_28839);
or U34069 (N_34069,N_26627,N_26641);
and U34070 (N_34070,N_27951,N_21453);
nand U34071 (N_34071,N_23823,N_20048);
xnor U34072 (N_34072,N_25656,N_28757);
and U34073 (N_34073,N_26828,N_26376);
or U34074 (N_34074,N_21654,N_26042);
or U34075 (N_34075,N_24319,N_20035);
nor U34076 (N_34076,N_26378,N_28707);
nand U34077 (N_34077,N_26885,N_22339);
nor U34078 (N_34078,N_20354,N_23911);
xor U34079 (N_34079,N_25237,N_21083);
or U34080 (N_34080,N_23522,N_24892);
and U34081 (N_34081,N_20965,N_20905);
nand U34082 (N_34082,N_29535,N_22297);
xor U34083 (N_34083,N_25621,N_26105);
and U34084 (N_34084,N_23362,N_24747);
nor U34085 (N_34085,N_28699,N_20595);
nor U34086 (N_34086,N_29875,N_28769);
nor U34087 (N_34087,N_21868,N_26784);
nand U34088 (N_34088,N_23678,N_20499);
or U34089 (N_34089,N_24709,N_24100);
or U34090 (N_34090,N_21790,N_24870);
nand U34091 (N_34091,N_23458,N_20635);
and U34092 (N_34092,N_23472,N_27706);
nand U34093 (N_34093,N_29175,N_25345);
or U34094 (N_34094,N_29794,N_22424);
nor U34095 (N_34095,N_25669,N_28214);
or U34096 (N_34096,N_29921,N_27960);
nand U34097 (N_34097,N_21251,N_20244);
or U34098 (N_34098,N_25365,N_29872);
and U34099 (N_34099,N_22386,N_27390);
or U34100 (N_34100,N_29179,N_28864);
or U34101 (N_34101,N_25075,N_23545);
or U34102 (N_34102,N_20114,N_29280);
or U34103 (N_34103,N_26460,N_20328);
xnor U34104 (N_34104,N_20925,N_26603);
nor U34105 (N_34105,N_26724,N_28902);
nand U34106 (N_34106,N_20064,N_24384);
and U34107 (N_34107,N_28478,N_20668);
xnor U34108 (N_34108,N_20995,N_23074);
nand U34109 (N_34109,N_24193,N_21200);
or U34110 (N_34110,N_20910,N_25359);
nand U34111 (N_34111,N_27562,N_29761);
and U34112 (N_34112,N_26025,N_27109);
or U34113 (N_34113,N_23231,N_24429);
and U34114 (N_34114,N_26356,N_22748);
and U34115 (N_34115,N_23368,N_25667);
and U34116 (N_34116,N_20921,N_24165);
or U34117 (N_34117,N_20545,N_20029);
nor U34118 (N_34118,N_29652,N_20896);
nand U34119 (N_34119,N_28607,N_20432);
and U34120 (N_34120,N_29093,N_28806);
nand U34121 (N_34121,N_29902,N_23725);
nor U34122 (N_34122,N_23526,N_22252);
and U34123 (N_34123,N_25513,N_20570);
xor U34124 (N_34124,N_22815,N_21396);
and U34125 (N_34125,N_20141,N_28023);
and U34126 (N_34126,N_24245,N_24654);
nor U34127 (N_34127,N_28457,N_25016);
and U34128 (N_34128,N_29744,N_26337);
xnor U34129 (N_34129,N_28501,N_28087);
nor U34130 (N_34130,N_26344,N_24325);
and U34131 (N_34131,N_24341,N_22323);
or U34132 (N_34132,N_24947,N_22263);
nand U34133 (N_34133,N_23929,N_25605);
or U34134 (N_34134,N_21288,N_24506);
xor U34135 (N_34135,N_26192,N_24745);
nor U34136 (N_34136,N_23116,N_28173);
nor U34137 (N_34137,N_21620,N_24301);
or U34138 (N_34138,N_23740,N_27987);
and U34139 (N_34139,N_27134,N_20268);
or U34140 (N_34140,N_24864,N_24941);
or U34141 (N_34141,N_21451,N_25127);
and U34142 (N_34142,N_24638,N_20640);
and U34143 (N_34143,N_27949,N_21044);
nand U34144 (N_34144,N_21930,N_22146);
or U34145 (N_34145,N_22932,N_22513);
nand U34146 (N_34146,N_26217,N_20824);
nand U34147 (N_34147,N_20898,N_29388);
nand U34148 (N_34148,N_23221,N_28697);
or U34149 (N_34149,N_23303,N_20847);
or U34150 (N_34150,N_29422,N_27416);
xor U34151 (N_34151,N_29080,N_23608);
nor U34152 (N_34152,N_20713,N_29587);
or U34153 (N_34153,N_27037,N_29793);
nor U34154 (N_34154,N_22990,N_25423);
and U34155 (N_34155,N_28531,N_28140);
nand U34156 (N_34156,N_21641,N_23977);
nor U34157 (N_34157,N_26314,N_29543);
nand U34158 (N_34158,N_22989,N_20105);
or U34159 (N_34159,N_23634,N_22652);
or U34160 (N_34160,N_20089,N_28029);
and U34161 (N_34161,N_27211,N_23933);
or U34162 (N_34162,N_27364,N_24846);
nor U34163 (N_34163,N_26779,N_23177);
xor U34164 (N_34164,N_20734,N_22860);
or U34165 (N_34165,N_25728,N_20480);
nand U34166 (N_34166,N_23239,N_23331);
and U34167 (N_34167,N_21459,N_25508);
nor U34168 (N_34168,N_22359,N_27493);
nor U34169 (N_34169,N_23406,N_26379);
and U34170 (N_34170,N_22429,N_22210);
nor U34171 (N_34171,N_24123,N_27318);
or U34172 (N_34172,N_21658,N_23300);
and U34173 (N_34173,N_29409,N_26646);
nand U34174 (N_34174,N_26194,N_26297);
nor U34175 (N_34175,N_21347,N_27201);
nand U34176 (N_34176,N_20185,N_29650);
nand U34177 (N_34177,N_29888,N_25783);
or U34178 (N_34178,N_23329,N_27538);
and U34179 (N_34179,N_27089,N_29905);
xnor U34180 (N_34180,N_29288,N_28209);
nor U34181 (N_34181,N_29038,N_23892);
xnor U34182 (N_34182,N_22658,N_20099);
nor U34183 (N_34183,N_24121,N_20127);
xor U34184 (N_34184,N_26769,N_22115);
or U34185 (N_34185,N_21510,N_28042);
nor U34186 (N_34186,N_22193,N_22615);
nor U34187 (N_34187,N_20700,N_20260);
and U34188 (N_34188,N_26236,N_26751);
or U34189 (N_34189,N_23346,N_27246);
nor U34190 (N_34190,N_23087,N_24284);
nor U34191 (N_34191,N_22487,N_25158);
nand U34192 (N_34192,N_22287,N_20715);
or U34193 (N_34193,N_29200,N_22607);
and U34194 (N_34194,N_22171,N_23812);
nor U34195 (N_34195,N_23647,N_23319);
and U34196 (N_34196,N_22213,N_23635);
or U34197 (N_34197,N_29555,N_22490);
nor U34198 (N_34198,N_22180,N_21491);
xor U34199 (N_34199,N_22924,N_25671);
or U34200 (N_34200,N_29827,N_21689);
nor U34201 (N_34201,N_26131,N_29618);
and U34202 (N_34202,N_28985,N_24256);
and U34203 (N_34203,N_22526,N_25407);
and U34204 (N_34204,N_20214,N_25503);
or U34205 (N_34205,N_27806,N_21972);
and U34206 (N_34206,N_21027,N_21719);
or U34207 (N_34207,N_21461,N_20377);
and U34208 (N_34208,N_26193,N_22107);
or U34209 (N_34209,N_21452,N_29787);
nor U34210 (N_34210,N_28528,N_20227);
nand U34211 (N_34211,N_23923,N_28444);
and U34212 (N_34212,N_21317,N_26031);
or U34213 (N_34213,N_28706,N_21422);
and U34214 (N_34214,N_26135,N_29832);
nand U34215 (N_34215,N_22041,N_29168);
or U34216 (N_34216,N_28947,N_22319);
nand U34217 (N_34217,N_28040,N_20221);
nand U34218 (N_34218,N_21878,N_22960);
or U34219 (N_34219,N_25548,N_29178);
nor U34220 (N_34220,N_27428,N_23604);
or U34221 (N_34221,N_25173,N_29662);
or U34222 (N_34222,N_25327,N_21162);
or U34223 (N_34223,N_25214,N_29188);
xor U34224 (N_34224,N_24111,N_29198);
and U34225 (N_34225,N_25693,N_25611);
nor U34226 (N_34226,N_29859,N_23578);
nand U34227 (N_34227,N_28327,N_21885);
or U34228 (N_34228,N_21071,N_24321);
nand U34229 (N_34229,N_29174,N_23968);
and U34230 (N_34230,N_21261,N_24216);
nor U34231 (N_34231,N_22257,N_21084);
nor U34232 (N_34232,N_22682,N_24406);
nand U34233 (N_34233,N_24612,N_22222);
nand U34234 (N_34234,N_21011,N_25894);
nand U34235 (N_34235,N_27901,N_20917);
nor U34236 (N_34236,N_20854,N_25305);
nand U34237 (N_34237,N_21052,N_24472);
or U34238 (N_34238,N_24101,N_21846);
nor U34239 (N_34239,N_27231,N_25650);
or U34240 (N_34240,N_21153,N_23622);
and U34241 (N_34241,N_26032,N_26743);
or U34242 (N_34242,N_27702,N_24443);
or U34243 (N_34243,N_26188,N_25707);
nand U34244 (N_34244,N_24913,N_25364);
nor U34245 (N_34245,N_21522,N_22805);
nand U34246 (N_34246,N_27501,N_21355);
nor U34247 (N_34247,N_28028,N_29089);
and U34248 (N_34248,N_24543,N_27804);
and U34249 (N_34249,N_20110,N_29997);
nand U34250 (N_34250,N_22494,N_21874);
nor U34251 (N_34251,N_28789,N_24628);
xor U34252 (N_34252,N_20128,N_23191);
or U34253 (N_34253,N_29983,N_26477);
nand U34254 (N_34254,N_29129,N_28036);
nand U34255 (N_34255,N_26498,N_28786);
nand U34256 (N_34256,N_28511,N_21278);
xor U34257 (N_34257,N_27472,N_21989);
nand U34258 (N_34258,N_23955,N_23484);
xor U34259 (N_34259,N_28664,N_20961);
nor U34260 (N_34260,N_20928,N_20446);
and U34261 (N_34261,N_29762,N_28576);
or U34262 (N_34262,N_21098,N_23888);
or U34263 (N_34263,N_23361,N_28124);
nor U34264 (N_34264,N_25933,N_25473);
and U34265 (N_34265,N_23404,N_25440);
nand U34266 (N_34266,N_20685,N_29562);
xnor U34267 (N_34267,N_27214,N_27761);
or U34268 (N_34268,N_21605,N_26016);
and U34269 (N_34269,N_29584,N_26543);
and U34270 (N_34270,N_27456,N_29849);
nand U34271 (N_34271,N_22914,N_22644);
and U34272 (N_34272,N_23713,N_27588);
nand U34273 (N_34273,N_23135,N_24861);
nor U34274 (N_34274,N_28072,N_27797);
nor U34275 (N_34275,N_23295,N_20346);
and U34276 (N_34276,N_23217,N_29140);
nand U34277 (N_34277,N_23399,N_21828);
nor U34278 (N_34278,N_26880,N_25951);
or U34279 (N_34279,N_26250,N_20054);
nor U34280 (N_34280,N_25439,N_21610);
or U34281 (N_34281,N_23228,N_25712);
nor U34282 (N_34282,N_20468,N_23772);
nor U34283 (N_34283,N_27856,N_20386);
nor U34284 (N_34284,N_20158,N_27135);
xnor U34285 (N_34285,N_24667,N_24686);
or U34286 (N_34286,N_24504,N_27258);
nor U34287 (N_34287,N_20371,N_23957);
nor U34288 (N_34288,N_29204,N_21819);
nand U34289 (N_34289,N_26216,N_22595);
or U34290 (N_34290,N_22951,N_29868);
xnor U34291 (N_34291,N_21936,N_28855);
or U34292 (N_34292,N_21625,N_20681);
nand U34293 (N_34293,N_25999,N_29682);
or U34294 (N_34294,N_26332,N_23115);
nand U34295 (N_34295,N_22639,N_27839);
nand U34296 (N_34296,N_23795,N_26184);
xnor U34297 (N_34297,N_29833,N_24968);
nor U34298 (N_34298,N_25724,N_26588);
and U34299 (N_34299,N_22853,N_24609);
or U34300 (N_34300,N_24032,N_26320);
and U34301 (N_34301,N_22637,N_29632);
and U34302 (N_34302,N_22149,N_27123);
nor U34303 (N_34303,N_26903,N_27986);
nand U34304 (N_34304,N_22201,N_24930);
or U34305 (N_34305,N_26569,N_29220);
or U34306 (N_34306,N_27595,N_21694);
and U34307 (N_34307,N_24163,N_22211);
nor U34308 (N_34308,N_23235,N_22552);
nor U34309 (N_34309,N_22823,N_26660);
nor U34310 (N_34310,N_22450,N_21785);
nand U34311 (N_34311,N_28423,N_27008);
or U34312 (N_34312,N_24034,N_24481);
or U34313 (N_34313,N_26152,N_22571);
nor U34314 (N_34314,N_28052,N_22366);
nand U34315 (N_34315,N_26853,N_23501);
nor U34316 (N_34316,N_21463,N_28811);
or U34317 (N_34317,N_26868,N_28018);
nor U34318 (N_34318,N_23091,N_24717);
and U34319 (N_34319,N_27198,N_28962);
nand U34320 (N_34320,N_22245,N_26235);
nand U34321 (N_34321,N_20440,N_29791);
or U34322 (N_34322,N_24354,N_27291);
or U34323 (N_34323,N_27018,N_24250);
and U34324 (N_34324,N_20322,N_29936);
xor U34325 (N_34325,N_27895,N_20358);
and U34326 (N_34326,N_26116,N_21154);
nor U34327 (N_34327,N_20205,N_26821);
nor U34328 (N_34328,N_23165,N_24559);
nor U34329 (N_34329,N_28556,N_23757);
nand U34330 (N_34330,N_28070,N_21369);
or U34331 (N_34331,N_21843,N_28653);
nor U34332 (N_34332,N_21316,N_20484);
and U34333 (N_34333,N_20978,N_21684);
or U34334 (N_34334,N_26839,N_22054);
or U34335 (N_34335,N_21935,N_24118);
nor U34336 (N_34336,N_26370,N_26921);
and U34337 (N_34337,N_24746,N_22931);
nand U34338 (N_34338,N_22104,N_23814);
or U34339 (N_34339,N_26656,N_20539);
and U34340 (N_34340,N_20300,N_23949);
nor U34341 (N_34341,N_20540,N_29265);
or U34342 (N_34342,N_22901,N_25458);
nand U34343 (N_34343,N_23910,N_27044);
nor U34344 (N_34344,N_23594,N_29068);
nand U34345 (N_34345,N_23586,N_28066);
and U34346 (N_34346,N_21856,N_20112);
nand U34347 (N_34347,N_26039,N_26954);
nor U34348 (N_34348,N_24014,N_27304);
xor U34349 (N_34349,N_29738,N_21580);
nand U34350 (N_34350,N_24982,N_28217);
and U34351 (N_34351,N_25170,N_25569);
nor U34352 (N_34352,N_29518,N_26556);
and U34353 (N_34353,N_28822,N_26413);
or U34354 (N_34354,N_25749,N_25389);
or U34355 (N_34355,N_28585,N_24206);
or U34356 (N_34356,N_24883,N_23560);
nand U34357 (N_34357,N_29602,N_22797);
or U34358 (N_34358,N_27171,N_23467);
xnor U34359 (N_34359,N_24624,N_23899);
or U34360 (N_34360,N_29352,N_28601);
xnor U34361 (N_34361,N_25956,N_23477);
or U34362 (N_34362,N_24646,N_23436);
nand U34363 (N_34363,N_20784,N_25032);
or U34364 (N_34364,N_26696,N_25921);
nor U34365 (N_34365,N_27785,N_21193);
nor U34366 (N_34366,N_20081,N_26106);
and U34367 (N_34367,N_22242,N_20673);
nor U34368 (N_34368,N_23365,N_27977);
or U34369 (N_34369,N_20353,N_23618);
and U34370 (N_34370,N_22283,N_28671);
xor U34371 (N_34371,N_20000,N_21568);
nor U34372 (N_34372,N_25499,N_20135);
nor U34373 (N_34373,N_20169,N_28046);
or U34374 (N_34374,N_20474,N_29334);
nand U34375 (N_34375,N_23871,N_28343);
and U34376 (N_34376,N_28995,N_26509);
nor U34377 (N_34377,N_27429,N_23632);
nor U34378 (N_34378,N_22546,N_29934);
and U34379 (N_34379,N_22012,N_21225);
nor U34380 (N_34380,N_25677,N_25333);
or U34381 (N_34381,N_22255,N_21287);
and U34382 (N_34382,N_20782,N_29304);
xor U34383 (N_34383,N_27248,N_23905);
or U34384 (N_34384,N_21583,N_21033);
and U34385 (N_34385,N_29251,N_27740);
nand U34386 (N_34386,N_25441,N_23330);
nand U34387 (N_34387,N_23834,N_29199);
or U34388 (N_34388,N_25162,N_20663);
or U34389 (N_34389,N_21132,N_28734);
nor U34390 (N_34390,N_25563,N_21292);
nor U34391 (N_34391,N_24047,N_20625);
or U34392 (N_34392,N_20343,N_22414);
nand U34393 (N_34393,N_27594,N_20731);
and U34394 (N_34394,N_29488,N_20053);
or U34395 (N_34395,N_26086,N_23479);
and U34396 (N_34396,N_22254,N_23384);
nand U34397 (N_34397,N_29521,N_23951);
and U34398 (N_34398,N_23689,N_25822);
and U34399 (N_34399,N_24817,N_25852);
or U34400 (N_34400,N_28911,N_22134);
nor U34401 (N_34401,N_29137,N_26538);
xnor U34402 (N_34402,N_27830,N_26426);
nor U34403 (N_34403,N_24642,N_24134);
nor U34404 (N_34404,N_22178,N_29506);
nor U34405 (N_34405,N_25109,N_24831);
nor U34406 (N_34406,N_21862,N_24236);
and U34407 (N_34407,N_22978,N_24442);
and U34408 (N_34408,N_22522,N_26843);
xnor U34409 (N_34409,N_21655,N_21458);
xnor U34410 (N_34410,N_25815,N_20733);
nand U34411 (N_34411,N_20060,N_25362);
nand U34412 (N_34412,N_27370,N_23989);
or U34413 (N_34413,N_25546,N_23385);
xor U34414 (N_34414,N_22714,N_20765);
nand U34415 (N_34415,N_21197,N_25101);
nor U34416 (N_34416,N_21925,N_27763);
nor U34417 (N_34417,N_28892,N_29869);
or U34418 (N_34418,N_22585,N_27828);
nand U34419 (N_34419,N_21409,N_25748);
or U34420 (N_34420,N_28346,N_24028);
and U34421 (N_34421,N_27579,N_27745);
nor U34422 (N_34422,N_28196,N_28884);
or U34423 (N_34423,N_27020,N_20330);
or U34424 (N_34424,N_28232,N_20401);
xor U34425 (N_34425,N_22643,N_20769);
nor U34426 (N_34426,N_21656,N_23358);
or U34427 (N_34427,N_29624,N_24676);
or U34428 (N_34428,N_29381,N_27156);
nand U34429 (N_34429,N_25947,N_20047);
nand U34430 (N_34430,N_21650,N_26725);
nand U34431 (N_34431,N_28270,N_23680);
xor U34432 (N_34432,N_22067,N_29781);
nor U34433 (N_34433,N_23173,N_21855);
xnor U34434 (N_34434,N_29299,N_23051);
xnor U34435 (N_34435,N_23797,N_26968);
and U34436 (N_34436,N_21612,N_29644);
xor U34437 (N_34437,N_29881,N_29309);
or U34438 (N_34438,N_21407,N_20908);
nand U34439 (N_34439,N_28926,N_20629);
and U34440 (N_34440,N_29149,N_22794);
and U34441 (N_34441,N_28547,N_24871);
or U34442 (N_34442,N_20574,N_22759);
and U34443 (N_34443,N_23897,N_21762);
nand U34444 (N_34444,N_28047,N_21050);
xnor U34445 (N_34445,N_20033,N_21820);
or U34446 (N_34446,N_29804,N_21318);
or U34447 (N_34447,N_23374,N_24617);
or U34448 (N_34448,N_22926,N_21581);
nor U34449 (N_34449,N_25076,N_24049);
nand U34450 (N_34450,N_25936,N_24291);
nand U34451 (N_34451,N_26857,N_23563);
or U34452 (N_34452,N_21341,N_29018);
or U34453 (N_34453,N_20490,N_24517);
nor U34454 (N_34454,N_20295,N_22666);
or U34455 (N_34455,N_25142,N_21134);
nand U34456 (N_34456,N_24602,N_28693);
nand U34457 (N_34457,N_20251,N_27708);
xnor U34458 (N_34458,N_22580,N_26537);
nand U34459 (N_34459,N_28130,N_23682);
nand U34460 (N_34460,N_28560,N_24791);
and U34461 (N_34461,N_22330,N_24639);
xnor U34462 (N_34462,N_25987,N_27386);
and U34463 (N_34463,N_27110,N_23410);
or U34464 (N_34464,N_27829,N_23640);
nor U34465 (N_34465,N_29522,N_22532);
or U34466 (N_34466,N_28579,N_29308);
or U34467 (N_34467,N_22002,N_28942);
nand U34468 (N_34468,N_23127,N_27011);
nor U34469 (N_34469,N_29956,N_22650);
or U34470 (N_34470,N_20563,N_27312);
and U34471 (N_34471,N_28543,N_24457);
nor U34472 (N_34472,N_24675,N_24434);
and U34473 (N_34473,N_26187,N_20395);
nand U34474 (N_34474,N_27522,N_29303);
nor U34475 (N_34475,N_22876,N_25241);
or U34476 (N_34476,N_21639,N_27048);
nor U34477 (N_34477,N_27820,N_20204);
nor U34478 (N_34478,N_25491,N_20329);
nand U34479 (N_34479,N_22066,N_22157);
nor U34480 (N_34480,N_21029,N_20764);
nor U34481 (N_34481,N_24175,N_21099);
and U34482 (N_34482,N_25579,N_25573);
or U34483 (N_34483,N_27208,N_20877);
nor U34484 (N_34484,N_29013,N_22673);
nor U34485 (N_34485,N_20151,N_28919);
nand U34486 (N_34486,N_24630,N_22278);
or U34487 (N_34487,N_29218,N_23783);
and U34488 (N_34488,N_25330,N_28090);
nor U34489 (N_34489,N_29947,N_24607);
or U34490 (N_34490,N_20034,N_21728);
or U34491 (N_34491,N_23820,N_21307);
and U34492 (N_34492,N_27154,N_28420);
nand U34493 (N_34493,N_27686,N_27762);
and U34494 (N_34494,N_22023,N_23688);
and U34495 (N_34495,N_24771,N_23836);
nand U34496 (N_34496,N_21095,N_24450);
nor U34497 (N_34497,N_23731,N_22663);
and U34498 (N_34498,N_22627,N_26726);
or U34499 (N_34499,N_29325,N_28907);
xor U34500 (N_34500,N_25119,N_24090);
nand U34501 (N_34501,N_27049,N_25268);
and U34502 (N_34502,N_29651,N_20614);
or U34503 (N_34503,N_25456,N_23735);
nand U34504 (N_34504,N_21832,N_22403);
or U34505 (N_34505,N_26653,N_26738);
or U34506 (N_34506,N_20812,N_22390);
or U34507 (N_34507,N_23238,N_21221);
and U34508 (N_34508,N_25015,N_25449);
nand U34509 (N_34509,N_29026,N_22076);
nor U34510 (N_34510,N_23155,N_21740);
nor U34511 (N_34511,N_27778,N_29754);
nand U34512 (N_34512,N_26088,N_29191);
xor U34513 (N_34513,N_29053,N_28407);
or U34514 (N_34514,N_20436,N_24377);
nor U34515 (N_34515,N_21679,N_20441);
xor U34516 (N_34516,N_22929,N_22326);
nand U34517 (N_34517,N_22616,N_23973);
nor U34518 (N_34518,N_23831,N_26447);
nand U34519 (N_34519,N_20375,N_23219);
and U34520 (N_34520,N_28692,N_28135);
and U34521 (N_34521,N_26923,N_23035);
nor U34522 (N_34522,N_29115,N_28742);
and U34523 (N_34523,N_21096,N_22537);
nand U34524 (N_34524,N_23601,N_28290);
and U34525 (N_34525,N_24343,N_24383);
nand U34526 (N_34526,N_29083,N_21478);
and U34527 (N_34527,N_25774,N_27183);
xnor U34528 (N_34528,N_27831,N_27765);
nor U34529 (N_34529,N_28101,N_20837);
or U34530 (N_34530,N_21725,N_23366);
nor U34531 (N_34531,N_27086,N_27954);
xnor U34532 (N_34532,N_23540,N_20411);
nor U34533 (N_34533,N_27843,N_28887);
nand U34534 (N_34534,N_25981,N_22151);
and U34535 (N_34535,N_24286,N_28208);
nor U34536 (N_34536,N_28339,N_29553);
nor U34537 (N_34537,N_24665,N_25030);
or U34538 (N_34538,N_20502,N_26478);
nand U34539 (N_34539,N_24185,N_23896);
nor U34540 (N_34540,N_22835,N_22993);
and U34541 (N_34541,N_20994,N_25293);
or U34542 (N_34542,N_24964,N_25580);
nand U34543 (N_34543,N_28752,N_24141);
and U34544 (N_34544,N_25813,N_20407);
and U34545 (N_34545,N_24842,N_20101);
or U34546 (N_34546,N_29582,N_22018);
and U34547 (N_34547,N_22137,N_28665);
or U34548 (N_34548,N_29444,N_25272);
or U34549 (N_34549,N_21647,N_24820);
xnor U34550 (N_34550,N_29346,N_22005);
and U34551 (N_34551,N_25300,N_22102);
or U34552 (N_34552,N_29964,N_29423);
and U34553 (N_34553,N_28043,N_28592);
nand U34554 (N_34554,N_23001,N_21553);
and U34555 (N_34555,N_26299,N_28411);
and U34556 (N_34556,N_28274,N_25583);
nand U34557 (N_34557,N_22562,N_21918);
nand U34558 (N_34558,N_28862,N_23026);
nor U34559 (N_34559,N_27094,N_28432);
and U34560 (N_34560,N_28616,N_29683);
or U34561 (N_34561,N_27529,N_22731);
or U34562 (N_34562,N_23027,N_21713);
and U34563 (N_34563,N_28446,N_29063);
nor U34564 (N_34564,N_24788,N_26260);
nand U34565 (N_34565,N_28698,N_22286);
and U34566 (N_34566,N_28296,N_26328);
nand U34567 (N_34567,N_27091,N_25551);
nand U34568 (N_34568,N_28668,N_26854);
xor U34569 (N_34569,N_26974,N_20189);
xor U34570 (N_34570,N_24942,N_24625);
or U34571 (N_34571,N_29235,N_28702);
nand U34572 (N_34572,N_29059,N_28394);
nand U34573 (N_34573,N_26701,N_21315);
nand U34574 (N_34574,N_21064,N_21956);
nor U34575 (N_34575,N_22307,N_23439);
and U34576 (N_34576,N_25130,N_24244);
nor U34577 (N_34577,N_27287,N_29958);
nor U34578 (N_34578,N_20552,N_20388);
nor U34579 (N_34579,N_22849,N_21112);
and U34580 (N_34580,N_29513,N_24853);
nand U34581 (N_34581,N_24830,N_23162);
and U34582 (N_34582,N_27661,N_25872);
or U34583 (N_34583,N_27962,N_27414);
and U34584 (N_34584,N_22030,N_28388);
xnor U34585 (N_34585,N_28010,N_20834);
nor U34586 (N_34586,N_20942,N_27223);
or U34587 (N_34587,N_28044,N_26381);
nor U34588 (N_34588,N_24785,N_20548);
nor U34589 (N_34589,N_20728,N_21971);
and U34590 (N_34590,N_27012,N_23627);
nor U34591 (N_34591,N_22753,N_25787);
and U34592 (N_34592,N_22499,N_26612);
nor U34593 (N_34593,N_24274,N_28770);
nand U34594 (N_34594,N_28602,N_25495);
nand U34595 (N_34595,N_28437,N_26811);
nor U34596 (N_34596,N_20758,N_25483);
or U34597 (N_34597,N_29126,N_26252);
nor U34598 (N_34598,N_22640,N_24584);
nor U34599 (N_34599,N_22619,N_20026);
nor U34600 (N_34600,N_22087,N_20527);
and U34601 (N_34601,N_21036,N_27933);
nor U34602 (N_34602,N_25963,N_27673);
or U34603 (N_34603,N_29354,N_21551);
nand U34604 (N_34604,N_29606,N_22719);
and U34605 (N_34605,N_22225,N_28836);
nand U34606 (N_34606,N_27358,N_26730);
nor U34607 (N_34607,N_24891,N_22109);
xor U34608 (N_34608,N_21115,N_26832);
and U34609 (N_34609,N_22545,N_22895);
nor U34610 (N_34610,N_24798,N_24977);
or U34611 (N_34611,N_28083,N_26163);
xor U34612 (N_34612,N_21739,N_24951);
or U34613 (N_34613,N_29763,N_28390);
nand U34614 (N_34614,N_22525,N_27578);
nor U34615 (N_34615,N_22638,N_26468);
nor U34616 (N_34616,N_21750,N_22878);
nor U34617 (N_34617,N_21523,N_28891);
and U34618 (N_34618,N_27793,N_29739);
and U34619 (N_34619,N_29969,N_25628);
and U34620 (N_34620,N_22275,N_28332);
and U34621 (N_34621,N_21490,N_27729);
xor U34622 (N_34622,N_26112,N_22756);
nand U34623 (N_34623,N_29328,N_28943);
nand U34624 (N_34624,N_24249,N_27734);
xor U34625 (N_34625,N_27335,N_26842);
and U34626 (N_34626,N_27757,N_20191);
nand U34627 (N_34627,N_24682,N_26119);
or U34628 (N_34628,N_21336,N_20010);
nand U34629 (N_34629,N_28933,N_20514);
and U34630 (N_34630,N_23363,N_29377);
nor U34631 (N_34631,N_28748,N_22466);
xnor U34632 (N_34632,N_24742,N_29167);
nor U34633 (N_34633,N_24340,N_22795);
nand U34634 (N_34634,N_29813,N_23268);
and U34635 (N_34635,N_20722,N_26975);
or U34636 (N_34636,N_21213,N_29098);
nand U34637 (N_34637,N_20773,N_23588);
nor U34638 (N_34638,N_29383,N_24916);
nand U34639 (N_34639,N_24744,N_25429);
or U34640 (N_34640,N_26896,N_23402);
nand U34641 (N_34641,N_24770,N_24151);
or U34642 (N_34642,N_20437,N_24521);
or U34643 (N_34643,N_24348,N_23269);
nor U34644 (N_34644,N_26582,N_26000);
nor U34645 (N_34645,N_20272,N_22944);
or U34646 (N_34646,N_25759,N_23591);
and U34647 (N_34647,N_21324,N_20841);
and U34648 (N_34648,N_23256,N_23210);
or U34649 (N_34649,N_25068,N_27664);
nand U34650 (N_34650,N_26387,N_22127);
nor U34651 (N_34651,N_25242,N_26268);
nor U34652 (N_34652,N_25838,N_20338);
nand U34653 (N_34653,N_28137,N_24939);
nand U34654 (N_34654,N_29728,N_29949);
xor U34655 (N_34655,N_26396,N_27115);
and U34656 (N_34656,N_25273,N_20689);
nand U34657 (N_34657,N_28190,N_28790);
nor U34658 (N_34658,N_25179,N_24358);
nor U34659 (N_34659,N_29850,N_21056);
or U34660 (N_34660,N_29416,N_23987);
xnor U34661 (N_34661,N_25326,N_28853);
xnor U34662 (N_34662,N_27204,N_26995);
nor U34663 (N_34663,N_28001,N_26373);
and U34664 (N_34664,N_28464,N_29550);
nor U34665 (N_34665,N_21723,N_25615);
or U34666 (N_34666,N_20962,N_26800);
nor U34667 (N_34667,N_23252,N_28380);
and U34668 (N_34668,N_29036,N_21091);
nor U34669 (N_34669,N_27010,N_28112);
and U34670 (N_34670,N_23782,N_29740);
and U34671 (N_34671,N_24066,N_20296);
nor U34672 (N_34672,N_23076,N_20190);
nor U34673 (N_34673,N_28905,N_22743);
nor U34674 (N_34674,N_23415,N_22243);
nor U34675 (N_34675,N_25058,N_21330);
nor U34676 (N_34676,N_20266,N_26171);
nand U34677 (N_34677,N_25753,N_26798);
nand U34678 (N_34678,N_27305,N_29970);
xnor U34679 (N_34679,N_20875,N_20926);
nand U34680 (N_34680,N_25567,N_27174);
xor U34681 (N_34681,N_28603,N_27045);
nand U34682 (N_34682,N_26436,N_21417);
xor U34683 (N_34683,N_20232,N_24275);
nor U34684 (N_34684,N_24421,N_28237);
or U34685 (N_34685,N_28056,N_23889);
nand U34686 (N_34686,N_25596,N_26403);
or U34687 (N_34687,N_21795,N_21353);
nor U34688 (N_34688,N_24807,N_24092);
and U34689 (N_34689,N_24407,N_29156);
nor U34690 (N_34690,N_24782,N_22200);
and U34691 (N_34691,N_22226,N_27836);
nand U34692 (N_34692,N_20553,N_28674);
nand U34693 (N_34693,N_23282,N_21771);
xor U34694 (N_34694,N_25311,N_25140);
nand U34695 (N_34695,N_28835,N_27787);
xor U34696 (N_34696,N_22021,N_29623);
nand U34697 (N_34697,N_21444,N_27343);
and U34698 (N_34698,N_24691,N_25805);
or U34699 (N_34699,N_24437,N_21183);
or U34700 (N_34700,N_20104,N_24522);
nor U34701 (N_34701,N_23240,N_21299);
and U34702 (N_34702,N_26609,N_29795);
or U34703 (N_34703,N_28882,N_20170);
xor U34704 (N_34704,N_28893,N_21904);
xor U34705 (N_34705,N_27103,N_28026);
or U34706 (N_34706,N_25572,N_21090);
nand U34707 (N_34707,N_22472,N_22573);
nand U34708 (N_34708,N_25920,N_25504);
xor U34709 (N_34709,N_25526,N_29931);
nor U34710 (N_34710,N_28147,N_27446);
or U34711 (N_34711,N_22885,N_29333);
and U34712 (N_34712,N_26310,N_29046);
xnor U34713 (N_34713,N_26684,N_23551);
nor U34714 (N_34714,N_24413,N_26744);
or U34715 (N_34715,N_22775,N_21168);
or U34716 (N_34716,N_20609,N_28623);
or U34717 (N_34717,N_28506,N_21450);
nand U34718 (N_34718,N_20378,N_23828);
nand U34719 (N_34719,N_28477,N_29467);
nand U34720 (N_34720,N_20471,N_20473);
nand U34721 (N_34721,N_26860,N_23576);
nor U34722 (N_34722,N_27517,N_23003);
nor U34723 (N_34723,N_25174,N_25662);
and U34724 (N_34724,N_22763,N_21101);
nand U34725 (N_34725,N_27622,N_22196);
xnor U34726 (N_34726,N_24850,N_27653);
or U34727 (N_34727,N_22934,N_27144);
xor U34728 (N_34728,N_22862,N_27652);
nor U34729 (N_34729,N_24550,N_26826);
nand U34730 (N_34730,N_27194,N_24145);
or U34731 (N_34731,N_28964,N_21053);
and U34732 (N_34732,N_25226,N_28416);
and U34733 (N_34733,N_27095,N_21087);
nor U34734 (N_34734,N_24080,N_25117);
xor U34735 (N_34735,N_20524,N_29245);
nor U34736 (N_34736,N_20435,N_24253);
nand U34737 (N_34737,N_21075,N_25172);
and U34738 (N_34738,N_22810,N_23900);
nor U34739 (N_34739,N_23665,N_24519);
nand U34740 (N_34740,N_28615,N_23830);
nor U34741 (N_34741,N_24396,N_24303);
xnor U34742 (N_34742,N_23585,N_29326);
or U34743 (N_34743,N_24052,N_29400);
and U34744 (N_34744,N_21877,N_20621);
nor U34745 (N_34745,N_21700,N_28204);
and U34746 (N_34746,N_22247,N_29228);
and U34747 (N_34747,N_25256,N_26439);
nor U34748 (N_34748,N_21184,N_24347);
nand U34749 (N_34749,N_26531,N_23736);
nand U34750 (N_34750,N_29694,N_28696);
or U34751 (N_34751,N_21519,N_21487);
nor U34752 (N_34752,N_27620,N_22138);
nor U34753 (N_34753,N_29608,N_28094);
xor U34754 (N_34754,N_25844,N_23639);
nor U34755 (N_34755,N_24563,N_24069);
and U34756 (N_34756,N_20333,N_20711);
nor U34757 (N_34757,N_27249,N_21710);
nor U34758 (N_34758,N_26926,N_25797);
or U34759 (N_34759,N_29669,N_28401);
nand U34760 (N_34760,N_22322,N_23970);
nor U34761 (N_34761,N_27670,N_22259);
or U34762 (N_34762,N_29032,N_21313);
and U34763 (N_34763,N_27473,N_29537);
nor U34764 (N_34764,N_26637,N_22367);
or U34765 (N_34765,N_21748,N_25212);
or U34766 (N_34766,N_25034,N_23984);
nor U34767 (N_34767,N_29672,N_23037);
or U34768 (N_34768,N_22870,N_25041);
xnor U34769 (N_34769,N_21496,N_22345);
nor U34770 (N_34770,N_24478,N_20312);
or U34771 (N_34771,N_20858,N_25839);
or U34772 (N_34772,N_23367,N_24393);
nand U34773 (N_34773,N_28885,N_27973);
xnor U34774 (N_34774,N_25227,N_25934);
nor U34775 (N_34775,N_26634,N_26950);
or U34776 (N_34776,N_25094,N_20277);
and U34777 (N_34777,N_21932,N_29374);
nor U34778 (N_34778,N_26795,N_20840);
or U34779 (N_34779,N_22145,N_29435);
and U34780 (N_34780,N_20529,N_26546);
nand U34781 (N_34781,N_25738,N_29384);
and U34782 (N_34782,N_20763,N_20756);
and U34783 (N_34783,N_28348,N_28609);
xnor U34784 (N_34784,N_26295,N_21019);
nor U34785 (N_34785,N_28889,N_27388);
nand U34786 (N_34786,N_26404,N_21787);
nor U34787 (N_34787,N_21010,N_24659);
nor U34788 (N_34788,N_24243,N_28435);
and U34789 (N_34789,N_21135,N_29120);
nor U34790 (N_34790,N_27028,N_22274);
nor U34791 (N_34791,N_29237,N_28909);
xnor U34792 (N_34792,N_25950,N_20370);
nor U34793 (N_34793,N_20787,N_25144);
nand U34794 (N_34794,N_27053,N_22949);
or U34795 (N_34795,N_26071,N_23700);
and U34796 (N_34796,N_27041,N_22485);
nor U34797 (N_34797,N_20182,N_28523);
and U34798 (N_34798,N_22348,N_28751);
nor U34799 (N_34799,N_24008,N_26005);
or U34800 (N_34800,N_29704,N_25840);
xor U34801 (N_34801,N_21582,N_26234);
nand U34802 (N_34802,N_24415,N_27756);
or U34803 (N_34803,N_28162,N_21547);
or U34804 (N_34804,N_29236,N_20607);
nand U34805 (N_34805,N_22718,N_20241);
nand U34806 (N_34806,N_24992,N_27679);
or U34807 (N_34807,N_27834,N_23873);
nand U34808 (N_34808,N_26294,N_27377);
nand U34809 (N_34809,N_27445,N_20690);
and U34810 (N_34810,N_25164,N_28353);
nand U34811 (N_34811,N_23936,N_24664);
and U34812 (N_34812,N_25524,N_25318);
or U34813 (N_34813,N_21383,N_21917);
or U34814 (N_34814,N_23262,N_26560);
nor U34815 (N_34815,N_22316,N_29247);
xor U34816 (N_34816,N_22328,N_23714);
or U34817 (N_34817,N_20107,N_23000);
nor U34818 (N_34818,N_27170,N_29342);
and U34819 (N_34819,N_20002,N_26307);
nand U34820 (N_34820,N_26672,N_21711);
or U34821 (N_34821,N_23877,N_26869);
nor U34822 (N_34822,N_24777,N_22379);
nand U34823 (N_34823,N_20583,N_22542);
nor U34824 (N_34824,N_29282,N_22434);
nor U34825 (N_34825,N_27978,N_24595);
nand U34826 (N_34826,N_22346,N_22528);
and U34827 (N_34827,N_21013,N_24862);
nor U34828 (N_34828,N_27419,N_23199);
nand U34829 (N_34829,N_21483,N_26398);
and U34830 (N_34830,N_29990,N_26292);
nand U34831 (N_34831,N_20202,N_27870);
and U34832 (N_34832,N_27282,N_24497);
xnor U34833 (N_34833,N_26322,N_27635);
and U34834 (N_34834,N_28267,N_25447);
and U34835 (N_34835,N_24526,N_22460);
nand U34836 (N_34836,N_26029,N_25031);
and U34837 (N_34837,N_24501,N_25571);
or U34838 (N_34838,N_22468,N_24778);
nand U34839 (N_34839,N_25477,N_25043);
nor U34840 (N_34840,N_20571,N_24181);
nand U34841 (N_34841,N_21617,N_25252);
nand U34842 (N_34842,N_21464,N_26692);
and U34843 (N_34843,N_20117,N_23886);
nor U34844 (N_34844,N_27203,N_20453);
and U34845 (N_34845,N_29439,N_28733);
nand U34846 (N_34846,N_22891,N_21001);
nor U34847 (N_34847,N_25020,N_28076);
xnor U34848 (N_34848,N_25785,N_23986);
xor U34849 (N_34849,N_24483,N_26279);
xnor U34850 (N_34850,N_20431,N_21408);
nor U34851 (N_34851,N_20727,N_26423);
or U34852 (N_34852,N_20321,N_24433);
or U34853 (N_34853,N_24740,N_21705);
nor U34854 (N_34854,N_24935,N_29287);
nand U34855 (N_34855,N_29995,N_24403);
or U34856 (N_34856,N_21631,N_25135);
nand U34857 (N_34857,N_25328,N_21105);
nor U34858 (N_34858,N_28344,N_28170);
and U34859 (N_34859,N_21873,N_22459);
nor U34860 (N_34860,N_21179,N_27739);
xor U34861 (N_34861,N_25459,N_26334);
and U34862 (N_34862,N_27093,N_25059);
or U34863 (N_34863,N_28033,N_24025);
or U34864 (N_34864,N_29851,N_20348);
and U34865 (N_34865,N_20121,N_21445);
nor U34866 (N_34866,N_29873,N_27619);
nand U34867 (N_34867,N_20936,N_26658);
or U34868 (N_34868,N_27323,N_21894);
nand U34869 (N_34869,N_28260,N_29633);
nor U34870 (N_34870,N_28793,N_27320);
nand U34871 (N_34871,N_21008,N_22783);
or U34872 (N_34872,N_26323,N_25989);
nor U34873 (N_34873,N_26245,N_25363);
nand U34874 (N_34874,N_20413,N_23457);
or U34875 (N_34875,N_28381,N_25896);
nand U34876 (N_34876,N_24912,N_26607);
nand U34877 (N_34877,N_21630,N_28035);
and U34878 (N_34878,N_21428,N_27738);
nor U34879 (N_34879,N_21913,N_20664);
nand U34880 (N_34880,N_22488,N_20871);
or U34881 (N_34881,N_26388,N_27311);
xor U34882 (N_34882,N_20253,N_26745);
xnor U34883 (N_34883,N_21626,N_20147);
or U34884 (N_34884,N_24623,N_23373);
nor U34885 (N_34885,N_21279,N_20929);
and U34886 (N_34886,N_25616,N_23565);
and U34887 (N_34887,N_21028,N_24338);
xor U34888 (N_34888,N_24674,N_25915);
or U34889 (N_34889,N_21163,N_20380);
nor U34890 (N_34890,N_23041,N_27486);
or U34891 (N_34891,N_23314,N_29163);
or U34892 (N_34892,N_25129,N_26733);
nand U34893 (N_34893,N_28364,N_25733);
nand U34894 (N_34894,N_27662,N_26835);
and U34895 (N_34895,N_29563,N_26602);
nor U34896 (N_34896,N_20085,N_22597);
nand U34897 (N_34897,N_22576,N_25342);
nor U34898 (N_34898,N_21114,N_25866);
or U34899 (N_34899,N_20578,N_24897);
nand U34900 (N_34900,N_29215,N_22770);
nor U34901 (N_34901,N_20143,N_20390);
xnor U34902 (N_34902,N_25206,N_29961);
and U34903 (N_34903,N_21870,N_29912);
and U34904 (N_34904,N_24398,N_25303);
and U34905 (N_34905,N_28251,N_24756);
and U34906 (N_34906,N_20018,N_26385);
and U34907 (N_34907,N_27727,N_24099);
or U34908 (N_34908,N_20181,N_28227);
and U34909 (N_34909,N_25482,N_26987);
or U34910 (N_34910,N_25806,N_24555);
xnor U34911 (N_34911,N_26475,N_20257);
nor U34912 (N_34912,N_28629,N_28871);
and U34913 (N_34913,N_21104,N_27556);
nor U34914 (N_34914,N_28979,N_26231);
xnor U34915 (N_34915,N_21627,N_27074);
or U34916 (N_34916,N_25908,N_26605);
or U34917 (N_34917,N_25412,N_29504);
or U34918 (N_34918,N_29166,N_23260);
nor U34919 (N_34919,N_21435,N_20184);
and U34920 (N_34920,N_20352,N_27993);
nand U34921 (N_34921,N_27205,N_28873);
nor U34922 (N_34922,N_23953,N_26830);
nand U34923 (N_34923,N_25228,N_24310);
xnor U34924 (N_34924,N_24448,N_28286);
and U34925 (N_34925,N_23017,N_23528);
and U34926 (N_34926,N_23574,N_26929);
and U34927 (N_34927,N_25465,N_29196);
nand U34928 (N_34928,N_21908,N_27932);
and U34929 (N_34929,N_23884,N_29864);
or U34930 (N_34930,N_27647,N_25828);
nor U34931 (N_34931,N_23304,N_27817);
nand U34932 (N_34932,N_25550,N_20070);
xor U34933 (N_34933,N_21593,N_22746);
or U34934 (N_34934,N_22984,N_29061);
nand U34935 (N_34935,N_24649,N_29021);
nand U34936 (N_34936,N_28230,N_26971);
nor U34937 (N_34937,N_25754,N_24993);
nand U34938 (N_34938,N_22502,N_27448);
nand U34939 (N_34939,N_25959,N_21329);
or U34940 (N_34940,N_20909,N_27908);
nand U34941 (N_34941,N_26661,N_24081);
nor U34942 (N_34942,N_21926,N_21802);
nor U34943 (N_34943,N_28308,N_28171);
nor U34944 (N_34944,N_23438,N_21290);
nor U34945 (N_34945,N_21722,N_29242);
nand U34946 (N_34946,N_22456,N_28544);
nor U34947 (N_34947,N_20977,N_24115);
nand U34948 (N_34948,N_21068,N_26114);
nor U34949 (N_34949,N_22564,N_28368);
and U34950 (N_34950,N_27380,N_26140);
nor U34951 (N_34951,N_22121,N_25654);
nand U34952 (N_34952,N_28483,N_29777);
xor U34953 (N_34953,N_21473,N_27655);
nor U34954 (N_34954,N_27923,N_24781);
and U34955 (N_34955,N_23113,N_22735);
nor U34956 (N_34956,N_27939,N_24021);
or U34957 (N_34957,N_28050,N_21858);
nor U34958 (N_34958,N_28982,N_26559);
and U34959 (N_34959,N_28582,N_27454);
and U34960 (N_34960,N_24068,N_29339);
nand U34961 (N_34961,N_27769,N_29443);
nor U34962 (N_34962,N_27776,N_24677);
or U34963 (N_34963,N_26918,N_27469);
or U34964 (N_34964,N_22156,N_23197);
xnor U34965 (N_34965,N_23818,N_25035);
or U34966 (N_34966,N_21822,N_28418);
or U34967 (N_34967,N_22290,N_20522);
and U34968 (N_34968,N_24738,N_21986);
nor U34969 (N_34969,N_21089,N_23296);
nor U34970 (N_34970,N_29392,N_23279);
nor U34971 (N_34971,N_29125,N_27863);
or U34972 (N_34972,N_21702,N_29278);
nand U34973 (N_34973,N_27272,N_23263);
or U34974 (N_34974,N_27559,N_21962);
or U34975 (N_34975,N_26773,N_25545);
or U34976 (N_34976,N_27182,N_20149);
nand U34977 (N_34977,N_21546,N_29846);
or U34978 (N_34978,N_28879,N_24125);
nor U34979 (N_34979,N_25536,N_20360);
or U34980 (N_34980,N_21781,N_26117);
nor U34981 (N_34981,N_29173,N_20317);
or U34982 (N_34982,N_27404,N_24567);
and U34983 (N_34983,N_25651,N_24105);
xor U34984 (N_34984,N_29315,N_24182);
or U34985 (N_34985,N_20886,N_29520);
and U34986 (N_34986,N_26783,N_27680);
nand U34987 (N_34987,N_29802,N_26103);
nor U34988 (N_34988,N_28827,N_25315);
nor U34989 (N_34989,N_23161,N_27909);
nand U34990 (N_34990,N_29695,N_22645);
or U34991 (N_34991,N_24059,N_28796);
and U34992 (N_34992,N_26151,N_27067);
nand U34993 (N_34993,N_24737,N_23408);
nor U34994 (N_34994,N_28293,N_24002);
or U34995 (N_34995,N_27896,N_22368);
xor U34996 (N_34996,N_22762,N_26056);
and U34997 (N_34997,N_25613,N_28447);
nor U34998 (N_34998,N_22507,N_23132);
or U34999 (N_34999,N_24222,N_25875);
nor U35000 (N_35000,N_23870,N_21920);
or U35001 (N_35001,N_22775,N_20211);
nor U35002 (N_35002,N_27487,N_20669);
nor U35003 (N_35003,N_22612,N_28558);
or U35004 (N_35004,N_22791,N_21424);
nor U35005 (N_35005,N_27228,N_20308);
or U35006 (N_35006,N_25766,N_23050);
or U35007 (N_35007,N_20939,N_26282);
nor U35008 (N_35008,N_24743,N_23295);
or U35009 (N_35009,N_28244,N_21486);
nor U35010 (N_35010,N_25250,N_26852);
and U35011 (N_35011,N_27341,N_28757);
and U35012 (N_35012,N_25436,N_21544);
nor U35013 (N_35013,N_26748,N_25998);
nand U35014 (N_35014,N_22251,N_20656);
nand U35015 (N_35015,N_25995,N_21791);
and U35016 (N_35016,N_23248,N_23668);
and U35017 (N_35017,N_27090,N_21834);
and U35018 (N_35018,N_28924,N_23303);
nand U35019 (N_35019,N_24877,N_28795);
nor U35020 (N_35020,N_24966,N_26851);
or U35021 (N_35021,N_24247,N_20744);
and U35022 (N_35022,N_21583,N_25507);
and U35023 (N_35023,N_23453,N_22419);
xor U35024 (N_35024,N_24525,N_20205);
nand U35025 (N_35025,N_25703,N_22885);
xor U35026 (N_35026,N_26232,N_22191);
nor U35027 (N_35027,N_26186,N_21429);
or U35028 (N_35028,N_21725,N_22599);
nor U35029 (N_35029,N_24619,N_26738);
nand U35030 (N_35030,N_24284,N_28253);
and U35031 (N_35031,N_22837,N_29131);
and U35032 (N_35032,N_20516,N_26194);
and U35033 (N_35033,N_27906,N_28666);
nor U35034 (N_35034,N_23029,N_23464);
and U35035 (N_35035,N_20910,N_21168);
nor U35036 (N_35036,N_28408,N_20080);
or U35037 (N_35037,N_29547,N_26831);
and U35038 (N_35038,N_22359,N_25096);
nor U35039 (N_35039,N_20569,N_22962);
and U35040 (N_35040,N_23787,N_26527);
or U35041 (N_35041,N_23179,N_29432);
nor U35042 (N_35042,N_27015,N_29615);
or U35043 (N_35043,N_24761,N_27969);
and U35044 (N_35044,N_20601,N_28744);
nand U35045 (N_35045,N_22913,N_21558);
or U35046 (N_35046,N_25249,N_26430);
nand U35047 (N_35047,N_23251,N_24915);
and U35048 (N_35048,N_26676,N_24718);
nor U35049 (N_35049,N_23720,N_25894);
nand U35050 (N_35050,N_22243,N_23555);
nand U35051 (N_35051,N_21795,N_20728);
and U35052 (N_35052,N_28630,N_23726);
xor U35053 (N_35053,N_29054,N_20070);
or U35054 (N_35054,N_20870,N_24334);
nand U35055 (N_35055,N_24363,N_24596);
and U35056 (N_35056,N_21512,N_24569);
or U35057 (N_35057,N_28338,N_28913);
nor U35058 (N_35058,N_26711,N_21283);
or U35059 (N_35059,N_22492,N_20595);
or U35060 (N_35060,N_23494,N_20908);
or U35061 (N_35061,N_21130,N_21006);
nor U35062 (N_35062,N_20316,N_21648);
nor U35063 (N_35063,N_28446,N_26299);
or U35064 (N_35064,N_25922,N_24941);
and U35065 (N_35065,N_28521,N_27560);
and U35066 (N_35066,N_27721,N_21281);
and U35067 (N_35067,N_27209,N_29293);
or U35068 (N_35068,N_24592,N_24006);
and U35069 (N_35069,N_29005,N_28985);
and U35070 (N_35070,N_29197,N_26500);
and U35071 (N_35071,N_23440,N_22967);
nor U35072 (N_35072,N_28304,N_26485);
nand U35073 (N_35073,N_29050,N_22159);
and U35074 (N_35074,N_27001,N_21664);
xnor U35075 (N_35075,N_28442,N_23924);
or U35076 (N_35076,N_24166,N_23955);
nand U35077 (N_35077,N_21838,N_24664);
nand U35078 (N_35078,N_29867,N_26768);
nand U35079 (N_35079,N_28621,N_28958);
and U35080 (N_35080,N_26122,N_27643);
nor U35081 (N_35081,N_29575,N_24096);
xor U35082 (N_35082,N_24154,N_27710);
or U35083 (N_35083,N_29678,N_28519);
nor U35084 (N_35084,N_22605,N_28064);
nor U35085 (N_35085,N_21340,N_21232);
nor U35086 (N_35086,N_23764,N_20270);
nor U35087 (N_35087,N_27946,N_24176);
xnor U35088 (N_35088,N_22376,N_21708);
nand U35089 (N_35089,N_25293,N_24986);
nor U35090 (N_35090,N_21513,N_21123);
nand U35091 (N_35091,N_20746,N_23142);
nand U35092 (N_35092,N_20415,N_29717);
nor U35093 (N_35093,N_21302,N_23777);
nand U35094 (N_35094,N_22332,N_29939);
or U35095 (N_35095,N_27922,N_29058);
xnor U35096 (N_35096,N_25933,N_23284);
nand U35097 (N_35097,N_20510,N_27444);
and U35098 (N_35098,N_21421,N_21058);
nor U35099 (N_35099,N_20445,N_21114);
nor U35100 (N_35100,N_25320,N_20980);
and U35101 (N_35101,N_21641,N_28815);
xor U35102 (N_35102,N_24643,N_22667);
and U35103 (N_35103,N_26101,N_24428);
nor U35104 (N_35104,N_28342,N_22175);
nand U35105 (N_35105,N_24786,N_28413);
nand U35106 (N_35106,N_25405,N_24395);
or U35107 (N_35107,N_21688,N_28312);
or U35108 (N_35108,N_22081,N_29467);
nand U35109 (N_35109,N_26200,N_26880);
nor U35110 (N_35110,N_20702,N_25850);
and U35111 (N_35111,N_28122,N_26797);
nand U35112 (N_35112,N_27306,N_21519);
nand U35113 (N_35113,N_27126,N_28562);
and U35114 (N_35114,N_22272,N_24954);
nand U35115 (N_35115,N_29910,N_22776);
nor U35116 (N_35116,N_29120,N_24941);
nand U35117 (N_35117,N_24735,N_21887);
or U35118 (N_35118,N_29126,N_25476);
nor U35119 (N_35119,N_26341,N_27938);
nor U35120 (N_35120,N_24614,N_28831);
and U35121 (N_35121,N_21480,N_22235);
and U35122 (N_35122,N_28840,N_29875);
or U35123 (N_35123,N_22614,N_27022);
nand U35124 (N_35124,N_29592,N_26906);
and U35125 (N_35125,N_27533,N_26722);
nor U35126 (N_35126,N_21225,N_28883);
nor U35127 (N_35127,N_21488,N_28233);
or U35128 (N_35128,N_20445,N_20284);
or U35129 (N_35129,N_24196,N_28002);
nor U35130 (N_35130,N_27938,N_24048);
and U35131 (N_35131,N_29811,N_25289);
nand U35132 (N_35132,N_24660,N_20801);
or U35133 (N_35133,N_21089,N_29961);
or U35134 (N_35134,N_27712,N_28706);
or U35135 (N_35135,N_28125,N_27164);
and U35136 (N_35136,N_26864,N_21193);
or U35137 (N_35137,N_24261,N_25578);
or U35138 (N_35138,N_29650,N_26671);
nor U35139 (N_35139,N_22547,N_21920);
and U35140 (N_35140,N_26915,N_23559);
nor U35141 (N_35141,N_23767,N_21351);
or U35142 (N_35142,N_20180,N_26123);
or U35143 (N_35143,N_20781,N_29294);
nor U35144 (N_35144,N_27071,N_27749);
nor U35145 (N_35145,N_20255,N_23503);
xor U35146 (N_35146,N_20410,N_21752);
nor U35147 (N_35147,N_22674,N_24607);
nand U35148 (N_35148,N_24601,N_22220);
and U35149 (N_35149,N_27557,N_20213);
nor U35150 (N_35150,N_28814,N_29156);
and U35151 (N_35151,N_23099,N_23693);
nor U35152 (N_35152,N_22877,N_20446);
nand U35153 (N_35153,N_23065,N_20776);
nor U35154 (N_35154,N_22112,N_23413);
or U35155 (N_35155,N_20032,N_25302);
nand U35156 (N_35156,N_21751,N_20108);
and U35157 (N_35157,N_20435,N_27125);
xor U35158 (N_35158,N_21594,N_22917);
or U35159 (N_35159,N_21227,N_28905);
xnor U35160 (N_35160,N_24728,N_23292);
nand U35161 (N_35161,N_22502,N_24354);
and U35162 (N_35162,N_26566,N_28344);
xor U35163 (N_35163,N_29491,N_28204);
nand U35164 (N_35164,N_27094,N_28717);
xnor U35165 (N_35165,N_22156,N_26842);
nor U35166 (N_35166,N_21805,N_29687);
nand U35167 (N_35167,N_28330,N_28069);
nor U35168 (N_35168,N_27389,N_24800);
nor U35169 (N_35169,N_23122,N_20957);
xnor U35170 (N_35170,N_24647,N_27727);
nand U35171 (N_35171,N_25654,N_27585);
nor U35172 (N_35172,N_22434,N_21742);
nor U35173 (N_35173,N_29128,N_25052);
xor U35174 (N_35174,N_25154,N_29658);
nor U35175 (N_35175,N_20335,N_25652);
and U35176 (N_35176,N_27630,N_20971);
or U35177 (N_35177,N_21719,N_24046);
nand U35178 (N_35178,N_23534,N_24760);
nor U35179 (N_35179,N_26654,N_25430);
nand U35180 (N_35180,N_25016,N_21481);
nand U35181 (N_35181,N_26649,N_28387);
nor U35182 (N_35182,N_29897,N_21346);
and U35183 (N_35183,N_21956,N_25539);
nor U35184 (N_35184,N_27484,N_25070);
nor U35185 (N_35185,N_29888,N_25656);
nand U35186 (N_35186,N_21080,N_26840);
xnor U35187 (N_35187,N_26058,N_26775);
and U35188 (N_35188,N_29124,N_22672);
or U35189 (N_35189,N_21083,N_23546);
nand U35190 (N_35190,N_26140,N_21259);
or U35191 (N_35191,N_20849,N_21285);
or U35192 (N_35192,N_20266,N_29004);
or U35193 (N_35193,N_28021,N_29302);
nand U35194 (N_35194,N_29521,N_23211);
nor U35195 (N_35195,N_25824,N_26711);
or U35196 (N_35196,N_27638,N_27870);
and U35197 (N_35197,N_22520,N_21645);
and U35198 (N_35198,N_29152,N_21365);
and U35199 (N_35199,N_27348,N_28149);
nand U35200 (N_35200,N_20039,N_26910);
and U35201 (N_35201,N_20991,N_22816);
and U35202 (N_35202,N_22780,N_21548);
or U35203 (N_35203,N_21211,N_26277);
nand U35204 (N_35204,N_25509,N_24643);
and U35205 (N_35205,N_24516,N_28511);
nor U35206 (N_35206,N_21530,N_28816);
nand U35207 (N_35207,N_20326,N_21193);
nor U35208 (N_35208,N_28708,N_22927);
or U35209 (N_35209,N_21069,N_22708);
nand U35210 (N_35210,N_24374,N_23241);
nand U35211 (N_35211,N_24541,N_22599);
nand U35212 (N_35212,N_26281,N_22506);
nor U35213 (N_35213,N_20287,N_29513);
nor U35214 (N_35214,N_21783,N_26190);
and U35215 (N_35215,N_26830,N_29762);
nor U35216 (N_35216,N_23118,N_24012);
xor U35217 (N_35217,N_25644,N_26387);
nor U35218 (N_35218,N_27257,N_28436);
and U35219 (N_35219,N_21472,N_22978);
or U35220 (N_35220,N_28751,N_25354);
nor U35221 (N_35221,N_23692,N_23827);
or U35222 (N_35222,N_20235,N_25194);
or U35223 (N_35223,N_26643,N_23253);
xor U35224 (N_35224,N_25769,N_20769);
nor U35225 (N_35225,N_20237,N_21590);
or U35226 (N_35226,N_26632,N_23850);
and U35227 (N_35227,N_24486,N_23592);
nand U35228 (N_35228,N_24589,N_23383);
nand U35229 (N_35229,N_27913,N_22808);
nor U35230 (N_35230,N_28366,N_29683);
nor U35231 (N_35231,N_24350,N_27805);
xnor U35232 (N_35232,N_21099,N_24677);
nor U35233 (N_35233,N_22473,N_26313);
or U35234 (N_35234,N_28870,N_28138);
nand U35235 (N_35235,N_24166,N_27078);
or U35236 (N_35236,N_26936,N_26379);
nor U35237 (N_35237,N_20054,N_22237);
nor U35238 (N_35238,N_26190,N_24285);
xnor U35239 (N_35239,N_26605,N_23917);
nor U35240 (N_35240,N_20772,N_25525);
nand U35241 (N_35241,N_25640,N_21279);
or U35242 (N_35242,N_27799,N_22747);
or U35243 (N_35243,N_24601,N_20082);
nand U35244 (N_35244,N_26523,N_23447);
and U35245 (N_35245,N_23871,N_22740);
and U35246 (N_35246,N_23827,N_29977);
or U35247 (N_35247,N_24886,N_23430);
and U35248 (N_35248,N_23584,N_22553);
nand U35249 (N_35249,N_24177,N_20903);
or U35250 (N_35250,N_26418,N_26067);
xor U35251 (N_35251,N_24735,N_23382);
xor U35252 (N_35252,N_25810,N_26145);
and U35253 (N_35253,N_22562,N_20803);
nand U35254 (N_35254,N_20799,N_23409);
nor U35255 (N_35255,N_20598,N_22431);
nor U35256 (N_35256,N_27184,N_25420);
and U35257 (N_35257,N_27594,N_29660);
or U35258 (N_35258,N_20298,N_20491);
nand U35259 (N_35259,N_23638,N_20950);
and U35260 (N_35260,N_21868,N_22195);
nand U35261 (N_35261,N_24322,N_22232);
nand U35262 (N_35262,N_28772,N_27164);
xor U35263 (N_35263,N_25199,N_29074);
or U35264 (N_35264,N_26906,N_24663);
nor U35265 (N_35265,N_29842,N_26202);
and U35266 (N_35266,N_25469,N_24059);
xnor U35267 (N_35267,N_24311,N_28459);
nor U35268 (N_35268,N_21256,N_26274);
and U35269 (N_35269,N_27540,N_29208);
nand U35270 (N_35270,N_21076,N_27705);
nor U35271 (N_35271,N_21861,N_24935);
nand U35272 (N_35272,N_28451,N_25639);
or U35273 (N_35273,N_21104,N_25574);
nor U35274 (N_35274,N_21384,N_22397);
nand U35275 (N_35275,N_22234,N_23415);
nand U35276 (N_35276,N_28737,N_26406);
nand U35277 (N_35277,N_27279,N_26418);
or U35278 (N_35278,N_20918,N_26764);
nor U35279 (N_35279,N_26623,N_24122);
nand U35280 (N_35280,N_23970,N_20053);
nor U35281 (N_35281,N_24371,N_23264);
nor U35282 (N_35282,N_23759,N_29935);
or U35283 (N_35283,N_25724,N_23661);
and U35284 (N_35284,N_27933,N_26848);
nor U35285 (N_35285,N_28640,N_24982);
nand U35286 (N_35286,N_20285,N_20158);
nand U35287 (N_35287,N_25033,N_22633);
and U35288 (N_35288,N_26004,N_29845);
or U35289 (N_35289,N_28799,N_27187);
and U35290 (N_35290,N_20492,N_24955);
and U35291 (N_35291,N_26090,N_26697);
nor U35292 (N_35292,N_20057,N_20788);
nand U35293 (N_35293,N_25284,N_21854);
or U35294 (N_35294,N_20469,N_20162);
nor U35295 (N_35295,N_27296,N_21917);
nor U35296 (N_35296,N_24940,N_23065);
nand U35297 (N_35297,N_27246,N_29726);
and U35298 (N_35298,N_22644,N_21651);
or U35299 (N_35299,N_29694,N_25330);
nand U35300 (N_35300,N_24530,N_22904);
or U35301 (N_35301,N_24670,N_26445);
nor U35302 (N_35302,N_28225,N_28729);
or U35303 (N_35303,N_22085,N_22332);
or U35304 (N_35304,N_24821,N_28970);
xor U35305 (N_35305,N_29821,N_22347);
nor U35306 (N_35306,N_24782,N_20323);
xnor U35307 (N_35307,N_23730,N_29813);
xnor U35308 (N_35308,N_21280,N_27175);
and U35309 (N_35309,N_21840,N_23890);
nand U35310 (N_35310,N_26275,N_20603);
nand U35311 (N_35311,N_29754,N_20206);
nand U35312 (N_35312,N_21078,N_25628);
and U35313 (N_35313,N_29726,N_29923);
nand U35314 (N_35314,N_28239,N_21212);
nor U35315 (N_35315,N_29265,N_20733);
xor U35316 (N_35316,N_28614,N_20876);
and U35317 (N_35317,N_23570,N_26813);
and U35318 (N_35318,N_21164,N_23603);
nand U35319 (N_35319,N_20918,N_27048);
or U35320 (N_35320,N_25194,N_24576);
and U35321 (N_35321,N_22080,N_27086);
nand U35322 (N_35322,N_20250,N_21079);
nand U35323 (N_35323,N_24861,N_22564);
nand U35324 (N_35324,N_29479,N_24942);
nand U35325 (N_35325,N_21800,N_27345);
and U35326 (N_35326,N_27657,N_27925);
nor U35327 (N_35327,N_26390,N_20292);
or U35328 (N_35328,N_20156,N_23161);
or U35329 (N_35329,N_22390,N_22379);
and U35330 (N_35330,N_24921,N_27302);
and U35331 (N_35331,N_24766,N_29245);
nand U35332 (N_35332,N_23075,N_29793);
and U35333 (N_35333,N_24273,N_20882);
and U35334 (N_35334,N_20890,N_26878);
nand U35335 (N_35335,N_28562,N_20610);
and U35336 (N_35336,N_22601,N_24325);
or U35337 (N_35337,N_28210,N_23096);
nor U35338 (N_35338,N_29567,N_23314);
or U35339 (N_35339,N_23393,N_21024);
xor U35340 (N_35340,N_20002,N_21785);
or U35341 (N_35341,N_28014,N_27346);
or U35342 (N_35342,N_26601,N_20113);
or U35343 (N_35343,N_26292,N_28934);
or U35344 (N_35344,N_29265,N_24724);
nor U35345 (N_35345,N_25532,N_23142);
nand U35346 (N_35346,N_25446,N_22057);
or U35347 (N_35347,N_20553,N_29467);
nand U35348 (N_35348,N_25883,N_28893);
nor U35349 (N_35349,N_23336,N_28272);
or U35350 (N_35350,N_29548,N_20734);
nor U35351 (N_35351,N_21913,N_29162);
nor U35352 (N_35352,N_25086,N_25137);
and U35353 (N_35353,N_24958,N_21666);
and U35354 (N_35354,N_22965,N_22771);
nand U35355 (N_35355,N_26152,N_23032);
nor U35356 (N_35356,N_20272,N_24910);
or U35357 (N_35357,N_26121,N_20501);
nand U35358 (N_35358,N_20778,N_28554);
or U35359 (N_35359,N_26360,N_21736);
and U35360 (N_35360,N_23766,N_23135);
or U35361 (N_35361,N_26947,N_28690);
xnor U35362 (N_35362,N_24324,N_20991);
and U35363 (N_35363,N_29369,N_29598);
nor U35364 (N_35364,N_22519,N_22905);
or U35365 (N_35365,N_21281,N_24237);
nor U35366 (N_35366,N_22685,N_25297);
or U35367 (N_35367,N_25370,N_23210);
nand U35368 (N_35368,N_22251,N_21742);
nor U35369 (N_35369,N_25843,N_27443);
nand U35370 (N_35370,N_27884,N_29543);
and U35371 (N_35371,N_22124,N_21323);
or U35372 (N_35372,N_27942,N_20376);
nand U35373 (N_35373,N_22027,N_25539);
xnor U35374 (N_35374,N_20111,N_29883);
or U35375 (N_35375,N_28355,N_28246);
nand U35376 (N_35376,N_27708,N_23322);
or U35377 (N_35377,N_24862,N_25359);
nor U35378 (N_35378,N_25964,N_25596);
or U35379 (N_35379,N_23258,N_27048);
or U35380 (N_35380,N_28432,N_21540);
and U35381 (N_35381,N_20294,N_26725);
nor U35382 (N_35382,N_27142,N_28689);
or U35383 (N_35383,N_29260,N_28334);
or U35384 (N_35384,N_26178,N_29764);
and U35385 (N_35385,N_22446,N_21013);
xnor U35386 (N_35386,N_24362,N_21552);
nor U35387 (N_35387,N_26143,N_24550);
or U35388 (N_35388,N_22425,N_22267);
nor U35389 (N_35389,N_27509,N_25923);
nor U35390 (N_35390,N_24686,N_28563);
and U35391 (N_35391,N_20759,N_22855);
nand U35392 (N_35392,N_21640,N_29612);
nand U35393 (N_35393,N_27589,N_20232);
nor U35394 (N_35394,N_29617,N_20171);
nor U35395 (N_35395,N_26414,N_29245);
or U35396 (N_35396,N_23257,N_20648);
or U35397 (N_35397,N_24517,N_23187);
or U35398 (N_35398,N_28572,N_21261);
nand U35399 (N_35399,N_24279,N_28629);
xnor U35400 (N_35400,N_24407,N_26523);
or U35401 (N_35401,N_20829,N_27651);
nor U35402 (N_35402,N_27630,N_21950);
and U35403 (N_35403,N_22147,N_21969);
xnor U35404 (N_35404,N_27182,N_24754);
nand U35405 (N_35405,N_25755,N_24335);
and U35406 (N_35406,N_25548,N_20015);
xnor U35407 (N_35407,N_28068,N_20795);
or U35408 (N_35408,N_24276,N_23256);
nand U35409 (N_35409,N_26614,N_27107);
or U35410 (N_35410,N_25304,N_20617);
or U35411 (N_35411,N_28392,N_23053);
and U35412 (N_35412,N_21598,N_27454);
nor U35413 (N_35413,N_27562,N_20152);
and U35414 (N_35414,N_21320,N_28833);
or U35415 (N_35415,N_25842,N_24708);
or U35416 (N_35416,N_21360,N_21990);
nor U35417 (N_35417,N_29279,N_26656);
nand U35418 (N_35418,N_25067,N_28267);
or U35419 (N_35419,N_24556,N_28114);
nor U35420 (N_35420,N_26649,N_22936);
and U35421 (N_35421,N_28298,N_27488);
or U35422 (N_35422,N_26541,N_20705);
or U35423 (N_35423,N_28583,N_25061);
nor U35424 (N_35424,N_27610,N_28915);
nand U35425 (N_35425,N_25303,N_20328);
xor U35426 (N_35426,N_26062,N_27969);
or U35427 (N_35427,N_21695,N_20134);
xor U35428 (N_35428,N_24257,N_21419);
nor U35429 (N_35429,N_24465,N_29464);
or U35430 (N_35430,N_27116,N_25448);
xor U35431 (N_35431,N_24505,N_22115);
or U35432 (N_35432,N_20580,N_20572);
or U35433 (N_35433,N_20671,N_27516);
and U35434 (N_35434,N_24185,N_21334);
nor U35435 (N_35435,N_21135,N_20241);
and U35436 (N_35436,N_26103,N_27744);
nor U35437 (N_35437,N_24224,N_20782);
or U35438 (N_35438,N_21781,N_25760);
nand U35439 (N_35439,N_27496,N_24291);
or U35440 (N_35440,N_22585,N_22789);
and U35441 (N_35441,N_29078,N_22594);
nor U35442 (N_35442,N_25240,N_27248);
nor U35443 (N_35443,N_28408,N_20473);
and U35444 (N_35444,N_27082,N_20592);
or U35445 (N_35445,N_26282,N_29658);
nor U35446 (N_35446,N_22564,N_29079);
nor U35447 (N_35447,N_27264,N_29078);
nor U35448 (N_35448,N_25982,N_20857);
nand U35449 (N_35449,N_20887,N_28519);
nor U35450 (N_35450,N_21246,N_26954);
xnor U35451 (N_35451,N_28136,N_25158);
nand U35452 (N_35452,N_21187,N_28814);
or U35453 (N_35453,N_28056,N_20975);
nand U35454 (N_35454,N_23180,N_23541);
nor U35455 (N_35455,N_23870,N_26073);
nand U35456 (N_35456,N_28911,N_23865);
xor U35457 (N_35457,N_24089,N_20055);
nand U35458 (N_35458,N_27838,N_23162);
or U35459 (N_35459,N_22500,N_27728);
or U35460 (N_35460,N_24017,N_27335);
and U35461 (N_35461,N_29776,N_28113);
or U35462 (N_35462,N_28246,N_26844);
nor U35463 (N_35463,N_29635,N_28422);
xor U35464 (N_35464,N_24464,N_28186);
nand U35465 (N_35465,N_22385,N_29148);
or U35466 (N_35466,N_20443,N_24170);
and U35467 (N_35467,N_27601,N_24896);
nor U35468 (N_35468,N_25971,N_23248);
nand U35469 (N_35469,N_21273,N_22041);
nor U35470 (N_35470,N_21426,N_22947);
nor U35471 (N_35471,N_29244,N_27552);
nand U35472 (N_35472,N_29824,N_20095);
nor U35473 (N_35473,N_26764,N_23890);
and U35474 (N_35474,N_29363,N_20825);
and U35475 (N_35475,N_21993,N_20697);
and U35476 (N_35476,N_21533,N_24686);
nor U35477 (N_35477,N_28591,N_27767);
nand U35478 (N_35478,N_22765,N_26807);
or U35479 (N_35479,N_22134,N_29635);
nor U35480 (N_35480,N_23517,N_26455);
or U35481 (N_35481,N_20689,N_20534);
and U35482 (N_35482,N_23970,N_22892);
nor U35483 (N_35483,N_29443,N_28964);
nand U35484 (N_35484,N_22341,N_26002);
nor U35485 (N_35485,N_28761,N_24980);
and U35486 (N_35486,N_20632,N_27165);
or U35487 (N_35487,N_23558,N_23274);
or U35488 (N_35488,N_29699,N_29466);
and U35489 (N_35489,N_20473,N_22252);
and U35490 (N_35490,N_26525,N_24098);
or U35491 (N_35491,N_22681,N_21642);
xnor U35492 (N_35492,N_21071,N_23594);
nor U35493 (N_35493,N_24174,N_22681);
nand U35494 (N_35494,N_20008,N_26196);
nand U35495 (N_35495,N_24370,N_27071);
and U35496 (N_35496,N_20622,N_24627);
nand U35497 (N_35497,N_21802,N_29962);
nor U35498 (N_35498,N_28436,N_23742);
xnor U35499 (N_35499,N_28326,N_29147);
nand U35500 (N_35500,N_25422,N_25552);
nand U35501 (N_35501,N_20667,N_21343);
xor U35502 (N_35502,N_27434,N_20809);
or U35503 (N_35503,N_26579,N_20542);
nand U35504 (N_35504,N_20668,N_20174);
and U35505 (N_35505,N_24437,N_20200);
nor U35506 (N_35506,N_26158,N_20684);
nand U35507 (N_35507,N_29872,N_25180);
or U35508 (N_35508,N_28084,N_25683);
nor U35509 (N_35509,N_27510,N_22512);
nor U35510 (N_35510,N_28612,N_21119);
or U35511 (N_35511,N_24698,N_27598);
nor U35512 (N_35512,N_20958,N_20530);
and U35513 (N_35513,N_24377,N_20785);
or U35514 (N_35514,N_22768,N_22113);
and U35515 (N_35515,N_29256,N_24457);
nand U35516 (N_35516,N_28246,N_22430);
or U35517 (N_35517,N_21228,N_26789);
and U35518 (N_35518,N_28787,N_24152);
nand U35519 (N_35519,N_24333,N_25586);
nor U35520 (N_35520,N_24813,N_21807);
and U35521 (N_35521,N_23590,N_28163);
xor U35522 (N_35522,N_20795,N_21258);
or U35523 (N_35523,N_26278,N_20120);
nor U35524 (N_35524,N_29352,N_23628);
nor U35525 (N_35525,N_24691,N_29965);
and U35526 (N_35526,N_29645,N_20800);
and U35527 (N_35527,N_27398,N_23331);
nand U35528 (N_35528,N_20291,N_22349);
or U35529 (N_35529,N_20969,N_23744);
or U35530 (N_35530,N_26511,N_28211);
and U35531 (N_35531,N_21207,N_20899);
nand U35532 (N_35532,N_21969,N_29040);
or U35533 (N_35533,N_29898,N_28749);
xor U35534 (N_35534,N_29235,N_24983);
and U35535 (N_35535,N_22451,N_28584);
or U35536 (N_35536,N_24542,N_26801);
xnor U35537 (N_35537,N_23380,N_21142);
and U35538 (N_35538,N_23228,N_23422);
or U35539 (N_35539,N_23200,N_24662);
or U35540 (N_35540,N_21661,N_25892);
nand U35541 (N_35541,N_26346,N_20117);
and U35542 (N_35542,N_29124,N_24960);
nand U35543 (N_35543,N_28603,N_24875);
or U35544 (N_35544,N_29666,N_23780);
nand U35545 (N_35545,N_24466,N_29219);
or U35546 (N_35546,N_21739,N_20769);
and U35547 (N_35547,N_29284,N_29720);
and U35548 (N_35548,N_29667,N_20887);
xor U35549 (N_35549,N_23150,N_24867);
and U35550 (N_35550,N_21439,N_24162);
nand U35551 (N_35551,N_24830,N_25118);
nor U35552 (N_35552,N_22058,N_27443);
nor U35553 (N_35553,N_22810,N_27045);
and U35554 (N_35554,N_25869,N_28606);
nand U35555 (N_35555,N_21284,N_27242);
xnor U35556 (N_35556,N_24308,N_20054);
nor U35557 (N_35557,N_21349,N_23522);
or U35558 (N_35558,N_21057,N_26760);
nand U35559 (N_35559,N_28400,N_27057);
and U35560 (N_35560,N_23128,N_20243);
xnor U35561 (N_35561,N_28402,N_29749);
nand U35562 (N_35562,N_24859,N_27546);
nor U35563 (N_35563,N_29705,N_20195);
nor U35564 (N_35564,N_20316,N_29431);
and U35565 (N_35565,N_23682,N_24612);
and U35566 (N_35566,N_26895,N_24893);
xnor U35567 (N_35567,N_20314,N_22305);
xnor U35568 (N_35568,N_24341,N_25395);
and U35569 (N_35569,N_22811,N_27885);
nor U35570 (N_35570,N_23220,N_23212);
nor U35571 (N_35571,N_23829,N_26328);
nand U35572 (N_35572,N_25444,N_26172);
or U35573 (N_35573,N_29138,N_23277);
or U35574 (N_35574,N_26579,N_26847);
nand U35575 (N_35575,N_22447,N_29522);
or U35576 (N_35576,N_29379,N_28772);
or U35577 (N_35577,N_24191,N_24474);
nor U35578 (N_35578,N_24310,N_26156);
or U35579 (N_35579,N_27695,N_24689);
nand U35580 (N_35580,N_23665,N_20302);
and U35581 (N_35581,N_20953,N_25373);
nor U35582 (N_35582,N_29319,N_27868);
and U35583 (N_35583,N_24283,N_20044);
nand U35584 (N_35584,N_23581,N_28759);
nand U35585 (N_35585,N_24917,N_20976);
nor U35586 (N_35586,N_22327,N_26339);
nand U35587 (N_35587,N_28768,N_28369);
or U35588 (N_35588,N_21783,N_28128);
or U35589 (N_35589,N_29454,N_24482);
and U35590 (N_35590,N_29232,N_21022);
or U35591 (N_35591,N_28113,N_24937);
and U35592 (N_35592,N_27630,N_21947);
or U35593 (N_35593,N_29695,N_24910);
nor U35594 (N_35594,N_24800,N_25998);
or U35595 (N_35595,N_22206,N_20070);
and U35596 (N_35596,N_29838,N_26966);
nor U35597 (N_35597,N_28564,N_23616);
nor U35598 (N_35598,N_27373,N_21825);
xor U35599 (N_35599,N_20609,N_29769);
nor U35600 (N_35600,N_28673,N_23762);
nand U35601 (N_35601,N_29212,N_27546);
or U35602 (N_35602,N_22802,N_29738);
nor U35603 (N_35603,N_24794,N_27643);
or U35604 (N_35604,N_28696,N_26998);
or U35605 (N_35605,N_21891,N_27744);
or U35606 (N_35606,N_23603,N_26759);
nor U35607 (N_35607,N_26410,N_29304);
nand U35608 (N_35608,N_20538,N_26900);
or U35609 (N_35609,N_24407,N_24360);
and U35610 (N_35610,N_27279,N_24531);
nand U35611 (N_35611,N_25938,N_29053);
and U35612 (N_35612,N_27881,N_24800);
nor U35613 (N_35613,N_22333,N_26574);
nor U35614 (N_35614,N_22951,N_23518);
xnor U35615 (N_35615,N_27292,N_21946);
and U35616 (N_35616,N_23130,N_23596);
nor U35617 (N_35617,N_28150,N_26504);
or U35618 (N_35618,N_28767,N_20209);
nor U35619 (N_35619,N_22548,N_24861);
or U35620 (N_35620,N_23717,N_26645);
nand U35621 (N_35621,N_25821,N_28023);
nor U35622 (N_35622,N_25935,N_23097);
nor U35623 (N_35623,N_26086,N_21067);
nand U35624 (N_35624,N_22181,N_29231);
and U35625 (N_35625,N_20562,N_21633);
nand U35626 (N_35626,N_23966,N_20639);
and U35627 (N_35627,N_23087,N_22932);
and U35628 (N_35628,N_29623,N_29905);
and U35629 (N_35629,N_29153,N_29235);
or U35630 (N_35630,N_28591,N_21634);
xnor U35631 (N_35631,N_26752,N_29854);
or U35632 (N_35632,N_23674,N_28870);
nand U35633 (N_35633,N_20573,N_29724);
nor U35634 (N_35634,N_25032,N_27775);
nand U35635 (N_35635,N_20887,N_24414);
nand U35636 (N_35636,N_26127,N_24746);
and U35637 (N_35637,N_28996,N_28846);
and U35638 (N_35638,N_22231,N_28333);
nand U35639 (N_35639,N_28055,N_28913);
nor U35640 (N_35640,N_24338,N_28105);
and U35641 (N_35641,N_20207,N_23647);
nor U35642 (N_35642,N_27255,N_22960);
and U35643 (N_35643,N_21923,N_22631);
nor U35644 (N_35644,N_24664,N_24148);
nand U35645 (N_35645,N_29700,N_21265);
xor U35646 (N_35646,N_23133,N_27930);
nor U35647 (N_35647,N_20133,N_27103);
and U35648 (N_35648,N_22194,N_21756);
or U35649 (N_35649,N_26109,N_29284);
xor U35650 (N_35650,N_20424,N_29228);
nand U35651 (N_35651,N_29349,N_22904);
and U35652 (N_35652,N_20970,N_26783);
and U35653 (N_35653,N_20236,N_25535);
nand U35654 (N_35654,N_22379,N_24872);
nor U35655 (N_35655,N_20967,N_29298);
nand U35656 (N_35656,N_26788,N_20788);
nor U35657 (N_35657,N_21854,N_27379);
or U35658 (N_35658,N_22329,N_24995);
or U35659 (N_35659,N_20044,N_20223);
xnor U35660 (N_35660,N_20772,N_26316);
and U35661 (N_35661,N_25739,N_26027);
and U35662 (N_35662,N_23220,N_23837);
and U35663 (N_35663,N_21167,N_24967);
or U35664 (N_35664,N_22343,N_23403);
and U35665 (N_35665,N_24480,N_27330);
and U35666 (N_35666,N_25528,N_23076);
nor U35667 (N_35667,N_21375,N_20900);
xor U35668 (N_35668,N_26144,N_26615);
nand U35669 (N_35669,N_22384,N_26501);
nor U35670 (N_35670,N_27273,N_27887);
or U35671 (N_35671,N_27402,N_29667);
nor U35672 (N_35672,N_23704,N_29533);
nor U35673 (N_35673,N_21954,N_23277);
or U35674 (N_35674,N_27925,N_29343);
nand U35675 (N_35675,N_24501,N_27737);
nor U35676 (N_35676,N_23818,N_22377);
nor U35677 (N_35677,N_23490,N_25462);
nor U35678 (N_35678,N_25298,N_24820);
nand U35679 (N_35679,N_21040,N_29317);
or U35680 (N_35680,N_29968,N_26837);
and U35681 (N_35681,N_28738,N_22718);
and U35682 (N_35682,N_25806,N_24764);
nand U35683 (N_35683,N_26821,N_25627);
nand U35684 (N_35684,N_25766,N_26862);
nor U35685 (N_35685,N_29039,N_27506);
and U35686 (N_35686,N_23476,N_29390);
xor U35687 (N_35687,N_23709,N_25224);
nor U35688 (N_35688,N_20318,N_26580);
xor U35689 (N_35689,N_25613,N_20420);
nand U35690 (N_35690,N_20602,N_27160);
xnor U35691 (N_35691,N_25073,N_24493);
and U35692 (N_35692,N_23239,N_22628);
and U35693 (N_35693,N_25990,N_26424);
nand U35694 (N_35694,N_25013,N_24586);
or U35695 (N_35695,N_28339,N_24020);
nand U35696 (N_35696,N_24554,N_24814);
or U35697 (N_35697,N_29551,N_25523);
or U35698 (N_35698,N_28325,N_21017);
nor U35699 (N_35699,N_22979,N_20676);
and U35700 (N_35700,N_27383,N_29307);
and U35701 (N_35701,N_24890,N_23524);
nor U35702 (N_35702,N_26331,N_20778);
or U35703 (N_35703,N_23110,N_28920);
nand U35704 (N_35704,N_28257,N_22758);
nand U35705 (N_35705,N_20799,N_25308);
or U35706 (N_35706,N_24441,N_27771);
and U35707 (N_35707,N_27341,N_27856);
or U35708 (N_35708,N_22168,N_21158);
xnor U35709 (N_35709,N_29222,N_27928);
or U35710 (N_35710,N_20748,N_21962);
nor U35711 (N_35711,N_28460,N_22932);
nand U35712 (N_35712,N_26582,N_26509);
nand U35713 (N_35713,N_25539,N_29355);
xor U35714 (N_35714,N_26604,N_25061);
or U35715 (N_35715,N_24389,N_26951);
and U35716 (N_35716,N_26113,N_25589);
nand U35717 (N_35717,N_20996,N_21262);
nand U35718 (N_35718,N_22937,N_27612);
and U35719 (N_35719,N_28306,N_28799);
nand U35720 (N_35720,N_24345,N_25801);
nand U35721 (N_35721,N_27782,N_29864);
nor U35722 (N_35722,N_29050,N_26884);
nand U35723 (N_35723,N_28936,N_24767);
nor U35724 (N_35724,N_24326,N_22680);
nand U35725 (N_35725,N_23465,N_25679);
xnor U35726 (N_35726,N_29130,N_21407);
xnor U35727 (N_35727,N_28451,N_28537);
nor U35728 (N_35728,N_28417,N_27475);
nand U35729 (N_35729,N_26820,N_27924);
or U35730 (N_35730,N_21260,N_25973);
nor U35731 (N_35731,N_28747,N_22255);
and U35732 (N_35732,N_27166,N_20363);
or U35733 (N_35733,N_29480,N_25695);
and U35734 (N_35734,N_26645,N_29124);
nor U35735 (N_35735,N_22748,N_22068);
nand U35736 (N_35736,N_22929,N_27668);
or U35737 (N_35737,N_26437,N_20537);
or U35738 (N_35738,N_29650,N_24700);
and U35739 (N_35739,N_27722,N_26927);
nand U35740 (N_35740,N_21705,N_28068);
nor U35741 (N_35741,N_23890,N_26610);
nand U35742 (N_35742,N_21412,N_22324);
xor U35743 (N_35743,N_23238,N_28388);
nor U35744 (N_35744,N_22386,N_20446);
and U35745 (N_35745,N_26729,N_28392);
nor U35746 (N_35746,N_27845,N_22987);
and U35747 (N_35747,N_25351,N_23559);
and U35748 (N_35748,N_27957,N_23567);
nand U35749 (N_35749,N_28723,N_25080);
or U35750 (N_35750,N_26066,N_25373);
nor U35751 (N_35751,N_21599,N_26637);
xor U35752 (N_35752,N_21642,N_28264);
and U35753 (N_35753,N_28228,N_23090);
nor U35754 (N_35754,N_26562,N_27467);
or U35755 (N_35755,N_22371,N_20808);
and U35756 (N_35756,N_27582,N_20733);
nor U35757 (N_35757,N_24184,N_22269);
nor U35758 (N_35758,N_28298,N_24152);
nor U35759 (N_35759,N_24962,N_25223);
nand U35760 (N_35760,N_26246,N_26929);
or U35761 (N_35761,N_27467,N_29977);
nand U35762 (N_35762,N_26293,N_24457);
and U35763 (N_35763,N_20300,N_28075);
xor U35764 (N_35764,N_26947,N_22894);
and U35765 (N_35765,N_23578,N_29624);
or U35766 (N_35766,N_29936,N_28958);
nand U35767 (N_35767,N_27240,N_21762);
or U35768 (N_35768,N_29693,N_21238);
or U35769 (N_35769,N_28435,N_20189);
or U35770 (N_35770,N_22445,N_20458);
nand U35771 (N_35771,N_29643,N_27206);
xor U35772 (N_35772,N_28064,N_25145);
nor U35773 (N_35773,N_20878,N_26790);
nor U35774 (N_35774,N_20419,N_21459);
or U35775 (N_35775,N_25806,N_22191);
xor U35776 (N_35776,N_25901,N_21296);
or U35777 (N_35777,N_21116,N_22253);
nand U35778 (N_35778,N_24461,N_20844);
nor U35779 (N_35779,N_28410,N_28111);
and U35780 (N_35780,N_25642,N_26914);
xor U35781 (N_35781,N_29487,N_20806);
nand U35782 (N_35782,N_25482,N_24631);
nand U35783 (N_35783,N_21579,N_21331);
nand U35784 (N_35784,N_29990,N_26592);
and U35785 (N_35785,N_24826,N_29399);
or U35786 (N_35786,N_26937,N_28531);
nor U35787 (N_35787,N_21576,N_23335);
nor U35788 (N_35788,N_26603,N_22810);
and U35789 (N_35789,N_24036,N_21899);
xor U35790 (N_35790,N_27750,N_21110);
xor U35791 (N_35791,N_28708,N_24856);
and U35792 (N_35792,N_23617,N_22980);
or U35793 (N_35793,N_26598,N_24628);
or U35794 (N_35794,N_24322,N_20547);
nor U35795 (N_35795,N_24552,N_27058);
xor U35796 (N_35796,N_26581,N_24683);
or U35797 (N_35797,N_25866,N_20237);
nor U35798 (N_35798,N_26998,N_25380);
xor U35799 (N_35799,N_28185,N_22113);
and U35800 (N_35800,N_26651,N_22770);
xor U35801 (N_35801,N_24579,N_21261);
and U35802 (N_35802,N_27522,N_28146);
nand U35803 (N_35803,N_24049,N_26511);
nand U35804 (N_35804,N_24592,N_21300);
or U35805 (N_35805,N_20016,N_25878);
or U35806 (N_35806,N_23657,N_28115);
and U35807 (N_35807,N_23124,N_29687);
nor U35808 (N_35808,N_28556,N_20708);
nor U35809 (N_35809,N_28722,N_28416);
nand U35810 (N_35810,N_25714,N_28297);
nor U35811 (N_35811,N_25951,N_26771);
and U35812 (N_35812,N_22806,N_27921);
nor U35813 (N_35813,N_26776,N_20244);
and U35814 (N_35814,N_23435,N_23857);
xnor U35815 (N_35815,N_20302,N_25033);
and U35816 (N_35816,N_28213,N_29793);
or U35817 (N_35817,N_29370,N_26649);
and U35818 (N_35818,N_21210,N_22221);
or U35819 (N_35819,N_27279,N_25310);
nand U35820 (N_35820,N_29327,N_23673);
nand U35821 (N_35821,N_21288,N_25626);
and U35822 (N_35822,N_27616,N_29692);
nand U35823 (N_35823,N_25260,N_21731);
nand U35824 (N_35824,N_29962,N_29486);
nor U35825 (N_35825,N_27072,N_21104);
or U35826 (N_35826,N_29942,N_27338);
nand U35827 (N_35827,N_29499,N_24435);
nand U35828 (N_35828,N_25393,N_24988);
and U35829 (N_35829,N_22972,N_20127);
xnor U35830 (N_35830,N_25888,N_28051);
and U35831 (N_35831,N_22286,N_28157);
nand U35832 (N_35832,N_29321,N_25767);
or U35833 (N_35833,N_20255,N_27857);
nand U35834 (N_35834,N_21661,N_28321);
and U35835 (N_35835,N_28963,N_23905);
xnor U35836 (N_35836,N_25963,N_24167);
or U35837 (N_35837,N_27750,N_24924);
nor U35838 (N_35838,N_28711,N_24411);
nor U35839 (N_35839,N_26708,N_26368);
nand U35840 (N_35840,N_27020,N_21973);
nand U35841 (N_35841,N_21391,N_23878);
nor U35842 (N_35842,N_28854,N_20049);
nand U35843 (N_35843,N_23499,N_20533);
nand U35844 (N_35844,N_25956,N_24103);
nand U35845 (N_35845,N_27307,N_27977);
and U35846 (N_35846,N_20491,N_29285);
nand U35847 (N_35847,N_26092,N_20356);
and U35848 (N_35848,N_21946,N_27272);
and U35849 (N_35849,N_24971,N_26280);
or U35850 (N_35850,N_20213,N_23075);
or U35851 (N_35851,N_21081,N_21125);
and U35852 (N_35852,N_28098,N_22808);
or U35853 (N_35853,N_27792,N_25802);
or U35854 (N_35854,N_23288,N_29589);
and U35855 (N_35855,N_29898,N_29985);
and U35856 (N_35856,N_29775,N_28246);
xnor U35857 (N_35857,N_28688,N_21547);
nand U35858 (N_35858,N_25106,N_26993);
nor U35859 (N_35859,N_20554,N_23289);
and U35860 (N_35860,N_29526,N_21004);
nand U35861 (N_35861,N_25556,N_20896);
nor U35862 (N_35862,N_25991,N_29859);
nor U35863 (N_35863,N_28894,N_27597);
and U35864 (N_35864,N_24758,N_23423);
and U35865 (N_35865,N_23547,N_22292);
and U35866 (N_35866,N_20847,N_22651);
and U35867 (N_35867,N_22906,N_21916);
nand U35868 (N_35868,N_25993,N_23387);
nor U35869 (N_35869,N_25508,N_28205);
or U35870 (N_35870,N_28904,N_24940);
and U35871 (N_35871,N_24064,N_29288);
nand U35872 (N_35872,N_20202,N_25402);
xnor U35873 (N_35873,N_26038,N_20109);
or U35874 (N_35874,N_24605,N_24683);
and U35875 (N_35875,N_27137,N_21046);
nand U35876 (N_35876,N_27870,N_27152);
and U35877 (N_35877,N_26322,N_24143);
xnor U35878 (N_35878,N_28339,N_22264);
nand U35879 (N_35879,N_27217,N_22037);
or U35880 (N_35880,N_22639,N_23720);
nor U35881 (N_35881,N_24335,N_27655);
and U35882 (N_35882,N_25409,N_25472);
or U35883 (N_35883,N_26843,N_22473);
and U35884 (N_35884,N_27899,N_28645);
or U35885 (N_35885,N_23194,N_25760);
nand U35886 (N_35886,N_28479,N_26460);
nor U35887 (N_35887,N_21217,N_29800);
nor U35888 (N_35888,N_21199,N_29191);
and U35889 (N_35889,N_20867,N_28257);
and U35890 (N_35890,N_22484,N_26037);
nand U35891 (N_35891,N_25248,N_25436);
nor U35892 (N_35892,N_26695,N_22830);
nor U35893 (N_35893,N_22152,N_21731);
and U35894 (N_35894,N_25399,N_25163);
and U35895 (N_35895,N_26994,N_29143);
or U35896 (N_35896,N_29068,N_29926);
or U35897 (N_35897,N_29471,N_20909);
xnor U35898 (N_35898,N_22299,N_24985);
nand U35899 (N_35899,N_26851,N_21374);
or U35900 (N_35900,N_29073,N_24904);
nand U35901 (N_35901,N_26582,N_24449);
or U35902 (N_35902,N_27285,N_26992);
xor U35903 (N_35903,N_20114,N_28006);
nor U35904 (N_35904,N_22298,N_28814);
xnor U35905 (N_35905,N_25145,N_21371);
xor U35906 (N_35906,N_25672,N_20810);
or U35907 (N_35907,N_21627,N_24493);
nor U35908 (N_35908,N_27036,N_27648);
nand U35909 (N_35909,N_21447,N_22035);
nor U35910 (N_35910,N_29064,N_21117);
or U35911 (N_35911,N_20588,N_29624);
and U35912 (N_35912,N_28387,N_24223);
xor U35913 (N_35913,N_28186,N_27592);
nor U35914 (N_35914,N_28158,N_25762);
and U35915 (N_35915,N_26176,N_27959);
nor U35916 (N_35916,N_21483,N_23521);
or U35917 (N_35917,N_24738,N_22231);
or U35918 (N_35918,N_24056,N_27606);
nand U35919 (N_35919,N_22678,N_26595);
nand U35920 (N_35920,N_27439,N_29356);
or U35921 (N_35921,N_28316,N_27488);
or U35922 (N_35922,N_21331,N_20776);
or U35923 (N_35923,N_28745,N_26324);
nor U35924 (N_35924,N_27857,N_24403);
nand U35925 (N_35925,N_29357,N_21842);
nand U35926 (N_35926,N_26201,N_22467);
or U35927 (N_35927,N_29593,N_28142);
or U35928 (N_35928,N_26085,N_27902);
nor U35929 (N_35929,N_29872,N_24141);
nor U35930 (N_35930,N_24251,N_22141);
or U35931 (N_35931,N_25092,N_20676);
xnor U35932 (N_35932,N_21971,N_26308);
nor U35933 (N_35933,N_22422,N_21096);
nor U35934 (N_35934,N_20080,N_28855);
or U35935 (N_35935,N_26165,N_22809);
nand U35936 (N_35936,N_23277,N_27474);
or U35937 (N_35937,N_21623,N_23223);
and U35938 (N_35938,N_20105,N_24979);
nor U35939 (N_35939,N_20707,N_22632);
nand U35940 (N_35940,N_22012,N_20204);
or U35941 (N_35941,N_21017,N_23805);
or U35942 (N_35942,N_24987,N_28820);
or U35943 (N_35943,N_23741,N_24072);
or U35944 (N_35944,N_29621,N_26937);
or U35945 (N_35945,N_22574,N_25643);
nor U35946 (N_35946,N_25506,N_23839);
nand U35947 (N_35947,N_21324,N_27097);
and U35948 (N_35948,N_27252,N_26447);
or U35949 (N_35949,N_24275,N_22061);
xor U35950 (N_35950,N_22852,N_29930);
and U35951 (N_35951,N_20873,N_24010);
or U35952 (N_35952,N_28560,N_24373);
and U35953 (N_35953,N_22717,N_21373);
nand U35954 (N_35954,N_28986,N_26345);
xor U35955 (N_35955,N_24458,N_22917);
nand U35956 (N_35956,N_25628,N_20731);
nand U35957 (N_35957,N_29798,N_24458);
or U35958 (N_35958,N_27543,N_21824);
nand U35959 (N_35959,N_20813,N_26153);
nand U35960 (N_35960,N_25170,N_28916);
or U35961 (N_35961,N_27847,N_29723);
nand U35962 (N_35962,N_26770,N_26195);
nor U35963 (N_35963,N_23770,N_22267);
nor U35964 (N_35964,N_28787,N_24348);
or U35965 (N_35965,N_26124,N_25421);
nand U35966 (N_35966,N_26812,N_27646);
nand U35967 (N_35967,N_23105,N_20651);
nand U35968 (N_35968,N_23367,N_29039);
nand U35969 (N_35969,N_28995,N_26182);
nand U35970 (N_35970,N_26004,N_21050);
or U35971 (N_35971,N_29996,N_22261);
nand U35972 (N_35972,N_23638,N_22893);
or U35973 (N_35973,N_21444,N_24300);
nor U35974 (N_35974,N_26370,N_23238);
nand U35975 (N_35975,N_27575,N_21835);
or U35976 (N_35976,N_25096,N_22869);
or U35977 (N_35977,N_28857,N_27816);
or U35978 (N_35978,N_28747,N_28042);
nand U35979 (N_35979,N_24806,N_28851);
nand U35980 (N_35980,N_25585,N_20118);
nand U35981 (N_35981,N_27805,N_21524);
or U35982 (N_35982,N_25488,N_29381);
or U35983 (N_35983,N_22600,N_29593);
nor U35984 (N_35984,N_20358,N_26875);
nor U35985 (N_35985,N_29294,N_22838);
or U35986 (N_35986,N_24391,N_27204);
and U35987 (N_35987,N_20138,N_21130);
nor U35988 (N_35988,N_22384,N_23884);
or U35989 (N_35989,N_27286,N_28887);
nand U35990 (N_35990,N_26185,N_28078);
and U35991 (N_35991,N_20478,N_23184);
or U35992 (N_35992,N_24858,N_21171);
nor U35993 (N_35993,N_28756,N_24505);
xnor U35994 (N_35994,N_20411,N_27625);
or U35995 (N_35995,N_20793,N_22038);
xor U35996 (N_35996,N_28294,N_27805);
and U35997 (N_35997,N_26008,N_20637);
or U35998 (N_35998,N_20272,N_28848);
xnor U35999 (N_35999,N_23235,N_26490);
and U36000 (N_36000,N_28575,N_29568);
nand U36001 (N_36001,N_25277,N_28054);
nor U36002 (N_36002,N_28765,N_22863);
nand U36003 (N_36003,N_26464,N_29963);
nand U36004 (N_36004,N_20781,N_20363);
and U36005 (N_36005,N_28744,N_20111);
or U36006 (N_36006,N_26709,N_22189);
or U36007 (N_36007,N_27679,N_22906);
xnor U36008 (N_36008,N_20862,N_27231);
xnor U36009 (N_36009,N_20709,N_24880);
nor U36010 (N_36010,N_20598,N_21478);
or U36011 (N_36011,N_21584,N_27290);
and U36012 (N_36012,N_20078,N_27618);
xor U36013 (N_36013,N_29202,N_20463);
or U36014 (N_36014,N_22970,N_29239);
xor U36015 (N_36015,N_21568,N_25276);
nand U36016 (N_36016,N_20439,N_21268);
nand U36017 (N_36017,N_20501,N_22324);
nand U36018 (N_36018,N_21767,N_27375);
nor U36019 (N_36019,N_21562,N_25655);
nand U36020 (N_36020,N_22469,N_21854);
and U36021 (N_36021,N_29199,N_20031);
nor U36022 (N_36022,N_28716,N_24753);
nor U36023 (N_36023,N_26012,N_24414);
nand U36024 (N_36024,N_22665,N_24464);
nor U36025 (N_36025,N_28565,N_24551);
nand U36026 (N_36026,N_28328,N_21219);
nand U36027 (N_36027,N_27672,N_21467);
nand U36028 (N_36028,N_20874,N_28724);
xor U36029 (N_36029,N_26053,N_23801);
nor U36030 (N_36030,N_23933,N_22966);
or U36031 (N_36031,N_21934,N_23480);
nor U36032 (N_36032,N_24626,N_22376);
or U36033 (N_36033,N_22829,N_24579);
and U36034 (N_36034,N_25660,N_28176);
nor U36035 (N_36035,N_26617,N_20546);
or U36036 (N_36036,N_25223,N_20560);
nand U36037 (N_36037,N_27211,N_20573);
xor U36038 (N_36038,N_29553,N_25562);
nor U36039 (N_36039,N_28722,N_28605);
nand U36040 (N_36040,N_27459,N_20070);
or U36041 (N_36041,N_26782,N_24101);
or U36042 (N_36042,N_22304,N_29381);
nand U36043 (N_36043,N_27279,N_28407);
nand U36044 (N_36044,N_27685,N_25397);
or U36045 (N_36045,N_23229,N_22888);
nand U36046 (N_36046,N_26572,N_20833);
nor U36047 (N_36047,N_22991,N_26774);
and U36048 (N_36048,N_27296,N_20155);
nand U36049 (N_36049,N_27002,N_26395);
or U36050 (N_36050,N_26409,N_20344);
and U36051 (N_36051,N_23648,N_23542);
nand U36052 (N_36052,N_29677,N_27026);
or U36053 (N_36053,N_29262,N_27975);
nand U36054 (N_36054,N_24576,N_25736);
nor U36055 (N_36055,N_24391,N_27501);
or U36056 (N_36056,N_26887,N_21441);
xor U36057 (N_36057,N_28857,N_20017);
or U36058 (N_36058,N_27373,N_29160);
nor U36059 (N_36059,N_28730,N_23815);
nor U36060 (N_36060,N_22288,N_29390);
or U36061 (N_36061,N_23284,N_24355);
nor U36062 (N_36062,N_26775,N_21612);
nor U36063 (N_36063,N_25252,N_27730);
xor U36064 (N_36064,N_29877,N_22471);
nand U36065 (N_36065,N_22623,N_26145);
nor U36066 (N_36066,N_22695,N_23521);
or U36067 (N_36067,N_27653,N_27730);
or U36068 (N_36068,N_26479,N_21967);
or U36069 (N_36069,N_28136,N_24908);
nand U36070 (N_36070,N_23239,N_20755);
nand U36071 (N_36071,N_21706,N_23697);
nand U36072 (N_36072,N_24394,N_24910);
nor U36073 (N_36073,N_29415,N_25461);
or U36074 (N_36074,N_26313,N_25144);
and U36075 (N_36075,N_23793,N_21907);
and U36076 (N_36076,N_21392,N_25550);
nor U36077 (N_36077,N_23491,N_21955);
and U36078 (N_36078,N_29263,N_21141);
and U36079 (N_36079,N_25040,N_23346);
and U36080 (N_36080,N_21507,N_25832);
and U36081 (N_36081,N_20991,N_24804);
or U36082 (N_36082,N_22348,N_25887);
nand U36083 (N_36083,N_26900,N_24455);
and U36084 (N_36084,N_28717,N_28415);
nand U36085 (N_36085,N_28359,N_20087);
nand U36086 (N_36086,N_20362,N_22031);
nor U36087 (N_36087,N_24397,N_23410);
nand U36088 (N_36088,N_24035,N_24276);
or U36089 (N_36089,N_20952,N_28442);
and U36090 (N_36090,N_27055,N_21740);
xor U36091 (N_36091,N_20285,N_27799);
and U36092 (N_36092,N_26713,N_22421);
or U36093 (N_36093,N_24693,N_20202);
or U36094 (N_36094,N_28806,N_21251);
nor U36095 (N_36095,N_24598,N_22677);
nand U36096 (N_36096,N_25287,N_26094);
nand U36097 (N_36097,N_24429,N_29411);
nand U36098 (N_36098,N_22402,N_25485);
and U36099 (N_36099,N_26458,N_26462);
nor U36100 (N_36100,N_28649,N_27567);
xor U36101 (N_36101,N_29841,N_28420);
or U36102 (N_36102,N_20032,N_22838);
nand U36103 (N_36103,N_20911,N_24969);
nor U36104 (N_36104,N_22791,N_21854);
and U36105 (N_36105,N_23618,N_21533);
nand U36106 (N_36106,N_21385,N_27509);
and U36107 (N_36107,N_29049,N_27289);
or U36108 (N_36108,N_24968,N_23249);
or U36109 (N_36109,N_29207,N_28185);
nand U36110 (N_36110,N_24052,N_23466);
nand U36111 (N_36111,N_26321,N_27489);
nor U36112 (N_36112,N_20990,N_21653);
or U36113 (N_36113,N_21887,N_22019);
nor U36114 (N_36114,N_29180,N_23908);
or U36115 (N_36115,N_27611,N_29152);
or U36116 (N_36116,N_20636,N_28745);
xnor U36117 (N_36117,N_25219,N_23510);
or U36118 (N_36118,N_23702,N_26112);
or U36119 (N_36119,N_25168,N_25033);
xnor U36120 (N_36120,N_24476,N_21694);
nand U36121 (N_36121,N_21593,N_22233);
xor U36122 (N_36122,N_21836,N_26029);
xor U36123 (N_36123,N_29532,N_23691);
and U36124 (N_36124,N_20425,N_26336);
nor U36125 (N_36125,N_24539,N_29444);
and U36126 (N_36126,N_20115,N_21096);
nor U36127 (N_36127,N_28433,N_22078);
or U36128 (N_36128,N_29212,N_29217);
nor U36129 (N_36129,N_21009,N_26690);
nor U36130 (N_36130,N_28765,N_22049);
and U36131 (N_36131,N_29617,N_21512);
and U36132 (N_36132,N_20840,N_29395);
and U36133 (N_36133,N_23084,N_24129);
or U36134 (N_36134,N_28289,N_24065);
nor U36135 (N_36135,N_24603,N_29763);
or U36136 (N_36136,N_28655,N_29116);
nand U36137 (N_36137,N_21239,N_29183);
and U36138 (N_36138,N_27335,N_22008);
nand U36139 (N_36139,N_24825,N_23132);
and U36140 (N_36140,N_27757,N_26579);
nand U36141 (N_36141,N_21523,N_24784);
nor U36142 (N_36142,N_26343,N_23880);
nand U36143 (N_36143,N_20637,N_27165);
nand U36144 (N_36144,N_22185,N_21352);
nand U36145 (N_36145,N_24375,N_25244);
nand U36146 (N_36146,N_21581,N_22759);
nor U36147 (N_36147,N_23583,N_24295);
nor U36148 (N_36148,N_28261,N_26754);
nand U36149 (N_36149,N_20872,N_26982);
xor U36150 (N_36150,N_20656,N_27851);
or U36151 (N_36151,N_28188,N_23147);
nor U36152 (N_36152,N_28627,N_28040);
nand U36153 (N_36153,N_27333,N_28352);
and U36154 (N_36154,N_21402,N_20410);
nand U36155 (N_36155,N_24523,N_20831);
or U36156 (N_36156,N_20149,N_20987);
xnor U36157 (N_36157,N_24535,N_29472);
nand U36158 (N_36158,N_23259,N_20632);
nand U36159 (N_36159,N_29916,N_27169);
and U36160 (N_36160,N_22754,N_21054);
or U36161 (N_36161,N_25851,N_22418);
nand U36162 (N_36162,N_29265,N_26234);
xnor U36163 (N_36163,N_24737,N_22837);
nand U36164 (N_36164,N_21705,N_27856);
nand U36165 (N_36165,N_24711,N_27268);
xnor U36166 (N_36166,N_21060,N_27234);
xor U36167 (N_36167,N_20624,N_20887);
and U36168 (N_36168,N_25165,N_22879);
nor U36169 (N_36169,N_25257,N_25402);
nand U36170 (N_36170,N_21753,N_20548);
and U36171 (N_36171,N_28556,N_23451);
xor U36172 (N_36172,N_29629,N_22340);
and U36173 (N_36173,N_27981,N_23932);
or U36174 (N_36174,N_21902,N_29334);
and U36175 (N_36175,N_23373,N_20110);
nand U36176 (N_36176,N_23411,N_28988);
and U36177 (N_36177,N_21838,N_28336);
or U36178 (N_36178,N_25784,N_27391);
and U36179 (N_36179,N_21857,N_22586);
or U36180 (N_36180,N_29255,N_20904);
nor U36181 (N_36181,N_29203,N_23986);
nand U36182 (N_36182,N_20157,N_29426);
or U36183 (N_36183,N_25320,N_27524);
xnor U36184 (N_36184,N_21232,N_21698);
and U36185 (N_36185,N_27142,N_23011);
and U36186 (N_36186,N_28667,N_20814);
and U36187 (N_36187,N_24571,N_22679);
and U36188 (N_36188,N_28451,N_29876);
and U36189 (N_36189,N_26900,N_21762);
or U36190 (N_36190,N_20041,N_24122);
and U36191 (N_36191,N_22951,N_21728);
or U36192 (N_36192,N_24419,N_27936);
nor U36193 (N_36193,N_22820,N_23134);
nand U36194 (N_36194,N_25460,N_21085);
xnor U36195 (N_36195,N_24161,N_24178);
or U36196 (N_36196,N_20444,N_22825);
and U36197 (N_36197,N_21828,N_22093);
or U36198 (N_36198,N_25177,N_27536);
or U36199 (N_36199,N_27739,N_26951);
and U36200 (N_36200,N_24128,N_29791);
xor U36201 (N_36201,N_25543,N_21215);
or U36202 (N_36202,N_20709,N_23949);
xnor U36203 (N_36203,N_27672,N_21469);
and U36204 (N_36204,N_29846,N_24398);
nor U36205 (N_36205,N_29214,N_24139);
or U36206 (N_36206,N_22144,N_22804);
and U36207 (N_36207,N_21557,N_23771);
nor U36208 (N_36208,N_23363,N_27957);
or U36209 (N_36209,N_29658,N_28281);
xor U36210 (N_36210,N_20432,N_26967);
nor U36211 (N_36211,N_28315,N_27060);
and U36212 (N_36212,N_26228,N_22899);
nand U36213 (N_36213,N_21595,N_22804);
and U36214 (N_36214,N_22754,N_21929);
and U36215 (N_36215,N_22176,N_20429);
nor U36216 (N_36216,N_27691,N_25203);
and U36217 (N_36217,N_22150,N_24091);
xnor U36218 (N_36218,N_24764,N_23710);
and U36219 (N_36219,N_29991,N_26304);
nand U36220 (N_36220,N_21400,N_23900);
nand U36221 (N_36221,N_23652,N_25886);
nor U36222 (N_36222,N_20804,N_24344);
xnor U36223 (N_36223,N_22856,N_27364);
nand U36224 (N_36224,N_28746,N_20552);
nand U36225 (N_36225,N_20388,N_24567);
and U36226 (N_36226,N_29419,N_27305);
or U36227 (N_36227,N_27610,N_22820);
nand U36228 (N_36228,N_21859,N_21672);
and U36229 (N_36229,N_27919,N_21574);
and U36230 (N_36230,N_24167,N_22554);
and U36231 (N_36231,N_24577,N_25588);
nor U36232 (N_36232,N_29481,N_29536);
nand U36233 (N_36233,N_21102,N_25117);
and U36234 (N_36234,N_25562,N_22162);
nor U36235 (N_36235,N_22736,N_26371);
nor U36236 (N_36236,N_22282,N_24248);
or U36237 (N_36237,N_29209,N_26561);
and U36238 (N_36238,N_26775,N_25811);
nor U36239 (N_36239,N_20001,N_26618);
or U36240 (N_36240,N_27569,N_20347);
and U36241 (N_36241,N_25171,N_22311);
or U36242 (N_36242,N_24240,N_21451);
and U36243 (N_36243,N_27121,N_21646);
and U36244 (N_36244,N_28427,N_24309);
or U36245 (N_36245,N_22553,N_28976);
and U36246 (N_36246,N_24393,N_26229);
nor U36247 (N_36247,N_21959,N_25833);
or U36248 (N_36248,N_21252,N_26780);
nor U36249 (N_36249,N_22401,N_26485);
or U36250 (N_36250,N_21628,N_29837);
and U36251 (N_36251,N_23720,N_23307);
or U36252 (N_36252,N_26534,N_28791);
and U36253 (N_36253,N_25511,N_25640);
nor U36254 (N_36254,N_23914,N_20886);
and U36255 (N_36255,N_23630,N_22324);
nand U36256 (N_36256,N_29616,N_21855);
xnor U36257 (N_36257,N_21890,N_29504);
nor U36258 (N_36258,N_24388,N_21685);
or U36259 (N_36259,N_23745,N_24874);
and U36260 (N_36260,N_29200,N_28522);
nor U36261 (N_36261,N_26557,N_24429);
or U36262 (N_36262,N_27510,N_22786);
or U36263 (N_36263,N_21392,N_21152);
nor U36264 (N_36264,N_25815,N_27151);
nor U36265 (N_36265,N_29606,N_25144);
or U36266 (N_36266,N_25596,N_24307);
or U36267 (N_36267,N_22600,N_21934);
and U36268 (N_36268,N_24063,N_29709);
or U36269 (N_36269,N_24573,N_22718);
xor U36270 (N_36270,N_21839,N_25180);
nor U36271 (N_36271,N_20305,N_29278);
and U36272 (N_36272,N_25682,N_28743);
xor U36273 (N_36273,N_21438,N_29942);
or U36274 (N_36274,N_25386,N_20363);
nor U36275 (N_36275,N_25561,N_26644);
and U36276 (N_36276,N_29848,N_27660);
and U36277 (N_36277,N_22326,N_23055);
or U36278 (N_36278,N_21578,N_26417);
nor U36279 (N_36279,N_23418,N_22422);
or U36280 (N_36280,N_29722,N_25314);
and U36281 (N_36281,N_26783,N_26866);
nor U36282 (N_36282,N_20836,N_21548);
and U36283 (N_36283,N_26214,N_28866);
or U36284 (N_36284,N_26403,N_29502);
nand U36285 (N_36285,N_25638,N_28759);
xnor U36286 (N_36286,N_25513,N_29350);
and U36287 (N_36287,N_29046,N_27655);
or U36288 (N_36288,N_21703,N_27993);
and U36289 (N_36289,N_25343,N_20578);
nand U36290 (N_36290,N_27580,N_20970);
and U36291 (N_36291,N_22320,N_27162);
nor U36292 (N_36292,N_26397,N_26681);
and U36293 (N_36293,N_28676,N_27355);
and U36294 (N_36294,N_20805,N_24380);
nand U36295 (N_36295,N_27920,N_29650);
or U36296 (N_36296,N_25315,N_26355);
and U36297 (N_36297,N_26953,N_26291);
nor U36298 (N_36298,N_22461,N_29755);
and U36299 (N_36299,N_27719,N_28049);
and U36300 (N_36300,N_21265,N_26516);
nand U36301 (N_36301,N_24892,N_29691);
or U36302 (N_36302,N_25708,N_29533);
and U36303 (N_36303,N_28094,N_22554);
or U36304 (N_36304,N_29534,N_26873);
or U36305 (N_36305,N_22254,N_24130);
and U36306 (N_36306,N_20444,N_29557);
and U36307 (N_36307,N_26348,N_25848);
nand U36308 (N_36308,N_22620,N_22053);
or U36309 (N_36309,N_21243,N_22916);
or U36310 (N_36310,N_21472,N_22179);
or U36311 (N_36311,N_25217,N_29391);
xnor U36312 (N_36312,N_22025,N_26171);
and U36313 (N_36313,N_29091,N_22451);
xnor U36314 (N_36314,N_25706,N_24755);
and U36315 (N_36315,N_23569,N_22608);
or U36316 (N_36316,N_22015,N_24999);
nor U36317 (N_36317,N_22146,N_27561);
xor U36318 (N_36318,N_21600,N_28426);
nor U36319 (N_36319,N_26604,N_25595);
nand U36320 (N_36320,N_20750,N_27792);
and U36321 (N_36321,N_22669,N_25731);
nand U36322 (N_36322,N_24006,N_25852);
nor U36323 (N_36323,N_29732,N_25266);
and U36324 (N_36324,N_24097,N_25112);
nand U36325 (N_36325,N_24958,N_28309);
nand U36326 (N_36326,N_26026,N_21631);
and U36327 (N_36327,N_21357,N_21343);
xor U36328 (N_36328,N_21591,N_26986);
xnor U36329 (N_36329,N_26640,N_22204);
and U36330 (N_36330,N_20995,N_27534);
or U36331 (N_36331,N_21690,N_22797);
or U36332 (N_36332,N_24455,N_26421);
nor U36333 (N_36333,N_22255,N_23813);
and U36334 (N_36334,N_25584,N_21778);
nand U36335 (N_36335,N_26628,N_22333);
or U36336 (N_36336,N_23496,N_27242);
nor U36337 (N_36337,N_20064,N_26938);
nand U36338 (N_36338,N_22503,N_27560);
xor U36339 (N_36339,N_28347,N_25075);
nand U36340 (N_36340,N_21488,N_23333);
or U36341 (N_36341,N_26531,N_22029);
or U36342 (N_36342,N_21013,N_21793);
nor U36343 (N_36343,N_24331,N_25796);
or U36344 (N_36344,N_29165,N_22481);
nor U36345 (N_36345,N_28943,N_25450);
nor U36346 (N_36346,N_25349,N_25977);
or U36347 (N_36347,N_29934,N_25169);
xor U36348 (N_36348,N_29428,N_27378);
nor U36349 (N_36349,N_28427,N_25899);
or U36350 (N_36350,N_26626,N_21797);
and U36351 (N_36351,N_25962,N_22795);
nand U36352 (N_36352,N_25583,N_22150);
nand U36353 (N_36353,N_29109,N_20323);
nand U36354 (N_36354,N_27382,N_21753);
nor U36355 (N_36355,N_29447,N_28624);
or U36356 (N_36356,N_26078,N_27862);
or U36357 (N_36357,N_28438,N_29992);
xor U36358 (N_36358,N_26304,N_27458);
or U36359 (N_36359,N_27133,N_23568);
nand U36360 (N_36360,N_26367,N_26563);
nand U36361 (N_36361,N_26466,N_22779);
xor U36362 (N_36362,N_29536,N_28942);
or U36363 (N_36363,N_21176,N_27294);
and U36364 (N_36364,N_26616,N_20282);
nor U36365 (N_36365,N_20452,N_24985);
and U36366 (N_36366,N_21647,N_20568);
nor U36367 (N_36367,N_29701,N_28705);
or U36368 (N_36368,N_22880,N_23041);
nor U36369 (N_36369,N_20706,N_29996);
and U36370 (N_36370,N_25339,N_24014);
or U36371 (N_36371,N_22072,N_29714);
xnor U36372 (N_36372,N_27824,N_22975);
nor U36373 (N_36373,N_25961,N_24863);
nand U36374 (N_36374,N_21916,N_22256);
nor U36375 (N_36375,N_21096,N_28943);
and U36376 (N_36376,N_22096,N_23838);
or U36377 (N_36377,N_29608,N_20336);
or U36378 (N_36378,N_21123,N_28615);
nor U36379 (N_36379,N_20616,N_23960);
nor U36380 (N_36380,N_27454,N_23373);
nand U36381 (N_36381,N_24757,N_23432);
or U36382 (N_36382,N_29038,N_23374);
xnor U36383 (N_36383,N_20179,N_21522);
and U36384 (N_36384,N_26403,N_25889);
or U36385 (N_36385,N_27876,N_27425);
or U36386 (N_36386,N_20985,N_28045);
nand U36387 (N_36387,N_26683,N_23276);
and U36388 (N_36388,N_21201,N_26919);
nor U36389 (N_36389,N_27528,N_23291);
or U36390 (N_36390,N_24627,N_28076);
and U36391 (N_36391,N_27346,N_28297);
nand U36392 (N_36392,N_20976,N_25448);
and U36393 (N_36393,N_29585,N_23844);
and U36394 (N_36394,N_27518,N_25695);
nor U36395 (N_36395,N_23608,N_22924);
nand U36396 (N_36396,N_22430,N_27917);
and U36397 (N_36397,N_22045,N_20926);
or U36398 (N_36398,N_27462,N_26394);
nand U36399 (N_36399,N_23817,N_24344);
and U36400 (N_36400,N_22496,N_25043);
nor U36401 (N_36401,N_28662,N_20184);
or U36402 (N_36402,N_23516,N_29751);
or U36403 (N_36403,N_25605,N_26284);
nor U36404 (N_36404,N_21404,N_25802);
nand U36405 (N_36405,N_24258,N_27418);
nand U36406 (N_36406,N_25940,N_20935);
nor U36407 (N_36407,N_23483,N_21938);
and U36408 (N_36408,N_21388,N_21916);
nand U36409 (N_36409,N_25038,N_28672);
nor U36410 (N_36410,N_26522,N_28589);
nor U36411 (N_36411,N_26661,N_22442);
nor U36412 (N_36412,N_22602,N_23477);
nand U36413 (N_36413,N_28790,N_21101);
nor U36414 (N_36414,N_27965,N_22196);
xor U36415 (N_36415,N_29007,N_22642);
or U36416 (N_36416,N_26613,N_20768);
and U36417 (N_36417,N_27131,N_24788);
nand U36418 (N_36418,N_29819,N_23648);
xor U36419 (N_36419,N_20691,N_29660);
or U36420 (N_36420,N_23404,N_24746);
nand U36421 (N_36421,N_22006,N_28218);
or U36422 (N_36422,N_29462,N_26551);
or U36423 (N_36423,N_21159,N_27175);
nor U36424 (N_36424,N_20692,N_22009);
nand U36425 (N_36425,N_24056,N_25733);
nand U36426 (N_36426,N_25658,N_26971);
or U36427 (N_36427,N_20646,N_21773);
or U36428 (N_36428,N_22475,N_26202);
or U36429 (N_36429,N_29584,N_21652);
or U36430 (N_36430,N_25773,N_26031);
and U36431 (N_36431,N_22693,N_24981);
nor U36432 (N_36432,N_25699,N_24627);
nor U36433 (N_36433,N_23454,N_25536);
nor U36434 (N_36434,N_22456,N_27725);
nand U36435 (N_36435,N_28032,N_23477);
and U36436 (N_36436,N_25589,N_24372);
nor U36437 (N_36437,N_27451,N_22185);
xor U36438 (N_36438,N_21116,N_21700);
or U36439 (N_36439,N_25074,N_25239);
and U36440 (N_36440,N_20955,N_27539);
and U36441 (N_36441,N_27247,N_26146);
or U36442 (N_36442,N_21978,N_24101);
nor U36443 (N_36443,N_25118,N_22046);
and U36444 (N_36444,N_20740,N_26840);
nor U36445 (N_36445,N_26548,N_26409);
or U36446 (N_36446,N_25144,N_27925);
and U36447 (N_36447,N_28410,N_20728);
xor U36448 (N_36448,N_28956,N_20269);
or U36449 (N_36449,N_27293,N_21978);
and U36450 (N_36450,N_28748,N_24433);
and U36451 (N_36451,N_24703,N_20271);
nor U36452 (N_36452,N_25165,N_27332);
and U36453 (N_36453,N_25509,N_28761);
or U36454 (N_36454,N_26219,N_21221);
xor U36455 (N_36455,N_29517,N_28708);
or U36456 (N_36456,N_25265,N_28109);
nand U36457 (N_36457,N_21416,N_21571);
nor U36458 (N_36458,N_25169,N_22223);
nand U36459 (N_36459,N_25651,N_27849);
or U36460 (N_36460,N_27145,N_24028);
or U36461 (N_36461,N_29691,N_22224);
and U36462 (N_36462,N_21231,N_21912);
nand U36463 (N_36463,N_24395,N_29752);
nor U36464 (N_36464,N_23436,N_25994);
nand U36465 (N_36465,N_25651,N_29965);
nand U36466 (N_36466,N_27954,N_27862);
and U36467 (N_36467,N_20439,N_23277);
nand U36468 (N_36468,N_29726,N_27289);
or U36469 (N_36469,N_22317,N_28647);
and U36470 (N_36470,N_27878,N_26694);
and U36471 (N_36471,N_22125,N_23965);
nand U36472 (N_36472,N_20912,N_21123);
nand U36473 (N_36473,N_26091,N_25958);
and U36474 (N_36474,N_28716,N_29172);
and U36475 (N_36475,N_25879,N_20992);
nor U36476 (N_36476,N_21697,N_21862);
nand U36477 (N_36477,N_27781,N_21341);
or U36478 (N_36478,N_27215,N_26159);
nand U36479 (N_36479,N_20527,N_27733);
nor U36480 (N_36480,N_25523,N_22765);
nand U36481 (N_36481,N_22908,N_23362);
xor U36482 (N_36482,N_20012,N_27282);
nor U36483 (N_36483,N_29360,N_24455);
nor U36484 (N_36484,N_27813,N_20409);
nand U36485 (N_36485,N_24760,N_22776);
nand U36486 (N_36486,N_26750,N_24409);
and U36487 (N_36487,N_28756,N_25259);
nor U36488 (N_36488,N_22022,N_24511);
and U36489 (N_36489,N_27238,N_22426);
nand U36490 (N_36490,N_28371,N_20368);
and U36491 (N_36491,N_22744,N_26256);
nor U36492 (N_36492,N_27041,N_29085);
nand U36493 (N_36493,N_26488,N_28113);
nor U36494 (N_36494,N_26566,N_21379);
xor U36495 (N_36495,N_25931,N_25853);
or U36496 (N_36496,N_23024,N_22544);
nand U36497 (N_36497,N_22597,N_22125);
and U36498 (N_36498,N_24755,N_26032);
nand U36499 (N_36499,N_21160,N_26873);
nor U36500 (N_36500,N_26006,N_21242);
or U36501 (N_36501,N_25301,N_21178);
and U36502 (N_36502,N_29068,N_21439);
and U36503 (N_36503,N_28163,N_27634);
nor U36504 (N_36504,N_24802,N_24837);
nor U36505 (N_36505,N_23519,N_25527);
nor U36506 (N_36506,N_24721,N_26531);
or U36507 (N_36507,N_29844,N_28516);
nor U36508 (N_36508,N_22710,N_22888);
and U36509 (N_36509,N_23464,N_26300);
nand U36510 (N_36510,N_26249,N_20145);
nor U36511 (N_36511,N_27360,N_24250);
nor U36512 (N_36512,N_24204,N_21100);
and U36513 (N_36513,N_28918,N_22993);
nor U36514 (N_36514,N_23734,N_20248);
or U36515 (N_36515,N_27273,N_20641);
and U36516 (N_36516,N_28423,N_28429);
nand U36517 (N_36517,N_27824,N_27657);
nor U36518 (N_36518,N_21495,N_25640);
xnor U36519 (N_36519,N_20428,N_20345);
nor U36520 (N_36520,N_24259,N_27667);
nand U36521 (N_36521,N_24162,N_21731);
or U36522 (N_36522,N_24037,N_25277);
nand U36523 (N_36523,N_25355,N_23235);
nand U36524 (N_36524,N_22858,N_23310);
nor U36525 (N_36525,N_22805,N_28416);
nor U36526 (N_36526,N_28770,N_21051);
or U36527 (N_36527,N_24425,N_22542);
nand U36528 (N_36528,N_29459,N_25791);
and U36529 (N_36529,N_25897,N_24236);
nor U36530 (N_36530,N_29832,N_24639);
nor U36531 (N_36531,N_21206,N_28134);
nor U36532 (N_36532,N_28825,N_23472);
or U36533 (N_36533,N_29125,N_21305);
or U36534 (N_36534,N_22231,N_24057);
or U36535 (N_36535,N_22160,N_27414);
nor U36536 (N_36536,N_29205,N_20476);
nor U36537 (N_36537,N_22835,N_27269);
and U36538 (N_36538,N_20618,N_27170);
and U36539 (N_36539,N_22226,N_21969);
and U36540 (N_36540,N_24326,N_27923);
or U36541 (N_36541,N_26305,N_25676);
nand U36542 (N_36542,N_29592,N_25780);
nand U36543 (N_36543,N_25014,N_26753);
nand U36544 (N_36544,N_24419,N_26562);
or U36545 (N_36545,N_22635,N_28528);
xnor U36546 (N_36546,N_28034,N_25466);
nand U36547 (N_36547,N_22602,N_27860);
and U36548 (N_36548,N_28682,N_29315);
or U36549 (N_36549,N_28591,N_21753);
and U36550 (N_36550,N_20946,N_25091);
or U36551 (N_36551,N_27435,N_24276);
nand U36552 (N_36552,N_23106,N_23203);
and U36553 (N_36553,N_28754,N_22198);
or U36554 (N_36554,N_29282,N_27455);
nor U36555 (N_36555,N_24006,N_29019);
and U36556 (N_36556,N_24849,N_28399);
xnor U36557 (N_36557,N_21846,N_25522);
and U36558 (N_36558,N_21159,N_29670);
nor U36559 (N_36559,N_25820,N_27614);
xnor U36560 (N_36560,N_28131,N_29801);
nand U36561 (N_36561,N_25012,N_24790);
or U36562 (N_36562,N_22974,N_24010);
nand U36563 (N_36563,N_21136,N_29042);
and U36564 (N_36564,N_24902,N_29351);
and U36565 (N_36565,N_28909,N_22525);
nand U36566 (N_36566,N_22942,N_29126);
or U36567 (N_36567,N_28072,N_24860);
xnor U36568 (N_36568,N_22492,N_22566);
or U36569 (N_36569,N_25860,N_24472);
nand U36570 (N_36570,N_24399,N_28247);
xnor U36571 (N_36571,N_27847,N_20614);
nand U36572 (N_36572,N_28176,N_28550);
nor U36573 (N_36573,N_28715,N_26693);
nand U36574 (N_36574,N_21461,N_25174);
and U36575 (N_36575,N_28949,N_29215);
nand U36576 (N_36576,N_27072,N_25887);
nand U36577 (N_36577,N_26550,N_20712);
nor U36578 (N_36578,N_22897,N_23343);
or U36579 (N_36579,N_20452,N_29725);
or U36580 (N_36580,N_26053,N_25831);
nor U36581 (N_36581,N_25737,N_24508);
nand U36582 (N_36582,N_22072,N_27421);
or U36583 (N_36583,N_27290,N_28387);
nand U36584 (N_36584,N_23656,N_23586);
and U36585 (N_36585,N_20888,N_22132);
and U36586 (N_36586,N_20567,N_23599);
nor U36587 (N_36587,N_28795,N_28823);
or U36588 (N_36588,N_24102,N_26273);
nor U36589 (N_36589,N_28807,N_23992);
nand U36590 (N_36590,N_21955,N_27743);
nor U36591 (N_36591,N_28336,N_24367);
nand U36592 (N_36592,N_29921,N_20424);
and U36593 (N_36593,N_26091,N_28595);
nand U36594 (N_36594,N_29835,N_27578);
nor U36595 (N_36595,N_25370,N_27514);
and U36596 (N_36596,N_28823,N_20381);
xnor U36597 (N_36597,N_26757,N_26415);
nor U36598 (N_36598,N_23337,N_29730);
nor U36599 (N_36599,N_20873,N_23841);
nor U36600 (N_36600,N_27735,N_28607);
or U36601 (N_36601,N_29639,N_27691);
nand U36602 (N_36602,N_26253,N_26352);
xor U36603 (N_36603,N_25996,N_21565);
xor U36604 (N_36604,N_23251,N_26256);
xnor U36605 (N_36605,N_29555,N_27721);
nor U36606 (N_36606,N_23706,N_20386);
and U36607 (N_36607,N_26099,N_27283);
and U36608 (N_36608,N_27270,N_23312);
and U36609 (N_36609,N_25512,N_26529);
or U36610 (N_36610,N_20382,N_26883);
nand U36611 (N_36611,N_24477,N_28148);
nor U36612 (N_36612,N_24062,N_22625);
nor U36613 (N_36613,N_23033,N_21793);
or U36614 (N_36614,N_26239,N_26807);
or U36615 (N_36615,N_23875,N_26524);
or U36616 (N_36616,N_25069,N_25133);
nand U36617 (N_36617,N_25343,N_27156);
and U36618 (N_36618,N_28885,N_26454);
nand U36619 (N_36619,N_24522,N_27661);
and U36620 (N_36620,N_22973,N_21030);
xnor U36621 (N_36621,N_21989,N_26796);
xnor U36622 (N_36622,N_29144,N_20352);
or U36623 (N_36623,N_27659,N_29299);
xnor U36624 (N_36624,N_27969,N_20494);
nand U36625 (N_36625,N_23143,N_20067);
and U36626 (N_36626,N_20859,N_25024);
nand U36627 (N_36627,N_27266,N_21177);
nand U36628 (N_36628,N_29989,N_29012);
nor U36629 (N_36629,N_23725,N_26424);
nand U36630 (N_36630,N_24430,N_22884);
nand U36631 (N_36631,N_24295,N_23820);
or U36632 (N_36632,N_25299,N_21345);
and U36633 (N_36633,N_28945,N_26896);
or U36634 (N_36634,N_22632,N_21683);
or U36635 (N_36635,N_28728,N_26363);
or U36636 (N_36636,N_26030,N_25493);
or U36637 (N_36637,N_29032,N_20184);
or U36638 (N_36638,N_29662,N_26770);
nor U36639 (N_36639,N_24711,N_25046);
xnor U36640 (N_36640,N_20005,N_22243);
or U36641 (N_36641,N_25950,N_20448);
nand U36642 (N_36642,N_26456,N_23538);
and U36643 (N_36643,N_24557,N_27753);
nor U36644 (N_36644,N_21941,N_27530);
or U36645 (N_36645,N_26733,N_20933);
or U36646 (N_36646,N_25801,N_21360);
nand U36647 (N_36647,N_23793,N_25520);
nor U36648 (N_36648,N_24601,N_26738);
and U36649 (N_36649,N_22729,N_26143);
nor U36650 (N_36650,N_21904,N_21800);
nand U36651 (N_36651,N_27129,N_22722);
nand U36652 (N_36652,N_21051,N_23530);
and U36653 (N_36653,N_24938,N_26566);
xnor U36654 (N_36654,N_22572,N_29131);
or U36655 (N_36655,N_21560,N_29506);
nand U36656 (N_36656,N_20608,N_27100);
nand U36657 (N_36657,N_27669,N_21423);
or U36658 (N_36658,N_23062,N_21457);
nand U36659 (N_36659,N_28625,N_21473);
nand U36660 (N_36660,N_20404,N_23225);
and U36661 (N_36661,N_24208,N_21955);
or U36662 (N_36662,N_20223,N_29518);
nor U36663 (N_36663,N_28507,N_27609);
or U36664 (N_36664,N_25302,N_28899);
nor U36665 (N_36665,N_27321,N_21175);
nor U36666 (N_36666,N_25175,N_20501);
or U36667 (N_36667,N_21454,N_29215);
nand U36668 (N_36668,N_26520,N_21355);
and U36669 (N_36669,N_20549,N_21618);
nand U36670 (N_36670,N_22034,N_23882);
and U36671 (N_36671,N_25309,N_24807);
nor U36672 (N_36672,N_26042,N_23095);
and U36673 (N_36673,N_27617,N_21597);
and U36674 (N_36674,N_27100,N_25963);
nand U36675 (N_36675,N_20408,N_25434);
nand U36676 (N_36676,N_28398,N_22356);
nor U36677 (N_36677,N_27220,N_23822);
or U36678 (N_36678,N_27182,N_29192);
or U36679 (N_36679,N_21082,N_27114);
nor U36680 (N_36680,N_24617,N_21045);
nand U36681 (N_36681,N_24788,N_23465);
and U36682 (N_36682,N_25655,N_26631);
nand U36683 (N_36683,N_20299,N_25942);
nand U36684 (N_36684,N_27677,N_21936);
or U36685 (N_36685,N_29151,N_26185);
nor U36686 (N_36686,N_25631,N_26245);
and U36687 (N_36687,N_25426,N_25815);
xor U36688 (N_36688,N_21319,N_20654);
nor U36689 (N_36689,N_25052,N_26628);
nand U36690 (N_36690,N_29328,N_24017);
nor U36691 (N_36691,N_25370,N_24600);
or U36692 (N_36692,N_27669,N_21569);
xor U36693 (N_36693,N_29158,N_24713);
nor U36694 (N_36694,N_24349,N_26088);
nor U36695 (N_36695,N_28640,N_23112);
or U36696 (N_36696,N_25743,N_26360);
xor U36697 (N_36697,N_20822,N_22254);
and U36698 (N_36698,N_28148,N_25640);
nor U36699 (N_36699,N_27935,N_25222);
xor U36700 (N_36700,N_25536,N_22265);
and U36701 (N_36701,N_21033,N_26659);
nor U36702 (N_36702,N_23841,N_28781);
nand U36703 (N_36703,N_29230,N_28090);
nor U36704 (N_36704,N_20415,N_27905);
and U36705 (N_36705,N_27808,N_28118);
nand U36706 (N_36706,N_23724,N_24075);
nor U36707 (N_36707,N_25363,N_24058);
and U36708 (N_36708,N_28922,N_26980);
nand U36709 (N_36709,N_21682,N_29927);
nand U36710 (N_36710,N_20473,N_29156);
nand U36711 (N_36711,N_20443,N_24794);
nand U36712 (N_36712,N_29580,N_20852);
nor U36713 (N_36713,N_20592,N_23188);
or U36714 (N_36714,N_25553,N_24294);
and U36715 (N_36715,N_21574,N_28305);
and U36716 (N_36716,N_29101,N_29798);
nor U36717 (N_36717,N_21696,N_22577);
or U36718 (N_36718,N_21465,N_28289);
and U36719 (N_36719,N_21084,N_28990);
or U36720 (N_36720,N_20900,N_20983);
xnor U36721 (N_36721,N_27032,N_23609);
nor U36722 (N_36722,N_29469,N_25234);
xnor U36723 (N_36723,N_27543,N_25178);
nand U36724 (N_36724,N_23954,N_23899);
and U36725 (N_36725,N_28715,N_23821);
or U36726 (N_36726,N_27815,N_25065);
and U36727 (N_36727,N_26694,N_23580);
and U36728 (N_36728,N_22280,N_28945);
nor U36729 (N_36729,N_29908,N_26991);
nand U36730 (N_36730,N_25104,N_23569);
nand U36731 (N_36731,N_26499,N_23648);
and U36732 (N_36732,N_27775,N_20673);
nor U36733 (N_36733,N_23494,N_27674);
and U36734 (N_36734,N_21654,N_29145);
nor U36735 (N_36735,N_21949,N_22967);
nand U36736 (N_36736,N_29039,N_29890);
nand U36737 (N_36737,N_23028,N_29442);
xnor U36738 (N_36738,N_20781,N_24036);
or U36739 (N_36739,N_25851,N_22910);
nand U36740 (N_36740,N_21191,N_22391);
nor U36741 (N_36741,N_23505,N_26780);
nand U36742 (N_36742,N_25785,N_21616);
nand U36743 (N_36743,N_29714,N_21466);
and U36744 (N_36744,N_28241,N_26781);
nor U36745 (N_36745,N_29502,N_20587);
nand U36746 (N_36746,N_21615,N_27841);
nand U36747 (N_36747,N_20128,N_26431);
and U36748 (N_36748,N_23137,N_28742);
nor U36749 (N_36749,N_22871,N_25823);
nor U36750 (N_36750,N_24174,N_29293);
nor U36751 (N_36751,N_23241,N_26139);
nand U36752 (N_36752,N_21313,N_28318);
or U36753 (N_36753,N_25119,N_20056);
or U36754 (N_36754,N_21145,N_24621);
and U36755 (N_36755,N_22551,N_20768);
and U36756 (N_36756,N_26207,N_27547);
nor U36757 (N_36757,N_27961,N_29201);
and U36758 (N_36758,N_23927,N_25210);
or U36759 (N_36759,N_28137,N_25381);
nor U36760 (N_36760,N_29008,N_22531);
nand U36761 (N_36761,N_24623,N_26339);
or U36762 (N_36762,N_26076,N_24480);
and U36763 (N_36763,N_22641,N_28326);
and U36764 (N_36764,N_22370,N_25846);
nor U36765 (N_36765,N_29129,N_20498);
or U36766 (N_36766,N_20849,N_28311);
nand U36767 (N_36767,N_25694,N_28605);
nand U36768 (N_36768,N_27823,N_28455);
xor U36769 (N_36769,N_25480,N_27031);
nand U36770 (N_36770,N_22482,N_29480);
xor U36771 (N_36771,N_29386,N_25394);
or U36772 (N_36772,N_27152,N_29651);
nor U36773 (N_36773,N_21213,N_20409);
nor U36774 (N_36774,N_23080,N_29283);
or U36775 (N_36775,N_23979,N_20097);
or U36776 (N_36776,N_28213,N_29218);
and U36777 (N_36777,N_23545,N_27121);
nand U36778 (N_36778,N_26821,N_22573);
or U36779 (N_36779,N_25511,N_21974);
and U36780 (N_36780,N_24575,N_29182);
nor U36781 (N_36781,N_25522,N_28359);
and U36782 (N_36782,N_20039,N_25554);
nor U36783 (N_36783,N_24733,N_21508);
and U36784 (N_36784,N_28864,N_28085);
and U36785 (N_36785,N_23109,N_26899);
nand U36786 (N_36786,N_21846,N_23146);
nor U36787 (N_36787,N_22436,N_21676);
and U36788 (N_36788,N_29369,N_26067);
or U36789 (N_36789,N_25567,N_20261);
and U36790 (N_36790,N_27184,N_24134);
and U36791 (N_36791,N_29662,N_21472);
nor U36792 (N_36792,N_27327,N_24508);
nor U36793 (N_36793,N_22778,N_20848);
or U36794 (N_36794,N_26677,N_23718);
nor U36795 (N_36795,N_27223,N_24014);
or U36796 (N_36796,N_24520,N_26842);
nor U36797 (N_36797,N_21303,N_21365);
nand U36798 (N_36798,N_22061,N_20565);
nand U36799 (N_36799,N_24323,N_29637);
or U36800 (N_36800,N_25883,N_22191);
nor U36801 (N_36801,N_28951,N_27514);
nand U36802 (N_36802,N_21367,N_24456);
and U36803 (N_36803,N_25741,N_21653);
or U36804 (N_36804,N_26988,N_29254);
nand U36805 (N_36805,N_28252,N_29668);
nor U36806 (N_36806,N_28297,N_27338);
nand U36807 (N_36807,N_21267,N_23135);
or U36808 (N_36808,N_27726,N_22719);
nor U36809 (N_36809,N_21814,N_26076);
and U36810 (N_36810,N_28702,N_20182);
nor U36811 (N_36811,N_20175,N_24012);
or U36812 (N_36812,N_21706,N_27621);
or U36813 (N_36813,N_28010,N_22577);
and U36814 (N_36814,N_26336,N_29154);
nor U36815 (N_36815,N_28739,N_25777);
nand U36816 (N_36816,N_26971,N_22209);
and U36817 (N_36817,N_25802,N_27483);
or U36818 (N_36818,N_22086,N_21681);
and U36819 (N_36819,N_20395,N_27174);
or U36820 (N_36820,N_22168,N_24869);
nand U36821 (N_36821,N_27523,N_26023);
xor U36822 (N_36822,N_24499,N_25345);
xor U36823 (N_36823,N_27265,N_25086);
xor U36824 (N_36824,N_21279,N_27801);
and U36825 (N_36825,N_25651,N_25349);
or U36826 (N_36826,N_22088,N_26674);
nor U36827 (N_36827,N_21313,N_27562);
or U36828 (N_36828,N_28858,N_20353);
nand U36829 (N_36829,N_22846,N_29967);
nor U36830 (N_36830,N_22676,N_25658);
nor U36831 (N_36831,N_27161,N_21105);
xor U36832 (N_36832,N_22824,N_24817);
nor U36833 (N_36833,N_24393,N_20110);
and U36834 (N_36834,N_23391,N_21382);
or U36835 (N_36835,N_22063,N_23451);
xor U36836 (N_36836,N_27699,N_27065);
nor U36837 (N_36837,N_27480,N_20447);
or U36838 (N_36838,N_27533,N_23464);
nor U36839 (N_36839,N_29253,N_20121);
and U36840 (N_36840,N_23233,N_26302);
or U36841 (N_36841,N_29887,N_24812);
nand U36842 (N_36842,N_22527,N_22851);
nand U36843 (N_36843,N_20296,N_23663);
nor U36844 (N_36844,N_21797,N_22828);
or U36845 (N_36845,N_26519,N_25549);
or U36846 (N_36846,N_25109,N_24184);
nand U36847 (N_36847,N_23489,N_20018);
nor U36848 (N_36848,N_27491,N_27790);
nand U36849 (N_36849,N_25489,N_22356);
nand U36850 (N_36850,N_29142,N_27662);
and U36851 (N_36851,N_24950,N_27718);
nor U36852 (N_36852,N_22939,N_24859);
and U36853 (N_36853,N_23817,N_28598);
nand U36854 (N_36854,N_23193,N_27483);
and U36855 (N_36855,N_21842,N_29973);
or U36856 (N_36856,N_21491,N_21820);
nor U36857 (N_36857,N_21345,N_27700);
xor U36858 (N_36858,N_20817,N_27652);
xnor U36859 (N_36859,N_24579,N_28981);
nor U36860 (N_36860,N_29087,N_23380);
and U36861 (N_36861,N_25601,N_27218);
and U36862 (N_36862,N_26147,N_26580);
or U36863 (N_36863,N_27710,N_25812);
nor U36864 (N_36864,N_26385,N_25060);
xnor U36865 (N_36865,N_22825,N_25745);
xor U36866 (N_36866,N_27875,N_27554);
or U36867 (N_36867,N_28645,N_22142);
or U36868 (N_36868,N_25148,N_22540);
xor U36869 (N_36869,N_28118,N_24397);
and U36870 (N_36870,N_26267,N_29630);
and U36871 (N_36871,N_22586,N_27395);
nor U36872 (N_36872,N_20591,N_27798);
and U36873 (N_36873,N_28399,N_25677);
and U36874 (N_36874,N_26985,N_28879);
xnor U36875 (N_36875,N_28909,N_20963);
or U36876 (N_36876,N_21834,N_25527);
nor U36877 (N_36877,N_25264,N_23226);
xnor U36878 (N_36878,N_22941,N_29954);
and U36879 (N_36879,N_28055,N_29968);
and U36880 (N_36880,N_22120,N_21978);
and U36881 (N_36881,N_27603,N_25793);
nand U36882 (N_36882,N_20025,N_23692);
and U36883 (N_36883,N_28749,N_22674);
nor U36884 (N_36884,N_25095,N_27855);
nand U36885 (N_36885,N_23860,N_29823);
or U36886 (N_36886,N_26695,N_20378);
nand U36887 (N_36887,N_26893,N_28191);
xor U36888 (N_36888,N_28876,N_23193);
or U36889 (N_36889,N_23678,N_22258);
nor U36890 (N_36890,N_20538,N_20003);
or U36891 (N_36891,N_23901,N_26384);
or U36892 (N_36892,N_25924,N_22275);
or U36893 (N_36893,N_29417,N_28326);
xnor U36894 (N_36894,N_25854,N_28640);
nand U36895 (N_36895,N_21286,N_20554);
and U36896 (N_36896,N_22870,N_28874);
and U36897 (N_36897,N_26835,N_27879);
nand U36898 (N_36898,N_23160,N_22329);
and U36899 (N_36899,N_24398,N_27883);
or U36900 (N_36900,N_26119,N_24014);
xnor U36901 (N_36901,N_27494,N_22878);
or U36902 (N_36902,N_26112,N_21690);
and U36903 (N_36903,N_23393,N_23407);
xnor U36904 (N_36904,N_25284,N_29423);
or U36905 (N_36905,N_26991,N_20494);
nor U36906 (N_36906,N_29270,N_29080);
and U36907 (N_36907,N_28802,N_20981);
or U36908 (N_36908,N_28266,N_22173);
and U36909 (N_36909,N_26428,N_26856);
nand U36910 (N_36910,N_24740,N_21564);
nand U36911 (N_36911,N_26515,N_28331);
or U36912 (N_36912,N_23799,N_24301);
and U36913 (N_36913,N_22664,N_25853);
or U36914 (N_36914,N_24559,N_28779);
xor U36915 (N_36915,N_24845,N_23060);
or U36916 (N_36916,N_28748,N_24604);
nand U36917 (N_36917,N_20979,N_26643);
or U36918 (N_36918,N_29403,N_24606);
and U36919 (N_36919,N_29982,N_21764);
nand U36920 (N_36920,N_21131,N_23010);
nor U36921 (N_36921,N_23483,N_25747);
nand U36922 (N_36922,N_25373,N_24382);
or U36923 (N_36923,N_25048,N_27754);
and U36924 (N_36924,N_24541,N_22186);
nand U36925 (N_36925,N_28456,N_20619);
and U36926 (N_36926,N_23185,N_23325);
xnor U36927 (N_36927,N_20015,N_21706);
and U36928 (N_36928,N_25874,N_22888);
or U36929 (N_36929,N_20857,N_28385);
nand U36930 (N_36930,N_20374,N_21152);
nor U36931 (N_36931,N_26865,N_21910);
or U36932 (N_36932,N_25883,N_29272);
nand U36933 (N_36933,N_22271,N_22433);
nor U36934 (N_36934,N_28672,N_22886);
or U36935 (N_36935,N_20958,N_22486);
and U36936 (N_36936,N_29252,N_22473);
xor U36937 (N_36937,N_29724,N_24346);
or U36938 (N_36938,N_20513,N_23472);
xor U36939 (N_36939,N_22415,N_21003);
nand U36940 (N_36940,N_28371,N_22230);
nor U36941 (N_36941,N_22933,N_27035);
or U36942 (N_36942,N_24562,N_27828);
or U36943 (N_36943,N_26601,N_25742);
nor U36944 (N_36944,N_27499,N_27397);
xor U36945 (N_36945,N_22929,N_24027);
nand U36946 (N_36946,N_20863,N_22334);
and U36947 (N_36947,N_21403,N_28077);
and U36948 (N_36948,N_28562,N_27245);
xnor U36949 (N_36949,N_24862,N_25103);
xnor U36950 (N_36950,N_26900,N_24882);
nand U36951 (N_36951,N_21030,N_25468);
and U36952 (N_36952,N_29239,N_26084);
nand U36953 (N_36953,N_24567,N_29582);
and U36954 (N_36954,N_22335,N_24102);
nor U36955 (N_36955,N_23469,N_28415);
and U36956 (N_36956,N_21753,N_26924);
and U36957 (N_36957,N_20731,N_28147);
or U36958 (N_36958,N_22283,N_24805);
and U36959 (N_36959,N_20085,N_22704);
nor U36960 (N_36960,N_20811,N_26176);
and U36961 (N_36961,N_27532,N_20186);
and U36962 (N_36962,N_22685,N_24821);
nand U36963 (N_36963,N_22836,N_20522);
and U36964 (N_36964,N_24512,N_21341);
and U36965 (N_36965,N_27903,N_26942);
nand U36966 (N_36966,N_27445,N_21843);
nor U36967 (N_36967,N_28465,N_26755);
or U36968 (N_36968,N_23608,N_29239);
or U36969 (N_36969,N_28954,N_24913);
or U36970 (N_36970,N_23206,N_21150);
or U36971 (N_36971,N_23849,N_24091);
and U36972 (N_36972,N_20065,N_24711);
and U36973 (N_36973,N_28358,N_20760);
and U36974 (N_36974,N_24819,N_24431);
nand U36975 (N_36975,N_24194,N_21198);
nor U36976 (N_36976,N_26724,N_20691);
nand U36977 (N_36977,N_24091,N_22817);
and U36978 (N_36978,N_21844,N_28599);
nor U36979 (N_36979,N_24812,N_26143);
or U36980 (N_36980,N_23105,N_25059);
and U36981 (N_36981,N_28002,N_20313);
and U36982 (N_36982,N_20872,N_28164);
or U36983 (N_36983,N_25005,N_23424);
nor U36984 (N_36984,N_26659,N_23048);
and U36985 (N_36985,N_21032,N_21261);
and U36986 (N_36986,N_29029,N_26780);
and U36987 (N_36987,N_29563,N_26888);
or U36988 (N_36988,N_23336,N_29900);
or U36989 (N_36989,N_24221,N_23546);
nor U36990 (N_36990,N_28092,N_27509);
or U36991 (N_36991,N_22859,N_24381);
nor U36992 (N_36992,N_29138,N_29534);
or U36993 (N_36993,N_25531,N_23950);
nand U36994 (N_36994,N_24263,N_26535);
nor U36995 (N_36995,N_27158,N_26200);
nand U36996 (N_36996,N_20787,N_21247);
nor U36997 (N_36997,N_24068,N_24811);
nand U36998 (N_36998,N_21198,N_27683);
or U36999 (N_36999,N_20589,N_26329);
nor U37000 (N_37000,N_28087,N_28639);
xor U37001 (N_37001,N_22066,N_28242);
or U37002 (N_37002,N_20116,N_21975);
and U37003 (N_37003,N_25474,N_27757);
and U37004 (N_37004,N_20905,N_23976);
nand U37005 (N_37005,N_21557,N_22983);
nor U37006 (N_37006,N_20254,N_21386);
or U37007 (N_37007,N_27623,N_22980);
or U37008 (N_37008,N_20178,N_27923);
nor U37009 (N_37009,N_24074,N_22774);
or U37010 (N_37010,N_27925,N_24255);
and U37011 (N_37011,N_28239,N_23729);
nor U37012 (N_37012,N_24163,N_21159);
nor U37013 (N_37013,N_25323,N_25889);
xor U37014 (N_37014,N_28342,N_27858);
or U37015 (N_37015,N_26773,N_22451);
or U37016 (N_37016,N_28507,N_20068);
nor U37017 (N_37017,N_20348,N_24875);
nor U37018 (N_37018,N_26151,N_23890);
or U37019 (N_37019,N_20123,N_25385);
nor U37020 (N_37020,N_20863,N_29368);
and U37021 (N_37021,N_26121,N_24848);
and U37022 (N_37022,N_28913,N_21991);
or U37023 (N_37023,N_28705,N_26424);
nand U37024 (N_37024,N_23005,N_25991);
nand U37025 (N_37025,N_25847,N_20604);
nand U37026 (N_37026,N_29665,N_29355);
nand U37027 (N_37027,N_23308,N_24265);
nor U37028 (N_37028,N_28412,N_22415);
or U37029 (N_37029,N_28243,N_21231);
or U37030 (N_37030,N_21151,N_28848);
xnor U37031 (N_37031,N_25022,N_20673);
and U37032 (N_37032,N_29900,N_24450);
nand U37033 (N_37033,N_24166,N_26695);
or U37034 (N_37034,N_29238,N_27756);
nand U37035 (N_37035,N_22470,N_21143);
nor U37036 (N_37036,N_21539,N_28595);
nor U37037 (N_37037,N_23077,N_25181);
nor U37038 (N_37038,N_29263,N_28654);
and U37039 (N_37039,N_21377,N_29816);
and U37040 (N_37040,N_21961,N_27602);
nand U37041 (N_37041,N_21639,N_25166);
nor U37042 (N_37042,N_27700,N_20476);
xor U37043 (N_37043,N_23694,N_23666);
or U37044 (N_37044,N_21498,N_20413);
or U37045 (N_37045,N_22803,N_21533);
xor U37046 (N_37046,N_22893,N_25884);
nand U37047 (N_37047,N_29693,N_28530);
or U37048 (N_37048,N_24266,N_21105);
and U37049 (N_37049,N_22202,N_29340);
and U37050 (N_37050,N_24519,N_23969);
and U37051 (N_37051,N_28615,N_28454);
nor U37052 (N_37052,N_28044,N_21688);
nand U37053 (N_37053,N_28663,N_27482);
nand U37054 (N_37054,N_22383,N_20696);
nor U37055 (N_37055,N_29059,N_27630);
and U37056 (N_37056,N_23940,N_21768);
nand U37057 (N_37057,N_22017,N_28264);
and U37058 (N_37058,N_21238,N_23923);
nor U37059 (N_37059,N_24125,N_26040);
nand U37060 (N_37060,N_24801,N_25512);
xnor U37061 (N_37061,N_29230,N_29560);
nand U37062 (N_37062,N_23682,N_22483);
nor U37063 (N_37063,N_26663,N_25939);
nand U37064 (N_37064,N_26876,N_28169);
nor U37065 (N_37065,N_29142,N_25601);
or U37066 (N_37066,N_21343,N_20808);
and U37067 (N_37067,N_29544,N_23426);
or U37068 (N_37068,N_20671,N_26858);
nor U37069 (N_37069,N_24559,N_22661);
and U37070 (N_37070,N_21630,N_26264);
nor U37071 (N_37071,N_23087,N_24417);
and U37072 (N_37072,N_25528,N_26785);
nand U37073 (N_37073,N_27648,N_26644);
nor U37074 (N_37074,N_28378,N_25639);
nand U37075 (N_37075,N_20496,N_22283);
and U37076 (N_37076,N_29454,N_28861);
nor U37077 (N_37077,N_21433,N_20289);
or U37078 (N_37078,N_22801,N_24464);
or U37079 (N_37079,N_27281,N_21571);
or U37080 (N_37080,N_25625,N_25626);
or U37081 (N_37081,N_21904,N_23946);
or U37082 (N_37082,N_22726,N_29872);
and U37083 (N_37083,N_25156,N_28345);
or U37084 (N_37084,N_24751,N_20326);
or U37085 (N_37085,N_20589,N_25251);
and U37086 (N_37086,N_29762,N_23999);
or U37087 (N_37087,N_26026,N_24409);
xnor U37088 (N_37088,N_29984,N_23078);
and U37089 (N_37089,N_23346,N_27211);
or U37090 (N_37090,N_24072,N_23090);
and U37091 (N_37091,N_21882,N_21773);
xor U37092 (N_37092,N_22226,N_22052);
nand U37093 (N_37093,N_28004,N_25415);
or U37094 (N_37094,N_28370,N_27029);
nor U37095 (N_37095,N_29670,N_24149);
nor U37096 (N_37096,N_22111,N_22539);
nand U37097 (N_37097,N_24996,N_26822);
nor U37098 (N_37098,N_23657,N_20191);
and U37099 (N_37099,N_29026,N_23057);
or U37100 (N_37100,N_29183,N_25257);
xor U37101 (N_37101,N_27433,N_26003);
or U37102 (N_37102,N_24408,N_25471);
nor U37103 (N_37103,N_24649,N_20012);
nor U37104 (N_37104,N_27363,N_21156);
and U37105 (N_37105,N_27942,N_22892);
and U37106 (N_37106,N_23366,N_23473);
nor U37107 (N_37107,N_25272,N_22943);
nor U37108 (N_37108,N_23793,N_28102);
nand U37109 (N_37109,N_26567,N_24210);
or U37110 (N_37110,N_26719,N_24836);
nor U37111 (N_37111,N_27619,N_23311);
nand U37112 (N_37112,N_25573,N_24509);
xor U37113 (N_37113,N_21499,N_20147);
nor U37114 (N_37114,N_24296,N_21383);
nor U37115 (N_37115,N_27314,N_22880);
xnor U37116 (N_37116,N_22760,N_27689);
nand U37117 (N_37117,N_24463,N_28715);
nor U37118 (N_37118,N_27761,N_28949);
or U37119 (N_37119,N_22814,N_29376);
or U37120 (N_37120,N_28279,N_23816);
or U37121 (N_37121,N_27729,N_20653);
nand U37122 (N_37122,N_27549,N_20242);
and U37123 (N_37123,N_20902,N_29208);
or U37124 (N_37124,N_27653,N_25176);
xnor U37125 (N_37125,N_23306,N_23939);
nor U37126 (N_37126,N_23621,N_25386);
nor U37127 (N_37127,N_25226,N_25279);
nor U37128 (N_37128,N_22633,N_23594);
nor U37129 (N_37129,N_21366,N_24993);
xnor U37130 (N_37130,N_20280,N_20902);
nor U37131 (N_37131,N_27334,N_25396);
nand U37132 (N_37132,N_25517,N_25176);
xnor U37133 (N_37133,N_20518,N_28824);
nor U37134 (N_37134,N_20251,N_28324);
nand U37135 (N_37135,N_24102,N_20303);
nor U37136 (N_37136,N_29893,N_20742);
nor U37137 (N_37137,N_24155,N_29338);
nand U37138 (N_37138,N_20033,N_20092);
or U37139 (N_37139,N_29074,N_27093);
and U37140 (N_37140,N_22409,N_27441);
nor U37141 (N_37141,N_23609,N_25007);
and U37142 (N_37142,N_24629,N_25454);
nand U37143 (N_37143,N_22345,N_20409);
nand U37144 (N_37144,N_26335,N_27420);
xnor U37145 (N_37145,N_25499,N_26299);
nand U37146 (N_37146,N_21375,N_27277);
nand U37147 (N_37147,N_27188,N_21032);
nor U37148 (N_37148,N_20593,N_21375);
nor U37149 (N_37149,N_24294,N_29577);
and U37150 (N_37150,N_26216,N_23588);
and U37151 (N_37151,N_24763,N_29170);
or U37152 (N_37152,N_26585,N_26483);
nor U37153 (N_37153,N_29648,N_26022);
xor U37154 (N_37154,N_29218,N_25550);
nand U37155 (N_37155,N_27168,N_22503);
nor U37156 (N_37156,N_23941,N_29035);
or U37157 (N_37157,N_27540,N_20818);
nand U37158 (N_37158,N_27959,N_23109);
xnor U37159 (N_37159,N_22785,N_20891);
nand U37160 (N_37160,N_23591,N_24540);
nor U37161 (N_37161,N_29676,N_22674);
nand U37162 (N_37162,N_23132,N_26994);
and U37163 (N_37163,N_24212,N_24225);
or U37164 (N_37164,N_22502,N_21122);
nand U37165 (N_37165,N_23663,N_25879);
or U37166 (N_37166,N_29045,N_28074);
and U37167 (N_37167,N_23460,N_26875);
nand U37168 (N_37168,N_25613,N_23177);
nor U37169 (N_37169,N_21528,N_26790);
nand U37170 (N_37170,N_29844,N_23447);
nor U37171 (N_37171,N_24716,N_20287);
and U37172 (N_37172,N_25368,N_22440);
nand U37173 (N_37173,N_20351,N_23076);
or U37174 (N_37174,N_22568,N_27006);
nand U37175 (N_37175,N_22906,N_21499);
or U37176 (N_37176,N_23423,N_20536);
xnor U37177 (N_37177,N_21016,N_25700);
nor U37178 (N_37178,N_23700,N_21981);
nor U37179 (N_37179,N_23005,N_26214);
nor U37180 (N_37180,N_29389,N_28570);
or U37181 (N_37181,N_26043,N_22274);
and U37182 (N_37182,N_26227,N_21602);
or U37183 (N_37183,N_24946,N_27535);
and U37184 (N_37184,N_25347,N_23245);
nand U37185 (N_37185,N_25446,N_22052);
or U37186 (N_37186,N_29519,N_26498);
nor U37187 (N_37187,N_21708,N_27338);
or U37188 (N_37188,N_22092,N_25201);
or U37189 (N_37189,N_20034,N_20384);
xnor U37190 (N_37190,N_27470,N_23334);
xor U37191 (N_37191,N_21995,N_25604);
nand U37192 (N_37192,N_25745,N_20406);
nand U37193 (N_37193,N_22224,N_24833);
nor U37194 (N_37194,N_21251,N_24312);
nor U37195 (N_37195,N_25752,N_26440);
xor U37196 (N_37196,N_27149,N_22031);
nor U37197 (N_37197,N_22296,N_26223);
nand U37198 (N_37198,N_26910,N_27738);
nand U37199 (N_37199,N_22868,N_23441);
and U37200 (N_37200,N_28085,N_22251);
nor U37201 (N_37201,N_25757,N_29631);
or U37202 (N_37202,N_23076,N_21666);
nor U37203 (N_37203,N_28491,N_25652);
and U37204 (N_37204,N_23778,N_27151);
xor U37205 (N_37205,N_28649,N_26620);
xnor U37206 (N_37206,N_27114,N_23500);
or U37207 (N_37207,N_28392,N_29213);
nand U37208 (N_37208,N_23902,N_24372);
and U37209 (N_37209,N_27435,N_23021);
nand U37210 (N_37210,N_29466,N_29479);
or U37211 (N_37211,N_22073,N_21867);
nor U37212 (N_37212,N_25407,N_26953);
nor U37213 (N_37213,N_25882,N_26044);
nand U37214 (N_37214,N_23789,N_27360);
and U37215 (N_37215,N_26897,N_27819);
nand U37216 (N_37216,N_24294,N_20033);
nor U37217 (N_37217,N_26014,N_29049);
and U37218 (N_37218,N_29042,N_21596);
nor U37219 (N_37219,N_23392,N_23329);
or U37220 (N_37220,N_20448,N_21529);
xnor U37221 (N_37221,N_26878,N_25041);
and U37222 (N_37222,N_21905,N_26377);
and U37223 (N_37223,N_21926,N_21575);
and U37224 (N_37224,N_27916,N_28863);
or U37225 (N_37225,N_24125,N_27882);
nand U37226 (N_37226,N_28262,N_26728);
nor U37227 (N_37227,N_29527,N_25221);
or U37228 (N_37228,N_24027,N_29807);
nor U37229 (N_37229,N_20213,N_28246);
nor U37230 (N_37230,N_24328,N_24013);
or U37231 (N_37231,N_27881,N_25385);
and U37232 (N_37232,N_27468,N_28840);
nor U37233 (N_37233,N_23607,N_21642);
or U37234 (N_37234,N_27134,N_25607);
nor U37235 (N_37235,N_25692,N_29722);
nand U37236 (N_37236,N_21024,N_29417);
and U37237 (N_37237,N_26219,N_24006);
nand U37238 (N_37238,N_29339,N_29444);
xor U37239 (N_37239,N_28818,N_20005);
nand U37240 (N_37240,N_23939,N_22254);
nand U37241 (N_37241,N_26377,N_22206);
and U37242 (N_37242,N_29250,N_21648);
nor U37243 (N_37243,N_25740,N_28217);
xor U37244 (N_37244,N_21755,N_22637);
and U37245 (N_37245,N_29251,N_27270);
and U37246 (N_37246,N_23337,N_20253);
nor U37247 (N_37247,N_27847,N_21478);
nor U37248 (N_37248,N_25410,N_24973);
or U37249 (N_37249,N_29032,N_24447);
nand U37250 (N_37250,N_20699,N_25063);
and U37251 (N_37251,N_25220,N_27502);
xor U37252 (N_37252,N_29988,N_27115);
xor U37253 (N_37253,N_24394,N_25706);
nor U37254 (N_37254,N_22718,N_29345);
and U37255 (N_37255,N_20449,N_29011);
nand U37256 (N_37256,N_24071,N_29933);
nand U37257 (N_37257,N_23556,N_28362);
nor U37258 (N_37258,N_26777,N_25346);
nand U37259 (N_37259,N_24300,N_25120);
nand U37260 (N_37260,N_25175,N_25270);
or U37261 (N_37261,N_25183,N_26404);
and U37262 (N_37262,N_29405,N_28948);
or U37263 (N_37263,N_27854,N_22652);
nand U37264 (N_37264,N_24193,N_26322);
and U37265 (N_37265,N_22672,N_21484);
nand U37266 (N_37266,N_21198,N_26505);
nor U37267 (N_37267,N_26327,N_22145);
and U37268 (N_37268,N_29963,N_27769);
xor U37269 (N_37269,N_22241,N_21666);
nor U37270 (N_37270,N_28114,N_24673);
or U37271 (N_37271,N_23358,N_23339);
nor U37272 (N_37272,N_28632,N_27914);
nor U37273 (N_37273,N_26769,N_22293);
nor U37274 (N_37274,N_21262,N_25411);
and U37275 (N_37275,N_29626,N_22981);
and U37276 (N_37276,N_27648,N_22657);
nor U37277 (N_37277,N_23165,N_21861);
or U37278 (N_37278,N_23328,N_27605);
and U37279 (N_37279,N_29398,N_28973);
nand U37280 (N_37280,N_29676,N_29361);
and U37281 (N_37281,N_26730,N_22633);
nand U37282 (N_37282,N_25224,N_26465);
or U37283 (N_37283,N_29480,N_23235);
xor U37284 (N_37284,N_22734,N_27356);
or U37285 (N_37285,N_21169,N_23580);
nor U37286 (N_37286,N_26094,N_20024);
or U37287 (N_37287,N_28643,N_22317);
nand U37288 (N_37288,N_22133,N_29090);
nor U37289 (N_37289,N_27474,N_29728);
nand U37290 (N_37290,N_26997,N_23114);
and U37291 (N_37291,N_21325,N_27520);
or U37292 (N_37292,N_23984,N_20280);
nand U37293 (N_37293,N_24799,N_20090);
or U37294 (N_37294,N_29427,N_22529);
nor U37295 (N_37295,N_28188,N_21840);
and U37296 (N_37296,N_26394,N_24361);
and U37297 (N_37297,N_24873,N_27672);
or U37298 (N_37298,N_24014,N_29980);
nor U37299 (N_37299,N_24966,N_24873);
nand U37300 (N_37300,N_23084,N_29064);
nand U37301 (N_37301,N_20025,N_29903);
xor U37302 (N_37302,N_27337,N_25418);
nand U37303 (N_37303,N_22915,N_28201);
and U37304 (N_37304,N_22560,N_27049);
or U37305 (N_37305,N_24598,N_28322);
or U37306 (N_37306,N_29236,N_29392);
or U37307 (N_37307,N_22358,N_25471);
or U37308 (N_37308,N_27586,N_29612);
xnor U37309 (N_37309,N_26390,N_25084);
and U37310 (N_37310,N_28159,N_23886);
or U37311 (N_37311,N_24938,N_24375);
and U37312 (N_37312,N_26012,N_24672);
xor U37313 (N_37313,N_29076,N_27578);
nor U37314 (N_37314,N_23696,N_23423);
or U37315 (N_37315,N_27967,N_24427);
nor U37316 (N_37316,N_23476,N_25395);
nand U37317 (N_37317,N_24632,N_24560);
nor U37318 (N_37318,N_21338,N_27079);
or U37319 (N_37319,N_22564,N_29207);
nand U37320 (N_37320,N_20354,N_21614);
and U37321 (N_37321,N_29123,N_26504);
xnor U37322 (N_37322,N_25835,N_29444);
nand U37323 (N_37323,N_25398,N_24614);
nor U37324 (N_37324,N_28474,N_27566);
or U37325 (N_37325,N_23172,N_29382);
nand U37326 (N_37326,N_28259,N_29430);
or U37327 (N_37327,N_28139,N_28317);
and U37328 (N_37328,N_20029,N_21467);
nand U37329 (N_37329,N_28557,N_29458);
nor U37330 (N_37330,N_26664,N_26530);
or U37331 (N_37331,N_25526,N_29452);
nand U37332 (N_37332,N_23228,N_28482);
nor U37333 (N_37333,N_24440,N_23053);
nor U37334 (N_37334,N_22748,N_22753);
and U37335 (N_37335,N_20323,N_21540);
or U37336 (N_37336,N_23587,N_27242);
or U37337 (N_37337,N_26179,N_23613);
and U37338 (N_37338,N_29578,N_22525);
nor U37339 (N_37339,N_28331,N_23060);
nand U37340 (N_37340,N_23859,N_25393);
and U37341 (N_37341,N_25478,N_28594);
nand U37342 (N_37342,N_25899,N_27508);
nand U37343 (N_37343,N_28176,N_20120);
nor U37344 (N_37344,N_28684,N_25235);
nand U37345 (N_37345,N_29009,N_28317);
nor U37346 (N_37346,N_27767,N_21850);
nand U37347 (N_37347,N_23196,N_29361);
or U37348 (N_37348,N_28687,N_25548);
nor U37349 (N_37349,N_26405,N_20135);
nor U37350 (N_37350,N_23220,N_27189);
nand U37351 (N_37351,N_22806,N_24607);
or U37352 (N_37352,N_28312,N_24461);
and U37353 (N_37353,N_20644,N_26287);
and U37354 (N_37354,N_26059,N_24596);
nand U37355 (N_37355,N_26249,N_25768);
xnor U37356 (N_37356,N_26948,N_21070);
and U37357 (N_37357,N_25520,N_26229);
nand U37358 (N_37358,N_24449,N_27930);
xnor U37359 (N_37359,N_28573,N_25071);
nand U37360 (N_37360,N_26582,N_22051);
and U37361 (N_37361,N_21425,N_22368);
or U37362 (N_37362,N_29074,N_20027);
or U37363 (N_37363,N_21159,N_23700);
nor U37364 (N_37364,N_25720,N_26456);
and U37365 (N_37365,N_27279,N_24379);
nor U37366 (N_37366,N_25827,N_22148);
xnor U37367 (N_37367,N_28865,N_28921);
nor U37368 (N_37368,N_21246,N_23676);
nor U37369 (N_37369,N_25592,N_20085);
nor U37370 (N_37370,N_27211,N_27396);
or U37371 (N_37371,N_25972,N_24242);
and U37372 (N_37372,N_24024,N_23377);
nand U37373 (N_37373,N_26756,N_27203);
xor U37374 (N_37374,N_24922,N_29787);
nand U37375 (N_37375,N_23693,N_27480);
or U37376 (N_37376,N_25673,N_22906);
nor U37377 (N_37377,N_26299,N_22728);
nand U37378 (N_37378,N_20784,N_29446);
nor U37379 (N_37379,N_26867,N_20275);
and U37380 (N_37380,N_29608,N_24975);
and U37381 (N_37381,N_20119,N_25826);
nand U37382 (N_37382,N_21069,N_26400);
nand U37383 (N_37383,N_27387,N_24058);
xor U37384 (N_37384,N_26686,N_22887);
nand U37385 (N_37385,N_27726,N_23533);
and U37386 (N_37386,N_22609,N_29831);
or U37387 (N_37387,N_29495,N_26169);
xnor U37388 (N_37388,N_25640,N_21687);
and U37389 (N_37389,N_20776,N_24581);
xnor U37390 (N_37390,N_24337,N_26975);
or U37391 (N_37391,N_29590,N_24775);
nand U37392 (N_37392,N_26399,N_27739);
or U37393 (N_37393,N_24506,N_24938);
xor U37394 (N_37394,N_20202,N_26887);
nor U37395 (N_37395,N_21486,N_27633);
or U37396 (N_37396,N_28434,N_22247);
nor U37397 (N_37397,N_24588,N_20160);
nand U37398 (N_37398,N_22509,N_27867);
and U37399 (N_37399,N_28459,N_24058);
nand U37400 (N_37400,N_23426,N_24323);
nor U37401 (N_37401,N_24824,N_23689);
nand U37402 (N_37402,N_24541,N_28852);
nand U37403 (N_37403,N_22539,N_20839);
and U37404 (N_37404,N_20184,N_20999);
or U37405 (N_37405,N_26087,N_25986);
xor U37406 (N_37406,N_25662,N_20634);
xnor U37407 (N_37407,N_25703,N_22390);
nor U37408 (N_37408,N_29455,N_29220);
and U37409 (N_37409,N_26113,N_20754);
or U37410 (N_37410,N_29067,N_24773);
xor U37411 (N_37411,N_28597,N_20847);
nand U37412 (N_37412,N_21572,N_25040);
nor U37413 (N_37413,N_27988,N_25313);
and U37414 (N_37414,N_24894,N_29465);
xor U37415 (N_37415,N_29815,N_24893);
or U37416 (N_37416,N_29983,N_21443);
and U37417 (N_37417,N_29727,N_27139);
nand U37418 (N_37418,N_29873,N_26676);
nor U37419 (N_37419,N_26751,N_22737);
or U37420 (N_37420,N_22457,N_29785);
nor U37421 (N_37421,N_23992,N_24049);
or U37422 (N_37422,N_23635,N_21002);
and U37423 (N_37423,N_22458,N_26417);
and U37424 (N_37424,N_29411,N_27100);
or U37425 (N_37425,N_22554,N_27628);
and U37426 (N_37426,N_20884,N_23216);
and U37427 (N_37427,N_27124,N_22666);
nor U37428 (N_37428,N_26800,N_21110);
xor U37429 (N_37429,N_21399,N_21548);
nand U37430 (N_37430,N_21739,N_29951);
and U37431 (N_37431,N_20050,N_23312);
nor U37432 (N_37432,N_20945,N_23999);
or U37433 (N_37433,N_29924,N_29157);
xor U37434 (N_37434,N_25942,N_20321);
xor U37435 (N_37435,N_23904,N_25001);
nand U37436 (N_37436,N_20752,N_29610);
nor U37437 (N_37437,N_26350,N_21782);
and U37438 (N_37438,N_21399,N_29554);
or U37439 (N_37439,N_27522,N_24359);
nor U37440 (N_37440,N_26270,N_22126);
xnor U37441 (N_37441,N_27673,N_24012);
nand U37442 (N_37442,N_26837,N_25809);
and U37443 (N_37443,N_23151,N_29349);
and U37444 (N_37444,N_25335,N_21020);
nand U37445 (N_37445,N_23440,N_20674);
xnor U37446 (N_37446,N_29936,N_21527);
nand U37447 (N_37447,N_24495,N_24020);
and U37448 (N_37448,N_21832,N_24643);
nand U37449 (N_37449,N_29046,N_23932);
nand U37450 (N_37450,N_27146,N_20931);
xnor U37451 (N_37451,N_29888,N_25234);
and U37452 (N_37452,N_23462,N_22795);
and U37453 (N_37453,N_26145,N_28134);
nor U37454 (N_37454,N_21362,N_25130);
nor U37455 (N_37455,N_21021,N_27905);
nor U37456 (N_37456,N_26756,N_24589);
or U37457 (N_37457,N_24880,N_24480);
or U37458 (N_37458,N_22212,N_29150);
nor U37459 (N_37459,N_22038,N_23692);
or U37460 (N_37460,N_29406,N_26436);
and U37461 (N_37461,N_29754,N_27664);
nand U37462 (N_37462,N_29142,N_25694);
nand U37463 (N_37463,N_22825,N_21824);
nand U37464 (N_37464,N_26672,N_24755);
nor U37465 (N_37465,N_20072,N_25140);
and U37466 (N_37466,N_22753,N_23028);
and U37467 (N_37467,N_23930,N_25818);
nand U37468 (N_37468,N_28405,N_20959);
nor U37469 (N_37469,N_23859,N_26229);
nor U37470 (N_37470,N_22058,N_28287);
nor U37471 (N_37471,N_23617,N_29851);
and U37472 (N_37472,N_22017,N_27683);
or U37473 (N_37473,N_22369,N_23973);
xnor U37474 (N_37474,N_22495,N_25711);
and U37475 (N_37475,N_24228,N_22019);
and U37476 (N_37476,N_20489,N_23721);
xor U37477 (N_37477,N_23838,N_27629);
nor U37478 (N_37478,N_20049,N_25316);
xnor U37479 (N_37479,N_29143,N_22726);
and U37480 (N_37480,N_26612,N_23906);
or U37481 (N_37481,N_22166,N_21601);
nand U37482 (N_37482,N_20350,N_24605);
nand U37483 (N_37483,N_28912,N_20089);
and U37484 (N_37484,N_28792,N_27703);
or U37485 (N_37485,N_21141,N_22493);
or U37486 (N_37486,N_24430,N_23046);
or U37487 (N_37487,N_28625,N_26201);
nand U37488 (N_37488,N_27067,N_29893);
nand U37489 (N_37489,N_27566,N_26187);
or U37490 (N_37490,N_28657,N_21848);
nand U37491 (N_37491,N_21567,N_23264);
nor U37492 (N_37492,N_22315,N_22998);
nor U37493 (N_37493,N_21759,N_24145);
or U37494 (N_37494,N_25553,N_24467);
and U37495 (N_37495,N_25675,N_20078);
and U37496 (N_37496,N_22979,N_26821);
nand U37497 (N_37497,N_26980,N_22794);
xor U37498 (N_37498,N_28733,N_23221);
and U37499 (N_37499,N_22890,N_25096);
or U37500 (N_37500,N_26918,N_27059);
or U37501 (N_37501,N_29742,N_22988);
xor U37502 (N_37502,N_23695,N_28978);
or U37503 (N_37503,N_23369,N_21246);
nand U37504 (N_37504,N_20085,N_26551);
and U37505 (N_37505,N_22381,N_25015);
nor U37506 (N_37506,N_27812,N_24604);
nand U37507 (N_37507,N_21742,N_29849);
nor U37508 (N_37508,N_29245,N_28235);
nor U37509 (N_37509,N_22687,N_21154);
or U37510 (N_37510,N_27432,N_21017);
nor U37511 (N_37511,N_23358,N_23067);
nand U37512 (N_37512,N_27293,N_21504);
or U37513 (N_37513,N_27572,N_25921);
and U37514 (N_37514,N_29014,N_26734);
and U37515 (N_37515,N_20153,N_29583);
and U37516 (N_37516,N_21799,N_29509);
nand U37517 (N_37517,N_20020,N_23780);
nor U37518 (N_37518,N_20404,N_25940);
nand U37519 (N_37519,N_20339,N_21876);
or U37520 (N_37520,N_20889,N_24698);
and U37521 (N_37521,N_29100,N_23793);
nand U37522 (N_37522,N_24169,N_23577);
nor U37523 (N_37523,N_22346,N_29887);
or U37524 (N_37524,N_23290,N_20908);
nor U37525 (N_37525,N_25810,N_24011);
nand U37526 (N_37526,N_22248,N_20201);
nor U37527 (N_37527,N_22796,N_25393);
nand U37528 (N_37528,N_25779,N_23271);
or U37529 (N_37529,N_22317,N_21424);
nor U37530 (N_37530,N_22598,N_27708);
nand U37531 (N_37531,N_22130,N_27237);
or U37532 (N_37532,N_23945,N_23806);
or U37533 (N_37533,N_29254,N_24778);
nor U37534 (N_37534,N_26259,N_28322);
nand U37535 (N_37535,N_24350,N_28228);
nand U37536 (N_37536,N_25801,N_22659);
or U37537 (N_37537,N_21873,N_21601);
or U37538 (N_37538,N_24593,N_20577);
nand U37539 (N_37539,N_24374,N_21134);
or U37540 (N_37540,N_21874,N_22342);
nand U37541 (N_37541,N_22666,N_22214);
xnor U37542 (N_37542,N_27883,N_22456);
nand U37543 (N_37543,N_20521,N_23451);
nor U37544 (N_37544,N_28847,N_24831);
xor U37545 (N_37545,N_27896,N_23259);
nand U37546 (N_37546,N_22268,N_24177);
and U37547 (N_37547,N_28522,N_26589);
and U37548 (N_37548,N_25523,N_29126);
xnor U37549 (N_37549,N_28682,N_27621);
xnor U37550 (N_37550,N_23512,N_26442);
and U37551 (N_37551,N_24066,N_26751);
or U37552 (N_37552,N_25757,N_29187);
nand U37553 (N_37553,N_29948,N_20953);
and U37554 (N_37554,N_27280,N_24360);
and U37555 (N_37555,N_23625,N_21746);
xnor U37556 (N_37556,N_22591,N_22208);
or U37557 (N_37557,N_22295,N_20860);
nand U37558 (N_37558,N_26425,N_20961);
nand U37559 (N_37559,N_27924,N_28801);
nor U37560 (N_37560,N_21523,N_24454);
and U37561 (N_37561,N_26264,N_27398);
and U37562 (N_37562,N_22494,N_22394);
and U37563 (N_37563,N_22273,N_20471);
nor U37564 (N_37564,N_23602,N_28906);
nor U37565 (N_37565,N_24035,N_24361);
xnor U37566 (N_37566,N_26792,N_21029);
and U37567 (N_37567,N_28341,N_21860);
nand U37568 (N_37568,N_22348,N_28958);
nand U37569 (N_37569,N_26453,N_25353);
nand U37570 (N_37570,N_23421,N_22732);
or U37571 (N_37571,N_27896,N_21429);
and U37572 (N_37572,N_21453,N_29406);
and U37573 (N_37573,N_21150,N_21458);
nand U37574 (N_37574,N_23339,N_23744);
nor U37575 (N_37575,N_26396,N_27923);
nand U37576 (N_37576,N_20120,N_28035);
or U37577 (N_37577,N_27724,N_22741);
nand U37578 (N_37578,N_20567,N_25835);
or U37579 (N_37579,N_27744,N_22836);
nand U37580 (N_37580,N_27707,N_22216);
nand U37581 (N_37581,N_23548,N_20392);
and U37582 (N_37582,N_29554,N_24153);
nand U37583 (N_37583,N_24911,N_26438);
and U37584 (N_37584,N_27770,N_22827);
xnor U37585 (N_37585,N_24747,N_29064);
xnor U37586 (N_37586,N_24632,N_25521);
or U37587 (N_37587,N_21409,N_25111);
and U37588 (N_37588,N_20818,N_20452);
or U37589 (N_37589,N_25995,N_20258);
or U37590 (N_37590,N_22266,N_29117);
or U37591 (N_37591,N_26847,N_27512);
nor U37592 (N_37592,N_21268,N_25736);
and U37593 (N_37593,N_21970,N_27838);
nor U37594 (N_37594,N_28432,N_24973);
nand U37595 (N_37595,N_20246,N_22779);
or U37596 (N_37596,N_25071,N_22424);
or U37597 (N_37597,N_22678,N_28754);
nand U37598 (N_37598,N_26512,N_23862);
or U37599 (N_37599,N_22427,N_28735);
xnor U37600 (N_37600,N_27334,N_27596);
and U37601 (N_37601,N_28790,N_27620);
or U37602 (N_37602,N_25746,N_29734);
nand U37603 (N_37603,N_20494,N_25434);
nand U37604 (N_37604,N_24731,N_27070);
and U37605 (N_37605,N_22986,N_26682);
xor U37606 (N_37606,N_29486,N_26744);
xor U37607 (N_37607,N_27052,N_23277);
nand U37608 (N_37608,N_22134,N_27912);
and U37609 (N_37609,N_24190,N_29939);
nand U37610 (N_37610,N_20740,N_23488);
and U37611 (N_37611,N_29765,N_26890);
xnor U37612 (N_37612,N_23193,N_23561);
xnor U37613 (N_37613,N_24261,N_20515);
nor U37614 (N_37614,N_20576,N_23643);
nand U37615 (N_37615,N_20721,N_28132);
nand U37616 (N_37616,N_25418,N_27463);
or U37617 (N_37617,N_21075,N_23603);
nand U37618 (N_37618,N_26101,N_24230);
nand U37619 (N_37619,N_25030,N_27537);
nor U37620 (N_37620,N_24052,N_29062);
nand U37621 (N_37621,N_28172,N_29099);
nor U37622 (N_37622,N_27248,N_21842);
or U37623 (N_37623,N_29169,N_24767);
xor U37624 (N_37624,N_21401,N_20532);
nor U37625 (N_37625,N_22040,N_24936);
and U37626 (N_37626,N_25285,N_24699);
or U37627 (N_37627,N_20279,N_26570);
or U37628 (N_37628,N_29834,N_27600);
and U37629 (N_37629,N_29911,N_24326);
xnor U37630 (N_37630,N_24839,N_29251);
and U37631 (N_37631,N_20620,N_24511);
xor U37632 (N_37632,N_27944,N_27984);
or U37633 (N_37633,N_25638,N_28441);
and U37634 (N_37634,N_22111,N_28656);
and U37635 (N_37635,N_21910,N_24960);
nand U37636 (N_37636,N_22890,N_28312);
xnor U37637 (N_37637,N_25619,N_25213);
and U37638 (N_37638,N_28754,N_20523);
xnor U37639 (N_37639,N_20633,N_28669);
xnor U37640 (N_37640,N_28551,N_21370);
or U37641 (N_37641,N_20310,N_27883);
nor U37642 (N_37642,N_27086,N_21784);
xor U37643 (N_37643,N_26097,N_24497);
and U37644 (N_37644,N_23206,N_28712);
nand U37645 (N_37645,N_25926,N_23859);
nor U37646 (N_37646,N_24239,N_24889);
or U37647 (N_37647,N_27985,N_27317);
or U37648 (N_37648,N_20253,N_29423);
nor U37649 (N_37649,N_25143,N_25529);
nand U37650 (N_37650,N_22907,N_21703);
nand U37651 (N_37651,N_25264,N_24654);
nor U37652 (N_37652,N_21283,N_20492);
nand U37653 (N_37653,N_29582,N_23262);
nand U37654 (N_37654,N_22254,N_23744);
nor U37655 (N_37655,N_24338,N_24743);
nor U37656 (N_37656,N_22586,N_21481);
and U37657 (N_37657,N_27578,N_25201);
xor U37658 (N_37658,N_26911,N_23973);
xor U37659 (N_37659,N_26712,N_25418);
nand U37660 (N_37660,N_24684,N_27614);
nand U37661 (N_37661,N_28942,N_24436);
and U37662 (N_37662,N_20729,N_24210);
or U37663 (N_37663,N_27230,N_24027);
nor U37664 (N_37664,N_22537,N_27784);
or U37665 (N_37665,N_24815,N_22250);
and U37666 (N_37666,N_28467,N_28266);
nand U37667 (N_37667,N_28613,N_27648);
and U37668 (N_37668,N_22167,N_20061);
or U37669 (N_37669,N_27675,N_23835);
or U37670 (N_37670,N_25750,N_20804);
or U37671 (N_37671,N_26697,N_21153);
or U37672 (N_37672,N_20037,N_23325);
or U37673 (N_37673,N_27119,N_24073);
or U37674 (N_37674,N_22085,N_24763);
nand U37675 (N_37675,N_29041,N_27865);
and U37676 (N_37676,N_28361,N_28682);
and U37677 (N_37677,N_25391,N_24640);
or U37678 (N_37678,N_25076,N_26376);
nand U37679 (N_37679,N_28568,N_28555);
or U37680 (N_37680,N_23428,N_20201);
nor U37681 (N_37681,N_24583,N_28121);
or U37682 (N_37682,N_25250,N_23640);
nor U37683 (N_37683,N_28078,N_28784);
nor U37684 (N_37684,N_22257,N_27096);
or U37685 (N_37685,N_21658,N_23858);
or U37686 (N_37686,N_26518,N_28951);
nor U37687 (N_37687,N_27914,N_23929);
and U37688 (N_37688,N_27426,N_24052);
nor U37689 (N_37689,N_20152,N_20620);
or U37690 (N_37690,N_23545,N_23593);
and U37691 (N_37691,N_24376,N_26830);
nand U37692 (N_37692,N_24854,N_21457);
xor U37693 (N_37693,N_29059,N_28024);
and U37694 (N_37694,N_25012,N_29200);
nand U37695 (N_37695,N_24071,N_23925);
xnor U37696 (N_37696,N_29424,N_26475);
xnor U37697 (N_37697,N_25106,N_20664);
xnor U37698 (N_37698,N_22392,N_23908);
nor U37699 (N_37699,N_28997,N_24800);
nand U37700 (N_37700,N_24996,N_25469);
nand U37701 (N_37701,N_24566,N_26795);
or U37702 (N_37702,N_20425,N_24402);
nor U37703 (N_37703,N_27411,N_24241);
nor U37704 (N_37704,N_26182,N_28499);
or U37705 (N_37705,N_25414,N_22926);
or U37706 (N_37706,N_28302,N_29666);
or U37707 (N_37707,N_29506,N_22339);
nand U37708 (N_37708,N_24677,N_28595);
or U37709 (N_37709,N_27769,N_22112);
nor U37710 (N_37710,N_25119,N_24489);
or U37711 (N_37711,N_23771,N_23720);
and U37712 (N_37712,N_25503,N_21452);
or U37713 (N_37713,N_26128,N_24585);
nand U37714 (N_37714,N_26147,N_20225);
and U37715 (N_37715,N_20092,N_26908);
and U37716 (N_37716,N_28810,N_28061);
xor U37717 (N_37717,N_25637,N_25458);
nand U37718 (N_37718,N_25200,N_22474);
nand U37719 (N_37719,N_25558,N_29094);
or U37720 (N_37720,N_25261,N_21324);
xnor U37721 (N_37721,N_22121,N_21517);
and U37722 (N_37722,N_28770,N_25200);
and U37723 (N_37723,N_23562,N_22220);
nor U37724 (N_37724,N_26339,N_20441);
and U37725 (N_37725,N_23534,N_26662);
nand U37726 (N_37726,N_24428,N_26501);
nor U37727 (N_37727,N_29228,N_22205);
xor U37728 (N_37728,N_26953,N_26349);
and U37729 (N_37729,N_26986,N_24307);
nand U37730 (N_37730,N_21354,N_27492);
nand U37731 (N_37731,N_23034,N_29491);
nor U37732 (N_37732,N_25374,N_22177);
and U37733 (N_37733,N_28494,N_24456);
nor U37734 (N_37734,N_27881,N_28537);
and U37735 (N_37735,N_22344,N_28024);
nand U37736 (N_37736,N_29975,N_25787);
nand U37737 (N_37737,N_24947,N_27419);
nor U37738 (N_37738,N_29759,N_27932);
and U37739 (N_37739,N_28903,N_20047);
nor U37740 (N_37740,N_23191,N_23231);
and U37741 (N_37741,N_28962,N_21534);
and U37742 (N_37742,N_20915,N_20448);
and U37743 (N_37743,N_26999,N_26637);
nand U37744 (N_37744,N_27518,N_21166);
xnor U37745 (N_37745,N_24167,N_25578);
xnor U37746 (N_37746,N_21144,N_26441);
nor U37747 (N_37747,N_23775,N_25895);
or U37748 (N_37748,N_23353,N_25528);
or U37749 (N_37749,N_29155,N_22634);
nor U37750 (N_37750,N_27891,N_29994);
or U37751 (N_37751,N_23533,N_22804);
nand U37752 (N_37752,N_20985,N_29436);
or U37753 (N_37753,N_28700,N_28040);
nand U37754 (N_37754,N_26306,N_24573);
nand U37755 (N_37755,N_23288,N_27391);
nand U37756 (N_37756,N_26678,N_26844);
nand U37757 (N_37757,N_24410,N_21190);
or U37758 (N_37758,N_23409,N_20016);
xor U37759 (N_37759,N_29162,N_23818);
nor U37760 (N_37760,N_28946,N_20344);
nor U37761 (N_37761,N_24303,N_26873);
or U37762 (N_37762,N_28503,N_20697);
xnor U37763 (N_37763,N_29362,N_21493);
nor U37764 (N_37764,N_21118,N_27371);
nor U37765 (N_37765,N_26314,N_28578);
and U37766 (N_37766,N_23877,N_25759);
xor U37767 (N_37767,N_20724,N_22355);
nand U37768 (N_37768,N_21159,N_29381);
nor U37769 (N_37769,N_20930,N_23074);
nand U37770 (N_37770,N_23108,N_20445);
or U37771 (N_37771,N_24715,N_21029);
nand U37772 (N_37772,N_24691,N_23439);
nor U37773 (N_37773,N_24188,N_27397);
and U37774 (N_37774,N_21504,N_22047);
and U37775 (N_37775,N_28223,N_29681);
nor U37776 (N_37776,N_29499,N_20737);
nand U37777 (N_37777,N_23544,N_25783);
or U37778 (N_37778,N_23239,N_27779);
or U37779 (N_37779,N_25930,N_22412);
or U37780 (N_37780,N_20662,N_29445);
nand U37781 (N_37781,N_29324,N_25298);
nand U37782 (N_37782,N_24209,N_20304);
and U37783 (N_37783,N_28034,N_23174);
nand U37784 (N_37784,N_28753,N_24858);
nand U37785 (N_37785,N_24649,N_20623);
nor U37786 (N_37786,N_28490,N_25798);
nor U37787 (N_37787,N_28937,N_22637);
nand U37788 (N_37788,N_25829,N_20483);
nor U37789 (N_37789,N_24842,N_29389);
nand U37790 (N_37790,N_28983,N_23400);
or U37791 (N_37791,N_23351,N_24502);
nor U37792 (N_37792,N_27628,N_23545);
or U37793 (N_37793,N_25762,N_24793);
and U37794 (N_37794,N_29277,N_28224);
nor U37795 (N_37795,N_27162,N_23692);
nor U37796 (N_37796,N_20937,N_20317);
nand U37797 (N_37797,N_26052,N_22506);
or U37798 (N_37798,N_22820,N_23626);
nand U37799 (N_37799,N_21239,N_28611);
nor U37800 (N_37800,N_26807,N_28975);
nand U37801 (N_37801,N_29268,N_27835);
and U37802 (N_37802,N_29786,N_22935);
or U37803 (N_37803,N_20602,N_29551);
nor U37804 (N_37804,N_23835,N_24933);
or U37805 (N_37805,N_29811,N_23935);
nor U37806 (N_37806,N_26366,N_25500);
nor U37807 (N_37807,N_24560,N_20291);
or U37808 (N_37808,N_28065,N_25766);
nand U37809 (N_37809,N_25812,N_21504);
nor U37810 (N_37810,N_29984,N_24962);
or U37811 (N_37811,N_29335,N_27969);
and U37812 (N_37812,N_29495,N_23898);
nand U37813 (N_37813,N_26434,N_28077);
nand U37814 (N_37814,N_22526,N_22278);
and U37815 (N_37815,N_29715,N_28332);
or U37816 (N_37816,N_27469,N_28250);
nor U37817 (N_37817,N_27628,N_27349);
nor U37818 (N_37818,N_25328,N_26439);
nand U37819 (N_37819,N_29374,N_21912);
or U37820 (N_37820,N_27188,N_21384);
nand U37821 (N_37821,N_20612,N_27328);
nor U37822 (N_37822,N_26523,N_27095);
and U37823 (N_37823,N_29602,N_29269);
or U37824 (N_37824,N_21069,N_20535);
nor U37825 (N_37825,N_24609,N_21973);
and U37826 (N_37826,N_21550,N_22354);
nand U37827 (N_37827,N_29045,N_29411);
and U37828 (N_37828,N_25415,N_22572);
nand U37829 (N_37829,N_29856,N_21411);
or U37830 (N_37830,N_25378,N_29785);
nand U37831 (N_37831,N_28083,N_24020);
nor U37832 (N_37832,N_21401,N_28518);
nand U37833 (N_37833,N_20556,N_22222);
nand U37834 (N_37834,N_20796,N_29699);
nand U37835 (N_37835,N_28940,N_20768);
and U37836 (N_37836,N_22113,N_22402);
nor U37837 (N_37837,N_24638,N_28783);
nor U37838 (N_37838,N_23032,N_28803);
or U37839 (N_37839,N_22034,N_23809);
or U37840 (N_37840,N_26665,N_21479);
or U37841 (N_37841,N_22398,N_24365);
nand U37842 (N_37842,N_24016,N_21301);
xor U37843 (N_37843,N_28065,N_23477);
nand U37844 (N_37844,N_20295,N_21612);
and U37845 (N_37845,N_28322,N_25911);
or U37846 (N_37846,N_24326,N_25396);
nand U37847 (N_37847,N_23275,N_25266);
xor U37848 (N_37848,N_25089,N_23489);
nand U37849 (N_37849,N_22691,N_23329);
or U37850 (N_37850,N_22381,N_22249);
nand U37851 (N_37851,N_21161,N_21670);
nor U37852 (N_37852,N_25508,N_24105);
nand U37853 (N_37853,N_28734,N_24845);
or U37854 (N_37854,N_22574,N_28584);
or U37855 (N_37855,N_27018,N_29932);
or U37856 (N_37856,N_22561,N_20043);
nand U37857 (N_37857,N_21435,N_25478);
or U37858 (N_37858,N_26381,N_25185);
nand U37859 (N_37859,N_29774,N_21477);
or U37860 (N_37860,N_21469,N_28666);
xor U37861 (N_37861,N_29359,N_23289);
nor U37862 (N_37862,N_25437,N_22004);
nand U37863 (N_37863,N_28002,N_26164);
and U37864 (N_37864,N_29392,N_23521);
and U37865 (N_37865,N_20359,N_22422);
nor U37866 (N_37866,N_22836,N_29984);
xnor U37867 (N_37867,N_25905,N_29708);
or U37868 (N_37868,N_27560,N_25303);
nor U37869 (N_37869,N_24663,N_24594);
nor U37870 (N_37870,N_27957,N_29778);
xor U37871 (N_37871,N_22162,N_21311);
or U37872 (N_37872,N_23667,N_21596);
nand U37873 (N_37873,N_29712,N_25485);
xnor U37874 (N_37874,N_27480,N_22026);
or U37875 (N_37875,N_28195,N_22472);
nor U37876 (N_37876,N_23801,N_20195);
and U37877 (N_37877,N_20210,N_27286);
nand U37878 (N_37878,N_22411,N_24624);
nand U37879 (N_37879,N_22792,N_28777);
and U37880 (N_37880,N_28971,N_21282);
nor U37881 (N_37881,N_27768,N_27829);
or U37882 (N_37882,N_29556,N_27437);
nor U37883 (N_37883,N_27791,N_21986);
nand U37884 (N_37884,N_20631,N_20893);
or U37885 (N_37885,N_28299,N_28790);
or U37886 (N_37886,N_20086,N_20096);
and U37887 (N_37887,N_27690,N_21786);
or U37888 (N_37888,N_21480,N_25443);
or U37889 (N_37889,N_27587,N_22804);
nor U37890 (N_37890,N_29895,N_21753);
or U37891 (N_37891,N_24253,N_25527);
or U37892 (N_37892,N_29106,N_22288);
nand U37893 (N_37893,N_25815,N_28311);
nand U37894 (N_37894,N_22203,N_23566);
or U37895 (N_37895,N_20720,N_21425);
or U37896 (N_37896,N_26271,N_27690);
and U37897 (N_37897,N_20136,N_25250);
xnor U37898 (N_37898,N_26564,N_27167);
nand U37899 (N_37899,N_27100,N_26742);
nor U37900 (N_37900,N_23910,N_28150);
or U37901 (N_37901,N_27982,N_25036);
nor U37902 (N_37902,N_24820,N_21104);
nor U37903 (N_37903,N_22401,N_22943);
or U37904 (N_37904,N_29803,N_24569);
and U37905 (N_37905,N_26649,N_20664);
or U37906 (N_37906,N_27869,N_21275);
or U37907 (N_37907,N_23261,N_20435);
nor U37908 (N_37908,N_25805,N_21177);
or U37909 (N_37909,N_24716,N_28869);
nand U37910 (N_37910,N_25736,N_26387);
or U37911 (N_37911,N_29090,N_27897);
nand U37912 (N_37912,N_26806,N_26503);
and U37913 (N_37913,N_21595,N_23846);
and U37914 (N_37914,N_28826,N_22363);
nor U37915 (N_37915,N_28247,N_25279);
and U37916 (N_37916,N_26049,N_27819);
xor U37917 (N_37917,N_29810,N_25239);
or U37918 (N_37918,N_25181,N_25966);
and U37919 (N_37919,N_22334,N_23461);
nor U37920 (N_37920,N_25168,N_24489);
nand U37921 (N_37921,N_28374,N_23012);
nor U37922 (N_37922,N_28846,N_25987);
xor U37923 (N_37923,N_24051,N_27923);
nand U37924 (N_37924,N_24698,N_23753);
xor U37925 (N_37925,N_28182,N_28128);
nor U37926 (N_37926,N_27849,N_26774);
or U37927 (N_37927,N_24510,N_24173);
and U37928 (N_37928,N_24574,N_22116);
or U37929 (N_37929,N_29757,N_25773);
or U37930 (N_37930,N_23345,N_21121);
and U37931 (N_37931,N_22596,N_25555);
xor U37932 (N_37932,N_24858,N_27744);
nor U37933 (N_37933,N_22856,N_28123);
nor U37934 (N_37934,N_29140,N_23714);
nor U37935 (N_37935,N_22271,N_22154);
xor U37936 (N_37936,N_27982,N_20302);
xnor U37937 (N_37937,N_20520,N_25586);
and U37938 (N_37938,N_27010,N_29357);
nor U37939 (N_37939,N_20406,N_27962);
nand U37940 (N_37940,N_29165,N_22095);
nor U37941 (N_37941,N_20679,N_27884);
or U37942 (N_37942,N_23548,N_20506);
nor U37943 (N_37943,N_29879,N_21709);
nand U37944 (N_37944,N_21173,N_29883);
xnor U37945 (N_37945,N_27086,N_20516);
nor U37946 (N_37946,N_23700,N_27958);
nor U37947 (N_37947,N_22759,N_21432);
or U37948 (N_37948,N_21326,N_22129);
nor U37949 (N_37949,N_24581,N_21194);
or U37950 (N_37950,N_24682,N_22161);
nand U37951 (N_37951,N_22165,N_21208);
or U37952 (N_37952,N_24602,N_23740);
nand U37953 (N_37953,N_24799,N_21398);
nand U37954 (N_37954,N_26932,N_20963);
xnor U37955 (N_37955,N_20654,N_22749);
and U37956 (N_37956,N_24541,N_22938);
nor U37957 (N_37957,N_24192,N_27666);
nand U37958 (N_37958,N_29580,N_28985);
or U37959 (N_37959,N_20369,N_29577);
or U37960 (N_37960,N_21058,N_29365);
nor U37961 (N_37961,N_28062,N_25234);
or U37962 (N_37962,N_20921,N_29222);
or U37963 (N_37963,N_27905,N_23772);
and U37964 (N_37964,N_23898,N_28435);
nand U37965 (N_37965,N_23191,N_21777);
nor U37966 (N_37966,N_29532,N_22011);
nand U37967 (N_37967,N_21349,N_29260);
nor U37968 (N_37968,N_21401,N_21358);
or U37969 (N_37969,N_21321,N_23495);
nand U37970 (N_37970,N_20075,N_28744);
nand U37971 (N_37971,N_20812,N_21475);
or U37972 (N_37972,N_29721,N_24274);
and U37973 (N_37973,N_28893,N_21870);
and U37974 (N_37974,N_29082,N_24136);
and U37975 (N_37975,N_26775,N_26580);
or U37976 (N_37976,N_20172,N_21139);
or U37977 (N_37977,N_28325,N_28309);
or U37978 (N_37978,N_27359,N_27499);
nand U37979 (N_37979,N_23778,N_26545);
nand U37980 (N_37980,N_24872,N_26123);
and U37981 (N_37981,N_25410,N_22464);
nand U37982 (N_37982,N_26413,N_26312);
nor U37983 (N_37983,N_25305,N_20713);
nand U37984 (N_37984,N_26298,N_25950);
and U37985 (N_37985,N_24419,N_27174);
or U37986 (N_37986,N_29868,N_24585);
nand U37987 (N_37987,N_21454,N_24190);
and U37988 (N_37988,N_20177,N_27183);
xnor U37989 (N_37989,N_26111,N_28296);
nand U37990 (N_37990,N_20692,N_29421);
xor U37991 (N_37991,N_25863,N_21101);
nand U37992 (N_37992,N_25550,N_28441);
and U37993 (N_37993,N_21865,N_23766);
or U37994 (N_37994,N_20283,N_24244);
or U37995 (N_37995,N_29541,N_25654);
or U37996 (N_37996,N_26248,N_29119);
nor U37997 (N_37997,N_24033,N_21902);
and U37998 (N_37998,N_23086,N_28903);
or U37999 (N_37999,N_27910,N_23218);
and U38000 (N_38000,N_22380,N_24113);
nand U38001 (N_38001,N_23132,N_29493);
and U38002 (N_38002,N_26256,N_23525);
or U38003 (N_38003,N_26990,N_23402);
and U38004 (N_38004,N_23310,N_22937);
nand U38005 (N_38005,N_24527,N_23217);
and U38006 (N_38006,N_23076,N_26364);
or U38007 (N_38007,N_23628,N_23932);
nand U38008 (N_38008,N_28098,N_29567);
nor U38009 (N_38009,N_25566,N_22296);
or U38010 (N_38010,N_26026,N_23190);
xor U38011 (N_38011,N_23279,N_29310);
nand U38012 (N_38012,N_23821,N_20643);
or U38013 (N_38013,N_20319,N_24240);
nor U38014 (N_38014,N_21583,N_24638);
or U38015 (N_38015,N_25553,N_27331);
nor U38016 (N_38016,N_27615,N_22444);
and U38017 (N_38017,N_29793,N_20820);
and U38018 (N_38018,N_24345,N_22988);
nand U38019 (N_38019,N_29943,N_25750);
and U38020 (N_38020,N_27686,N_26296);
nor U38021 (N_38021,N_26028,N_27204);
nor U38022 (N_38022,N_28867,N_28667);
and U38023 (N_38023,N_29817,N_29747);
nor U38024 (N_38024,N_28610,N_23596);
nand U38025 (N_38025,N_23615,N_20298);
and U38026 (N_38026,N_28559,N_25808);
nor U38027 (N_38027,N_26850,N_22268);
nor U38028 (N_38028,N_23366,N_20624);
nand U38029 (N_38029,N_25555,N_21068);
and U38030 (N_38030,N_20097,N_22252);
or U38031 (N_38031,N_21785,N_22160);
and U38032 (N_38032,N_26443,N_25507);
xnor U38033 (N_38033,N_26646,N_24898);
nor U38034 (N_38034,N_29067,N_21280);
and U38035 (N_38035,N_24781,N_20525);
nand U38036 (N_38036,N_24008,N_26301);
nor U38037 (N_38037,N_25953,N_22804);
xor U38038 (N_38038,N_22356,N_23123);
nand U38039 (N_38039,N_21175,N_23541);
nor U38040 (N_38040,N_23099,N_29065);
nand U38041 (N_38041,N_25332,N_24650);
nor U38042 (N_38042,N_29776,N_21486);
xnor U38043 (N_38043,N_27778,N_26712);
and U38044 (N_38044,N_22634,N_27669);
or U38045 (N_38045,N_29243,N_25816);
nand U38046 (N_38046,N_25259,N_26026);
and U38047 (N_38047,N_25422,N_26253);
nor U38048 (N_38048,N_25713,N_29221);
and U38049 (N_38049,N_20606,N_29407);
or U38050 (N_38050,N_29123,N_20722);
and U38051 (N_38051,N_21037,N_26414);
and U38052 (N_38052,N_25076,N_23743);
or U38053 (N_38053,N_28176,N_20480);
or U38054 (N_38054,N_22849,N_27374);
nor U38055 (N_38055,N_22198,N_24828);
nand U38056 (N_38056,N_24275,N_24226);
and U38057 (N_38057,N_20848,N_26927);
nor U38058 (N_38058,N_29174,N_23266);
xor U38059 (N_38059,N_23242,N_29659);
xor U38060 (N_38060,N_27085,N_24957);
or U38061 (N_38061,N_27390,N_23742);
or U38062 (N_38062,N_29273,N_22396);
and U38063 (N_38063,N_22183,N_29998);
xnor U38064 (N_38064,N_28141,N_29186);
nand U38065 (N_38065,N_20247,N_21687);
nand U38066 (N_38066,N_20762,N_28622);
nand U38067 (N_38067,N_20978,N_28011);
nor U38068 (N_38068,N_26170,N_20801);
or U38069 (N_38069,N_26689,N_24058);
nor U38070 (N_38070,N_23533,N_27742);
or U38071 (N_38071,N_26011,N_27170);
nand U38072 (N_38072,N_20036,N_25964);
and U38073 (N_38073,N_27238,N_27191);
nand U38074 (N_38074,N_27993,N_29658);
nor U38075 (N_38075,N_22208,N_23057);
nand U38076 (N_38076,N_20676,N_23236);
nand U38077 (N_38077,N_20908,N_23376);
or U38078 (N_38078,N_21842,N_28363);
xnor U38079 (N_38079,N_24086,N_27909);
or U38080 (N_38080,N_25044,N_23099);
or U38081 (N_38081,N_24813,N_22494);
xnor U38082 (N_38082,N_28995,N_21950);
and U38083 (N_38083,N_26229,N_25746);
nand U38084 (N_38084,N_22140,N_22157);
nor U38085 (N_38085,N_22823,N_28310);
nand U38086 (N_38086,N_22446,N_26257);
nand U38087 (N_38087,N_28109,N_21819);
nor U38088 (N_38088,N_20204,N_29955);
or U38089 (N_38089,N_20578,N_24939);
or U38090 (N_38090,N_27074,N_21785);
or U38091 (N_38091,N_20054,N_29943);
nand U38092 (N_38092,N_25686,N_22499);
nand U38093 (N_38093,N_29762,N_23014);
and U38094 (N_38094,N_21109,N_24080);
xor U38095 (N_38095,N_20743,N_26076);
or U38096 (N_38096,N_28548,N_28141);
nand U38097 (N_38097,N_28315,N_28336);
nand U38098 (N_38098,N_29241,N_26400);
or U38099 (N_38099,N_26964,N_21774);
and U38100 (N_38100,N_22956,N_26614);
or U38101 (N_38101,N_29350,N_22536);
or U38102 (N_38102,N_22072,N_28779);
nand U38103 (N_38103,N_29378,N_27482);
and U38104 (N_38104,N_20393,N_22217);
or U38105 (N_38105,N_28657,N_27369);
nand U38106 (N_38106,N_24929,N_22506);
nand U38107 (N_38107,N_21629,N_20272);
nor U38108 (N_38108,N_20445,N_22042);
and U38109 (N_38109,N_21757,N_26344);
and U38110 (N_38110,N_22019,N_26280);
or U38111 (N_38111,N_27128,N_28878);
or U38112 (N_38112,N_24304,N_22884);
nand U38113 (N_38113,N_25316,N_21283);
nor U38114 (N_38114,N_28511,N_28651);
nand U38115 (N_38115,N_29864,N_21535);
nand U38116 (N_38116,N_27792,N_25512);
or U38117 (N_38117,N_21427,N_26527);
xnor U38118 (N_38118,N_20560,N_20043);
nor U38119 (N_38119,N_29633,N_21709);
nand U38120 (N_38120,N_22493,N_22097);
or U38121 (N_38121,N_25935,N_21908);
nor U38122 (N_38122,N_29788,N_27201);
nand U38123 (N_38123,N_25828,N_26711);
xnor U38124 (N_38124,N_26438,N_21610);
nor U38125 (N_38125,N_21634,N_22461);
xor U38126 (N_38126,N_23074,N_26533);
nand U38127 (N_38127,N_29555,N_27899);
nor U38128 (N_38128,N_23066,N_28933);
nand U38129 (N_38129,N_26165,N_22093);
and U38130 (N_38130,N_26303,N_22354);
nor U38131 (N_38131,N_21444,N_20392);
nor U38132 (N_38132,N_22750,N_23417);
and U38133 (N_38133,N_25732,N_25286);
nand U38134 (N_38134,N_29433,N_24379);
or U38135 (N_38135,N_24640,N_28843);
and U38136 (N_38136,N_22684,N_29472);
nor U38137 (N_38137,N_24999,N_28844);
nand U38138 (N_38138,N_28527,N_24928);
or U38139 (N_38139,N_24775,N_20720);
nand U38140 (N_38140,N_28612,N_29928);
nand U38141 (N_38141,N_21169,N_21482);
nor U38142 (N_38142,N_22861,N_21097);
nand U38143 (N_38143,N_27787,N_21733);
nor U38144 (N_38144,N_25495,N_21042);
and U38145 (N_38145,N_28909,N_29215);
and U38146 (N_38146,N_28143,N_21533);
xor U38147 (N_38147,N_23676,N_25764);
and U38148 (N_38148,N_22136,N_28955);
xor U38149 (N_38149,N_21709,N_24697);
xnor U38150 (N_38150,N_26571,N_27636);
nor U38151 (N_38151,N_23517,N_25862);
nand U38152 (N_38152,N_23889,N_25785);
and U38153 (N_38153,N_20370,N_28874);
or U38154 (N_38154,N_21551,N_20770);
nand U38155 (N_38155,N_27511,N_24028);
xor U38156 (N_38156,N_24934,N_29515);
nor U38157 (N_38157,N_27390,N_25945);
or U38158 (N_38158,N_24520,N_20262);
or U38159 (N_38159,N_20840,N_29507);
nor U38160 (N_38160,N_20931,N_29934);
or U38161 (N_38161,N_23826,N_22583);
or U38162 (N_38162,N_28426,N_27286);
and U38163 (N_38163,N_23459,N_25412);
nand U38164 (N_38164,N_27473,N_22887);
and U38165 (N_38165,N_29246,N_21660);
and U38166 (N_38166,N_22720,N_29764);
nand U38167 (N_38167,N_27588,N_21083);
nor U38168 (N_38168,N_29057,N_28409);
and U38169 (N_38169,N_21853,N_28722);
xnor U38170 (N_38170,N_25539,N_22794);
and U38171 (N_38171,N_22520,N_25957);
nand U38172 (N_38172,N_29790,N_22587);
nand U38173 (N_38173,N_26276,N_29300);
xnor U38174 (N_38174,N_28647,N_20885);
nand U38175 (N_38175,N_25930,N_23208);
nor U38176 (N_38176,N_29827,N_20127);
nand U38177 (N_38177,N_24244,N_20545);
or U38178 (N_38178,N_20644,N_20212);
nand U38179 (N_38179,N_24191,N_29615);
nand U38180 (N_38180,N_21213,N_26929);
nand U38181 (N_38181,N_28161,N_26818);
xnor U38182 (N_38182,N_26528,N_29598);
and U38183 (N_38183,N_27297,N_20039);
and U38184 (N_38184,N_20118,N_27121);
xor U38185 (N_38185,N_28909,N_26124);
nand U38186 (N_38186,N_22096,N_26431);
xnor U38187 (N_38187,N_26522,N_28060);
nor U38188 (N_38188,N_29178,N_24504);
nand U38189 (N_38189,N_27507,N_20240);
and U38190 (N_38190,N_29177,N_27945);
nand U38191 (N_38191,N_26461,N_26500);
nor U38192 (N_38192,N_21677,N_26307);
nand U38193 (N_38193,N_26337,N_22694);
and U38194 (N_38194,N_26516,N_23183);
nor U38195 (N_38195,N_21399,N_24664);
nor U38196 (N_38196,N_22672,N_27894);
or U38197 (N_38197,N_23544,N_26042);
and U38198 (N_38198,N_28786,N_26597);
nor U38199 (N_38199,N_24371,N_26612);
nor U38200 (N_38200,N_23955,N_27785);
nand U38201 (N_38201,N_22928,N_21009);
or U38202 (N_38202,N_27482,N_29859);
and U38203 (N_38203,N_23769,N_26829);
nor U38204 (N_38204,N_21129,N_27101);
or U38205 (N_38205,N_28115,N_27401);
nand U38206 (N_38206,N_24581,N_20687);
or U38207 (N_38207,N_23005,N_28642);
nor U38208 (N_38208,N_20651,N_28237);
nand U38209 (N_38209,N_26128,N_26681);
nor U38210 (N_38210,N_21877,N_29298);
nor U38211 (N_38211,N_29536,N_20938);
or U38212 (N_38212,N_28759,N_20500);
nor U38213 (N_38213,N_26070,N_22373);
nor U38214 (N_38214,N_29247,N_20239);
nand U38215 (N_38215,N_26931,N_24511);
or U38216 (N_38216,N_27437,N_28529);
nor U38217 (N_38217,N_27717,N_22500);
nand U38218 (N_38218,N_24669,N_25519);
and U38219 (N_38219,N_21413,N_29345);
or U38220 (N_38220,N_23140,N_26569);
or U38221 (N_38221,N_22642,N_27542);
xor U38222 (N_38222,N_25936,N_22356);
nand U38223 (N_38223,N_28365,N_29482);
nor U38224 (N_38224,N_26635,N_24295);
xnor U38225 (N_38225,N_28713,N_21469);
nand U38226 (N_38226,N_21651,N_26736);
or U38227 (N_38227,N_29442,N_23977);
xnor U38228 (N_38228,N_28770,N_25443);
nor U38229 (N_38229,N_29093,N_24371);
nand U38230 (N_38230,N_23844,N_27417);
or U38231 (N_38231,N_24607,N_22013);
and U38232 (N_38232,N_26401,N_23554);
nand U38233 (N_38233,N_21162,N_27856);
xnor U38234 (N_38234,N_20691,N_27196);
and U38235 (N_38235,N_20494,N_20003);
or U38236 (N_38236,N_28032,N_20461);
or U38237 (N_38237,N_21372,N_22177);
and U38238 (N_38238,N_26662,N_23532);
and U38239 (N_38239,N_27100,N_24623);
and U38240 (N_38240,N_23983,N_24053);
nand U38241 (N_38241,N_21486,N_23943);
nor U38242 (N_38242,N_24686,N_20699);
and U38243 (N_38243,N_23787,N_25757);
and U38244 (N_38244,N_25262,N_28827);
xnor U38245 (N_38245,N_21826,N_26158);
nor U38246 (N_38246,N_24883,N_26714);
nor U38247 (N_38247,N_24546,N_27063);
xor U38248 (N_38248,N_24274,N_24551);
and U38249 (N_38249,N_27211,N_24921);
nand U38250 (N_38250,N_22997,N_21864);
nand U38251 (N_38251,N_25946,N_28587);
and U38252 (N_38252,N_23078,N_26710);
or U38253 (N_38253,N_26942,N_24173);
nand U38254 (N_38254,N_25992,N_20400);
or U38255 (N_38255,N_23704,N_22832);
nor U38256 (N_38256,N_28649,N_29315);
or U38257 (N_38257,N_27950,N_29722);
or U38258 (N_38258,N_24551,N_29446);
xnor U38259 (N_38259,N_25635,N_29261);
or U38260 (N_38260,N_25488,N_27874);
or U38261 (N_38261,N_25818,N_27200);
nand U38262 (N_38262,N_22294,N_22873);
and U38263 (N_38263,N_26218,N_28100);
or U38264 (N_38264,N_25555,N_29411);
or U38265 (N_38265,N_25123,N_24164);
and U38266 (N_38266,N_25272,N_24929);
and U38267 (N_38267,N_21564,N_28606);
and U38268 (N_38268,N_25597,N_24112);
nand U38269 (N_38269,N_28354,N_25367);
nor U38270 (N_38270,N_25127,N_28554);
nor U38271 (N_38271,N_26435,N_24113);
and U38272 (N_38272,N_26037,N_20261);
or U38273 (N_38273,N_25468,N_26030);
or U38274 (N_38274,N_22466,N_21415);
nor U38275 (N_38275,N_20888,N_22656);
nor U38276 (N_38276,N_21769,N_29319);
nand U38277 (N_38277,N_22082,N_27847);
or U38278 (N_38278,N_20385,N_21438);
and U38279 (N_38279,N_24784,N_22862);
nand U38280 (N_38280,N_29588,N_28138);
nand U38281 (N_38281,N_28804,N_29466);
nor U38282 (N_38282,N_23040,N_26678);
and U38283 (N_38283,N_27460,N_23000);
nand U38284 (N_38284,N_22194,N_20313);
or U38285 (N_38285,N_21213,N_28695);
and U38286 (N_38286,N_24429,N_24539);
nor U38287 (N_38287,N_22620,N_27440);
xnor U38288 (N_38288,N_21811,N_21579);
and U38289 (N_38289,N_24492,N_26084);
xnor U38290 (N_38290,N_21507,N_24374);
nand U38291 (N_38291,N_24597,N_22370);
nand U38292 (N_38292,N_23444,N_22044);
and U38293 (N_38293,N_23512,N_21803);
and U38294 (N_38294,N_23718,N_21489);
or U38295 (N_38295,N_29841,N_29010);
or U38296 (N_38296,N_27468,N_29842);
or U38297 (N_38297,N_28362,N_20548);
or U38298 (N_38298,N_26975,N_20143);
nand U38299 (N_38299,N_21717,N_27803);
nor U38300 (N_38300,N_29602,N_27704);
and U38301 (N_38301,N_23144,N_21049);
and U38302 (N_38302,N_22885,N_29921);
xor U38303 (N_38303,N_28699,N_20157);
nand U38304 (N_38304,N_29937,N_29162);
and U38305 (N_38305,N_21851,N_21049);
nand U38306 (N_38306,N_29605,N_21193);
nand U38307 (N_38307,N_29826,N_22990);
xor U38308 (N_38308,N_26646,N_26693);
nand U38309 (N_38309,N_27761,N_26819);
and U38310 (N_38310,N_29253,N_24266);
or U38311 (N_38311,N_27390,N_26742);
nand U38312 (N_38312,N_26559,N_29931);
and U38313 (N_38313,N_21881,N_21759);
nor U38314 (N_38314,N_23911,N_20455);
and U38315 (N_38315,N_22949,N_23425);
nand U38316 (N_38316,N_26744,N_22896);
and U38317 (N_38317,N_23646,N_26986);
or U38318 (N_38318,N_23115,N_25906);
nor U38319 (N_38319,N_22256,N_29600);
and U38320 (N_38320,N_23263,N_23051);
or U38321 (N_38321,N_28517,N_25403);
nand U38322 (N_38322,N_24567,N_22431);
xnor U38323 (N_38323,N_26697,N_28379);
nor U38324 (N_38324,N_21036,N_24801);
nand U38325 (N_38325,N_21934,N_28170);
nand U38326 (N_38326,N_24819,N_29718);
nor U38327 (N_38327,N_29376,N_22918);
and U38328 (N_38328,N_27622,N_29154);
xnor U38329 (N_38329,N_23860,N_20641);
nor U38330 (N_38330,N_28627,N_26499);
nand U38331 (N_38331,N_28641,N_25024);
and U38332 (N_38332,N_24071,N_21662);
and U38333 (N_38333,N_21512,N_22796);
and U38334 (N_38334,N_28305,N_23226);
xor U38335 (N_38335,N_24891,N_24776);
nor U38336 (N_38336,N_23071,N_28794);
nor U38337 (N_38337,N_24831,N_29480);
and U38338 (N_38338,N_23017,N_20650);
and U38339 (N_38339,N_28635,N_29378);
or U38340 (N_38340,N_21524,N_20992);
or U38341 (N_38341,N_24976,N_20409);
or U38342 (N_38342,N_29088,N_28419);
nor U38343 (N_38343,N_29987,N_24540);
nor U38344 (N_38344,N_28668,N_24999);
nor U38345 (N_38345,N_27330,N_23590);
or U38346 (N_38346,N_21450,N_28035);
nand U38347 (N_38347,N_23876,N_24896);
nand U38348 (N_38348,N_22025,N_28696);
or U38349 (N_38349,N_23511,N_22692);
nor U38350 (N_38350,N_24417,N_27599);
nand U38351 (N_38351,N_24179,N_22182);
nor U38352 (N_38352,N_28403,N_20195);
and U38353 (N_38353,N_28596,N_21848);
and U38354 (N_38354,N_20449,N_24944);
nand U38355 (N_38355,N_20269,N_21282);
or U38356 (N_38356,N_26009,N_29629);
nand U38357 (N_38357,N_23942,N_29961);
and U38358 (N_38358,N_29472,N_23143);
and U38359 (N_38359,N_22667,N_28207);
and U38360 (N_38360,N_28247,N_23403);
nor U38361 (N_38361,N_26450,N_28118);
nand U38362 (N_38362,N_27779,N_29911);
or U38363 (N_38363,N_21821,N_29164);
and U38364 (N_38364,N_25836,N_22726);
nand U38365 (N_38365,N_20569,N_20132);
nand U38366 (N_38366,N_21930,N_21314);
nor U38367 (N_38367,N_28742,N_22849);
xor U38368 (N_38368,N_23197,N_26289);
or U38369 (N_38369,N_29410,N_23775);
nor U38370 (N_38370,N_29060,N_26962);
and U38371 (N_38371,N_21929,N_29726);
nand U38372 (N_38372,N_26141,N_28226);
xnor U38373 (N_38373,N_23321,N_26599);
xnor U38374 (N_38374,N_22661,N_21901);
nor U38375 (N_38375,N_21847,N_21134);
nor U38376 (N_38376,N_20126,N_29570);
or U38377 (N_38377,N_27692,N_24925);
or U38378 (N_38378,N_20763,N_26628);
and U38379 (N_38379,N_29054,N_22481);
nor U38380 (N_38380,N_27880,N_21909);
or U38381 (N_38381,N_28051,N_26428);
nand U38382 (N_38382,N_26758,N_23614);
nand U38383 (N_38383,N_27328,N_27326);
or U38384 (N_38384,N_23327,N_24318);
or U38385 (N_38385,N_23145,N_28539);
nor U38386 (N_38386,N_27335,N_28038);
or U38387 (N_38387,N_21438,N_22248);
or U38388 (N_38388,N_27286,N_21466);
nand U38389 (N_38389,N_22488,N_21555);
or U38390 (N_38390,N_25152,N_24290);
nor U38391 (N_38391,N_28783,N_21549);
nor U38392 (N_38392,N_27767,N_27092);
or U38393 (N_38393,N_24867,N_24428);
nand U38394 (N_38394,N_24158,N_27549);
or U38395 (N_38395,N_20214,N_22077);
nor U38396 (N_38396,N_27170,N_27617);
or U38397 (N_38397,N_22634,N_24749);
or U38398 (N_38398,N_25452,N_26499);
or U38399 (N_38399,N_27539,N_22164);
nand U38400 (N_38400,N_24842,N_28343);
xnor U38401 (N_38401,N_25401,N_27019);
xnor U38402 (N_38402,N_29228,N_23519);
nand U38403 (N_38403,N_24265,N_24259);
nor U38404 (N_38404,N_20789,N_20139);
nor U38405 (N_38405,N_29347,N_24722);
nor U38406 (N_38406,N_24633,N_21769);
or U38407 (N_38407,N_22045,N_26350);
nor U38408 (N_38408,N_25776,N_20395);
and U38409 (N_38409,N_25773,N_29538);
or U38410 (N_38410,N_27103,N_29286);
nor U38411 (N_38411,N_26199,N_27186);
xnor U38412 (N_38412,N_24209,N_25688);
or U38413 (N_38413,N_20531,N_21614);
or U38414 (N_38414,N_20763,N_27806);
nand U38415 (N_38415,N_26623,N_24658);
or U38416 (N_38416,N_22814,N_26949);
xnor U38417 (N_38417,N_29007,N_25870);
nor U38418 (N_38418,N_26201,N_23272);
nand U38419 (N_38419,N_21062,N_29414);
or U38420 (N_38420,N_27051,N_24431);
and U38421 (N_38421,N_26799,N_28547);
nor U38422 (N_38422,N_21090,N_21963);
nand U38423 (N_38423,N_28378,N_28293);
nand U38424 (N_38424,N_24090,N_27875);
nand U38425 (N_38425,N_22741,N_28756);
nor U38426 (N_38426,N_22621,N_29030);
nand U38427 (N_38427,N_29030,N_25419);
or U38428 (N_38428,N_25295,N_21735);
or U38429 (N_38429,N_26596,N_23071);
nor U38430 (N_38430,N_25358,N_20209);
xnor U38431 (N_38431,N_27638,N_26968);
or U38432 (N_38432,N_23921,N_27024);
or U38433 (N_38433,N_27265,N_27015);
nand U38434 (N_38434,N_23462,N_28559);
or U38435 (N_38435,N_27630,N_22326);
or U38436 (N_38436,N_29469,N_27122);
nand U38437 (N_38437,N_24412,N_28091);
or U38438 (N_38438,N_27028,N_24893);
nor U38439 (N_38439,N_22031,N_28280);
nor U38440 (N_38440,N_25758,N_28739);
nor U38441 (N_38441,N_28017,N_28052);
nor U38442 (N_38442,N_23525,N_20350);
nand U38443 (N_38443,N_23184,N_27498);
and U38444 (N_38444,N_29305,N_21078);
or U38445 (N_38445,N_29960,N_21095);
and U38446 (N_38446,N_29058,N_21699);
and U38447 (N_38447,N_29044,N_27137);
nand U38448 (N_38448,N_29939,N_21366);
nor U38449 (N_38449,N_23828,N_27725);
nand U38450 (N_38450,N_24608,N_23118);
nor U38451 (N_38451,N_23502,N_27463);
nand U38452 (N_38452,N_27792,N_23179);
or U38453 (N_38453,N_27589,N_21224);
or U38454 (N_38454,N_22497,N_29432);
or U38455 (N_38455,N_26457,N_25573);
nand U38456 (N_38456,N_23799,N_26418);
and U38457 (N_38457,N_20670,N_24617);
nor U38458 (N_38458,N_23884,N_20638);
nand U38459 (N_38459,N_25195,N_22930);
and U38460 (N_38460,N_24006,N_20166);
xor U38461 (N_38461,N_28659,N_20675);
nor U38462 (N_38462,N_27590,N_24214);
xor U38463 (N_38463,N_20339,N_21285);
xor U38464 (N_38464,N_25132,N_22833);
and U38465 (N_38465,N_20990,N_25280);
nand U38466 (N_38466,N_21436,N_24034);
nand U38467 (N_38467,N_20436,N_26958);
and U38468 (N_38468,N_23492,N_20676);
nand U38469 (N_38469,N_28881,N_28801);
nand U38470 (N_38470,N_28113,N_22342);
nor U38471 (N_38471,N_25088,N_28688);
nand U38472 (N_38472,N_29028,N_22005);
xnor U38473 (N_38473,N_26496,N_22903);
nand U38474 (N_38474,N_29477,N_21171);
or U38475 (N_38475,N_24005,N_20976);
nor U38476 (N_38476,N_21063,N_27506);
nor U38477 (N_38477,N_22424,N_20114);
nor U38478 (N_38478,N_26912,N_29310);
nor U38479 (N_38479,N_27341,N_27137);
and U38480 (N_38480,N_21699,N_27169);
nor U38481 (N_38481,N_26752,N_26961);
xor U38482 (N_38482,N_29246,N_29391);
nor U38483 (N_38483,N_21101,N_21582);
and U38484 (N_38484,N_22320,N_26181);
xor U38485 (N_38485,N_20409,N_29677);
or U38486 (N_38486,N_25397,N_22106);
or U38487 (N_38487,N_22013,N_24070);
and U38488 (N_38488,N_22135,N_28366);
and U38489 (N_38489,N_25617,N_24761);
and U38490 (N_38490,N_27180,N_22689);
nand U38491 (N_38491,N_20935,N_26949);
nor U38492 (N_38492,N_29530,N_21998);
or U38493 (N_38493,N_23041,N_28821);
and U38494 (N_38494,N_23072,N_27914);
nand U38495 (N_38495,N_28706,N_23068);
xor U38496 (N_38496,N_21451,N_23289);
and U38497 (N_38497,N_25899,N_22890);
xor U38498 (N_38498,N_22659,N_21188);
and U38499 (N_38499,N_28578,N_20370);
nand U38500 (N_38500,N_20005,N_24617);
or U38501 (N_38501,N_28930,N_22908);
nand U38502 (N_38502,N_21112,N_22340);
xnor U38503 (N_38503,N_25795,N_22576);
and U38504 (N_38504,N_21601,N_26416);
or U38505 (N_38505,N_27869,N_29135);
or U38506 (N_38506,N_29529,N_25663);
or U38507 (N_38507,N_22238,N_26388);
nand U38508 (N_38508,N_21615,N_26546);
nor U38509 (N_38509,N_28112,N_28366);
and U38510 (N_38510,N_24253,N_21875);
or U38511 (N_38511,N_20537,N_21187);
nand U38512 (N_38512,N_23654,N_21893);
and U38513 (N_38513,N_25308,N_28347);
and U38514 (N_38514,N_20127,N_24034);
nand U38515 (N_38515,N_20743,N_26765);
and U38516 (N_38516,N_26267,N_22200);
nand U38517 (N_38517,N_27662,N_25544);
nand U38518 (N_38518,N_20845,N_29510);
nor U38519 (N_38519,N_25868,N_25539);
and U38520 (N_38520,N_26592,N_26478);
xnor U38521 (N_38521,N_29237,N_25617);
nand U38522 (N_38522,N_24524,N_24761);
nand U38523 (N_38523,N_28748,N_24368);
nor U38524 (N_38524,N_25326,N_27371);
or U38525 (N_38525,N_29571,N_28174);
or U38526 (N_38526,N_20573,N_29248);
xnor U38527 (N_38527,N_29977,N_28241);
nor U38528 (N_38528,N_25882,N_25085);
or U38529 (N_38529,N_23647,N_23394);
nor U38530 (N_38530,N_20162,N_26750);
and U38531 (N_38531,N_27069,N_29758);
and U38532 (N_38532,N_28138,N_21940);
or U38533 (N_38533,N_22012,N_21901);
or U38534 (N_38534,N_21748,N_24370);
xor U38535 (N_38535,N_26518,N_25280);
and U38536 (N_38536,N_25170,N_27251);
or U38537 (N_38537,N_20193,N_20891);
or U38538 (N_38538,N_26562,N_25054);
nand U38539 (N_38539,N_24525,N_28070);
nand U38540 (N_38540,N_28993,N_20328);
nand U38541 (N_38541,N_27049,N_21745);
nor U38542 (N_38542,N_28213,N_25533);
nand U38543 (N_38543,N_21978,N_29474);
xnor U38544 (N_38544,N_25228,N_26156);
or U38545 (N_38545,N_23578,N_20884);
nor U38546 (N_38546,N_21034,N_26361);
or U38547 (N_38547,N_25666,N_22104);
nor U38548 (N_38548,N_23486,N_29232);
and U38549 (N_38549,N_26328,N_27082);
and U38550 (N_38550,N_27310,N_24959);
and U38551 (N_38551,N_21571,N_27979);
or U38552 (N_38552,N_29590,N_22906);
nand U38553 (N_38553,N_28223,N_23672);
nor U38554 (N_38554,N_21474,N_20458);
or U38555 (N_38555,N_23466,N_23111);
xnor U38556 (N_38556,N_21093,N_23546);
or U38557 (N_38557,N_29445,N_22751);
nand U38558 (N_38558,N_21911,N_23106);
nand U38559 (N_38559,N_27928,N_29961);
nor U38560 (N_38560,N_21603,N_23386);
nor U38561 (N_38561,N_29842,N_29887);
nand U38562 (N_38562,N_20289,N_20210);
and U38563 (N_38563,N_23917,N_23482);
and U38564 (N_38564,N_27292,N_21364);
and U38565 (N_38565,N_25634,N_20318);
and U38566 (N_38566,N_28109,N_22018);
or U38567 (N_38567,N_23685,N_20868);
and U38568 (N_38568,N_22913,N_22713);
nand U38569 (N_38569,N_27007,N_25677);
nand U38570 (N_38570,N_29065,N_25714);
xor U38571 (N_38571,N_26131,N_24367);
and U38572 (N_38572,N_28992,N_28535);
and U38573 (N_38573,N_21121,N_27361);
or U38574 (N_38574,N_26406,N_23323);
nand U38575 (N_38575,N_22357,N_20290);
nand U38576 (N_38576,N_25294,N_21120);
or U38577 (N_38577,N_25386,N_21044);
or U38578 (N_38578,N_23229,N_26725);
nor U38579 (N_38579,N_24633,N_28519);
xnor U38580 (N_38580,N_24564,N_21197);
nor U38581 (N_38581,N_24385,N_20092);
and U38582 (N_38582,N_23386,N_22648);
nand U38583 (N_38583,N_21653,N_21112);
and U38584 (N_38584,N_22846,N_27135);
nor U38585 (N_38585,N_28881,N_22197);
or U38586 (N_38586,N_28253,N_22093);
nor U38587 (N_38587,N_20117,N_24590);
and U38588 (N_38588,N_24180,N_29766);
nand U38589 (N_38589,N_23527,N_20496);
or U38590 (N_38590,N_26841,N_26229);
nand U38591 (N_38591,N_29753,N_28310);
and U38592 (N_38592,N_24453,N_29966);
and U38593 (N_38593,N_23345,N_21373);
nand U38594 (N_38594,N_28167,N_20402);
and U38595 (N_38595,N_20362,N_27265);
nand U38596 (N_38596,N_24856,N_20659);
nor U38597 (N_38597,N_28929,N_22564);
and U38598 (N_38598,N_22666,N_22455);
and U38599 (N_38599,N_25621,N_28776);
or U38600 (N_38600,N_23862,N_27547);
or U38601 (N_38601,N_22499,N_26704);
nor U38602 (N_38602,N_21728,N_21558);
xor U38603 (N_38603,N_29614,N_29997);
nand U38604 (N_38604,N_26910,N_23275);
or U38605 (N_38605,N_23127,N_23043);
nand U38606 (N_38606,N_27752,N_20231);
nand U38607 (N_38607,N_22995,N_29189);
nor U38608 (N_38608,N_22227,N_29752);
nand U38609 (N_38609,N_20291,N_29762);
or U38610 (N_38610,N_24209,N_29317);
xnor U38611 (N_38611,N_20582,N_27449);
or U38612 (N_38612,N_26187,N_23316);
or U38613 (N_38613,N_28839,N_25246);
and U38614 (N_38614,N_24754,N_25805);
nor U38615 (N_38615,N_20171,N_28052);
nand U38616 (N_38616,N_22789,N_22037);
nor U38617 (N_38617,N_28870,N_25924);
and U38618 (N_38618,N_20036,N_25721);
nor U38619 (N_38619,N_21159,N_28514);
or U38620 (N_38620,N_25308,N_20992);
and U38621 (N_38621,N_22267,N_26540);
and U38622 (N_38622,N_25141,N_25186);
nor U38623 (N_38623,N_28717,N_21354);
or U38624 (N_38624,N_29040,N_24213);
nand U38625 (N_38625,N_20379,N_21846);
or U38626 (N_38626,N_25799,N_24640);
nand U38627 (N_38627,N_26522,N_20587);
nand U38628 (N_38628,N_27846,N_24250);
and U38629 (N_38629,N_26987,N_25081);
or U38630 (N_38630,N_29316,N_25949);
or U38631 (N_38631,N_22877,N_21543);
nor U38632 (N_38632,N_27577,N_20056);
xnor U38633 (N_38633,N_23388,N_26325);
and U38634 (N_38634,N_22298,N_28556);
and U38635 (N_38635,N_28321,N_25819);
and U38636 (N_38636,N_25865,N_29022);
or U38637 (N_38637,N_29934,N_23000);
or U38638 (N_38638,N_25257,N_25839);
nand U38639 (N_38639,N_21594,N_28821);
or U38640 (N_38640,N_25220,N_22938);
nand U38641 (N_38641,N_25150,N_27861);
nor U38642 (N_38642,N_26223,N_25723);
nand U38643 (N_38643,N_26289,N_26738);
nor U38644 (N_38644,N_20194,N_25231);
nor U38645 (N_38645,N_28468,N_21598);
nor U38646 (N_38646,N_20641,N_29194);
or U38647 (N_38647,N_22349,N_26546);
and U38648 (N_38648,N_28337,N_24290);
or U38649 (N_38649,N_21352,N_22024);
nand U38650 (N_38650,N_20921,N_23249);
xor U38651 (N_38651,N_26964,N_20806);
nor U38652 (N_38652,N_24492,N_24725);
and U38653 (N_38653,N_25521,N_29014);
nand U38654 (N_38654,N_27127,N_23244);
nor U38655 (N_38655,N_24870,N_25718);
nor U38656 (N_38656,N_24334,N_28097);
or U38657 (N_38657,N_23485,N_24315);
nor U38658 (N_38658,N_26402,N_24582);
nand U38659 (N_38659,N_27344,N_26095);
or U38660 (N_38660,N_26242,N_22944);
nor U38661 (N_38661,N_26942,N_22963);
nand U38662 (N_38662,N_20141,N_24051);
nand U38663 (N_38663,N_25914,N_29621);
or U38664 (N_38664,N_24236,N_24386);
and U38665 (N_38665,N_22942,N_25500);
and U38666 (N_38666,N_29020,N_21869);
and U38667 (N_38667,N_24748,N_20075);
or U38668 (N_38668,N_20848,N_23991);
nand U38669 (N_38669,N_26043,N_21875);
nor U38670 (N_38670,N_28722,N_28723);
nand U38671 (N_38671,N_21428,N_20597);
and U38672 (N_38672,N_23522,N_28467);
or U38673 (N_38673,N_25105,N_24703);
nor U38674 (N_38674,N_22510,N_29437);
or U38675 (N_38675,N_22975,N_21412);
and U38676 (N_38676,N_24528,N_21005);
and U38677 (N_38677,N_27404,N_27385);
nor U38678 (N_38678,N_25361,N_22630);
nor U38679 (N_38679,N_22891,N_24594);
and U38680 (N_38680,N_20253,N_23763);
xor U38681 (N_38681,N_26098,N_27049);
and U38682 (N_38682,N_28970,N_22616);
nand U38683 (N_38683,N_21107,N_23651);
nand U38684 (N_38684,N_24420,N_24174);
nor U38685 (N_38685,N_28136,N_24194);
nor U38686 (N_38686,N_26062,N_29632);
nor U38687 (N_38687,N_26206,N_26885);
or U38688 (N_38688,N_20942,N_23384);
and U38689 (N_38689,N_20970,N_26964);
nand U38690 (N_38690,N_23097,N_24213);
or U38691 (N_38691,N_27524,N_23118);
or U38692 (N_38692,N_23936,N_20897);
and U38693 (N_38693,N_21527,N_24057);
and U38694 (N_38694,N_29356,N_23822);
and U38695 (N_38695,N_29066,N_28063);
nand U38696 (N_38696,N_25632,N_29198);
nor U38697 (N_38697,N_24660,N_22901);
nand U38698 (N_38698,N_27135,N_20321);
and U38699 (N_38699,N_25594,N_29403);
nor U38700 (N_38700,N_27318,N_26074);
and U38701 (N_38701,N_21567,N_22787);
and U38702 (N_38702,N_20324,N_27845);
or U38703 (N_38703,N_20420,N_24131);
or U38704 (N_38704,N_26840,N_24273);
and U38705 (N_38705,N_27237,N_21657);
nand U38706 (N_38706,N_20558,N_27139);
nand U38707 (N_38707,N_24598,N_28748);
nor U38708 (N_38708,N_21439,N_21400);
or U38709 (N_38709,N_25215,N_22352);
or U38710 (N_38710,N_22039,N_26182);
nor U38711 (N_38711,N_20243,N_23386);
nand U38712 (N_38712,N_25290,N_25948);
or U38713 (N_38713,N_24113,N_22239);
and U38714 (N_38714,N_25566,N_20844);
xor U38715 (N_38715,N_25796,N_27099);
or U38716 (N_38716,N_24444,N_24540);
nand U38717 (N_38717,N_21576,N_23717);
and U38718 (N_38718,N_26742,N_28190);
nor U38719 (N_38719,N_21533,N_22481);
or U38720 (N_38720,N_20730,N_21490);
and U38721 (N_38721,N_25592,N_24306);
nand U38722 (N_38722,N_21465,N_23111);
or U38723 (N_38723,N_28253,N_26804);
xor U38724 (N_38724,N_27781,N_24897);
nand U38725 (N_38725,N_28982,N_25597);
nand U38726 (N_38726,N_28035,N_23463);
nor U38727 (N_38727,N_23154,N_21348);
nor U38728 (N_38728,N_21238,N_25987);
nand U38729 (N_38729,N_24656,N_26180);
or U38730 (N_38730,N_25530,N_25509);
xor U38731 (N_38731,N_25295,N_21783);
or U38732 (N_38732,N_29343,N_23526);
nand U38733 (N_38733,N_26901,N_25874);
nor U38734 (N_38734,N_28810,N_20347);
and U38735 (N_38735,N_24554,N_24302);
nand U38736 (N_38736,N_27769,N_28403);
or U38737 (N_38737,N_29781,N_28407);
nor U38738 (N_38738,N_20673,N_26922);
nor U38739 (N_38739,N_23121,N_27457);
nor U38740 (N_38740,N_28244,N_29979);
nand U38741 (N_38741,N_25106,N_23902);
and U38742 (N_38742,N_27410,N_29387);
nand U38743 (N_38743,N_29374,N_20334);
and U38744 (N_38744,N_25845,N_21574);
and U38745 (N_38745,N_27014,N_20648);
or U38746 (N_38746,N_21236,N_24474);
or U38747 (N_38747,N_26632,N_20271);
and U38748 (N_38748,N_27458,N_22509);
or U38749 (N_38749,N_26931,N_25759);
or U38750 (N_38750,N_25161,N_21651);
xnor U38751 (N_38751,N_27990,N_20224);
nand U38752 (N_38752,N_25648,N_20344);
xnor U38753 (N_38753,N_29947,N_21885);
nor U38754 (N_38754,N_23891,N_21152);
and U38755 (N_38755,N_23350,N_28698);
nand U38756 (N_38756,N_26557,N_28643);
and U38757 (N_38757,N_20342,N_22036);
nor U38758 (N_38758,N_28535,N_22710);
nor U38759 (N_38759,N_20649,N_24622);
or U38760 (N_38760,N_22211,N_23079);
nand U38761 (N_38761,N_25556,N_27784);
nor U38762 (N_38762,N_23444,N_26779);
and U38763 (N_38763,N_24949,N_24445);
nor U38764 (N_38764,N_28483,N_20929);
nand U38765 (N_38765,N_27741,N_23215);
or U38766 (N_38766,N_28639,N_26483);
xnor U38767 (N_38767,N_23380,N_24267);
xnor U38768 (N_38768,N_29588,N_29160);
nor U38769 (N_38769,N_27487,N_24199);
nand U38770 (N_38770,N_22202,N_27894);
nand U38771 (N_38771,N_29071,N_20400);
or U38772 (N_38772,N_24756,N_27320);
nand U38773 (N_38773,N_20122,N_21976);
or U38774 (N_38774,N_24255,N_26552);
nor U38775 (N_38775,N_26603,N_24266);
nand U38776 (N_38776,N_23121,N_25551);
and U38777 (N_38777,N_23502,N_29267);
nor U38778 (N_38778,N_21865,N_24473);
and U38779 (N_38779,N_25484,N_25330);
and U38780 (N_38780,N_23743,N_27722);
nor U38781 (N_38781,N_27133,N_26536);
nor U38782 (N_38782,N_22373,N_27500);
or U38783 (N_38783,N_22426,N_29511);
and U38784 (N_38784,N_20396,N_25802);
xor U38785 (N_38785,N_25764,N_22032);
nor U38786 (N_38786,N_20332,N_25922);
nor U38787 (N_38787,N_24255,N_24784);
nand U38788 (N_38788,N_27132,N_24858);
or U38789 (N_38789,N_29684,N_26463);
and U38790 (N_38790,N_23899,N_21299);
xor U38791 (N_38791,N_28977,N_23592);
xnor U38792 (N_38792,N_21314,N_25012);
nor U38793 (N_38793,N_28726,N_25138);
nand U38794 (N_38794,N_20113,N_28331);
nand U38795 (N_38795,N_27613,N_27707);
and U38796 (N_38796,N_29229,N_28316);
or U38797 (N_38797,N_24092,N_23365);
and U38798 (N_38798,N_26927,N_26221);
nand U38799 (N_38799,N_20924,N_26626);
nand U38800 (N_38800,N_27932,N_25849);
nand U38801 (N_38801,N_29313,N_26612);
nor U38802 (N_38802,N_29925,N_27632);
and U38803 (N_38803,N_24371,N_20293);
and U38804 (N_38804,N_28245,N_21183);
nor U38805 (N_38805,N_24908,N_23592);
or U38806 (N_38806,N_20028,N_23156);
or U38807 (N_38807,N_22289,N_29949);
and U38808 (N_38808,N_22532,N_26175);
and U38809 (N_38809,N_21981,N_22629);
nor U38810 (N_38810,N_25590,N_27463);
nand U38811 (N_38811,N_28127,N_22672);
xnor U38812 (N_38812,N_20893,N_23264);
and U38813 (N_38813,N_23570,N_21140);
nor U38814 (N_38814,N_23450,N_29990);
and U38815 (N_38815,N_22985,N_23171);
nand U38816 (N_38816,N_23576,N_23230);
or U38817 (N_38817,N_23200,N_21644);
nor U38818 (N_38818,N_25938,N_27641);
xnor U38819 (N_38819,N_28005,N_22917);
or U38820 (N_38820,N_26424,N_28211);
nand U38821 (N_38821,N_29311,N_26785);
or U38822 (N_38822,N_25777,N_25249);
xor U38823 (N_38823,N_20330,N_26006);
nor U38824 (N_38824,N_25945,N_21521);
or U38825 (N_38825,N_26792,N_27174);
nand U38826 (N_38826,N_24315,N_23245);
nor U38827 (N_38827,N_24121,N_21948);
xnor U38828 (N_38828,N_26559,N_23291);
nor U38829 (N_38829,N_26942,N_28858);
and U38830 (N_38830,N_24348,N_20825);
nand U38831 (N_38831,N_27383,N_24427);
and U38832 (N_38832,N_29244,N_25300);
xnor U38833 (N_38833,N_27291,N_26590);
and U38834 (N_38834,N_27253,N_20663);
nand U38835 (N_38835,N_24612,N_22297);
nor U38836 (N_38836,N_27435,N_28880);
xnor U38837 (N_38837,N_22269,N_27491);
and U38838 (N_38838,N_21663,N_27375);
and U38839 (N_38839,N_23717,N_25629);
nor U38840 (N_38840,N_25572,N_28492);
and U38841 (N_38841,N_22549,N_20241);
nor U38842 (N_38842,N_27808,N_26397);
nand U38843 (N_38843,N_26511,N_28095);
and U38844 (N_38844,N_26581,N_20162);
nor U38845 (N_38845,N_27656,N_22595);
nor U38846 (N_38846,N_27140,N_27704);
nand U38847 (N_38847,N_20546,N_25624);
and U38848 (N_38848,N_24775,N_25712);
or U38849 (N_38849,N_20533,N_22538);
nor U38850 (N_38850,N_23300,N_27775);
nor U38851 (N_38851,N_20024,N_22744);
and U38852 (N_38852,N_24549,N_27928);
nand U38853 (N_38853,N_24523,N_26714);
nand U38854 (N_38854,N_29410,N_29575);
nor U38855 (N_38855,N_29741,N_27226);
and U38856 (N_38856,N_25160,N_29970);
xnor U38857 (N_38857,N_23116,N_29058);
or U38858 (N_38858,N_22708,N_27514);
or U38859 (N_38859,N_24487,N_23807);
and U38860 (N_38860,N_20726,N_23622);
and U38861 (N_38861,N_27817,N_21183);
xor U38862 (N_38862,N_21122,N_28124);
or U38863 (N_38863,N_20188,N_21115);
nand U38864 (N_38864,N_26274,N_29467);
or U38865 (N_38865,N_22543,N_22076);
or U38866 (N_38866,N_20545,N_26003);
nand U38867 (N_38867,N_21417,N_22599);
and U38868 (N_38868,N_23260,N_26623);
nand U38869 (N_38869,N_28575,N_24771);
nor U38870 (N_38870,N_26611,N_28412);
nor U38871 (N_38871,N_22998,N_24148);
nand U38872 (N_38872,N_20442,N_29366);
nor U38873 (N_38873,N_22036,N_20472);
nand U38874 (N_38874,N_26964,N_23179);
xnor U38875 (N_38875,N_20645,N_27944);
and U38876 (N_38876,N_28283,N_25708);
or U38877 (N_38877,N_24156,N_27974);
nand U38878 (N_38878,N_23500,N_23427);
and U38879 (N_38879,N_22063,N_23943);
nor U38880 (N_38880,N_22492,N_27266);
and U38881 (N_38881,N_25070,N_27521);
and U38882 (N_38882,N_26094,N_28220);
and U38883 (N_38883,N_23342,N_21150);
nand U38884 (N_38884,N_26775,N_25217);
nor U38885 (N_38885,N_22657,N_27666);
xor U38886 (N_38886,N_20272,N_23725);
nand U38887 (N_38887,N_20529,N_23572);
or U38888 (N_38888,N_21887,N_29708);
nor U38889 (N_38889,N_20326,N_28589);
and U38890 (N_38890,N_28968,N_20444);
nor U38891 (N_38891,N_26404,N_25094);
nand U38892 (N_38892,N_22190,N_24668);
nor U38893 (N_38893,N_25874,N_21145);
and U38894 (N_38894,N_22252,N_29645);
nor U38895 (N_38895,N_20824,N_25692);
and U38896 (N_38896,N_20397,N_21041);
nand U38897 (N_38897,N_26912,N_25814);
nand U38898 (N_38898,N_24510,N_21921);
nor U38899 (N_38899,N_23215,N_25713);
nand U38900 (N_38900,N_28762,N_21811);
or U38901 (N_38901,N_21591,N_26275);
nand U38902 (N_38902,N_27584,N_24525);
or U38903 (N_38903,N_21686,N_26156);
nor U38904 (N_38904,N_23264,N_24648);
or U38905 (N_38905,N_29559,N_25670);
and U38906 (N_38906,N_23268,N_24501);
nor U38907 (N_38907,N_26710,N_29854);
nor U38908 (N_38908,N_25955,N_27772);
nor U38909 (N_38909,N_20082,N_26326);
nor U38910 (N_38910,N_29496,N_20252);
and U38911 (N_38911,N_29448,N_21767);
and U38912 (N_38912,N_28851,N_28798);
or U38913 (N_38913,N_22982,N_27190);
nand U38914 (N_38914,N_28139,N_20368);
and U38915 (N_38915,N_24804,N_28236);
and U38916 (N_38916,N_24277,N_20795);
nor U38917 (N_38917,N_22155,N_22403);
nor U38918 (N_38918,N_23963,N_24264);
nand U38919 (N_38919,N_23129,N_20074);
nor U38920 (N_38920,N_23470,N_29882);
nand U38921 (N_38921,N_20209,N_26334);
xor U38922 (N_38922,N_26356,N_22315);
nand U38923 (N_38923,N_28563,N_24818);
and U38924 (N_38924,N_20269,N_29624);
or U38925 (N_38925,N_27866,N_23640);
nor U38926 (N_38926,N_28348,N_22924);
and U38927 (N_38927,N_29193,N_22602);
nor U38928 (N_38928,N_26864,N_25389);
nor U38929 (N_38929,N_25780,N_29077);
nand U38930 (N_38930,N_27126,N_24871);
nor U38931 (N_38931,N_23630,N_23396);
and U38932 (N_38932,N_28150,N_22208);
and U38933 (N_38933,N_26739,N_22651);
and U38934 (N_38934,N_27975,N_25685);
nand U38935 (N_38935,N_24525,N_23410);
or U38936 (N_38936,N_28803,N_29590);
nor U38937 (N_38937,N_25626,N_20575);
or U38938 (N_38938,N_26513,N_26318);
or U38939 (N_38939,N_20206,N_27589);
nor U38940 (N_38940,N_29558,N_25610);
xnor U38941 (N_38941,N_28203,N_24392);
and U38942 (N_38942,N_21824,N_21187);
nand U38943 (N_38943,N_21221,N_22515);
nand U38944 (N_38944,N_21471,N_27073);
or U38945 (N_38945,N_29600,N_22912);
nand U38946 (N_38946,N_23890,N_26577);
nand U38947 (N_38947,N_26475,N_20198);
xnor U38948 (N_38948,N_27031,N_29963);
nand U38949 (N_38949,N_22100,N_21823);
and U38950 (N_38950,N_24475,N_25352);
or U38951 (N_38951,N_29124,N_24265);
nand U38952 (N_38952,N_29272,N_24370);
and U38953 (N_38953,N_23126,N_24113);
xnor U38954 (N_38954,N_22862,N_22031);
and U38955 (N_38955,N_29501,N_29255);
nand U38956 (N_38956,N_24134,N_29820);
nor U38957 (N_38957,N_29613,N_29129);
or U38958 (N_38958,N_22107,N_23354);
nor U38959 (N_38959,N_29706,N_24503);
and U38960 (N_38960,N_28728,N_26080);
nand U38961 (N_38961,N_26241,N_23794);
and U38962 (N_38962,N_23147,N_21214);
nor U38963 (N_38963,N_23595,N_25143);
and U38964 (N_38964,N_25474,N_23318);
nor U38965 (N_38965,N_26903,N_24469);
nand U38966 (N_38966,N_22506,N_23128);
and U38967 (N_38967,N_26542,N_20848);
nand U38968 (N_38968,N_28946,N_29200);
and U38969 (N_38969,N_29860,N_23218);
or U38970 (N_38970,N_24447,N_27028);
and U38971 (N_38971,N_28680,N_29840);
nand U38972 (N_38972,N_27651,N_28052);
and U38973 (N_38973,N_27629,N_24510);
or U38974 (N_38974,N_23594,N_26657);
xnor U38975 (N_38975,N_29048,N_28540);
and U38976 (N_38976,N_21932,N_24140);
xnor U38977 (N_38977,N_21487,N_26096);
and U38978 (N_38978,N_26751,N_21771);
nand U38979 (N_38979,N_21174,N_27629);
nand U38980 (N_38980,N_27805,N_26958);
and U38981 (N_38981,N_21390,N_21836);
nor U38982 (N_38982,N_28516,N_25206);
or U38983 (N_38983,N_28753,N_25537);
or U38984 (N_38984,N_22646,N_20077);
nand U38985 (N_38985,N_20976,N_24286);
nor U38986 (N_38986,N_25565,N_29994);
xnor U38987 (N_38987,N_21221,N_27394);
and U38988 (N_38988,N_27328,N_25652);
or U38989 (N_38989,N_21549,N_21821);
nor U38990 (N_38990,N_26575,N_21051);
and U38991 (N_38991,N_27555,N_27848);
and U38992 (N_38992,N_25053,N_28300);
or U38993 (N_38993,N_29819,N_23689);
or U38994 (N_38994,N_29903,N_27362);
nor U38995 (N_38995,N_28065,N_23749);
and U38996 (N_38996,N_25734,N_21581);
and U38997 (N_38997,N_25129,N_23306);
or U38998 (N_38998,N_27954,N_26965);
xnor U38999 (N_38999,N_21567,N_23013);
nor U39000 (N_39000,N_24064,N_22054);
and U39001 (N_39001,N_20925,N_21312);
and U39002 (N_39002,N_28114,N_20452);
nor U39003 (N_39003,N_20183,N_20107);
and U39004 (N_39004,N_20961,N_23864);
or U39005 (N_39005,N_24711,N_25027);
nor U39006 (N_39006,N_26846,N_20778);
xor U39007 (N_39007,N_24950,N_26133);
xor U39008 (N_39008,N_24467,N_29798);
xnor U39009 (N_39009,N_21292,N_23761);
and U39010 (N_39010,N_23343,N_25578);
nand U39011 (N_39011,N_26019,N_25249);
and U39012 (N_39012,N_25732,N_20980);
nand U39013 (N_39013,N_23054,N_26144);
and U39014 (N_39014,N_22624,N_29664);
nor U39015 (N_39015,N_21232,N_25464);
nand U39016 (N_39016,N_22726,N_24832);
nand U39017 (N_39017,N_21635,N_26569);
or U39018 (N_39018,N_23588,N_21121);
nor U39019 (N_39019,N_26906,N_28153);
nor U39020 (N_39020,N_29934,N_20707);
and U39021 (N_39021,N_21943,N_24604);
xor U39022 (N_39022,N_21188,N_20504);
nand U39023 (N_39023,N_28589,N_21183);
and U39024 (N_39024,N_23802,N_28022);
or U39025 (N_39025,N_25022,N_26371);
and U39026 (N_39026,N_22467,N_23012);
nand U39027 (N_39027,N_29875,N_26132);
nor U39028 (N_39028,N_25672,N_29681);
or U39029 (N_39029,N_21021,N_22582);
and U39030 (N_39030,N_21370,N_29942);
and U39031 (N_39031,N_20551,N_20440);
nor U39032 (N_39032,N_29576,N_26278);
and U39033 (N_39033,N_29697,N_27165);
nor U39034 (N_39034,N_29875,N_28609);
and U39035 (N_39035,N_28874,N_28717);
or U39036 (N_39036,N_29605,N_21797);
xnor U39037 (N_39037,N_26314,N_22977);
nor U39038 (N_39038,N_20727,N_27593);
and U39039 (N_39039,N_27767,N_23008);
nor U39040 (N_39040,N_27728,N_25031);
nand U39041 (N_39041,N_28248,N_25330);
or U39042 (N_39042,N_26363,N_20435);
nand U39043 (N_39043,N_23834,N_22101);
nor U39044 (N_39044,N_22821,N_26596);
and U39045 (N_39045,N_21021,N_25957);
nand U39046 (N_39046,N_24569,N_29074);
and U39047 (N_39047,N_27125,N_26661);
and U39048 (N_39048,N_29065,N_27661);
xor U39049 (N_39049,N_24051,N_28310);
nor U39050 (N_39050,N_22457,N_20319);
xnor U39051 (N_39051,N_28826,N_21281);
nor U39052 (N_39052,N_22817,N_21214);
nand U39053 (N_39053,N_28338,N_24651);
or U39054 (N_39054,N_28933,N_23187);
or U39055 (N_39055,N_29738,N_20201);
and U39056 (N_39056,N_29678,N_24299);
nand U39057 (N_39057,N_20089,N_28109);
or U39058 (N_39058,N_24955,N_25214);
nor U39059 (N_39059,N_25709,N_26558);
nand U39060 (N_39060,N_29166,N_22490);
nor U39061 (N_39061,N_22485,N_23918);
nand U39062 (N_39062,N_29461,N_21911);
or U39063 (N_39063,N_24807,N_27265);
or U39064 (N_39064,N_22339,N_28506);
and U39065 (N_39065,N_28561,N_26172);
and U39066 (N_39066,N_24393,N_24014);
nand U39067 (N_39067,N_23448,N_20613);
and U39068 (N_39068,N_28382,N_28747);
and U39069 (N_39069,N_23585,N_20849);
nand U39070 (N_39070,N_20095,N_25090);
nand U39071 (N_39071,N_25976,N_24778);
nor U39072 (N_39072,N_27472,N_28190);
or U39073 (N_39073,N_25380,N_26044);
xor U39074 (N_39074,N_29177,N_29680);
or U39075 (N_39075,N_26123,N_21866);
nand U39076 (N_39076,N_29202,N_29937);
xor U39077 (N_39077,N_29005,N_28884);
and U39078 (N_39078,N_23451,N_25062);
nand U39079 (N_39079,N_28676,N_28657);
and U39080 (N_39080,N_23444,N_24503);
xor U39081 (N_39081,N_24792,N_20347);
or U39082 (N_39082,N_27979,N_23469);
nor U39083 (N_39083,N_25370,N_22639);
or U39084 (N_39084,N_24682,N_25127);
nand U39085 (N_39085,N_26122,N_20486);
nand U39086 (N_39086,N_26964,N_26092);
and U39087 (N_39087,N_22512,N_23930);
nor U39088 (N_39088,N_26746,N_25481);
or U39089 (N_39089,N_26868,N_23903);
and U39090 (N_39090,N_23239,N_21652);
xnor U39091 (N_39091,N_26205,N_20161);
or U39092 (N_39092,N_23665,N_23659);
nor U39093 (N_39093,N_27431,N_22892);
nor U39094 (N_39094,N_24590,N_20290);
nand U39095 (N_39095,N_25905,N_27747);
xnor U39096 (N_39096,N_20836,N_20628);
nand U39097 (N_39097,N_24715,N_28014);
nor U39098 (N_39098,N_23615,N_22840);
nand U39099 (N_39099,N_27746,N_26651);
and U39100 (N_39100,N_23894,N_21481);
nand U39101 (N_39101,N_21747,N_24560);
nor U39102 (N_39102,N_24164,N_25042);
nor U39103 (N_39103,N_23066,N_28056);
nor U39104 (N_39104,N_28649,N_24497);
or U39105 (N_39105,N_24249,N_23668);
xnor U39106 (N_39106,N_22807,N_29405);
xnor U39107 (N_39107,N_29663,N_28104);
nor U39108 (N_39108,N_29745,N_23899);
nor U39109 (N_39109,N_25754,N_29432);
and U39110 (N_39110,N_26096,N_29766);
nor U39111 (N_39111,N_26428,N_29088);
nor U39112 (N_39112,N_20729,N_23355);
nor U39113 (N_39113,N_22584,N_25029);
nor U39114 (N_39114,N_25323,N_25733);
or U39115 (N_39115,N_20643,N_29340);
nor U39116 (N_39116,N_29086,N_20172);
and U39117 (N_39117,N_25749,N_29463);
and U39118 (N_39118,N_24494,N_29866);
and U39119 (N_39119,N_29901,N_22116);
and U39120 (N_39120,N_21521,N_22767);
xnor U39121 (N_39121,N_27108,N_25124);
xnor U39122 (N_39122,N_29539,N_29592);
xor U39123 (N_39123,N_26220,N_26783);
and U39124 (N_39124,N_22832,N_28229);
nand U39125 (N_39125,N_24823,N_29195);
nand U39126 (N_39126,N_24943,N_22484);
nand U39127 (N_39127,N_25987,N_22177);
and U39128 (N_39128,N_25515,N_29180);
and U39129 (N_39129,N_24799,N_27662);
nand U39130 (N_39130,N_28859,N_20976);
or U39131 (N_39131,N_28866,N_28086);
nand U39132 (N_39132,N_29304,N_22571);
or U39133 (N_39133,N_25326,N_29989);
xor U39134 (N_39134,N_25591,N_25928);
and U39135 (N_39135,N_26946,N_29051);
xor U39136 (N_39136,N_21930,N_22521);
nand U39137 (N_39137,N_20336,N_20497);
or U39138 (N_39138,N_21174,N_21208);
or U39139 (N_39139,N_24071,N_29856);
and U39140 (N_39140,N_21993,N_22864);
nor U39141 (N_39141,N_25996,N_22992);
nor U39142 (N_39142,N_27792,N_22803);
or U39143 (N_39143,N_29339,N_21027);
nand U39144 (N_39144,N_20957,N_22199);
and U39145 (N_39145,N_28389,N_22827);
xnor U39146 (N_39146,N_23407,N_27356);
or U39147 (N_39147,N_28234,N_23083);
nor U39148 (N_39148,N_26890,N_26737);
xnor U39149 (N_39149,N_20094,N_29858);
or U39150 (N_39150,N_26359,N_24669);
or U39151 (N_39151,N_25171,N_26471);
and U39152 (N_39152,N_21368,N_25721);
nor U39153 (N_39153,N_22605,N_22985);
xor U39154 (N_39154,N_29315,N_22433);
nand U39155 (N_39155,N_23355,N_24579);
and U39156 (N_39156,N_23226,N_28740);
nor U39157 (N_39157,N_21771,N_23116);
nor U39158 (N_39158,N_22287,N_28290);
nor U39159 (N_39159,N_25343,N_23587);
nor U39160 (N_39160,N_24300,N_29997);
and U39161 (N_39161,N_27837,N_23703);
nor U39162 (N_39162,N_20143,N_21967);
or U39163 (N_39163,N_24340,N_27929);
nand U39164 (N_39164,N_20620,N_23632);
nand U39165 (N_39165,N_20769,N_29523);
or U39166 (N_39166,N_29961,N_28548);
or U39167 (N_39167,N_27947,N_29840);
nor U39168 (N_39168,N_24720,N_22817);
nor U39169 (N_39169,N_29181,N_27450);
or U39170 (N_39170,N_20054,N_22619);
and U39171 (N_39171,N_26498,N_26574);
and U39172 (N_39172,N_23496,N_25541);
nor U39173 (N_39173,N_27200,N_24992);
and U39174 (N_39174,N_27631,N_23697);
or U39175 (N_39175,N_23902,N_20618);
or U39176 (N_39176,N_20643,N_25869);
or U39177 (N_39177,N_26496,N_28357);
and U39178 (N_39178,N_29397,N_25506);
nand U39179 (N_39179,N_25273,N_28482);
nand U39180 (N_39180,N_25862,N_29150);
or U39181 (N_39181,N_21888,N_29630);
nand U39182 (N_39182,N_27355,N_27482);
and U39183 (N_39183,N_20746,N_21685);
nand U39184 (N_39184,N_27548,N_27593);
nand U39185 (N_39185,N_21213,N_27032);
or U39186 (N_39186,N_20016,N_24391);
or U39187 (N_39187,N_21992,N_25069);
nor U39188 (N_39188,N_24439,N_27361);
nand U39189 (N_39189,N_25697,N_24794);
and U39190 (N_39190,N_26777,N_23919);
nand U39191 (N_39191,N_21683,N_20272);
xor U39192 (N_39192,N_26933,N_23438);
nand U39193 (N_39193,N_25498,N_21585);
or U39194 (N_39194,N_28549,N_20594);
nor U39195 (N_39195,N_21946,N_26829);
nor U39196 (N_39196,N_20060,N_27139);
and U39197 (N_39197,N_22692,N_29756);
nor U39198 (N_39198,N_27324,N_27933);
and U39199 (N_39199,N_27041,N_20808);
xor U39200 (N_39200,N_27204,N_26781);
or U39201 (N_39201,N_21108,N_28658);
or U39202 (N_39202,N_22677,N_22876);
and U39203 (N_39203,N_23199,N_25387);
or U39204 (N_39204,N_29730,N_27163);
or U39205 (N_39205,N_24930,N_24288);
nand U39206 (N_39206,N_26117,N_27847);
nand U39207 (N_39207,N_20607,N_25802);
and U39208 (N_39208,N_23140,N_27077);
nor U39209 (N_39209,N_21975,N_20790);
nand U39210 (N_39210,N_28380,N_25515);
nand U39211 (N_39211,N_25499,N_23515);
nand U39212 (N_39212,N_29302,N_25684);
nor U39213 (N_39213,N_28598,N_22208);
xnor U39214 (N_39214,N_24602,N_23357);
nor U39215 (N_39215,N_23239,N_28539);
and U39216 (N_39216,N_24119,N_27491);
nand U39217 (N_39217,N_28453,N_24880);
nand U39218 (N_39218,N_25435,N_27745);
and U39219 (N_39219,N_20952,N_25672);
nand U39220 (N_39220,N_25340,N_22967);
xnor U39221 (N_39221,N_27863,N_24637);
or U39222 (N_39222,N_21128,N_23164);
nor U39223 (N_39223,N_28878,N_25327);
nand U39224 (N_39224,N_28858,N_29815);
or U39225 (N_39225,N_28454,N_20841);
nand U39226 (N_39226,N_26886,N_20431);
or U39227 (N_39227,N_24694,N_23728);
xnor U39228 (N_39228,N_23475,N_20725);
and U39229 (N_39229,N_22019,N_26748);
nand U39230 (N_39230,N_27665,N_23340);
nand U39231 (N_39231,N_20384,N_20463);
and U39232 (N_39232,N_23973,N_28389);
and U39233 (N_39233,N_27149,N_24247);
or U39234 (N_39234,N_20344,N_25401);
nor U39235 (N_39235,N_26250,N_28963);
nand U39236 (N_39236,N_24266,N_23552);
or U39237 (N_39237,N_21138,N_28962);
nor U39238 (N_39238,N_21074,N_22828);
and U39239 (N_39239,N_26415,N_24192);
xor U39240 (N_39240,N_24818,N_21453);
and U39241 (N_39241,N_25131,N_29450);
nand U39242 (N_39242,N_26004,N_21707);
and U39243 (N_39243,N_24086,N_22783);
nor U39244 (N_39244,N_20699,N_20640);
or U39245 (N_39245,N_25141,N_23733);
nor U39246 (N_39246,N_27079,N_21311);
nor U39247 (N_39247,N_27121,N_25128);
and U39248 (N_39248,N_21986,N_21492);
and U39249 (N_39249,N_26729,N_24675);
xnor U39250 (N_39250,N_23589,N_20881);
nand U39251 (N_39251,N_22695,N_27315);
or U39252 (N_39252,N_21304,N_29711);
and U39253 (N_39253,N_29103,N_20013);
nor U39254 (N_39254,N_28365,N_20962);
nor U39255 (N_39255,N_27982,N_21354);
or U39256 (N_39256,N_27763,N_23672);
nand U39257 (N_39257,N_20011,N_22087);
nand U39258 (N_39258,N_25275,N_20095);
nor U39259 (N_39259,N_29540,N_26978);
or U39260 (N_39260,N_21483,N_21531);
or U39261 (N_39261,N_24576,N_25505);
nor U39262 (N_39262,N_21184,N_21667);
or U39263 (N_39263,N_29914,N_23193);
and U39264 (N_39264,N_29356,N_25046);
or U39265 (N_39265,N_21158,N_28557);
nor U39266 (N_39266,N_20830,N_29959);
and U39267 (N_39267,N_24105,N_27358);
nand U39268 (N_39268,N_24826,N_27432);
nor U39269 (N_39269,N_28341,N_28937);
and U39270 (N_39270,N_25904,N_24093);
and U39271 (N_39271,N_24459,N_24889);
nand U39272 (N_39272,N_26449,N_27753);
and U39273 (N_39273,N_20198,N_28781);
and U39274 (N_39274,N_21020,N_29933);
nor U39275 (N_39275,N_21049,N_24159);
and U39276 (N_39276,N_20280,N_25990);
xor U39277 (N_39277,N_23668,N_25419);
and U39278 (N_39278,N_26411,N_28493);
or U39279 (N_39279,N_29372,N_24276);
nand U39280 (N_39280,N_29209,N_27296);
nor U39281 (N_39281,N_29258,N_29648);
or U39282 (N_39282,N_22938,N_23487);
and U39283 (N_39283,N_20513,N_29721);
or U39284 (N_39284,N_29946,N_22054);
or U39285 (N_39285,N_27185,N_29717);
nand U39286 (N_39286,N_26336,N_26569);
and U39287 (N_39287,N_27862,N_24877);
or U39288 (N_39288,N_20225,N_28758);
xor U39289 (N_39289,N_28214,N_29434);
nand U39290 (N_39290,N_26477,N_23592);
and U39291 (N_39291,N_28072,N_23289);
nor U39292 (N_39292,N_23378,N_22444);
xor U39293 (N_39293,N_28568,N_27792);
xor U39294 (N_39294,N_21303,N_20820);
or U39295 (N_39295,N_25714,N_20780);
nand U39296 (N_39296,N_25327,N_27219);
nor U39297 (N_39297,N_27612,N_28479);
xnor U39298 (N_39298,N_22064,N_25424);
nand U39299 (N_39299,N_28402,N_23625);
xor U39300 (N_39300,N_26639,N_20179);
nor U39301 (N_39301,N_22329,N_22689);
or U39302 (N_39302,N_29857,N_20872);
or U39303 (N_39303,N_23723,N_23137);
and U39304 (N_39304,N_27142,N_27437);
or U39305 (N_39305,N_24549,N_28900);
nor U39306 (N_39306,N_28291,N_28270);
or U39307 (N_39307,N_29516,N_23557);
nand U39308 (N_39308,N_26893,N_20042);
and U39309 (N_39309,N_28873,N_28625);
nor U39310 (N_39310,N_25888,N_21927);
or U39311 (N_39311,N_26109,N_24603);
xor U39312 (N_39312,N_23167,N_24614);
nor U39313 (N_39313,N_24940,N_28176);
and U39314 (N_39314,N_21664,N_28358);
and U39315 (N_39315,N_22119,N_23626);
nand U39316 (N_39316,N_21732,N_29800);
nor U39317 (N_39317,N_23881,N_29253);
and U39318 (N_39318,N_25245,N_23028);
or U39319 (N_39319,N_26966,N_28911);
xor U39320 (N_39320,N_23410,N_29469);
nand U39321 (N_39321,N_25116,N_25934);
nor U39322 (N_39322,N_26690,N_27285);
and U39323 (N_39323,N_26065,N_21218);
and U39324 (N_39324,N_23070,N_25921);
and U39325 (N_39325,N_26474,N_21389);
nor U39326 (N_39326,N_21573,N_25351);
xnor U39327 (N_39327,N_26552,N_29312);
nand U39328 (N_39328,N_21771,N_26325);
nor U39329 (N_39329,N_20529,N_25849);
nand U39330 (N_39330,N_20744,N_20336);
nand U39331 (N_39331,N_21313,N_25739);
xor U39332 (N_39332,N_25481,N_24326);
or U39333 (N_39333,N_21053,N_28862);
nor U39334 (N_39334,N_25075,N_25896);
nand U39335 (N_39335,N_24472,N_20375);
nor U39336 (N_39336,N_23741,N_25399);
or U39337 (N_39337,N_28923,N_20090);
and U39338 (N_39338,N_22132,N_29342);
xnor U39339 (N_39339,N_28562,N_23144);
nand U39340 (N_39340,N_23073,N_22122);
nand U39341 (N_39341,N_25933,N_22011);
and U39342 (N_39342,N_25586,N_24122);
nor U39343 (N_39343,N_21912,N_27155);
nor U39344 (N_39344,N_22011,N_26532);
nand U39345 (N_39345,N_26483,N_25307);
nand U39346 (N_39346,N_24276,N_23274);
nand U39347 (N_39347,N_21706,N_26691);
or U39348 (N_39348,N_24280,N_21928);
nand U39349 (N_39349,N_25430,N_25876);
or U39350 (N_39350,N_20433,N_22281);
or U39351 (N_39351,N_22058,N_25762);
nor U39352 (N_39352,N_28091,N_29863);
nor U39353 (N_39353,N_20924,N_22350);
or U39354 (N_39354,N_29299,N_20622);
or U39355 (N_39355,N_26013,N_25378);
nor U39356 (N_39356,N_24117,N_21083);
nor U39357 (N_39357,N_28848,N_23565);
xor U39358 (N_39358,N_29642,N_28440);
or U39359 (N_39359,N_22678,N_20147);
or U39360 (N_39360,N_25273,N_27486);
nand U39361 (N_39361,N_21117,N_25690);
or U39362 (N_39362,N_24379,N_21325);
or U39363 (N_39363,N_27341,N_28697);
nor U39364 (N_39364,N_20914,N_29390);
nor U39365 (N_39365,N_28799,N_29318);
nor U39366 (N_39366,N_28297,N_26978);
xor U39367 (N_39367,N_28183,N_24141);
xor U39368 (N_39368,N_26954,N_25686);
and U39369 (N_39369,N_28579,N_21218);
or U39370 (N_39370,N_22161,N_23332);
nand U39371 (N_39371,N_29317,N_21098);
xor U39372 (N_39372,N_20609,N_29984);
nor U39373 (N_39373,N_29106,N_23971);
nor U39374 (N_39374,N_29429,N_22119);
or U39375 (N_39375,N_25854,N_28289);
nand U39376 (N_39376,N_20376,N_28041);
or U39377 (N_39377,N_20867,N_21417);
and U39378 (N_39378,N_23717,N_24885);
or U39379 (N_39379,N_27888,N_23223);
and U39380 (N_39380,N_28738,N_24338);
nand U39381 (N_39381,N_27476,N_27283);
and U39382 (N_39382,N_21506,N_23839);
nand U39383 (N_39383,N_21148,N_24118);
xor U39384 (N_39384,N_28802,N_26479);
nand U39385 (N_39385,N_25296,N_25556);
and U39386 (N_39386,N_29659,N_22194);
nand U39387 (N_39387,N_27088,N_29200);
nor U39388 (N_39388,N_26860,N_21765);
and U39389 (N_39389,N_29457,N_29126);
or U39390 (N_39390,N_27125,N_29282);
or U39391 (N_39391,N_27504,N_21364);
nor U39392 (N_39392,N_28454,N_26173);
nand U39393 (N_39393,N_23141,N_22039);
nor U39394 (N_39394,N_29806,N_20450);
and U39395 (N_39395,N_23609,N_20465);
nand U39396 (N_39396,N_25411,N_22916);
and U39397 (N_39397,N_21644,N_27671);
xor U39398 (N_39398,N_29738,N_25779);
or U39399 (N_39399,N_25191,N_24114);
or U39400 (N_39400,N_27573,N_23820);
and U39401 (N_39401,N_21856,N_23810);
and U39402 (N_39402,N_25821,N_21505);
nor U39403 (N_39403,N_20526,N_21129);
and U39404 (N_39404,N_22849,N_25641);
nor U39405 (N_39405,N_21254,N_22982);
nor U39406 (N_39406,N_26398,N_27981);
xnor U39407 (N_39407,N_20642,N_29031);
or U39408 (N_39408,N_24522,N_25239);
and U39409 (N_39409,N_27930,N_23129);
nor U39410 (N_39410,N_24127,N_28636);
nor U39411 (N_39411,N_20726,N_21591);
and U39412 (N_39412,N_23101,N_21834);
nor U39413 (N_39413,N_22865,N_22920);
or U39414 (N_39414,N_23372,N_28595);
and U39415 (N_39415,N_24623,N_20881);
nor U39416 (N_39416,N_24719,N_20652);
nor U39417 (N_39417,N_28811,N_29505);
and U39418 (N_39418,N_28127,N_25249);
or U39419 (N_39419,N_22612,N_27896);
nor U39420 (N_39420,N_29880,N_20069);
nand U39421 (N_39421,N_20314,N_24471);
or U39422 (N_39422,N_23049,N_22109);
or U39423 (N_39423,N_26424,N_26374);
nor U39424 (N_39424,N_20498,N_26226);
nand U39425 (N_39425,N_20798,N_21230);
nand U39426 (N_39426,N_21004,N_29949);
and U39427 (N_39427,N_20835,N_25615);
nor U39428 (N_39428,N_22548,N_23817);
and U39429 (N_39429,N_25683,N_26817);
nand U39430 (N_39430,N_20884,N_29960);
and U39431 (N_39431,N_22277,N_24990);
or U39432 (N_39432,N_24646,N_29262);
or U39433 (N_39433,N_20204,N_25102);
or U39434 (N_39434,N_25469,N_29243);
or U39435 (N_39435,N_23398,N_20154);
nand U39436 (N_39436,N_20868,N_21442);
xor U39437 (N_39437,N_21582,N_28503);
nand U39438 (N_39438,N_27386,N_27449);
and U39439 (N_39439,N_24915,N_29499);
nor U39440 (N_39440,N_26936,N_22226);
or U39441 (N_39441,N_20962,N_24204);
nor U39442 (N_39442,N_24381,N_20298);
and U39443 (N_39443,N_25298,N_27521);
nand U39444 (N_39444,N_20321,N_20518);
nor U39445 (N_39445,N_27533,N_23032);
nor U39446 (N_39446,N_20632,N_24107);
xnor U39447 (N_39447,N_28527,N_28472);
and U39448 (N_39448,N_27635,N_26602);
xnor U39449 (N_39449,N_27754,N_24340);
or U39450 (N_39450,N_20309,N_24656);
nand U39451 (N_39451,N_24983,N_21335);
xnor U39452 (N_39452,N_28905,N_24125);
nand U39453 (N_39453,N_20437,N_29729);
and U39454 (N_39454,N_28721,N_27102);
or U39455 (N_39455,N_22964,N_21754);
xor U39456 (N_39456,N_25093,N_22093);
and U39457 (N_39457,N_21640,N_22916);
nand U39458 (N_39458,N_25956,N_29796);
or U39459 (N_39459,N_29484,N_23821);
or U39460 (N_39460,N_27385,N_28932);
or U39461 (N_39461,N_27667,N_25843);
xnor U39462 (N_39462,N_29334,N_26769);
or U39463 (N_39463,N_20378,N_22646);
nand U39464 (N_39464,N_25145,N_20612);
nand U39465 (N_39465,N_23188,N_20448);
or U39466 (N_39466,N_29763,N_21393);
or U39467 (N_39467,N_24710,N_29288);
nand U39468 (N_39468,N_25963,N_20312);
nor U39469 (N_39469,N_26974,N_26181);
and U39470 (N_39470,N_21825,N_20137);
nor U39471 (N_39471,N_21420,N_28232);
nand U39472 (N_39472,N_23027,N_24731);
and U39473 (N_39473,N_23321,N_21267);
and U39474 (N_39474,N_20758,N_22989);
nor U39475 (N_39475,N_23500,N_25106);
nand U39476 (N_39476,N_25728,N_21713);
xor U39477 (N_39477,N_20787,N_28629);
nand U39478 (N_39478,N_21048,N_21357);
nor U39479 (N_39479,N_26609,N_22580);
nor U39480 (N_39480,N_25712,N_29265);
nor U39481 (N_39481,N_25749,N_20821);
or U39482 (N_39482,N_22676,N_27428);
xor U39483 (N_39483,N_22492,N_29350);
xor U39484 (N_39484,N_24823,N_25103);
nor U39485 (N_39485,N_29163,N_24887);
nand U39486 (N_39486,N_26005,N_28056);
nand U39487 (N_39487,N_22140,N_28287);
or U39488 (N_39488,N_26807,N_24289);
and U39489 (N_39489,N_23547,N_21180);
nand U39490 (N_39490,N_21737,N_20156);
nor U39491 (N_39491,N_26992,N_23711);
nor U39492 (N_39492,N_22211,N_20661);
nor U39493 (N_39493,N_29353,N_20353);
and U39494 (N_39494,N_21283,N_25318);
nand U39495 (N_39495,N_21783,N_25329);
xnor U39496 (N_39496,N_20505,N_25863);
nand U39497 (N_39497,N_22324,N_27374);
nand U39498 (N_39498,N_22581,N_20629);
nand U39499 (N_39499,N_22392,N_27437);
nor U39500 (N_39500,N_20738,N_23088);
and U39501 (N_39501,N_26848,N_23176);
or U39502 (N_39502,N_23804,N_23044);
xor U39503 (N_39503,N_24919,N_27079);
or U39504 (N_39504,N_23052,N_23036);
nand U39505 (N_39505,N_27005,N_25091);
nor U39506 (N_39506,N_27266,N_22936);
xor U39507 (N_39507,N_20772,N_23329);
nor U39508 (N_39508,N_29721,N_29756);
and U39509 (N_39509,N_25635,N_24601);
xor U39510 (N_39510,N_20785,N_23269);
and U39511 (N_39511,N_28316,N_20903);
or U39512 (N_39512,N_29654,N_25222);
nor U39513 (N_39513,N_25026,N_24975);
or U39514 (N_39514,N_27396,N_23856);
nor U39515 (N_39515,N_25791,N_28303);
nand U39516 (N_39516,N_22801,N_23354);
nor U39517 (N_39517,N_28005,N_26240);
and U39518 (N_39518,N_21426,N_26498);
nor U39519 (N_39519,N_26304,N_24842);
or U39520 (N_39520,N_28240,N_21274);
xor U39521 (N_39521,N_26138,N_21319);
and U39522 (N_39522,N_28211,N_25809);
nand U39523 (N_39523,N_24544,N_25501);
or U39524 (N_39524,N_26359,N_20587);
nor U39525 (N_39525,N_22108,N_21830);
nand U39526 (N_39526,N_25029,N_29109);
nand U39527 (N_39527,N_25031,N_21347);
or U39528 (N_39528,N_22845,N_20317);
nor U39529 (N_39529,N_28851,N_23991);
and U39530 (N_39530,N_29511,N_26744);
and U39531 (N_39531,N_20292,N_23281);
or U39532 (N_39532,N_23346,N_20513);
and U39533 (N_39533,N_25820,N_29838);
nand U39534 (N_39534,N_23923,N_27710);
nor U39535 (N_39535,N_25073,N_25524);
nor U39536 (N_39536,N_22206,N_27117);
or U39537 (N_39537,N_25129,N_28597);
nand U39538 (N_39538,N_23535,N_29360);
or U39539 (N_39539,N_25809,N_20573);
xor U39540 (N_39540,N_22968,N_20726);
xnor U39541 (N_39541,N_25758,N_28217);
nor U39542 (N_39542,N_25862,N_26950);
and U39543 (N_39543,N_28444,N_28187);
xor U39544 (N_39544,N_26964,N_21772);
or U39545 (N_39545,N_27889,N_24864);
nand U39546 (N_39546,N_25974,N_22023);
nand U39547 (N_39547,N_20895,N_29596);
nor U39548 (N_39548,N_23352,N_22325);
and U39549 (N_39549,N_25393,N_29670);
and U39550 (N_39550,N_20132,N_28442);
xnor U39551 (N_39551,N_22287,N_23845);
or U39552 (N_39552,N_21861,N_27371);
and U39553 (N_39553,N_26921,N_25992);
or U39554 (N_39554,N_22748,N_25650);
nand U39555 (N_39555,N_22843,N_21286);
or U39556 (N_39556,N_29129,N_20102);
nand U39557 (N_39557,N_23084,N_26345);
nand U39558 (N_39558,N_29066,N_29833);
nand U39559 (N_39559,N_27323,N_24479);
nand U39560 (N_39560,N_28263,N_20239);
nand U39561 (N_39561,N_28503,N_24995);
nand U39562 (N_39562,N_23826,N_28877);
and U39563 (N_39563,N_23429,N_28576);
nand U39564 (N_39564,N_20713,N_27833);
or U39565 (N_39565,N_26659,N_22829);
nand U39566 (N_39566,N_22308,N_22411);
nand U39567 (N_39567,N_25508,N_28832);
nor U39568 (N_39568,N_26985,N_27369);
and U39569 (N_39569,N_22416,N_26018);
nand U39570 (N_39570,N_22011,N_22300);
or U39571 (N_39571,N_26279,N_24521);
and U39572 (N_39572,N_21590,N_21232);
and U39573 (N_39573,N_23786,N_21635);
or U39574 (N_39574,N_26395,N_28835);
nand U39575 (N_39575,N_24829,N_25327);
and U39576 (N_39576,N_24393,N_26902);
or U39577 (N_39577,N_27339,N_24816);
or U39578 (N_39578,N_25432,N_22186);
or U39579 (N_39579,N_21143,N_25490);
nor U39580 (N_39580,N_26652,N_20068);
nand U39581 (N_39581,N_26757,N_23644);
and U39582 (N_39582,N_20321,N_24402);
nor U39583 (N_39583,N_24298,N_26512);
or U39584 (N_39584,N_23854,N_23033);
and U39585 (N_39585,N_20790,N_26298);
nand U39586 (N_39586,N_22809,N_29222);
nor U39587 (N_39587,N_27269,N_28346);
and U39588 (N_39588,N_27911,N_24256);
or U39589 (N_39589,N_28851,N_25587);
or U39590 (N_39590,N_23380,N_28875);
and U39591 (N_39591,N_25054,N_27462);
and U39592 (N_39592,N_26759,N_20459);
nand U39593 (N_39593,N_27376,N_28239);
nand U39594 (N_39594,N_26170,N_24053);
and U39595 (N_39595,N_21552,N_26612);
nor U39596 (N_39596,N_26475,N_28423);
nand U39597 (N_39597,N_29147,N_28615);
nand U39598 (N_39598,N_21714,N_24143);
xor U39599 (N_39599,N_28905,N_21868);
nor U39600 (N_39600,N_20692,N_25600);
nor U39601 (N_39601,N_22083,N_22182);
and U39602 (N_39602,N_26503,N_24403);
or U39603 (N_39603,N_25585,N_21925);
xor U39604 (N_39604,N_27599,N_20119);
or U39605 (N_39605,N_20953,N_22285);
xnor U39606 (N_39606,N_29355,N_22819);
xnor U39607 (N_39607,N_24686,N_23313);
nor U39608 (N_39608,N_21989,N_22689);
or U39609 (N_39609,N_22064,N_23969);
or U39610 (N_39610,N_22834,N_20060);
and U39611 (N_39611,N_29699,N_24199);
nand U39612 (N_39612,N_24345,N_25086);
nand U39613 (N_39613,N_22719,N_28875);
xnor U39614 (N_39614,N_21502,N_29115);
and U39615 (N_39615,N_20602,N_28575);
and U39616 (N_39616,N_29850,N_28896);
or U39617 (N_39617,N_23405,N_26714);
nand U39618 (N_39618,N_27140,N_29124);
nand U39619 (N_39619,N_26193,N_24105);
nand U39620 (N_39620,N_26439,N_28874);
xor U39621 (N_39621,N_21773,N_23911);
nor U39622 (N_39622,N_21270,N_23601);
nand U39623 (N_39623,N_28368,N_20415);
or U39624 (N_39624,N_23830,N_24421);
nor U39625 (N_39625,N_26387,N_24323);
or U39626 (N_39626,N_27759,N_25925);
and U39627 (N_39627,N_28541,N_20592);
or U39628 (N_39628,N_21249,N_29957);
or U39629 (N_39629,N_24542,N_25943);
or U39630 (N_39630,N_28274,N_26597);
and U39631 (N_39631,N_29428,N_29192);
xor U39632 (N_39632,N_22333,N_26073);
or U39633 (N_39633,N_21791,N_29325);
nor U39634 (N_39634,N_20616,N_27097);
nand U39635 (N_39635,N_24965,N_20329);
nor U39636 (N_39636,N_20991,N_24498);
nor U39637 (N_39637,N_22959,N_21419);
nor U39638 (N_39638,N_29589,N_29207);
nand U39639 (N_39639,N_25479,N_28106);
or U39640 (N_39640,N_22015,N_28629);
nand U39641 (N_39641,N_25161,N_25419);
and U39642 (N_39642,N_21826,N_20664);
or U39643 (N_39643,N_22081,N_28623);
and U39644 (N_39644,N_22515,N_20740);
nor U39645 (N_39645,N_20019,N_25346);
and U39646 (N_39646,N_26837,N_23260);
and U39647 (N_39647,N_27826,N_27130);
and U39648 (N_39648,N_26504,N_26145);
and U39649 (N_39649,N_23158,N_23884);
or U39650 (N_39650,N_26609,N_23280);
and U39651 (N_39651,N_28882,N_27384);
nand U39652 (N_39652,N_24770,N_22281);
nor U39653 (N_39653,N_20702,N_21499);
or U39654 (N_39654,N_24561,N_20818);
nand U39655 (N_39655,N_27459,N_27465);
nand U39656 (N_39656,N_23350,N_23869);
and U39657 (N_39657,N_27272,N_24026);
nor U39658 (N_39658,N_23944,N_29942);
nor U39659 (N_39659,N_24498,N_26064);
and U39660 (N_39660,N_28457,N_24532);
nor U39661 (N_39661,N_27851,N_20465);
or U39662 (N_39662,N_26885,N_26002);
nor U39663 (N_39663,N_29685,N_26668);
and U39664 (N_39664,N_28493,N_24272);
or U39665 (N_39665,N_24386,N_21943);
or U39666 (N_39666,N_26509,N_25535);
and U39667 (N_39667,N_24252,N_22584);
nor U39668 (N_39668,N_27721,N_25816);
and U39669 (N_39669,N_25350,N_23368);
or U39670 (N_39670,N_27865,N_29311);
and U39671 (N_39671,N_20135,N_27249);
and U39672 (N_39672,N_20197,N_23766);
or U39673 (N_39673,N_26475,N_26807);
and U39674 (N_39674,N_28235,N_28895);
and U39675 (N_39675,N_26254,N_26212);
or U39676 (N_39676,N_28373,N_27208);
or U39677 (N_39677,N_26624,N_21965);
or U39678 (N_39678,N_28790,N_26461);
nor U39679 (N_39679,N_28100,N_23217);
nand U39680 (N_39680,N_21313,N_24389);
nand U39681 (N_39681,N_22930,N_29784);
xor U39682 (N_39682,N_26583,N_27426);
and U39683 (N_39683,N_21543,N_25943);
or U39684 (N_39684,N_27632,N_21217);
and U39685 (N_39685,N_25045,N_28106);
or U39686 (N_39686,N_23054,N_23943);
nor U39687 (N_39687,N_28686,N_26415);
and U39688 (N_39688,N_22477,N_24111);
or U39689 (N_39689,N_23906,N_28430);
or U39690 (N_39690,N_25811,N_22024);
xnor U39691 (N_39691,N_29540,N_29029);
nand U39692 (N_39692,N_22840,N_21224);
and U39693 (N_39693,N_21776,N_22932);
nand U39694 (N_39694,N_22738,N_29353);
and U39695 (N_39695,N_21697,N_29370);
and U39696 (N_39696,N_23532,N_21143);
or U39697 (N_39697,N_26370,N_24012);
or U39698 (N_39698,N_21393,N_25812);
and U39699 (N_39699,N_20841,N_20097);
and U39700 (N_39700,N_21022,N_21764);
nor U39701 (N_39701,N_27128,N_28069);
nor U39702 (N_39702,N_27984,N_29205);
nand U39703 (N_39703,N_29030,N_21843);
or U39704 (N_39704,N_27167,N_25496);
nor U39705 (N_39705,N_27793,N_24124);
xor U39706 (N_39706,N_27960,N_22928);
and U39707 (N_39707,N_24950,N_28804);
nand U39708 (N_39708,N_29391,N_28178);
and U39709 (N_39709,N_20987,N_29844);
or U39710 (N_39710,N_23351,N_24386);
nor U39711 (N_39711,N_28084,N_29917);
or U39712 (N_39712,N_29626,N_25889);
and U39713 (N_39713,N_26696,N_20976);
and U39714 (N_39714,N_21972,N_26938);
nor U39715 (N_39715,N_25550,N_22586);
and U39716 (N_39716,N_21055,N_20746);
nor U39717 (N_39717,N_26741,N_20179);
or U39718 (N_39718,N_29880,N_27427);
xnor U39719 (N_39719,N_21600,N_20270);
and U39720 (N_39720,N_27005,N_24667);
nand U39721 (N_39721,N_22079,N_23643);
and U39722 (N_39722,N_25503,N_24898);
and U39723 (N_39723,N_22008,N_22176);
nand U39724 (N_39724,N_26670,N_28801);
or U39725 (N_39725,N_25600,N_28061);
and U39726 (N_39726,N_26768,N_21461);
and U39727 (N_39727,N_21862,N_24541);
or U39728 (N_39728,N_28141,N_25068);
or U39729 (N_39729,N_27381,N_28230);
and U39730 (N_39730,N_20649,N_24763);
and U39731 (N_39731,N_21501,N_25344);
nand U39732 (N_39732,N_27086,N_20939);
or U39733 (N_39733,N_21533,N_22031);
xor U39734 (N_39734,N_23961,N_21766);
or U39735 (N_39735,N_23009,N_25719);
nor U39736 (N_39736,N_25845,N_29618);
and U39737 (N_39737,N_27011,N_28476);
and U39738 (N_39738,N_26717,N_27715);
or U39739 (N_39739,N_27620,N_26291);
and U39740 (N_39740,N_26534,N_28836);
and U39741 (N_39741,N_20413,N_23518);
and U39742 (N_39742,N_20866,N_20366);
nand U39743 (N_39743,N_25370,N_20865);
and U39744 (N_39744,N_28979,N_26414);
or U39745 (N_39745,N_26891,N_25703);
nor U39746 (N_39746,N_28732,N_25354);
or U39747 (N_39747,N_29363,N_24496);
and U39748 (N_39748,N_24153,N_20439);
nand U39749 (N_39749,N_28816,N_22362);
xor U39750 (N_39750,N_24986,N_27110);
nand U39751 (N_39751,N_29630,N_24005);
or U39752 (N_39752,N_21468,N_28769);
xnor U39753 (N_39753,N_28528,N_24179);
nand U39754 (N_39754,N_23107,N_25044);
nor U39755 (N_39755,N_29700,N_25479);
nor U39756 (N_39756,N_20579,N_22168);
and U39757 (N_39757,N_24618,N_29960);
nor U39758 (N_39758,N_26973,N_29780);
or U39759 (N_39759,N_29804,N_27252);
nand U39760 (N_39760,N_20326,N_28079);
nand U39761 (N_39761,N_24628,N_26900);
nand U39762 (N_39762,N_25968,N_28185);
or U39763 (N_39763,N_24853,N_22897);
nand U39764 (N_39764,N_22672,N_25778);
and U39765 (N_39765,N_26998,N_21152);
nor U39766 (N_39766,N_22788,N_27228);
and U39767 (N_39767,N_22490,N_25398);
or U39768 (N_39768,N_27764,N_20164);
nand U39769 (N_39769,N_20718,N_23015);
or U39770 (N_39770,N_22423,N_29035);
and U39771 (N_39771,N_27509,N_20618);
nor U39772 (N_39772,N_24364,N_21849);
or U39773 (N_39773,N_27877,N_29469);
xnor U39774 (N_39774,N_23038,N_26154);
nor U39775 (N_39775,N_27625,N_20622);
or U39776 (N_39776,N_20333,N_29346);
nand U39777 (N_39777,N_21701,N_23204);
nand U39778 (N_39778,N_27197,N_21898);
and U39779 (N_39779,N_23609,N_26092);
nand U39780 (N_39780,N_28045,N_26746);
nor U39781 (N_39781,N_25801,N_21904);
nand U39782 (N_39782,N_23848,N_23197);
nor U39783 (N_39783,N_29421,N_20468);
nand U39784 (N_39784,N_24899,N_26862);
or U39785 (N_39785,N_29632,N_29992);
and U39786 (N_39786,N_20240,N_23291);
or U39787 (N_39787,N_26601,N_27198);
or U39788 (N_39788,N_24999,N_25102);
xnor U39789 (N_39789,N_23842,N_20601);
and U39790 (N_39790,N_28514,N_25539);
and U39791 (N_39791,N_28335,N_26174);
nand U39792 (N_39792,N_28421,N_24086);
nand U39793 (N_39793,N_21950,N_21751);
nand U39794 (N_39794,N_26874,N_29252);
xor U39795 (N_39795,N_29299,N_25995);
and U39796 (N_39796,N_21404,N_24052);
and U39797 (N_39797,N_28083,N_27307);
nand U39798 (N_39798,N_21182,N_24849);
nand U39799 (N_39799,N_23318,N_21312);
nand U39800 (N_39800,N_25439,N_25569);
or U39801 (N_39801,N_24108,N_24319);
or U39802 (N_39802,N_23426,N_20911);
or U39803 (N_39803,N_26120,N_27664);
or U39804 (N_39804,N_29140,N_24129);
nand U39805 (N_39805,N_20890,N_29568);
xor U39806 (N_39806,N_23508,N_26104);
and U39807 (N_39807,N_29048,N_25731);
nand U39808 (N_39808,N_25869,N_26641);
nor U39809 (N_39809,N_20817,N_29807);
and U39810 (N_39810,N_26056,N_23781);
and U39811 (N_39811,N_29872,N_21161);
or U39812 (N_39812,N_22124,N_23245);
or U39813 (N_39813,N_26361,N_20570);
nor U39814 (N_39814,N_20741,N_26343);
or U39815 (N_39815,N_23274,N_22853);
nand U39816 (N_39816,N_25029,N_27974);
xor U39817 (N_39817,N_20880,N_23151);
nor U39818 (N_39818,N_23547,N_24582);
and U39819 (N_39819,N_24262,N_22401);
nor U39820 (N_39820,N_25765,N_26199);
and U39821 (N_39821,N_22892,N_29154);
xor U39822 (N_39822,N_22865,N_27203);
or U39823 (N_39823,N_26318,N_28933);
xor U39824 (N_39824,N_28001,N_26825);
and U39825 (N_39825,N_21795,N_22087);
nand U39826 (N_39826,N_20957,N_28953);
nor U39827 (N_39827,N_23469,N_27339);
and U39828 (N_39828,N_25912,N_20816);
nor U39829 (N_39829,N_23787,N_29846);
nand U39830 (N_39830,N_23035,N_21719);
nand U39831 (N_39831,N_28508,N_26166);
nor U39832 (N_39832,N_20575,N_22372);
or U39833 (N_39833,N_21674,N_26055);
nand U39834 (N_39834,N_20291,N_23017);
nand U39835 (N_39835,N_22428,N_25304);
and U39836 (N_39836,N_29548,N_23977);
nor U39837 (N_39837,N_25753,N_28173);
or U39838 (N_39838,N_23562,N_20908);
and U39839 (N_39839,N_22039,N_23698);
nor U39840 (N_39840,N_22125,N_27585);
and U39841 (N_39841,N_23673,N_20682);
nand U39842 (N_39842,N_29956,N_20275);
nand U39843 (N_39843,N_28595,N_27386);
xor U39844 (N_39844,N_27870,N_21523);
or U39845 (N_39845,N_25511,N_26765);
nand U39846 (N_39846,N_25741,N_29284);
nor U39847 (N_39847,N_24689,N_23478);
xor U39848 (N_39848,N_24011,N_28281);
xor U39849 (N_39849,N_29014,N_23011);
nor U39850 (N_39850,N_23060,N_21506);
nand U39851 (N_39851,N_23848,N_21664);
or U39852 (N_39852,N_25748,N_21622);
nand U39853 (N_39853,N_23729,N_21049);
or U39854 (N_39854,N_28175,N_27173);
or U39855 (N_39855,N_28867,N_26025);
nor U39856 (N_39856,N_23247,N_21945);
or U39857 (N_39857,N_27097,N_21318);
and U39858 (N_39858,N_20890,N_24802);
or U39859 (N_39859,N_26855,N_25936);
and U39860 (N_39860,N_27639,N_20268);
nor U39861 (N_39861,N_24076,N_22353);
or U39862 (N_39862,N_24122,N_20796);
nand U39863 (N_39863,N_28009,N_22879);
or U39864 (N_39864,N_21531,N_24627);
xor U39865 (N_39865,N_28242,N_20105);
or U39866 (N_39866,N_20561,N_29629);
nand U39867 (N_39867,N_20634,N_20007);
nor U39868 (N_39868,N_21970,N_27023);
nor U39869 (N_39869,N_20225,N_25643);
nor U39870 (N_39870,N_26051,N_25727);
nor U39871 (N_39871,N_23764,N_27333);
nand U39872 (N_39872,N_24893,N_28804);
nor U39873 (N_39873,N_26083,N_27863);
or U39874 (N_39874,N_28793,N_27309);
nor U39875 (N_39875,N_27632,N_21192);
nand U39876 (N_39876,N_21594,N_22214);
or U39877 (N_39877,N_27068,N_22921);
nand U39878 (N_39878,N_29727,N_20700);
and U39879 (N_39879,N_20229,N_20993);
or U39880 (N_39880,N_22826,N_27646);
or U39881 (N_39881,N_25831,N_21484);
nand U39882 (N_39882,N_25108,N_29480);
nand U39883 (N_39883,N_23137,N_23340);
or U39884 (N_39884,N_29788,N_20076);
xor U39885 (N_39885,N_29036,N_20209);
nand U39886 (N_39886,N_27621,N_20846);
nor U39887 (N_39887,N_25359,N_22395);
nor U39888 (N_39888,N_24790,N_24241);
xnor U39889 (N_39889,N_21212,N_25533);
nor U39890 (N_39890,N_20442,N_24926);
or U39891 (N_39891,N_23642,N_22943);
nand U39892 (N_39892,N_24582,N_28956);
xor U39893 (N_39893,N_25486,N_22701);
nor U39894 (N_39894,N_28097,N_27266);
xnor U39895 (N_39895,N_20540,N_27572);
nor U39896 (N_39896,N_29486,N_22349);
and U39897 (N_39897,N_28722,N_26196);
xnor U39898 (N_39898,N_21285,N_20631);
nor U39899 (N_39899,N_27949,N_26062);
nor U39900 (N_39900,N_26710,N_20554);
nor U39901 (N_39901,N_21316,N_25482);
or U39902 (N_39902,N_27134,N_20922);
nand U39903 (N_39903,N_24929,N_28454);
or U39904 (N_39904,N_21036,N_25795);
xnor U39905 (N_39905,N_26640,N_29460);
or U39906 (N_39906,N_23822,N_22244);
and U39907 (N_39907,N_27669,N_23467);
nor U39908 (N_39908,N_26436,N_28853);
or U39909 (N_39909,N_25349,N_24624);
or U39910 (N_39910,N_20270,N_25592);
nand U39911 (N_39911,N_21947,N_29554);
nand U39912 (N_39912,N_25053,N_22948);
xor U39913 (N_39913,N_29526,N_22004);
or U39914 (N_39914,N_23768,N_24578);
or U39915 (N_39915,N_25760,N_20780);
or U39916 (N_39916,N_25559,N_23133);
and U39917 (N_39917,N_29769,N_25595);
xor U39918 (N_39918,N_28525,N_22443);
nor U39919 (N_39919,N_21183,N_22261);
xnor U39920 (N_39920,N_28762,N_28048);
nand U39921 (N_39921,N_29339,N_25321);
nand U39922 (N_39922,N_21405,N_22232);
xnor U39923 (N_39923,N_25328,N_29222);
and U39924 (N_39924,N_20898,N_29861);
nand U39925 (N_39925,N_20538,N_26744);
xor U39926 (N_39926,N_26571,N_28196);
nand U39927 (N_39927,N_29222,N_20665);
xnor U39928 (N_39928,N_29928,N_21728);
nor U39929 (N_39929,N_24615,N_22096);
nand U39930 (N_39930,N_27416,N_29013);
nor U39931 (N_39931,N_22020,N_22921);
and U39932 (N_39932,N_24770,N_24738);
or U39933 (N_39933,N_26342,N_27696);
nand U39934 (N_39934,N_25035,N_25926);
and U39935 (N_39935,N_25971,N_20381);
nand U39936 (N_39936,N_28577,N_27086);
and U39937 (N_39937,N_23499,N_29876);
and U39938 (N_39938,N_20850,N_23293);
nand U39939 (N_39939,N_23651,N_23943);
nand U39940 (N_39940,N_25923,N_22927);
nand U39941 (N_39941,N_27073,N_28183);
or U39942 (N_39942,N_22621,N_27510);
and U39943 (N_39943,N_26057,N_23076);
or U39944 (N_39944,N_21927,N_21006);
or U39945 (N_39945,N_29738,N_20905);
nand U39946 (N_39946,N_29728,N_25796);
and U39947 (N_39947,N_24151,N_27384);
nor U39948 (N_39948,N_28003,N_25222);
nor U39949 (N_39949,N_28042,N_27415);
and U39950 (N_39950,N_25623,N_29911);
and U39951 (N_39951,N_26458,N_22934);
nand U39952 (N_39952,N_25181,N_28158);
nand U39953 (N_39953,N_29922,N_20707);
or U39954 (N_39954,N_23288,N_20718);
and U39955 (N_39955,N_24332,N_27567);
and U39956 (N_39956,N_24492,N_25658);
xnor U39957 (N_39957,N_24111,N_25503);
or U39958 (N_39958,N_25513,N_25432);
nor U39959 (N_39959,N_29611,N_29320);
or U39960 (N_39960,N_24545,N_22640);
and U39961 (N_39961,N_27105,N_29435);
nor U39962 (N_39962,N_26246,N_27228);
nor U39963 (N_39963,N_28797,N_24942);
nor U39964 (N_39964,N_21668,N_27803);
or U39965 (N_39965,N_25023,N_26517);
nor U39966 (N_39966,N_27427,N_28415);
or U39967 (N_39967,N_21376,N_24605);
nand U39968 (N_39968,N_20022,N_21642);
nor U39969 (N_39969,N_20162,N_28998);
xnor U39970 (N_39970,N_26665,N_24861);
nand U39971 (N_39971,N_26580,N_21450);
nand U39972 (N_39972,N_28303,N_20779);
or U39973 (N_39973,N_26289,N_27681);
and U39974 (N_39974,N_25600,N_20386);
or U39975 (N_39975,N_20513,N_27316);
and U39976 (N_39976,N_25996,N_24358);
nor U39977 (N_39977,N_29559,N_28422);
or U39978 (N_39978,N_28339,N_29737);
and U39979 (N_39979,N_20727,N_22518);
nor U39980 (N_39980,N_26663,N_25262);
or U39981 (N_39981,N_25102,N_28519);
nand U39982 (N_39982,N_24016,N_24683);
xnor U39983 (N_39983,N_23301,N_27635);
nand U39984 (N_39984,N_28836,N_25768);
and U39985 (N_39985,N_21725,N_26584);
nor U39986 (N_39986,N_28402,N_21438);
nand U39987 (N_39987,N_28182,N_22457);
or U39988 (N_39988,N_22602,N_29962);
and U39989 (N_39989,N_27793,N_25042);
or U39990 (N_39990,N_27826,N_29801);
nand U39991 (N_39991,N_20357,N_29624);
or U39992 (N_39992,N_28304,N_28356);
nand U39993 (N_39993,N_24415,N_29870);
nor U39994 (N_39994,N_26995,N_25538);
and U39995 (N_39995,N_23831,N_24919);
xor U39996 (N_39996,N_20563,N_21837);
nor U39997 (N_39997,N_29487,N_21093);
nor U39998 (N_39998,N_24396,N_25401);
nand U39999 (N_39999,N_29696,N_27473);
and U40000 (N_40000,N_30035,N_37375);
and U40001 (N_40001,N_34431,N_38330);
xor U40002 (N_40002,N_31013,N_30096);
and U40003 (N_40003,N_39521,N_32413);
nor U40004 (N_40004,N_36512,N_31270);
xnor U40005 (N_40005,N_35078,N_34411);
nor U40006 (N_40006,N_35017,N_32963);
nand U40007 (N_40007,N_32591,N_36131);
nor U40008 (N_40008,N_35836,N_31561);
nor U40009 (N_40009,N_31656,N_39483);
and U40010 (N_40010,N_31077,N_39164);
nor U40011 (N_40011,N_32682,N_38600);
xor U40012 (N_40012,N_35179,N_34438);
nand U40013 (N_40013,N_39095,N_30954);
nor U40014 (N_40014,N_32848,N_35526);
xor U40015 (N_40015,N_30131,N_34576);
nand U40016 (N_40016,N_35421,N_32106);
nor U40017 (N_40017,N_32240,N_35853);
and U40018 (N_40018,N_32687,N_31367);
or U40019 (N_40019,N_33303,N_35290);
or U40020 (N_40020,N_32596,N_37632);
or U40021 (N_40021,N_30106,N_31518);
or U40022 (N_40022,N_33708,N_34009);
nor U40023 (N_40023,N_32501,N_35630);
and U40024 (N_40024,N_38019,N_30217);
or U40025 (N_40025,N_33137,N_32298);
and U40026 (N_40026,N_33512,N_34304);
nand U40027 (N_40027,N_38265,N_34098);
or U40028 (N_40028,N_30143,N_39413);
nand U40029 (N_40029,N_31749,N_32456);
nor U40030 (N_40030,N_30592,N_33686);
nor U40031 (N_40031,N_36344,N_35164);
or U40032 (N_40032,N_36024,N_35690);
nand U40033 (N_40033,N_35909,N_38456);
and U40034 (N_40034,N_37137,N_36036);
or U40035 (N_40035,N_33481,N_39859);
xnor U40036 (N_40036,N_32764,N_36665);
or U40037 (N_40037,N_34151,N_33764);
nor U40038 (N_40038,N_32688,N_37393);
nor U40039 (N_40039,N_30620,N_32400);
and U40040 (N_40040,N_31381,N_37761);
nor U40041 (N_40041,N_32485,N_30610);
or U40042 (N_40042,N_38131,N_35639);
nand U40043 (N_40043,N_38542,N_32968);
nand U40044 (N_40044,N_31395,N_31993);
and U40045 (N_40045,N_30761,N_39353);
nor U40046 (N_40046,N_39469,N_38531);
or U40047 (N_40047,N_34114,N_31611);
and U40048 (N_40048,N_36772,N_37127);
nand U40049 (N_40049,N_32639,N_36763);
and U40050 (N_40050,N_38002,N_37297);
nor U40051 (N_40051,N_31834,N_38700);
or U40052 (N_40052,N_34000,N_35759);
and U40053 (N_40053,N_33462,N_37420);
and U40054 (N_40054,N_35934,N_37454);
nand U40055 (N_40055,N_30898,N_37073);
or U40056 (N_40056,N_30079,N_30296);
nand U40057 (N_40057,N_36566,N_37503);
nand U40058 (N_40058,N_30179,N_32630);
or U40059 (N_40059,N_32251,N_37923);
and U40060 (N_40060,N_35650,N_30308);
nor U40061 (N_40061,N_36474,N_39274);
nor U40062 (N_40062,N_31891,N_32593);
xor U40063 (N_40063,N_33328,N_39454);
nand U40064 (N_40064,N_37017,N_39330);
nand U40065 (N_40065,N_30501,N_33584);
nand U40066 (N_40066,N_36522,N_38721);
nor U40067 (N_40067,N_34691,N_33738);
or U40068 (N_40068,N_31553,N_33919);
nand U40069 (N_40069,N_35349,N_33711);
or U40070 (N_40070,N_38776,N_39770);
and U40071 (N_40071,N_33236,N_30187);
nor U40072 (N_40072,N_35578,N_32859);
nand U40073 (N_40073,N_39262,N_33573);
nand U40074 (N_40074,N_38029,N_34405);
xnor U40075 (N_40075,N_32262,N_31816);
or U40076 (N_40076,N_35027,N_33253);
xnor U40077 (N_40077,N_30137,N_35373);
nor U40078 (N_40078,N_33639,N_32601);
nor U40079 (N_40079,N_39529,N_39855);
and U40080 (N_40080,N_30013,N_39049);
and U40081 (N_40081,N_39899,N_34048);
and U40082 (N_40082,N_34131,N_38780);
xor U40083 (N_40083,N_36739,N_36765);
nor U40084 (N_40084,N_36506,N_39810);
nor U40085 (N_40085,N_37005,N_34232);
and U40086 (N_40086,N_39293,N_34121);
nand U40087 (N_40087,N_38098,N_32358);
nor U40088 (N_40088,N_31990,N_30981);
or U40089 (N_40089,N_33426,N_32884);
nor U40090 (N_40090,N_30684,N_35675);
or U40091 (N_40091,N_39908,N_30430);
and U40092 (N_40092,N_30972,N_39984);
nor U40093 (N_40093,N_30003,N_39787);
or U40094 (N_40094,N_39311,N_36050);
nand U40095 (N_40095,N_39923,N_39971);
nand U40096 (N_40096,N_32678,N_35080);
nand U40097 (N_40097,N_30538,N_36212);
or U40098 (N_40098,N_37765,N_34944);
nand U40099 (N_40099,N_36793,N_31578);
and U40100 (N_40100,N_33214,N_35165);
nand U40101 (N_40101,N_37576,N_33940);
or U40102 (N_40102,N_38351,N_39386);
nor U40103 (N_40103,N_37623,N_35978);
nor U40104 (N_40104,N_33716,N_30286);
nand U40105 (N_40105,N_33184,N_38285);
nor U40106 (N_40106,N_32081,N_37291);
or U40107 (N_40107,N_30568,N_30061);
nand U40108 (N_40108,N_32399,N_39786);
nor U40109 (N_40109,N_34979,N_31281);
nor U40110 (N_40110,N_37522,N_37519);
and U40111 (N_40111,N_36632,N_31681);
nor U40112 (N_40112,N_31564,N_36611);
and U40113 (N_40113,N_34213,N_38641);
xor U40114 (N_40114,N_38834,N_32608);
and U40115 (N_40115,N_31207,N_35443);
or U40116 (N_40116,N_34991,N_30253);
nand U40117 (N_40117,N_30526,N_39423);
xor U40118 (N_40118,N_31256,N_30313);
and U40119 (N_40119,N_32158,N_30085);
or U40120 (N_40120,N_30874,N_33801);
nand U40121 (N_40121,N_37965,N_31980);
nor U40122 (N_40122,N_30589,N_36752);
or U40123 (N_40123,N_36390,N_35167);
and U40124 (N_40124,N_39146,N_34189);
xor U40125 (N_40125,N_34473,N_36549);
or U40126 (N_40126,N_35082,N_35045);
nand U40127 (N_40127,N_37081,N_37372);
nand U40128 (N_40128,N_31677,N_33208);
nor U40129 (N_40129,N_36931,N_37777);
nor U40130 (N_40130,N_35730,N_35516);
nand U40131 (N_40131,N_36110,N_36424);
xor U40132 (N_40132,N_36247,N_36456);
and U40133 (N_40133,N_34280,N_34165);
and U40134 (N_40134,N_34519,N_36278);
nor U40135 (N_40135,N_34034,N_33658);
nand U40136 (N_40136,N_30181,N_31360);
nor U40137 (N_40137,N_32188,N_38473);
and U40138 (N_40138,N_37483,N_36238);
xor U40139 (N_40139,N_32294,N_34076);
or U40140 (N_40140,N_36400,N_33581);
or U40141 (N_40141,N_30897,N_30836);
or U40142 (N_40142,N_30483,N_32973);
nor U40143 (N_40143,N_30166,N_38913);
or U40144 (N_40144,N_38137,N_38328);
xnor U40145 (N_40145,N_30019,N_38711);
or U40146 (N_40146,N_38548,N_39410);
and U40147 (N_40147,N_31575,N_34770);
or U40148 (N_40148,N_36296,N_36918);
and U40149 (N_40149,N_38078,N_34577);
xor U40150 (N_40150,N_31587,N_34238);
and U40151 (N_40151,N_37129,N_35847);
xnor U40152 (N_40152,N_33792,N_38570);
and U40153 (N_40153,N_30361,N_33307);
nor U40154 (N_40154,N_37685,N_37424);
nand U40155 (N_40155,N_32161,N_38068);
nand U40156 (N_40156,N_37226,N_35766);
nor U40157 (N_40157,N_36115,N_30277);
xor U40158 (N_40158,N_38888,N_37981);
or U40159 (N_40159,N_34490,N_39734);
and U40160 (N_40160,N_34722,N_39664);
and U40161 (N_40161,N_35555,N_34790);
nor U40162 (N_40162,N_31524,N_36414);
and U40163 (N_40163,N_36147,N_37971);
xnor U40164 (N_40164,N_35928,N_34509);
or U40165 (N_40165,N_34791,N_32911);
nor U40166 (N_40166,N_35661,N_30665);
and U40167 (N_40167,N_35959,N_36286);
and U40168 (N_40168,N_33650,N_39148);
xor U40169 (N_40169,N_36895,N_39357);
and U40170 (N_40170,N_32722,N_33619);
or U40171 (N_40171,N_34475,N_39533);
nor U40172 (N_40172,N_36623,N_36649);
and U40173 (N_40173,N_39071,N_37224);
nand U40174 (N_40174,N_39507,N_30506);
nor U40175 (N_40175,N_36737,N_34161);
nand U40176 (N_40176,N_39307,N_30550);
nand U40177 (N_40177,N_31496,N_38490);
and U40178 (N_40178,N_35243,N_35037);
xnor U40179 (N_40179,N_39597,N_33321);
xnor U40180 (N_40180,N_31279,N_30698);
and U40181 (N_40181,N_33252,N_38237);
and U40182 (N_40182,N_37809,N_36472);
nand U40183 (N_40183,N_32763,N_39970);
nor U40184 (N_40184,N_31145,N_33380);
or U40185 (N_40185,N_37996,N_30237);
nand U40186 (N_40186,N_31512,N_34681);
xnor U40187 (N_40187,N_38587,N_38759);
or U40188 (N_40188,N_36799,N_37513);
and U40189 (N_40189,N_30261,N_31764);
and U40190 (N_40190,N_34402,N_37053);
or U40191 (N_40191,N_34983,N_31184);
and U40192 (N_40192,N_37292,N_37589);
and U40193 (N_40193,N_32468,N_39775);
nor U40194 (N_40194,N_32482,N_39047);
nor U40195 (N_40195,N_33829,N_33857);
nand U40196 (N_40196,N_36722,N_39061);
or U40197 (N_40197,N_30733,N_35881);
nand U40198 (N_40198,N_33483,N_33780);
nand U40199 (N_40199,N_38819,N_32843);
nor U40200 (N_40200,N_34541,N_33762);
or U40201 (N_40201,N_39150,N_39826);
nor U40202 (N_40202,N_36721,N_31300);
nand U40203 (N_40203,N_39275,N_35546);
nand U40204 (N_40204,N_36349,N_32786);
nor U40205 (N_40205,N_38563,N_32738);
or U40206 (N_40206,N_39869,N_38356);
xnor U40207 (N_40207,N_31694,N_30622);
nand U40208 (N_40208,N_30976,N_39324);
nand U40209 (N_40209,N_38442,N_36155);
nand U40210 (N_40210,N_38282,N_36294);
nor U40211 (N_40211,N_33398,N_38509);
nor U40212 (N_40212,N_34903,N_36425);
nor U40213 (N_40213,N_31495,N_36468);
nand U40214 (N_40214,N_37395,N_34959);
nand U40215 (N_40215,N_39480,N_38554);
and U40216 (N_40216,N_38879,N_34685);
and U40217 (N_40217,N_38872,N_31795);
or U40218 (N_40218,N_36555,N_36984);
nor U40219 (N_40219,N_32931,N_31594);
or U40220 (N_40220,N_30386,N_36006);
xor U40221 (N_40221,N_32905,N_35299);
nor U40222 (N_40222,N_34248,N_34588);
and U40223 (N_40223,N_32723,N_37075);
or U40224 (N_40224,N_39137,N_34228);
nor U40225 (N_40225,N_38412,N_33117);
and U40226 (N_40226,N_36987,N_35343);
and U40227 (N_40227,N_30887,N_36967);
or U40228 (N_40228,N_32919,N_39259);
nand U40229 (N_40229,N_31447,N_33505);
or U40230 (N_40230,N_32493,N_31627);
or U40231 (N_40231,N_34115,N_38231);
or U40232 (N_40232,N_34557,N_30011);
or U40233 (N_40233,N_38314,N_30616);
xnor U40234 (N_40234,N_31063,N_33926);
nor U40235 (N_40235,N_34286,N_39958);
or U40236 (N_40236,N_37662,N_32868);
and U40237 (N_40237,N_33977,N_39067);
or U40238 (N_40238,N_39182,N_35237);
or U40239 (N_40239,N_38226,N_34635);
nand U40240 (N_40240,N_38826,N_39607);
or U40241 (N_40241,N_39288,N_35742);
and U40242 (N_40242,N_34130,N_34297);
or U40243 (N_40243,N_33496,N_37116);
or U40244 (N_40244,N_36751,N_35328);
and U40245 (N_40245,N_37265,N_32010);
nand U40246 (N_40246,N_35529,N_38414);
nand U40247 (N_40247,N_39669,N_35034);
nor U40248 (N_40248,N_36417,N_37628);
nor U40249 (N_40249,N_39070,N_32402);
and U40250 (N_40250,N_33779,N_38470);
and U40251 (N_40251,N_31242,N_30212);
nand U40252 (N_40252,N_38153,N_32794);
nor U40253 (N_40253,N_35747,N_38723);
or U40254 (N_40254,N_33828,N_34057);
nor U40255 (N_40255,N_31630,N_34898);
and U40256 (N_40256,N_35504,N_33622);
nor U40257 (N_40257,N_30279,N_30602);
or U40258 (N_40258,N_32210,N_32088);
nand U40259 (N_40259,N_36143,N_38283);
nor U40260 (N_40260,N_30458,N_38033);
and U40261 (N_40261,N_34712,N_32713);
or U40262 (N_40262,N_31723,N_32921);
and U40263 (N_40263,N_38573,N_39737);
and U40264 (N_40264,N_35713,N_32724);
or U40265 (N_40265,N_37376,N_32005);
and U40266 (N_40266,N_33185,N_31193);
or U40267 (N_40267,N_38457,N_33114);
or U40268 (N_40268,N_37888,N_30224);
and U40269 (N_40269,N_30312,N_39983);
nor U40270 (N_40270,N_39955,N_32292);
and U40271 (N_40271,N_36373,N_35607);
and U40272 (N_40272,N_31782,N_34615);
xnor U40273 (N_40273,N_31756,N_38064);
nand U40274 (N_40274,N_37221,N_30696);
or U40275 (N_40275,N_34016,N_34579);
nor U40276 (N_40276,N_39181,N_35732);
or U40277 (N_40277,N_32053,N_34327);
or U40278 (N_40278,N_37550,N_32375);
or U40279 (N_40279,N_31180,N_35790);
nor U40280 (N_40280,N_33673,N_34124);
nor U40281 (N_40281,N_31415,N_32389);
or U40282 (N_40282,N_35401,N_33823);
nand U40283 (N_40283,N_34224,N_36406);
nand U40284 (N_40284,N_31220,N_36090);
and U40285 (N_40285,N_30210,N_35022);
nand U40286 (N_40286,N_31488,N_39938);
nand U40287 (N_40287,N_36377,N_39657);
or U40288 (N_40288,N_39271,N_33778);
or U40289 (N_40289,N_34520,N_31954);
or U40290 (N_40290,N_31781,N_32462);
or U40291 (N_40291,N_35880,N_30334);
nand U40292 (N_40292,N_33286,N_30203);
nor U40293 (N_40293,N_34351,N_35266);
nand U40294 (N_40294,N_30243,N_39084);
or U40295 (N_40295,N_32404,N_37054);
and U40296 (N_40296,N_35685,N_30080);
nor U40297 (N_40297,N_34760,N_31039);
and U40298 (N_40298,N_31282,N_33702);
nand U40299 (N_40299,N_35883,N_33467);
and U40300 (N_40300,N_38762,N_33485);
nor U40301 (N_40301,N_37274,N_39997);
or U40302 (N_40302,N_34994,N_37910);
nand U40303 (N_40303,N_32187,N_32508);
or U40304 (N_40304,N_36114,N_39540);
nor U40305 (N_40305,N_34394,N_31659);
and U40306 (N_40306,N_33032,N_39765);
or U40307 (N_40307,N_37964,N_33938);
and U40308 (N_40308,N_30030,N_31854);
or U40309 (N_40309,N_39819,N_34245);
and U40310 (N_40310,N_37658,N_34060);
nand U40311 (N_40311,N_34075,N_39270);
nor U40312 (N_40312,N_36317,N_35293);
nor U40313 (N_40313,N_35859,N_37686);
or U40314 (N_40314,N_30824,N_30051);
xnor U40315 (N_40315,N_38656,N_36943);
nor U40316 (N_40316,N_35274,N_32787);
or U40317 (N_40317,N_39823,N_39717);
nand U40318 (N_40318,N_33074,N_33067);
xor U40319 (N_40319,N_38169,N_39367);
and U40320 (N_40320,N_39728,N_30452);
and U40321 (N_40321,N_38165,N_35162);
and U40322 (N_40322,N_38520,N_31684);
and U40323 (N_40323,N_39509,N_38427);
nand U40324 (N_40324,N_38949,N_37443);
xor U40325 (N_40325,N_39013,N_36808);
and U40326 (N_40326,N_39566,N_38950);
nand U40327 (N_40327,N_31427,N_30886);
nand U40328 (N_40328,N_30453,N_31002);
nor U40329 (N_40329,N_37230,N_33755);
nand U40330 (N_40330,N_38448,N_30326);
and U40331 (N_40331,N_32539,N_30401);
nor U40332 (N_40332,N_39650,N_35550);
and U40333 (N_40333,N_33900,N_33627);
and U40334 (N_40334,N_30941,N_36382);
nand U40335 (N_40335,N_36375,N_39914);
nand U40336 (N_40336,N_35579,N_36378);
and U40337 (N_40337,N_39282,N_36308);
and U40338 (N_40338,N_37485,N_35355);
xor U40339 (N_40339,N_31176,N_30125);
and U40340 (N_40340,N_34477,N_39986);
and U40341 (N_40341,N_37323,N_32168);
xor U40342 (N_40342,N_32633,N_30147);
nor U40343 (N_40343,N_34470,N_33883);
and U40344 (N_40344,N_32813,N_33172);
or U40345 (N_40345,N_35851,N_37568);
xor U40346 (N_40346,N_32385,N_36023);
nand U40347 (N_40347,N_31419,N_30764);
xnor U40348 (N_40348,N_39504,N_33547);
nand U40349 (N_40349,N_37653,N_31346);
or U40350 (N_40350,N_39021,N_35007);
or U40351 (N_40351,N_39172,N_39045);
xor U40352 (N_40352,N_38049,N_35030);
or U40353 (N_40353,N_34779,N_38239);
nand U40354 (N_40354,N_31321,N_30017);
and U40355 (N_40355,N_34456,N_37931);
or U40356 (N_40356,N_33843,N_39940);
nand U40357 (N_40357,N_39985,N_39881);
xor U40358 (N_40358,N_31972,N_37937);
or U40359 (N_40359,N_38758,N_39860);
xor U40360 (N_40360,N_32094,N_39889);
or U40361 (N_40361,N_37108,N_34739);
or U40362 (N_40362,N_35569,N_32906);
and U40363 (N_40363,N_36591,N_30488);
nor U40364 (N_40364,N_34601,N_31956);
or U40365 (N_40365,N_38280,N_35760);
nand U40366 (N_40366,N_36836,N_34489);
or U40367 (N_40367,N_32904,N_30491);
nor U40368 (N_40368,N_34278,N_38610);
and U40369 (N_40369,N_38751,N_37115);
or U40370 (N_40370,N_36438,N_39924);
nand U40371 (N_40371,N_37235,N_32397);
and U40372 (N_40372,N_39063,N_34073);
and U40373 (N_40373,N_31873,N_35321);
nor U40374 (N_40374,N_33712,N_32945);
or U40375 (N_40375,N_39605,N_33125);
and U40376 (N_40376,N_35455,N_35564);
xnor U40377 (N_40377,N_39265,N_39694);
xor U40378 (N_40378,N_39600,N_39455);
and U40379 (N_40379,N_39651,N_39906);
nor U40380 (N_40380,N_32204,N_35408);
nor U40381 (N_40381,N_38901,N_32825);
nand U40382 (N_40382,N_39012,N_38404);
and U40383 (N_40383,N_34525,N_39493);
xnor U40384 (N_40384,N_30177,N_37110);
and U40385 (N_40385,N_35374,N_35895);
nor U40386 (N_40386,N_38316,N_31239);
or U40387 (N_40387,N_30412,N_38381);
nand U40388 (N_40388,N_32167,N_33341);
nand U40389 (N_40389,N_32257,N_37881);
or U40390 (N_40390,N_38774,N_38887);
or U40391 (N_40391,N_36507,N_36600);
nand U40392 (N_40392,N_37473,N_35496);
or U40393 (N_40393,N_35268,N_34293);
xor U40394 (N_40394,N_30427,N_38478);
nor U40395 (N_40395,N_37798,N_33043);
or U40396 (N_40396,N_30123,N_38366);
nor U40397 (N_40397,N_36015,N_39750);
or U40398 (N_40398,N_33265,N_37247);
and U40399 (N_40399,N_37864,N_39263);
or U40400 (N_40400,N_37456,N_36633);
and U40401 (N_40401,N_39977,N_34140);
nor U40402 (N_40402,N_37835,N_36051);
nor U40403 (N_40403,N_35036,N_34564);
nor U40404 (N_40404,N_37386,N_38468);
xnor U40405 (N_40405,N_34428,N_39705);
and U40406 (N_40406,N_33661,N_30970);
nor U40407 (N_40407,N_37228,N_38869);
or U40408 (N_40408,N_30160,N_38926);
or U40409 (N_40409,N_35269,N_30282);
nor U40410 (N_40410,N_37222,N_33081);
nor U40411 (N_40411,N_39348,N_31820);
nor U40412 (N_40412,N_30877,N_36666);
nand U40413 (N_40413,N_38865,N_32083);
nand U40414 (N_40414,N_39671,N_31964);
nor U40415 (N_40415,N_31821,N_30745);
and U40416 (N_40416,N_30033,N_36654);
nor U40417 (N_40417,N_30194,N_34384);
or U40418 (N_40418,N_35271,N_34782);
nor U40419 (N_40419,N_37079,N_32225);
and U40420 (N_40420,N_38939,N_30139);
and U40421 (N_40421,N_31500,N_37878);
nor U40422 (N_40422,N_35427,N_38584);
nor U40423 (N_40423,N_31535,N_33934);
nor U40424 (N_40424,N_34247,N_30206);
nand U40425 (N_40425,N_39406,N_30182);
or U40426 (N_40426,N_32031,N_37242);
xor U40427 (N_40427,N_31453,N_31895);
nor U40428 (N_40428,N_37409,N_38281);
nand U40429 (N_40429,N_38270,N_36615);
nor U40430 (N_40430,N_31464,N_34697);
and U40431 (N_40431,N_39018,N_35768);
nor U40432 (N_40432,N_32135,N_34409);
or U40433 (N_40433,N_35485,N_30278);
and U40434 (N_40434,N_30374,N_37250);
or U40435 (N_40435,N_32234,N_35326);
nand U40436 (N_40436,N_34330,N_33066);
nand U40437 (N_40437,N_32394,N_37870);
nor U40438 (N_40438,N_37603,N_33723);
or U40439 (N_40439,N_31605,N_39450);
nand U40440 (N_40440,N_32506,N_30032);
nor U40441 (N_40441,N_35971,N_34605);
and U40442 (N_40442,N_35175,N_34969);
or U40443 (N_40443,N_34391,N_37970);
nand U40444 (N_40444,N_38529,N_37924);
or U40445 (N_40445,N_34480,N_35081);
and U40446 (N_40446,N_31084,N_30964);
or U40447 (N_40447,N_38426,N_35487);
or U40448 (N_40448,N_38824,N_38208);
nor U40449 (N_40449,N_33869,N_32245);
nor U40450 (N_40450,N_36769,N_31865);
or U40451 (N_40451,N_39967,N_34478);
nor U40452 (N_40452,N_39690,N_31966);
and U40453 (N_40453,N_38747,N_38012);
nor U40454 (N_40454,N_35296,N_31758);
and U40455 (N_40455,N_38923,N_35762);
or U40456 (N_40456,N_37731,N_31014);
nand U40457 (N_40457,N_38393,N_30633);
or U40458 (N_40458,N_39277,N_32272);
and U40459 (N_40459,N_30304,N_38632);
nor U40460 (N_40460,N_32524,N_33620);
xor U40461 (N_40461,N_35926,N_36476);
or U40462 (N_40462,N_36441,N_30405);
nor U40463 (N_40463,N_37355,N_36260);
nor U40464 (N_40464,N_35594,N_39165);
and U40465 (N_40465,N_35581,N_37308);
or U40466 (N_40466,N_31460,N_38555);
or U40467 (N_40467,N_37548,N_39517);
nand U40468 (N_40468,N_30801,N_39851);
nor U40469 (N_40469,N_38994,N_32479);
nor U40470 (N_40470,N_33083,N_31499);
nor U40471 (N_40471,N_37669,N_32387);
and U40472 (N_40472,N_35478,N_32130);
nand U40473 (N_40473,N_30482,N_30196);
nand U40474 (N_40474,N_31147,N_36081);
nor U40475 (N_40475,N_36599,N_33490);
or U40476 (N_40476,N_38942,N_33082);
and U40477 (N_40477,N_38532,N_30363);
nand U40478 (N_40478,N_36239,N_32883);
xnor U40479 (N_40479,N_31296,N_34925);
nor U40480 (N_40480,N_34479,N_31451);
nand U40481 (N_40481,N_36264,N_36069);
or U40482 (N_40482,N_31588,N_35431);
and U40483 (N_40483,N_31910,N_32636);
and U40484 (N_40484,N_34310,N_33211);
and U40485 (N_40485,N_31958,N_34665);
or U40486 (N_40486,N_34290,N_30800);
nor U40487 (N_40487,N_31526,N_32316);
or U40488 (N_40488,N_37943,N_37905);
and U40489 (N_40489,N_36647,N_31480);
nand U40490 (N_40490,N_37883,N_37190);
or U40491 (N_40491,N_39863,N_33478);
nand U40492 (N_40492,N_39171,N_38032);
or U40493 (N_40493,N_32638,N_39833);
or U40494 (N_40494,N_32138,N_35003);
nand U40495 (N_40495,N_30846,N_31201);
xnor U40496 (N_40496,N_37067,N_37392);
or U40497 (N_40497,N_31770,N_35043);
or U40498 (N_40498,N_36053,N_34381);
or U40499 (N_40499,N_38562,N_32237);
or U40500 (N_40500,N_34938,N_30343);
xor U40501 (N_40501,N_35962,N_33429);
nand U40502 (N_40502,N_37475,N_36078);
xnor U40503 (N_40503,N_36746,N_36126);
or U40504 (N_40504,N_37026,N_36891);
nand U40505 (N_40505,N_33930,N_30664);
or U40506 (N_40506,N_37369,N_35014);
xor U40507 (N_40507,N_36650,N_30931);
nor U40508 (N_40508,N_37098,N_31604);
or U40509 (N_40509,N_35388,N_37529);
nand U40510 (N_40510,N_35955,N_33128);
nor U40511 (N_40511,N_32957,N_30637);
or U40512 (N_40512,N_30925,N_34641);
and U40513 (N_40513,N_33342,N_36004);
nand U40514 (N_40514,N_34514,N_39805);
nand U40515 (N_40515,N_33245,N_31926);
xnor U40516 (N_40516,N_31102,N_32747);
or U40517 (N_40517,N_33442,N_35429);
and U40518 (N_40518,N_35131,N_31273);
or U40519 (N_40519,N_31338,N_33713);
nand U40520 (N_40520,N_35907,N_35552);
nand U40521 (N_40521,N_36365,N_39407);
nor U40522 (N_40522,N_30345,N_30226);
or U40523 (N_40523,N_33155,N_38850);
nand U40524 (N_40524,N_39228,N_32117);
and U40525 (N_40525,N_30805,N_32829);
and U40526 (N_40526,N_38685,N_32132);
nor U40527 (N_40527,N_37799,N_35674);
and U40528 (N_40528,N_34112,N_37492);
nor U40529 (N_40529,N_30070,N_33873);
or U40530 (N_40530,N_32147,N_39359);
nand U40531 (N_40531,N_30281,N_35994);
and U40532 (N_40532,N_30650,N_35451);
xnor U40533 (N_40533,N_34550,N_33129);
xor U40534 (N_40534,N_38228,N_39317);
nand U40535 (N_40535,N_33048,N_38255);
nand U40536 (N_40536,N_34415,N_33116);
nor U40537 (N_40537,N_35277,N_33413);
nor U40538 (N_40538,N_35954,N_37215);
nand U40539 (N_40539,N_34659,N_35310);
nand U40540 (N_40540,N_32249,N_37240);
nor U40541 (N_40541,N_31371,N_33021);
and U40542 (N_40542,N_33008,N_32112);
or U40543 (N_40543,N_35035,N_33835);
and U40544 (N_40544,N_39088,N_36869);
or U40545 (N_40545,N_36258,N_39168);
or U40546 (N_40546,N_36451,N_30913);
nor U40547 (N_40547,N_36782,N_36346);
or U40548 (N_40548,N_39388,N_34045);
nor U40549 (N_40549,N_31301,N_35775);
or U40550 (N_40550,N_33529,N_30499);
or U40551 (N_40551,N_37408,N_36343);
or U40552 (N_40552,N_38771,N_34137);
or U40553 (N_40553,N_37212,N_31863);
nand U40554 (N_40554,N_32808,N_35459);
and U40555 (N_40555,N_33097,N_30197);
nor U40556 (N_40556,N_33545,N_37299);
xor U40557 (N_40557,N_32109,N_34718);
nand U40558 (N_40558,N_31101,N_37004);
nand U40559 (N_40559,N_33502,N_38207);
or U40560 (N_40560,N_35830,N_36152);
and U40561 (N_40561,N_31051,N_30344);
xor U40562 (N_40562,N_33501,N_30697);
or U40563 (N_40563,N_30702,N_37122);
xnor U40564 (N_40564,N_39877,N_37402);
or U40565 (N_40565,N_35769,N_32324);
nor U40566 (N_40566,N_39094,N_39358);
or U40567 (N_40567,N_32562,N_38586);
and U40568 (N_40568,N_32996,N_37302);
nand U40569 (N_40569,N_30302,N_39815);
or U40570 (N_40570,N_38968,N_34393);
or U40571 (N_40571,N_37535,N_39489);
and U40572 (N_40572,N_38161,N_37480);
xor U40573 (N_40573,N_31421,N_35272);
or U40574 (N_40574,N_37705,N_30722);
nand U40575 (N_40575,N_33663,N_32208);
xor U40576 (N_40576,N_32431,N_39552);
nor U40577 (N_40577,N_34963,N_39204);
or U40578 (N_40578,N_34754,N_31787);
nand U40579 (N_40579,N_35450,N_31801);
nor U40580 (N_40580,N_34007,N_37332);
nor U40581 (N_40581,N_34933,N_36690);
nand U40582 (N_40582,N_37739,N_39890);
and U40583 (N_40583,N_37734,N_39156);
nor U40584 (N_40584,N_39804,N_30958);
and U40585 (N_40585,N_39485,N_39347);
nand U40586 (N_40586,N_36289,N_30882);
or U40587 (N_40587,N_36055,N_34749);
and U40588 (N_40588,N_39298,N_31846);
and U40589 (N_40589,N_38992,N_30821);
or U40590 (N_40590,N_37146,N_32785);
or U40591 (N_40591,N_37521,N_37134);
nor U40592 (N_40592,N_38648,N_36319);
nor U40593 (N_40593,N_31040,N_37732);
nand U40594 (N_40594,N_31823,N_31602);
and U40595 (N_40595,N_39355,N_38638);
and U40596 (N_40596,N_33258,N_34709);
or U40597 (N_40597,N_32133,N_36059);
nor U40598 (N_40598,N_36563,N_34485);
or U40599 (N_40599,N_38243,N_32614);
nor U40600 (N_40600,N_34631,N_30256);
xor U40601 (N_40601,N_36983,N_35643);
and U40602 (N_40602,N_31502,N_33741);
and U40603 (N_40603,N_34211,N_31023);
nand U40604 (N_40604,N_39046,N_35028);
or U40605 (N_40605,N_33243,N_39640);
nand U40606 (N_40606,N_35291,N_32391);
nor U40607 (N_40607,N_34690,N_39539);
or U40608 (N_40608,N_34798,N_38496);
xor U40609 (N_40609,N_33968,N_31977);
or U40610 (N_40610,N_38545,N_34044);
xnor U40611 (N_40611,N_32664,N_37565);
nand U40612 (N_40612,N_35996,N_33783);
nor U40613 (N_40613,N_35869,N_32617);
or U40614 (N_40614,N_32801,N_38793);
or U40615 (N_40615,N_30672,N_33308);
nor U40616 (N_40616,N_37484,N_32836);
or U40617 (N_40617,N_39594,N_35542);
or U40618 (N_40618,N_35322,N_31728);
nor U40619 (N_40619,N_34314,N_34939);
nor U40620 (N_40620,N_30817,N_30744);
xor U40621 (N_40621,N_30849,N_38825);
nor U40622 (N_40622,N_30456,N_31329);
nand U40623 (N_40623,N_32733,N_33476);
or U40624 (N_40624,N_30460,N_34276);
nand U40625 (N_40625,N_31725,N_32611);
or U40626 (N_40626,N_32333,N_33434);
and U40627 (N_40627,N_32612,N_32929);
nand U40628 (N_40628,N_33012,N_35843);
and U40629 (N_40629,N_37326,N_36327);
or U40630 (N_40630,N_37135,N_34176);
and U40631 (N_40631,N_39767,N_35927);
and U40632 (N_40632,N_31845,N_37237);
and U40633 (N_40633,N_30539,N_31547);
xor U40634 (N_40634,N_31697,N_34664);
nand U40635 (N_40635,N_31736,N_31112);
nand U40636 (N_40636,N_38498,N_35295);
and U40637 (N_40637,N_34464,N_36538);
nor U40638 (N_40638,N_30251,N_35763);
and U40639 (N_40639,N_38295,N_31332);
nand U40640 (N_40640,N_33244,N_39237);
nor U40641 (N_40641,N_33503,N_35456);
or U40642 (N_40642,N_36577,N_38315);
and U40643 (N_40643,N_39989,N_35882);
xor U40644 (N_40644,N_34856,N_30792);
xnor U40645 (N_40645,N_37341,N_35966);
nor U40646 (N_40646,N_33039,N_37432);
nor U40647 (N_40647,N_38904,N_33385);
nand U40648 (N_40648,N_34323,N_35124);
nand U40649 (N_40649,N_32903,N_30000);
or U40650 (N_40650,N_34708,N_36570);
and U40651 (N_40651,N_36908,N_38508);
nand U40652 (N_40652,N_37902,N_37678);
nand U40653 (N_40653,N_39755,N_38613);
or U40654 (N_40654,N_39523,N_39167);
nand U40655 (N_40655,N_31456,N_33862);
xnor U40656 (N_40656,N_32365,N_37159);
nor U40657 (N_40657,N_35508,N_32232);
and U40658 (N_40658,N_34325,N_34077);
nand U40659 (N_40659,N_38201,N_39617);
and U40660 (N_40660,N_39127,N_30202);
or U40661 (N_40661,N_32100,N_33696);
or U40662 (N_40662,N_36035,N_35866);
xnor U40663 (N_40663,N_35292,N_37404);
nor U40664 (N_40664,N_34780,N_39720);
or U40665 (N_40665,N_34349,N_32725);
nand U40666 (N_40666,N_33087,N_39404);
or U40667 (N_40667,N_33844,N_30815);
nor U40668 (N_40668,N_31818,N_36704);
or U40669 (N_40669,N_33532,N_31142);
nor U40670 (N_40670,N_33292,N_33352);
or U40671 (N_40671,N_32831,N_34899);
or U40672 (N_40672,N_34904,N_37197);
xor U40673 (N_40673,N_38370,N_35621);
nor U40674 (N_40674,N_35090,N_36061);
and U40675 (N_40675,N_37904,N_36339);
nand U40676 (N_40676,N_35094,N_39223);
nor U40677 (N_40677,N_33974,N_38832);
nor U40678 (N_40678,N_35446,N_39788);
nor U40679 (N_40679,N_33774,N_36528);
nor U40680 (N_40680,N_34504,N_39588);
and U40681 (N_40681,N_32975,N_31850);
and U40682 (N_40682,N_33516,N_35772);
or U40683 (N_40683,N_36355,N_31640);
or U40684 (N_40684,N_30752,N_39211);
nor U40685 (N_40685,N_37216,N_36307);
nand U40686 (N_40686,N_37433,N_30566);
nor U40687 (N_40687,N_36466,N_32499);
xor U40688 (N_40688,N_34965,N_33717);
xnor U40689 (N_40689,N_33431,N_38856);
xor U40690 (N_40690,N_38848,N_35117);
and U40691 (N_40691,N_31260,N_39299);
nand U40692 (N_40692,N_37014,N_39030);
nor U40693 (N_40693,N_38059,N_38769);
and U40694 (N_40694,N_32940,N_33917);
and U40695 (N_40695,N_30227,N_31025);
or U40696 (N_40696,N_33405,N_38090);
and U40697 (N_40697,N_34862,N_32422);
nor U40698 (N_40698,N_36246,N_34460);
and U40699 (N_40699,N_30642,N_30574);
or U40700 (N_40700,N_32148,N_39460);
nor U40701 (N_40701,N_39898,N_35976);
nand U40702 (N_40702,N_33313,N_36595);
and U40703 (N_40703,N_34813,N_34420);
nand U40704 (N_40704,N_32806,N_31079);
or U40705 (N_40705,N_39696,N_30789);
or U40706 (N_40706,N_30741,N_30813);
nand U40707 (N_40707,N_33633,N_34955);
nand U40708 (N_40708,N_33446,N_30373);
or U40709 (N_40709,N_33302,N_30400);
nand U40710 (N_40710,N_38670,N_31652);
or U40711 (N_40711,N_36293,N_30023);
nand U40712 (N_40712,N_37142,N_34821);
xor U40713 (N_40713,N_38013,N_38698);
nor U40714 (N_40714,N_39139,N_33205);
and U40715 (N_40715,N_38911,N_30221);
and U40716 (N_40716,N_34972,N_32980);
nand U40717 (N_40717,N_38331,N_30284);
or U40718 (N_40718,N_33336,N_33075);
or U40719 (N_40719,N_36785,N_35749);
nand U40720 (N_40720,N_33450,N_33776);
and U40721 (N_40721,N_35188,N_30447);
nor U40722 (N_40722,N_36399,N_36454);
nor U40723 (N_40723,N_31716,N_31730);
nor U40724 (N_40724,N_33579,N_34296);
and U40725 (N_40725,N_34922,N_30324);
nor U40726 (N_40726,N_35780,N_38277);
nor U40727 (N_40727,N_34387,N_36240);
or U40728 (N_40728,N_38660,N_37549);
and U40729 (N_40729,N_36262,N_37874);
nand U40730 (N_40730,N_35437,N_35683);
or U40731 (N_40731,N_32475,N_34199);
or U40732 (N_40732,N_37940,N_39853);
nor U40733 (N_40733,N_36448,N_35734);
and U40734 (N_40734,N_30749,N_32832);
or U40735 (N_40735,N_37317,N_33850);
xnor U40736 (N_40736,N_34181,N_33894);
and U40737 (N_40737,N_39871,N_31059);
nor U40738 (N_40738,N_34989,N_37130);
nand U40739 (N_40739,N_37232,N_30442);
or U40740 (N_40740,N_37551,N_35577);
xor U40741 (N_40741,N_36612,N_33745);
or U40742 (N_40742,N_31223,N_32822);
or U40743 (N_40743,N_36826,N_37394);
or U40744 (N_40744,N_30119,N_33034);
nand U40745 (N_40745,N_32091,N_33599);
or U40746 (N_40746,N_38608,N_33424);
or U40747 (N_40747,N_39373,N_35362);
or U40748 (N_40748,N_38775,N_33720);
nand U40749 (N_40749,N_32882,N_34350);
nand U40750 (N_40750,N_36844,N_35612);
nor U40751 (N_40751,N_30659,N_32407);
xnor U40752 (N_40752,N_38307,N_36877);
or U40753 (N_40753,N_32648,N_36726);
nand U40754 (N_40754,N_35492,N_31890);
and U40755 (N_40755,N_30683,N_35916);
xnor U40756 (N_40756,N_36837,N_35828);
nor U40757 (N_40757,N_30480,N_31959);
or U40758 (N_40758,N_31856,N_34833);
nor U40759 (N_40759,N_30330,N_30393);
nand U40760 (N_40760,N_30057,N_30036);
xor U40761 (N_40761,N_34303,N_32338);
and U40762 (N_40762,N_38273,N_30703);
nor U40763 (N_40763,N_36594,N_37561);
nor U40764 (N_40764,N_34871,N_38804);
nor U40765 (N_40765,N_38664,N_30979);
xor U40766 (N_40766,N_35040,N_37198);
nand U40767 (N_40767,N_31937,N_36708);
or U40768 (N_40768,N_39099,N_33156);
nand U40769 (N_40769,N_31864,N_37806);
nand U40770 (N_40770,N_31635,N_34607);
nand U40771 (N_40771,N_39442,N_36149);
and U40772 (N_40772,N_39609,N_30149);
nor U40773 (N_40773,N_37337,N_39051);
or U40774 (N_40774,N_36927,N_30779);
nand U40775 (N_40775,N_38162,N_37173);
or U40776 (N_40776,N_37637,N_32477);
and U40777 (N_40777,N_38640,N_36700);
nor U40778 (N_40778,N_39350,N_38261);
nor U40779 (N_40779,N_38768,N_34295);
nand U40780 (N_40780,N_35434,N_39698);
and U40781 (N_40781,N_33173,N_31246);
and U40782 (N_40782,N_37241,N_34715);
nor U40783 (N_40783,N_37987,N_39474);
or U40784 (N_40784,N_33445,N_33528);
nor U40785 (N_40785,N_37692,N_32190);
nand U40786 (N_40786,N_38245,N_32784);
nor U40787 (N_40787,N_32156,N_35096);
nor U40788 (N_40788,N_36284,N_35309);
xnor U40789 (N_40789,N_33560,N_34229);
or U40790 (N_40790,N_36854,N_31747);
nor U40791 (N_40791,N_34670,N_33339);
or U40792 (N_40792,N_35778,N_36741);
and U40793 (N_40793,N_33928,N_35941);
nor U40794 (N_40794,N_38108,N_30780);
or U40795 (N_40795,N_32932,N_39843);
and U40796 (N_40796,N_35347,N_32029);
and U40797 (N_40797,N_32509,N_36960);
nand U40798 (N_40798,N_30729,N_39557);
and U40799 (N_40799,N_33559,N_33152);
and U40800 (N_40800,N_36010,N_39300);
and U40801 (N_40801,N_31359,N_35099);
nand U40802 (N_40802,N_34988,N_31546);
nor U40803 (N_40803,N_39463,N_36495);
xor U40804 (N_40804,N_30364,N_35826);
nand U40805 (N_40805,N_35327,N_34454);
or U40806 (N_40806,N_33188,N_32051);
or U40807 (N_40807,N_31508,N_39949);
nor U40808 (N_40808,N_33147,N_30375);
nand U40809 (N_40809,N_31600,N_37664);
nor U40810 (N_40810,N_39117,N_33605);
or U40811 (N_40811,N_37751,N_33903);
nor U40812 (N_40812,N_34164,N_39255);
and U40813 (N_40813,N_39092,N_34561);
or U40814 (N_40814,N_32283,N_33159);
nor U40815 (N_40815,N_31309,N_36883);
nand U40816 (N_40816,N_38881,N_35653);
or U40817 (N_40817,N_31898,N_32655);
and U40818 (N_40818,N_34103,N_33407);
and U40819 (N_40819,N_32511,N_35754);
or U40820 (N_40820,N_32126,N_34866);
or U40821 (N_40821,N_33914,N_31094);
and U40822 (N_40822,N_35886,N_39937);
or U40823 (N_40823,N_39361,N_30992);
and U40824 (N_40824,N_33488,N_30311);
or U40825 (N_40825,N_36613,N_33520);
nand U40826 (N_40826,N_34049,N_38061);
or U40827 (N_40827,N_39528,N_39935);
nor U40828 (N_40828,N_34653,N_33969);
or U40829 (N_40829,N_33606,N_30946);
xor U40830 (N_40830,N_39132,N_34037);
and U40831 (N_40831,N_36865,N_34182);
and U40832 (N_40832,N_38560,N_37536);
and U40833 (N_40833,N_35898,N_37357);
nor U40834 (N_40834,N_31516,N_34855);
nand U40835 (N_40835,N_33575,N_33091);
xnor U40836 (N_40836,N_36430,N_33314);
nor U40837 (N_40837,N_32544,N_38649);
xor U40838 (N_40838,N_35764,N_39880);
nand U40839 (N_40839,N_31325,N_31886);
or U40840 (N_40840,N_30810,N_31981);
and U40841 (N_40841,N_38304,N_38401);
and U40842 (N_40842,N_35797,N_34548);
nand U40843 (N_40843,N_33667,N_37507);
nand U40844 (N_40844,N_39443,N_38629);
nor U40845 (N_40845,N_34240,N_31775);
nor U40846 (N_40846,N_37306,N_39028);
nor U40847 (N_40847,N_34740,N_32307);
nand U40848 (N_40848,N_35056,N_32698);
nor U40849 (N_40849,N_31987,N_39456);
nand U40850 (N_40850,N_30916,N_37755);
xor U40851 (N_40851,N_30366,N_33199);
nor U40852 (N_40852,N_37969,N_33346);
nor U40853 (N_40853,N_38017,N_36652);
nand U40854 (N_40854,N_33127,N_31311);
or U40855 (N_40855,N_33798,N_33187);
nor U40856 (N_40856,N_39170,N_34800);
nand U40857 (N_40857,N_35918,N_31061);
nand U40858 (N_40858,N_32780,N_37677);
nor U40859 (N_40859,N_34643,N_34616);
and U40860 (N_40860,N_37416,N_32576);
or U40861 (N_40861,N_31996,N_38707);
nand U40862 (N_40862,N_34651,N_35260);
xor U40863 (N_40863,N_32287,N_34654);
nor U40864 (N_40864,N_32671,N_35284);
and U40865 (N_40865,N_36778,N_37151);
and U40866 (N_40866,N_33000,N_32683);
or U40867 (N_40867,N_33090,N_37626);
or U40868 (N_40868,N_36881,N_37253);
or U40869 (N_40869,N_30262,N_35925);
or U40870 (N_40870,N_36151,N_31336);
nor U40871 (N_40871,N_31024,N_32987);
nor U40872 (N_40872,N_31998,N_39603);
nand U40873 (N_40873,N_33811,N_39424);
xnor U40874 (N_40874,N_39105,N_38653);
nand U40875 (N_40875,N_35923,N_32068);
nand U40876 (N_40876,N_32119,N_31240);
or U40877 (N_40877,N_38871,N_38781);
or U40878 (N_40878,N_36391,N_37158);
and U40879 (N_40879,N_34015,N_31433);
and U40880 (N_40880,N_35225,N_31377);
or U40881 (N_40881,N_38658,N_32065);
nor U40882 (N_40882,N_32581,N_30504);
and U40883 (N_40883,N_38524,N_35795);
or U40884 (N_40884,N_34701,N_39356);
xor U40885 (N_40885,N_32271,N_31324);
xnor U40886 (N_40886,N_30287,N_30360);
nand U40887 (N_40887,N_32326,N_32924);
nor U40888 (N_40888,N_30930,N_32652);
nand U40889 (N_40889,N_30248,N_37699);
nand U40890 (N_40890,N_39554,N_36907);
nand U40891 (N_40891,N_38845,N_30638);
nand U40892 (N_40892,N_37907,N_35329);
or U40893 (N_40893,N_31933,N_32030);
or U40894 (N_40894,N_34743,N_39993);
nand U40895 (N_40895,N_31532,N_37205);
xor U40896 (N_40896,N_34021,N_39661);
xor U40897 (N_40897,N_38297,N_36887);
xor U40898 (N_40898,N_35738,N_35285);
or U40899 (N_40899,N_39441,N_30188);
nor U40900 (N_40900,N_36292,N_39128);
or U40901 (N_40901,N_38748,N_35313);
nor U40902 (N_40902,N_33094,N_33255);
nand U40903 (N_40903,N_33585,N_31394);
nand U40904 (N_40904,N_32626,N_38571);
nor U40905 (N_40905,N_39005,N_32420);
xor U40906 (N_40906,N_32052,N_39672);
nand U40907 (N_40907,N_33316,N_37153);
nand U40908 (N_40908,N_30632,N_30490);
nor U40909 (N_40909,N_30753,N_39447);
and U40910 (N_40910,N_32125,N_37175);
nor U40911 (N_40911,N_34817,N_32595);
nor U40912 (N_40912,N_33001,N_37103);
nor U40913 (N_40913,N_32571,N_38249);
xor U40914 (N_40914,N_37657,N_34522);
nand U40915 (N_40915,N_37783,N_31050);
xnor U40916 (N_40916,N_38892,N_35378);
nand U40917 (N_40917,N_36602,N_35518);
or U40918 (N_40918,N_34929,N_36054);
nor U40919 (N_40919,N_33115,N_32299);
or U40920 (N_40920,N_30865,N_34594);
nand U40921 (N_40921,N_30593,N_36221);
nand U40922 (N_40922,N_32111,N_31673);
and U40923 (N_40923,N_31724,N_39119);
nand U40924 (N_40924,N_39791,N_33109);
and U40925 (N_40925,N_39294,N_31667);
nor U40926 (N_40926,N_39905,N_33854);
or U40927 (N_40927,N_30514,N_38674);
and U40928 (N_40928,N_39152,N_30860);
or U40929 (N_40929,N_37199,N_34734);
xor U40930 (N_40930,N_32011,N_32536);
xor U40931 (N_40931,N_37763,N_36386);
nand U40932 (N_40932,N_30339,N_36223);
nand U40933 (N_40933,N_35619,N_36465);
and U40934 (N_40934,N_34311,N_39238);
or U40935 (N_40935,N_36331,N_38526);
or U40936 (N_40936,N_36838,N_31141);
or U40937 (N_40937,N_31169,N_37608);
and U40938 (N_40938,N_33274,N_35143);
nand U40939 (N_40939,N_38518,N_32563);
nand U40940 (N_40940,N_35058,N_37049);
nor U40941 (N_40941,N_32853,N_35116);
and U40942 (N_40942,N_36271,N_33694);
or U40943 (N_40943,N_32529,N_37973);
nand U40944 (N_40944,N_32640,N_31278);
and U40945 (N_40945,N_38242,N_34626);
and U40946 (N_40946,N_31137,N_37210);
and U40947 (N_40947,N_35668,N_35656);
nor U40948 (N_40948,N_39658,N_31151);
or U40949 (N_40949,N_37715,N_31041);
and U40950 (N_40950,N_36121,N_33383);
nand U40951 (N_40951,N_34656,N_31352);
nand U40952 (N_40952,N_38020,N_34756);
and U40953 (N_40953,N_37446,N_37155);
nand U40954 (N_40954,N_30688,N_30839);
nand U40955 (N_40955,N_31417,N_33951);
or U40956 (N_40956,N_30838,N_33197);
and U40957 (N_40957,N_38836,N_32691);
or U40958 (N_40958,N_34491,N_30863);
xnor U40959 (N_40959,N_35498,N_31235);
nand U40960 (N_40960,N_30320,N_33871);
or U40961 (N_40961,N_39968,N_35915);
or U40962 (N_40962,N_34095,N_33912);
and U40963 (N_40963,N_30398,N_35039);
nor U40964 (N_40964,N_34158,N_31289);
or U40965 (N_40965,N_37149,N_35534);
and U40966 (N_40966,N_33347,N_32770);
and U40967 (N_40967,N_38772,N_31204);
or U40968 (N_40968,N_38301,N_34326);
and U40969 (N_40969,N_36236,N_34439);
and U40970 (N_40970,N_31889,N_31772);
nand U40971 (N_40971,N_38699,N_36302);
and U40972 (N_40972,N_37572,N_33733);
nor U40973 (N_40973,N_36658,N_32114);
nand U40974 (N_40974,N_35527,N_34356);
or U40975 (N_40975,N_33080,N_31767);
xor U40976 (N_40976,N_37911,N_36300);
nand U40977 (N_40977,N_37919,N_36871);
nor U40978 (N_40978,N_32433,N_38990);
nor U40979 (N_40979,N_37555,N_33310);
xor U40980 (N_40980,N_30965,N_32959);
and U40981 (N_40981,N_34166,N_30674);
or U40982 (N_40982,N_34678,N_37817);
xor U40983 (N_40983,N_36464,N_33604);
xor U40984 (N_40984,N_33271,N_37562);
nor U40985 (N_40985,N_34066,N_38801);
nor U40986 (N_40986,N_36995,N_37820);
nand U40987 (N_40987,N_34687,N_38953);
and U40988 (N_40988,N_35525,N_36884);
xnor U40989 (N_40989,N_33574,N_38127);
and U40990 (N_40990,N_33363,N_30485);
or U40991 (N_40991,N_37021,N_38432);
and U40992 (N_40992,N_34258,N_32543);
or U40993 (N_40993,N_33732,N_38603);
nand U40994 (N_40994,N_37472,N_33452);
nor U40995 (N_40995,N_38734,N_38737);
nor U40996 (N_40996,N_30403,N_30171);
and U40997 (N_40997,N_31861,N_33978);
or U40998 (N_40998,N_36132,N_32258);
nand U40999 (N_40999,N_30540,N_33656);
and U41000 (N_41000,N_39797,N_32878);
and U41001 (N_41001,N_33838,N_37064);
nand U41002 (N_41002,N_38910,N_33088);
or U41003 (N_41003,N_35572,N_34667);
nand U41004 (N_41004,N_30392,N_35103);
or U41005 (N_41005,N_39798,N_32685);
nor U41006 (N_41006,N_37450,N_34555);
or U41007 (N_41007,N_38784,N_37309);
or U41008 (N_41008,N_35820,N_33787);
nor U41009 (N_41009,N_31623,N_38588);
and U41010 (N_41010,N_37690,N_37660);
nand U41011 (N_41011,N_38040,N_38170);
and U41012 (N_41012,N_33964,N_39740);
xor U41013 (N_41013,N_32067,N_33851);
nor U41014 (N_41014,N_30594,N_38175);
nor U41015 (N_41015,N_30861,N_31689);
and U41016 (N_41016,N_32007,N_32495);
nor U41017 (N_41017,N_33884,N_31152);
or U41018 (N_41018,N_38877,N_38868);
and U41019 (N_41019,N_36526,N_39586);
nor U41020 (N_41020,N_33819,N_36235);
or U41021 (N_41021,N_30128,N_33987);
nand U41022 (N_41022,N_36760,N_36222);
nor U41023 (N_41023,N_30939,N_35665);
nor U41024 (N_41024,N_37333,N_33158);
or U41025 (N_41025,N_37353,N_32790);
and U41026 (N_41026,N_31477,N_38047);
xor U41027 (N_41027,N_32075,N_35109);
nand U41028 (N_41028,N_38305,N_35879);
nand U41029 (N_41029,N_35465,N_38864);
or U41030 (N_41030,N_32070,N_35802);
nor U41031 (N_41031,N_34256,N_33932);
nor U41032 (N_41032,N_30331,N_39942);
and U41033 (N_41033,N_35151,N_30900);
nor U41034 (N_41034,N_30257,N_30655);
nand U41035 (N_41035,N_36056,N_37368);
and U41036 (N_41036,N_35114,N_38113);
nand U41037 (N_41037,N_35472,N_39218);
nor U41038 (N_41038,N_37354,N_35387);
or U41039 (N_41039,N_39157,N_34212);
nand U41040 (N_41040,N_33726,N_37769);
or U41041 (N_41041,N_33818,N_33037);
and U41042 (N_41042,N_36076,N_39260);
nand U41043 (N_41043,N_37076,N_32935);
xor U41044 (N_41044,N_38541,N_32746);
or U41045 (N_41045,N_31654,N_38447);
nor U41046 (N_41046,N_31906,N_37042);
nor U41047 (N_41047,N_34999,N_34368);
nor U41048 (N_41048,N_32552,N_39943);
nor U41049 (N_41049,N_38657,N_31073);
and U41050 (N_41050,N_34863,N_33830);
nor U41051 (N_41051,N_31560,N_34403);
nand U41052 (N_41052,N_34352,N_36449);
nor U41053 (N_41053,N_31842,N_37627);
and U41054 (N_41054,N_34465,N_33078);
and U41055 (N_41055,N_36175,N_32050);
and U41056 (N_41056,N_30899,N_31306);
nand U41057 (N_41057,N_33956,N_36587);
nor U41058 (N_41058,N_34187,N_39327);
and U41059 (N_41059,N_37511,N_38465);
nor U41060 (N_41060,N_37546,N_35726);
and U41061 (N_41061,N_31115,N_34155);
nor U41062 (N_41062,N_30500,N_37436);
nand U41063 (N_41063,N_38348,N_30681);
or U41064 (N_41064,N_31323,N_36241);
or U41065 (N_41065,N_35210,N_33396);
nor U41066 (N_41066,N_34252,N_38917);
nand U41067 (N_41067,N_38324,N_33768);
nor U41068 (N_41068,N_38533,N_30045);
nor U41069 (N_41069,N_33348,N_33123);
nor U41070 (N_41070,N_31335,N_30738);
nand U41071 (N_41071,N_31732,N_30639);
or U41072 (N_41072,N_37361,N_31658);
and U41073 (N_41073,N_33729,N_33868);
or U41074 (N_41074,N_30394,N_39337);
and U41075 (N_41075,N_38176,N_30072);
nand U41076 (N_41076,N_33058,N_34752);
nand U41077 (N_41077,N_30441,N_33180);
nor U41078 (N_41078,N_38512,N_34320);
nor U41079 (N_41079,N_31457,N_35344);
nand U41080 (N_41080,N_30678,N_36824);
xor U41081 (N_41081,N_38680,N_30960);
or U41082 (N_41082,N_32202,N_33174);
nand U41083 (N_41083,N_33061,N_38344);
nor U41084 (N_41084,N_30883,N_35561);
and U41085 (N_41085,N_37800,N_34370);
nand U41086 (N_41086,N_34637,N_37364);
nor U41087 (N_41087,N_33744,N_35688);
or U41088 (N_41088,N_31701,N_36431);
and U41089 (N_41089,N_37597,N_39655);
or U41090 (N_41090,N_34723,N_36873);
nand U41091 (N_41091,N_38407,N_34401);
nor U41092 (N_41092,N_39000,N_31721);
or U41093 (N_41093,N_39595,N_36379);
and U41094 (N_41094,N_33130,N_31138);
xor U41095 (N_41095,N_36797,N_32374);
and U41096 (N_41096,N_31387,N_32057);
or U41097 (N_41097,N_38177,N_34916);
and U41098 (N_41098,N_32760,N_30444);
or U41099 (N_41099,N_36484,N_34171);
xor U41100 (N_41100,N_32141,N_34162);
nand U41101 (N_41101,N_35132,N_35892);
nand U41102 (N_41102,N_31493,N_30766);
and U41103 (N_41103,N_34110,N_38217);
and U41104 (N_41104,N_35625,N_38712);
or U41105 (N_41105,N_32756,N_38765);
xnor U41106 (N_41106,N_37217,N_39585);
and U41107 (N_41107,N_36195,N_33468);
nor U41108 (N_41108,N_38937,N_39623);
xor U41109 (N_41109,N_35816,N_30693);
nor U41110 (N_41110,N_35933,N_32486);
or U41111 (N_41111,N_34090,N_39048);
nand U41112 (N_41112,N_30701,N_36080);
or U41113 (N_41113,N_39835,N_31363);
nand U41114 (N_41114,N_33228,N_37272);
nand U41115 (N_41115,N_34397,N_37666);
nor U41116 (N_41116,N_38627,N_36434);
nor U41117 (N_41117,N_39897,N_37659);
or U41118 (N_41118,N_34116,N_32557);
or U41119 (N_41119,N_32344,N_30997);
nand U41120 (N_41120,N_36959,N_36217);
and U41121 (N_41121,N_34508,N_38349);
or U41122 (N_41122,N_33943,N_30434);
and U41123 (N_41123,N_37262,N_39766);
nand U41124 (N_41124,N_33556,N_34600);
or U41125 (N_41125,N_33587,N_35366);
nor U41126 (N_41126,N_34755,N_36203);
or U41127 (N_41127,N_36154,N_32918);
nor U41128 (N_41128,N_30159,N_33531);
and U41129 (N_41129,N_33709,N_33576);
xor U41130 (N_41130,N_30109,N_36672);
nand U41131 (N_41131,N_34823,N_35801);
or U41132 (N_41132,N_34324,N_36815);
nor U41133 (N_41133,N_36040,N_32938);
nand U41134 (N_41134,N_32710,N_37052);
nand U41135 (N_41135,N_32192,N_35986);
nand U41136 (N_41136,N_30317,N_30907);
nand U41137 (N_41137,N_31813,N_32327);
and U41138 (N_41138,N_33670,N_30358);
nor U41139 (N_41139,N_39857,N_33765);
and U41140 (N_41140,N_33132,N_33534);
and U41141 (N_41141,N_34812,N_35250);
xor U41142 (N_41142,N_31866,N_30044);
and U41143 (N_41143,N_30829,N_33541);
or U41144 (N_41144,N_39104,N_36201);
nand U41145 (N_41145,N_37462,N_32597);
or U41146 (N_41146,N_30338,N_32473);
and U41147 (N_41147,N_32049,N_38523);
or U41148 (N_41148,N_31651,N_39969);
and U41149 (N_41149,N_30948,N_35091);
nand U41150 (N_41150,N_38667,N_35589);
xnor U41151 (N_41151,N_35708,N_34699);
nand U41152 (N_41152,N_39618,N_37346);
nand U41153 (N_41153,N_34388,N_37945);
and U41154 (N_41154,N_37460,N_34987);
xnor U41155 (N_41155,N_39966,N_30435);
and U41156 (N_41156,N_30335,N_34885);
nor U41157 (N_41157,N_32766,N_33758);
and U41158 (N_41158,N_37714,N_32994);
or U41159 (N_41159,N_31344,N_32531);
nand U41160 (N_41160,N_31042,N_33084);
or U41161 (N_41161,N_37704,N_31181);
or U41162 (N_41162,N_34275,N_30018);
nand U41163 (N_41163,N_30726,N_37266);
nor U41164 (N_41164,N_32018,N_35112);
or U41165 (N_41165,N_34551,N_39642);
nor U41166 (N_41166,N_38851,N_34872);
nor U41167 (N_41167,N_38089,N_38206);
and U41168 (N_41168,N_34763,N_34319);
xor U41169 (N_41169,N_34802,N_34775);
nand U41170 (N_41170,N_33009,N_39091);
nand U41171 (N_41171,N_32983,N_36897);
nand U41172 (N_41172,N_39637,N_33535);
or U41173 (N_41173,N_35604,N_30687);
and U41174 (N_41174,N_36896,N_34068);
or U41175 (N_41175,N_35441,N_37500);
xor U41176 (N_41176,N_31186,N_30020);
nor U41177 (N_41177,N_38957,N_39757);
and U41178 (N_41178,N_39065,N_36639);
nor U41179 (N_41179,N_30967,N_33710);
nor U41180 (N_41180,N_33704,N_33133);
xor U41181 (N_41181,N_33861,N_31400);
xor U41182 (N_41182,N_32357,N_30940);
xnor U41183 (N_41183,N_30735,N_37625);
xor U41184 (N_41184,N_39464,N_34759);
nor U41185 (N_41185,N_39315,N_36757);
or U41186 (N_41186,N_36833,N_33063);
nand U41187 (N_41187,N_38452,N_30309);
and U41188 (N_41188,N_32096,N_38250);
or U41189 (N_41189,N_38822,N_30881);
nand U41190 (N_41190,N_31700,N_33897);
and U41191 (N_41191,N_35733,N_35553);
or U41192 (N_41192,N_32979,N_33719);
or U41193 (N_41193,N_35715,N_33418);
or U41194 (N_41194,N_30117,N_35019);
nor U41195 (N_41195,N_30933,N_37470);
or U41196 (N_41196,N_39758,N_34560);
and U41197 (N_41197,N_36118,N_36106);
nor U41198 (N_41198,N_37344,N_32851);
nand U41199 (N_41199,N_35106,N_35319);
nor U41200 (N_41200,N_38569,N_35667);
xnor U41201 (N_41201,N_34259,N_36210);
nor U41202 (N_41202,N_30834,N_35052);
and U41203 (N_41203,N_35246,N_35381);
and U41204 (N_41204,N_32735,N_39278);
or U41205 (N_41205,N_39726,N_36017);
or U41206 (N_41206,N_36494,N_33183);
and U41207 (N_41207,N_33646,N_37160);
nand U41208 (N_41208,N_38703,N_36020);
or U41209 (N_41209,N_31908,N_30859);
xor U41210 (N_41210,N_35724,N_39719);
nand U41211 (N_41211,N_30321,N_31276);
and U41212 (N_41212,N_36361,N_32528);
or U41213 (N_41213,N_34713,N_31704);
nand U41214 (N_41214,N_36252,N_35307);
nor U41215 (N_41215,N_36248,N_35560);
or U41216 (N_41216,N_33998,N_30475);
nor U41217 (N_41217,N_38572,N_31285);
or U41218 (N_41218,N_35010,N_38360);
and U41219 (N_41219,N_33112,N_32941);
nor U41220 (N_41220,N_32913,N_31948);
or U41221 (N_41221,N_35316,N_35689);
nand U41222 (N_41222,N_37651,N_32016);
nand U41223 (N_41223,N_31434,N_30541);
nand U41224 (N_41224,N_35539,N_33825);
xor U41225 (N_41225,N_30852,N_33809);
or U41226 (N_41226,N_35753,N_39343);
nand U41227 (N_41227,N_32663,N_32414);
nor U41228 (N_41228,N_30785,N_39107);
nand U41229 (N_41229,N_30189,N_35111);
and U41230 (N_41230,N_38731,N_31274);
nand U41231 (N_41231,N_34507,N_33406);
xnor U41232 (N_41232,N_30365,N_31714);
nor U41233 (N_41233,N_30420,N_35937);
nand U41234 (N_41234,N_38984,N_34337);
or U41235 (N_41235,N_34089,N_30162);
xor U41236 (N_41236,N_30873,N_39007);
and U41237 (N_41237,N_32410,N_30102);
and U41238 (N_41238,N_32026,N_34035);
xnor U41239 (N_41239,N_36303,N_34453);
nor U41240 (N_41240,N_31979,N_39014);
or U41241 (N_41241,N_37387,N_32525);
or U41242 (N_41242,N_31662,N_38773);
nor U41243 (N_41243,N_31672,N_36250);
nor U41244 (N_41244,N_35230,N_38815);
and U41245 (N_41245,N_33403,N_39496);
xnor U41246 (N_41246,N_36868,N_33421);
or U41247 (N_41247,N_33555,N_38253);
nor U41248 (N_41248,N_30569,N_32762);
nor U41249 (N_41249,N_34696,N_37476);
and U41250 (N_41250,N_36958,N_36717);
nand U41251 (N_41251,N_33748,N_37925);
nor U41252 (N_41252,N_32054,N_35651);
or U41253 (N_41253,N_31214,N_33946);
nand U41254 (N_41254,N_39124,N_36939);
and U41255 (N_41255,N_36809,N_31615);
nand U41256 (N_41256,N_31660,N_38976);
nor U41257 (N_41257,N_35288,N_31165);
or U41258 (N_41258,N_32471,N_39918);
nand U41259 (N_41259,N_31290,N_38193);
xor U41260 (N_41260,N_30848,N_36188);
and U41261 (N_41261,N_38727,N_37972);
xor U41262 (N_41262,N_39649,N_31641);
and U41263 (N_41263,N_39112,N_31462);
nor U41264 (N_41264,N_37793,N_37822);
nand U41265 (N_41265,N_35335,N_30487);
or U41266 (N_41266,N_31302,N_34529);
or U41267 (N_41267,N_39090,N_30588);
nand U41268 (N_41268,N_38783,N_34544);
nor U41269 (N_41269,N_32396,N_33297);
nand U41270 (N_41270,N_39473,N_31286);
xnor U41271 (N_41271,N_32992,N_38514);
nand U41272 (N_41272,N_34907,N_35963);
xnor U41273 (N_41273,N_38549,N_35752);
or U41274 (N_41274,N_36281,N_34745);
or U41275 (N_41275,N_35608,N_30446);
and U41276 (N_41276,N_34673,N_32191);
or U41277 (N_41277,N_37245,N_33784);
and U41278 (N_41278,N_36044,N_31268);
or U41279 (N_41279,N_38124,N_35814);
xnor U41280 (N_41280,N_35294,N_34222);
or U41281 (N_41281,N_35482,N_34107);
nand U41282 (N_41282,N_33590,N_31162);
and U41283 (N_41283,N_32280,N_30986);
or U41284 (N_41284,N_30362,N_38591);
or U41285 (N_41285,N_33796,N_32446);
nand U41286 (N_41286,N_30353,N_31771);
nor U41287 (N_41287,N_35187,N_33027);
and U41288 (N_41288,N_34455,N_32438);
xor U41289 (N_41289,N_33947,N_34893);
nand U41290 (N_41290,N_37569,N_31712);
nor U41291 (N_41291,N_32481,N_30244);
nand U41292 (N_41292,N_31267,N_31096);
nor U41293 (N_41293,N_31874,N_35702);
and U41294 (N_41294,N_36277,N_36974);
nor U41295 (N_41295,N_39659,N_30998);
nor U41296 (N_41296,N_33821,N_36353);
nand U41297 (N_41297,N_34145,N_32632);
and U41298 (N_41298,N_33589,N_34769);
nand U41299 (N_41299,N_36364,N_30656);
or U41300 (N_41300,N_36113,N_38322);
nor U41301 (N_41301,N_31669,N_33060);
or U41302 (N_41302,N_30451,N_37957);
or U41303 (N_41303,N_38598,N_35119);
nand U41304 (N_41304,N_35224,N_36380);
nor U41305 (N_41305,N_39858,N_37676);
nor U41306 (N_41306,N_35275,N_32063);
or U41307 (N_41307,N_35050,N_38706);
nor U41308 (N_41308,N_37278,N_36511);
or U41309 (N_41309,N_35306,N_34549);
xnor U41310 (N_41310,N_31707,N_30250);
and U41311 (N_41311,N_39196,N_32348);
or U41312 (N_41312,N_34534,N_36042);
or U41313 (N_41313,N_38916,N_32902);
and U41314 (N_41314,N_31529,N_31737);
nor U41315 (N_41315,N_30522,N_31955);
and U41316 (N_41316,N_35068,N_37766);
nand U41317 (N_41317,N_30854,N_37260);
or U41318 (N_41318,N_33817,N_39520);
nor U41319 (N_41319,N_39368,N_36539);
nor U41320 (N_41320,N_39780,N_35696);
and U41321 (N_41321,N_32817,N_35480);
nand U41322 (N_41322,N_37811,N_34100);
nand U41323 (N_41323,N_33455,N_36428);
nor U41324 (N_41324,N_38296,N_37351);
or U41325 (N_41325,N_39840,N_39547);
or U41326 (N_41326,N_32332,N_31001);
or U41327 (N_41327,N_33989,N_37675);
nand U41328 (N_41328,N_36068,N_37389);
and U41329 (N_41329,N_37812,N_34152);
nor U41330 (N_41330,N_39207,N_35989);
nand U41331 (N_41331,N_38495,N_31247);
or U41332 (N_41332,N_32353,N_32491);
nor U41333 (N_41333,N_31288,N_37069);
or U41334 (N_41334,N_30455,N_38275);
nand U41335 (N_41335,N_30316,N_36163);
and U41336 (N_41336,N_38424,N_38025);
or U41337 (N_41337,N_36376,N_30110);
nor U41338 (N_41338,N_37913,N_33393);
and U41339 (N_41339,N_32566,N_38436);
and U41340 (N_41340,N_36590,N_31680);
and U41341 (N_41341,N_33318,N_36579);
or U41342 (N_41342,N_32949,N_37072);
and U41343 (N_41343,N_35283,N_36182);
nand U41344 (N_41344,N_36903,N_36713);
nand U41345 (N_41345,N_39718,N_34031);
or U41346 (N_41346,N_36429,N_38419);
nor U41347 (N_41347,N_33195,N_32551);
or U41348 (N_41348,N_31264,N_34639);
nand U41349 (N_41349,N_37463,N_30468);
nor U41350 (N_41350,N_32550,N_32217);
or U41351 (N_41351,N_36543,N_31506);
or U41352 (N_41352,N_33025,N_35244);
xnor U41353 (N_41353,N_35556,N_38863);
and U41354 (N_41354,N_39202,N_31815);
and U41355 (N_41355,N_33002,N_38071);
and U41356 (N_41356,N_33135,N_39987);
and U41357 (N_41357,N_33944,N_34026);
and U41358 (N_41358,N_30532,N_32140);
nor U41359 (N_41359,N_34414,N_33986);
nor U41360 (N_41360,N_37828,N_32498);
nand U41361 (N_41361,N_33570,N_35400);
and U41362 (N_41362,N_33395,N_35323);
nand U41363 (N_41363,N_33311,N_39199);
xor U41364 (N_41364,N_35305,N_35488);
and U41365 (N_41365,N_37789,N_30369);
and U41366 (N_41366,N_39703,N_39593);
or U41367 (N_41367,N_30627,N_35838);
nand U41368 (N_41368,N_30700,N_38637);
or U41369 (N_41369,N_31942,N_34299);
xor U41370 (N_41370,N_38310,N_39822);
nand U41371 (N_41371,N_33546,N_36694);
nand U41372 (N_41372,N_38174,N_30523);
nor U41373 (N_41373,N_33414,N_35357);
nand U41374 (N_41374,N_34334,N_35832);
and U41375 (N_41375,N_38889,N_37850);
or U41376 (N_41376,N_31384,N_30265);
and U41377 (N_41377,N_34056,N_32346);
and U41378 (N_41378,N_38321,N_34559);
xor U41379 (N_41379,N_30164,N_39596);
and U41380 (N_41380,N_35059,N_31322);
nor U41381 (N_41381,N_30417,N_35193);
nand U41382 (N_41382,N_38233,N_36440);
or U41383 (N_41383,N_32984,N_36981);
nand U41384 (N_41384,N_36846,N_33272);
xnor U41385 (N_41385,N_35201,N_36671);
and U41386 (N_41386,N_31859,N_32505);
and U41387 (N_41387,N_37985,N_32345);
nand U41388 (N_41388,N_32504,N_30346);
or U41389 (N_41389,N_35587,N_32815);
or U41390 (N_41390,N_39242,N_32754);
nand U41391 (N_41391,N_36545,N_30495);
or U41392 (N_41392,N_35807,N_31638);
or U41393 (N_41393,N_35717,N_31099);
nand U41394 (N_41394,N_31722,N_36806);
or U41395 (N_41395,N_39747,N_31206);
and U41396 (N_41396,N_34784,N_31154);
nand U41397 (N_41397,N_37602,N_31159);
and U41398 (N_41398,N_38689,N_34888);
nand U41399 (N_41399,N_31830,N_30381);
xnor U41400 (N_41400,N_39543,N_31963);
nand U41401 (N_41401,N_37301,N_32750);
nand U41402 (N_41402,N_38500,N_34694);
or U41403 (N_41403,N_38580,N_32110);
nor U41404 (N_41404,N_36697,N_36554);
and U41405 (N_41405,N_32635,N_31389);
nor U41406 (N_41406,N_35416,N_30195);
or U41407 (N_41407,N_38798,N_30558);
and U41408 (N_41408,N_30151,N_31396);
or U41409 (N_41409,N_30133,N_38862);
nor U41410 (N_41410,N_30484,N_32285);
nor U41411 (N_41411,N_39711,N_32673);
nor U41412 (N_41412,N_32909,N_38340);
nand U41413 (N_41413,N_36437,N_36929);
and U41414 (N_41414,N_35813,N_30094);
and U41415 (N_41415,N_34515,N_35827);
nand U41416 (N_41416,N_35855,N_31251);
nand U41417 (N_41417,N_35515,N_33549);
and U41418 (N_41418,N_39574,N_37488);
and U41419 (N_41419,N_37951,N_35658);
or U41420 (N_41420,N_36948,N_39570);
and U41421 (N_41421,N_36874,N_37380);
nand U41422 (N_41422,N_33984,N_39086);
xnor U41423 (N_41423,N_30534,N_38121);
or U41424 (N_41424,N_33761,N_33449);
and U41425 (N_41425,N_36926,N_38739);
nor U41426 (N_41426,N_38899,N_34890);
nand U41427 (N_41427,N_33293,N_35890);
nor U41428 (N_41428,N_32861,N_38128);
xnor U41429 (N_41429,N_36937,N_37554);
xnor U41430 (N_41430,N_32535,N_37702);
and U41431 (N_41431,N_33108,N_34700);
nor U41432 (N_41432,N_37545,N_38437);
nor U41433 (N_41433,N_32153,N_38466);
and U41434 (N_41434,N_35189,N_35532);
xor U41435 (N_41435,N_35258,N_33752);
or U41436 (N_41436,N_39561,N_38048);
nor U41437 (N_41437,N_32439,N_39777);
nand U41438 (N_41438,N_39229,N_34587);
and U41439 (N_41439,N_30754,N_37901);
nor U41440 (N_41440,N_36487,N_33929);
and U41441 (N_41441,N_31903,N_31185);
and U41442 (N_41442,N_34826,N_37862);
xor U41443 (N_41443,N_37875,N_37873);
nor U41444 (N_41444,N_33482,N_38853);
or U41445 (N_41445,N_34072,N_31189);
and U41446 (N_41446,N_32082,N_36552);
nand U41447 (N_41447,N_39743,N_34880);
or U41448 (N_41448,N_34553,N_37764);
nor U41449 (N_41449,N_39764,N_39198);
or U41450 (N_41450,N_37890,N_37638);
nor U41451 (N_41451,N_35227,N_30802);
xor U41452 (N_41452,N_39188,N_31989);
nand U41453 (N_41453,N_34783,N_36133);
nand U41454 (N_41454,N_39511,N_30075);
nand U41455 (N_41455,N_31548,N_38909);
and U41456 (N_41456,N_38062,N_36614);
nand U41457 (N_41457,N_30796,N_36048);
or U41458 (N_41458,N_33003,N_32181);
xor U41459 (N_41459,N_35391,N_32613);
and U41460 (N_41460,N_34197,N_36681);
and U41461 (N_41461,N_35728,N_36384);
nand U41462 (N_41462,N_33795,N_35596);
nor U41463 (N_41463,N_39701,N_34841);
nand U41464 (N_41464,N_33221,N_30853);
xor U41465 (N_41465,N_38527,N_30969);
nor U41466 (N_41466,N_33759,N_38030);
and U41467 (N_41467,N_31157,N_38492);
xnor U41468 (N_41468,N_30126,N_30572);
nor U41469 (N_41469,N_34886,N_35372);
xor U41470 (N_41470,N_37435,N_34424);
nand U41471 (N_41471,N_34061,N_37070);
or U41472 (N_41472,N_30717,N_38623);
and U41473 (N_41473,N_35170,N_37810);
xnor U41474 (N_41474,N_33444,N_39130);
nor U41475 (N_41475,N_36502,N_32317);
or U41476 (N_41476,N_34847,N_38397);
and U41477 (N_41477,N_39508,N_30101);
or U41478 (N_41478,N_32680,N_38515);
or U41479 (N_41479,N_30778,N_31800);
xor U41480 (N_41480,N_37474,N_31649);
and U41481 (N_41481,N_34183,N_35251);
xor U41482 (N_41482,N_38978,N_34554);
or U41483 (N_41483,N_39017,N_36901);
nand U41484 (N_41484,N_37015,N_39363);
or U41485 (N_41485,N_35449,N_39306);
and U41486 (N_41486,N_33714,N_36978);
nor U41487 (N_41487,N_34119,N_33054);
or U41488 (N_41488,N_37838,N_39679);
or U41489 (N_41489,N_35842,N_39619);
or U41490 (N_41490,N_33909,N_38744);
and U41491 (N_41491,N_35130,N_33269);
and U41492 (N_41492,N_35098,N_37983);
nor U41493 (N_41493,N_34284,N_34170);
nand U41494 (N_41494,N_30508,N_38799);
nor U41495 (N_41495,N_37518,N_30669);
nor U41496 (N_41496,N_34316,N_38184);
or U41497 (N_41497,N_34977,N_34157);
nand U41498 (N_41498,N_39578,N_30367);
or U41499 (N_41499,N_37390,N_33026);
or U41500 (N_41500,N_39565,N_30545);
nand U41501 (N_41501,N_30428,N_30524);
and U41502 (N_41502,N_31616,N_32238);
and U41503 (N_41503,N_32584,N_34346);
or U41504 (N_41504,N_35679,N_30507);
or U41505 (N_41505,N_35166,N_38220);
xor U41506 (N_41506,N_33402,N_34995);
nor U41507 (N_41507,N_30734,N_35077);
xnor U41508 (N_41508,N_39016,N_32642);
and U41509 (N_41509,N_35943,N_37537);
nor U41510 (N_41510,N_36157,N_31601);
or U41511 (N_41511,N_31570,N_30583);
and U41512 (N_41512,N_35265,N_32235);
and U41513 (N_41513,N_35848,N_38037);
nand U41514 (N_41514,N_31740,N_32540);
xnor U41515 (N_41515,N_30552,N_31612);
nor U41516 (N_41516,N_33614,N_35544);
and U41517 (N_41517,N_30832,N_30271);
nor U41518 (N_41518,N_36325,N_35590);
nand U41519 (N_41519,N_38770,N_33356);
or U41520 (N_41520,N_31272,N_35575);
and U41521 (N_41521,N_37490,N_38139);
and U41522 (N_41522,N_32206,N_31897);
nand U41523 (N_41523,N_37837,N_39173);
and U41524 (N_41524,N_32072,N_36755);
or U41525 (N_41525,N_32812,N_32448);
nor U41526 (N_41526,N_35018,N_37842);
and U41527 (N_41527,N_36957,N_32175);
or U41528 (N_41528,N_31245,N_39622);
or U41529 (N_41529,N_39996,N_35364);
nor U41530 (N_41530,N_39678,N_33626);
and U41531 (N_41531,N_32854,N_39670);
nand U41532 (N_41532,N_37641,N_34706);
or U41533 (N_41533,N_33176,N_38290);
nand U41534 (N_41534,N_30058,N_37152);
nor U41535 (N_41535,N_31916,N_36783);
or U41536 (N_41536,N_32826,N_35719);
or U41537 (N_41537,N_39147,N_30716);
or U41538 (N_41538,N_30155,N_34406);
or U41539 (N_41539,N_39549,N_31370);
and U41540 (N_41540,N_38357,N_37171);
or U41541 (N_41541,N_33494,N_33945);
and U41542 (N_41542,N_32306,N_37293);
and U41543 (N_41543,N_32594,N_36388);
nor U41544 (N_41544,N_35592,N_34106);
or U41545 (N_41545,N_38719,N_39790);
or U41546 (N_41546,N_31655,N_37847);
nor U41547 (N_41547,N_39852,N_37606);
and U41548 (N_41548,N_33677,N_30186);
or U41549 (N_41549,N_33618,N_31341);
nand U41550 (N_41550,N_32502,N_31303);
nand U41551 (N_41551,N_38477,N_37065);
and U41552 (N_41552,N_30906,N_35798);
or U41553 (N_41553,N_30290,N_36923);
or U41554 (N_41554,N_35932,N_33777);
nand U41555 (N_41555,N_36814,N_34574);
nor U41556 (N_41556,N_37670,N_32516);
nor U41557 (N_41557,N_36518,N_35536);
and U41558 (N_41558,N_33793,N_38491);
and U41559 (N_41559,N_34133,N_39297);
nor U41560 (N_41560,N_31244,N_31442);
and U41561 (N_41561,N_33260,N_35998);
or U41562 (N_41562,N_31190,N_36489);
nor U41563 (N_41563,N_39209,N_35875);
xnor U41564 (N_41564,N_35235,N_37033);
or U41565 (N_41565,N_35140,N_35141);
nand U41566 (N_41566,N_31682,N_35977);
nor U41567 (N_41567,N_39809,N_31342);
nor U41568 (N_41568,N_30956,N_35803);
or U41569 (N_41569,N_39573,N_32105);
and U41570 (N_41570,N_34201,N_33301);
or U41571 (N_41571,N_33192,N_32842);
nand U41572 (N_41572,N_37691,N_38429);
or U41573 (N_41573,N_35389,N_39039);
and U41574 (N_41574,N_35521,N_32734);
nor U41575 (N_41575,N_35558,N_33550);
or U41576 (N_41576,N_37440,N_36033);
nand U41577 (N_41577,N_32553,N_32835);
or U41578 (N_41578,N_37960,N_39318);
xor U41579 (N_41579,N_39795,N_33867);
and U41580 (N_41580,N_37866,N_38044);
and U41581 (N_41581,N_36839,N_32121);
nor U41582 (N_41582,N_32943,N_36677);
nor U41583 (N_41583,N_38126,N_33141);
nor U41584 (N_41584,N_36146,N_37434);
xor U41585 (N_41585,N_35253,N_32549);
nand U41586 (N_41586,N_34680,N_39834);
nand U41587 (N_41587,N_35385,N_31317);
nand U41588 (N_41588,N_30502,N_37726);
nor U41589 (N_41589,N_36795,N_37844);
nor U41590 (N_41590,N_39952,N_36213);
xnor U41591 (N_41591,N_30239,N_37867);
xor U41592 (N_41592,N_33595,N_38298);
xnor U41593 (N_41593,N_36546,N_38185);
or U41594 (N_41594,N_36422,N_31852);
nor U41595 (N_41595,N_39185,N_36811);
nor U41596 (N_41596,N_36829,N_37729);
and U41597 (N_41597,N_38198,N_30982);
nor U41598 (N_41598,N_35704,N_32946);
or U41599 (N_41599,N_35634,N_36525);
and U41600 (N_41600,N_34180,N_31439);
nor U41601 (N_41601,N_34602,N_30843);
nand U41602 (N_41602,N_32782,N_38095);
or U41603 (N_41603,N_35939,N_34377);
xnor U41604 (N_41604,N_34840,N_33210);
or U41605 (N_41605,N_33430,N_30844);
nor U41606 (N_41606,N_34382,N_35255);
or U41607 (N_41607,N_38167,N_30082);
and U41608 (N_41608,N_39909,N_31333);
nand U41609 (N_41609,N_38927,N_30535);
nor U41610 (N_41610,N_34985,N_33168);
or U41611 (N_41611,N_30791,N_31536);
and U41612 (N_41612,N_38846,N_37172);
or U41613 (N_41613,N_32522,N_30714);
xnor U41614 (N_41614,N_35538,N_30847);
nand U41615 (N_41615,N_38103,N_31887);
and U41616 (N_41616,N_33564,N_30554);
and U41617 (N_41617,N_36964,N_32449);
nand U41618 (N_41618,N_39393,N_30040);
and U41619 (N_41619,N_38914,N_34207);
or U41620 (N_41620,N_31835,N_30457);
or U41621 (N_41621,N_33309,N_35439);
nor U41622 (N_41622,N_32554,N_30450);
nand U41623 (N_41623,N_36727,N_30370);
and U41624 (N_41624,N_38014,N_38852);
nor U41625 (N_41625,N_30356,N_30571);
and U41626 (N_41626,N_30962,N_39579);
xor U41627 (N_41627,N_30211,N_35914);
nand U41628 (N_41628,N_32164,N_38462);
xor U41629 (N_41629,N_30915,N_34028);
nor U41630 (N_41630,N_37084,N_37236);
nand U41631 (N_41631,N_36767,N_32239);
and U41632 (N_41632,N_30640,N_36813);
nand U41633 (N_41633,N_32887,N_31210);
nor U41634 (N_41634,N_36703,N_34676);
nor U41635 (N_41635,N_31832,N_37311);
nor U41636 (N_41636,N_33162,N_36994);
nand U41637 (N_41637,N_32441,N_32605);
and U41638 (N_41638,N_38558,N_35992);
nor U41639 (N_41639,N_38695,N_31173);
or U41640 (N_41640,N_30768,N_37950);
nor U41641 (N_41641,N_30419,N_35428);
and U41642 (N_41642,N_30258,N_35823);
and U41643 (N_41643,N_33305,N_32086);
xor U41644 (N_41644,N_34022,N_34174);
nand U41645 (N_41645,N_38009,N_38517);
nand U41646 (N_41646,N_39079,N_37815);
and U41647 (N_41647,N_37499,N_38566);
and U41648 (N_41648,N_36731,N_31555);
or U41649 (N_41649,N_31741,N_37824);
or U41650 (N_41650,N_37656,N_33621);
or U41651 (N_41651,N_35447,N_35758);
nor U41652 (N_41652,N_37271,N_34785);
nor U41653 (N_41653,N_34374,N_38816);
nand U41654 (N_41654,N_35524,N_32017);
and U41655 (N_41655,N_35318,N_37176);
nor U41656 (N_41656,N_38755,N_36941);
and U41657 (N_41657,N_33300,N_31398);
nand U41658 (N_41658,N_31855,N_38254);
or U41659 (N_41659,N_39213,N_37505);
and U41660 (N_41660,N_30043,N_34271);
nand U41661 (N_41661,N_37861,N_35163);
and U41662 (N_41662,N_33993,N_39342);
xor U41663 (N_41663,N_33948,N_36707);
nand U41664 (N_41664,N_35092,N_37962);
nor U41665 (N_41665,N_38893,N_33957);
nor U41666 (N_41666,N_34921,N_38413);
nor U41667 (N_41667,N_34122,N_33772);
nor U41668 (N_41668,N_34634,N_36226);
xnor U41669 (N_41669,N_34218,N_33086);
nor U41670 (N_41670,N_31664,N_33425);
or U41671 (N_41671,N_31837,N_33222);
and U41672 (N_41672,N_33865,N_30299);
or U41673 (N_41673,N_39291,N_34934);
and U41674 (N_41674,N_34444,N_38010);
or U41675 (N_41675,N_32840,N_30644);
nand U41676 (N_41676,N_34265,N_37277);
and U41677 (N_41677,N_31229,N_35513);
or U41678 (N_41678,N_37469,N_34867);
nor U41679 (N_41679,N_30548,N_39273);
nor U41680 (N_41680,N_36097,N_38192);
nor U41681 (N_41681,N_34495,N_32538);
nor U41682 (N_41682,N_38668,N_33580);
nand U41683 (N_41683,N_32178,N_30919);
nand U41684 (N_41684,N_33015,N_33182);
or U41685 (N_41685,N_36913,N_35042);
and U41686 (N_41686,N_36095,N_36496);
nand U41687 (N_41687,N_31060,N_34154);
nand U41688 (N_41688,N_36904,N_31710);
or U41689 (N_41689,N_36089,N_34787);
and U41690 (N_41690,N_37772,N_37886);
nand U41691 (N_41691,N_32165,N_38417);
xor U41692 (N_41692,N_37975,N_33106);
or U41693 (N_41693,N_33836,N_30347);
or U41694 (N_41694,N_36626,N_35256);
nor U41695 (N_41695,N_38480,N_36046);
nand U41696 (N_41696,N_35833,N_39776);
nand U41697 (N_41697,N_31975,N_33770);
nand U41698 (N_41698,N_31062,N_34950);
xnor U41699 (N_41699,N_32160,N_37863);
or U41700 (N_41700,N_34716,N_32720);
or U41701 (N_41701,N_38023,N_39556);
nor U41702 (N_41702,N_39505,N_38214);
xor U41703 (N_41703,N_38585,N_38561);
or U41704 (N_41704,N_38605,N_31999);
or U41705 (N_41705,N_31590,N_39825);
nor U41706 (N_41706,N_35808,N_37370);
or U41707 (N_41707,N_35376,N_39625);
nor U41708 (N_41708,N_32585,N_32574);
nand U41709 (N_41709,N_31543,N_38979);
or U41710 (N_41710,N_37032,N_36542);
nand U41711 (N_41711,N_36500,N_36588);
or U41712 (N_41712,N_36274,N_38196);
or U41713 (N_41713,N_34492,N_34836);
or U41714 (N_41714,N_39638,N_36753);
and U41715 (N_41715,N_39285,N_33567);
nor U41716 (N_41716,N_37697,N_35423);
and U41717 (N_41717,N_39081,N_36270);
and U41718 (N_41718,N_39627,N_38156);
nor U41719 (N_41719,N_30601,N_38666);
nor U41720 (N_41720,N_30557,N_32989);
nand U41721 (N_41721,N_30641,N_39944);
and U41722 (N_41722,N_35215,N_33887);
nor U41723 (N_41723,N_37136,N_35896);
and U41724 (N_41724,N_36413,N_39830);
nor U41725 (N_41725,N_34850,N_39402);
nor U41726 (N_41726,N_35687,N_32429);
nand U41727 (N_41727,N_32379,N_32231);
nand U41728 (N_41728,N_33607,N_31802);
nand U41729 (N_41729,N_38342,N_34523);
nor U41730 (N_41730,N_36657,N_39261);
nand U41731 (N_41731,N_38857,N_30216);
and U41732 (N_41732,N_39850,N_30084);
nand U41733 (N_41733,N_34721,N_34747);
nand U41734 (N_41734,N_35070,N_34178);
nand U41735 (N_41735,N_30657,N_36025);
and U41736 (N_41736,N_33409,N_35402);
or U41737 (N_41737,N_33721,N_36679);
and U41738 (N_41738,N_33273,N_39608);
nor U41739 (N_41739,N_33433,N_38785);
nand U41740 (N_41740,N_35159,N_32666);
nand U41741 (N_41741,N_30543,N_35616);
or U41742 (N_41742,N_31016,N_36820);
and U41743 (N_41743,N_30570,N_30966);
nor U41744 (N_41744,N_34143,N_38814);
nor U41745 (N_41745,N_38760,N_30097);
and U41746 (N_41746,N_31107,N_37914);
or U41747 (N_41747,N_31130,N_36791);
or U41748 (N_41748,N_39564,N_31312);
and U41749 (N_41749,N_34457,N_34793);
and U41750 (N_41750,N_32797,N_34868);
nor U41751 (N_41751,N_32886,N_30628);
or U41752 (N_41752,N_36104,N_38829);
and U41753 (N_41753,N_30994,N_30233);
and U41754 (N_41754,N_36916,N_37352);
or U41755 (N_41755,N_39475,N_31883);
and U41756 (N_41756,N_36381,N_37117);
xor U41757 (N_41757,N_36748,N_39468);
nor U41758 (N_41758,N_35858,N_32496);
and U41759 (N_41759,N_34472,N_36150);
nand U41760 (N_41760,N_39817,N_31056);
or U41761 (N_41761,N_34434,N_35102);
nor U41762 (N_41762,N_37527,N_32923);
nor U41763 (N_41763,N_39184,N_30961);
and U41764 (N_41764,N_32542,N_38581);
xnor U41765 (N_41765,N_38248,N_35620);
nand U41766 (N_41766,N_31794,N_33428);
and U41767 (N_41767,N_32699,N_34824);
or U41768 (N_41768,N_32289,N_31709);
nand U41769 (N_41769,N_31598,N_31430);
and U41770 (N_41770,N_30875,N_39641);
xnor U41771 (N_41771,N_32037,N_38963);
xor U41772 (N_41772,N_37191,N_38550);
and U41773 (N_41773,N_34169,N_36779);
and U41774 (N_41774,N_31735,N_37514);
or U41775 (N_41775,N_36408,N_34047);
or U41776 (N_41776,N_34317,N_33104);
or U41777 (N_41777,N_37616,N_39753);
xor U41778 (N_41778,N_38743,N_33175);
nor U41779 (N_41779,N_38692,N_37495);
and U41780 (N_41780,N_34013,N_37544);
xor U41781 (N_41781,N_39239,N_30732);
nor U41782 (N_41782,N_35346,N_39654);
nand U41783 (N_41783,N_38187,N_31123);
and U41784 (N_41784,N_38483,N_31822);
nand U41785 (N_41785,N_39864,N_34849);
nor U41786 (N_41786,N_38981,N_33568);
and U41787 (N_41787,N_35686,N_36461);
nand U41788 (N_41788,N_37588,N_32649);
or U41789 (N_41789,N_30348,N_37464);
and U41790 (N_41790,N_33148,N_37698);
nor U41791 (N_41791,N_33906,N_31461);
and U41792 (N_41792,N_37384,N_39289);
nor U41793 (N_41793,N_34483,N_32343);
nand U41794 (N_41794,N_37321,N_33359);
or U41795 (N_41795,N_37051,N_35226);
or U41796 (N_41796,N_36609,N_38320);
xnor U41797 (N_41797,N_36514,N_30074);
or U41798 (N_41798,N_30774,N_31792);
nand U41799 (N_41799,N_35186,N_34511);
and U41800 (N_41800,N_31166,N_33921);
nand U41801 (N_41801,N_37929,N_30636);
and U41802 (N_41802,N_30340,N_33072);
and U41803 (N_41803,N_34064,N_39280);
nand U41804 (N_41804,N_36352,N_35029);
or U41805 (N_41805,N_36950,N_38675);
xor U41806 (N_41806,N_35174,N_39335);
nand U41807 (N_41807,N_39774,N_31049);
nor U41808 (N_41808,N_36699,N_35598);
nand U41809 (N_41809,N_32820,N_35691);
or U41810 (N_41810,N_34462,N_31271);
nor U41811 (N_41811,N_38503,N_38827);
xor U41812 (N_41812,N_30826,N_38024);
and U41813 (N_41813,N_39258,N_32526);
and U41814 (N_41814,N_36045,N_34976);
xnor U41815 (N_41815,N_35403,N_30319);
or U41816 (N_41816,N_34425,N_30130);
nand U41817 (N_41817,N_34679,N_37501);
and U41818 (N_41818,N_32650,N_36524);
nor U41819 (N_41819,N_31868,N_36467);
and U41820 (N_41820,N_30607,N_38716);
xnor U41821 (N_41821,N_33609,N_35681);
and U41822 (N_41822,N_34209,N_38352);
or U41823 (N_41823,N_32603,N_36857);
nand U41824 (N_41824,N_39487,N_32008);
nand U41825 (N_41825,N_39389,N_32534);
and U41826 (N_41826,N_34683,N_35212);
and U41827 (N_41827,N_30943,N_31613);
nand U41828 (N_41828,N_35888,N_33572);
nor U41829 (N_41829,N_32180,N_32694);
xnor U41830 (N_41830,N_35422,N_36673);
and U41831 (N_41831,N_34926,N_33493);
xor U41832 (N_41832,N_31545,N_35333);
nand U41833 (N_41833,N_39838,N_37516);
or U41834 (N_41834,N_30283,N_37760);
nor U41835 (N_41835,N_37794,N_38808);
nor U41836 (N_41836,N_37267,N_39803);
nor U41837 (N_41837,N_38511,N_32541);
or U41838 (N_41838,N_35911,N_37060);
and U41839 (N_41839,N_36885,N_34186);
nand U41840 (N_41840,N_33181,N_30989);
nand U41841 (N_41841,N_35436,N_38493);
or U41842 (N_41842,N_37497,N_34126);
or U41843 (N_41843,N_35363,N_38001);
or U41844 (N_41844,N_34177,N_35392);
nor U41845 (N_41845,N_32647,N_35195);
and U41846 (N_41846,N_39778,N_31205);
nand U41847 (N_41847,N_30205,N_38097);
and U41848 (N_41848,N_38488,N_37980);
or U41849 (N_41849,N_35947,N_32701);
or U41850 (N_41850,N_30049,N_37421);
or U41851 (N_41851,N_31878,N_38662);
nand U41852 (N_41852,N_30046,N_35216);
nand U41853 (N_41853,N_30124,N_38087);
nand U41854 (N_41854,N_31851,N_30464);
nand U41855 (N_41855,N_34837,N_38200);
nand U41856 (N_41856,N_31087,N_39831);
or U41857 (N_41857,N_31379,N_30673);
and U41858 (N_41858,N_33515,N_34947);
or U41859 (N_41859,N_36773,N_35805);
nand U41860 (N_41860,N_35236,N_34827);
nor U41861 (N_41861,N_34603,N_31125);
or U41862 (N_41862,N_35142,N_37596);
nor U41863 (N_41863,N_39158,N_31780);
nand U41864 (N_41864,N_36736,N_32035);
and U41865 (N_41865,N_32197,N_38831);
nor U41866 (N_41866,N_35676,N_30750);
nand U41867 (N_41867,N_38390,N_33655);
or U41868 (N_41868,N_39611,N_31857);
or U41869 (N_41869,N_36705,N_32775);
or U41870 (N_41870,N_31117,N_34030);
or U41871 (N_41871,N_34852,N_31422);
or U41872 (N_41872,N_39981,N_33256);
nand U41873 (N_41873,N_31470,N_34139);
and U41874 (N_41874,N_33053,N_32118);
xor U41875 (N_41875,N_31718,N_36403);
and U41876 (N_41876,N_39418,N_34065);
xor U41877 (N_41877,N_36597,N_34198);
and U41878 (N_41878,N_37414,N_30368);
and U41879 (N_41879,N_33239,N_31763);
and U41880 (N_41880,N_39372,N_35468);
and U41881 (N_41881,N_38371,N_30896);
nor U41882 (N_41882,N_39628,N_30537);
nor U41883 (N_41883,N_32331,N_37022);
nor U41884 (N_41884,N_32356,N_35783);
nand U41885 (N_41885,N_35999,N_30567);
nand U41886 (N_41886,N_37563,N_37574);
nand U41887 (N_41887,N_33279,N_39844);
nand U41888 (N_41888,N_37855,N_34225);
and U41889 (N_41889,N_38336,N_39708);
and U41890 (N_41890,N_31110,N_32403);
nor U41891 (N_41891,N_39142,N_31653);
xor U41892 (N_41892,N_38210,N_32741);
or U41893 (N_41893,N_38264,N_36012);
nand U41894 (N_41894,N_33226,N_36139);
nor U41895 (N_41895,N_34175,N_37944);
and U41896 (N_41896,N_37834,N_38647);
nor U41897 (N_41897,N_34733,N_36214);
nor U41898 (N_41898,N_35263,N_39250);
xnor U41899 (N_41899,N_37897,N_34301);
and U41900 (N_41900,N_35011,N_39575);
nand U41901 (N_41901,N_32849,N_33959);
nand U41902 (N_41902,N_33855,N_37746);
nand U41903 (N_41903,N_39212,N_33519);
nand U41904 (N_41904,N_32388,N_37790);
and U41905 (N_41905,N_37526,N_36460);
nor U41906 (N_41906,N_35396,N_36998);
nor U41907 (N_41907,N_33329,N_36893);
or U41908 (N_41908,N_38501,N_35238);
or U41909 (N_41909,N_33140,N_39629);
or U41910 (N_41910,N_30065,N_31739);
and U41911 (N_41911,N_33358,N_37833);
nand U41912 (N_41912,N_31469,N_38235);
xor U41913 (N_41913,N_35382,N_34081);
nor U41914 (N_41914,N_39072,N_35342);
and U41915 (N_41915,N_34487,N_36021);
xnor U41916 (N_41916,N_36674,N_32668);
nand U41917 (N_41917,N_31423,N_36305);
or U41918 (N_41918,N_34820,N_39592);
xor U41919 (N_41919,N_37349,N_36003);
nor U41920 (N_41920,N_31036,N_34274);
or U41921 (N_41921,N_35300,N_38204);
nand U41922 (N_41922,N_31098,N_31092);
nor U41923 (N_41923,N_31053,N_36661);
nand U41924 (N_41924,N_33457,N_30520);
and U41925 (N_41925,N_30840,N_37063);
or U41926 (N_41926,N_33615,N_31297);
nand U41927 (N_41927,N_30025,N_35469);
and U41928 (N_41928,N_38858,N_31086);
nor U41929 (N_41929,N_38642,N_38416);
or U41930 (N_41930,N_34505,N_39772);
or U41931 (N_41931,N_33014,N_36455);
xnor U41932 (N_41932,N_35818,N_35910);
and U41933 (N_41933,N_32759,N_39002);
nor U41934 (N_41934,N_37896,N_38230);
or U41935 (N_41935,N_30894,N_32149);
nor U41936 (N_41936,N_33955,N_38702);
or U41937 (N_41937,N_39166,N_38039);
nand U41938 (N_41938,N_39411,N_34117);
xor U41939 (N_41939,N_37782,N_30169);
or U41940 (N_41940,N_38341,N_38837);
and U41941 (N_41941,N_36367,N_30436);
nand U41942 (N_41942,N_39121,N_34958);
nor U41943 (N_41943,N_36696,N_33361);
xor U41944 (N_41944,N_39988,N_38980);
nor U41945 (N_41945,N_34448,N_39057);
nor U41946 (N_41946,N_35973,N_32322);
and U41947 (N_41947,N_32185,N_31932);
xnor U41948 (N_41948,N_38959,N_31985);
and U41949 (N_41949,N_31702,N_32810);
and U41950 (N_41950,N_35514,N_38812);
nand U41951 (N_41951,N_36099,N_32034);
and U41952 (N_41952,N_34636,N_31751);
nand U41953 (N_41953,N_32833,N_37227);
and U41954 (N_41954,N_32246,N_31241);
xor U41955 (N_41955,N_39748,N_35885);
or U41956 (N_41956,N_37577,N_37989);
and U41957 (N_41957,N_38604,N_32325);
nand U41958 (N_41958,N_39518,N_34050);
nand U41959 (N_41959,N_36669,N_36603);
nand U41960 (N_41960,N_32489,N_30034);
and U41961 (N_41961,N_36074,N_30757);
and U41962 (N_41962,N_31647,N_38684);
nand U41963 (N_41963,N_37946,N_31118);
and U41964 (N_41964,N_32777,N_39832);
nand U41965 (N_41965,N_34291,N_39001);
and U41966 (N_41966,N_30384,N_36582);
or U41967 (N_41967,N_32355,N_30531);
nor U41968 (N_41968,N_36077,N_33312);
or U41969 (N_41969,N_35418,N_34918);
or U41970 (N_41970,N_38313,N_33699);
nand U41971 (N_41971,N_39793,N_33023);
nand U41972 (N_41972,N_39829,N_33706);
and U41973 (N_41973,N_37452,N_34250);
and U41974 (N_41974,N_33167,N_30086);
or U41975 (N_41975,N_36683,N_33389);
and U41976 (N_41976,N_35506,N_32745);
nor U41977 (N_41977,N_34727,N_39686);
or U41978 (N_41978,N_38903,N_39383);
nor U41979 (N_41979,N_37830,N_37915);
xor U41980 (N_41980,N_34753,N_37594);
nor U41981 (N_41981,N_38409,N_35360);
or U41982 (N_41982,N_33766,N_35041);
and U41983 (N_41983,N_32828,N_38797);
or U41984 (N_41984,N_30260,N_36784);
nand U41985 (N_41985,N_36130,N_37415);
or U41986 (N_41986,N_35093,N_31893);
nand U41987 (N_41987,N_32730,N_37599);
and U41988 (N_41988,N_37307,N_38240);
and U41989 (N_41989,N_32527,N_30087);
or U41990 (N_41990,N_39839,N_37733);
xor U41991 (N_41991,N_39378,N_32150);
xor U41992 (N_41992,N_38828,N_34408);
nor U41993 (N_41993,N_33518,N_32087);
and U41994 (N_41994,N_38988,N_35176);
and U41995 (N_41995,N_36019,N_32871);
and U41996 (N_41996,N_33571,N_38948);
nand U41997 (N_41997,N_36166,N_30031);
nand U41998 (N_41998,N_39589,N_35325);
nand U41999 (N_41999,N_32430,N_33971);
or U42000 (N_42000,N_33905,N_32993);
and U42001 (N_42001,N_31750,N_36124);
or U42002 (N_42002,N_39396,N_36199);
or U42003 (N_42003,N_39479,N_30512);
nand U42004 (N_42004,N_30841,N_32991);
xnor U42005 (N_42005,N_36497,N_33668);
or U42006 (N_42006,N_37825,N_35705);
or U42007 (N_42007,N_38050,N_33813);
or U42008 (N_42008,N_38620,N_39854);
nor U42009 (N_42009,N_35574,N_39558);
nand U42010 (N_42010,N_37774,N_38339);
nand U42011 (N_42011,N_38593,N_39309);
xor U42012 (N_42012,N_34497,N_32384);
or U42013 (N_42013,N_31058,N_30878);
xor U42014 (N_42014,N_38900,N_38678);
or U42015 (N_42015,N_39580,N_38293);
and U42016 (N_42016,N_36415,N_32252);
nor U42017 (N_42017,N_35950,N_34935);
nand U42018 (N_42018,N_33261,N_32302);
nor U42019 (N_42019,N_33164,N_30385);
nand U42020 (N_42020,N_33150,N_36301);
nor U42021 (N_42021,N_39387,N_36387);
xor U42022 (N_42022,N_36008,N_31589);
and U42023 (N_42023,N_33248,N_34822);
nor U42024 (N_42024,N_37688,N_37024);
nand U42025 (N_42025,N_38238,N_35203);
or U42026 (N_42026,N_33557,N_39870);
xnor U42027 (N_42027,N_38075,N_35085);
nand U42028 (N_42028,N_32947,N_38288);
and U42029 (N_42029,N_37208,N_39417);
or U42030 (N_42030,N_33267,N_38150);
nor U42031 (N_42031,N_33224,N_39488);
or U42032 (N_42032,N_33317,N_30517);
nand U42033 (N_42033,N_37023,N_37858);
or U42034 (N_42034,N_38408,N_37379);
nor U42035 (N_42035,N_33814,N_37872);
nand U42036 (N_42036,N_35379,N_30449);
or U42037 (N_42037,N_36625,N_33725);
nand U42038 (N_42038,N_33931,N_39796);
nor U42039 (N_42039,N_31944,N_35698);
or U42040 (N_42040,N_35627,N_33178);
nand U42041 (N_42041,N_33791,N_33924);
nor U42042 (N_42042,N_33169,N_34859);
nand U42043 (N_42043,N_38564,N_37517);
and U42044 (N_42044,N_34025,N_30944);
and U42045 (N_42045,N_33538,N_39693);
nor U42046 (N_42046,N_38178,N_39601);
nand U42047 (N_42047,N_35302,N_39240);
or U42048 (N_42048,N_32804,N_32876);
nand U42049 (N_42049,N_38933,N_35457);
nor U42050 (N_42050,N_30470,N_37477);
or U42051 (N_42051,N_35974,N_36220);
nand U42052 (N_42052,N_38973,N_33370);
xor U42053 (N_42053,N_39516,N_32964);
and U42054 (N_42054,N_35695,N_32095);
nor U42055 (N_42055,N_34019,N_30577);
or U42056 (N_42056,N_31586,N_36675);
and U42057 (N_42057,N_35788,N_36920);
nor U42058 (N_42058,N_37979,N_34788);
nor U42059 (N_42059,N_32512,N_34001);
nand U42060 (N_42060,N_39401,N_31275);
and U42061 (N_42061,N_35198,N_39226);
or U42062 (N_42062,N_35061,N_36174);
or U42063 (N_42063,N_30396,N_31179);
nor U42064 (N_42064,N_30559,N_33249);
nor U42065 (N_42065,N_32865,N_39187);
or U42066 (N_42066,N_38740,N_36259);
or U42067 (N_42067,N_31020,N_38736);
and U42068 (N_42068,N_36872,N_34744);
or U42069 (N_42069,N_36847,N_32962);
nor U42070 (N_42070,N_36227,N_34502);
nor U42071 (N_42071,N_30652,N_36109);
nand U42072 (N_42072,N_39200,N_31657);
or U42073 (N_42073,N_32013,N_35642);
xnor U42074 (N_42074,N_32129,N_32607);
and U42075 (N_42075,N_37020,N_33506);
nand U42076 (N_42076,N_34435,N_38147);
or U42077 (N_42077,N_30288,N_35499);
and U42078 (N_42078,N_37634,N_39769);
and U42079 (N_42079,N_33477,N_33139);
nand U42080 (N_42080,N_38474,N_38058);
nor U42081 (N_42081,N_36204,N_32196);
nor U42082 (N_42082,N_34646,N_38578);
and U42083 (N_42083,N_36323,N_38317);
and U42084 (N_42084,N_36758,N_34932);
nor U42085 (N_42085,N_34191,N_38634);
nand U42086 (N_42086,N_34443,N_34144);
or U42087 (N_42087,N_35920,N_36453);
or U42088 (N_42088,N_35617,N_37868);
or U42089 (N_42089,N_39736,N_36723);
and U42090 (N_42090,N_36394,N_35282);
nand U42091 (N_42091,N_39956,N_30489);
xnor U42092 (N_42092,N_35113,N_33103);
and U42093 (N_42093,N_38358,N_37041);
nand U42094 (N_42094,N_34231,N_33730);
nor U42095 (N_42095,N_31556,N_38982);
and U42096 (N_42096,N_31103,N_33427);
nand U42097 (N_42097,N_37453,N_36185);
nor U42098 (N_42098,N_35995,N_34148);
xor U42099 (N_42099,N_39559,N_30922);
nand U42100 (N_42100,N_34254,N_31836);
or U42101 (N_42101,N_32721,N_37949);
xor U42102 (N_42102,N_30910,N_37030);
nor U42103 (N_42103,N_30712,N_36917);
or U42104 (N_42104,N_31583,N_32494);
and U42105 (N_42105,N_39034,N_36619);
nor U42106 (N_42106,N_38519,N_35308);
nor U42107 (N_42107,N_39453,N_30519);
and U42108 (N_42108,N_33561,N_30666);
nor U42109 (N_42109,N_31385,N_32885);
nand U42110 (N_42110,N_36634,N_31727);
and U42111 (N_42111,N_31131,N_37148);
or U42112 (N_42112,N_39201,N_37895);
nand U42113 (N_42113,N_30055,N_30721);
nor U42114 (N_42114,N_34960,N_33201);
nand U42115 (N_42115,N_37932,N_30579);
nor U42116 (N_42116,N_30624,N_32219);
and U42117 (N_42117,N_37547,N_37487);
xnor U42118 (N_42118,N_35849,N_36232);
nand U42119 (N_42119,N_33612,N_38896);
nand U42120 (N_42120,N_38882,N_36764);
nand U42121 (N_42121,N_36608,N_30830);
xor U42122 (N_42122,N_35232,N_31382);
or U42123 (N_42123,N_30993,N_39916);
nand U42124 (N_42124,N_30518,N_37315);
and U42125 (N_42125,N_38395,N_38779);
xnor U42126 (N_42126,N_38576,N_30988);
nand U42127 (N_42127,N_34920,N_38803);
nor U42128 (N_42128,N_35278,N_36065);
and U42129 (N_42129,N_37090,N_39220);
and U42130 (N_42130,N_38983,N_39008);
nand U42131 (N_42131,N_36774,N_36867);
or U42132 (N_42132,N_33456,N_36393);
or U42133 (N_42133,N_31650,N_35720);
nand U42134 (N_42134,N_31645,N_32952);
nand U42135 (N_42135,N_37556,N_33800);
or U42136 (N_42136,N_36585,N_39264);
nand U42137 (N_42137,N_31187,N_32709);
and U42138 (N_42138,N_33740,N_35107);
or U42139 (N_42139,N_36982,N_39992);
nand U42140 (N_42140,N_31817,N_34879);
nand U42141 (N_42141,N_32247,N_36870);
nand U42142 (N_42142,N_35979,N_38223);
or U42143 (N_42143,N_38860,N_37036);
nand U42144 (N_42144,N_39744,N_38995);
nand U42145 (N_42145,N_31695,N_33231);
nand U42146 (N_42146,N_30140,N_32350);
and U42147 (N_42147,N_33875,N_37196);
nand U42148 (N_42148,N_32706,N_37101);
or U42149 (N_42149,N_32205,N_31784);
and U42150 (N_42150,N_37493,N_31443);
nor U42151 (N_42151,N_32103,N_37582);
or U42152 (N_42152,N_37377,N_33767);
nor U42153 (N_42153,N_30782,N_33381);
nor U42154 (N_42154,N_37995,N_32731);
and U42155 (N_42155,N_39883,N_31066);
nor U42156 (N_42156,N_37649,N_34366);
xnor U42157 (N_42157,N_34761,N_31976);
or U42158 (N_42158,N_35961,N_30204);
xnor U42159 (N_42159,N_36789,N_36620);
nor U42160 (N_42160,N_37120,N_36930);
or U42161 (N_42161,N_37885,N_30008);
nor U42162 (N_42162,N_39269,N_36037);
or U42163 (N_42163,N_31729,N_34604);
xor U42164 (N_42164,N_31678,N_39965);
and U42165 (N_42165,N_36979,N_39636);
xor U42166 (N_42166,N_37280,N_37423);
nor U42167 (N_42167,N_39425,N_36641);
nand U42168 (N_42168,N_31231,N_37180);
and U42169 (N_42169,N_35196,N_31743);
and U42170 (N_42170,N_32214,N_30777);
and U42171 (N_42171,N_38782,N_37665);
nand U42172 (N_42172,N_37124,N_37999);
nor U42173 (N_42173,N_38347,N_39267);
nor U42174 (N_42174,N_38854,N_37238);
nor U42175 (N_42175,N_35972,N_38018);
nand U42176 (N_42176,N_39490,N_32248);
xor U42177 (N_42177,N_31759,N_34843);
nor U42178 (N_42178,N_36544,N_32606);
and U42179 (N_42179,N_30775,N_39249);
or U42180 (N_42180,N_39486,N_37016);
and U42181 (N_42181,N_31199,N_38867);
or U42182 (N_42182,N_33065,N_30553);
or U42183 (N_42183,N_33544,N_31774);
nor U42184 (N_42184,N_32677,N_38486);
or U42185 (N_42185,N_38306,N_36057);
nand U42186 (N_42186,N_32515,N_37832);
and U42187 (N_42187,N_30781,N_36822);
nand U42188 (N_42188,N_37700,N_38599);
or U42189 (N_42189,N_30605,N_34055);
or U42190 (N_42190,N_39183,N_30295);
nor U42191 (N_42191,N_31257,N_38902);
nand U42192 (N_42192,N_34273,N_36976);
nor U42193 (N_42193,N_37431,N_31982);
and U42194 (N_42194,N_36747,N_37104);
or U42195 (N_42195,N_34583,N_33898);
nor U42196 (N_42196,N_37059,N_34786);
or U42197 (N_42197,N_39807,N_32821);
and U42198 (N_42198,N_34725,N_32757);
or U42199 (N_42199,N_32243,N_37163);
nand U42200 (N_42200,N_33785,N_32015);
nand U42201 (N_42201,N_30285,N_39043);
xnor U42202 (N_42202,N_35065,N_37748);
nor U42203 (N_42203,N_32816,N_31080);
and U42204 (N_42204,N_30653,N_39836);
and U42205 (N_42205,N_35845,N_30917);
nor U42206 (N_42206,N_32888,N_35217);
nor U42207 (N_42207,N_30765,N_34063);
nor U42208 (N_42208,N_30769,N_32143);
and U42209 (N_42209,N_33876,N_31675);
xnor U42210 (N_42210,N_30259,N_35591);
nand U42211 (N_42211,N_36374,N_38763);
xor U42212 (N_42212,N_31927,N_36060);
nor U42213 (N_42213,N_31046,N_34524);
xor U42214 (N_42214,N_33040,N_32467);
nor U42215 (N_42215,N_33513,N_31211);
nand U42216 (N_42216,N_38367,N_35712);
and U42217 (N_42217,N_38000,N_37682);
or U42218 (N_42218,N_39901,N_37926);
and U42219 (N_42219,N_34912,N_32349);
nand U42220 (N_42220,N_36605,N_31596);
xor U42221 (N_42221,N_35899,N_35641);
and U42222 (N_42222,N_36470,N_32483);
and U42223 (N_42223,N_38383,N_34942);
xnor U42224 (N_42224,N_34897,N_36985);
nor U42225 (N_42225,N_37290,N_33591);
and U42226 (N_42226,N_32300,N_37407);
nand U42227 (N_42227,N_39712,N_31901);
and U42228 (N_42228,N_35771,N_33241);
xor U42229 (N_42229,N_39336,N_39582);
or U42230 (N_42230,N_31991,N_38861);
xor U42231 (N_42231,N_32019,N_35944);
nor U42232 (N_42232,N_32978,N_37852);
or U42233 (N_42233,N_33337,N_36397);
nor U42234 (N_42234,N_39153,N_34657);
nor U42235 (N_42235,N_36117,N_34895);
nand U42236 (N_42236,N_30818,N_33608);
or U42237 (N_42237,N_38908,N_32056);
nand U42238 (N_42238,N_36266,N_30619);
nand U42239 (N_42239,N_33059,N_33196);
nor U42240 (N_42240,N_38072,N_34531);
and U42241 (N_42241,N_30851,N_33435);
and U42242 (N_42242,N_31514,N_33690);
or U42243 (N_42243,N_33465,N_39284);
nor U42244 (N_42244,N_39700,N_30329);
nor U42245 (N_42245,N_30111,N_39848);
nor U42246 (N_42246,N_35233,N_30723);
or U42247 (N_42247,N_37071,N_36085);
nand U42248 (N_42248,N_30790,N_36462);
nand U42249 (N_42249,N_33602,N_39313);
and U42250 (N_42250,N_36194,N_34202);
xnor U42251 (N_42251,N_30737,N_38977);
nor U42252 (N_42252,N_32604,N_33461);
nand U42253 (N_42253,N_31796,N_34599);
nor U42254 (N_42254,N_34237,N_32213);
and U42255 (N_42255,N_31307,N_37003);
xor U42256 (N_42256,N_33371,N_39646);
and U42257 (N_42257,N_32609,N_39964);
or U42258 (N_42258,N_36183,N_34662);
or U42259 (N_42259,N_30866,N_30325);
or U42260 (N_42260,N_37575,N_37427);
nor U42261 (N_42261,N_39886,N_30142);
or U42262 (N_42262,N_39915,N_31091);
nor U42263 (N_42263,N_33517,N_38691);
and U42264 (N_42264,N_31249,N_35507);
or U42265 (N_42265,N_38140,N_39370);
or U42266 (N_42266,N_32352,N_36845);
and U42267 (N_42267,N_39420,N_36780);
nor U42268 (N_42268,N_39382,N_31478);
nor U42269 (N_42269,N_34973,N_31634);
xor U42270 (N_42270,N_30867,N_33343);
xnor U42271 (N_42271,N_39362,N_34404);
nor U42272 (N_42272,N_31473,N_31595);
nand U42273 (N_42273,N_36038,N_39773);
or U42274 (N_42274,N_35837,N_37338);
xor U42275 (N_42275,N_39888,N_38284);
and U42276 (N_42276,N_36105,N_36287);
and U42277 (N_42277,N_34219,N_33983);
nor U42278 (N_42278,N_31448,N_36604);
and U42279 (N_42279,N_36618,N_30337);
nand U42280 (N_42280,N_32703,N_33386);
nand U42281 (N_42281,N_36862,N_39208);
nor U42282 (N_42282,N_39645,N_38669);
nand U42283 (N_42283,N_39098,N_34141);
and U42284 (N_42284,N_32672,N_31994);
or U42285 (N_42285,N_37595,N_37993);
or U42286 (N_42286,N_37717,N_34305);
and U42287 (N_42287,N_32107,N_32653);
nor U42288 (N_42288,N_33443,N_36616);
and U42289 (N_42289,N_39452,N_39438);
nor U42290 (N_42290,N_37645,N_33131);
and U42291 (N_42291,N_32880,N_36645);
nand U42292 (N_42292,N_38035,N_31943);
or U42293 (N_42293,N_31592,N_35707);
nand U42294 (N_42294,N_39662,N_32917);
nand U42295 (N_42295,N_33374,N_30215);
and U42296 (N_42296,N_36490,N_31047);
or U42297 (N_42297,N_37504,N_35477);
nand U42298 (N_42298,N_32064,N_31026);
nor U42299 (N_42299,N_31314,N_39445);
and U42300 (N_42300,N_31706,N_32858);
nand U42301 (N_42301,N_31128,N_33976);
and U42302 (N_42302,N_39257,N_38359);
and U42303 (N_42303,N_30172,N_32415);
nand U42304 (N_42304,N_30949,N_34003);
nor U42305 (N_42305,N_36858,N_31406);
or U42306 (N_42306,N_34993,N_38053);
and U42307 (N_42307,N_34536,N_36314);
or U42308 (N_42308,N_31929,N_32942);
and U42309 (N_42309,N_36951,N_34876);
and U42310 (N_42310,N_34458,N_34390);
and U42311 (N_42311,N_37256,N_39639);
nand U42312 (N_42312,N_32290,N_35779);
nand U42313 (N_42313,N_31805,N_38148);
xnor U42314 (N_42314,N_35714,N_36178);
xnor U42315 (N_42315,N_31253,N_39887);
or U42316 (N_42316,N_38687,N_31666);
nand U42317 (N_42317,N_33935,N_38876);
nand U42318 (N_42318,N_34376,N_32260);
or U42319 (N_42319,N_36505,N_34869);
and U42320 (N_42320,N_37243,N_30770);
nor U42321 (N_42321,N_39415,N_31365);
and U42322 (N_42322,N_32768,N_33879);
and U42323 (N_42323,N_37615,N_33790);
xor U42324 (N_42324,N_33464,N_35015);
and U42325 (N_42325,N_31498,N_35139);
and U42326 (N_42326,N_31776,N_39397);
nor U42327 (N_42327,N_34707,N_34379);
and U42328 (N_42328,N_32297,N_35864);
and U42329 (N_42329,N_39233,N_32484);
nor U42330 (N_42330,N_35917,N_37385);
and U42331 (N_42331,N_30691,N_38403);
nand U42332 (N_42332,N_38880,N_32590);
nor U42333 (N_42333,N_30021,N_30315);
or U42334 (N_42334,N_35334,N_39999);
and U42335 (N_42335,N_38999,N_31078);
nand U42336 (N_42336,N_31779,N_33749);
nor U42337 (N_42337,N_37621,N_36709);
nor U42338 (N_42338,N_33526,N_35902);
nor U42339 (N_42339,N_33357,N_31437);
xor U42340 (N_42340,N_30671,N_37534);
xnor U42341 (N_42341,N_34675,N_36433);
or U42342 (N_42342,N_33229,N_33474);
and U42343 (N_42343,N_36285,N_31313);
and U42344 (N_42344,N_36066,N_38384);
and U42345 (N_42345,N_38622,N_38439);
or U42346 (N_42346,N_30787,N_30440);
xor U42347 (N_42347,N_36402,N_36311);
or U42348 (N_42348,N_37706,N_39800);
nor U42349 (N_42349,N_35736,N_39426);
xor U42350 (N_42350,N_34810,N_31484);
nor U42351 (N_42351,N_34589,N_37963);
or U42352 (N_42352,N_36562,N_33105);
or U42353 (N_42353,N_32337,N_34277);
xnor U42354 (N_42354,N_31778,N_30156);
nor U42355 (N_42355,N_32222,N_37223);
and U42356 (N_42356,N_39302,N_34127);
or U42357 (N_42357,N_35024,N_36627);
nor U42358 (N_42358,N_37119,N_39584);
and U42359 (N_42359,N_37792,N_38924);
or U42360 (N_42360,N_31549,N_34307);
and U42361 (N_42361,N_37849,N_34797);
xnor U42362 (N_42362,N_36719,N_34943);
nand U42363 (N_42363,N_36676,N_37713);
nand U42364 (N_42364,N_31554,N_34563);
nor U42365 (N_42365,N_38485,N_37419);
or U42366 (N_42366,N_31161,N_36075);
and U42367 (N_42367,N_38682,N_34450);
or U42368 (N_42368,N_30268,N_34036);
or U42369 (N_42369,N_38866,N_33682);
and U42370 (N_42370,N_32999,N_36660);
or U42371 (N_42371,N_30341,N_34773);
or U42372 (N_42372,N_38376,N_38830);
nand U42373 (N_42373,N_37668,N_34829);
or U42374 (N_42374,N_33965,N_36452);
or U42375 (N_42375,N_33834,N_35438);
and U42376 (N_42376,N_37305,N_32847);
nor U42377 (N_42377,N_39197,N_33294);
xor U42378 (N_42378,N_36831,N_32201);
nor U42379 (N_42379,N_36668,N_38906);
nand U42380 (N_42380,N_36670,N_33644);
or U42381 (N_42381,N_34846,N_36047);
nand U42382 (N_42382,N_33136,N_32277);
xnor U42383 (N_42383,N_39907,N_35264);
xnor U42384 (N_42384,N_37935,N_31075);
or U42385 (N_42385,N_38278,N_33990);
xnor U42386 (N_42386,N_37918,N_37092);
nor U42387 (N_42387,N_33332,N_33523);
xor U42388 (N_42388,N_37725,N_38133);
nor U42389 (N_42389,N_38639,N_33291);
nand U42390 (N_42390,N_31917,N_33509);
nor U42391 (N_42391,N_38730,N_36898);
and U42392 (N_42392,N_37251,N_35765);
and U42393 (N_42393,N_36111,N_34590);
and U42394 (N_42394,N_38343,N_32411);
and U42395 (N_42395,N_39882,N_38227);
nand U42396 (N_42396,N_31127,N_34714);
nand U42397 (N_42397,N_31482,N_36596);
and U42398 (N_42398,N_30437,N_31327);
nor U42399 (N_42399,N_32182,N_39031);
nor U42400 (N_42400,N_35194,N_34159);
nor U42401 (N_42401,N_34185,N_32451);
nor U42402 (N_42402,N_36005,N_37683);
or U42403 (N_42403,N_35371,N_36802);
nor U42404 (N_42404,N_39419,N_32457);
or U42405 (N_42405,N_39562,N_37123);
or U42406 (N_42406,N_32179,N_30598);
nor U42407 (N_42407,N_30746,N_35261);
or U42408 (N_42408,N_39902,N_32323);
nor U42409 (N_42409,N_35509,N_36179);
and U42410 (N_42410,N_31713,N_39113);
and U42411 (N_42411,N_35568,N_39022);
and U42412 (N_42412,N_32427,N_34518);
nor U42413 (N_42413,N_35454,N_30903);
nor U42414 (N_42414,N_37128,N_32027);
and U42415 (N_42415,N_33499,N_33952);
nor U42416 (N_42416,N_31925,N_39395);
nor U42417 (N_42417,N_33073,N_36628);
nand U42418 (N_42418,N_37283,N_31633);
nand U42419 (N_42419,N_33901,N_32875);
and U42420 (N_42420,N_35722,N_38735);
nand U42421 (N_42421,N_30647,N_34794);
and U42422 (N_42422,N_38619,N_36389);
nor U42423 (N_42423,N_38659,N_38216);
or U42424 (N_42424,N_36636,N_32631);
nor U42425 (N_42425,N_39606,N_37336);
nor U42426 (N_42426,N_34234,N_36481);
or U42427 (N_42427,N_32922,N_36249);
or U42428 (N_42428,N_39041,N_33975);
nand U42429 (N_42429,N_35083,N_34512);
and U42430 (N_42430,N_35350,N_32926);
xor U42431 (N_42431,N_32009,N_39231);
and U42432 (N_42432,N_33033,N_35033);
nand U42433 (N_42433,N_35461,N_36875);
nand U42434 (N_42434,N_33480,N_38875);
and U42435 (N_42435,N_37091,N_34528);
xor U42436 (N_42436,N_38654,N_36244);
nor U42437 (N_42437,N_34570,N_39354);
nor U42438 (N_42438,N_39077,N_33436);
or U42439 (N_42439,N_34260,N_31065);
nand U42440 (N_42440,N_37854,N_37417);
nand U42441 (N_42441,N_30880,N_38258);
nand U42442 (N_42442,N_39875,N_32367);
nor U42443 (N_42443,N_36209,N_37082);
or U42444 (N_42444,N_31221,N_30715);
nand U42445 (N_42445,N_34053,N_35026);
nor U42446 (N_42446,N_34446,N_33492);
nand U42447 (N_42447,N_37322,N_36812);
nand U42448 (N_42448,N_38609,N_37491);
nor U42449 (N_42449,N_36689,N_35202);
and U42450 (N_42450,N_33284,N_37034);
nand U42451 (N_42451,N_37229,N_32803);
nand U42452 (N_42452,N_33338,N_33628);
or U42453 (N_42453,N_37342,N_30725);
nor U42454 (N_42454,N_31676,N_37094);
nand U42455 (N_42455,N_37619,N_39004);
nand U42456 (N_42456,N_39303,N_30612);
and U42457 (N_42457,N_34451,N_33124);
nor U42458 (N_42458,N_35279,N_35134);
nand U42459 (N_42459,N_34371,N_39247);
nand U42460 (N_42460,N_33355,N_38489);
and U42461 (N_42461,N_31621,N_34768);
xor U42462 (N_42462,N_38955,N_31139);
and U42463 (N_42463,N_32779,N_37984);
or U42464 (N_42464,N_31259,N_39812);
and U42465 (N_42465,N_32173,N_36176);
and U42466 (N_42466,N_36716,N_37348);
nor U42467 (N_42467,N_36177,N_33207);
and U42468 (N_42468,N_38543,N_39169);
and U42469 (N_42469,N_39272,N_35793);
nand U42470 (N_42470,N_31715,N_30547);
or U42471 (N_42471,N_32910,N_33872);
xor U42472 (N_42472,N_34342,N_38112);
nand U42473 (N_42473,N_38334,N_31939);
and U42474 (N_42474,N_34611,N_32660);
nor U42475 (N_42475,N_34263,N_33852);
or U42476 (N_42476,N_30909,N_34692);
nor U42477 (N_42477,N_37667,N_37107);
and U42478 (N_42478,N_30564,N_39689);
nor U42479 (N_42479,N_31904,N_39304);
or U42480 (N_42480,N_36482,N_31008);
nor U42481 (N_42481,N_34923,N_31000);
nor U42482 (N_42482,N_35505,N_36371);
nor U42483 (N_42483,N_31277,N_34586);
nand U42484 (N_42484,N_33095,N_34816);
or U42485 (N_42485,N_35983,N_33739);
nand U42486 (N_42486,N_33632,N_34623);
and U42487 (N_42487,N_36924,N_35297);
nor U42488 (N_42488,N_33533,N_33548);
or U42489 (N_42489,N_34468,N_32824);
nor U42490 (N_42490,N_33290,N_37720);
or U42491 (N_42491,N_30872,N_39551);
and U42492 (N_42492,N_34179,N_30561);
and U42493 (N_42493,N_37942,N_31225);
or U42494 (N_42494,N_30377,N_35145);
and U42495 (N_42495,N_32478,N_37270);
nor U42496 (N_42496,N_36792,N_31768);
or U42497 (N_42497,N_37007,N_39217);
nand U42498 (N_42498,N_33922,N_38787);
and U42499 (N_42499,N_31458,N_31995);
and U42500 (N_42500,N_32602,N_31032);
xnor U42501 (N_42501,N_36578,N_35684);
nor U42502 (N_42502,N_35448,N_30410);
nor U42503 (N_42503,N_36607,N_30573);
nand U42504 (N_42504,N_34023,N_35161);
and U42505 (N_42505,N_36392,N_34246);
nand U42506 (N_42506,N_34367,N_34204);
and U42507 (N_42507,N_37780,N_32728);
xor U42508 (N_42508,N_32998,N_35088);
nor U42509 (N_42509,N_39276,N_35407);
nand U42510 (N_42510,N_32044,N_30448);
or U42511 (N_42511,N_32791,N_39205);
nand U42512 (N_42512,N_33727,N_37711);
nor U42513 (N_42513,N_31391,N_35067);
xnor U42514 (N_42514,N_39394,N_32654);
nor U42515 (N_42515,N_39221,N_35835);
nor U42516 (N_42516,N_39060,N_39571);
and U42517 (N_42517,N_31038,N_37894);
and U42518 (N_42518,N_38754,N_37164);
or U42519 (N_42519,N_37592,N_37776);
nand U42520 (N_42520,N_31870,N_30200);
or U42521 (N_42521,N_39894,N_33882);
or U42522 (N_42522,N_37742,N_34488);
nand U42523 (N_42523,N_39360,N_32490);
nand U42524 (N_42524,N_35125,N_37796);
and U42525 (N_42525,N_31374,N_30476);
nor U42526 (N_42526,N_34208,N_39522);
nor U42527 (N_42527,N_30651,N_37193);
or U42528 (N_42528,N_38085,N_32667);
and U42529 (N_42529,N_34720,N_34894);
and U42530 (N_42530,N_35123,N_37652);
nand U42531 (N_42531,N_33044,N_34526);
nand U42532 (N_42532,N_36520,N_33432);
nor U42533 (N_42533,N_35987,N_34251);
and U42534 (N_42534,N_38215,N_34217);
or U42535 (N_42535,N_36276,N_39287);
xor U42536 (N_42536,N_38528,N_36475);
nand U42537 (N_42537,N_36322,N_36161);
or U42538 (N_42538,N_39461,N_32560);
nor U42539 (N_42539,N_38224,N_34535);
nand U42540 (N_42540,N_39926,N_30225);
nand U42541 (N_42541,N_38450,N_31228);
nor U42542 (N_42542,N_38989,N_31911);
nor U42543 (N_42543,N_31109,N_30307);
nand U42544 (N_42544,N_36698,N_39075);
and U42545 (N_42545,N_37936,N_36354);
nand U42546 (N_42546,N_31019,N_39033);
or U42547 (N_42547,N_38946,N_35905);
and U42548 (N_42548,N_30006,N_30220);
nor U42549 (N_42549,N_38392,N_35053);
nor U42550 (N_42550,N_39234,N_39332);
or U42551 (N_42551,N_37289,N_30727);
and U42552 (N_42552,N_31961,N_32556);
or U42553 (N_42553,N_37756,N_34369);
or U42554 (N_42554,N_34648,N_34385);
or U42555 (N_42555,N_33915,N_37264);
nand U42556 (N_42556,N_32423,N_34108);
nor U42557 (N_42557,N_31953,N_36018);
nand U42558 (N_42558,N_39295,N_38120);
xor U42559 (N_42559,N_35930,N_32465);
nand U42560 (N_42560,N_38362,N_32048);
nor U42561 (N_42561,N_31576,N_32752);
nand U42562 (N_42562,N_33611,N_38272);
and U42563 (N_42563,N_34236,N_36574);
nor U42564 (N_42564,N_37512,N_31580);
and U42565 (N_42565,N_33982,N_37459);
nand U42566 (N_42566,N_35383,N_34805);
nand U42567 (N_42567,N_36567,N_34344);
or U42568 (N_42568,N_33209,N_34584);
nor U42569 (N_42569,N_35245,N_32425);
nand U42570 (N_42570,N_32308,N_32085);
and U42571 (N_42571,N_37457,N_39254);
and U42572 (N_42572,N_33120,N_33881);
xnor U42573 (N_42573,N_32152,N_39610);
or U42574 (N_42574,N_39087,N_36291);
and U42575 (N_42575,N_31950,N_30706);
or U42576 (N_42576,N_38236,N_35699);
xor U42577 (N_42577,N_36892,N_34200);
and U42578 (N_42578,N_35815,N_36079);
or U42579 (N_42579,N_32879,N_34196);
xnor U42580 (N_42580,N_37520,N_36267);
nand U42581 (N_42581,N_32436,N_33807);
nor U42582 (N_42582,N_34608,N_30835);
nor U42583 (N_42583,N_33693,N_35426);
nand U42584 (N_42584,N_35573,N_35120);
and U42585 (N_42585,N_36030,N_38101);
and U42586 (N_42586,N_32341,N_32915);
nor U42587 (N_42587,N_33895,N_35425);
xnor U42588 (N_42588,N_30511,N_37058);
or U42589 (N_42589,N_37213,N_32533);
xnor U42590 (N_42590,N_35054,N_30190);
and U42591 (N_42591,N_32069,N_36687);
nor U42592 (N_42592,N_35136,N_39009);
or U42593 (N_42593,N_32689,N_34215);
and U42594 (N_42594,N_38919,N_30354);
or U42595 (N_42595,N_37930,N_34285);
nor U42596 (N_42596,N_30555,N_36031);
nand U42597 (N_42597,N_31445,N_32936);
or U42598 (N_42598,N_38382,N_30209);
and U42599 (N_42599,N_39847,N_34069);
and U42600 (N_42600,N_31610,N_36488);
nand U42601 (N_42601,N_39245,N_33251);
nand U42602 (N_42602,N_30975,N_35397);
nand U42603 (N_42603,N_31789,N_36027);
nand U42604 (N_42604,N_33453,N_35635);
xnor U42605 (N_42605,N_31907,N_38369);
or U42606 (N_42606,N_33703,N_31474);
nor U42607 (N_42607,N_38794,N_39616);
nand U42608 (N_42608,N_31884,N_33803);
and U42609 (N_42609,N_38449,N_32460);
nand U42610 (N_42610,N_32301,N_34975);
nand U42611 (N_42611,N_30920,N_38589);
or U42612 (N_42612,N_31479,N_36164);
nor U42613 (N_42613,N_33896,N_31918);
or U42614 (N_42614,N_31326,N_33558);
and U42615 (N_42615,N_35173,N_31315);
nand U42616 (N_42616,N_30617,N_39727);
nand U42617 (N_42617,N_35610,N_31938);
or U42618 (N_42618,N_34633,N_39866);
or U42619 (N_42619,N_36825,N_31291);
nand U42620 (N_42620,N_38884,N_36306);
nor U42621 (N_42621,N_38709,N_37618);
nand U42622 (N_42622,N_36559,N_38951);
xnor U42623 (N_42623,N_35229,N_32749);
xnor U42624 (N_42624,N_33049,N_33651);
or U42625 (N_42625,N_39006,N_30266);
nor U42626 (N_42626,N_34815,N_31373);
or U42627 (N_42627,N_31237,N_37178);
or U42628 (N_42628,N_30015,N_39745);
nor U42629 (N_42629,N_35467,N_32452);
nor U42630 (N_42630,N_37411,N_39991);
xor U42631 (N_42631,N_33757,N_32071);
or U42632 (N_42632,N_38329,N_37382);
nor U42633 (N_42633,N_30064,N_32620);
xor U42634 (N_42634,N_32274,N_35386);
and U42635 (N_42635,N_37209,N_38636);
and U42636 (N_42636,N_34123,N_37001);
xnor U42637 (N_42637,N_37162,N_35490);
nand U42638 (N_42638,N_39995,N_36359);
or U42639 (N_42639,N_35624,N_34058);
nand U42640 (N_42640,N_35314,N_37327);
nor U42641 (N_42641,N_31424,N_38070);
nor U42642 (N_42642,N_32665,N_36664);
nand U42643 (N_42643,N_35252,N_38003);
or U42644 (N_42644,N_30901,N_37640);
or U42645 (N_42645,N_38507,N_38960);
nand U42646 (N_42646,N_30496,N_34416);
nor U42647 (N_42647,N_32645,N_38807);
nor U42648 (N_42648,N_30580,N_31603);
nand U42649 (N_42649,N_37331,N_33634);
xor U42650 (N_42650,N_35990,N_38446);
nor U42651 (N_42651,N_32712,N_32898);
nor U42652 (N_42652,N_37934,N_36318);
nor U42653 (N_42653,N_32004,N_33242);
nor U42654 (N_42654,N_39538,N_33996);
and U42655 (N_42655,N_30183,N_36261);
nand U42656 (N_42656,N_31806,N_38821);
nor U42657 (N_42657,N_30076,N_30952);
nor U42658 (N_42658,N_35100,N_30983);
or U42659 (N_42659,N_37334,N_32521);
or U42660 (N_42660,N_31869,N_38673);
nand U42661 (N_42661,N_39019,N_31418);
and U42662 (N_42662,N_36432,N_36801);
nand U42663 (N_42663,N_34481,N_33050);
and U42664 (N_42664,N_31219,N_36823);
and U42665 (N_42665,N_33280,N_35458);
nor U42666 (N_42666,N_38652,N_36503);
or U42667 (N_42667,N_31331,N_38244);
and U42668 (N_42668,N_33320,N_35584);
nor U42669 (N_42669,N_30812,N_33047);
nand U42670 (N_42670,N_36642,N_37316);
or U42671 (N_42671,N_34206,N_38766);
nor U42672 (N_42672,N_35375,N_37184);
or U42673 (N_42673,N_36745,N_36410);
nor U42674 (N_42674,N_39827,N_31033);
and U42675 (N_42675,N_34998,N_30141);
xnor U42676 (N_42676,N_34262,N_39560);
and U42677 (N_42677,N_38720,N_35940);
nor U42678 (N_42678,N_30811,N_39500);
and U42679 (N_42679,N_36986,N_32193);
nand U42680 (N_42680,N_39954,N_32329);
or U42681 (N_42681,N_31349,N_38625);
nor U42682 (N_42682,N_39466,N_36781);
nor U42683 (N_42683,N_31420,N_35936);
or U42684 (N_42684,N_35301,N_36295);
or U42685 (N_42685,N_38624,N_37401);
nor U42686 (N_42686,N_36992,N_38510);
and U42687 (N_42687,N_37458,N_36733);
nand U42688 (N_42688,N_39590,N_37612);
and U42689 (N_42689,N_32461,N_32113);
or U42690 (N_42690,N_33593,N_37836);
nor U42691 (N_42691,N_31468,N_36216);
or U42692 (N_42692,N_34088,N_32559);
nor U42693 (N_42693,N_30977,N_31194);
nor U42694 (N_42694,N_30590,N_32656);
nand U42695 (N_42695,N_32841,N_38451);
nand U42696 (N_42696,N_39224,N_31472);
and U42697 (N_42697,N_37581,N_37099);
nor U42698 (N_42698,N_30024,N_31825);
and U42699 (N_42699,N_34742,N_31148);
nand U42700 (N_42700,N_35682,N_39097);
or U42701 (N_42701,N_35452,N_30677);
nor U42702 (N_42702,N_34567,N_36233);
xor U42703 (N_42703,N_33098,N_31896);
or U42704 (N_42704,N_36663,N_38338);
xnor U42705 (N_42705,N_33629,N_36859);
or U42706 (N_42706,N_34661,N_33697);
nand U42707 (N_42707,N_36446,N_32586);
nor U42708 (N_42708,N_30783,N_31708);
and U42709 (N_42709,N_34427,N_37816);
nor U42710 (N_42710,N_39680,N_37631);
or U42711 (N_42711,N_35304,N_36835);
nand U42712 (N_42712,N_39713,N_31248);
and U42713 (N_42713,N_33071,N_37363);
nand U42714 (N_42714,N_34292,N_30704);
or U42715 (N_42715,N_35723,N_32055);
or U42716 (N_42716,N_30466,N_35660);
nand U42717 (N_42717,N_30167,N_30556);
nor U42718 (N_42718,N_30991,N_38323);
nand U42719 (N_42719,N_35782,N_30300);
nand U42720 (N_42720,N_35991,N_38838);
or U42721 (N_42721,N_37506,N_34216);
and U42722 (N_42722,N_37050,N_32514);
and U42723 (N_42723,N_33397,N_36202);
and U42724 (N_42724,N_37179,N_33186);
and U42725 (N_42725,N_36409,N_35097);
nor U42726 (N_42726,N_31507,N_32227);
and U42727 (N_42727,N_33423,N_31345);
nor U42728 (N_42728,N_30213,N_32259);
and U42729 (N_42729,N_30328,N_30469);
xnor U42730 (N_42730,N_38568,N_39634);
nor U42731 (N_42731,N_33893,N_34877);
xnor U42732 (N_42732,N_38795,N_31238);
or U42733 (N_42733,N_38380,N_30391);
xor U42734 (N_42734,N_32971,N_33672);
nor U42735 (N_42735,N_34203,N_31364);
xor U42736 (N_42736,N_35975,N_37846);
xor U42737 (N_42737,N_37745,N_32041);
nor U42738 (N_42738,N_30481,N_33422);
or U42739 (N_42739,N_36680,N_32310);
or U42740 (N_42740,N_30760,N_33908);
xnor U42741 (N_42741,N_37254,N_34698);
or U42742 (N_42742,N_36899,N_37156);
xnor U42743 (N_42743,N_32950,N_35207);
and U42744 (N_42744,N_32318,N_33369);
nor U42745 (N_42745,N_37418,N_33920);
nor U42746 (N_42746,N_31386,N_38144);
or U42747 (N_42747,N_36807,N_33889);
nor U42748 (N_42748,N_39900,N_34809);
and U42749 (N_42749,N_38171,N_32061);
nand U42750 (N_42750,N_32334,N_37593);
nand U42751 (N_42751,N_34244,N_38241);
and U42752 (N_42752,N_30736,N_33750);
and U42753 (N_42753,N_38274,N_34071);
nand U42754 (N_42754,N_37648,N_38428);
nor U42755 (N_42755,N_39364,N_36830);
nand U42756 (N_42756,N_38499,N_34545);
or U42757 (N_42757,N_37687,N_35562);
nand U42758 (N_42758,N_31762,N_39377);
xnor U42759 (N_42759,N_39710,N_32416);
or U42760 (N_42760,N_38849,N_37011);
or U42761 (N_42761,N_34704,N_34243);
and U42762 (N_42762,N_33470,N_33885);
or U42763 (N_42763,N_31885,N_33469);
or U42764 (N_42764,N_38327,N_37367);
nor U42765 (N_42765,N_37530,N_39080);
xor U42766 (N_42766,N_34517,N_35756);
nor U42767 (N_42767,N_38905,N_33257);
nand U42768 (N_42768,N_35413,N_30711);
nor U42769 (N_42769,N_35817,N_36279);
nor U42770 (N_42770,N_33235,N_33420);
and U42771 (N_42771,N_33659,N_36041);
or U42772 (N_42772,N_34565,N_31661);
nand U42773 (N_42773,N_31045,N_32233);
nor U42774 (N_42774,N_37779,N_38309);
or U42775 (N_42775,N_32228,N_31521);
and U42776 (N_42776,N_32097,N_35153);
nand U42777 (N_42777,N_31624,N_31557);
nor U42778 (N_42778,N_39203,N_31606);
and U42779 (N_42779,N_32469,N_35632);
or U42780 (N_42780,N_32046,N_30389);
or U42781 (N_42781,N_36573,N_36396);
nor U42782 (N_42782,N_39524,N_34644);
and U42783 (N_42783,N_31284,N_36648);
nor U42784 (N_42784,N_36804,N_37257);
xor U42785 (N_42785,N_31044,N_37982);
and U42786 (N_42786,N_31209,N_38125);
nand U42787 (N_42787,N_33138,N_38878);
or U42788 (N_42788,N_31622,N_31810);
nand U42789 (N_42789,N_33486,N_31539);
and U42790 (N_42790,N_35777,N_33524);
and U42791 (N_42791,N_34266,N_30276);
nand U42792 (N_42792,N_32039,N_31501);
or U42793 (N_42793,N_39175,N_39179);
nor U42794 (N_42794,N_33782,N_32058);
nor U42795 (N_42795,N_31280,N_37771);
xor U42796 (N_42796,N_33266,N_31585);
and U42797 (N_42797,N_39032,N_39856);
nand U42798 (N_42798,N_32908,N_38202);
nand U42799 (N_42799,N_36761,N_39116);
and U42800 (N_42800,N_38912,N_35152);
and U42801 (N_42801,N_35240,N_36329);
xor U42802 (N_42802,N_38052,N_32309);
or U42803 (N_42803,N_36254,N_39163);
and U42804 (N_42804,N_37388,N_34825);
nor U42805 (N_42805,N_30978,N_39714);
xnor U42806 (N_42806,N_32974,N_30048);
xor U42807 (N_42807,N_30660,N_37374);
xor U42808 (N_42808,N_34372,N_37383);
or U42809 (N_42809,N_38547,N_34771);
or U42810 (N_42810,N_37781,N_33160);
xnor U42811 (N_42811,N_39216,N_37165);
nor U42812 (N_42812,N_38962,N_35785);
and U42813 (N_42813,N_30690,N_33660);
and U42814 (N_42814,N_33958,N_38732);
or U42815 (N_42815,N_35952,N_35727);
or U42816 (N_42816,N_39648,N_36439);
nand U42817 (N_42817,N_36324,N_39314);
or U42818 (N_42818,N_30240,N_39371);
nor U42819 (N_42819,N_36141,N_30629);
and U42820 (N_42820,N_30728,N_35032);
nand U42821 (N_42821,N_39244,N_33815);
nand U42822 (N_42822,N_31797,N_34741);
or U42823 (N_42823,N_32564,N_33441);
nor U42824 (N_42824,N_39920,N_36933);
nand U42825 (N_42825,N_36062,N_30053);
or U42826 (N_42826,N_34313,N_34136);
and U42827 (N_42827,N_39024,N_38057);
and U42828 (N_42828,N_33647,N_36770);
and U42829 (N_42829,N_34889,N_35799);
nand U42830 (N_42830,N_33076,N_31913);
nor U42831 (N_42831,N_30497,N_39936);
nand U42832 (N_42832,N_32255,N_34329);
nand U42833 (N_42833,N_31076,N_33751);
and U42834 (N_42834,N_32939,N_37624);
nor U42835 (N_42835,N_30388,N_33458);
and U42836 (N_42836,N_39374,N_31441);
nand U42837 (N_42837,N_30615,N_37328);
and U42838 (N_42838,N_38455,N_36480);
nor U42839 (N_42839,N_34808,N_30404);
xnor U42840 (N_42840,N_35317,N_36208);
xor U42841 (N_42841,N_36395,N_33812);
and U42842 (N_42842,N_31283,N_31354);
nand U42843 (N_42843,N_38006,N_31573);
and U42844 (N_42844,N_39760,N_31844);
or U42845 (N_42845,N_38897,N_32470);
or U42846 (N_42846,N_38168,N_39782);
xnor U42847 (N_42847,N_35956,N_36342);
nor U42848 (N_42848,N_36127,N_36678);
or U42849 (N_42849,N_37365,N_35104);
nand U42850 (N_42850,N_35796,N_34471);
and U42851 (N_42851,N_35463,N_38159);
xnor U42852 (N_42852,N_39036,N_39946);
and U42853 (N_42853,N_35494,N_37921);
nand U42854 (N_42854,N_38800,N_36052);
or U42855 (N_42855,N_39161,N_30462);
or U42856 (N_42856,N_36935,N_38063);
nand U42857 (N_42857,N_31997,N_34884);
nand U42858 (N_42858,N_38894,N_35172);
or U42859 (N_42859,N_32955,N_31738);
and U42860 (N_42860,N_38590,N_32362);
nor U42861 (N_42861,N_30516,N_34389);
nand U42862 (N_42862,N_34328,N_30575);
or U42863 (N_42863,N_32169,N_39015);
or U42864 (N_42864,N_30264,N_35557);
or U42865 (N_42865,N_36968,N_36483);
nor U42866 (N_42866,N_36197,N_39674);
and U42867 (N_42867,N_34658,N_35409);
nand U42868 (N_42868,N_32578,N_37444);
or U42869 (N_42869,N_39390,N_38626);
nand U42870 (N_42870,N_30893,N_30676);
or U42871 (N_42871,N_37941,N_38805);
xor U42872 (N_42872,N_31006,N_38817);
nor U42873 (N_42873,N_38299,N_32264);
nor U42874 (N_42874,N_33472,N_36786);
xor U42875 (N_42875,N_33282,N_35739);
and U42876 (N_42876,N_33588,N_39162);
nor U42877 (N_42877,N_38183,N_37826);
and U42878 (N_42878,N_35377,N_37111);
nor U42879 (N_42879,N_34915,N_34997);
nand U42880 (N_42880,N_32697,N_34163);
xor U42881 (N_42881,N_33775,N_39959);
or U42882 (N_42882,N_34135,N_37478);
nand U42883 (N_42883,N_33375,N_36624);
nor U42884 (N_42884,N_35239,N_34622);
nand U42885 (N_42885,N_38164,N_30415);
and U42886 (N_42886,N_32744,N_31967);
nand U42887 (N_42887,N_36756,N_34373);
nand U42888 (N_42888,N_34253,N_38967);
and U42889 (N_42889,N_34851,N_30542);
or U42890 (N_42890,N_32028,N_33412);
xnor U42891 (N_42891,N_31067,N_35670);
xor U42892 (N_42892,N_36598,N_30891);
nand U42893 (N_42893,N_37013,N_38681);
and U42894 (N_42894,N_38505,N_36938);
or U42895 (N_42895,N_30747,N_38410);
or U42896 (N_42896,N_37709,N_32783);
and U42897 (N_42897,N_35563,N_32899);
and U42898 (N_42898,N_37953,N_35231);
or U42899 (N_42899,N_33042,N_33454);
nor U42900 (N_42900,N_30219,N_39990);
or U42901 (N_42901,N_35597,N_37939);
and U42902 (N_42902,N_31265,N_38056);
nor U42903 (N_42903,N_39794,N_32408);
xnor U42904 (N_42904,N_36832,N_38402);
and U42905 (N_42905,N_35850,N_38038);
nor U42906 (N_42906,N_39140,N_35055);
nand U42907 (N_42907,N_33489,N_38118);
or U42908 (N_42908,N_33238,N_34806);
nor U42909 (N_42909,N_30816,N_37112);
nor U42910 (N_42910,N_38333,N_31411);
nor U42911 (N_42911,N_34193,N_36547);
nor U42912 (N_42912,N_34878,N_34083);
nor U42913 (N_42913,N_31489,N_31824);
or U42914 (N_42914,N_37673,N_37586);
or U42915 (N_42915,N_34002,N_31809);
and U42916 (N_42916,N_32223,N_30148);
and U42917 (N_42917,N_31599,N_37821);
and U42918 (N_42918,N_39096,N_30950);
and U42919 (N_42919,N_31129,N_34167);
and U42920 (N_42920,N_38463,N_34858);
xnor U42921 (N_42921,N_36347,N_33504);
nor U42922 (N_42922,N_31733,N_32695);
or U42923 (N_42923,N_31487,N_31233);
xnor U42924 (N_42924,N_32761,N_36253);
xnor U42925 (N_42925,N_35781,N_37109);
nor U42926 (N_42926,N_39103,N_36100);
nand U42927 (N_42927,N_36828,N_36122);
or U42928 (N_42928,N_36067,N_38363);
and U42929 (N_42929,N_31826,N_35605);
nor U42930 (N_42930,N_39210,N_33562);
nor U42931 (N_42931,N_34580,N_35677);
or U42932 (N_42932,N_36533,N_31698);
nor U42933 (N_42933,N_30091,N_32377);
nor U42934 (N_42934,N_38745,N_32226);
nand U42935 (N_42935,N_38688,N_35351);
nor U42936 (N_42936,N_39035,N_39872);
nand U42937 (N_42937,N_36309,N_37859);
or U42938 (N_42938,N_38031,N_38958);
nand U42939 (N_42939,N_34010,N_30439);
or U42940 (N_42940,N_37721,N_34776);
xnor U42941 (N_42941,N_34040,N_37358);
and U42942 (N_42942,N_31494,N_31719);
nand U42943 (N_42943,N_30658,N_33771);
nor U42944 (N_42944,N_31337,N_32330);
or U42945 (N_42945,N_39076,N_38742);
or U42946 (N_42946,N_33698,N_31308);
xor U42947 (N_42947,N_31392,N_37400);
and U42948 (N_42948,N_38956,N_32589);
nand U42949 (N_42949,N_31444,N_38060);
or U42950 (N_42950,N_39189,N_39837);
or U42951 (N_42951,N_33603,N_31692);
and U42952 (N_42952,N_34184,N_33831);
nand U42953 (N_42953,N_31467,N_34474);
and U42954 (N_42954,N_33118,N_32719);
or U42955 (N_42955,N_34764,N_35337);
nand U42956 (N_42956,N_30336,N_34011);
and U42957 (N_42957,N_37754,N_35341);
xor U42958 (N_42958,N_30515,N_39053);
nand U42959 (N_42959,N_38676,N_38444);
nand U42960 (N_42960,N_31665,N_39878);
xor U42961 (N_42961,N_30828,N_37002);
or U42962 (N_42962,N_37722,N_30807);
nand U42963 (N_42963,N_37803,N_36447);
nor U42964 (N_42964,N_34105,N_30306);
nand U42965 (N_42965,N_36275,N_39555);
xor U42966 (N_42966,N_38839,N_30957);
and U42967 (N_42967,N_33910,N_33643);
nand U42968 (N_42968,N_35884,N_35860);
nor U42969 (N_42969,N_38388,N_39497);
and U42970 (N_42970,N_30804,N_33099);
or U42971 (N_42971,N_34573,N_38400);
nand U42972 (N_42972,N_31007,N_38022);
and U42973 (N_42973,N_36682,N_35353);
or U42974 (N_42974,N_35824,N_30719);
nor U42975 (N_42975,N_39439,N_31788);
or U42976 (N_42976,N_33126,N_36714);
and U42977 (N_42977,N_32363,N_33592);
and U42978 (N_42978,N_38308,N_39471);
or U42979 (N_42979,N_34482,N_37613);
nand U42980 (N_42980,N_32890,N_35503);
and U42981 (N_42981,N_30214,N_34671);
nand U42982 (N_42982,N_38579,N_37531);
nor U42983 (N_42983,N_38129,N_38936);
nand U42984 (N_42984,N_35287,N_36922);
or U42985 (N_42985,N_33388,N_34625);
nand U42986 (N_42986,N_38672,N_39715);
xor U42987 (N_42987,N_31734,N_31334);
nand U42988 (N_42988,N_37642,N_32870);
nand U42989 (N_42989,N_32690,N_33890);
and U42990 (N_42990,N_37362,N_31292);
and U42991 (N_42991,N_35171,N_31843);
nand U42992 (N_42992,N_34078,N_36477);
nand U42993 (N_42993,N_37105,N_30918);
nor U42994 (N_42994,N_33789,N_34547);
xnor U42995 (N_42995,N_38026,N_39215);
and U42996 (N_42996,N_39243,N_31571);
nor U42997 (N_42997,N_38704,N_37977);
and U42998 (N_42998,N_36420,N_33177);
nand U42999 (N_42999,N_39962,N_32792);
and U43000 (N_43000,N_35411,N_39895);
nand U43001 (N_43001,N_34046,N_33217);
nand U43002 (N_43002,N_34024,N_38841);
and U43003 (N_43003,N_37591,N_36977);
and U43004 (N_43004,N_39682,N_36103);
nand U43005 (N_43005,N_39979,N_32850);
or U43006 (N_43006,N_30551,N_33206);
and U43007 (N_43007,N_39421,N_33913);
xor U43008 (N_43008,N_32409,N_35784);
nor U43009 (N_43009,N_33939,N_33057);
or U43010 (N_43010,N_34150,N_39994);
and U43011 (N_43011,N_33401,N_33232);
nor U43012 (N_43012,N_37263,N_39799);
xor U43013 (N_43013,N_30885,N_31639);
or U43014 (N_43014,N_36556,N_39742);
and U43015 (N_43015,N_33392,N_36651);
nor U43016 (N_43016,N_30739,N_36427);
xnor U43017 (N_43017,N_30985,N_36363);
nand U43018 (N_43018,N_39470,N_39821);
nand U43019 (N_43019,N_36643,N_32881);
and U43020 (N_43020,N_36637,N_33005);
nor U43021 (N_43021,N_31140,N_38438);
nand U43022 (N_43022,N_32426,N_32497);
or U43023 (N_43023,N_36622,N_38199);
nand U43024 (N_43024,N_32296,N_36192);
nand U43025 (N_43025,N_30819,N_37954);
or U43026 (N_43026,N_38107,N_30443);
nor U43027 (N_43027,N_37738,N_39506);
nor U43028 (N_43028,N_34596,N_36335);
and U43029 (N_43029,N_37605,N_30528);
nor U43030 (N_43030,N_39283,N_35662);
or U43031 (N_43031,N_33415,N_38302);
nor U43032 (N_43032,N_31648,N_33093);
or U43033 (N_43033,N_37219,N_37611);
or U43034 (N_43034,N_37952,N_30902);
and U43035 (N_43035,N_33157,N_32802);
nand U43036 (N_43036,N_33408,N_39101);
or U43037 (N_43037,N_31766,N_38269);
or U43038 (N_43038,N_34609,N_30301);
nand U43039 (N_43039,N_32643,N_37259);
nand U43040 (N_43040,N_30416,N_36730);
nor U43041 (N_43041,N_36991,N_32154);
nor U43042 (N_43042,N_33306,N_34684);
nand U43043 (N_43043,N_35774,N_35648);
or U43044 (N_43044,N_33918,N_33007);
or U43045 (N_43045,N_35336,N_37998);
xor U43046 (N_43046,N_36026,N_34521);
or U43047 (N_43047,N_37823,N_35089);
nand U43048 (N_43048,N_37802,N_36450);
xor U43049 (N_43049,N_32618,N_32798);
nand U43050 (N_43050,N_34361,N_36458);
xor U43051 (N_43051,N_30429,N_32116);
nor U43052 (N_43052,N_32474,N_35751);
nor U43053 (N_43053,N_36880,N_33031);
nand U43054 (N_43054,N_34940,N_35073);
and U43055 (N_43055,N_35549,N_32718);
nor U43056 (N_43056,N_31428,N_33521);
nand U43057 (N_43057,N_31399,N_32373);
or U43058 (N_43058,N_33988,N_32093);
nand U43059 (N_43059,N_39100,N_38332);
xnor U43060 (N_43060,N_31252,N_39154);
or U43061 (N_43061,N_35367,N_33278);
xor U43062 (N_43062,N_39660,N_37086);
and U43063 (N_43063,N_38186,N_38663);
nand U43064 (N_43064,N_33684,N_34765);
xnor U43065 (N_43065,N_34924,N_31068);
xnor U43066 (N_43066,N_33154,N_38553);
xnor U43067 (N_43067,N_30730,N_34832);
nor U43068 (N_43068,N_33411,N_39133);
and U43069 (N_43069,N_38915,N_33950);
or U43070 (N_43070,N_39123,N_30937);
nand U43071 (N_43071,N_37880,N_39042);
nor U43072 (N_43072,N_36635,N_36092);
or U43073 (N_43073,N_37410,N_36357);
nand U43074 (N_43074,N_39621,N_30409);
xnor U43075 (N_43075,N_30823,N_39026);
and U43076 (N_43076,N_37412,N_34974);
nor U43077 (N_43077,N_32172,N_32776);
xor U43078 (N_43078,N_30433,N_30924);
and U43079 (N_43079,N_30176,N_35829);
nand U43080 (N_43080,N_34595,N_39449);
nor U43081 (N_43081,N_33530,N_30078);
xor U43082 (N_43082,N_35965,N_30809);
xnor U43083 (N_43083,N_36775,N_33536);
and U43084 (N_43084,N_34194,N_39422);
nor U43085 (N_43085,N_36548,N_32500);
or U43086 (N_43086,N_33963,N_33582);
xnor U43087 (N_43087,N_38092,N_31790);
and U43088 (N_43088,N_39512,N_31671);
and U43089 (N_43089,N_32319,N_36715);
and U43090 (N_43090,N_33805,N_35545);
and U43091 (N_43091,N_38728,N_33707);
and U43092 (N_43092,N_30270,N_31510);
or U43093 (N_43093,N_31378,N_30349);
or U43094 (N_43094,N_37947,N_34618);
or U43095 (N_43095,N_32022,N_34264);
nor U43096 (N_43096,N_31305,N_37831);
and U43097 (N_43097,N_30073,N_34459);
xor U43098 (N_43098,N_36416,N_30529);
nor U43099 (N_43099,N_37448,N_37143);
and U43100 (N_43100,N_30797,N_30599);
and U43101 (N_43101,N_32624,N_31017);
nor U43102 (N_43102,N_32084,N_37471);
nor U43103 (N_43103,N_33145,N_33666);
nor U43104 (N_43104,N_35530,N_34835);
or U43105 (N_43105,N_36180,N_31799);
and U43106 (N_43106,N_34214,N_33016);
xnor U43107 (N_43107,N_32773,N_39059);
or U43108 (N_43108,N_32284,N_32774);
nand U43109 (N_43109,N_33122,N_32463);
or U43110 (N_43110,N_33596,N_38034);
and U43111 (N_43111,N_36358,N_34501);
nand U43112 (N_43112,N_32313,N_30395);
or U43113 (N_43113,N_36580,N_30022);
nand U43114 (N_43114,N_39268,N_37288);
and U43115 (N_43115,N_31579,N_35206);
or U43116 (N_43116,N_31083,N_35158);
nand U43117 (N_43117,N_39050,N_32863);
nand U43118 (N_43118,N_32200,N_36905);
xor U43119 (N_43119,N_39599,N_31401);
nor U43120 (N_43120,N_33979,N_35964);
or U43121 (N_43121,N_32715,N_35384);
nor U43122 (N_43122,N_30928,N_34242);
or U43123 (N_43123,N_39527,N_34628);
or U43124 (N_43124,N_36702,N_36701);
nor U43125 (N_43125,N_31366,N_31814);
nand U43126 (N_43126,N_32328,N_39903);
or U43127 (N_43127,N_36218,N_31748);
nand U43128 (N_43128,N_36366,N_35126);
and U43129 (N_43129,N_32145,N_30581);
or U43130 (N_43130,N_36742,N_32800);
and U43131 (N_43131,N_30503,N_38454);
nand U43132 (N_43132,N_38389,N_35473);
nand U43133 (N_43133,N_30560,N_32361);
nor U43134 (N_43134,N_39739,N_38303);
nor U43135 (N_43135,N_31452,N_33036);
nor U43136 (N_43136,N_38602,N_33100);
or U43137 (N_43137,N_38134,N_39055);
and U43138 (N_43138,N_30184,N_37920);
and U43139 (N_43139,N_39465,N_38975);
xor U43140 (N_43140,N_31563,N_36341);
and U43141 (N_43141,N_37903,N_36070);
nor U43142 (N_43142,N_37284,N_39537);
nand U43143 (N_43143,N_37009,N_39344);
nor U43144 (N_43144,N_36656,N_33365);
or U43145 (N_43145,N_35750,N_32440);
nand U43146 (N_43146,N_30510,N_34845);
nand U43147 (N_43147,N_36693,N_36876);
or U43148 (N_43148,N_31833,N_39948);
xnor U43149 (N_43149,N_37466,N_39532);
and U43150 (N_43150,N_32437,N_35901);
nand U43151 (N_43151,N_31879,N_33569);
nand U43152 (N_43152,N_37787,N_34339);
nand U43153 (N_43153,N_36321,N_36834);
nor U43154 (N_43154,N_34724,N_34928);
nand U43155 (N_43155,N_36659,N_35794);
and U43156 (N_43156,N_33824,N_37590);
nor U43157 (N_43157,N_30303,N_33149);
and U43158 (N_43158,N_34945,N_38708);
or U43159 (N_43159,N_37125,N_30748);
or U43160 (N_43160,N_37557,N_32953);
nand U43161 (N_43161,N_32137,N_38792);
and U43162 (N_43162,N_37927,N_31491);
or U43163 (N_43163,N_35528,N_37728);
and U43164 (N_43164,N_31037,N_34927);
nor U43165 (N_43165,N_36290,N_30586);
nand U43166 (N_43166,N_33866,N_30892);
and U43167 (N_43167,N_30218,N_38621);
and U43168 (N_43168,N_33324,N_36039);
nand U43169 (N_43169,N_36360,N_35601);
or U43170 (N_43170,N_39286,N_33911);
xnor U43171 (N_43171,N_34363,N_31537);
and U43172 (N_43172,N_38079,N_31010);
nand U43173 (N_43173,N_36686,N_31934);
and U43174 (N_43174,N_32809,N_37296);
xnor U43175 (N_43175,N_39525,N_36771);
xor U43176 (N_43176,N_37429,N_38530);
xnor U43177 (N_43177,N_38791,N_39683);
and U43178 (N_43178,N_34606,N_32627);
or U43179 (N_43179,N_39054,N_31409);
and U43180 (N_43180,N_39136,N_33179);
or U43181 (N_43181,N_39481,N_36617);
xnor U43182 (N_43182,N_30431,N_39675);
or U43183 (N_43183,N_35770,N_32778);
and U43184 (N_43184,N_30904,N_38365);
or U43185 (N_43185,N_32079,N_35394);
xnor U43186 (N_43186,N_38453,N_39891);
or U43187 (N_43187,N_31408,N_34312);
nand U43188 (N_43188,N_37558,N_32897);
nor U43189 (N_43189,N_31090,N_33794);
or U43190 (N_43190,N_38630,N_36910);
or U43191 (N_43191,N_35200,N_32089);
and U43192 (N_43192,N_35908,N_37133);
and U43193 (N_43193,N_33754,N_31974);
xnor U43194 (N_43194,N_34828,N_31607);
and U43195 (N_43195,N_37573,N_30608);
nand U43196 (N_43196,N_37655,N_34870);
and U43197 (N_43197,N_38487,N_37990);
and U43198 (N_43198,N_35002,N_36949);
and U43199 (N_43199,N_36890,N_35981);
nor U43200 (N_43200,N_35906,N_35440);
nand U43201 (N_43201,N_39545,N_37093);
or U43202 (N_43202,N_34407,N_30527);
and U43203 (N_43203,N_34956,N_30120);
nand U43204 (N_43204,N_35412,N_30724);
nand U43205 (N_43205,N_31232,N_39531);
or U43206 (N_43206,N_33237,N_36491);
and U43207 (N_43207,N_31330,N_39384);
nand U43208 (N_43208,N_31957,N_32455);
nand U43209 (N_43209,N_30806,N_33594);
nand U43210 (N_43210,N_32751,N_30038);
or U43211 (N_43211,N_33816,N_35511);
and U43212 (N_43212,N_32930,N_35222);
nand U43213 (N_43213,N_39323,N_36443);
and U43214 (N_43214,N_39432,N_38110);
or U43215 (N_43215,N_33287,N_31230);
nand U43216 (N_43216,N_36158,N_36198);
nand U43217 (N_43217,N_38813,N_36313);
and U43218 (N_43218,N_31644,N_36471);
nor U43219 (N_43219,N_39159,N_36936);
nor U43220 (N_43220,N_33788,N_32371);
and U43221 (N_43221,N_37893,N_32453);
nor U43222 (N_43222,N_31636,N_36169);
or U43223 (N_43223,N_37019,N_31620);
nand U43224 (N_43224,N_30689,N_34908);
xnor U43225 (N_43225,N_35878,N_34688);
nand U43226 (N_43226,N_33637,N_35834);
and U43227 (N_43227,N_31497,N_33276);
or U43228 (N_43228,N_39879,N_37066);
and U43229 (N_43229,N_39919,N_30168);
xor U43230 (N_43230,N_34795,N_30758);
nand U43231 (N_43231,N_33166,N_36102);
nor U43232 (N_43232,N_36551,N_32372);
nand U43233 (N_43233,N_31269,N_34235);
and U43234 (N_43234,N_38612,N_37181);
xnor U43235 (N_43235,N_36646,N_35865);
nand U43236 (N_43236,N_36952,N_37689);
nand U43237 (N_43237,N_30963,N_37200);
or U43238 (N_43238,N_35792,N_37737);
nor U43239 (N_43239,N_35433,N_34957);
or U43240 (N_43240,N_39365,N_35565);
and U43241 (N_43241,N_34335,N_34321);
or U43242 (N_43242,N_33864,N_38152);
or U43243 (N_43243,N_32428,N_39930);
xor U43244 (N_43244,N_33540,N_32390);
nor U43245 (N_43245,N_38920,N_37630);
or U43246 (N_43246,N_36644,N_33285);
and U43247 (N_43247,N_38004,N_32708);
nor U43248 (N_43248,N_31213,N_33085);
nor U43249 (N_43249,N_39732,N_38163);
and U43250 (N_43250,N_38997,N_35444);
and U43251 (N_43251,N_35654,N_33345);
and U43252 (N_43252,N_39656,N_35177);
xor U43253 (N_43253,N_35101,N_35315);
nand U43254 (N_43254,N_33194,N_33216);
nor U43255 (N_43255,N_33017,N_34677);
xor U43256 (N_43256,N_39536,N_36853);
nand U43257 (N_43257,N_35405,N_39138);
xnor U43258 (N_43258,N_37898,N_38076);
nor U43259 (N_43259,N_33289,N_30606);
nor U43260 (N_43260,N_32263,N_35481);
nor U43261 (N_43261,N_35205,N_36921);
nor U43262 (N_43262,N_33669,N_30280);
nand U43263 (N_43263,N_37442,N_30731);
and U43264 (N_43264,N_39414,N_36970);
and U43265 (N_43265,N_37892,N_34099);
and U43266 (N_43266,N_37515,N_31608);
nand U43267 (N_43267,N_33275,N_31827);
nor U43268 (N_43268,N_35602,N_34668);
and U43269 (N_43269,N_37195,N_34440);
xnor U43270 (N_43270,N_37553,N_34347);
nand U43271 (N_43271,N_31328,N_37373);
nand U43272 (N_43272,N_32279,N_30921);
xor U43273 (N_43273,N_31113,N_31754);
or U43274 (N_43274,N_31591,N_36167);
nand U43275 (N_43275,N_38431,N_38694);
or U43276 (N_43276,N_31920,N_35228);
nand U43277 (N_43277,N_39349,N_35606);
nor U43278 (N_43278,N_31674,N_34930);
nand U43279 (N_43279,N_37057,N_34674);
or U43280 (N_43280,N_32261,N_34496);
and U43281 (N_43281,N_31459,N_36000);
and U43282 (N_43282,N_33826,N_36550);
nand U43283 (N_43283,N_38582,N_39023);
nand U43284 (N_43284,N_30493,N_33688);
and U43285 (N_43285,N_30837,N_32711);
nor U43286 (N_43286,N_38211,N_34738);
and U43287 (N_43287,N_31690,N_31449);
nand U43288 (N_43288,N_36457,N_34919);
nor U43289 (N_43289,N_39752,N_39884);
or U43290 (N_43290,N_32900,N_32781);
nand U43291 (N_43291,N_36255,N_31350);
nor U43292 (N_43292,N_31388,N_38119);
nor U43293 (N_43293,N_33991,N_39457);
nor U43294 (N_43294,N_30662,N_34591);
nor U43295 (N_43295,N_33143,N_39192);
or U43296 (N_43296,N_34445,N_39814);
or U43297 (N_43297,N_37038,N_39120);
and U43298 (N_43298,N_31004,N_31351);
nand U43299 (N_43299,N_34111,N_38077);
or U43300 (N_43300,N_33387,N_38300);
and U43301 (N_43301,N_37663,N_36231);
nor U43302 (N_43302,N_32146,N_31358);
or U43303 (N_43303,N_32043,N_37233);
or U43304 (N_43304,N_37168,N_39716);
nor U43305 (N_43305,N_31785,N_37617);
and U43306 (N_43306,N_36569,N_39572);
nor U43307 (N_43307,N_34874,N_35512);
or U43308 (N_43308,N_36129,N_30603);
or U43309 (N_43309,N_31965,N_36972);
nand U43310 (N_43310,N_36584,N_34091);
nor U43311 (N_43311,N_33679,N_37399);
and U43312 (N_43312,N_37564,N_30788);
nand U43313 (N_43313,N_35671,N_36557);
nor U43314 (N_43314,N_39102,N_31216);
and U43315 (N_43315,N_36385,N_35709);
nand U43316 (N_43316,N_35013,N_31742);
nand U43317 (N_43317,N_32986,N_30911);
nand U43318 (N_43318,N_34413,N_31156);
or U43319 (N_43319,N_31167,N_34128);
or U43320 (N_43320,N_30751,N_33475);
xnor U43321 (N_43321,N_34052,N_39143);
nand U43322 (N_43322,N_39957,N_39392);
xnor U43323 (N_43323,N_36856,N_31100);
or U43324 (N_43324,N_31438,N_32958);
and U43325 (N_43325,N_32789,N_30298);
nand U43326 (N_43326,N_33254,N_34210);
or U43327 (N_43327,N_36263,N_32793);
nor U43328 (N_43328,N_30699,N_34386);
and U43329 (N_43329,N_30833,N_33737);
or U43330 (N_43330,N_32099,N_38525);
nand U43331 (N_43331,N_37684,N_34896);
and U43332 (N_43332,N_33551,N_35178);
nand U43333 (N_43333,N_35669,N_37479);
and U43334 (N_43334,N_36088,N_39784);
and U43335 (N_43335,N_37571,N_31150);
nand U43336 (N_43336,N_38481,N_32291);
nor U43337 (N_43337,N_38475,N_38143);
xor U43338 (N_43338,N_35148,N_35673);
and U43339 (N_43339,N_34205,N_38141);
or U43340 (N_43340,N_35247,N_30010);
nand U43341 (N_43341,N_31018,N_37268);
and U43342 (N_43342,N_36852,N_35289);
nand U43343 (N_43343,N_36768,N_30793);
and U43344 (N_43344,N_30135,N_38041);
xor U43345 (N_43345,N_32378,N_38934);
nor U43346 (N_43346,N_35711,N_33376);
nor U43347 (N_43347,N_32814,N_35066);
nand U43348 (N_43348,N_34612,N_32925);
and U43349 (N_43349,N_30630,N_34552);
nor U43350 (N_43350,N_32447,N_39913);
nand U43351 (N_43351,N_30192,N_38396);
and U43352 (N_43352,N_39266,N_37784);
and U43353 (N_43353,N_33377,N_31919);
nor U43354 (N_43354,N_34085,N_34059);
nor U43355 (N_43355,N_35912,N_34322);
nor U43356 (N_43356,N_39375,N_38415);
and U43357 (N_43357,N_38286,N_36098);
xnor U43358 (N_43358,N_32062,N_30382);
nand U43359 (N_43359,N_37261,N_31295);
nor U43360 (N_43360,N_34597,N_32266);
nand U43361 (N_43361,N_38705,N_39941);
or U43362 (N_43362,N_35861,N_39976);
nor U43363 (N_43363,N_33892,N_33554);
nor U43364 (N_43364,N_34172,N_39321);
and U43365 (N_43365,N_36101,N_31565);
nand U43366 (N_43366,N_30494,N_37609);
nor U43367 (N_43367,N_33552,N_37095);
or U43368 (N_43368,N_30332,N_35559);
nand U43369 (N_43369,N_32155,N_32417);
and U43370 (N_43370,N_37439,N_33797);
nor U43371 (N_43371,N_33052,N_32466);
or U43372 (N_43372,N_36965,N_30163);
or U43373 (N_43373,N_33070,N_38411);
nor U43374 (N_43374,N_39230,N_37275);
nor U43375 (N_43375,N_34147,N_38180);
nand U43376 (N_43376,N_39723,N_37633);
and U43377 (N_43377,N_35257,N_35365);
and U43378 (N_43378,N_32646,N_39587);
or U43379 (N_43379,N_32818,N_39569);
nand U43380 (N_43380,N_39845,N_33200);
nor U43381 (N_43381,N_38741,N_30799);
nor U43382 (N_43382,N_35147,N_38538);
and U43383 (N_43383,N_38686,N_34838);
nand U43384 (N_43384,N_31376,N_32487);
and U43385 (N_43385,N_33625,N_33204);
xnor U43386 (N_43386,N_37183,N_38074);
xnor U43387 (N_43387,N_39312,N_37037);
or U43388 (N_43388,N_35701,N_37671);
nand U43389 (N_43389,N_33121,N_36073);
or U43390 (N_43390,N_36200,N_33344);
nand U43391 (N_43391,N_32166,N_35520);
nor U43392 (N_43392,N_34729,N_32707);
xnor U43393 (N_43393,N_39155,N_38890);
nor U43394 (N_43394,N_34533,N_39316);
nand U43395 (N_43395,N_32060,N_38943);
nand U43396 (N_43396,N_36980,N_32198);
nand U43397 (N_43397,N_35743,N_39868);
xor U43398 (N_43398,N_37185,N_37759);
xor U43399 (N_43399,N_32405,N_30845);
xor U43400 (N_43400,N_32714,N_30438);
or U43401 (N_43401,N_30372,N_37584);
xor U43402 (N_43402,N_36165,N_37343);
and U43403 (N_43403,N_35500,N_33227);
nand U43404 (N_43404,N_33923,N_34748);
nor U43405 (N_43405,N_31544,N_32684);
and U43406 (N_43406,N_36142,N_35889);
xnor U43407 (N_43407,N_30682,N_36072);
nor U43408 (N_43408,N_35442,N_30402);
nor U43409 (N_43409,N_31541,N_37403);
nand U43410 (N_43410,N_32622,N_30951);
nor U43411 (N_43411,N_30756,N_35108);
or U43412 (N_43412,N_31696,N_33662);
nor U43413 (N_43413,N_35312,N_31356);
nand U43414 (N_43414,N_38346,N_37524);
nor U43415 (N_43415,N_37804,N_36553);
and U43416 (N_43416,N_30987,N_37437);
and U43417 (N_43417,N_36251,N_35370);
nand U43418 (N_43418,N_35841,N_30228);
and U43419 (N_43419,N_38938,N_39403);
and U43420 (N_43420,N_30771,N_34663);
or U43421 (N_43421,N_32265,N_32916);
xnor U43422 (N_43422,N_34621,N_38574);
or U43423 (N_43423,N_30486,N_37083);
or U43424 (N_43424,N_38809,N_32127);
and U43425 (N_43425,N_31450,N_30850);
nor U43426 (N_43426,N_32003,N_34762);
nor U43427 (N_43427,N_36368,N_39369);
xor U43428 (N_43428,N_30007,N_35957);
nand U43429 (N_43429,N_32418,N_39333);
and U43430 (N_43430,N_38099,N_30635);
nor U43431 (N_43431,N_38291,N_38422);
and U43432 (N_43432,N_31872,N_36688);
nor U43433 (N_43433,N_36629,N_35931);
or U43434 (N_43434,N_39109,N_39577);
nand U43435 (N_43435,N_31011,N_36086);
or U43436 (N_43436,N_39972,N_31628);
nor U43437 (N_43437,N_37329,N_32740);
nor U43438 (N_43438,N_32572,N_34598);
nand U43439 (N_43439,N_31984,N_34437);
or U43440 (N_43440,N_34705,N_34399);
nor U43441 (N_43441,N_38996,N_30201);
and U43442 (N_43442,N_36191,N_37744);
nand U43443 (N_43443,N_32159,N_36138);
nand U43444 (N_43444,N_32892,N_37062);
nor U43445 (N_43445,N_37405,N_33400);
or U43446 (N_43446,N_39598,N_30905);
nand U43447 (N_43447,N_31208,N_37860);
and U43448 (N_43448,N_35571,N_34241);
or U43449 (N_43449,N_36014,N_34134);
xor U43450 (N_43450,N_39510,N_32380);
or U43451 (N_43451,N_33839,N_36187);
and U43452 (N_43452,N_32370,N_34283);
nor U43453 (N_43453,N_32716,N_30959);
nor U43454 (N_43454,N_31745,N_38718);
nand U43455 (N_43455,N_35623,N_34572);
and U43456 (N_43456,N_31533,N_35786);
nor U43457 (N_43457,N_32954,N_36942);
nand U43458 (N_43458,N_36640,N_34268);
or U43459 (N_43459,N_34527,N_38011);
and U43460 (N_43460,N_32765,N_33299);
nor U43461 (N_43461,N_34961,N_37853);
or U43462 (N_43462,N_31538,N_30173);
nor U43463 (N_43463,N_37465,N_31853);
nor U43464 (N_43464,N_32567,N_34410);
nor U43465 (N_43465,N_38502,N_39085);
or U43466 (N_43466,N_38595,N_31095);
nor U43467 (N_43467,N_35649,N_33645);
and U43468 (N_43468,N_38430,N_39681);
or U43469 (N_43469,N_31126,N_38374);
nor U43470 (N_43470,N_38082,N_39643);
or U43471 (N_43471,N_34308,N_38820);
and U43472 (N_43472,N_32616,N_33880);
and U43473 (N_43473,N_39542,N_38067);
nand U43474 (N_43474,N_35084,N_37961);
nor U43475 (N_43475,N_32139,N_30387);
nand U43476 (N_43476,N_33404,N_39010);
nand U43477 (N_43477,N_39615,N_35234);
nand U43478 (N_43478,N_33010,N_36790);
and U43479 (N_43479,N_33029,N_34581);
and U43480 (N_43480,N_39476,N_38534);
and U43481 (N_43481,N_33636,N_33888);
and U43482 (N_43482,N_31492,N_31517);
nor U43483 (N_43483,N_36841,N_32424);
xnor U43484 (N_43484,N_32981,N_36685);
or U43485 (N_43485,N_30027,N_35725);
or U43486 (N_43486,N_30884,N_34610);
and U43487 (N_43487,N_32002,N_36499);
or U43488 (N_43488,N_33333,N_30713);
nor U43489 (N_43489,N_37693,N_33437);
and U43490 (N_43490,N_37061,N_33641);
xnor U43491 (N_43491,N_35298,N_34331);
nand U43492 (N_43492,N_39472,N_35745);
xor U43493 (N_43493,N_35001,N_38260);
or U43494 (N_43494,N_36519,N_37114);
nand U43495 (N_43495,N_39939,N_36206);
and U43496 (N_43496,N_35737,N_39612);
and U43497 (N_43497,N_37938,N_33820);
nor U43498 (N_43498,N_34655,N_33247);
nor U43499 (N_43499,N_38631,N_38115);
and U43500 (N_43500,N_39873,N_34964);
nand U43501 (N_43501,N_33522,N_34702);
and U43502 (N_43502,N_30803,N_34558);
and U43503 (N_43503,N_32679,N_33323);
nor U43504 (N_43504,N_34652,N_30081);
and U43505 (N_43505,N_34249,N_30825);
and U43506 (N_43506,N_30513,N_36710);
and U43507 (N_43507,N_35839,N_32857);
or U43508 (N_43508,N_36421,N_38921);
and U43509 (N_43509,N_32948,N_34429);
nor U43510 (N_43510,N_33270,N_32575);
and U43511 (N_43511,N_33246,N_37909);
and U43512 (N_43512,N_32038,N_36265);
and U43513 (N_43513,N_31340,N_38405);
nor U43514 (N_43514,N_32901,N_36517);
and U43515 (N_43515,N_30584,N_38205);
and U43516 (N_43516,N_34986,N_30351);
and U43517 (N_43517,N_30062,N_39604);
and U43518 (N_43518,N_36273,N_34539);
nand U43519 (N_43519,N_33046,N_38633);
or U43520 (N_43520,N_34067,N_36558);
or U43521 (N_43521,N_33391,N_34074);
xor U43522 (N_43522,N_37177,N_33994);
nand U43523 (N_43523,N_34970,N_31668);
nor U43524 (N_43524,N_32513,N_30245);
and U43525 (N_43525,N_36485,N_34948);
and U43526 (N_43526,N_34758,N_32464);
xor U43527 (N_43527,N_34910,N_33954);
and U43528 (N_43528,N_30333,N_32144);
or U43529 (N_43529,N_34710,N_32059);
or U43530 (N_43530,N_35729,N_36667);
and U43531 (N_43531,N_38928,N_36029);
or U43532 (N_43532,N_35997,N_39322);
xnor U43533 (N_43533,N_36571,N_33340);
xnor U43534 (N_43534,N_33351,N_32737);
or U43535 (N_43535,N_39176,N_33877);
and U43536 (N_43536,N_34039,N_39892);
and U43537 (N_43537,N_37310,N_32236);
or U43538 (N_43538,N_32839,N_32336);
or U43539 (N_43539,N_38086,N_31089);
or U43540 (N_43540,N_39345,N_36016);
and U43541 (N_43541,N_31005,N_32914);
nand U43542 (N_43542,N_31254,N_30974);
nand U43543 (N_43543,N_32547,N_32692);
or U43544 (N_43544,N_34695,N_38964);
or U43545 (N_43545,N_34839,N_34092);
or U43546 (N_43546,N_34892,N_35655);
xnor U43547 (N_43547,N_31941,N_31121);
or U43548 (N_43548,N_30294,N_35531);
and U43549 (N_43549,N_37560,N_34358);
nand U43550 (N_43550,N_37978,N_35262);
nand U43551 (N_43551,N_35254,N_31552);
nand U43552 (N_43552,N_37031,N_38337);
nand U43553 (N_43553,N_36821,N_34735);
or U43554 (N_43554,N_37203,N_32386);
nand U43555 (N_43555,N_37144,N_34430);
and U43556 (N_43556,N_35551,N_32736);
and U43557 (N_43557,N_30914,N_39477);
nand U43558 (N_43558,N_35970,N_34510);
nand U43559 (N_43559,N_38516,N_31009);
and U43560 (N_43560,N_37356,N_36372);
or U43561 (N_43561,N_30305,N_38213);
or U43562 (N_43562,N_36879,N_34353);
nor U43563 (N_43563,N_31082,N_37851);
nand U43564 (N_43564,N_36063,N_33373);
xnor U43565 (N_43565,N_30098,N_34542);
xnor U43566 (N_43566,N_35424,N_33760);
and U43567 (N_43567,N_33858,N_38810);
nor U43568 (N_43568,N_36193,N_37600);
nor U43569 (N_43569,N_36134,N_36350);
nand U43570 (N_43570,N_39482,N_36589);
nor U43571 (N_43571,N_38083,N_35664);
xor U43572 (N_43572,N_31119,N_33500);
nand U43573 (N_43573,N_31429,N_32845);
and U43574 (N_43574,N_33631,N_36819);
nand U43575 (N_43575,N_35844,N_31952);
nor U43576 (N_43576,N_38987,N_32920);
or U43577 (N_43577,N_35710,N_39444);
nand U43578 (N_43578,N_36850,N_30054);
or U43579 (N_43579,N_35223,N_34901);
xor U43580 (N_43580,N_39073,N_36788);
xnor U43581 (N_43581,N_34624,N_39526);
nor U43582 (N_43582,N_35064,N_32927);
and U43583 (N_43583,N_32216,N_30596);
and U43584 (N_43584,N_39399,N_32577);
xnor U43585 (N_43585,N_30069,N_32224);
nand U43586 (N_43586,N_37174,N_39824);
nor U43587 (N_43587,N_34452,N_30505);
nand U43588 (N_43588,N_37255,N_37889);
and U43589 (N_43589,N_35489,N_38484);
nor U43590 (N_43590,N_30634,N_36504);
nor U43591 (N_43591,N_36245,N_34461);
or U43592 (N_43592,N_37933,N_39118);
or U43593 (N_43593,N_32796,N_37740);
and U43594 (N_43594,N_34830,N_31614);
nand U43595 (N_43595,N_38373,N_32856);
or U43596 (N_43596,N_30157,N_31812);
or U43597 (N_43597,N_39448,N_32889);
nand U43598 (N_43598,N_34287,N_37583);
xnor U43599 (N_43599,N_30654,N_33170);
or U43600 (N_43600,N_30459,N_32997);
nand U43601 (N_43601,N_32000,N_38859);
nand U43602 (N_43602,N_34146,N_38945);
nand U43603 (N_43603,N_33539,N_32558);
nand U43604 (N_43604,N_38870,N_35182);
nand U43605 (N_43605,N_38262,N_31255);
or U43606 (N_43606,N_30174,N_32855);
or U43607 (N_43607,N_36043,N_31691);
nor U43608 (N_43608,N_35023,N_33315);
or U43609 (N_43609,N_34269,N_34467);
and U43610 (N_43610,N_32696,N_30379);
nor U43611 (N_43611,N_32742,N_36369);
xor U43612 (N_43612,N_30623,N_36173);
nor U43613 (N_43613,N_31867,N_39801);
nor U43614 (N_43614,N_31946,N_39982);
nor U43615 (N_43615,N_35415,N_38007);
nor U43616 (N_43616,N_30103,N_37234);
nand U43617 (N_43617,N_33806,N_34104);
and U43618 (N_43618,N_39376,N_32321);
or U43619 (N_43619,N_38635,N_39647);
and U43620 (N_43620,N_30352,N_35988);
and U43621 (N_43621,N_31769,N_36148);
and U43622 (N_43622,N_33941,N_31765);
or U43623 (N_43623,N_34619,N_30842);
and U43624 (N_43624,N_34638,N_38197);
nor U43625 (N_43625,N_34804,N_37182);
nor U43626 (N_43626,N_36096,N_37077);
nor U43627 (N_43627,N_35324,N_34288);
nand U43628 (N_43628,N_35000,N_33372);
nor U43629 (N_43629,N_30247,N_33985);
nand U43630 (N_43630,N_38895,N_37451);
nor U43631 (N_43631,N_37614,N_31811);
or U43632 (N_43632,N_34355,N_33487);
and U43633 (N_43633,N_32177,N_38016);
or U43634 (N_43634,N_32078,N_39494);
and U43635 (N_43635,N_32788,N_30037);
or U43636 (N_43636,N_36492,N_30582);
and U43637 (N_43637,N_32221,N_32014);
or U43638 (N_43638,N_32686,N_32860);
xnor U43639 (N_43639,N_31106,N_33322);
nor U43640 (N_43640,N_35072,N_33652);
and U43641 (N_43641,N_34566,N_31503);
or U43642 (N_43642,N_37829,N_39756);
or U43643 (N_43643,N_30359,N_38387);
or U43644 (N_43644,N_36153,N_37528);
or U43645 (N_43645,N_38714,N_32658);
nor U43646 (N_43646,N_39673,N_38145);
nand U43647 (N_43647,N_38786,N_38312);
or U43648 (N_43648,N_36515,N_38080);
nor U43649 (N_43649,N_31572,N_35395);
nand U43650 (N_43650,N_36137,N_34173);
nor U43651 (N_43651,N_32830,N_36521);
and U43652 (N_43652,N_33623,N_31504);
nor U43653 (N_43653,N_31266,N_30121);
nor U43654 (N_43654,N_31643,N_32753);
or U43655 (N_43655,N_34730,N_38289);
and U43656 (N_43656,N_38537,N_37788);
nor U43657 (N_43657,N_36338,N_32582);
nand U43658 (N_43658,N_34617,N_33102);
nand U43659 (N_43659,N_32092,N_35566);
nand U43660 (N_43660,N_32340,N_34101);
and U43661 (N_43661,N_31446,N_30477);
nor U43662 (N_43662,N_31551,N_38935);
and U43663 (N_43663,N_33146,N_33018);
nand U43664 (N_43664,N_30050,N_33563);
or U43665 (N_43665,N_33268,N_36816);
or U43666 (N_43666,N_37819,N_32120);
or U43667 (N_43667,N_34719,N_33715);
nor U43668 (N_43668,N_34168,N_34865);
nand U43669 (N_43669,N_33681,N_31054);
and U43670 (N_43670,N_37287,N_35812);
and U43671 (N_43671,N_38885,N_33907);
or U43672 (N_43672,N_38246,N_30232);
and U43673 (N_43673,N_35213,N_32933);
or U43674 (N_43674,N_31339,N_37795);
and U43675 (N_43675,N_35636,N_39125);
and U43676 (N_43676,N_32748,N_39178);
or U43677 (N_43677,N_38385,N_31848);
nor U43678 (N_43678,N_32115,N_33583);
nor U43679 (N_43679,N_37988,N_34949);
nand U43680 (N_43680,N_36170,N_36971);
or U43681 (N_43681,N_30114,N_32755);
and U43682 (N_43682,N_32278,N_32583);
nand U43683 (N_43683,N_32811,N_33111);
and U43684 (N_43684,N_30685,N_37871);
and U43685 (N_43685,N_39174,N_37467);
nor U43686 (N_43686,N_35846,N_38361);
and U43687 (N_43687,N_39738,N_34032);
nor U43688 (N_43688,N_39126,N_35281);
or U43689 (N_43689,N_31880,N_39763);
and U43690 (N_43690,N_33298,N_32211);
and U43691 (N_43691,N_34941,N_38399);
and U43692 (N_43692,N_36541,N_36963);
or U43693 (N_43693,N_32020,N_34426);
and U43694 (N_43694,N_30763,N_31471);
nor U43695 (N_43695,N_35303,N_30759);
nor U43696 (N_43696,N_30990,N_31558);
nor U43697 (N_43697,N_38738,N_35009);
or U43698 (N_43698,N_35248,N_30597);
or U43699 (N_43699,N_38833,N_37543);
or U43700 (N_43700,N_35672,N_39066);
nand U43701 (N_43701,N_38051,N_32131);
and U43702 (N_43702,N_33264,N_30643);
nor U43703 (N_43703,N_33675,N_38065);
or U43704 (N_43704,N_38335,N_31757);
and U43705 (N_43705,N_35535,N_32304);
nand U43706 (N_43706,N_34004,N_36513);
or U43707 (N_43707,N_37413,N_34632);
nand U43708 (N_43708,N_35806,N_39934);
nand U43709 (N_43709,N_33937,N_38472);
nand U43710 (N_43710,N_33687,N_33416);
or U43711 (N_43711,N_35967,N_35476);
and U43712 (N_43712,N_35740,N_34306);
nand U43713 (N_43713,N_35938,N_32548);
or U43714 (N_43714,N_34129,N_38628);
xnor U43715 (N_43715,N_39725,N_38104);
nor U43716 (N_43716,N_31646,N_30089);
nand U43717 (N_43717,N_37282,N_32275);
and U43718 (N_43718,N_31858,N_39541);
xor U43719 (N_43719,N_34070,N_32305);
nand U43720 (N_43720,N_31849,N_31120);
or U43721 (N_43721,N_33471,N_35286);
or U43722 (N_43722,N_39025,N_38093);
nor U43723 (N_43723,N_38713,N_37126);
nor U43724 (N_43724,N_34476,N_37097);
nor U43725 (N_43725,N_32176,N_31172);
and U43726 (N_43726,N_33283,N_36230);
nor U43727 (N_43727,N_33019,N_34593);
and U43728 (N_43728,N_38818,N_33353);
and U43729 (N_43729,N_35453,N_36610);
nand U43730 (N_43730,N_30145,N_39998);
and U43731 (N_43731,N_36510,N_37928);
and U43732 (N_43732,N_37967,N_38433);
xor U43733 (N_43733,N_37585,N_33390);
nand U43734 (N_43734,N_35984,N_38539);
or U43735 (N_43735,N_30426,N_34113);
nand U43736 (N_43736,N_34383,N_38263);
and U43737 (N_43737,N_30600,N_37857);
nand U43738 (N_43738,N_32163,N_32393);
and U43739 (N_43739,N_39535,N_30231);
and U43740 (N_43740,N_32600,N_34281);
or U43741 (N_43741,N_38106,N_37814);
nor U43742 (N_43742,N_33700,N_33577);
or U43743 (N_43743,N_35410,N_30773);
nor U43744 (N_43744,N_36744,N_34540);
nand U43745 (N_43745,N_34267,N_30591);
and U43746 (N_43746,N_36463,N_35404);
or U43747 (N_43747,N_32951,N_37724);
nor U43748 (N_43748,N_30342,N_36159);
nand U43749 (N_43749,N_35110,N_37147);
nand U43750 (N_43750,N_34359,N_39697);
nor U43751 (N_43751,N_34818,N_31153);
nand U43752 (N_43752,N_36112,N_35359);
and U43753 (N_43753,N_31183,N_33724);
or U43754 (N_43754,N_32241,N_30831);
and U43755 (N_43755,N_37438,N_31372);
or U43756 (N_43756,N_31263,N_32644);
nor U43757 (N_43757,N_38319,N_38898);
and U43758 (N_43758,N_31074,N_35419);
nand U43759 (N_43759,N_39816,N_37747);
and U43760 (N_43760,N_32392,N_37426);
nand U43761 (N_43761,N_32123,N_38661);
nand U43762 (N_43762,N_33860,N_34221);
nand U43763 (N_43763,N_37768,N_36196);
nand U43764 (N_43764,N_33035,N_31819);
nor U43765 (N_43765,N_37187,N_32819);
and U43766 (N_43766,N_31928,N_31838);
nand U43767 (N_43767,N_32555,N_33856);
nand U43768 (N_43768,N_35870,N_35887);
nand U43769 (N_43769,N_37797,N_38425);
or U43770 (N_43770,N_31035,N_38717);
and U43771 (N_43771,N_36032,N_35168);
nor U43772 (N_43772,N_35757,N_37096);
nand U43773 (N_43773,N_36954,N_33223);
or U43774 (N_43774,N_33022,N_35221);
nor U43775 (N_43775,N_39530,N_31353);
or U43776 (N_43776,N_36691,N_35038);
nor U43777 (N_43777,N_33810,N_38567);
nor U43778 (N_43778,N_38130,N_35946);
or U43779 (N_43779,N_37188,N_31720);
and U43780 (N_43780,N_35731,N_31513);
and U43781 (N_43781,N_38046,N_31978);
or U43782 (N_43782,N_30864,N_30263);
nor U43783 (N_43783,N_36184,N_34333);
nand U43784 (N_43784,N_37430,N_38094);
and U43785 (N_43785,N_39191,N_30947);
and U43786 (N_43786,N_32215,N_36961);
nor U43787 (N_43787,N_30879,N_31476);
nand U43788 (N_43788,N_30929,N_31192);
or U43789 (N_43789,N_31413,N_35613);
and U43790 (N_43790,N_34079,N_39478);
nor U43791 (N_43791,N_35626,N_35486);
and U43792 (N_43792,N_39515,N_36955);
nor U43793 (N_43793,N_34592,N_30692);
xor U43794 (N_43794,N_38645,N_30474);
and U43795 (N_43795,N_30720,N_39929);
or U43796 (N_43796,N_32580,N_36034);
xor U43797 (N_43797,N_39141,N_32503);
nand U43798 (N_43798,N_31567,N_38391);
nor U43799 (N_43799,N_32024,N_36888);
and U43800 (N_43800,N_31881,N_30093);
or U43801 (N_43801,N_34766,N_31218);
and U43802 (N_43802,N_30626,N_31483);
nor U43803 (N_43803,N_30694,N_31525);
and U43804 (N_43804,N_35352,N_32151);
nor U43805 (N_43805,N_30014,N_30808);
or U43806 (N_43806,N_36162,N_38212);
and U43807 (N_43807,N_34156,N_33638);
nor U43808 (N_43808,N_35800,N_37141);
nor U43809 (N_43809,N_35479,N_31466);
and U43810 (N_43810,N_34298,N_34996);
and U43811 (N_43811,N_34486,N_38268);
and U43812 (N_43812,N_31222,N_35517);
or U43813 (N_43813,N_30012,N_36532);
or U43814 (N_43814,N_34190,N_31703);
nor U43815 (N_43815,N_38643,N_38752);
and U43816 (N_43816,N_30525,N_34614);
or U43817 (N_43817,N_35903,N_37646);
nor U43818 (N_43818,N_38435,N_32230);
and U43819 (N_43819,N_39225,N_35593);
xor U43820 (N_43820,N_30418,N_33833);
nor U43821 (N_43821,N_31191,N_31970);
nor U43822 (N_43822,N_33191,N_37161);
or U43823 (N_43823,N_39093,N_39862);
xor U43824 (N_43824,N_30193,N_34686);
and U43825 (N_43825,N_31505,N_31945);
nand U43826 (N_43826,N_38840,N_31132);
nand U43827 (N_43827,N_36740,N_36219);
nor U43828 (N_43828,N_36592,N_35873);
or U43829 (N_43829,N_32124,N_30293);
or U43830 (N_43830,N_35049,N_34255);
or U43831 (N_43831,N_31234,N_35958);
and U43832 (N_43832,N_30026,N_38583);
or U43833 (N_43833,N_30478,N_31164);
or U43834 (N_43834,N_31577,N_39232);
nor U43835 (N_43835,N_34027,N_36058);
nor U43836 (N_43836,N_36720,N_38965);
nor U43837 (N_43837,N_30129,N_35982);
nor U43838 (N_43838,N_36593,N_30327);
nand U43839 (N_43839,N_38985,N_30705);
or U43840 (N_43840,N_35155,N_36711);
nor U43841 (N_43841,N_39896,N_31454);
and U43842 (N_43842,N_35789,N_37865);
nand U43843 (N_43843,N_37533,N_34669);
nand U43844 (N_43844,N_30675,N_39980);
xor U43845 (N_43845,N_38151,N_38954);
nor U43846 (N_43846,N_39513,N_37917);
xnor U43847 (N_43847,N_31921,N_38096);
and U43848 (N_43848,N_36692,N_33096);
nor U43849 (N_43849,N_31670,N_33325);
nand U43850 (N_43850,N_38710,N_37010);
nor U43851 (N_43851,N_39668,N_32376);
or U43852 (N_43852,N_36282,N_31027);
nand U43853 (N_43853,N_37045,N_35267);
nand U43854 (N_43854,N_39256,N_38459);
xnor U43855 (N_43855,N_33763,N_30090);
and U43856 (N_43856,N_33304,N_36631);
or U43857 (N_43857,N_34380,N_39334);
nand U43858 (N_43858,N_32827,N_34980);
xor U43859 (N_43859,N_33878,N_30645);
nor U43860 (N_43860,N_31828,N_36944);
and U43861 (N_43861,N_31629,N_30136);
nor U43862 (N_43862,N_38644,N_31034);
nor U43863 (N_43863,N_31158,N_35985);
or U43864 (N_43864,N_34503,N_38594);
or U43865 (N_43865,N_39434,N_31791);
or U43866 (N_43866,N_37298,N_35533);
nor U43867 (N_43867,N_30357,N_32587);
xor U43868 (N_43868,N_33410,N_36269);
or U43869 (N_43869,N_31755,N_39691);
nor U43870 (N_43870,N_37325,N_31261);
xor U43871 (N_43871,N_39893,N_35502);
nand U43872 (N_43872,N_37239,N_31631);
and U43873 (N_43873,N_38406,N_36087);
and U43874 (N_43874,N_30223,N_35741);
nor U43875 (N_43875,N_34814,N_30663);
nand U43876 (N_43876,N_30230,N_35048);
and U43877 (N_43877,N_33746,N_31369);
nand U43878 (N_43878,N_32012,N_31227);
nand U43879 (N_43879,N_32368,N_32045);
and U43880 (N_43880,N_36990,N_33151);
and U43881 (N_43881,N_32347,N_35393);
and U43882 (N_43882,N_33062,N_31550);
and U43883 (N_43883,N_39702,N_34844);
and U43884 (N_43884,N_37695,N_38540);
or U43885 (N_43885,N_34270,N_39381);
xor U43886 (N_43886,N_33379,N_35464);
and U43887 (N_43887,N_30786,N_31402);
nand U43888 (N_43888,N_39553,N_37876);
or U43889 (N_43889,N_31528,N_39818);
and U43890 (N_43890,N_36565,N_30926);
and U43891 (N_43891,N_33198,N_34546);
xnor U43892 (N_43892,N_30107,N_38173);
nor U43893 (N_43893,N_38577,N_32104);
or U43894 (N_43894,N_33837,N_30585);
nor U43895 (N_43895,N_32967,N_31841);
or U43896 (N_43896,N_33804,N_34556);
nand U43897 (N_43897,N_39620,N_32339);
or U43898 (N_43898,N_38088,N_31632);
xnor U43899 (N_43899,N_34819,N_34992);
or U43900 (N_43900,N_36743,N_36093);
nor U43901 (N_43901,N_33107,N_34966);
nand U43902 (N_43902,N_35156,N_34233);
nor U43903 (N_43903,N_31699,N_31197);
or U43904 (N_43904,N_34803,N_39754);
or U43905 (N_43905,N_34689,N_34018);
or U43906 (N_43906,N_35345,N_38494);
or U43907 (N_43907,N_30544,N_37879);
nor U43908 (N_43908,N_36621,N_34853);
or U43909 (N_43909,N_34096,N_38683);
nand U43910 (N_43910,N_34831,N_37018);
and U43911 (N_43911,N_34530,N_37422);
and U43912 (N_43912,N_31619,N_39921);
nand U43913 (N_43913,N_38802,N_30423);
nor U43914 (N_43914,N_32561,N_30679);
and U43915 (N_43915,N_34978,N_36975);
nor U43916 (N_43916,N_36734,N_35857);
nand U43917 (N_43917,N_39768,N_36989);
xor U43918 (N_43918,N_35980,N_37974);
xor U43919 (N_43919,N_33378,N_35220);
nor U43920 (N_43920,N_34537,N_32592);
nand U43921 (N_43921,N_38835,N_39145);
nor U43922 (N_43922,N_31522,N_38251);
and U43923 (N_43923,N_39624,N_31432);
xor U43924 (N_43924,N_38234,N_39626);
nor U43925 (N_43925,N_32476,N_31746);
or U43926 (N_43926,N_35095,N_30742);
xnor U43927 (N_43927,N_31136,N_38873);
nand U43928 (N_43928,N_31688,N_36509);
nor U43929 (N_43929,N_39911,N_34364);
nor U43930 (N_43930,N_38811,N_35646);
xnor U43931 (N_43931,N_34883,N_39380);
nor U43932 (N_43932,N_37276,N_35868);
or U43933 (N_43933,N_34726,N_32419);
nor U43934 (N_43934,N_36855,N_38575);
nand U43935 (N_43935,N_30432,N_39110);
nand U43936 (N_43936,N_31304,N_38551);
and U43937 (N_43937,N_37607,N_38191);
nand U43938 (N_43938,N_35748,N_34365);
nand U43939 (N_43939,N_37869,N_31022);
nand U43940 (N_43940,N_37958,N_37396);
or U43941 (N_43941,N_37785,N_37840);
xnor U43942 (N_43942,N_33484,N_37211);
and U43943 (N_43943,N_33020,N_33846);
or U43944 (N_43944,N_38066,N_35044);
or U43945 (N_43945,N_37248,N_30646);
or U43946 (N_43946,N_39405,N_34900);
or U43947 (N_43947,N_33653,N_33473);
nor U43948 (N_43948,N_35358,N_31455);
and U43949 (N_43949,N_39391,N_30322);
and U43950 (N_43950,N_38287,N_32517);
nand U43951 (N_43951,N_36800,N_32364);
nor U43952 (N_43952,N_30613,N_38504);
nor U43953 (N_43953,N_33649,N_37884);
and U43954 (N_43954,N_39781,N_38259);
and U43955 (N_43955,N_35209,N_35522);
or U43956 (N_43956,N_32281,N_34982);
nor U43957 (N_43957,N_35694,N_35204);
nand U43958 (N_43958,N_38114,N_37899);
nand U43959 (N_43959,N_36945,N_37703);
and U43960 (N_43960,N_30077,N_37791);
xnor U43961 (N_43961,N_35369,N_33360);
or U43962 (N_43962,N_33144,N_37244);
nand U43963 (N_43963,N_37997,N_37968);
xor U43964 (N_43964,N_35105,N_30414);
and U43965 (N_43965,N_39704,N_31531);
nor U43966 (N_43966,N_35703,N_33648);
nor U43967 (N_43967,N_37508,N_32912);
nand U43968 (N_43968,N_37801,N_35211);
and U43969 (N_43969,N_37225,N_36123);
and U43970 (N_43970,N_35270,N_30822);
or U43971 (N_43971,N_32312,N_32293);
and U43972 (N_43972,N_32893,N_33600);
nor U43973 (N_43973,N_37157,N_36083);
and U43974 (N_43974,N_31343,N_38947);
and U43975 (N_43975,N_32171,N_37397);
nor U43976 (N_43976,N_31839,N_31808);
and U43977 (N_43977,N_36912,N_34012);
or U43978 (N_43978,N_37680,N_33678);
nor U43979 (N_43979,N_31753,N_32545);
and U43980 (N_43980,N_38166,N_31093);
or U43981 (N_43981,N_33514,N_32288);
and U43982 (N_43982,N_35825,N_31840);
and U43983 (N_43983,N_38918,N_30314);
xor U43984 (N_43984,N_31871,N_35582);
and U43985 (N_43985,N_35773,N_31860);
nand U43986 (N_43986,N_34642,N_35628);
and U43987 (N_43987,N_39802,N_35340);
and U43988 (N_43988,N_31807,N_37068);
nor U43989 (N_43989,N_35700,N_31383);
nand U43990 (N_43990,N_37269,N_35128);
and U43991 (N_43991,N_33527,N_34449);
nor U43992 (N_43992,N_39062,N_38398);
nor U43993 (N_43993,N_35951,N_34094);
and U43994 (N_43994,N_37672,N_35122);
xor U43995 (N_43995,N_34279,N_39846);
nand U43996 (N_43996,N_30002,N_34120);
and U43997 (N_43997,N_30399,N_36946);
xor U43998 (N_43998,N_32705,N_30604);
and U43999 (N_43999,N_35063,N_33925);
nand U44000 (N_44000,N_36334,N_31475);
and U44001 (N_44001,N_39310,N_38232);
nor U44002 (N_44002,N_39699,N_31405);
nor U44003 (N_44003,N_35311,N_39632);
or U44004 (N_44004,N_38132,N_36953);
nor U44005 (N_44005,N_31174,N_30465);
nor U44006 (N_44006,N_33537,N_36735);
nor U44007 (N_44007,N_31711,N_31188);
nand U44008 (N_44008,N_38386,N_32960);
and U44009 (N_44009,N_36894,N_38842);
and U44010 (N_44010,N_31055,N_38069);
or U44011 (N_44011,N_30144,N_36940);
and U44012 (N_44012,N_31923,N_36712);
nand U44013 (N_44013,N_30134,N_37359);
and U44014 (N_44014,N_30105,N_33665);
and U44015 (N_44015,N_30820,N_34649);
xor U44016 (N_44016,N_33543,N_39331);
nand U44017 (N_44017,N_37012,N_30104);
and U44018 (N_44018,N_32990,N_39761);
nor U44019 (N_44019,N_38172,N_31986);
or U44020 (N_44020,N_36310,N_32599);
nand U44021 (N_44021,N_35913,N_39122);
or U44022 (N_44022,N_36473,N_32573);
xor U44023 (N_44023,N_36288,N_33089);
xnor U44024 (N_44024,N_30595,N_33438);
nand U44025 (N_44025,N_37566,N_36333);
and U44026 (N_44026,N_34423,N_37959);
nor U44027 (N_44027,N_34097,N_36140);
and U44028 (N_44028,N_36866,N_39614);
and U44029 (N_44029,N_30463,N_39186);
or U44030 (N_44030,N_38651,N_34220);
or U44031 (N_44031,N_30710,N_35160);
nand U44032 (N_44032,N_32066,N_39111);
or U44033 (N_44033,N_34953,N_36754);
nor U44034 (N_44034,N_32077,N_32080);
nor U44035 (N_44035,N_39114,N_33997);
nand U44036 (N_44036,N_31894,N_33262);
nand U44037 (N_44037,N_36084,N_39106);
nand U44038 (N_44038,N_31124,N_34660);
nor U44039 (N_44039,N_35197,N_38843);
nand U44040 (N_44040,N_36863,N_34118);
or U44041 (N_44041,N_37194,N_36537);
nand U44042 (N_44042,N_30932,N_33362);
or U44043 (N_44043,N_35060,N_32976);
or U44044 (N_44044,N_39961,N_39534);
and U44045 (N_44045,N_34006,N_38460);
nand U44046 (N_44046,N_30936,N_35588);
nand U44047 (N_44047,N_33832,N_35609);
nor U44048 (N_44048,N_32891,N_30029);
nand U44049 (N_44049,N_38318,N_39912);
and U44050 (N_44050,N_30755,N_38778);
or U44051 (N_44051,N_35493,N_33233);
or U44052 (N_44052,N_30380,N_36351);
and U44053 (N_44053,N_39563,N_38565);
or U44054 (N_44054,N_30180,N_33447);
nand U44055 (N_44055,N_38368,N_38907);
nand U44056 (N_44056,N_32988,N_31829);
xnor U44057 (N_44057,N_38546,N_31146);
nand U44058 (N_44058,N_33220,N_35471);
or U44059 (N_44059,N_31581,N_34102);
or U44060 (N_44060,N_31250,N_33942);
or U44061 (N_44061,N_31224,N_39433);
or U44062 (N_44062,N_37620,N_31195);
and U44063 (N_44063,N_38940,N_34041);
nand U44064 (N_44064,N_35491,N_39431);
or U44065 (N_44065,N_34499,N_36581);
and U44066 (N_44066,N_34223,N_36956);
and U44067 (N_44067,N_35474,N_31215);
nor U44068 (N_44068,N_35208,N_32134);
and U44069 (N_44069,N_33840,N_35004);
or U44070 (N_44070,N_32628,N_31029);
and U44071 (N_44071,N_34834,N_35942);
nand U44072 (N_44072,N_39917,N_32568);
nor U44073 (N_44073,N_36934,N_38100);
nor U44074 (N_44074,N_35330,N_34398);
xnor U44075 (N_44075,N_37956,N_30445);
nor U44076 (N_44076,N_30631,N_31831);
nor U44077 (N_44077,N_36561,N_32101);
and U44078 (N_44078,N_34751,N_39978);
and U44079 (N_44079,N_31534,N_32700);
nand U44080 (N_44080,N_30762,N_34029);
or U44081 (N_44081,N_30113,N_33701);
nor U44082 (N_44082,N_31960,N_38931);
xor U44083 (N_44083,N_36418,N_33891);
or U44084 (N_44084,N_33163,N_39751);
nor U44085 (N_44085,N_39222,N_30112);
nor U44086 (N_44086,N_38941,N_33630);
and U44087 (N_44087,N_33874,N_38105);
or U44088 (N_44088,N_34436,N_30095);
and U44089 (N_44089,N_37167,N_38257);
and U44090 (N_44090,N_31876,N_31320);
and U44091 (N_44091,N_33319,N_33848);
xor U44092 (N_44092,N_33161,N_35118);
nand U44093 (N_44093,N_30709,N_36272);
or U44094 (N_44094,N_38136,N_39953);
or U44095 (N_44095,N_30467,N_38671);
or U44096 (N_44096,N_36320,N_31731);
nor U44097 (N_44097,N_37877,N_32675);
nor U44098 (N_44098,N_37080,N_31726);
or U44099 (N_44099,N_38991,N_33859);
and U44100 (N_44100,N_31915,N_30888);
nor U44101 (N_44101,N_36851,N_35854);
or U44102 (N_44102,N_33508,N_36071);
and U44103 (N_44103,N_30066,N_31520);
nand U44104 (N_44104,N_36116,N_31584);
and U44105 (N_44105,N_34630,N_35214);
or U44106 (N_44106,N_34500,N_37494);
nor U44107 (N_44107,N_30272,N_34913);
and U44108 (N_44108,N_38469,N_36128);
nand U44109 (N_44109,N_31752,N_37976);
or U44110 (N_44110,N_34728,N_39340);
or U44111 (N_44111,N_36501,N_36426);
nor U44112 (N_44112,N_30234,N_30718);
xor U44113 (N_44113,N_34441,N_35368);
or U44114 (N_44114,N_36729,N_35585);
and U44115 (N_44115,N_36370,N_38181);
or U44116 (N_44116,N_35924,N_38179);
xor U44117 (N_44117,N_33902,N_35121);
nor U44118 (N_44118,N_39437,N_36684);
and U44119 (N_44119,N_38696,N_32184);
or U44120 (N_44120,N_34613,N_34620);
nand U44121 (N_44121,N_37366,N_31562);
and U44122 (N_44122,N_32186,N_37398);
xnor U44123 (N_44123,N_32335,N_32023);
or U44124 (N_44124,N_35484,N_33498);
nand U44125 (N_44125,N_36119,N_34336);
nor U44126 (N_44126,N_34043,N_35900);
nor U44127 (N_44127,N_34936,N_34038);
xnor U44128 (N_44128,N_32570,N_39874);
nor U44129 (N_44129,N_39652,N_38042);
nor U44130 (N_44130,N_32194,N_31783);
nor U44131 (N_44131,N_30862,N_31048);
or U44132 (N_44132,N_37089,N_32651);
nor U44133 (N_44133,N_38084,N_38796);
or U44134 (N_44134,N_32662,N_38855);
nand U44135 (N_44135,N_37371,N_31931);
or U44136 (N_44136,N_34188,N_36827);
nor U44137 (N_44137,N_32961,N_31177);
or U44138 (N_44138,N_35706,N_34778);
nor U44139 (N_44139,N_36091,N_31108);
xnor U44140 (N_44140,N_36993,N_34360);
xnor U44141 (N_44141,N_30667,N_35893);
nor U44142 (N_44142,N_37991,N_35086);
nor U44143 (N_44143,N_33466,N_32342);
or U44144 (N_44144,N_37214,N_39068);
and U44145 (N_44145,N_33980,N_31519);
or U44146 (N_44146,N_34911,N_33215);
nand U44147 (N_44147,N_30318,N_34300);
and U44148 (N_44148,N_30099,N_35356);
nor U44149 (N_44149,N_38974,N_35548);
or U44150 (N_44150,N_37207,N_39325);
nand U44151 (N_44151,N_30009,N_36316);
nor U44152 (N_44152,N_37468,N_34469);
nor U44153 (N_44153,N_31072,N_33970);
nand U44154 (N_44154,N_31361,N_39038);
or U44155 (N_44155,N_36947,N_30565);
nor U44156 (N_44156,N_31319,N_31436);
nor U44157 (N_44157,N_38972,N_32406);
or U44158 (N_44158,N_38522,N_32837);
and U44159 (N_44159,N_37381,N_38746);
xor U44160 (N_44160,N_35693,N_32209);
nand U44161 (N_44161,N_35953,N_35076);
or U44162 (N_44162,N_30267,N_32443);
and U44163 (N_44163,N_31902,N_34891);
xor U44164 (N_44164,N_37712,N_30154);
and U44165 (N_44165,N_34732,N_36653);
nor U44166 (N_44166,N_30649,N_38326);
or U44167 (N_44167,N_32681,N_33981);
or U44168 (N_44168,N_34400,N_34905);
or U44169 (N_44169,N_31983,N_37636);
and U44170 (N_44170,N_30955,N_39813);
and U44171 (N_44171,N_33134,N_36840);
or U44172 (N_44172,N_31888,N_36001);
nor U44173 (N_44173,N_39319,N_35332);
nor U44174 (N_44174,N_32532,N_34421);
or U44175 (N_44175,N_32598,N_37312);
xnor U44176 (N_44176,N_35008,N_36268);
nand U44177 (N_44177,N_32772,N_30648);
or U44178 (N_44178,N_33110,N_32421);
xnor U44179 (N_44179,N_32862,N_34419);
or U44180 (N_44180,N_34138,N_37314);
and U44181 (N_44181,N_31043,N_39427);
nand U44182 (N_44182,N_32969,N_33960);
nand U44183 (N_44183,N_31940,N_39927);
nand U44184 (N_44184,N_30161,N_33024);
nor U44185 (N_44185,N_31357,N_31202);
xnor U44186 (N_44186,N_39729,N_31310);
and U44187 (N_44187,N_33808,N_35876);
or U44188 (N_44188,N_37206,N_38209);
nand U44189 (N_44189,N_31134,N_30889);
nor U44190 (N_44190,N_32872,N_33565);
or U44191 (N_44191,N_30858,N_32398);
nand U44192 (N_44192,N_32042,N_34954);
nand U44193 (N_44193,N_33743,N_33870);
or U44194 (N_44194,N_33417,N_35280);
nor U44195 (N_44195,N_32704,N_35021);
or U44196 (N_44196,N_33695,N_32928);
or U44197 (N_44197,N_30707,N_36022);
nor U44198 (N_44198,N_31988,N_34109);
nor U44199 (N_44199,N_34418,N_32937);
nand U44200 (N_44200,N_36136,N_37629);
and U44201 (N_44201,N_37908,N_37000);
or U44202 (N_44202,N_39069,N_39462);
nand U44203 (N_44203,N_34917,N_32032);
nor U44204 (N_44204,N_33853,N_38559);
and U44205 (N_44205,N_30827,N_39583);
nand U44206 (N_44206,N_35115,N_36493);
or U44207 (N_44207,N_35005,N_39484);
xor U44208 (N_44208,N_38355,N_34711);
or U44209 (N_44209,N_39865,N_38823);
and U44210 (N_44210,N_30876,N_32320);
nor U44211 (N_44211,N_33966,N_31393);
nor U44212 (N_44212,N_38753,N_36738);
xnor U44213 (N_44213,N_36889,N_33685);
nand U44214 (N_44214,N_34532,N_37805);
or U44215 (N_44215,N_36886,N_34463);
and U44216 (N_44216,N_32771,N_33234);
nand U44217 (N_44217,N_36234,N_39305);
xnor U44218 (N_44218,N_38440,N_38160);
nor U44219 (N_44219,N_38073,N_35618);
nand U44220 (N_44220,N_30254,N_33439);
and U44221 (N_44221,N_34569,N_35380);
xnor U44222 (N_44222,N_33440,N_33250);
nand U44223 (N_44223,N_38650,N_32693);
xor U44224 (N_44224,N_38777,N_39706);
nand U44225 (N_44225,N_36996,N_34582);
xnor U44226 (N_44226,N_39925,N_31625);
and U44227 (N_44227,N_31875,N_37986);
nand U44228 (N_44228,N_37285,N_31760);
nand U44229 (N_44229,N_32869,N_30138);
nand U44230 (N_44230,N_35599,N_39193);
and U44231 (N_44231,N_31617,N_37523);
and U44232 (N_44232,N_33331,N_32183);
and U44233 (N_44233,N_32864,N_39904);
nand U44234 (N_44234,N_32254,N_37339);
or U44235 (N_44235,N_39279,N_35863);
and U44236 (N_44236,N_33553,N_35320);
xnor U44237 (N_44237,N_39435,N_36906);
or U44238 (N_44238,N_35398,N_38535);
xnor U44239 (N_44239,N_34014,N_36925);
and U44240 (N_44240,N_30390,N_37252);
and U44241 (N_44241,N_30059,N_35652);
or U44242 (N_44242,N_33038,N_33597);
and U44243 (N_44243,N_39044,N_30999);
and U44244 (N_44244,N_33756,N_37428);
nand U44245 (N_44245,N_35414,N_30004);
and U44246 (N_44246,N_36107,N_35338);
or U44247 (N_44247,N_31905,N_33841);
nand U44248 (N_44248,N_35586,N_38353);
nand U44249 (N_44249,N_31705,N_35659);
and U44250 (N_44250,N_37542,N_37106);
nor U44251 (N_44251,N_35718,N_36144);
and U44252 (N_44252,N_31203,N_38008);
or U44253 (N_44253,N_38722,N_39135);
or U44254 (N_44254,N_37567,N_36423);
nor U44255 (N_44255,N_33671,N_36575);
nand U44256 (N_44256,N_37587,N_30001);
nor U44257 (N_44257,N_31262,N_37154);
and U44258 (N_44258,N_37808,N_39666);
nor U44259 (N_44259,N_35657,N_38441);
and U44260 (N_44260,N_38311,N_38434);
xor U44261 (N_44261,N_39214,N_31530);
or U44262 (N_44262,N_32519,N_37679);
or U44263 (N_44263,N_31178,N_33281);
nand U44264 (N_44264,N_35051,N_30871);
or U44265 (N_44265,N_33616,N_30740);
or U44266 (N_44266,N_38294,N_30857);
nor U44267 (N_44267,N_32625,N_36777);
or U44268 (N_44268,N_34860,N_30115);
xnor U44269 (N_44269,N_32743,N_37345);
nand U44270 (N_44270,N_34042,N_38045);
xnor U44271 (N_44271,N_39811,N_35904);
nor U44272 (N_44272,N_31485,N_36280);
nand U44273 (N_44273,N_37300,N_31465);
nand U44274 (N_44274,N_31414,N_38266);
nand U44275 (N_44275,N_36383,N_39501);
nor U44276 (N_44276,N_36527,N_39546);
or U44277 (N_44277,N_33295,N_30191);
xnor U44278 (N_44278,N_37202,N_35079);
xor U44279 (N_44279,N_37887,N_39064);
and U44280 (N_44280,N_34731,N_39398);
or U44281 (N_44281,N_33028,N_33624);
or U44282 (N_44282,N_38749,N_37708);
nand U44283 (N_44283,N_39320,N_32359);
nor U44284 (N_44284,N_34736,N_37727);
and U44285 (N_44285,N_33995,N_36442);
nand U44286 (N_44286,N_33213,N_36766);
nand U44287 (N_44287,N_32767,N_30942);
nand U44288 (N_44288,N_38733,N_33219);
and U44289 (N_44289,N_30938,N_37750);
nand U44290 (N_44290,N_33691,N_31962);
and U44291 (N_44291,N_35129,N_31435);
or U44292 (N_44292,N_37258,N_32510);
nand U44293 (N_44293,N_30100,N_31877);
nor U44294 (N_44294,N_38847,N_38091);
nor U44295 (N_44295,N_36283,N_37246);
and U44296 (N_44296,N_32972,N_33972);
or U44297 (N_44297,N_32303,N_30923);
nand U44298 (N_44298,N_37948,N_35475);
nand U44299 (N_44299,N_36125,N_33734);
xor U44300 (N_44300,N_39416,N_30625);
nor U44301 (N_44301,N_38479,N_35615);
or U44302 (N_44302,N_39663,N_36298);
nor U44303 (N_44303,N_34737,N_33495);
nor U44304 (N_44304,N_34811,N_37204);
nand U44305 (N_44305,N_33006,N_33566);
nor U44306 (N_44306,N_30536,N_31114);
or U44307 (N_44307,N_32726,N_38544);
and U44308 (N_44308,N_38372,N_33899);
nor U44309 (N_44309,N_30934,N_33973);
and U44310 (N_44310,N_34767,N_30578);
nand U44311 (N_44311,N_31111,N_32268);
nand U44312 (N_44312,N_38276,N_30170);
xor U44313 (N_44313,N_36534,N_38138);
and U44314 (N_44314,N_33731,N_38952);
nor U44315 (N_44315,N_36606,N_35541);
or U44316 (N_44316,N_39945,N_32896);
nor U44317 (N_44317,N_33171,N_35420);
xor U44318 (N_44318,N_32136,N_35645);
nand U44319 (N_44319,N_39458,N_31347);
and U44320 (N_44320,N_36583,N_37718);
nand U44321 (N_44321,N_35576,N_35603);
and U44322 (N_44322,N_34493,N_30323);
and U44323 (N_44323,N_39876,N_38219);
nor U44324 (N_44324,N_36108,N_30238);
and U44325 (N_44325,N_32033,N_30611);
or U44326 (N_44326,N_31412,N_37220);
nor U44327 (N_44327,N_35852,N_39206);
or U44328 (N_44328,N_33728,N_36326);
nand U44329 (N_44329,N_36211,N_38614);
nor U44330 (N_44330,N_36662,N_34887);
and U44331 (N_44331,N_38203,N_37139);
or U44332 (N_44332,N_38102,N_34937);
xor U44333 (N_44333,N_34432,N_37295);
nor U44334 (N_44334,N_39928,N_36498);
xnor U44335 (N_44335,N_39366,N_35135);
nor U44336 (N_44336,N_34962,N_32569);
nor U44337 (N_44337,N_34395,N_38158);
nor U44338 (N_44338,N_34282,N_36256);
nand U44339 (N_44339,N_30236,N_36915);
or U44340 (N_44340,N_31803,N_32907);
nand U44341 (N_44341,N_37601,N_38616);
nand U44342 (N_44342,N_31426,N_32610);
or U44343 (N_44343,N_34153,N_35180);
and U44344 (N_44344,N_36796,N_36186);
nor U44345 (N_44345,N_34396,N_31404);
or U44346 (N_44346,N_32518,N_34020);
nand U44347 (N_44347,N_39329,N_30150);
nor U44348 (N_44348,N_31104,N_34774);
or U44349 (N_44349,N_31992,N_33640);
nand U44350 (N_44350,N_34340,N_39058);
nor U44351 (N_44351,N_39020,N_30185);
nor U44352 (N_44352,N_34082,N_33399);
nor U44353 (N_44353,N_31683,N_31686);
nor U44354 (N_44354,N_34417,N_33330);
or U44355 (N_44355,N_35570,N_39436);
nand U44356 (N_44356,N_39089,N_31574);
nor U44357 (N_44357,N_32629,N_35157);
xor U44358 (N_44358,N_39326,N_35432);
and U44359 (N_44359,N_35242,N_37449);
xor U44360 (N_44360,N_38757,N_32432);
nand U44361 (N_44361,N_32360,N_37701);
nand U44362 (N_44362,N_35181,N_30092);
nor U44363 (N_44363,N_39027,N_34981);
nand U44364 (N_44364,N_37335,N_36445);
and U44365 (N_44365,N_39241,N_36340);
and U44366 (N_44366,N_39235,N_30397);
nor U44367 (N_44367,N_32076,N_32641);
nand U44368 (N_44368,N_37598,N_38552);
or U44369 (N_44369,N_31212,N_38596);
and U44370 (N_44370,N_35891,N_36805);
or U44371 (N_44371,N_31160,N_33497);
nand U44372 (N_44372,N_30255,N_30533);
or U44373 (N_44373,N_30563,N_38618);
and U44374 (N_44374,N_36229,N_32073);
nor U44375 (N_44375,N_37102,N_35537);
or U44376 (N_44376,N_39514,N_38445);
nand U44377 (N_44377,N_39341,N_39408);
or U44378 (N_44378,N_37654,N_39252);
and U44379 (N_44379,N_35637,N_38111);
nand U44380 (N_44380,N_39195,N_36299);
or U44381 (N_44381,N_30471,N_38930);
or U44382 (N_44382,N_35462,N_30869);
or U44383 (N_44383,N_34857,N_38806);
nor U44384 (N_44384,N_39975,N_32276);
nand U44385 (N_44385,N_34087,N_30890);
nor U44386 (N_44386,N_38271,N_36718);
nand U44387 (N_44387,N_39144,N_30269);
xnor U44388 (N_44388,N_32995,N_31930);
or U44389 (N_44389,N_38188,N_37218);
nor U44390 (N_44390,N_37922,N_30071);
nand U44391 (N_44391,N_39502,N_36007);
nor U44392 (N_44392,N_37169,N_39078);
nor U44393 (N_44393,N_39741,N_32867);
nand U44394 (N_44394,N_32846,N_31133);
nand U44395 (N_44395,N_34585,N_32295);
nor U44396 (N_44396,N_36168,N_30371);
or U44397 (N_44397,N_37039,N_32944);
nand U44398 (N_44398,N_32795,N_39746);
or U44399 (N_44399,N_31105,N_32273);
and U44400 (N_44400,N_37661,N_31892);
and U44401 (N_44401,N_37047,N_31030);
or U44402 (N_44402,N_38969,N_38279);
and U44403 (N_44403,N_39867,N_33448);
nand U44404 (N_44404,N_34051,N_32621);
or U44405 (N_44405,N_37752,N_39709);
nand U44406 (N_44406,N_37710,N_36516);
nor U44407 (N_44407,N_36332,N_38142);
or U44408 (N_44408,N_30355,N_32242);
and U44409 (N_44409,N_32873,N_35767);
or U44410 (N_44410,N_36297,N_31243);
nor U44411 (N_44411,N_39400,N_36638);
nand U44412 (N_44412,N_38497,N_34378);
or U44413 (N_44413,N_37681,N_39806);
and U44414 (N_44414,N_38993,N_36762);
nor U44415 (N_44415,N_31163,N_37035);
nor U44416 (N_44416,N_38189,N_36028);
xnor U44417 (N_44417,N_36878,N_36328);
nor U44418 (N_44418,N_33368,N_35945);
or U44419 (N_44419,N_36999,N_38225);
or U44420 (N_44420,N_30249,N_32434);
and U44421 (N_44421,N_34881,N_36601);
nor U44422 (N_44422,N_34005,N_37318);
and U44423 (N_44423,N_34343,N_32021);
and U44424 (N_44424,N_31593,N_31582);
nand U44425 (N_44425,N_34951,N_30039);
nand U44426 (N_44426,N_32934,N_38536);
or U44427 (N_44427,N_34272,N_30971);
nor U44428 (N_44428,N_33683,N_38005);
or U44429 (N_44429,N_31882,N_39947);
or U44430 (N_44430,N_33212,N_30005);
nand U44431 (N_44431,N_34789,N_31935);
nor U44432 (N_44432,N_38247,N_30461);
nor U44433 (N_44433,N_39685,N_39440);
nand U44434 (N_44434,N_33101,N_33011);
and U44435 (N_44435,N_30995,N_32729);
or U44436 (N_44436,N_31637,N_37818);
nand U44437 (N_44437,N_33680,N_35692);
nand U44438 (N_44438,N_30028,N_36530);
nand U44439 (N_44439,N_33479,N_31744);
or U44440 (N_44440,N_33165,N_33491);
nand U44441 (N_44441,N_39190,N_35877);
or U44442 (N_44442,N_36435,N_31626);
xor U44443 (N_44443,N_33886,N_39544);
and U44444 (N_44444,N_31293,N_34160);
xnor U44445 (N_44445,N_37445,N_39631);
and U44446 (N_44446,N_38190,N_39762);
nor U44447 (N_44447,N_38521,N_37118);
and U44448 (N_44448,N_35840,N_38998);
nand U44449 (N_44449,N_34345,N_32412);
and U44450 (N_44450,N_37778,N_35062);
and U44451 (N_44451,N_31777,N_31511);
and U44452 (N_44452,N_36966,N_37391);
and U44453 (N_44453,N_39721,N_39029);
or U44454 (N_44454,N_37425,N_37150);
or U44455 (N_44455,N_37757,N_39581);
and U44456 (N_44456,N_39037,N_34568);
xnor U44457 (N_44457,N_33664,N_30870);
xor U44458 (N_44458,N_34693,N_33045);
nor U44459 (N_44459,N_32895,N_33735);
xnor U44460 (N_44460,N_36135,N_36401);
and U44461 (N_44461,N_37121,N_33601);
and U44462 (N_44462,N_36009,N_39328);
nor U44463 (N_44463,N_37559,N_32229);
or U44464 (N_44464,N_38421,N_30153);
and U44465 (N_44465,N_34192,N_38028);
nand U44466 (N_44466,N_39351,N_33676);
nand U44467 (N_44467,N_32956,N_33747);
nand U44468 (N_44468,N_39724,N_36225);
or U44469 (N_44469,N_37313,N_32838);
nor U44470 (N_44470,N_33354,N_32314);
nand U44471 (N_44471,N_38015,N_31509);
nor U44472 (N_44472,N_35071,N_38054);
or U44473 (N_44473,N_39667,N_34864);
nor U44474 (N_44474,N_35580,N_36919);
nand U44475 (N_44475,N_33586,N_31914);
nand U44476 (N_44476,N_30116,N_38055);
or U44477 (N_44477,N_31566,N_37044);
and U44478 (N_44478,N_37078,N_30473);
or U44479 (N_44479,N_31052,N_31380);
and U44480 (N_44480,N_37040,N_30175);
nor U44481 (N_44481,N_39974,N_31287);
nand U44482 (N_44482,N_30246,N_31793);
nor U44483 (N_44483,N_37378,N_34354);
nor U44484 (N_44484,N_37635,N_37749);
and U44485 (N_44485,N_37743,N_39692);
or U44486 (N_44486,N_37622,N_35647);
nor U44487 (N_44487,N_39308,N_36787);
and U44488 (N_44488,N_33992,N_39467);
or U44489 (N_44489,N_33069,N_37131);
or U44490 (N_44490,N_37916,N_35922);
nor U44491 (N_44491,N_35138,N_38364);
or U44492 (N_44492,N_32458,N_30406);
nand U44493 (N_44493,N_39301,N_39550);
or U44494 (N_44494,N_31416,N_37166);
nor U44495 (N_44495,N_32537,N_36560);
or U44496 (N_44496,N_37906,N_35470);
and U44497 (N_44497,N_32270,N_30056);
or U44498 (N_44498,N_32001,N_38123);
xor U44499 (N_44499,N_31200,N_38292);
nor U44500 (N_44500,N_35540,N_37900);
xor U44501 (N_44501,N_37340,N_35755);
and U44502 (N_44502,N_39003,N_34484);
nor U44503 (N_44503,N_33327,N_37525);
and U44504 (N_44504,N_32866,N_34746);
xnor U44505 (N_44505,N_38267,N_37741);
xnor U44506 (N_44506,N_35919,N_33218);
or U44507 (N_44507,N_35025,N_31355);
nand U44508 (N_44508,N_32174,N_34750);
and U44509 (N_44509,N_32758,N_30273);
nor U44510 (N_44510,N_33542,N_36848);
and U44511 (N_44511,N_30973,N_38883);
or U44512 (N_44512,N_31609,N_36818);
nand U44513 (N_44513,N_30621,N_37570);
nor U44514 (N_44514,N_30492,N_34571);
or U44515 (N_44515,N_35600,N_39459);
nor U44516 (N_44516,N_38844,N_33349);
nor U44517 (N_44517,N_39134,N_35871);
or U44518 (N_44518,N_37192,N_39630);
xor U44519 (N_44519,N_39731,N_34084);
xnor U44520 (N_44520,N_38116,N_33030);
nand U44521 (N_44521,N_35276,N_39346);
and U44522 (N_44522,N_36529,N_38222);
nor U44523 (N_44523,N_35069,N_37088);
and U44524 (N_44524,N_32286,N_31217);
nand U44525 (N_44525,N_33119,N_31407);
nand U44526 (N_44526,N_36568,N_30772);
or U44527 (N_44527,N_31318,N_34842);
and U44528 (N_44528,N_32102,N_33451);
xor U44529 (N_44529,N_37360,N_30041);
or U44530 (N_44530,N_37170,N_39687);
and U44531 (N_44531,N_32250,N_35006);
nand U44532 (N_44532,N_34315,N_33842);
nor U44533 (N_44533,N_39695,N_34682);
nor U44534 (N_44534,N_31070,N_31523);
and U44535 (N_44535,N_39056,N_32894);
nor U44536 (N_44536,N_32579,N_35510);
nand U44537 (N_44537,N_34543,N_37455);
nand U44538 (N_44538,N_30670,N_34466);
nand U44539 (N_44539,N_36842,N_37604);
nand U44540 (N_44540,N_39491,N_36864);
nor U44541 (N_44541,N_37912,N_34498);
or U44542 (N_44542,N_31568,N_37579);
and U44543 (N_44543,N_30587,N_39083);
nand U44544 (N_44544,N_34357,N_34033);
or U44545 (N_44545,N_33366,N_31949);
nand U44546 (N_44546,N_31687,N_30945);
nand U44547 (N_44547,N_35460,N_39430);
nor U44548 (N_44548,N_38146,N_31425);
nand U44549 (N_44549,N_37841,N_34777);
xor U44550 (N_44550,N_39576,N_33394);
nor U44551 (N_44551,N_32244,N_36120);
nor U44552 (N_44552,N_38379,N_37281);
xnor U44553 (N_44553,N_30274,N_32170);
nor U44554 (N_44554,N_33092,N_39633);
xnor U44555 (N_44555,N_36337,N_32282);
or U44556 (N_44556,N_38764,N_34906);
xor U44557 (N_44557,N_39950,N_38155);
xnor U44558 (N_44558,N_30680,N_30165);
or U44559 (N_44559,N_30953,N_35874);
or U44560 (N_44560,N_32212,N_32444);
xor U44561 (N_44561,N_37694,N_31597);
nand U44562 (N_44562,N_32382,N_30984);
nor U44563 (N_44563,N_35339,N_30708);
and U44564 (N_44564,N_35192,N_39849);
or U44565 (N_44565,N_39759,N_32507);
and U44566 (N_44566,N_33936,N_32676);
nand U44567 (N_44567,N_38790,N_30927);
and U44568 (N_44568,N_38195,N_35259);
or U44569 (N_44569,N_35993,N_31642);
nor U44570 (N_44570,N_34640,N_36911);
nand U44571 (N_44571,N_38043,N_31515);
or U44572 (N_44572,N_35012,N_35354);
nor U44573 (N_44573,N_31542,N_34772);
and U44574 (N_44574,N_33827,N_39412);
and U44575 (N_44575,N_31569,N_37502);
and U44576 (N_44576,N_36304,N_30383);
or U44577 (N_44577,N_38464,N_36160);
nand U44578 (N_44578,N_39602,N_37730);
xnor U44579 (N_44579,N_35949,N_38154);
nor U44580 (N_44580,N_38986,N_38756);
nor U44581 (N_44581,N_37786,N_33288);
nand U44582 (N_44582,N_33510,N_34909);
and U44583 (N_44583,N_35417,N_35185);
or U44584 (N_44584,N_30222,N_34294);
nor U44585 (N_44585,N_35016,N_38443);
nand U44586 (N_44586,N_38655,N_38482);
and U44587 (N_44587,N_32256,N_35638);
or U44588 (N_44588,N_33459,N_34239);
nor U44589 (N_44589,N_35822,N_38036);
and U44590 (N_44590,N_38697,N_38932);
or U44591 (N_44591,N_37639,N_37845);
and U44592 (N_44592,N_30158,N_31182);
xnor U44593 (N_44593,N_34703,N_33781);
or U44594 (N_44594,N_37087,N_30454);
and U44595 (N_44595,N_32520,N_36882);
and U44596 (N_44596,N_35680,N_31069);
or U44597 (N_44597,N_39735,N_38461);
xnor U44598 (N_44598,N_39498,N_30198);
and U44599 (N_44599,N_31922,N_37856);
nand U44600 (N_44600,N_33753,N_38925);
and U44601 (N_44601,N_36145,N_32025);
nor U44602 (N_44602,N_36412,N_37643);
nor U44603 (N_44603,N_34261,N_39548);
and U44604 (N_44604,N_32732,N_39248);
xor U44605 (N_44605,N_30968,N_34807);
nand U44606 (N_44606,N_35716,N_39177);
nor U44607 (N_44607,N_36655,N_33962);
and U44608 (N_44608,N_30207,N_36630);
nor U44609 (N_44609,N_30252,N_34931);
and U44610 (N_44610,N_34302,N_35872);
xor U44611 (N_44611,N_39219,N_37489);
and U44612 (N_44612,N_38157,N_39789);
and U44613 (N_44613,N_32702,N_31679);
nor U44614 (N_44614,N_34494,N_32128);
nand U44615 (N_44615,N_39251,N_30407);
nor U44616 (N_44616,N_35948,N_33113);
nor U44617 (N_44617,N_37539,N_38476);
and U44618 (N_44618,N_32383,N_33068);
or U44619 (N_44619,N_36362,N_33742);
nand U44620 (N_44620,N_36172,N_37441);
nor U44621 (N_44621,N_35787,N_32074);
and U44622 (N_44622,N_35744,N_38194);
or U44623 (N_44623,N_39841,N_34422);
nor U44624 (N_44624,N_30297,N_36002);
nor U44625 (N_44625,N_34289,N_39785);
xor U44626 (N_44626,N_36064,N_35721);
or U44627 (N_44627,N_35821,N_35445);
nand U44628 (N_44628,N_38767,N_32142);
xor U44629 (N_44629,N_31773,N_31936);
nand U44630 (N_44630,N_31149,N_33916);
nand U44631 (N_44631,N_32040,N_33263);
nor U44632 (N_44632,N_31015,N_32442);
xnor U44633 (N_44633,N_32670,N_37482);
or U44634 (N_44634,N_36586,N_39733);
and U44635 (N_44635,N_32727,N_39379);
nor U44636 (N_44636,N_36082,N_38350);
xor U44637 (N_44637,N_37303,N_36411);
nor U44638 (N_44638,N_39082,N_37509);
nand U44639 (N_44639,N_39885,N_39933);
or U44640 (N_44640,N_30235,N_35483);
and U44641 (N_44641,N_34348,N_34672);
or U44642 (N_44642,N_33845,N_31693);
nand U44643 (N_44643,N_30122,N_35746);
nand U44644 (N_44644,N_36776,N_36171);
nand U44645 (N_44645,N_31294,N_38378);
nand U44646 (N_44646,N_34447,N_35810);
or U44647 (N_44647,N_33296,N_33460);
and U44648 (N_44648,N_35897,N_36914);
nor U44649 (N_44649,N_34757,N_39842);
or U44650 (N_44650,N_32047,N_36486);
and U44651 (N_44651,N_30242,N_35567);
nand U44652 (N_44652,N_36749,N_36843);
nand U44653 (N_44653,N_36215,N_36902);
nor U44654 (N_44654,N_36803,N_34062);
or U44655 (N_44655,N_32162,N_35184);
and U44656 (N_44656,N_34132,N_37762);
nor U44657 (N_44657,N_35348,N_34717);
nor U44658 (N_44658,N_33654,N_35273);
nor U44659 (N_44659,N_32098,N_39653);
nand U44660 (N_44660,N_33904,N_39783);
or U44661 (N_44661,N_37773,N_32189);
and U44662 (N_44662,N_35929,N_38375);
nand U44663 (N_44663,N_37532,N_36695);
and U44664 (N_44664,N_30776,N_36962);
xor U44665 (N_44665,N_39446,N_30576);
and U44666 (N_44666,N_39503,N_38874);
nand U44667 (N_44667,N_34967,N_32965);
or U44668 (N_44668,N_39290,N_35583);
or U44669 (N_44669,N_36572,N_39749);
or U44670 (N_44670,N_30668,N_30814);
nand U44671 (N_44671,N_30378,N_34647);
nor U44672 (N_44672,N_31196,N_37994);
or U44673 (N_44673,N_39730,N_31258);
or U44674 (N_44674,N_38109,N_37486);
or U44675 (N_44675,N_33367,N_39352);
nor U44676 (N_44676,N_37140,N_32472);
nand U44677 (N_44677,N_38420,N_39960);
nor U44678 (N_44678,N_35399,N_39808);
nor U44679 (N_44679,N_39131,N_39246);
nand U44680 (N_44680,N_37650,N_32661);
and U44681 (N_44681,N_39492,N_39567);
or U44682 (N_44682,N_31947,N_35547);
nor U44683 (N_44683,N_36407,N_38256);
nor U44684 (N_44684,N_38557,N_37249);
nor U44685 (N_44685,N_39499,N_39820);
and U44686 (N_44686,N_37775,N_36849);
nand U44687 (N_44687,N_31527,N_31397);
or U44688 (N_44688,N_38725,N_39495);
or U44689 (N_44689,N_31924,N_32381);
xor U44690 (N_44690,N_33079,N_32090);
nor U44691 (N_44691,N_31440,N_30856);
nor U44692 (N_44692,N_35761,N_30127);
or U44693 (N_44693,N_39149,N_38513);
and U44694 (N_44694,N_37008,N_36156);
nand U44695 (N_44695,N_32874,N_35057);
or U44696 (N_44696,N_32195,N_32805);
or U44697 (N_44697,N_35154,N_31559);
and U44698 (N_44698,N_34338,N_38677);
or U44699 (N_44699,N_34513,N_36508);
or U44700 (N_44700,N_36345,N_39129);
nand U44701 (N_44701,N_33203,N_38726);
and U44702 (N_44702,N_35241,N_38601);
nand U44703 (N_44703,N_38218,N_31490);
nand U44704 (N_44704,N_37578,N_30118);
and U44705 (N_44705,N_30047,N_32459);
nor U44706 (N_44706,N_35390,N_36732);
nand U44707 (N_44707,N_30661,N_35935);
xor U44708 (N_44708,N_39951,N_36860);
or U44709 (N_44709,N_35523,N_30411);
xnor U44710 (N_44710,N_34575,N_30686);
and U44711 (N_44711,N_36725,N_32657);
and U44712 (N_44712,N_38922,N_39932);
nand U44713 (N_44713,N_36312,N_30421);
or U44714 (N_44714,N_38693,N_33013);
nand U44715 (N_44715,N_33961,N_38423);
nand U44716 (N_44716,N_37540,N_30795);
nor U44717 (N_44717,N_38701,N_39451);
and U44718 (N_44718,N_32488,N_34375);
nand U44719 (N_44719,N_31717,N_38081);
xnor U44720 (N_44720,N_34562,N_32435);
nor U44721 (N_44721,N_38394,N_30521);
and U44722 (N_44722,N_33225,N_31299);
nor U44723 (N_44723,N_34318,N_30289);
xnor U44724 (N_44724,N_38679,N_33718);
nor U44725 (N_44725,N_35169,N_33507);
nand U44726 (N_44726,N_38592,N_35149);
nand U44727 (N_44727,N_33849,N_39771);
nand U44728 (N_44728,N_35629,N_34952);
and U44729 (N_44729,N_37029,N_39074);
nand U44730 (N_44730,N_32852,N_33736);
nand U44731 (N_44731,N_38607,N_35735);
nand U44732 (N_44732,N_30241,N_30908);
nor U44733 (N_44733,N_31081,N_39688);
and U44734 (N_44734,N_39684,N_36478);
and U44735 (N_44735,N_37767,N_30498);
and U44736 (N_44736,N_30413,N_36049);
or U44737 (N_44737,N_38788,N_39644);
xnor U44738 (N_44738,N_31097,N_38252);
nand U44739 (N_44739,N_37696,N_39052);
nor U44740 (N_44740,N_31198,N_36479);
nor U44741 (N_44741,N_36997,N_39281);
and U44742 (N_44742,N_33689,N_31618);
and U44743 (N_44743,N_35867,N_33189);
or U44744 (N_44744,N_34017,N_34332);
or U44745 (N_44745,N_33999,N_34914);
nand U44746 (N_44746,N_34990,N_32218);
nand U44747 (N_44747,N_30509,N_32588);
and U44748 (N_44748,N_30178,N_37753);
xnor U44749 (N_44749,N_33773,N_37304);
and U44750 (N_44750,N_34086,N_37610);
nand U44751 (N_44751,N_31057,N_34627);
and U44752 (N_44752,N_34230,N_39591);
xor U44753 (N_44753,N_37056,N_37498);
nand U44754 (N_44754,N_39338,N_33927);
nand U44755 (N_44755,N_30868,N_30935);
or U44756 (N_44756,N_31481,N_30895);
nand U44757 (N_44757,N_30549,N_37496);
or U44758 (N_44758,N_32877,N_34578);
nand U44759 (N_44759,N_31951,N_36794);
xor U44760 (N_44760,N_39963,N_35331);
nor U44761 (N_44761,N_38966,N_31685);
and U44762 (N_44762,N_36242,N_38617);
nand U44763 (N_44763,N_34506,N_33055);
nand U44764 (N_44764,N_36817,N_36750);
nand U44765 (N_44765,N_36398,N_31798);
nor U44766 (N_44766,N_39194,N_33610);
and U44767 (N_44767,N_39296,N_32366);
or U44768 (N_44768,N_30310,N_39792);
or U44769 (N_44769,N_33933,N_30980);
nor U44770 (N_44770,N_39115,N_35075);
nand U44771 (N_44771,N_30016,N_33822);
nor U44772 (N_44772,N_36444,N_37132);
xor U44773 (N_44773,N_37043,N_33525);
and U44774 (N_44774,N_36909,N_32269);
or U44775 (N_44775,N_36728,N_31170);
nand U44776 (N_44776,N_34195,N_36900);
and U44777 (N_44777,N_33722,N_37891);
or U44778 (N_44778,N_35137,N_37843);
or U44779 (N_44779,N_31116,N_36404);
xor U44780 (N_44780,N_34971,N_32199);
or U44781 (N_44781,N_33064,N_38761);
or U44782 (N_44782,N_38970,N_36405);
and U44783 (N_44783,N_37273,N_37286);
and U44784 (N_44784,N_31122,N_36189);
xor U44785 (N_44785,N_31969,N_38467);
or U44786 (N_44786,N_33334,N_31912);
or U44787 (N_44787,N_38221,N_35133);
nor U44788 (N_44788,N_30695,N_30609);
and U44789 (N_44789,N_36315,N_37201);
xor U44790 (N_44790,N_38971,N_30052);
or U44791 (N_44791,N_33802,N_35183);
nand U44792 (N_44792,N_38789,N_37461);
nor U44793 (N_44793,N_37347,N_36798);
or U44794 (N_44794,N_37145,N_33419);
nand U44795 (N_44795,N_35831,N_32445);
or U44796 (N_44796,N_38229,N_31362);
nand U44797 (N_44797,N_34054,N_32207);
and U44798 (N_44798,N_38471,N_30614);
and U44799 (N_44799,N_31900,N_31899);
nand U44800 (N_44800,N_38961,N_35495);
and U44801 (N_44801,N_38345,N_32669);
and U44802 (N_44802,N_34854,N_39722);
or U44803 (N_44803,N_34309,N_30912);
nor U44804 (N_44804,N_36181,N_37100);
and U44805 (N_44805,N_38117,N_35894);
or U44806 (N_44806,N_32674,N_36348);
and U44807 (N_44807,N_32492,N_36469);
and U44808 (N_44808,N_39973,N_39861);
and U44809 (N_44809,N_37319,N_34149);
and U44810 (N_44810,N_33202,N_37770);
nor U44811 (N_44811,N_31761,N_30562);
and U44812 (N_44812,N_34412,N_32970);
nor U44813 (N_44813,N_37350,N_33364);
and U44814 (N_44814,N_31804,N_39108);
nor U44815 (N_44815,N_39676,N_37882);
and U44816 (N_44816,N_37707,N_36243);
and U44817 (N_44817,N_39922,N_37552);
or U44818 (N_44818,N_31973,N_38556);
nand U44819 (N_44819,N_35430,N_30060);
or U44820 (N_44820,N_38611,N_31909);
nor U44821 (N_44821,N_35501,N_38886);
and U44822 (N_44822,N_33786,N_32157);
nand U44823 (N_44823,N_38506,N_37481);
nor U44824 (N_44824,N_31348,N_30132);
or U44825 (N_44825,N_31012,N_32799);
nand U44826 (N_44826,N_38182,N_33193);
nor U44827 (N_44827,N_34650,N_33077);
nor U44828 (N_44828,N_38418,N_38646);
xor U44829 (N_44829,N_32769,N_32565);
nor U44830 (N_44830,N_38665,N_38122);
nand U44831 (N_44831,N_30767,N_39160);
or U44832 (N_44832,N_35554,N_37085);
nor U44833 (N_44833,N_39180,N_38606);
or U44834 (N_44834,N_39707,N_35199);
nor U44835 (N_44835,N_39151,N_34080);
or U44836 (N_44836,N_38021,N_35921);
nand U44837 (N_44837,N_37644,N_39665);
and U44838 (N_44838,N_34125,N_37048);
xnor U44839 (N_44839,N_31003,N_33230);
or U44840 (N_44840,N_30530,N_30067);
nor U44841 (N_44841,N_30229,N_32369);
nor U44842 (N_44842,N_32480,N_36224);
nor U44843 (N_44843,N_35640,N_37027);
or U44844 (N_44844,N_39828,N_32823);
xor U44845 (N_44845,N_33511,N_37716);
nand U44846 (N_44846,N_37541,N_34442);
nand U44847 (N_44847,N_30425,N_37025);
nand U44848 (N_44848,N_32203,N_32619);
nor U44849 (N_44849,N_33635,N_36531);
or U44850 (N_44850,N_34362,N_31031);
and U44851 (N_44851,N_33578,N_33051);
nor U44852 (N_44852,N_39779,N_33692);
nor U44853 (N_44853,N_35644,N_35678);
nor U44854 (N_44854,N_31968,N_35614);
and U44855 (N_44855,N_30408,N_32977);
and U44856 (N_44856,N_37827,N_31144);
nor U44857 (N_44857,N_35595,N_34799);
or U44858 (N_44858,N_34792,N_34629);
nor U44859 (N_44859,N_33642,N_34433);
nor U44860 (N_44860,N_32717,N_31403);
nor U44861 (N_44861,N_36011,N_31143);
or U44862 (N_44862,N_38729,N_33674);
and U44863 (N_44863,N_32354,N_32530);
xor U44864 (N_44864,N_34008,N_35435);
xnor U44865 (N_44865,N_33769,N_37647);
xor U44866 (N_44866,N_33153,N_39931);
and U44867 (N_44867,N_35804,N_34902);
nor U44868 (N_44868,N_36810,N_36988);
xnor U44869 (N_44869,N_31786,N_33463);
nand U44870 (N_44870,N_31431,N_34142);
nand U44871 (N_44871,N_36336,N_30422);
nor U44872 (N_44872,N_35856,N_39568);
nor U44873 (N_44873,N_37447,N_34875);
xor U44874 (N_44874,N_30996,N_36932);
nor U44875 (N_44875,N_39910,N_36540);
nand U44876 (N_44876,N_31410,N_35074);
nor U44877 (N_44877,N_36419,N_32315);
and U44878 (N_44878,N_36969,N_34861);
or U44879 (N_44879,N_36759,N_38715);
and U44880 (N_44880,N_36928,N_32036);
or U44881 (N_44881,N_30784,N_35127);
xor U44882 (N_44882,N_38027,N_36094);
and U44883 (N_44883,N_38354,N_35960);
nor U44884 (N_44884,N_35862,N_34984);
and U44885 (N_44885,N_37028,N_30424);
or U44886 (N_44886,N_30152,N_37330);
or U44887 (N_44887,N_38149,N_36523);
nand U44888 (N_44888,N_38724,N_37186);
and U44889 (N_44889,N_33705,N_32253);
or U44890 (N_44890,N_39253,N_37674);
and U44891 (N_44891,N_35031,N_39385);
or U44892 (N_44892,N_34227,N_37719);
nor U44893 (N_44893,N_31862,N_32659);
and U44894 (N_44894,N_32739,N_37813);
nand U44895 (N_44895,N_33259,N_33967);
and U44896 (N_44896,N_31135,N_39429);
nor U44897 (N_44897,N_38597,N_33277);
or U44898 (N_44898,N_35466,N_30063);
nand U44899 (N_44899,N_39428,N_36973);
and U44900 (N_44900,N_34781,N_34666);
nand U44901 (N_44901,N_30068,N_34226);
nor U44902 (N_44902,N_39519,N_35811);
and U44903 (N_44903,N_37055,N_39011);
or U44904 (N_44904,N_32108,N_35249);
and U44905 (N_44905,N_30292,N_33382);
nor U44906 (N_44906,N_34873,N_36459);
and U44907 (N_44907,N_37758,N_32311);
nand U44908 (N_44908,N_33041,N_31155);
or U44909 (N_44909,N_32623,N_35219);
or U44910 (N_44910,N_33863,N_30794);
nor U44911 (N_44911,N_31463,N_31375);
or U44912 (N_44912,N_37735,N_34946);
and U44913 (N_44913,N_30042,N_35631);
and U44914 (N_44914,N_35968,N_36257);
or U44915 (N_44915,N_36237,N_38944);
nor U44916 (N_44916,N_31226,N_32122);
and U44917 (N_44917,N_30855,N_30798);
or U44918 (N_44918,N_38929,N_35218);
nand U44919 (N_44919,N_32615,N_35666);
or U44920 (N_44920,N_35190,N_33847);
and U44921 (N_44921,N_35361,N_30199);
nor U44922 (N_44922,N_37324,N_35087);
or U44923 (N_44923,N_35969,N_36576);
or U44924 (N_44924,N_36535,N_32546);
and U44925 (N_44925,N_31085,N_34801);
nor U44926 (N_44926,N_38135,N_37279);
and U44927 (N_44927,N_30546,N_35809);
xor U44928 (N_44928,N_38750,N_35047);
xor U44929 (N_44929,N_39409,N_39236);
nor U44930 (N_44930,N_31071,N_30618);
or U44931 (N_44931,N_32220,N_33190);
nand U44932 (N_44932,N_31175,N_33953);
xor U44933 (N_44933,N_35144,N_39635);
or U44934 (N_44934,N_32985,N_33598);
and U44935 (N_44935,N_35497,N_33335);
or U44936 (N_44936,N_32401,N_34093);
nor U44937 (N_44937,N_30350,N_31971);
and U44938 (N_44938,N_31486,N_35406);
nor U44939 (N_44939,N_31663,N_36536);
and U44940 (N_44940,N_35663,N_38377);
nand U44941 (N_44941,N_32834,N_38891);
nor U44942 (N_44942,N_36190,N_30479);
and U44943 (N_44943,N_31088,N_33799);
xnor U44944 (N_44944,N_30208,N_31298);
and U44945 (N_44945,N_37006,N_30472);
or U44946 (N_44946,N_32006,N_37966);
xnor U44947 (N_44947,N_30376,N_38615);
nand U44948 (N_44948,N_34392,N_34882);
nand U44949 (N_44949,N_38690,N_37406);
nor U44950 (N_44950,N_33613,N_31540);
nand U44951 (N_44951,N_31064,N_36205);
or U44952 (N_44952,N_36564,N_36436);
xnor U44953 (N_44953,N_35791,N_37955);
and U44954 (N_44954,N_36861,N_31847);
nor U44955 (N_44955,N_31028,N_37510);
or U44956 (N_44956,N_32807,N_37046);
nand U44957 (N_44957,N_39227,N_31368);
nor U44958 (N_44958,N_35020,N_36228);
or U44959 (N_44959,N_36013,N_33657);
or U44960 (N_44960,N_37320,N_31316);
and U44961 (N_44961,N_37138,N_34968);
or U44962 (N_44962,N_31021,N_30291);
and U44963 (N_44963,N_36724,N_34516);
nor U44964 (N_44964,N_35519,N_30108);
and U44965 (N_44965,N_37736,N_39339);
and U44966 (N_44966,N_37113,N_33142);
and U44967 (N_44967,N_39292,N_35697);
nand U44968 (N_44968,N_32523,N_30083);
nor U44969 (N_44969,N_37294,N_35191);
and U44970 (N_44970,N_34796,N_39613);
or U44971 (N_44971,N_30275,N_35150);
or U44972 (N_44972,N_31236,N_33617);
and U44973 (N_44973,N_30088,N_32351);
or U44974 (N_44974,N_33949,N_32982);
nand U44975 (N_44975,N_37848,N_36207);
and U44976 (N_44976,N_32450,N_36356);
or U44977 (N_44977,N_35046,N_31390);
and U44978 (N_44978,N_37807,N_32966);
or U44979 (N_44979,N_32637,N_31171);
nor U44980 (N_44980,N_39677,N_35633);
or U44981 (N_44981,N_37580,N_37723);
nor U44982 (N_44982,N_35819,N_37538);
nor U44983 (N_44983,N_32844,N_33004);
and U44984 (N_44984,N_37189,N_32454);
and U44985 (N_44985,N_34341,N_39040);
and U44986 (N_44986,N_35776,N_32634);
nor U44987 (N_44987,N_33240,N_37074);
and U44988 (N_44988,N_34257,N_30146);
nor U44989 (N_44989,N_36706,N_31168);
and U44990 (N_44990,N_33056,N_34538);
nor U44991 (N_44991,N_32267,N_36330);
or U44992 (N_44992,N_33326,N_33384);
and U44993 (N_44993,N_35622,N_35146);
and U44994 (N_44994,N_37992,N_37231);
and U44995 (N_44995,N_38325,N_38458);
nand U44996 (N_44996,N_33350,N_35543);
or U44997 (N_44997,N_32395,N_30743);
or U44998 (N_44998,N_37839,N_35611);
nor U44999 (N_44999,N_34645,N_34848);
and U45000 (N_45000,N_35983,N_34788);
nand U45001 (N_45001,N_34214,N_37633);
nand U45002 (N_45002,N_33849,N_38819);
nor U45003 (N_45003,N_38390,N_39459);
and U45004 (N_45004,N_38155,N_36500);
or U45005 (N_45005,N_34749,N_37462);
or U45006 (N_45006,N_38980,N_34466);
nand U45007 (N_45007,N_35950,N_38796);
and U45008 (N_45008,N_31042,N_34354);
and U45009 (N_45009,N_32911,N_31111);
xnor U45010 (N_45010,N_31329,N_31025);
or U45011 (N_45011,N_37225,N_39078);
nor U45012 (N_45012,N_39371,N_36878);
or U45013 (N_45013,N_39388,N_30719);
and U45014 (N_45014,N_39807,N_33780);
nor U45015 (N_45015,N_34947,N_30794);
xnor U45016 (N_45016,N_31912,N_38851);
nand U45017 (N_45017,N_33938,N_37865);
nor U45018 (N_45018,N_38163,N_34305);
nor U45019 (N_45019,N_31490,N_34338);
nand U45020 (N_45020,N_37120,N_37861);
or U45021 (N_45021,N_38756,N_30405);
and U45022 (N_45022,N_32102,N_31573);
nand U45023 (N_45023,N_32208,N_38948);
or U45024 (N_45024,N_34224,N_31805);
and U45025 (N_45025,N_31260,N_37930);
or U45026 (N_45026,N_31271,N_33202);
xnor U45027 (N_45027,N_33928,N_38251);
nor U45028 (N_45028,N_32793,N_30431);
nand U45029 (N_45029,N_34225,N_39032);
nor U45030 (N_45030,N_32673,N_37679);
nand U45031 (N_45031,N_37087,N_39729);
nand U45032 (N_45032,N_35118,N_35647);
nor U45033 (N_45033,N_33125,N_36017);
nand U45034 (N_45034,N_30970,N_34191);
nor U45035 (N_45035,N_34628,N_34342);
or U45036 (N_45036,N_31731,N_33815);
and U45037 (N_45037,N_31881,N_32170);
and U45038 (N_45038,N_36191,N_35727);
xor U45039 (N_45039,N_37999,N_39455);
nor U45040 (N_45040,N_32146,N_36064);
and U45041 (N_45041,N_35838,N_34062);
or U45042 (N_45042,N_34662,N_38186);
nand U45043 (N_45043,N_36194,N_39262);
and U45044 (N_45044,N_38148,N_31318);
or U45045 (N_45045,N_36084,N_33203);
xor U45046 (N_45046,N_30995,N_38949);
and U45047 (N_45047,N_30122,N_38816);
or U45048 (N_45048,N_35893,N_30890);
nand U45049 (N_45049,N_36110,N_39193);
nand U45050 (N_45050,N_36484,N_31143);
nand U45051 (N_45051,N_36723,N_35543);
or U45052 (N_45052,N_34402,N_30267);
and U45053 (N_45053,N_39444,N_32490);
nand U45054 (N_45054,N_36408,N_34163);
nand U45055 (N_45055,N_30886,N_39160);
nor U45056 (N_45056,N_37577,N_34047);
and U45057 (N_45057,N_38991,N_39287);
nor U45058 (N_45058,N_39992,N_34859);
xnor U45059 (N_45059,N_39368,N_36075);
nand U45060 (N_45060,N_33978,N_30620);
nor U45061 (N_45061,N_32993,N_34236);
xnor U45062 (N_45062,N_34869,N_39077);
xor U45063 (N_45063,N_30287,N_38637);
xor U45064 (N_45064,N_33018,N_30400);
nor U45065 (N_45065,N_33978,N_30018);
nand U45066 (N_45066,N_31946,N_31099);
nor U45067 (N_45067,N_36487,N_31939);
nand U45068 (N_45068,N_33750,N_38788);
xnor U45069 (N_45069,N_32692,N_34266);
nand U45070 (N_45070,N_37517,N_34657);
nor U45071 (N_45071,N_38987,N_36390);
xnor U45072 (N_45072,N_38684,N_38578);
and U45073 (N_45073,N_37568,N_35410);
and U45074 (N_45074,N_30774,N_33538);
nor U45075 (N_45075,N_36266,N_36468);
or U45076 (N_45076,N_35540,N_36843);
and U45077 (N_45077,N_34497,N_32368);
nor U45078 (N_45078,N_37034,N_38297);
or U45079 (N_45079,N_33997,N_33811);
or U45080 (N_45080,N_35310,N_33472);
xor U45081 (N_45081,N_36223,N_32687);
or U45082 (N_45082,N_39559,N_38164);
nand U45083 (N_45083,N_30775,N_36415);
or U45084 (N_45084,N_31915,N_34504);
nor U45085 (N_45085,N_39605,N_34019);
nor U45086 (N_45086,N_39496,N_36345);
or U45087 (N_45087,N_34737,N_36079);
and U45088 (N_45088,N_31446,N_34016);
xor U45089 (N_45089,N_34209,N_31426);
nor U45090 (N_45090,N_33591,N_32651);
and U45091 (N_45091,N_37536,N_33750);
and U45092 (N_45092,N_33521,N_30871);
nor U45093 (N_45093,N_38512,N_34620);
nor U45094 (N_45094,N_37392,N_37696);
or U45095 (N_45095,N_32273,N_36584);
nand U45096 (N_45096,N_35892,N_38861);
nor U45097 (N_45097,N_36846,N_30009);
nor U45098 (N_45098,N_37196,N_31581);
and U45099 (N_45099,N_30044,N_33931);
nor U45100 (N_45100,N_37748,N_32816);
and U45101 (N_45101,N_30410,N_34547);
nand U45102 (N_45102,N_36104,N_36323);
and U45103 (N_45103,N_34484,N_30870);
nand U45104 (N_45104,N_33861,N_30303);
nand U45105 (N_45105,N_31900,N_32212);
and U45106 (N_45106,N_31745,N_30473);
or U45107 (N_45107,N_36917,N_32443);
nor U45108 (N_45108,N_37016,N_39933);
and U45109 (N_45109,N_31919,N_35825);
nand U45110 (N_45110,N_32013,N_39404);
nor U45111 (N_45111,N_38455,N_34588);
and U45112 (N_45112,N_33385,N_38748);
or U45113 (N_45113,N_32760,N_37458);
nand U45114 (N_45114,N_33945,N_39839);
nand U45115 (N_45115,N_39967,N_37653);
nor U45116 (N_45116,N_32892,N_31503);
nand U45117 (N_45117,N_35724,N_34115);
nor U45118 (N_45118,N_39324,N_37459);
or U45119 (N_45119,N_34716,N_33178);
nor U45120 (N_45120,N_31654,N_32798);
nand U45121 (N_45121,N_35403,N_37749);
or U45122 (N_45122,N_35834,N_36669);
nor U45123 (N_45123,N_37114,N_38929);
or U45124 (N_45124,N_32541,N_38383);
nand U45125 (N_45125,N_32756,N_37575);
and U45126 (N_45126,N_38098,N_36044);
and U45127 (N_45127,N_33977,N_36168);
or U45128 (N_45128,N_31788,N_34313);
nand U45129 (N_45129,N_31896,N_32544);
nor U45130 (N_45130,N_36489,N_33462);
and U45131 (N_45131,N_33180,N_36280);
and U45132 (N_45132,N_32835,N_30716);
nand U45133 (N_45133,N_39698,N_39161);
nor U45134 (N_45134,N_38098,N_31289);
nor U45135 (N_45135,N_34277,N_31082);
or U45136 (N_45136,N_32252,N_32011);
nand U45137 (N_45137,N_34333,N_39971);
or U45138 (N_45138,N_33322,N_38830);
nor U45139 (N_45139,N_35439,N_33104);
and U45140 (N_45140,N_36807,N_32913);
or U45141 (N_45141,N_35991,N_38383);
nor U45142 (N_45142,N_37172,N_35385);
and U45143 (N_45143,N_33212,N_33079);
nand U45144 (N_45144,N_37986,N_37749);
or U45145 (N_45145,N_38341,N_38711);
nor U45146 (N_45146,N_30026,N_34618);
or U45147 (N_45147,N_31564,N_31908);
nor U45148 (N_45148,N_35244,N_35635);
nor U45149 (N_45149,N_33964,N_33141);
nor U45150 (N_45150,N_34061,N_38861);
and U45151 (N_45151,N_37560,N_35316);
nor U45152 (N_45152,N_37135,N_35300);
nor U45153 (N_45153,N_35759,N_37633);
and U45154 (N_45154,N_34273,N_34317);
xor U45155 (N_45155,N_39558,N_30606);
nor U45156 (N_45156,N_34354,N_38819);
and U45157 (N_45157,N_37034,N_38576);
nand U45158 (N_45158,N_34546,N_36121);
and U45159 (N_45159,N_31509,N_33761);
or U45160 (N_45160,N_33393,N_32642);
or U45161 (N_45161,N_35668,N_37958);
nand U45162 (N_45162,N_37378,N_38961);
nor U45163 (N_45163,N_31350,N_37144);
nand U45164 (N_45164,N_33243,N_31258);
nand U45165 (N_45165,N_34365,N_34388);
or U45166 (N_45166,N_36830,N_36258);
or U45167 (N_45167,N_30880,N_30687);
nor U45168 (N_45168,N_34711,N_37263);
and U45169 (N_45169,N_31945,N_37709);
nand U45170 (N_45170,N_32451,N_33357);
and U45171 (N_45171,N_31409,N_34870);
nor U45172 (N_45172,N_30254,N_34240);
nor U45173 (N_45173,N_37375,N_35479);
and U45174 (N_45174,N_37430,N_31891);
nor U45175 (N_45175,N_33993,N_35542);
and U45176 (N_45176,N_32780,N_39824);
or U45177 (N_45177,N_32679,N_39614);
nand U45178 (N_45178,N_32331,N_32587);
nand U45179 (N_45179,N_37391,N_38257);
or U45180 (N_45180,N_36460,N_34826);
xnor U45181 (N_45181,N_33022,N_35635);
and U45182 (N_45182,N_36281,N_31067);
nor U45183 (N_45183,N_32937,N_36935);
and U45184 (N_45184,N_31101,N_34356);
or U45185 (N_45185,N_38663,N_37772);
and U45186 (N_45186,N_36545,N_30212);
nand U45187 (N_45187,N_31750,N_37404);
xor U45188 (N_45188,N_36414,N_35831);
nor U45189 (N_45189,N_35034,N_35063);
or U45190 (N_45190,N_34655,N_36345);
or U45191 (N_45191,N_39497,N_34146);
and U45192 (N_45192,N_32220,N_31899);
nor U45193 (N_45193,N_39813,N_32423);
and U45194 (N_45194,N_37818,N_38791);
and U45195 (N_45195,N_39966,N_34035);
or U45196 (N_45196,N_30830,N_32133);
or U45197 (N_45197,N_35009,N_35876);
and U45198 (N_45198,N_34042,N_37319);
nor U45199 (N_45199,N_38253,N_37390);
or U45200 (N_45200,N_35735,N_30187);
nand U45201 (N_45201,N_32976,N_30490);
nand U45202 (N_45202,N_38048,N_39913);
nand U45203 (N_45203,N_31267,N_33334);
nand U45204 (N_45204,N_39798,N_39810);
nor U45205 (N_45205,N_39887,N_34789);
nand U45206 (N_45206,N_30084,N_35333);
nor U45207 (N_45207,N_30004,N_33765);
or U45208 (N_45208,N_31379,N_39568);
and U45209 (N_45209,N_30113,N_31698);
nor U45210 (N_45210,N_33287,N_31838);
nand U45211 (N_45211,N_34695,N_34987);
nor U45212 (N_45212,N_38963,N_38894);
nor U45213 (N_45213,N_34364,N_30186);
and U45214 (N_45214,N_39443,N_33479);
nand U45215 (N_45215,N_31726,N_35219);
nor U45216 (N_45216,N_39931,N_37127);
or U45217 (N_45217,N_33102,N_34227);
nor U45218 (N_45218,N_36241,N_39995);
or U45219 (N_45219,N_31376,N_30464);
xnor U45220 (N_45220,N_38757,N_38029);
or U45221 (N_45221,N_32616,N_33987);
or U45222 (N_45222,N_36058,N_34183);
or U45223 (N_45223,N_30394,N_37928);
nor U45224 (N_45224,N_30930,N_32064);
nand U45225 (N_45225,N_39871,N_31427);
nand U45226 (N_45226,N_30100,N_39500);
nand U45227 (N_45227,N_37119,N_38304);
nand U45228 (N_45228,N_33480,N_34506);
and U45229 (N_45229,N_35105,N_31943);
nor U45230 (N_45230,N_32173,N_33090);
xor U45231 (N_45231,N_31714,N_34071);
nor U45232 (N_45232,N_30773,N_34109);
nor U45233 (N_45233,N_32804,N_30753);
nand U45234 (N_45234,N_33970,N_33010);
nor U45235 (N_45235,N_38743,N_36461);
or U45236 (N_45236,N_31894,N_36237);
nand U45237 (N_45237,N_39538,N_36110);
or U45238 (N_45238,N_32012,N_39817);
nand U45239 (N_45239,N_31217,N_30327);
nand U45240 (N_45240,N_35152,N_31184);
nor U45241 (N_45241,N_38775,N_35590);
nor U45242 (N_45242,N_34648,N_34507);
or U45243 (N_45243,N_38012,N_32732);
nand U45244 (N_45244,N_38662,N_36534);
and U45245 (N_45245,N_31241,N_30077);
xor U45246 (N_45246,N_34019,N_32149);
and U45247 (N_45247,N_31062,N_38238);
nand U45248 (N_45248,N_38736,N_35873);
and U45249 (N_45249,N_33729,N_36404);
or U45250 (N_45250,N_35928,N_33494);
or U45251 (N_45251,N_38828,N_39063);
and U45252 (N_45252,N_35281,N_30468);
or U45253 (N_45253,N_32771,N_33158);
nor U45254 (N_45254,N_39637,N_35965);
or U45255 (N_45255,N_34663,N_36646);
nor U45256 (N_45256,N_39571,N_31159);
and U45257 (N_45257,N_38814,N_32044);
and U45258 (N_45258,N_38351,N_31082);
and U45259 (N_45259,N_31224,N_35100);
nor U45260 (N_45260,N_38519,N_37180);
or U45261 (N_45261,N_33847,N_32003);
and U45262 (N_45262,N_31720,N_36660);
and U45263 (N_45263,N_34558,N_34618);
nor U45264 (N_45264,N_31602,N_35894);
or U45265 (N_45265,N_38818,N_32868);
or U45266 (N_45266,N_37674,N_33349);
and U45267 (N_45267,N_33904,N_37541);
and U45268 (N_45268,N_31778,N_36119);
nor U45269 (N_45269,N_35074,N_34226);
and U45270 (N_45270,N_33065,N_35303);
or U45271 (N_45271,N_32174,N_31374);
and U45272 (N_45272,N_30033,N_39389);
nand U45273 (N_45273,N_33450,N_37613);
nand U45274 (N_45274,N_35264,N_36334);
and U45275 (N_45275,N_34409,N_30474);
or U45276 (N_45276,N_34973,N_30011);
and U45277 (N_45277,N_34226,N_37701);
and U45278 (N_45278,N_34977,N_33613);
nand U45279 (N_45279,N_36730,N_37932);
xnor U45280 (N_45280,N_34139,N_34862);
nor U45281 (N_45281,N_33713,N_33142);
xnor U45282 (N_45282,N_35512,N_37258);
and U45283 (N_45283,N_31878,N_37009);
nand U45284 (N_45284,N_31310,N_30004);
or U45285 (N_45285,N_37715,N_35218);
and U45286 (N_45286,N_37672,N_37012);
nand U45287 (N_45287,N_30460,N_33145);
nor U45288 (N_45288,N_38743,N_33130);
and U45289 (N_45289,N_37611,N_32472);
xor U45290 (N_45290,N_34552,N_31673);
nand U45291 (N_45291,N_35050,N_30134);
nand U45292 (N_45292,N_38483,N_39454);
xnor U45293 (N_45293,N_35206,N_34292);
and U45294 (N_45294,N_30209,N_37522);
or U45295 (N_45295,N_37276,N_35768);
nor U45296 (N_45296,N_37985,N_31077);
nand U45297 (N_45297,N_33195,N_34082);
and U45298 (N_45298,N_32629,N_35927);
or U45299 (N_45299,N_34629,N_33684);
nor U45300 (N_45300,N_33188,N_30039);
xor U45301 (N_45301,N_34976,N_38409);
nor U45302 (N_45302,N_36356,N_35593);
and U45303 (N_45303,N_32646,N_36384);
nand U45304 (N_45304,N_38202,N_35325);
nor U45305 (N_45305,N_30706,N_36348);
nor U45306 (N_45306,N_39632,N_34191);
nand U45307 (N_45307,N_31289,N_32092);
nand U45308 (N_45308,N_32516,N_36445);
xnor U45309 (N_45309,N_39643,N_36720);
nor U45310 (N_45310,N_39645,N_33978);
or U45311 (N_45311,N_30297,N_38687);
or U45312 (N_45312,N_35039,N_38427);
nand U45313 (N_45313,N_33057,N_35836);
and U45314 (N_45314,N_33959,N_35148);
and U45315 (N_45315,N_36974,N_32518);
xnor U45316 (N_45316,N_31553,N_33203);
and U45317 (N_45317,N_34725,N_36938);
and U45318 (N_45318,N_37706,N_37070);
nor U45319 (N_45319,N_39097,N_32115);
or U45320 (N_45320,N_30492,N_30663);
or U45321 (N_45321,N_30763,N_38678);
and U45322 (N_45322,N_32228,N_30301);
xnor U45323 (N_45323,N_37810,N_30420);
nor U45324 (N_45324,N_31283,N_32787);
nand U45325 (N_45325,N_30367,N_39381);
nor U45326 (N_45326,N_37357,N_35673);
or U45327 (N_45327,N_35604,N_30013);
and U45328 (N_45328,N_30643,N_31833);
and U45329 (N_45329,N_37935,N_32233);
and U45330 (N_45330,N_39020,N_35632);
or U45331 (N_45331,N_39923,N_39704);
nor U45332 (N_45332,N_37869,N_36053);
or U45333 (N_45333,N_32413,N_31475);
and U45334 (N_45334,N_38778,N_34261);
and U45335 (N_45335,N_37158,N_35401);
or U45336 (N_45336,N_39083,N_32407);
or U45337 (N_45337,N_37712,N_37366);
nand U45338 (N_45338,N_35479,N_33919);
nor U45339 (N_45339,N_39925,N_39337);
nor U45340 (N_45340,N_39908,N_30425);
nand U45341 (N_45341,N_32894,N_36421);
and U45342 (N_45342,N_32301,N_31101);
or U45343 (N_45343,N_30733,N_38902);
or U45344 (N_45344,N_37845,N_36758);
or U45345 (N_45345,N_33755,N_36460);
xor U45346 (N_45346,N_35333,N_31105);
nand U45347 (N_45347,N_33866,N_35470);
or U45348 (N_45348,N_36373,N_39809);
or U45349 (N_45349,N_33886,N_39499);
nor U45350 (N_45350,N_34278,N_34053);
and U45351 (N_45351,N_39389,N_37117);
or U45352 (N_45352,N_32391,N_37433);
nor U45353 (N_45353,N_37519,N_32208);
and U45354 (N_45354,N_39784,N_36280);
or U45355 (N_45355,N_35287,N_38789);
nor U45356 (N_45356,N_34069,N_35623);
nor U45357 (N_45357,N_31638,N_34260);
and U45358 (N_45358,N_39116,N_38885);
nor U45359 (N_45359,N_34624,N_33892);
xor U45360 (N_45360,N_30448,N_30994);
nor U45361 (N_45361,N_38148,N_34183);
nor U45362 (N_45362,N_35695,N_38812);
or U45363 (N_45363,N_37993,N_38003);
nor U45364 (N_45364,N_33931,N_34046);
nor U45365 (N_45365,N_38514,N_38918);
nand U45366 (N_45366,N_36505,N_31216);
nand U45367 (N_45367,N_35059,N_38747);
nor U45368 (N_45368,N_38768,N_34248);
nand U45369 (N_45369,N_31186,N_34943);
and U45370 (N_45370,N_38228,N_33625);
or U45371 (N_45371,N_35653,N_37373);
nand U45372 (N_45372,N_34295,N_37244);
or U45373 (N_45373,N_34035,N_30164);
xnor U45374 (N_45374,N_38899,N_37082);
nand U45375 (N_45375,N_38232,N_33542);
xnor U45376 (N_45376,N_36675,N_37859);
nand U45377 (N_45377,N_38271,N_38380);
nand U45378 (N_45378,N_34440,N_31887);
xnor U45379 (N_45379,N_31142,N_39450);
nand U45380 (N_45380,N_35266,N_33412);
or U45381 (N_45381,N_31865,N_32310);
nand U45382 (N_45382,N_31009,N_33886);
nand U45383 (N_45383,N_32472,N_39247);
nor U45384 (N_45384,N_31701,N_36611);
nand U45385 (N_45385,N_33187,N_34437);
xnor U45386 (N_45386,N_37366,N_37872);
nor U45387 (N_45387,N_36241,N_36049);
or U45388 (N_45388,N_38250,N_33691);
and U45389 (N_45389,N_33393,N_38401);
and U45390 (N_45390,N_39740,N_39835);
nand U45391 (N_45391,N_31560,N_35042);
nand U45392 (N_45392,N_37558,N_38847);
or U45393 (N_45393,N_32725,N_36163);
xnor U45394 (N_45394,N_32159,N_37679);
nor U45395 (N_45395,N_37929,N_36425);
or U45396 (N_45396,N_31317,N_38776);
nor U45397 (N_45397,N_39123,N_32006);
and U45398 (N_45398,N_36072,N_39732);
nand U45399 (N_45399,N_39762,N_36990);
nand U45400 (N_45400,N_39382,N_35685);
nand U45401 (N_45401,N_33989,N_38493);
and U45402 (N_45402,N_33957,N_31110);
and U45403 (N_45403,N_32831,N_34454);
or U45404 (N_45404,N_35114,N_35330);
and U45405 (N_45405,N_32130,N_35466);
nor U45406 (N_45406,N_33901,N_31768);
or U45407 (N_45407,N_38735,N_31542);
and U45408 (N_45408,N_37298,N_30265);
or U45409 (N_45409,N_38330,N_33287);
nand U45410 (N_45410,N_37970,N_33519);
and U45411 (N_45411,N_31581,N_36012);
nand U45412 (N_45412,N_32481,N_30650);
nand U45413 (N_45413,N_32542,N_37825);
or U45414 (N_45414,N_30194,N_31580);
or U45415 (N_45415,N_30817,N_37016);
and U45416 (N_45416,N_39421,N_34131);
nor U45417 (N_45417,N_33971,N_38199);
nand U45418 (N_45418,N_35670,N_30946);
or U45419 (N_45419,N_31226,N_35210);
or U45420 (N_45420,N_30029,N_32842);
nand U45421 (N_45421,N_39305,N_36773);
nand U45422 (N_45422,N_33412,N_33771);
nor U45423 (N_45423,N_39228,N_37444);
or U45424 (N_45424,N_39351,N_36646);
nor U45425 (N_45425,N_35791,N_35390);
and U45426 (N_45426,N_30718,N_31176);
nand U45427 (N_45427,N_36873,N_30876);
or U45428 (N_45428,N_34327,N_33840);
xor U45429 (N_45429,N_34824,N_37209);
and U45430 (N_45430,N_35160,N_37050);
nand U45431 (N_45431,N_39402,N_34529);
and U45432 (N_45432,N_36176,N_36560);
and U45433 (N_45433,N_37114,N_35270);
nor U45434 (N_45434,N_33700,N_32939);
nor U45435 (N_45435,N_31072,N_35267);
nand U45436 (N_45436,N_31430,N_37699);
or U45437 (N_45437,N_32114,N_33832);
and U45438 (N_45438,N_38462,N_38234);
nand U45439 (N_45439,N_37783,N_32757);
nand U45440 (N_45440,N_36485,N_32763);
nor U45441 (N_45441,N_32374,N_36781);
nor U45442 (N_45442,N_35998,N_32813);
or U45443 (N_45443,N_33484,N_34872);
nand U45444 (N_45444,N_36010,N_36959);
or U45445 (N_45445,N_36641,N_31403);
nand U45446 (N_45446,N_32222,N_38719);
xor U45447 (N_45447,N_35909,N_36088);
or U45448 (N_45448,N_36535,N_37591);
nand U45449 (N_45449,N_39409,N_32016);
and U45450 (N_45450,N_35827,N_31205);
nand U45451 (N_45451,N_38085,N_38523);
nor U45452 (N_45452,N_30400,N_36471);
and U45453 (N_45453,N_35725,N_37614);
and U45454 (N_45454,N_32973,N_31413);
or U45455 (N_45455,N_36460,N_31337);
nor U45456 (N_45456,N_33079,N_38612);
nand U45457 (N_45457,N_39094,N_39783);
and U45458 (N_45458,N_38995,N_32267);
or U45459 (N_45459,N_33318,N_34078);
nand U45460 (N_45460,N_37093,N_33470);
nand U45461 (N_45461,N_33987,N_32678);
nand U45462 (N_45462,N_39847,N_34162);
nand U45463 (N_45463,N_38739,N_30644);
and U45464 (N_45464,N_33095,N_39927);
nand U45465 (N_45465,N_35008,N_34771);
nor U45466 (N_45466,N_31760,N_33723);
nand U45467 (N_45467,N_34593,N_33862);
xor U45468 (N_45468,N_34387,N_38390);
and U45469 (N_45469,N_39353,N_30128);
nor U45470 (N_45470,N_39969,N_35290);
nand U45471 (N_45471,N_39700,N_39206);
nor U45472 (N_45472,N_34123,N_34449);
nand U45473 (N_45473,N_35016,N_39312);
nand U45474 (N_45474,N_33115,N_33137);
nor U45475 (N_45475,N_38832,N_34264);
xnor U45476 (N_45476,N_31538,N_30325);
and U45477 (N_45477,N_31618,N_36597);
and U45478 (N_45478,N_39265,N_37563);
nor U45479 (N_45479,N_36958,N_31308);
or U45480 (N_45480,N_31008,N_32655);
xor U45481 (N_45481,N_37349,N_31063);
nor U45482 (N_45482,N_38717,N_35306);
or U45483 (N_45483,N_31718,N_36736);
nor U45484 (N_45484,N_38974,N_33171);
nand U45485 (N_45485,N_30328,N_32142);
xnor U45486 (N_45486,N_37547,N_33831);
and U45487 (N_45487,N_35410,N_33220);
nor U45488 (N_45488,N_38841,N_35414);
and U45489 (N_45489,N_36491,N_34634);
and U45490 (N_45490,N_38587,N_33484);
xor U45491 (N_45491,N_30637,N_39810);
and U45492 (N_45492,N_35815,N_37540);
or U45493 (N_45493,N_38877,N_37715);
xnor U45494 (N_45494,N_35490,N_36513);
nor U45495 (N_45495,N_36751,N_31130);
and U45496 (N_45496,N_31678,N_39971);
nor U45497 (N_45497,N_32633,N_35067);
nor U45498 (N_45498,N_39498,N_37129);
xor U45499 (N_45499,N_37580,N_37158);
and U45500 (N_45500,N_33826,N_39775);
or U45501 (N_45501,N_33064,N_35729);
nor U45502 (N_45502,N_31853,N_31561);
nor U45503 (N_45503,N_34832,N_38358);
and U45504 (N_45504,N_39076,N_30535);
or U45505 (N_45505,N_38200,N_33422);
nor U45506 (N_45506,N_34639,N_30882);
xnor U45507 (N_45507,N_32599,N_31387);
or U45508 (N_45508,N_33223,N_32880);
nor U45509 (N_45509,N_33692,N_37618);
or U45510 (N_45510,N_37561,N_34767);
or U45511 (N_45511,N_35476,N_30240);
and U45512 (N_45512,N_34417,N_38624);
or U45513 (N_45513,N_39028,N_33436);
nor U45514 (N_45514,N_33929,N_34394);
or U45515 (N_45515,N_32883,N_32005);
or U45516 (N_45516,N_37415,N_38623);
nand U45517 (N_45517,N_30593,N_33113);
and U45518 (N_45518,N_33975,N_33789);
or U45519 (N_45519,N_38255,N_32306);
or U45520 (N_45520,N_36955,N_33364);
xnor U45521 (N_45521,N_30452,N_35158);
or U45522 (N_45522,N_32915,N_30470);
nor U45523 (N_45523,N_38561,N_35344);
and U45524 (N_45524,N_32487,N_33782);
and U45525 (N_45525,N_39037,N_31614);
nor U45526 (N_45526,N_30439,N_30205);
nand U45527 (N_45527,N_35840,N_36858);
or U45528 (N_45528,N_38944,N_33204);
nand U45529 (N_45529,N_31541,N_37530);
or U45530 (N_45530,N_34089,N_39249);
or U45531 (N_45531,N_37839,N_30833);
xor U45532 (N_45532,N_33449,N_30926);
and U45533 (N_45533,N_34145,N_30546);
nor U45534 (N_45534,N_36042,N_31496);
or U45535 (N_45535,N_32354,N_33225);
nand U45536 (N_45536,N_30824,N_39564);
or U45537 (N_45537,N_31443,N_39127);
and U45538 (N_45538,N_33080,N_35586);
nor U45539 (N_45539,N_31593,N_35738);
nand U45540 (N_45540,N_39388,N_30180);
and U45541 (N_45541,N_38125,N_30304);
or U45542 (N_45542,N_33292,N_30931);
or U45543 (N_45543,N_37568,N_33310);
and U45544 (N_45544,N_33799,N_37059);
nor U45545 (N_45545,N_35891,N_37208);
nand U45546 (N_45546,N_33889,N_36745);
nand U45547 (N_45547,N_32378,N_30081);
or U45548 (N_45548,N_39603,N_37136);
or U45549 (N_45549,N_31277,N_30346);
or U45550 (N_45550,N_39636,N_31720);
or U45551 (N_45551,N_32777,N_36231);
nand U45552 (N_45552,N_37949,N_33329);
and U45553 (N_45553,N_33594,N_38149);
nor U45554 (N_45554,N_35545,N_38101);
nor U45555 (N_45555,N_35995,N_33067);
nor U45556 (N_45556,N_33739,N_39890);
nor U45557 (N_45557,N_35034,N_34907);
nand U45558 (N_45558,N_33163,N_39888);
and U45559 (N_45559,N_35107,N_32557);
or U45560 (N_45560,N_34430,N_38689);
xor U45561 (N_45561,N_39651,N_37397);
nor U45562 (N_45562,N_35460,N_39568);
nor U45563 (N_45563,N_37764,N_39969);
or U45564 (N_45564,N_36875,N_34315);
and U45565 (N_45565,N_33766,N_37341);
nor U45566 (N_45566,N_37342,N_31959);
nor U45567 (N_45567,N_33787,N_34478);
or U45568 (N_45568,N_31086,N_38005);
or U45569 (N_45569,N_34802,N_35167);
or U45570 (N_45570,N_33931,N_38739);
xor U45571 (N_45571,N_32686,N_39163);
nor U45572 (N_45572,N_31372,N_36806);
xnor U45573 (N_45573,N_33244,N_33381);
or U45574 (N_45574,N_31356,N_37018);
xnor U45575 (N_45575,N_33385,N_32606);
xor U45576 (N_45576,N_34018,N_37428);
or U45577 (N_45577,N_35890,N_33292);
or U45578 (N_45578,N_33993,N_35743);
nand U45579 (N_45579,N_30213,N_31560);
and U45580 (N_45580,N_33340,N_32153);
or U45581 (N_45581,N_39562,N_37358);
nand U45582 (N_45582,N_35375,N_31429);
or U45583 (N_45583,N_37517,N_33548);
nand U45584 (N_45584,N_32424,N_37254);
nor U45585 (N_45585,N_35033,N_36472);
nor U45586 (N_45586,N_38786,N_32237);
nand U45587 (N_45587,N_39205,N_33698);
or U45588 (N_45588,N_30879,N_30675);
nor U45589 (N_45589,N_32811,N_31603);
xnor U45590 (N_45590,N_37697,N_33129);
or U45591 (N_45591,N_35302,N_33652);
nor U45592 (N_45592,N_35804,N_34877);
nand U45593 (N_45593,N_30922,N_33036);
or U45594 (N_45594,N_35235,N_33533);
or U45595 (N_45595,N_31164,N_35283);
nor U45596 (N_45596,N_34806,N_33379);
nand U45597 (N_45597,N_35854,N_33824);
and U45598 (N_45598,N_33407,N_32596);
or U45599 (N_45599,N_32868,N_32167);
xor U45600 (N_45600,N_36950,N_39933);
or U45601 (N_45601,N_33224,N_30555);
and U45602 (N_45602,N_33063,N_30545);
and U45603 (N_45603,N_34375,N_31906);
nand U45604 (N_45604,N_30012,N_34237);
and U45605 (N_45605,N_36678,N_36659);
nor U45606 (N_45606,N_30762,N_38802);
and U45607 (N_45607,N_39993,N_34041);
nand U45608 (N_45608,N_35912,N_37406);
nor U45609 (N_45609,N_32631,N_38558);
and U45610 (N_45610,N_39220,N_33110);
xnor U45611 (N_45611,N_30726,N_39222);
xnor U45612 (N_45612,N_33710,N_37890);
or U45613 (N_45613,N_38207,N_38819);
nor U45614 (N_45614,N_34206,N_39856);
nand U45615 (N_45615,N_33846,N_36495);
or U45616 (N_45616,N_37572,N_32559);
or U45617 (N_45617,N_31605,N_38067);
nor U45618 (N_45618,N_32203,N_37601);
and U45619 (N_45619,N_33562,N_33174);
nand U45620 (N_45620,N_30501,N_38241);
nor U45621 (N_45621,N_36253,N_30529);
xor U45622 (N_45622,N_36425,N_37035);
and U45623 (N_45623,N_34255,N_31916);
nor U45624 (N_45624,N_38256,N_37424);
and U45625 (N_45625,N_38596,N_31164);
nor U45626 (N_45626,N_37871,N_32564);
nand U45627 (N_45627,N_31540,N_38219);
nand U45628 (N_45628,N_30368,N_34584);
nand U45629 (N_45629,N_30448,N_38650);
or U45630 (N_45630,N_34084,N_36519);
xnor U45631 (N_45631,N_35253,N_39867);
xnor U45632 (N_45632,N_36909,N_33029);
or U45633 (N_45633,N_30740,N_32077);
or U45634 (N_45634,N_37720,N_35453);
nand U45635 (N_45635,N_32583,N_31359);
or U45636 (N_45636,N_30722,N_30140);
nor U45637 (N_45637,N_36754,N_34497);
nor U45638 (N_45638,N_34078,N_32172);
xor U45639 (N_45639,N_39886,N_38326);
and U45640 (N_45640,N_38072,N_32004);
nor U45641 (N_45641,N_34461,N_37816);
nor U45642 (N_45642,N_34182,N_30060);
nor U45643 (N_45643,N_38427,N_34551);
nand U45644 (N_45644,N_34096,N_33151);
and U45645 (N_45645,N_30320,N_34229);
or U45646 (N_45646,N_35846,N_35148);
nand U45647 (N_45647,N_38892,N_37005);
nand U45648 (N_45648,N_34972,N_36177);
and U45649 (N_45649,N_34440,N_34568);
and U45650 (N_45650,N_39580,N_33465);
xnor U45651 (N_45651,N_34749,N_34894);
and U45652 (N_45652,N_36860,N_34205);
and U45653 (N_45653,N_31158,N_34561);
nor U45654 (N_45654,N_33794,N_34866);
nor U45655 (N_45655,N_34727,N_38877);
nand U45656 (N_45656,N_32859,N_36564);
nand U45657 (N_45657,N_30442,N_39183);
nand U45658 (N_45658,N_35430,N_39094);
nand U45659 (N_45659,N_30125,N_37636);
and U45660 (N_45660,N_37208,N_36673);
nor U45661 (N_45661,N_30694,N_30905);
and U45662 (N_45662,N_37943,N_38941);
xor U45663 (N_45663,N_37490,N_36301);
nor U45664 (N_45664,N_33538,N_38884);
nor U45665 (N_45665,N_32855,N_35844);
and U45666 (N_45666,N_34848,N_35867);
nand U45667 (N_45667,N_33471,N_32856);
nand U45668 (N_45668,N_37758,N_33925);
and U45669 (N_45669,N_36605,N_38230);
or U45670 (N_45670,N_32631,N_33349);
or U45671 (N_45671,N_31334,N_35207);
nand U45672 (N_45672,N_36506,N_39794);
nand U45673 (N_45673,N_39696,N_35879);
or U45674 (N_45674,N_36434,N_34057);
or U45675 (N_45675,N_34757,N_31868);
or U45676 (N_45676,N_34750,N_31309);
nor U45677 (N_45677,N_30943,N_38574);
nor U45678 (N_45678,N_39296,N_32574);
nand U45679 (N_45679,N_38825,N_36276);
or U45680 (N_45680,N_39116,N_31143);
and U45681 (N_45681,N_35606,N_32580);
nor U45682 (N_45682,N_36345,N_34615);
nand U45683 (N_45683,N_39142,N_38493);
nand U45684 (N_45684,N_31627,N_33879);
and U45685 (N_45685,N_39119,N_39107);
and U45686 (N_45686,N_37641,N_31586);
nand U45687 (N_45687,N_37235,N_32170);
nand U45688 (N_45688,N_32809,N_32735);
nor U45689 (N_45689,N_34810,N_35564);
or U45690 (N_45690,N_35758,N_36093);
or U45691 (N_45691,N_31079,N_33778);
nand U45692 (N_45692,N_38418,N_34104);
xor U45693 (N_45693,N_33188,N_30231);
nor U45694 (N_45694,N_30158,N_34106);
and U45695 (N_45695,N_37560,N_31291);
or U45696 (N_45696,N_37033,N_37543);
or U45697 (N_45697,N_32978,N_31457);
and U45698 (N_45698,N_37302,N_31947);
nand U45699 (N_45699,N_34667,N_37083);
nor U45700 (N_45700,N_36936,N_32756);
xor U45701 (N_45701,N_31716,N_37940);
or U45702 (N_45702,N_30278,N_33961);
or U45703 (N_45703,N_39465,N_30930);
and U45704 (N_45704,N_32391,N_33056);
and U45705 (N_45705,N_31449,N_33931);
nor U45706 (N_45706,N_32844,N_30131);
nand U45707 (N_45707,N_34972,N_34702);
and U45708 (N_45708,N_35014,N_32861);
nor U45709 (N_45709,N_38034,N_38512);
nand U45710 (N_45710,N_33396,N_38372);
nand U45711 (N_45711,N_32778,N_36633);
nand U45712 (N_45712,N_32538,N_32490);
nor U45713 (N_45713,N_37663,N_36703);
nor U45714 (N_45714,N_38133,N_38691);
nor U45715 (N_45715,N_31593,N_37266);
or U45716 (N_45716,N_35181,N_30906);
nor U45717 (N_45717,N_39099,N_30467);
nor U45718 (N_45718,N_37252,N_35370);
and U45719 (N_45719,N_31807,N_37837);
nand U45720 (N_45720,N_35459,N_36091);
or U45721 (N_45721,N_39387,N_38535);
xor U45722 (N_45722,N_35685,N_37468);
nand U45723 (N_45723,N_33331,N_39472);
and U45724 (N_45724,N_39831,N_37301);
nand U45725 (N_45725,N_33194,N_34316);
or U45726 (N_45726,N_39886,N_32724);
nand U45727 (N_45727,N_32781,N_33825);
xnor U45728 (N_45728,N_30872,N_36895);
and U45729 (N_45729,N_35565,N_38803);
nand U45730 (N_45730,N_36934,N_33291);
or U45731 (N_45731,N_33918,N_32692);
nor U45732 (N_45732,N_35648,N_30017);
nand U45733 (N_45733,N_38501,N_30541);
or U45734 (N_45734,N_32830,N_38257);
nor U45735 (N_45735,N_32540,N_31717);
nor U45736 (N_45736,N_31299,N_38454);
and U45737 (N_45737,N_33221,N_31355);
xnor U45738 (N_45738,N_39153,N_35726);
or U45739 (N_45739,N_31378,N_32967);
xnor U45740 (N_45740,N_36202,N_32445);
nor U45741 (N_45741,N_30318,N_34604);
or U45742 (N_45742,N_38553,N_38726);
or U45743 (N_45743,N_31487,N_36605);
and U45744 (N_45744,N_31645,N_39915);
nand U45745 (N_45745,N_36093,N_39988);
nand U45746 (N_45746,N_30135,N_32165);
or U45747 (N_45747,N_31636,N_31889);
and U45748 (N_45748,N_39626,N_32892);
nand U45749 (N_45749,N_30981,N_39894);
nor U45750 (N_45750,N_31743,N_39346);
and U45751 (N_45751,N_38200,N_34328);
and U45752 (N_45752,N_35691,N_32537);
and U45753 (N_45753,N_34991,N_34948);
nand U45754 (N_45754,N_37277,N_34713);
nand U45755 (N_45755,N_38473,N_30274);
nand U45756 (N_45756,N_32896,N_36215);
nand U45757 (N_45757,N_37427,N_32346);
or U45758 (N_45758,N_36415,N_31516);
xor U45759 (N_45759,N_35668,N_36134);
xor U45760 (N_45760,N_31741,N_37853);
and U45761 (N_45761,N_38558,N_32113);
and U45762 (N_45762,N_30092,N_31953);
xnor U45763 (N_45763,N_39062,N_34251);
xor U45764 (N_45764,N_39175,N_39410);
nand U45765 (N_45765,N_33067,N_33227);
nand U45766 (N_45766,N_37815,N_33360);
nor U45767 (N_45767,N_30647,N_38923);
nor U45768 (N_45768,N_39719,N_32391);
xor U45769 (N_45769,N_37891,N_35037);
or U45770 (N_45770,N_34304,N_35365);
and U45771 (N_45771,N_30415,N_31805);
and U45772 (N_45772,N_37220,N_33636);
or U45773 (N_45773,N_32972,N_38123);
nand U45774 (N_45774,N_34457,N_38316);
nor U45775 (N_45775,N_39143,N_36490);
and U45776 (N_45776,N_32143,N_31602);
and U45777 (N_45777,N_39149,N_34052);
nor U45778 (N_45778,N_31341,N_31513);
or U45779 (N_45779,N_35737,N_34322);
and U45780 (N_45780,N_32848,N_33576);
nand U45781 (N_45781,N_31351,N_33980);
or U45782 (N_45782,N_37222,N_36302);
or U45783 (N_45783,N_32715,N_39654);
nor U45784 (N_45784,N_34421,N_33989);
nand U45785 (N_45785,N_35815,N_30784);
nand U45786 (N_45786,N_39096,N_30825);
nand U45787 (N_45787,N_38452,N_32312);
nand U45788 (N_45788,N_30621,N_37942);
nand U45789 (N_45789,N_35033,N_38708);
nor U45790 (N_45790,N_39296,N_39169);
or U45791 (N_45791,N_30089,N_36132);
and U45792 (N_45792,N_30375,N_32558);
or U45793 (N_45793,N_35863,N_36230);
nand U45794 (N_45794,N_34801,N_31179);
nand U45795 (N_45795,N_31173,N_36229);
nand U45796 (N_45796,N_33149,N_38416);
nor U45797 (N_45797,N_31028,N_32292);
and U45798 (N_45798,N_33061,N_37599);
nand U45799 (N_45799,N_39338,N_31313);
or U45800 (N_45800,N_30960,N_33574);
or U45801 (N_45801,N_38182,N_34482);
nand U45802 (N_45802,N_31634,N_38260);
or U45803 (N_45803,N_33953,N_36393);
xnor U45804 (N_45804,N_37106,N_30555);
nand U45805 (N_45805,N_30692,N_30316);
and U45806 (N_45806,N_38057,N_36405);
and U45807 (N_45807,N_34329,N_36420);
or U45808 (N_45808,N_32517,N_38760);
nand U45809 (N_45809,N_30257,N_34482);
or U45810 (N_45810,N_30059,N_32218);
xnor U45811 (N_45811,N_39970,N_30638);
nor U45812 (N_45812,N_30222,N_35131);
or U45813 (N_45813,N_39456,N_33481);
or U45814 (N_45814,N_37060,N_36045);
and U45815 (N_45815,N_35958,N_34054);
nor U45816 (N_45816,N_36490,N_37964);
nand U45817 (N_45817,N_39348,N_37636);
nor U45818 (N_45818,N_33886,N_36293);
nor U45819 (N_45819,N_31099,N_36338);
nand U45820 (N_45820,N_32654,N_32964);
nand U45821 (N_45821,N_37014,N_33600);
or U45822 (N_45822,N_34825,N_34549);
nand U45823 (N_45823,N_39367,N_33445);
nor U45824 (N_45824,N_32237,N_37501);
and U45825 (N_45825,N_34848,N_38990);
nand U45826 (N_45826,N_31497,N_31982);
or U45827 (N_45827,N_30987,N_34295);
nand U45828 (N_45828,N_34487,N_34942);
xor U45829 (N_45829,N_30978,N_33008);
and U45830 (N_45830,N_38208,N_37416);
and U45831 (N_45831,N_35794,N_35250);
nor U45832 (N_45832,N_34674,N_38531);
and U45833 (N_45833,N_30737,N_35344);
nor U45834 (N_45834,N_31260,N_30672);
nor U45835 (N_45835,N_33121,N_31933);
xor U45836 (N_45836,N_37199,N_34848);
or U45837 (N_45837,N_33856,N_34726);
nand U45838 (N_45838,N_36803,N_39562);
or U45839 (N_45839,N_37236,N_34665);
or U45840 (N_45840,N_36158,N_38408);
nand U45841 (N_45841,N_34140,N_37343);
nor U45842 (N_45842,N_34387,N_33036);
nor U45843 (N_45843,N_39258,N_34591);
or U45844 (N_45844,N_30133,N_36868);
nand U45845 (N_45845,N_38260,N_38200);
nor U45846 (N_45846,N_33180,N_35215);
nor U45847 (N_45847,N_34315,N_33927);
or U45848 (N_45848,N_30458,N_32698);
or U45849 (N_45849,N_37906,N_32700);
nand U45850 (N_45850,N_39758,N_36944);
nor U45851 (N_45851,N_31089,N_38290);
nor U45852 (N_45852,N_39191,N_36118);
nor U45853 (N_45853,N_38370,N_35454);
nor U45854 (N_45854,N_30595,N_34437);
nor U45855 (N_45855,N_37240,N_30969);
nor U45856 (N_45856,N_30162,N_35691);
or U45857 (N_45857,N_39387,N_32744);
nor U45858 (N_45858,N_31671,N_31006);
and U45859 (N_45859,N_35708,N_33347);
xnor U45860 (N_45860,N_34887,N_32367);
nand U45861 (N_45861,N_35291,N_33477);
and U45862 (N_45862,N_39759,N_32960);
and U45863 (N_45863,N_37714,N_34384);
nand U45864 (N_45864,N_36404,N_30108);
nand U45865 (N_45865,N_37158,N_33432);
xor U45866 (N_45866,N_39966,N_34849);
nand U45867 (N_45867,N_31807,N_30669);
nand U45868 (N_45868,N_36968,N_31007);
xor U45869 (N_45869,N_32693,N_35755);
nor U45870 (N_45870,N_33270,N_33638);
and U45871 (N_45871,N_36314,N_36310);
nand U45872 (N_45872,N_37234,N_32927);
or U45873 (N_45873,N_38535,N_33690);
nand U45874 (N_45874,N_39673,N_32529);
nor U45875 (N_45875,N_39711,N_32780);
nand U45876 (N_45876,N_36842,N_38617);
nor U45877 (N_45877,N_36192,N_34575);
and U45878 (N_45878,N_34781,N_32489);
nor U45879 (N_45879,N_39691,N_31911);
and U45880 (N_45880,N_33273,N_37570);
nor U45881 (N_45881,N_31548,N_31380);
nand U45882 (N_45882,N_38893,N_32132);
and U45883 (N_45883,N_39635,N_37141);
or U45884 (N_45884,N_30227,N_36607);
or U45885 (N_45885,N_31194,N_34587);
nand U45886 (N_45886,N_31582,N_31616);
or U45887 (N_45887,N_36859,N_37037);
and U45888 (N_45888,N_39751,N_39009);
and U45889 (N_45889,N_36349,N_37288);
and U45890 (N_45890,N_37167,N_38863);
nor U45891 (N_45891,N_33645,N_30583);
or U45892 (N_45892,N_32416,N_35819);
nor U45893 (N_45893,N_36718,N_39431);
and U45894 (N_45894,N_38355,N_30183);
nor U45895 (N_45895,N_30225,N_32002);
and U45896 (N_45896,N_34039,N_37283);
nand U45897 (N_45897,N_35514,N_37222);
and U45898 (N_45898,N_31113,N_31157);
or U45899 (N_45899,N_33176,N_30245);
or U45900 (N_45900,N_34824,N_34713);
or U45901 (N_45901,N_30227,N_37213);
and U45902 (N_45902,N_39645,N_35237);
nor U45903 (N_45903,N_32231,N_38980);
nor U45904 (N_45904,N_32683,N_37211);
nand U45905 (N_45905,N_30669,N_34178);
or U45906 (N_45906,N_33954,N_31912);
xnor U45907 (N_45907,N_38052,N_39377);
or U45908 (N_45908,N_39818,N_38647);
nor U45909 (N_45909,N_33240,N_36025);
nor U45910 (N_45910,N_33512,N_32312);
nand U45911 (N_45911,N_36441,N_34268);
or U45912 (N_45912,N_37069,N_33968);
and U45913 (N_45913,N_35089,N_38229);
xor U45914 (N_45914,N_32033,N_37494);
or U45915 (N_45915,N_38448,N_30060);
or U45916 (N_45916,N_30645,N_37474);
and U45917 (N_45917,N_36065,N_38224);
and U45918 (N_45918,N_31026,N_35442);
and U45919 (N_45919,N_39511,N_35334);
nor U45920 (N_45920,N_31689,N_37769);
or U45921 (N_45921,N_35346,N_33579);
nor U45922 (N_45922,N_34586,N_30110);
or U45923 (N_45923,N_34368,N_33999);
xor U45924 (N_45924,N_36231,N_35508);
nor U45925 (N_45925,N_31451,N_30077);
or U45926 (N_45926,N_33539,N_36963);
nor U45927 (N_45927,N_31827,N_39639);
or U45928 (N_45928,N_36335,N_32825);
nand U45929 (N_45929,N_31398,N_30572);
xor U45930 (N_45930,N_39752,N_33445);
xor U45931 (N_45931,N_37955,N_37109);
or U45932 (N_45932,N_35312,N_39760);
and U45933 (N_45933,N_39000,N_36964);
and U45934 (N_45934,N_36083,N_32235);
or U45935 (N_45935,N_32856,N_38407);
and U45936 (N_45936,N_36427,N_31602);
and U45937 (N_45937,N_30861,N_37241);
nor U45938 (N_45938,N_39532,N_31367);
and U45939 (N_45939,N_34406,N_39732);
xor U45940 (N_45940,N_36043,N_30828);
and U45941 (N_45941,N_38331,N_31462);
or U45942 (N_45942,N_36338,N_39027);
and U45943 (N_45943,N_34144,N_35591);
nand U45944 (N_45944,N_33956,N_35012);
nor U45945 (N_45945,N_30799,N_36935);
nor U45946 (N_45946,N_34112,N_37949);
or U45947 (N_45947,N_32880,N_35899);
nor U45948 (N_45948,N_33319,N_32830);
nor U45949 (N_45949,N_39458,N_39159);
xnor U45950 (N_45950,N_35375,N_38542);
nand U45951 (N_45951,N_35591,N_34535);
or U45952 (N_45952,N_31952,N_37673);
nor U45953 (N_45953,N_35764,N_38635);
nor U45954 (N_45954,N_33403,N_30187);
xnor U45955 (N_45955,N_35892,N_36043);
nand U45956 (N_45956,N_36357,N_37693);
or U45957 (N_45957,N_34365,N_37919);
or U45958 (N_45958,N_30795,N_31544);
and U45959 (N_45959,N_30244,N_34462);
or U45960 (N_45960,N_30825,N_32694);
and U45961 (N_45961,N_32403,N_33484);
or U45962 (N_45962,N_31965,N_37839);
and U45963 (N_45963,N_34351,N_33614);
nand U45964 (N_45964,N_34067,N_30598);
or U45965 (N_45965,N_32943,N_36300);
and U45966 (N_45966,N_31657,N_30192);
or U45967 (N_45967,N_35777,N_35590);
or U45968 (N_45968,N_36713,N_37239);
nand U45969 (N_45969,N_39433,N_38627);
xor U45970 (N_45970,N_30768,N_38811);
and U45971 (N_45971,N_37226,N_31653);
nor U45972 (N_45972,N_34710,N_39228);
xnor U45973 (N_45973,N_39023,N_34184);
or U45974 (N_45974,N_35808,N_38469);
or U45975 (N_45975,N_38547,N_35016);
and U45976 (N_45976,N_30153,N_31598);
or U45977 (N_45977,N_35135,N_34626);
nor U45978 (N_45978,N_36334,N_32124);
nor U45979 (N_45979,N_34351,N_35862);
nor U45980 (N_45980,N_33175,N_39380);
or U45981 (N_45981,N_38984,N_30990);
or U45982 (N_45982,N_37123,N_33136);
or U45983 (N_45983,N_37388,N_35861);
nor U45984 (N_45984,N_35004,N_35553);
and U45985 (N_45985,N_32065,N_36755);
or U45986 (N_45986,N_31330,N_34623);
nand U45987 (N_45987,N_38279,N_31975);
nand U45988 (N_45988,N_31907,N_37549);
and U45989 (N_45989,N_30270,N_30255);
or U45990 (N_45990,N_37739,N_30325);
nor U45991 (N_45991,N_33644,N_38510);
or U45992 (N_45992,N_37036,N_30255);
or U45993 (N_45993,N_38170,N_36921);
and U45994 (N_45994,N_36989,N_37242);
nand U45995 (N_45995,N_31755,N_34631);
xor U45996 (N_45996,N_32521,N_34693);
nand U45997 (N_45997,N_31174,N_38884);
nand U45998 (N_45998,N_39803,N_34693);
xnor U45999 (N_45999,N_30437,N_31453);
or U46000 (N_46000,N_34374,N_33532);
xor U46001 (N_46001,N_38931,N_36438);
or U46002 (N_46002,N_32302,N_35540);
nand U46003 (N_46003,N_38550,N_35291);
or U46004 (N_46004,N_34306,N_32816);
and U46005 (N_46005,N_31429,N_32308);
and U46006 (N_46006,N_36905,N_38650);
nor U46007 (N_46007,N_33481,N_34938);
nor U46008 (N_46008,N_32571,N_37717);
nand U46009 (N_46009,N_36753,N_34228);
and U46010 (N_46010,N_39418,N_30423);
nor U46011 (N_46011,N_36171,N_36545);
or U46012 (N_46012,N_31943,N_34198);
or U46013 (N_46013,N_32839,N_32624);
nand U46014 (N_46014,N_39852,N_34359);
and U46015 (N_46015,N_32954,N_37237);
xnor U46016 (N_46016,N_34845,N_39861);
and U46017 (N_46017,N_36836,N_33925);
and U46018 (N_46018,N_35171,N_31346);
nand U46019 (N_46019,N_34293,N_33106);
nor U46020 (N_46020,N_30864,N_31955);
nor U46021 (N_46021,N_32288,N_39595);
and U46022 (N_46022,N_39680,N_37364);
and U46023 (N_46023,N_37984,N_39982);
xnor U46024 (N_46024,N_31821,N_36737);
nor U46025 (N_46025,N_33466,N_34500);
nand U46026 (N_46026,N_35795,N_30417);
nor U46027 (N_46027,N_35935,N_35503);
nor U46028 (N_46028,N_31839,N_31596);
nand U46029 (N_46029,N_31940,N_35616);
xor U46030 (N_46030,N_33108,N_33775);
nor U46031 (N_46031,N_37755,N_37795);
and U46032 (N_46032,N_35556,N_37141);
and U46033 (N_46033,N_38711,N_39644);
nand U46034 (N_46034,N_37797,N_39835);
and U46035 (N_46035,N_31886,N_39152);
xnor U46036 (N_46036,N_31605,N_38650);
and U46037 (N_46037,N_30712,N_38897);
or U46038 (N_46038,N_35498,N_35394);
nor U46039 (N_46039,N_30132,N_39645);
and U46040 (N_46040,N_31217,N_39923);
and U46041 (N_46041,N_32285,N_35390);
and U46042 (N_46042,N_34085,N_38357);
nand U46043 (N_46043,N_36753,N_30292);
nor U46044 (N_46044,N_30584,N_34511);
nor U46045 (N_46045,N_35761,N_37895);
and U46046 (N_46046,N_30580,N_35822);
and U46047 (N_46047,N_34510,N_36100);
nand U46048 (N_46048,N_35580,N_32754);
nand U46049 (N_46049,N_34885,N_37645);
xor U46050 (N_46050,N_31498,N_31768);
or U46051 (N_46051,N_35517,N_32101);
nor U46052 (N_46052,N_35955,N_30875);
nor U46053 (N_46053,N_35836,N_33615);
nand U46054 (N_46054,N_32074,N_33472);
or U46055 (N_46055,N_35589,N_31001);
and U46056 (N_46056,N_32956,N_32914);
and U46057 (N_46057,N_33877,N_35835);
nor U46058 (N_46058,N_30664,N_30947);
and U46059 (N_46059,N_36268,N_38651);
nor U46060 (N_46060,N_36177,N_37164);
nand U46061 (N_46061,N_36454,N_37632);
nand U46062 (N_46062,N_38667,N_32609);
nor U46063 (N_46063,N_30311,N_39453);
and U46064 (N_46064,N_34915,N_35635);
xnor U46065 (N_46065,N_35152,N_31159);
xor U46066 (N_46066,N_33077,N_35813);
and U46067 (N_46067,N_33336,N_36761);
or U46068 (N_46068,N_36800,N_33597);
nand U46069 (N_46069,N_38187,N_38817);
and U46070 (N_46070,N_39960,N_34318);
nand U46071 (N_46071,N_35754,N_36027);
nor U46072 (N_46072,N_33065,N_36097);
or U46073 (N_46073,N_37333,N_33046);
nor U46074 (N_46074,N_30134,N_39426);
or U46075 (N_46075,N_38107,N_32106);
and U46076 (N_46076,N_32872,N_36606);
and U46077 (N_46077,N_34927,N_37703);
or U46078 (N_46078,N_32747,N_33098);
nor U46079 (N_46079,N_38919,N_33144);
nand U46080 (N_46080,N_37769,N_31054);
nor U46081 (N_46081,N_34299,N_32673);
nor U46082 (N_46082,N_36063,N_33325);
nor U46083 (N_46083,N_33173,N_31942);
or U46084 (N_46084,N_30658,N_32144);
xor U46085 (N_46085,N_35928,N_39480);
xor U46086 (N_46086,N_37525,N_33397);
and U46087 (N_46087,N_34157,N_34260);
nor U46088 (N_46088,N_33781,N_31395);
nor U46089 (N_46089,N_32398,N_38181);
or U46090 (N_46090,N_37385,N_30248);
or U46091 (N_46091,N_38527,N_31845);
or U46092 (N_46092,N_38032,N_36490);
nor U46093 (N_46093,N_35206,N_30070);
nor U46094 (N_46094,N_32364,N_39006);
nor U46095 (N_46095,N_38974,N_30375);
nand U46096 (N_46096,N_33688,N_30434);
or U46097 (N_46097,N_38035,N_32896);
nand U46098 (N_46098,N_37334,N_37145);
or U46099 (N_46099,N_37734,N_30595);
nor U46100 (N_46100,N_35938,N_37325);
nor U46101 (N_46101,N_36836,N_33720);
nor U46102 (N_46102,N_34176,N_37755);
nor U46103 (N_46103,N_32065,N_33950);
nor U46104 (N_46104,N_38379,N_35902);
or U46105 (N_46105,N_38084,N_31587);
or U46106 (N_46106,N_31761,N_38071);
nand U46107 (N_46107,N_39328,N_36627);
or U46108 (N_46108,N_34962,N_38895);
nor U46109 (N_46109,N_33194,N_32347);
nand U46110 (N_46110,N_33649,N_35654);
nor U46111 (N_46111,N_39817,N_38625);
nor U46112 (N_46112,N_35105,N_36476);
nand U46113 (N_46113,N_30660,N_35390);
and U46114 (N_46114,N_34331,N_39682);
or U46115 (N_46115,N_39866,N_34796);
nand U46116 (N_46116,N_37341,N_30444);
or U46117 (N_46117,N_36719,N_32257);
nand U46118 (N_46118,N_30402,N_34045);
nand U46119 (N_46119,N_37136,N_38538);
or U46120 (N_46120,N_34555,N_32712);
or U46121 (N_46121,N_30845,N_34074);
or U46122 (N_46122,N_35322,N_32263);
nor U46123 (N_46123,N_30958,N_38122);
nand U46124 (N_46124,N_39043,N_36918);
xor U46125 (N_46125,N_34779,N_36939);
and U46126 (N_46126,N_30981,N_32322);
nor U46127 (N_46127,N_32516,N_38667);
and U46128 (N_46128,N_31591,N_32211);
nor U46129 (N_46129,N_34351,N_32045);
nor U46130 (N_46130,N_39628,N_34880);
xor U46131 (N_46131,N_37285,N_37559);
nand U46132 (N_46132,N_34402,N_34449);
and U46133 (N_46133,N_36813,N_35035);
or U46134 (N_46134,N_36323,N_32290);
nor U46135 (N_46135,N_31305,N_32338);
and U46136 (N_46136,N_30042,N_36131);
or U46137 (N_46137,N_34919,N_39876);
nor U46138 (N_46138,N_39791,N_33859);
or U46139 (N_46139,N_33990,N_33723);
or U46140 (N_46140,N_35895,N_30194);
or U46141 (N_46141,N_35824,N_37982);
and U46142 (N_46142,N_38112,N_34887);
and U46143 (N_46143,N_38318,N_33256);
nand U46144 (N_46144,N_31692,N_39024);
nand U46145 (N_46145,N_34767,N_33299);
nand U46146 (N_46146,N_35374,N_33725);
nor U46147 (N_46147,N_36516,N_39271);
xnor U46148 (N_46148,N_34072,N_30302);
nand U46149 (N_46149,N_30688,N_32575);
and U46150 (N_46150,N_34379,N_38000);
and U46151 (N_46151,N_36435,N_38889);
nor U46152 (N_46152,N_34891,N_37326);
xor U46153 (N_46153,N_31602,N_35807);
and U46154 (N_46154,N_35828,N_31412);
nand U46155 (N_46155,N_36026,N_30156);
nand U46156 (N_46156,N_37958,N_32989);
nand U46157 (N_46157,N_35310,N_32953);
nor U46158 (N_46158,N_33880,N_33674);
nand U46159 (N_46159,N_33044,N_31485);
and U46160 (N_46160,N_38750,N_35233);
or U46161 (N_46161,N_30479,N_36976);
xnor U46162 (N_46162,N_30430,N_38760);
and U46163 (N_46163,N_36631,N_36643);
or U46164 (N_46164,N_33461,N_31926);
nand U46165 (N_46165,N_39128,N_39630);
or U46166 (N_46166,N_31128,N_39970);
or U46167 (N_46167,N_37434,N_31173);
and U46168 (N_46168,N_33681,N_36563);
nor U46169 (N_46169,N_36181,N_32670);
and U46170 (N_46170,N_37304,N_39193);
nor U46171 (N_46171,N_38830,N_32837);
or U46172 (N_46172,N_39712,N_35150);
and U46173 (N_46173,N_31310,N_39099);
xor U46174 (N_46174,N_31344,N_35774);
and U46175 (N_46175,N_33876,N_31989);
xnor U46176 (N_46176,N_30020,N_36989);
or U46177 (N_46177,N_38675,N_33186);
nor U46178 (N_46178,N_35947,N_37936);
and U46179 (N_46179,N_35127,N_39439);
nand U46180 (N_46180,N_33899,N_33404);
xor U46181 (N_46181,N_34943,N_37981);
nand U46182 (N_46182,N_36810,N_35187);
nand U46183 (N_46183,N_31029,N_32224);
nand U46184 (N_46184,N_35121,N_39243);
and U46185 (N_46185,N_30285,N_37223);
and U46186 (N_46186,N_33045,N_32806);
and U46187 (N_46187,N_30171,N_36763);
xnor U46188 (N_46188,N_39926,N_34904);
nand U46189 (N_46189,N_35581,N_37139);
nor U46190 (N_46190,N_33756,N_37498);
or U46191 (N_46191,N_38864,N_33938);
nand U46192 (N_46192,N_38001,N_33256);
nand U46193 (N_46193,N_36860,N_30597);
or U46194 (N_46194,N_35175,N_32747);
nor U46195 (N_46195,N_34695,N_38199);
nand U46196 (N_46196,N_38397,N_36573);
nor U46197 (N_46197,N_34085,N_31500);
nor U46198 (N_46198,N_30395,N_32522);
nor U46199 (N_46199,N_37585,N_33492);
nand U46200 (N_46200,N_36504,N_34580);
or U46201 (N_46201,N_34820,N_34897);
xor U46202 (N_46202,N_37835,N_37741);
and U46203 (N_46203,N_32857,N_37457);
nand U46204 (N_46204,N_35498,N_35728);
and U46205 (N_46205,N_33737,N_36938);
nor U46206 (N_46206,N_30087,N_34193);
nor U46207 (N_46207,N_37663,N_35808);
xor U46208 (N_46208,N_32537,N_39844);
nor U46209 (N_46209,N_32743,N_30987);
xnor U46210 (N_46210,N_30217,N_38015);
xnor U46211 (N_46211,N_31105,N_39680);
xnor U46212 (N_46212,N_36306,N_38370);
nor U46213 (N_46213,N_35167,N_38759);
xor U46214 (N_46214,N_33832,N_36166);
nor U46215 (N_46215,N_35948,N_38215);
and U46216 (N_46216,N_31418,N_36490);
nand U46217 (N_46217,N_37053,N_34366);
and U46218 (N_46218,N_37754,N_37479);
nor U46219 (N_46219,N_31596,N_39922);
and U46220 (N_46220,N_34004,N_34073);
or U46221 (N_46221,N_34379,N_36322);
and U46222 (N_46222,N_30035,N_34121);
or U46223 (N_46223,N_36173,N_37164);
or U46224 (N_46224,N_33075,N_37845);
nand U46225 (N_46225,N_36579,N_38738);
and U46226 (N_46226,N_30391,N_39729);
and U46227 (N_46227,N_34317,N_34209);
nand U46228 (N_46228,N_31264,N_38070);
and U46229 (N_46229,N_32665,N_32967);
nand U46230 (N_46230,N_32561,N_33237);
and U46231 (N_46231,N_36366,N_39890);
nand U46232 (N_46232,N_39193,N_37532);
nor U46233 (N_46233,N_30753,N_33951);
nand U46234 (N_46234,N_38450,N_36216);
nand U46235 (N_46235,N_36184,N_36032);
nor U46236 (N_46236,N_39013,N_38646);
or U46237 (N_46237,N_37208,N_31362);
xor U46238 (N_46238,N_32520,N_32699);
and U46239 (N_46239,N_31802,N_36778);
and U46240 (N_46240,N_37515,N_37873);
and U46241 (N_46241,N_38382,N_32886);
or U46242 (N_46242,N_31067,N_34567);
nand U46243 (N_46243,N_32827,N_30150);
and U46244 (N_46244,N_37789,N_37257);
or U46245 (N_46245,N_38157,N_32222);
nand U46246 (N_46246,N_33857,N_34741);
nand U46247 (N_46247,N_30493,N_30877);
and U46248 (N_46248,N_38257,N_30288);
and U46249 (N_46249,N_36149,N_37593);
nor U46250 (N_46250,N_31410,N_35223);
or U46251 (N_46251,N_37296,N_30819);
nor U46252 (N_46252,N_37726,N_36359);
nand U46253 (N_46253,N_30638,N_36211);
and U46254 (N_46254,N_31867,N_35734);
nand U46255 (N_46255,N_37804,N_39255);
nor U46256 (N_46256,N_34601,N_31894);
nand U46257 (N_46257,N_37080,N_33881);
and U46258 (N_46258,N_33399,N_33488);
nand U46259 (N_46259,N_37695,N_38253);
or U46260 (N_46260,N_34511,N_39011);
nor U46261 (N_46261,N_37801,N_30975);
xor U46262 (N_46262,N_36409,N_32756);
or U46263 (N_46263,N_31150,N_32392);
or U46264 (N_46264,N_32511,N_36892);
and U46265 (N_46265,N_30051,N_39581);
or U46266 (N_46266,N_39037,N_38925);
or U46267 (N_46267,N_34459,N_31359);
nand U46268 (N_46268,N_30773,N_36876);
and U46269 (N_46269,N_32259,N_34410);
xor U46270 (N_46270,N_38854,N_39697);
nand U46271 (N_46271,N_37502,N_35668);
nor U46272 (N_46272,N_38752,N_32532);
nand U46273 (N_46273,N_31225,N_32471);
nor U46274 (N_46274,N_37016,N_34174);
nor U46275 (N_46275,N_36592,N_39650);
or U46276 (N_46276,N_39861,N_36472);
nand U46277 (N_46277,N_33200,N_32500);
nor U46278 (N_46278,N_38633,N_33770);
or U46279 (N_46279,N_33714,N_34319);
nor U46280 (N_46280,N_33170,N_37989);
or U46281 (N_46281,N_32756,N_35983);
nand U46282 (N_46282,N_37263,N_32839);
or U46283 (N_46283,N_36333,N_33944);
nand U46284 (N_46284,N_31148,N_39360);
nor U46285 (N_46285,N_35384,N_34569);
nor U46286 (N_46286,N_34924,N_38906);
or U46287 (N_46287,N_39725,N_39163);
nor U46288 (N_46288,N_34207,N_37872);
and U46289 (N_46289,N_30357,N_31312);
and U46290 (N_46290,N_38802,N_39170);
or U46291 (N_46291,N_32267,N_33058);
and U46292 (N_46292,N_30655,N_39336);
xnor U46293 (N_46293,N_37908,N_35717);
or U46294 (N_46294,N_34110,N_32678);
or U46295 (N_46295,N_33151,N_35865);
nor U46296 (N_46296,N_33383,N_36541);
and U46297 (N_46297,N_31596,N_31285);
nor U46298 (N_46298,N_31680,N_39826);
or U46299 (N_46299,N_30021,N_34297);
nand U46300 (N_46300,N_34712,N_39826);
and U46301 (N_46301,N_37669,N_36834);
and U46302 (N_46302,N_34407,N_34191);
xnor U46303 (N_46303,N_32104,N_30184);
nor U46304 (N_46304,N_31623,N_32233);
and U46305 (N_46305,N_34110,N_37020);
nand U46306 (N_46306,N_33977,N_38765);
nor U46307 (N_46307,N_36373,N_38010);
and U46308 (N_46308,N_34655,N_31679);
or U46309 (N_46309,N_39558,N_33950);
or U46310 (N_46310,N_32458,N_38601);
and U46311 (N_46311,N_36928,N_35316);
and U46312 (N_46312,N_36207,N_35096);
and U46313 (N_46313,N_33528,N_34593);
nand U46314 (N_46314,N_31683,N_30533);
xor U46315 (N_46315,N_35496,N_35456);
nor U46316 (N_46316,N_32679,N_36520);
xor U46317 (N_46317,N_35640,N_38820);
nor U46318 (N_46318,N_32328,N_31626);
nand U46319 (N_46319,N_37419,N_33446);
xnor U46320 (N_46320,N_36629,N_34432);
and U46321 (N_46321,N_36749,N_39915);
xor U46322 (N_46322,N_33556,N_38933);
nor U46323 (N_46323,N_36615,N_36984);
nor U46324 (N_46324,N_37358,N_37916);
and U46325 (N_46325,N_35137,N_30933);
nand U46326 (N_46326,N_33929,N_37184);
nand U46327 (N_46327,N_32955,N_35856);
and U46328 (N_46328,N_35948,N_36786);
xor U46329 (N_46329,N_38006,N_30198);
and U46330 (N_46330,N_36123,N_32803);
or U46331 (N_46331,N_39461,N_33170);
nor U46332 (N_46332,N_32650,N_35533);
nand U46333 (N_46333,N_35340,N_33313);
nand U46334 (N_46334,N_30904,N_36735);
nand U46335 (N_46335,N_37397,N_30392);
nand U46336 (N_46336,N_30476,N_38019);
and U46337 (N_46337,N_35588,N_30541);
and U46338 (N_46338,N_31485,N_39179);
or U46339 (N_46339,N_33514,N_37924);
xnor U46340 (N_46340,N_39307,N_38844);
xnor U46341 (N_46341,N_35426,N_36247);
or U46342 (N_46342,N_37262,N_32995);
nor U46343 (N_46343,N_34729,N_33919);
nand U46344 (N_46344,N_39442,N_37625);
or U46345 (N_46345,N_34526,N_34620);
xnor U46346 (N_46346,N_34373,N_34068);
nand U46347 (N_46347,N_36545,N_37572);
or U46348 (N_46348,N_33522,N_33126);
and U46349 (N_46349,N_34788,N_35447);
or U46350 (N_46350,N_36000,N_36690);
nor U46351 (N_46351,N_38648,N_34290);
xor U46352 (N_46352,N_35409,N_34738);
or U46353 (N_46353,N_33721,N_38934);
nand U46354 (N_46354,N_32848,N_35069);
or U46355 (N_46355,N_38550,N_31029);
and U46356 (N_46356,N_35239,N_32587);
xor U46357 (N_46357,N_37980,N_30063);
nor U46358 (N_46358,N_34167,N_35778);
and U46359 (N_46359,N_32813,N_33072);
nor U46360 (N_46360,N_38600,N_38349);
or U46361 (N_46361,N_39116,N_34398);
and U46362 (N_46362,N_34084,N_31110);
nand U46363 (N_46363,N_38818,N_39797);
and U46364 (N_46364,N_33914,N_34699);
nor U46365 (N_46365,N_38318,N_38231);
or U46366 (N_46366,N_37715,N_38633);
or U46367 (N_46367,N_35382,N_32190);
nand U46368 (N_46368,N_39644,N_38115);
nand U46369 (N_46369,N_32883,N_33222);
xor U46370 (N_46370,N_30180,N_36584);
and U46371 (N_46371,N_35352,N_39812);
nand U46372 (N_46372,N_32795,N_38215);
nand U46373 (N_46373,N_37421,N_31202);
nor U46374 (N_46374,N_30375,N_32756);
or U46375 (N_46375,N_34433,N_36673);
or U46376 (N_46376,N_30981,N_39415);
nand U46377 (N_46377,N_30918,N_38150);
nand U46378 (N_46378,N_32861,N_33609);
and U46379 (N_46379,N_34056,N_39609);
or U46380 (N_46380,N_30736,N_34159);
or U46381 (N_46381,N_38264,N_37896);
and U46382 (N_46382,N_39407,N_36437);
nand U46383 (N_46383,N_30109,N_36684);
and U46384 (N_46384,N_32861,N_37774);
nor U46385 (N_46385,N_37871,N_31112);
nand U46386 (N_46386,N_34754,N_32715);
nand U46387 (N_46387,N_38864,N_37382);
and U46388 (N_46388,N_33226,N_30673);
or U46389 (N_46389,N_33423,N_36298);
nor U46390 (N_46390,N_31725,N_33366);
nand U46391 (N_46391,N_34479,N_32069);
or U46392 (N_46392,N_39110,N_35363);
nor U46393 (N_46393,N_31184,N_33927);
xor U46394 (N_46394,N_31355,N_32128);
nand U46395 (N_46395,N_34202,N_31733);
and U46396 (N_46396,N_30396,N_30546);
xor U46397 (N_46397,N_30520,N_37165);
or U46398 (N_46398,N_31686,N_31257);
nand U46399 (N_46399,N_36663,N_38568);
nand U46400 (N_46400,N_32132,N_37187);
and U46401 (N_46401,N_39557,N_36430);
nor U46402 (N_46402,N_35352,N_38948);
nor U46403 (N_46403,N_38829,N_36046);
and U46404 (N_46404,N_33330,N_32438);
or U46405 (N_46405,N_30543,N_35786);
and U46406 (N_46406,N_38223,N_34288);
and U46407 (N_46407,N_33578,N_34979);
and U46408 (N_46408,N_35740,N_36746);
and U46409 (N_46409,N_37815,N_38498);
nor U46410 (N_46410,N_35245,N_30156);
nand U46411 (N_46411,N_30486,N_36193);
or U46412 (N_46412,N_36219,N_37513);
xor U46413 (N_46413,N_32616,N_31731);
xor U46414 (N_46414,N_31204,N_38596);
and U46415 (N_46415,N_36763,N_32772);
and U46416 (N_46416,N_33801,N_35192);
and U46417 (N_46417,N_36767,N_38062);
or U46418 (N_46418,N_32111,N_39097);
and U46419 (N_46419,N_30418,N_31010);
nor U46420 (N_46420,N_36607,N_34296);
and U46421 (N_46421,N_36814,N_31052);
or U46422 (N_46422,N_30239,N_38262);
and U46423 (N_46423,N_31544,N_34668);
and U46424 (N_46424,N_39530,N_34943);
and U46425 (N_46425,N_30521,N_30201);
nand U46426 (N_46426,N_31422,N_35204);
xor U46427 (N_46427,N_37057,N_33053);
xnor U46428 (N_46428,N_32375,N_36589);
and U46429 (N_46429,N_30231,N_39427);
or U46430 (N_46430,N_33173,N_38511);
nor U46431 (N_46431,N_35975,N_39762);
nand U46432 (N_46432,N_39042,N_32661);
and U46433 (N_46433,N_30362,N_38146);
xnor U46434 (N_46434,N_30855,N_31671);
or U46435 (N_46435,N_35492,N_30801);
and U46436 (N_46436,N_33433,N_34531);
nor U46437 (N_46437,N_37863,N_32732);
or U46438 (N_46438,N_35690,N_31176);
nor U46439 (N_46439,N_36548,N_36925);
or U46440 (N_46440,N_33565,N_37750);
and U46441 (N_46441,N_38721,N_33046);
and U46442 (N_46442,N_39646,N_38134);
nand U46443 (N_46443,N_31369,N_32299);
and U46444 (N_46444,N_30967,N_31252);
xnor U46445 (N_46445,N_39711,N_34125);
nor U46446 (N_46446,N_31033,N_39356);
nor U46447 (N_46447,N_34291,N_32342);
nor U46448 (N_46448,N_33177,N_35047);
nand U46449 (N_46449,N_33307,N_31268);
nand U46450 (N_46450,N_30941,N_39862);
or U46451 (N_46451,N_30810,N_38713);
and U46452 (N_46452,N_39860,N_38054);
or U46453 (N_46453,N_39660,N_34088);
nor U46454 (N_46454,N_37758,N_36684);
or U46455 (N_46455,N_32973,N_37673);
or U46456 (N_46456,N_38194,N_38066);
and U46457 (N_46457,N_38431,N_35872);
or U46458 (N_46458,N_30523,N_36431);
and U46459 (N_46459,N_33944,N_30277);
nor U46460 (N_46460,N_35843,N_39772);
nand U46461 (N_46461,N_32846,N_36534);
or U46462 (N_46462,N_33390,N_34336);
nand U46463 (N_46463,N_38798,N_39087);
xnor U46464 (N_46464,N_36359,N_33110);
xor U46465 (N_46465,N_35026,N_33749);
nor U46466 (N_46466,N_30076,N_39003);
nand U46467 (N_46467,N_36075,N_36196);
nor U46468 (N_46468,N_39783,N_34835);
or U46469 (N_46469,N_30689,N_31538);
and U46470 (N_46470,N_31223,N_37650);
or U46471 (N_46471,N_33299,N_34610);
and U46472 (N_46472,N_38424,N_34670);
nand U46473 (N_46473,N_39118,N_39487);
and U46474 (N_46474,N_37690,N_36549);
or U46475 (N_46475,N_38296,N_34796);
nand U46476 (N_46476,N_39725,N_30579);
or U46477 (N_46477,N_38617,N_36716);
nor U46478 (N_46478,N_32525,N_37357);
or U46479 (N_46479,N_30576,N_34779);
or U46480 (N_46480,N_38853,N_32969);
or U46481 (N_46481,N_30728,N_34574);
nand U46482 (N_46482,N_33322,N_32611);
xnor U46483 (N_46483,N_34059,N_38743);
and U46484 (N_46484,N_32068,N_34124);
nor U46485 (N_46485,N_31430,N_36201);
nand U46486 (N_46486,N_39465,N_35407);
and U46487 (N_46487,N_39043,N_30535);
and U46488 (N_46488,N_33631,N_36797);
and U46489 (N_46489,N_37254,N_34920);
nor U46490 (N_46490,N_39110,N_37617);
nor U46491 (N_46491,N_30348,N_33124);
nand U46492 (N_46492,N_32602,N_31969);
and U46493 (N_46493,N_31015,N_39764);
or U46494 (N_46494,N_31096,N_38647);
nor U46495 (N_46495,N_30043,N_30988);
or U46496 (N_46496,N_31827,N_36682);
nor U46497 (N_46497,N_33835,N_32585);
or U46498 (N_46498,N_32395,N_36337);
and U46499 (N_46499,N_32738,N_38609);
or U46500 (N_46500,N_35435,N_35845);
and U46501 (N_46501,N_35825,N_30637);
or U46502 (N_46502,N_33693,N_37088);
nand U46503 (N_46503,N_33230,N_37625);
nor U46504 (N_46504,N_30904,N_32335);
and U46505 (N_46505,N_33930,N_30389);
and U46506 (N_46506,N_31923,N_38402);
nand U46507 (N_46507,N_32253,N_33852);
or U46508 (N_46508,N_35980,N_30788);
nor U46509 (N_46509,N_31070,N_32176);
nand U46510 (N_46510,N_34145,N_31431);
and U46511 (N_46511,N_39967,N_30487);
and U46512 (N_46512,N_30589,N_33377);
or U46513 (N_46513,N_38128,N_36173);
nor U46514 (N_46514,N_37557,N_37463);
and U46515 (N_46515,N_37680,N_34761);
nand U46516 (N_46516,N_36084,N_38278);
and U46517 (N_46517,N_39216,N_35743);
or U46518 (N_46518,N_38563,N_36563);
nand U46519 (N_46519,N_37910,N_34692);
nand U46520 (N_46520,N_39030,N_36238);
and U46521 (N_46521,N_37289,N_39543);
nand U46522 (N_46522,N_32904,N_37553);
xnor U46523 (N_46523,N_32623,N_35576);
or U46524 (N_46524,N_37929,N_30021);
nand U46525 (N_46525,N_38685,N_35935);
and U46526 (N_46526,N_36149,N_39210);
xnor U46527 (N_46527,N_35786,N_34880);
nor U46528 (N_46528,N_37266,N_38405);
nor U46529 (N_46529,N_36214,N_37185);
and U46530 (N_46530,N_34418,N_39490);
nand U46531 (N_46531,N_30490,N_35371);
and U46532 (N_46532,N_36219,N_30854);
or U46533 (N_46533,N_37334,N_30415);
nand U46534 (N_46534,N_33187,N_31372);
nand U46535 (N_46535,N_33275,N_38650);
or U46536 (N_46536,N_34242,N_38682);
nand U46537 (N_46537,N_35191,N_37384);
nor U46538 (N_46538,N_36215,N_35092);
and U46539 (N_46539,N_33788,N_32330);
and U46540 (N_46540,N_37325,N_30811);
and U46541 (N_46541,N_34863,N_35666);
or U46542 (N_46542,N_32359,N_34437);
nand U46543 (N_46543,N_34339,N_36969);
nor U46544 (N_46544,N_34534,N_34377);
and U46545 (N_46545,N_30221,N_30352);
nand U46546 (N_46546,N_32417,N_39350);
nor U46547 (N_46547,N_32234,N_31488);
or U46548 (N_46548,N_34011,N_33696);
nor U46549 (N_46549,N_34346,N_36524);
or U46550 (N_46550,N_36877,N_39897);
and U46551 (N_46551,N_34207,N_38227);
nand U46552 (N_46552,N_34895,N_36596);
and U46553 (N_46553,N_31364,N_38400);
and U46554 (N_46554,N_34899,N_30101);
nand U46555 (N_46555,N_36839,N_33576);
or U46556 (N_46556,N_30526,N_37113);
and U46557 (N_46557,N_32916,N_39314);
and U46558 (N_46558,N_35037,N_34788);
and U46559 (N_46559,N_33379,N_36039);
nand U46560 (N_46560,N_33464,N_30307);
nor U46561 (N_46561,N_31919,N_32404);
or U46562 (N_46562,N_37107,N_34147);
nand U46563 (N_46563,N_38825,N_35187);
nand U46564 (N_46564,N_34727,N_36325);
and U46565 (N_46565,N_32401,N_37409);
nand U46566 (N_46566,N_39217,N_37803);
and U46567 (N_46567,N_38204,N_31155);
or U46568 (N_46568,N_31736,N_37801);
nand U46569 (N_46569,N_33996,N_39546);
and U46570 (N_46570,N_31231,N_34337);
and U46571 (N_46571,N_38359,N_39425);
xor U46572 (N_46572,N_31263,N_30189);
or U46573 (N_46573,N_30441,N_31179);
and U46574 (N_46574,N_31871,N_32138);
nor U46575 (N_46575,N_32979,N_38326);
nand U46576 (N_46576,N_31377,N_32133);
nand U46577 (N_46577,N_35373,N_33948);
nand U46578 (N_46578,N_34622,N_38033);
nand U46579 (N_46579,N_33047,N_38111);
nor U46580 (N_46580,N_35394,N_33090);
and U46581 (N_46581,N_39124,N_34404);
and U46582 (N_46582,N_32726,N_36958);
or U46583 (N_46583,N_38121,N_31118);
nor U46584 (N_46584,N_39229,N_32645);
or U46585 (N_46585,N_39079,N_34112);
or U46586 (N_46586,N_36052,N_39214);
xor U46587 (N_46587,N_35202,N_35642);
and U46588 (N_46588,N_32112,N_34507);
and U46589 (N_46589,N_35839,N_36481);
or U46590 (N_46590,N_35154,N_34238);
xor U46591 (N_46591,N_35870,N_37488);
nand U46592 (N_46592,N_35890,N_39855);
nor U46593 (N_46593,N_34479,N_38177);
or U46594 (N_46594,N_33659,N_30228);
xnor U46595 (N_46595,N_33375,N_36408);
or U46596 (N_46596,N_31915,N_39502);
nand U46597 (N_46597,N_35866,N_37458);
and U46598 (N_46598,N_35466,N_32434);
and U46599 (N_46599,N_30024,N_37921);
xnor U46600 (N_46600,N_37527,N_38464);
xor U46601 (N_46601,N_39903,N_33128);
and U46602 (N_46602,N_32240,N_34361);
or U46603 (N_46603,N_36790,N_39696);
nand U46604 (N_46604,N_36769,N_31759);
nor U46605 (N_46605,N_36619,N_31736);
and U46606 (N_46606,N_37978,N_30689);
xor U46607 (N_46607,N_34779,N_34631);
or U46608 (N_46608,N_37593,N_30053);
and U46609 (N_46609,N_33180,N_38765);
and U46610 (N_46610,N_39976,N_34785);
nand U46611 (N_46611,N_36804,N_37758);
or U46612 (N_46612,N_32323,N_39351);
or U46613 (N_46613,N_39095,N_39807);
nor U46614 (N_46614,N_35620,N_30751);
nand U46615 (N_46615,N_32440,N_39014);
or U46616 (N_46616,N_34025,N_36086);
and U46617 (N_46617,N_39035,N_38580);
nor U46618 (N_46618,N_33864,N_35988);
and U46619 (N_46619,N_33291,N_35736);
or U46620 (N_46620,N_36224,N_32277);
nand U46621 (N_46621,N_36768,N_38010);
nor U46622 (N_46622,N_35106,N_31234);
nand U46623 (N_46623,N_37470,N_39274);
or U46624 (N_46624,N_34204,N_32281);
nand U46625 (N_46625,N_35170,N_32180);
and U46626 (N_46626,N_36967,N_38240);
nor U46627 (N_46627,N_30439,N_31072);
or U46628 (N_46628,N_37865,N_32273);
or U46629 (N_46629,N_36222,N_30715);
nor U46630 (N_46630,N_34916,N_36783);
and U46631 (N_46631,N_36833,N_32259);
and U46632 (N_46632,N_38182,N_35021);
nor U46633 (N_46633,N_35479,N_34181);
and U46634 (N_46634,N_30733,N_38841);
nor U46635 (N_46635,N_39267,N_30956);
nand U46636 (N_46636,N_36332,N_32546);
and U46637 (N_46637,N_37513,N_38515);
and U46638 (N_46638,N_39012,N_36449);
or U46639 (N_46639,N_39566,N_30654);
nand U46640 (N_46640,N_30770,N_37626);
or U46641 (N_46641,N_32541,N_33047);
nor U46642 (N_46642,N_30720,N_30996);
or U46643 (N_46643,N_39336,N_39340);
nor U46644 (N_46644,N_34554,N_34852);
and U46645 (N_46645,N_39523,N_36566);
nor U46646 (N_46646,N_31681,N_33356);
or U46647 (N_46647,N_34669,N_39992);
or U46648 (N_46648,N_34526,N_39912);
nand U46649 (N_46649,N_38647,N_31027);
and U46650 (N_46650,N_37766,N_32466);
or U46651 (N_46651,N_32883,N_36911);
nor U46652 (N_46652,N_33624,N_36072);
xnor U46653 (N_46653,N_35988,N_30331);
and U46654 (N_46654,N_35289,N_30631);
nor U46655 (N_46655,N_34671,N_35537);
and U46656 (N_46656,N_36661,N_31509);
nor U46657 (N_46657,N_31008,N_33072);
or U46658 (N_46658,N_35731,N_32541);
nor U46659 (N_46659,N_31085,N_34486);
and U46660 (N_46660,N_36133,N_36071);
or U46661 (N_46661,N_34614,N_30106);
or U46662 (N_46662,N_30213,N_32117);
or U46663 (N_46663,N_30992,N_39580);
and U46664 (N_46664,N_32811,N_36209);
nand U46665 (N_46665,N_35684,N_32165);
nand U46666 (N_46666,N_39180,N_33431);
or U46667 (N_46667,N_33512,N_38996);
nor U46668 (N_46668,N_33372,N_32374);
and U46669 (N_46669,N_39889,N_33831);
nand U46670 (N_46670,N_30478,N_30328);
nor U46671 (N_46671,N_30516,N_33347);
nand U46672 (N_46672,N_36740,N_33460);
nor U46673 (N_46673,N_37478,N_39533);
nor U46674 (N_46674,N_35311,N_34320);
xnor U46675 (N_46675,N_32302,N_38707);
or U46676 (N_46676,N_35226,N_34810);
nor U46677 (N_46677,N_35852,N_36003);
nor U46678 (N_46678,N_33700,N_30628);
and U46679 (N_46679,N_38060,N_39644);
or U46680 (N_46680,N_36067,N_37521);
nor U46681 (N_46681,N_38780,N_31856);
nor U46682 (N_46682,N_39042,N_32577);
or U46683 (N_46683,N_39332,N_31402);
or U46684 (N_46684,N_39591,N_32132);
or U46685 (N_46685,N_38206,N_34404);
or U46686 (N_46686,N_35367,N_34845);
nand U46687 (N_46687,N_32153,N_38342);
or U46688 (N_46688,N_30182,N_33423);
nor U46689 (N_46689,N_32620,N_32756);
or U46690 (N_46690,N_33863,N_36508);
xor U46691 (N_46691,N_39714,N_35014);
nor U46692 (N_46692,N_35376,N_34166);
nand U46693 (N_46693,N_32202,N_31934);
or U46694 (N_46694,N_37288,N_33621);
nand U46695 (N_46695,N_33884,N_31541);
xor U46696 (N_46696,N_37506,N_34290);
and U46697 (N_46697,N_35371,N_36672);
nor U46698 (N_46698,N_33450,N_36850);
nor U46699 (N_46699,N_30420,N_32230);
and U46700 (N_46700,N_36505,N_38326);
nor U46701 (N_46701,N_32245,N_33626);
nand U46702 (N_46702,N_38812,N_33481);
and U46703 (N_46703,N_36811,N_39260);
nor U46704 (N_46704,N_37074,N_36972);
or U46705 (N_46705,N_35594,N_32989);
xnor U46706 (N_46706,N_36510,N_38831);
nand U46707 (N_46707,N_30008,N_35909);
nor U46708 (N_46708,N_39017,N_36647);
or U46709 (N_46709,N_37261,N_37807);
nor U46710 (N_46710,N_34625,N_38916);
and U46711 (N_46711,N_35901,N_30475);
xnor U46712 (N_46712,N_35418,N_37266);
or U46713 (N_46713,N_30917,N_35505);
nor U46714 (N_46714,N_30175,N_38002);
and U46715 (N_46715,N_38874,N_39155);
and U46716 (N_46716,N_32859,N_37768);
and U46717 (N_46717,N_39783,N_37884);
or U46718 (N_46718,N_36400,N_37027);
or U46719 (N_46719,N_33894,N_36880);
nand U46720 (N_46720,N_38700,N_30807);
and U46721 (N_46721,N_39922,N_33085);
or U46722 (N_46722,N_33620,N_31817);
xnor U46723 (N_46723,N_38143,N_30433);
nor U46724 (N_46724,N_33820,N_32846);
nor U46725 (N_46725,N_36197,N_34219);
nand U46726 (N_46726,N_31406,N_33165);
and U46727 (N_46727,N_34361,N_39190);
and U46728 (N_46728,N_37260,N_30529);
xor U46729 (N_46729,N_30615,N_38834);
nand U46730 (N_46730,N_36182,N_39996);
nand U46731 (N_46731,N_37704,N_34762);
and U46732 (N_46732,N_34739,N_31285);
nor U46733 (N_46733,N_34112,N_30228);
and U46734 (N_46734,N_32253,N_36500);
and U46735 (N_46735,N_36547,N_35213);
and U46736 (N_46736,N_31800,N_32128);
nor U46737 (N_46737,N_37886,N_36029);
and U46738 (N_46738,N_36598,N_30417);
xnor U46739 (N_46739,N_39091,N_39452);
nor U46740 (N_46740,N_36191,N_35193);
and U46741 (N_46741,N_38276,N_33796);
nor U46742 (N_46742,N_35018,N_34924);
or U46743 (N_46743,N_39402,N_36315);
nand U46744 (N_46744,N_34985,N_36020);
and U46745 (N_46745,N_39361,N_30111);
nand U46746 (N_46746,N_36058,N_38673);
or U46747 (N_46747,N_32869,N_30495);
and U46748 (N_46748,N_38421,N_33131);
xnor U46749 (N_46749,N_33686,N_35614);
nand U46750 (N_46750,N_33568,N_36389);
or U46751 (N_46751,N_33132,N_38162);
xor U46752 (N_46752,N_31430,N_37285);
nand U46753 (N_46753,N_38297,N_33559);
or U46754 (N_46754,N_32440,N_32308);
or U46755 (N_46755,N_35861,N_36083);
nor U46756 (N_46756,N_38704,N_39928);
or U46757 (N_46757,N_34732,N_38253);
nor U46758 (N_46758,N_36784,N_33084);
and U46759 (N_46759,N_35964,N_30338);
and U46760 (N_46760,N_31155,N_32269);
nor U46761 (N_46761,N_38785,N_37941);
or U46762 (N_46762,N_33840,N_32877);
nor U46763 (N_46763,N_33547,N_37235);
nor U46764 (N_46764,N_35273,N_33030);
or U46765 (N_46765,N_37821,N_34421);
and U46766 (N_46766,N_35364,N_31672);
nor U46767 (N_46767,N_36523,N_39901);
and U46768 (N_46768,N_31518,N_34933);
nor U46769 (N_46769,N_35507,N_31855);
or U46770 (N_46770,N_34683,N_32679);
nor U46771 (N_46771,N_33558,N_34051);
or U46772 (N_46772,N_35610,N_38299);
nor U46773 (N_46773,N_32410,N_34547);
or U46774 (N_46774,N_34325,N_37867);
or U46775 (N_46775,N_32595,N_38383);
or U46776 (N_46776,N_30358,N_32305);
xnor U46777 (N_46777,N_39869,N_36012);
nor U46778 (N_46778,N_31091,N_30868);
nor U46779 (N_46779,N_35529,N_36724);
nand U46780 (N_46780,N_38108,N_38934);
or U46781 (N_46781,N_36180,N_30798);
nor U46782 (N_46782,N_32568,N_33968);
and U46783 (N_46783,N_31689,N_33274);
nand U46784 (N_46784,N_33911,N_35598);
and U46785 (N_46785,N_31997,N_32635);
or U46786 (N_46786,N_34442,N_34505);
nor U46787 (N_46787,N_32213,N_39918);
nor U46788 (N_46788,N_35843,N_34053);
nor U46789 (N_46789,N_36780,N_33700);
nor U46790 (N_46790,N_36087,N_31734);
xnor U46791 (N_46791,N_32647,N_30147);
nand U46792 (N_46792,N_37627,N_35288);
nor U46793 (N_46793,N_35811,N_38367);
nand U46794 (N_46794,N_32139,N_33697);
and U46795 (N_46795,N_34852,N_37469);
and U46796 (N_46796,N_30027,N_37130);
nand U46797 (N_46797,N_37361,N_39027);
or U46798 (N_46798,N_37964,N_30052);
and U46799 (N_46799,N_33522,N_37923);
nor U46800 (N_46800,N_31868,N_36281);
xor U46801 (N_46801,N_33294,N_37140);
and U46802 (N_46802,N_36796,N_35824);
or U46803 (N_46803,N_33440,N_37236);
nor U46804 (N_46804,N_31393,N_33957);
nand U46805 (N_46805,N_37625,N_38028);
nor U46806 (N_46806,N_35342,N_39492);
or U46807 (N_46807,N_32102,N_33226);
nor U46808 (N_46808,N_34329,N_36032);
and U46809 (N_46809,N_32795,N_36624);
xor U46810 (N_46810,N_37521,N_33227);
nor U46811 (N_46811,N_30900,N_35825);
or U46812 (N_46812,N_37638,N_32481);
nand U46813 (N_46813,N_36025,N_34396);
or U46814 (N_46814,N_33597,N_30908);
nand U46815 (N_46815,N_39613,N_30211);
nand U46816 (N_46816,N_34276,N_30732);
and U46817 (N_46817,N_33164,N_32092);
nor U46818 (N_46818,N_39901,N_35861);
and U46819 (N_46819,N_38590,N_35375);
or U46820 (N_46820,N_34329,N_34072);
nor U46821 (N_46821,N_30587,N_36859);
nand U46822 (N_46822,N_32743,N_33747);
or U46823 (N_46823,N_33204,N_31121);
nor U46824 (N_46824,N_31824,N_34437);
and U46825 (N_46825,N_30280,N_31185);
nand U46826 (N_46826,N_37337,N_31423);
nor U46827 (N_46827,N_39391,N_31072);
and U46828 (N_46828,N_35370,N_37627);
nand U46829 (N_46829,N_39957,N_31450);
nor U46830 (N_46830,N_38302,N_37587);
nor U46831 (N_46831,N_30772,N_34467);
and U46832 (N_46832,N_33033,N_39160);
nand U46833 (N_46833,N_31334,N_33059);
nor U46834 (N_46834,N_39421,N_35877);
xor U46835 (N_46835,N_35439,N_35109);
or U46836 (N_46836,N_34825,N_34492);
or U46837 (N_46837,N_34524,N_36844);
or U46838 (N_46838,N_38143,N_39670);
nor U46839 (N_46839,N_38186,N_39216);
nor U46840 (N_46840,N_39485,N_31082);
nand U46841 (N_46841,N_38040,N_36072);
nor U46842 (N_46842,N_38008,N_34064);
nor U46843 (N_46843,N_36029,N_31840);
nor U46844 (N_46844,N_30450,N_30420);
nor U46845 (N_46845,N_32903,N_31028);
nand U46846 (N_46846,N_38264,N_32579);
and U46847 (N_46847,N_32734,N_33684);
or U46848 (N_46848,N_35803,N_37796);
or U46849 (N_46849,N_39947,N_33487);
nor U46850 (N_46850,N_37869,N_36982);
xor U46851 (N_46851,N_30822,N_34590);
nor U46852 (N_46852,N_38099,N_37348);
or U46853 (N_46853,N_36599,N_32941);
nand U46854 (N_46854,N_36955,N_36130);
nand U46855 (N_46855,N_38585,N_34431);
or U46856 (N_46856,N_35093,N_36585);
nor U46857 (N_46857,N_32551,N_34872);
nand U46858 (N_46858,N_31715,N_37498);
or U46859 (N_46859,N_33496,N_37577);
nand U46860 (N_46860,N_30119,N_37064);
or U46861 (N_46861,N_39569,N_38356);
and U46862 (N_46862,N_39013,N_31335);
nand U46863 (N_46863,N_33142,N_37557);
nand U46864 (N_46864,N_35273,N_37186);
xor U46865 (N_46865,N_36522,N_36064);
or U46866 (N_46866,N_31394,N_38750);
and U46867 (N_46867,N_34103,N_38700);
nor U46868 (N_46868,N_39732,N_38563);
nor U46869 (N_46869,N_37033,N_35068);
nand U46870 (N_46870,N_32817,N_38808);
nor U46871 (N_46871,N_32260,N_33510);
and U46872 (N_46872,N_31724,N_32514);
nor U46873 (N_46873,N_31029,N_33732);
xor U46874 (N_46874,N_35336,N_38928);
nor U46875 (N_46875,N_39078,N_39846);
nor U46876 (N_46876,N_31755,N_33235);
nor U46877 (N_46877,N_30835,N_32731);
nand U46878 (N_46878,N_38670,N_37040);
nand U46879 (N_46879,N_30702,N_30286);
nor U46880 (N_46880,N_34879,N_37091);
nand U46881 (N_46881,N_34041,N_32148);
xnor U46882 (N_46882,N_33981,N_32256);
nor U46883 (N_46883,N_33947,N_38552);
or U46884 (N_46884,N_33407,N_33444);
nor U46885 (N_46885,N_34110,N_39567);
nand U46886 (N_46886,N_32901,N_30813);
nor U46887 (N_46887,N_39908,N_32062);
or U46888 (N_46888,N_35737,N_33258);
and U46889 (N_46889,N_31870,N_36777);
and U46890 (N_46890,N_38510,N_36582);
or U46891 (N_46891,N_39627,N_36759);
nand U46892 (N_46892,N_39872,N_32029);
nor U46893 (N_46893,N_37440,N_39153);
xor U46894 (N_46894,N_35882,N_39371);
nor U46895 (N_46895,N_38768,N_39064);
xnor U46896 (N_46896,N_31565,N_38800);
nand U46897 (N_46897,N_39247,N_34329);
nor U46898 (N_46898,N_31596,N_39051);
xor U46899 (N_46899,N_39659,N_34657);
or U46900 (N_46900,N_39010,N_31843);
nor U46901 (N_46901,N_38113,N_37224);
or U46902 (N_46902,N_35155,N_39207);
nor U46903 (N_46903,N_36037,N_30174);
or U46904 (N_46904,N_31227,N_36950);
nand U46905 (N_46905,N_31248,N_33921);
nand U46906 (N_46906,N_39006,N_38236);
nor U46907 (N_46907,N_30773,N_39488);
or U46908 (N_46908,N_38965,N_37517);
or U46909 (N_46909,N_38908,N_32497);
nand U46910 (N_46910,N_35329,N_33942);
and U46911 (N_46911,N_36621,N_30516);
nor U46912 (N_46912,N_34194,N_35220);
and U46913 (N_46913,N_35847,N_36342);
nand U46914 (N_46914,N_38588,N_31329);
nor U46915 (N_46915,N_36808,N_34922);
and U46916 (N_46916,N_36741,N_33297);
or U46917 (N_46917,N_31353,N_35464);
nor U46918 (N_46918,N_39839,N_31075);
xnor U46919 (N_46919,N_39491,N_35936);
nor U46920 (N_46920,N_39224,N_32144);
or U46921 (N_46921,N_33384,N_36866);
nand U46922 (N_46922,N_37998,N_33788);
xnor U46923 (N_46923,N_30949,N_39820);
and U46924 (N_46924,N_38214,N_35053);
and U46925 (N_46925,N_35329,N_38381);
or U46926 (N_46926,N_30631,N_30079);
nor U46927 (N_46927,N_34934,N_36346);
or U46928 (N_46928,N_30298,N_34180);
xor U46929 (N_46929,N_39732,N_38443);
nor U46930 (N_46930,N_34490,N_30259);
xnor U46931 (N_46931,N_33729,N_32927);
nand U46932 (N_46932,N_37956,N_31868);
nor U46933 (N_46933,N_35885,N_32996);
nand U46934 (N_46934,N_33646,N_32362);
nor U46935 (N_46935,N_39431,N_33543);
xnor U46936 (N_46936,N_38403,N_33253);
nand U46937 (N_46937,N_34228,N_31803);
nand U46938 (N_46938,N_30183,N_31032);
nor U46939 (N_46939,N_38327,N_33180);
or U46940 (N_46940,N_31737,N_39217);
nor U46941 (N_46941,N_36455,N_37156);
nor U46942 (N_46942,N_31225,N_35124);
or U46943 (N_46943,N_39849,N_31480);
nor U46944 (N_46944,N_33028,N_39386);
nor U46945 (N_46945,N_37709,N_33334);
and U46946 (N_46946,N_38238,N_30363);
and U46947 (N_46947,N_30732,N_37587);
nand U46948 (N_46948,N_32383,N_32607);
xnor U46949 (N_46949,N_34905,N_34784);
nand U46950 (N_46950,N_34114,N_36320);
and U46951 (N_46951,N_37382,N_39732);
nand U46952 (N_46952,N_37070,N_37509);
or U46953 (N_46953,N_32221,N_38575);
nand U46954 (N_46954,N_35010,N_36376);
nor U46955 (N_46955,N_36557,N_36465);
or U46956 (N_46956,N_39010,N_38338);
nor U46957 (N_46957,N_30246,N_36525);
or U46958 (N_46958,N_36282,N_32906);
nor U46959 (N_46959,N_32001,N_34505);
or U46960 (N_46960,N_38963,N_30468);
nand U46961 (N_46961,N_32966,N_30810);
or U46962 (N_46962,N_31422,N_30479);
and U46963 (N_46963,N_34502,N_30137);
nand U46964 (N_46964,N_34831,N_34004);
xor U46965 (N_46965,N_38903,N_30766);
and U46966 (N_46966,N_37606,N_37738);
and U46967 (N_46967,N_31212,N_32462);
and U46968 (N_46968,N_35766,N_30312);
and U46969 (N_46969,N_31512,N_32416);
nor U46970 (N_46970,N_32234,N_33206);
and U46971 (N_46971,N_32093,N_37324);
or U46972 (N_46972,N_32996,N_36255);
nor U46973 (N_46973,N_37777,N_33238);
and U46974 (N_46974,N_37430,N_35863);
nor U46975 (N_46975,N_37693,N_31354);
nor U46976 (N_46976,N_32504,N_31986);
and U46977 (N_46977,N_30585,N_33297);
nor U46978 (N_46978,N_37951,N_33137);
or U46979 (N_46979,N_32768,N_37172);
xnor U46980 (N_46980,N_33672,N_32184);
xnor U46981 (N_46981,N_37885,N_38857);
nand U46982 (N_46982,N_37521,N_31782);
and U46983 (N_46983,N_38233,N_37835);
nand U46984 (N_46984,N_31405,N_33841);
or U46985 (N_46985,N_36448,N_33817);
and U46986 (N_46986,N_35719,N_39874);
nor U46987 (N_46987,N_38687,N_32254);
and U46988 (N_46988,N_38005,N_30159);
and U46989 (N_46989,N_37304,N_34975);
xnor U46990 (N_46990,N_30562,N_32160);
and U46991 (N_46991,N_30198,N_31271);
and U46992 (N_46992,N_39970,N_31092);
nor U46993 (N_46993,N_36295,N_38916);
or U46994 (N_46994,N_34167,N_33829);
and U46995 (N_46995,N_34067,N_39642);
nor U46996 (N_46996,N_32836,N_36013);
nand U46997 (N_46997,N_39758,N_39913);
nor U46998 (N_46998,N_35879,N_37114);
and U46999 (N_46999,N_33419,N_36952);
and U47000 (N_47000,N_32026,N_30072);
nor U47001 (N_47001,N_36746,N_35454);
nand U47002 (N_47002,N_31055,N_37080);
or U47003 (N_47003,N_30460,N_39618);
xnor U47004 (N_47004,N_37622,N_34019);
xnor U47005 (N_47005,N_38935,N_35513);
and U47006 (N_47006,N_32565,N_34147);
nor U47007 (N_47007,N_38028,N_38703);
xnor U47008 (N_47008,N_37856,N_36094);
and U47009 (N_47009,N_30350,N_37435);
and U47010 (N_47010,N_39810,N_30879);
nand U47011 (N_47011,N_39933,N_38058);
or U47012 (N_47012,N_34392,N_31626);
and U47013 (N_47013,N_36971,N_36385);
nor U47014 (N_47014,N_37466,N_35620);
nor U47015 (N_47015,N_39571,N_30685);
nor U47016 (N_47016,N_30164,N_38161);
and U47017 (N_47017,N_38715,N_32317);
and U47018 (N_47018,N_34723,N_31712);
nand U47019 (N_47019,N_39280,N_30481);
nand U47020 (N_47020,N_32904,N_31409);
or U47021 (N_47021,N_38917,N_31851);
and U47022 (N_47022,N_33266,N_34584);
nand U47023 (N_47023,N_35333,N_30792);
and U47024 (N_47024,N_39797,N_35793);
or U47025 (N_47025,N_37095,N_34365);
and U47026 (N_47026,N_37032,N_39512);
nand U47027 (N_47027,N_38218,N_30928);
and U47028 (N_47028,N_32870,N_34680);
nand U47029 (N_47029,N_32882,N_35073);
and U47030 (N_47030,N_32528,N_30671);
and U47031 (N_47031,N_39794,N_30344);
and U47032 (N_47032,N_36326,N_35822);
or U47033 (N_47033,N_39736,N_34947);
nand U47034 (N_47034,N_37956,N_37836);
and U47035 (N_47035,N_39283,N_32280);
nand U47036 (N_47036,N_38333,N_36769);
and U47037 (N_47037,N_33761,N_31612);
or U47038 (N_47038,N_34609,N_39786);
nand U47039 (N_47039,N_36791,N_30027);
nor U47040 (N_47040,N_31161,N_31819);
xor U47041 (N_47041,N_31829,N_30656);
nand U47042 (N_47042,N_31723,N_36390);
nor U47043 (N_47043,N_36171,N_38499);
xnor U47044 (N_47044,N_38143,N_33324);
nor U47045 (N_47045,N_38365,N_33098);
nand U47046 (N_47046,N_30227,N_34544);
or U47047 (N_47047,N_36825,N_35402);
nand U47048 (N_47048,N_37118,N_30785);
or U47049 (N_47049,N_35825,N_31277);
nor U47050 (N_47050,N_33451,N_37258);
nand U47051 (N_47051,N_31023,N_36927);
and U47052 (N_47052,N_34358,N_39275);
and U47053 (N_47053,N_36556,N_36677);
or U47054 (N_47054,N_32738,N_34874);
and U47055 (N_47055,N_33424,N_37612);
nor U47056 (N_47056,N_30757,N_39290);
nand U47057 (N_47057,N_38166,N_37970);
xor U47058 (N_47058,N_34247,N_31967);
and U47059 (N_47059,N_33417,N_38544);
and U47060 (N_47060,N_39106,N_35192);
nand U47061 (N_47061,N_30848,N_33144);
and U47062 (N_47062,N_30068,N_31604);
and U47063 (N_47063,N_39930,N_38983);
nor U47064 (N_47064,N_37188,N_32865);
and U47065 (N_47065,N_33013,N_38068);
and U47066 (N_47066,N_35007,N_30590);
or U47067 (N_47067,N_36660,N_34789);
and U47068 (N_47068,N_36151,N_39028);
and U47069 (N_47069,N_34081,N_38758);
nand U47070 (N_47070,N_33436,N_35654);
nand U47071 (N_47071,N_33394,N_33595);
nand U47072 (N_47072,N_33266,N_31614);
xor U47073 (N_47073,N_33717,N_31223);
or U47074 (N_47074,N_32518,N_31895);
or U47075 (N_47075,N_39989,N_30728);
nand U47076 (N_47076,N_32442,N_37622);
nor U47077 (N_47077,N_39885,N_37085);
nand U47078 (N_47078,N_36152,N_32054);
nand U47079 (N_47079,N_32151,N_32602);
and U47080 (N_47080,N_37230,N_36449);
or U47081 (N_47081,N_34380,N_34447);
and U47082 (N_47082,N_33328,N_31278);
nor U47083 (N_47083,N_36454,N_30309);
or U47084 (N_47084,N_32295,N_30875);
and U47085 (N_47085,N_39385,N_38889);
or U47086 (N_47086,N_38075,N_31326);
and U47087 (N_47087,N_31967,N_39994);
xor U47088 (N_47088,N_39692,N_36727);
xnor U47089 (N_47089,N_36629,N_33133);
and U47090 (N_47090,N_32364,N_34547);
and U47091 (N_47091,N_36336,N_39356);
nand U47092 (N_47092,N_36086,N_30314);
xnor U47093 (N_47093,N_37580,N_39112);
or U47094 (N_47094,N_35165,N_30075);
or U47095 (N_47095,N_31306,N_32507);
nand U47096 (N_47096,N_39022,N_36758);
nand U47097 (N_47097,N_35608,N_33529);
nand U47098 (N_47098,N_34155,N_39005);
and U47099 (N_47099,N_38631,N_39891);
or U47100 (N_47100,N_33051,N_37653);
and U47101 (N_47101,N_36103,N_36687);
xor U47102 (N_47102,N_34654,N_33859);
or U47103 (N_47103,N_30719,N_37577);
and U47104 (N_47104,N_31767,N_39802);
nor U47105 (N_47105,N_35934,N_31238);
and U47106 (N_47106,N_35999,N_39312);
and U47107 (N_47107,N_34273,N_36064);
xnor U47108 (N_47108,N_34147,N_38883);
nor U47109 (N_47109,N_38611,N_32003);
nand U47110 (N_47110,N_39817,N_33740);
nor U47111 (N_47111,N_33349,N_30863);
or U47112 (N_47112,N_38743,N_34508);
xnor U47113 (N_47113,N_31426,N_35698);
and U47114 (N_47114,N_39431,N_38976);
or U47115 (N_47115,N_33660,N_33268);
nand U47116 (N_47116,N_37537,N_39123);
and U47117 (N_47117,N_30449,N_30994);
nand U47118 (N_47118,N_33250,N_39069);
or U47119 (N_47119,N_36158,N_39039);
or U47120 (N_47120,N_35248,N_34971);
and U47121 (N_47121,N_35605,N_37190);
or U47122 (N_47122,N_38904,N_37840);
or U47123 (N_47123,N_38606,N_33371);
nand U47124 (N_47124,N_39181,N_37412);
nand U47125 (N_47125,N_33020,N_32443);
nand U47126 (N_47126,N_34137,N_32498);
and U47127 (N_47127,N_38763,N_34049);
and U47128 (N_47128,N_32212,N_33549);
nand U47129 (N_47129,N_30440,N_31266);
and U47130 (N_47130,N_31360,N_30953);
or U47131 (N_47131,N_34664,N_34989);
nor U47132 (N_47132,N_34638,N_31535);
nor U47133 (N_47133,N_30915,N_32845);
nand U47134 (N_47134,N_38788,N_36436);
and U47135 (N_47135,N_38522,N_34668);
nand U47136 (N_47136,N_31782,N_36278);
nor U47137 (N_47137,N_33602,N_36928);
and U47138 (N_47138,N_37764,N_34190);
nor U47139 (N_47139,N_37290,N_37773);
and U47140 (N_47140,N_35960,N_39672);
or U47141 (N_47141,N_34850,N_31673);
nor U47142 (N_47142,N_38751,N_39535);
nor U47143 (N_47143,N_36179,N_35160);
xnor U47144 (N_47144,N_37114,N_33003);
or U47145 (N_47145,N_31739,N_36515);
nor U47146 (N_47146,N_37859,N_32858);
xor U47147 (N_47147,N_38634,N_31762);
nand U47148 (N_47148,N_30827,N_38325);
nor U47149 (N_47149,N_35248,N_38468);
nor U47150 (N_47150,N_35950,N_36238);
xnor U47151 (N_47151,N_30211,N_31971);
and U47152 (N_47152,N_36990,N_31819);
or U47153 (N_47153,N_36182,N_30655);
or U47154 (N_47154,N_33487,N_39094);
nor U47155 (N_47155,N_39224,N_36895);
nor U47156 (N_47156,N_33983,N_32798);
nor U47157 (N_47157,N_33434,N_30741);
nand U47158 (N_47158,N_30121,N_39492);
nor U47159 (N_47159,N_33715,N_35033);
nand U47160 (N_47160,N_33294,N_31268);
and U47161 (N_47161,N_36060,N_39642);
or U47162 (N_47162,N_37323,N_33041);
xor U47163 (N_47163,N_32961,N_35201);
xor U47164 (N_47164,N_39001,N_39519);
nor U47165 (N_47165,N_37209,N_37523);
xnor U47166 (N_47166,N_35979,N_34299);
and U47167 (N_47167,N_30273,N_33692);
xor U47168 (N_47168,N_31559,N_33114);
nor U47169 (N_47169,N_37487,N_37282);
nand U47170 (N_47170,N_33241,N_31181);
or U47171 (N_47171,N_31542,N_34256);
and U47172 (N_47172,N_39267,N_30442);
and U47173 (N_47173,N_34157,N_30766);
nor U47174 (N_47174,N_39083,N_32409);
or U47175 (N_47175,N_33487,N_30268);
or U47176 (N_47176,N_38890,N_30459);
or U47177 (N_47177,N_32994,N_33461);
or U47178 (N_47178,N_35327,N_35034);
xnor U47179 (N_47179,N_33393,N_33836);
nor U47180 (N_47180,N_32116,N_33765);
nand U47181 (N_47181,N_32302,N_35649);
xnor U47182 (N_47182,N_30572,N_33779);
and U47183 (N_47183,N_36302,N_36279);
or U47184 (N_47184,N_30800,N_33642);
or U47185 (N_47185,N_36763,N_34294);
nor U47186 (N_47186,N_38943,N_35965);
nand U47187 (N_47187,N_36650,N_36083);
or U47188 (N_47188,N_30138,N_36781);
or U47189 (N_47189,N_38405,N_37146);
and U47190 (N_47190,N_38973,N_34544);
nor U47191 (N_47191,N_30191,N_32270);
xor U47192 (N_47192,N_35781,N_38017);
and U47193 (N_47193,N_37049,N_35041);
or U47194 (N_47194,N_34450,N_34583);
nor U47195 (N_47195,N_33658,N_35627);
nand U47196 (N_47196,N_31286,N_39434);
and U47197 (N_47197,N_39116,N_32797);
and U47198 (N_47198,N_39350,N_33068);
and U47199 (N_47199,N_39832,N_38562);
nor U47200 (N_47200,N_34235,N_34370);
nand U47201 (N_47201,N_39733,N_31206);
and U47202 (N_47202,N_34282,N_38827);
xnor U47203 (N_47203,N_30676,N_33771);
and U47204 (N_47204,N_38754,N_33066);
nand U47205 (N_47205,N_35365,N_38800);
nand U47206 (N_47206,N_38326,N_32973);
nand U47207 (N_47207,N_37309,N_30946);
nand U47208 (N_47208,N_37025,N_37297);
nor U47209 (N_47209,N_32045,N_30632);
or U47210 (N_47210,N_38268,N_39356);
xor U47211 (N_47211,N_36597,N_33265);
or U47212 (N_47212,N_37714,N_39310);
and U47213 (N_47213,N_37781,N_31558);
and U47214 (N_47214,N_31178,N_38025);
and U47215 (N_47215,N_39891,N_39221);
nor U47216 (N_47216,N_33173,N_35158);
xor U47217 (N_47217,N_34154,N_35348);
and U47218 (N_47218,N_32782,N_33283);
xnor U47219 (N_47219,N_31245,N_31473);
and U47220 (N_47220,N_35485,N_30929);
nor U47221 (N_47221,N_31573,N_36706);
nor U47222 (N_47222,N_31531,N_33855);
nand U47223 (N_47223,N_35679,N_39511);
nand U47224 (N_47224,N_34170,N_31015);
and U47225 (N_47225,N_36575,N_38166);
nand U47226 (N_47226,N_38439,N_34441);
or U47227 (N_47227,N_36877,N_35641);
nand U47228 (N_47228,N_34267,N_30524);
or U47229 (N_47229,N_34020,N_38340);
xor U47230 (N_47230,N_34050,N_34658);
nand U47231 (N_47231,N_30965,N_31235);
nor U47232 (N_47232,N_31199,N_38304);
nand U47233 (N_47233,N_38933,N_35607);
nor U47234 (N_47234,N_35762,N_33815);
and U47235 (N_47235,N_39457,N_34592);
xnor U47236 (N_47236,N_33365,N_32531);
nand U47237 (N_47237,N_31037,N_34403);
or U47238 (N_47238,N_39894,N_39393);
nor U47239 (N_47239,N_37793,N_34849);
and U47240 (N_47240,N_34205,N_30945);
or U47241 (N_47241,N_30580,N_35777);
or U47242 (N_47242,N_37061,N_34332);
nor U47243 (N_47243,N_37332,N_33132);
xor U47244 (N_47244,N_34237,N_33247);
or U47245 (N_47245,N_35551,N_32762);
or U47246 (N_47246,N_35480,N_39817);
nand U47247 (N_47247,N_36471,N_36375);
nand U47248 (N_47248,N_37426,N_38553);
nor U47249 (N_47249,N_30707,N_32831);
nand U47250 (N_47250,N_32945,N_38025);
nand U47251 (N_47251,N_34119,N_36094);
or U47252 (N_47252,N_31319,N_31374);
nor U47253 (N_47253,N_33822,N_34860);
or U47254 (N_47254,N_31522,N_35181);
nand U47255 (N_47255,N_37353,N_32465);
nand U47256 (N_47256,N_31677,N_38825);
xnor U47257 (N_47257,N_30793,N_38036);
and U47258 (N_47258,N_35258,N_35198);
and U47259 (N_47259,N_30046,N_36162);
xor U47260 (N_47260,N_33431,N_37216);
nand U47261 (N_47261,N_30639,N_32647);
nor U47262 (N_47262,N_36258,N_36581);
xnor U47263 (N_47263,N_31087,N_34157);
nor U47264 (N_47264,N_36928,N_38436);
nand U47265 (N_47265,N_31172,N_30544);
and U47266 (N_47266,N_39050,N_36204);
and U47267 (N_47267,N_34352,N_32544);
nor U47268 (N_47268,N_32854,N_30102);
nand U47269 (N_47269,N_37127,N_32062);
nor U47270 (N_47270,N_36102,N_31923);
and U47271 (N_47271,N_34635,N_37099);
or U47272 (N_47272,N_35673,N_37033);
nor U47273 (N_47273,N_35596,N_31910);
nor U47274 (N_47274,N_38468,N_35511);
and U47275 (N_47275,N_32217,N_39742);
nand U47276 (N_47276,N_33265,N_34017);
or U47277 (N_47277,N_30080,N_34638);
nand U47278 (N_47278,N_32912,N_38857);
or U47279 (N_47279,N_34350,N_39625);
nor U47280 (N_47280,N_37819,N_33843);
nand U47281 (N_47281,N_34265,N_33594);
or U47282 (N_47282,N_30280,N_32027);
nor U47283 (N_47283,N_38465,N_36640);
or U47284 (N_47284,N_30688,N_33309);
xor U47285 (N_47285,N_31335,N_34609);
and U47286 (N_47286,N_34433,N_30298);
xnor U47287 (N_47287,N_32979,N_36652);
and U47288 (N_47288,N_37956,N_38657);
or U47289 (N_47289,N_33221,N_32208);
nor U47290 (N_47290,N_38584,N_39520);
or U47291 (N_47291,N_35198,N_36957);
nand U47292 (N_47292,N_37123,N_33391);
and U47293 (N_47293,N_39975,N_39110);
nor U47294 (N_47294,N_31841,N_37594);
or U47295 (N_47295,N_30055,N_37730);
and U47296 (N_47296,N_38976,N_33680);
or U47297 (N_47297,N_31094,N_37217);
xnor U47298 (N_47298,N_33837,N_34089);
nor U47299 (N_47299,N_36109,N_36787);
or U47300 (N_47300,N_39237,N_36019);
or U47301 (N_47301,N_33437,N_33310);
or U47302 (N_47302,N_38585,N_36606);
xnor U47303 (N_47303,N_36609,N_37490);
xor U47304 (N_47304,N_37285,N_38323);
or U47305 (N_47305,N_32528,N_37757);
and U47306 (N_47306,N_34336,N_32607);
or U47307 (N_47307,N_34852,N_33145);
and U47308 (N_47308,N_35639,N_35113);
or U47309 (N_47309,N_36814,N_36878);
nor U47310 (N_47310,N_33122,N_31171);
or U47311 (N_47311,N_38146,N_39583);
and U47312 (N_47312,N_39693,N_30804);
nand U47313 (N_47313,N_31613,N_33088);
nor U47314 (N_47314,N_33310,N_36857);
or U47315 (N_47315,N_36429,N_35987);
xnor U47316 (N_47316,N_33656,N_39766);
and U47317 (N_47317,N_35841,N_35756);
nor U47318 (N_47318,N_35436,N_38603);
nand U47319 (N_47319,N_34029,N_35835);
nor U47320 (N_47320,N_33399,N_32016);
xor U47321 (N_47321,N_36381,N_31243);
nand U47322 (N_47322,N_35074,N_37800);
nand U47323 (N_47323,N_33346,N_36932);
or U47324 (N_47324,N_30234,N_33936);
nand U47325 (N_47325,N_33587,N_39247);
or U47326 (N_47326,N_39679,N_39125);
nand U47327 (N_47327,N_36069,N_33256);
or U47328 (N_47328,N_37785,N_36407);
or U47329 (N_47329,N_38683,N_34634);
nor U47330 (N_47330,N_34682,N_37620);
xnor U47331 (N_47331,N_36675,N_34990);
and U47332 (N_47332,N_38314,N_38819);
nor U47333 (N_47333,N_38795,N_32989);
and U47334 (N_47334,N_35673,N_38400);
and U47335 (N_47335,N_32776,N_35093);
nand U47336 (N_47336,N_30097,N_35829);
and U47337 (N_47337,N_30636,N_38592);
nand U47338 (N_47338,N_37968,N_36994);
nor U47339 (N_47339,N_30270,N_37665);
or U47340 (N_47340,N_36131,N_36893);
nand U47341 (N_47341,N_36765,N_37139);
nand U47342 (N_47342,N_39970,N_35633);
and U47343 (N_47343,N_30390,N_34611);
nor U47344 (N_47344,N_38864,N_35883);
and U47345 (N_47345,N_30839,N_31255);
nor U47346 (N_47346,N_32165,N_39159);
or U47347 (N_47347,N_37682,N_35449);
nand U47348 (N_47348,N_32812,N_34149);
xnor U47349 (N_47349,N_33123,N_36449);
xor U47350 (N_47350,N_38324,N_35409);
or U47351 (N_47351,N_32732,N_37994);
and U47352 (N_47352,N_30928,N_35759);
nor U47353 (N_47353,N_36449,N_36726);
or U47354 (N_47354,N_32625,N_34606);
xnor U47355 (N_47355,N_37164,N_31471);
nand U47356 (N_47356,N_37291,N_33577);
nor U47357 (N_47357,N_34873,N_31146);
or U47358 (N_47358,N_31720,N_36813);
nand U47359 (N_47359,N_31537,N_31761);
nor U47360 (N_47360,N_34424,N_35210);
nand U47361 (N_47361,N_35049,N_36620);
or U47362 (N_47362,N_33682,N_38768);
nor U47363 (N_47363,N_37533,N_32878);
and U47364 (N_47364,N_32929,N_38038);
or U47365 (N_47365,N_31534,N_35831);
xnor U47366 (N_47366,N_36434,N_36011);
nand U47367 (N_47367,N_39430,N_37237);
nor U47368 (N_47368,N_39490,N_36637);
or U47369 (N_47369,N_38528,N_38594);
or U47370 (N_47370,N_39741,N_30643);
or U47371 (N_47371,N_38432,N_31264);
and U47372 (N_47372,N_30730,N_31895);
xor U47373 (N_47373,N_36577,N_33178);
and U47374 (N_47374,N_35732,N_34635);
nand U47375 (N_47375,N_36739,N_30137);
or U47376 (N_47376,N_34438,N_30308);
xnor U47377 (N_47377,N_30706,N_38698);
and U47378 (N_47378,N_31279,N_36166);
nand U47379 (N_47379,N_37435,N_38659);
or U47380 (N_47380,N_33930,N_32225);
nand U47381 (N_47381,N_32093,N_32589);
or U47382 (N_47382,N_30493,N_39698);
nor U47383 (N_47383,N_32326,N_37985);
and U47384 (N_47384,N_32521,N_38916);
nand U47385 (N_47385,N_34634,N_39339);
nor U47386 (N_47386,N_38363,N_35700);
xnor U47387 (N_47387,N_32269,N_38450);
and U47388 (N_47388,N_37253,N_32008);
or U47389 (N_47389,N_36225,N_30972);
nor U47390 (N_47390,N_36235,N_34805);
and U47391 (N_47391,N_32961,N_32095);
nor U47392 (N_47392,N_39926,N_31079);
and U47393 (N_47393,N_32537,N_39553);
nor U47394 (N_47394,N_36733,N_34031);
or U47395 (N_47395,N_30978,N_39452);
nand U47396 (N_47396,N_31810,N_31792);
or U47397 (N_47397,N_34279,N_33905);
nor U47398 (N_47398,N_33529,N_32316);
nand U47399 (N_47399,N_34999,N_36860);
or U47400 (N_47400,N_32016,N_37195);
and U47401 (N_47401,N_32458,N_34573);
nor U47402 (N_47402,N_33680,N_39804);
nor U47403 (N_47403,N_31398,N_38010);
and U47404 (N_47404,N_39327,N_31597);
nand U47405 (N_47405,N_38733,N_39255);
or U47406 (N_47406,N_36463,N_30799);
nand U47407 (N_47407,N_33500,N_34745);
or U47408 (N_47408,N_33256,N_34140);
nand U47409 (N_47409,N_35200,N_38718);
or U47410 (N_47410,N_36734,N_38643);
nand U47411 (N_47411,N_34778,N_30180);
nor U47412 (N_47412,N_32819,N_36482);
nor U47413 (N_47413,N_38156,N_36784);
nor U47414 (N_47414,N_34106,N_32639);
and U47415 (N_47415,N_36904,N_34900);
xor U47416 (N_47416,N_32683,N_39679);
or U47417 (N_47417,N_35044,N_39191);
or U47418 (N_47418,N_35826,N_36770);
nand U47419 (N_47419,N_31787,N_37095);
and U47420 (N_47420,N_32783,N_36494);
nand U47421 (N_47421,N_31567,N_33572);
or U47422 (N_47422,N_30055,N_34158);
nand U47423 (N_47423,N_39264,N_35490);
and U47424 (N_47424,N_33586,N_32581);
and U47425 (N_47425,N_38861,N_32206);
or U47426 (N_47426,N_31553,N_33571);
and U47427 (N_47427,N_35327,N_33499);
and U47428 (N_47428,N_31717,N_31002);
or U47429 (N_47429,N_39504,N_38495);
or U47430 (N_47430,N_31645,N_39497);
or U47431 (N_47431,N_34748,N_39604);
nor U47432 (N_47432,N_31264,N_36369);
or U47433 (N_47433,N_30047,N_38042);
or U47434 (N_47434,N_39944,N_36856);
nor U47435 (N_47435,N_32839,N_34941);
nand U47436 (N_47436,N_38810,N_38180);
and U47437 (N_47437,N_30050,N_36050);
and U47438 (N_47438,N_31767,N_30611);
nor U47439 (N_47439,N_32753,N_35229);
and U47440 (N_47440,N_31615,N_35309);
nor U47441 (N_47441,N_38030,N_34708);
nand U47442 (N_47442,N_38446,N_35308);
or U47443 (N_47443,N_33467,N_31795);
or U47444 (N_47444,N_32174,N_31497);
nand U47445 (N_47445,N_38139,N_32500);
nor U47446 (N_47446,N_36681,N_35694);
or U47447 (N_47447,N_33766,N_30274);
or U47448 (N_47448,N_30757,N_37462);
xnor U47449 (N_47449,N_34288,N_36301);
or U47450 (N_47450,N_31000,N_36198);
nand U47451 (N_47451,N_31368,N_34420);
nand U47452 (N_47452,N_32058,N_31792);
nand U47453 (N_47453,N_33485,N_30800);
and U47454 (N_47454,N_34025,N_36029);
and U47455 (N_47455,N_38103,N_35817);
nor U47456 (N_47456,N_39082,N_36071);
nand U47457 (N_47457,N_34073,N_30354);
nand U47458 (N_47458,N_34137,N_38847);
and U47459 (N_47459,N_37649,N_32527);
nor U47460 (N_47460,N_35151,N_39018);
and U47461 (N_47461,N_30358,N_35888);
nand U47462 (N_47462,N_38670,N_31057);
nor U47463 (N_47463,N_33011,N_36243);
nor U47464 (N_47464,N_37561,N_37863);
nor U47465 (N_47465,N_34723,N_37037);
nor U47466 (N_47466,N_36510,N_39973);
or U47467 (N_47467,N_36110,N_30191);
nor U47468 (N_47468,N_35009,N_33957);
xnor U47469 (N_47469,N_36838,N_38378);
or U47470 (N_47470,N_34441,N_35959);
nor U47471 (N_47471,N_38026,N_38511);
or U47472 (N_47472,N_34741,N_34689);
nor U47473 (N_47473,N_32514,N_36593);
nor U47474 (N_47474,N_31620,N_38927);
or U47475 (N_47475,N_39700,N_34916);
or U47476 (N_47476,N_33674,N_30132);
and U47477 (N_47477,N_37977,N_37802);
nor U47478 (N_47478,N_31499,N_34601);
xor U47479 (N_47479,N_37272,N_37874);
or U47480 (N_47480,N_36506,N_34893);
xor U47481 (N_47481,N_31014,N_37766);
nand U47482 (N_47482,N_37202,N_32088);
or U47483 (N_47483,N_32898,N_36019);
and U47484 (N_47484,N_33019,N_37611);
and U47485 (N_47485,N_39745,N_30147);
nor U47486 (N_47486,N_31163,N_38832);
or U47487 (N_47487,N_35779,N_34684);
nor U47488 (N_47488,N_38213,N_33103);
or U47489 (N_47489,N_36496,N_32338);
xor U47490 (N_47490,N_33650,N_32841);
nor U47491 (N_47491,N_39582,N_33214);
xnor U47492 (N_47492,N_36192,N_37059);
or U47493 (N_47493,N_34013,N_33727);
and U47494 (N_47494,N_30964,N_32808);
nor U47495 (N_47495,N_38968,N_39588);
or U47496 (N_47496,N_32782,N_36132);
and U47497 (N_47497,N_30651,N_36050);
xor U47498 (N_47498,N_39188,N_30333);
nor U47499 (N_47499,N_39276,N_39535);
nor U47500 (N_47500,N_36537,N_37182);
or U47501 (N_47501,N_38885,N_38309);
xnor U47502 (N_47502,N_32187,N_35055);
or U47503 (N_47503,N_36548,N_33131);
xor U47504 (N_47504,N_37965,N_38247);
and U47505 (N_47505,N_30649,N_31852);
nor U47506 (N_47506,N_32411,N_39101);
xnor U47507 (N_47507,N_32858,N_30698);
or U47508 (N_47508,N_34818,N_32309);
nand U47509 (N_47509,N_30261,N_34519);
nor U47510 (N_47510,N_39526,N_34918);
and U47511 (N_47511,N_34051,N_39031);
and U47512 (N_47512,N_33208,N_33841);
nand U47513 (N_47513,N_37256,N_30626);
and U47514 (N_47514,N_31104,N_38628);
and U47515 (N_47515,N_34474,N_38959);
or U47516 (N_47516,N_30128,N_32445);
nand U47517 (N_47517,N_32086,N_34676);
nand U47518 (N_47518,N_39366,N_30668);
xnor U47519 (N_47519,N_31798,N_33145);
nand U47520 (N_47520,N_30970,N_36577);
xnor U47521 (N_47521,N_39492,N_31322);
or U47522 (N_47522,N_35848,N_31114);
or U47523 (N_47523,N_31561,N_39559);
nor U47524 (N_47524,N_33271,N_37062);
or U47525 (N_47525,N_32279,N_34451);
or U47526 (N_47526,N_31172,N_36645);
and U47527 (N_47527,N_31839,N_38639);
nor U47528 (N_47528,N_37975,N_31526);
nor U47529 (N_47529,N_39941,N_38762);
nor U47530 (N_47530,N_32401,N_32041);
or U47531 (N_47531,N_36318,N_39769);
nand U47532 (N_47532,N_37948,N_39899);
nor U47533 (N_47533,N_32601,N_34929);
or U47534 (N_47534,N_39050,N_35096);
and U47535 (N_47535,N_35417,N_33784);
nor U47536 (N_47536,N_33771,N_33099);
and U47537 (N_47537,N_38574,N_37663);
xnor U47538 (N_47538,N_35211,N_32681);
nor U47539 (N_47539,N_32184,N_38111);
nor U47540 (N_47540,N_33239,N_33466);
nor U47541 (N_47541,N_35486,N_32950);
xnor U47542 (N_47542,N_36457,N_35755);
or U47543 (N_47543,N_34730,N_36566);
nor U47544 (N_47544,N_34706,N_33068);
nand U47545 (N_47545,N_39544,N_33274);
and U47546 (N_47546,N_33742,N_39779);
xor U47547 (N_47547,N_38622,N_39828);
or U47548 (N_47548,N_39738,N_35385);
xor U47549 (N_47549,N_39187,N_31902);
nand U47550 (N_47550,N_34849,N_33843);
or U47551 (N_47551,N_37346,N_36752);
xnor U47552 (N_47552,N_33977,N_38437);
nand U47553 (N_47553,N_39766,N_37698);
and U47554 (N_47554,N_31569,N_31177);
or U47555 (N_47555,N_31331,N_35306);
or U47556 (N_47556,N_34691,N_33817);
and U47557 (N_47557,N_30427,N_35142);
nor U47558 (N_47558,N_39552,N_34340);
nor U47559 (N_47559,N_31232,N_33126);
or U47560 (N_47560,N_31328,N_30546);
xnor U47561 (N_47561,N_34172,N_31131);
or U47562 (N_47562,N_33092,N_37450);
nor U47563 (N_47563,N_33149,N_38968);
and U47564 (N_47564,N_36243,N_32034);
xnor U47565 (N_47565,N_38633,N_37658);
nand U47566 (N_47566,N_36621,N_38891);
xnor U47567 (N_47567,N_36707,N_36459);
or U47568 (N_47568,N_33255,N_39711);
nor U47569 (N_47569,N_30744,N_30538);
nand U47570 (N_47570,N_30775,N_34698);
nand U47571 (N_47571,N_31286,N_37670);
and U47572 (N_47572,N_37826,N_32792);
and U47573 (N_47573,N_33754,N_39733);
or U47574 (N_47574,N_38818,N_31920);
or U47575 (N_47575,N_33390,N_31704);
nor U47576 (N_47576,N_31270,N_38725);
nand U47577 (N_47577,N_33272,N_35999);
nor U47578 (N_47578,N_39883,N_32094);
nor U47579 (N_47579,N_38415,N_35994);
or U47580 (N_47580,N_37086,N_37206);
nor U47581 (N_47581,N_36458,N_34911);
and U47582 (N_47582,N_33412,N_39656);
nand U47583 (N_47583,N_32164,N_30018);
xor U47584 (N_47584,N_30875,N_31232);
or U47585 (N_47585,N_38897,N_33704);
nor U47586 (N_47586,N_31369,N_39503);
or U47587 (N_47587,N_38180,N_34047);
nand U47588 (N_47588,N_39087,N_30530);
nor U47589 (N_47589,N_36278,N_34729);
or U47590 (N_47590,N_31420,N_35687);
nand U47591 (N_47591,N_38341,N_35143);
nor U47592 (N_47592,N_37688,N_34838);
nand U47593 (N_47593,N_33573,N_31191);
nand U47594 (N_47594,N_38776,N_38108);
or U47595 (N_47595,N_31727,N_33929);
nor U47596 (N_47596,N_33477,N_32403);
or U47597 (N_47597,N_32253,N_32086);
and U47598 (N_47598,N_39697,N_35264);
or U47599 (N_47599,N_33436,N_32541);
or U47600 (N_47600,N_32753,N_37097);
and U47601 (N_47601,N_35484,N_37318);
or U47602 (N_47602,N_36756,N_36413);
xor U47603 (N_47603,N_39519,N_39869);
nor U47604 (N_47604,N_36331,N_34309);
nor U47605 (N_47605,N_39063,N_30399);
nor U47606 (N_47606,N_38458,N_34573);
or U47607 (N_47607,N_32413,N_35535);
nor U47608 (N_47608,N_36959,N_37043);
nand U47609 (N_47609,N_39419,N_34926);
nor U47610 (N_47610,N_36834,N_37456);
nor U47611 (N_47611,N_31382,N_31391);
or U47612 (N_47612,N_36680,N_37269);
nor U47613 (N_47613,N_32512,N_35897);
or U47614 (N_47614,N_36608,N_39048);
or U47615 (N_47615,N_36024,N_32755);
nand U47616 (N_47616,N_32002,N_30344);
nand U47617 (N_47617,N_33006,N_34552);
or U47618 (N_47618,N_34381,N_31090);
or U47619 (N_47619,N_30657,N_34410);
or U47620 (N_47620,N_38103,N_37735);
or U47621 (N_47621,N_34525,N_33449);
nor U47622 (N_47622,N_32675,N_32409);
or U47623 (N_47623,N_37056,N_32454);
nand U47624 (N_47624,N_34627,N_32741);
or U47625 (N_47625,N_33425,N_36844);
xor U47626 (N_47626,N_33720,N_34228);
or U47627 (N_47627,N_31324,N_38894);
and U47628 (N_47628,N_30985,N_33460);
or U47629 (N_47629,N_33163,N_36553);
nor U47630 (N_47630,N_39551,N_38803);
nor U47631 (N_47631,N_38314,N_36730);
or U47632 (N_47632,N_36591,N_34605);
nand U47633 (N_47633,N_37421,N_31810);
nor U47634 (N_47634,N_34728,N_33480);
nand U47635 (N_47635,N_39414,N_30139);
nand U47636 (N_47636,N_35196,N_38051);
nor U47637 (N_47637,N_36767,N_31419);
and U47638 (N_47638,N_37538,N_34511);
nand U47639 (N_47639,N_31153,N_33692);
or U47640 (N_47640,N_30875,N_31590);
nor U47641 (N_47641,N_31595,N_39803);
nor U47642 (N_47642,N_31926,N_36641);
nor U47643 (N_47643,N_38844,N_31249);
or U47644 (N_47644,N_37267,N_36564);
nand U47645 (N_47645,N_34763,N_34109);
or U47646 (N_47646,N_37658,N_36578);
nor U47647 (N_47647,N_33790,N_35627);
and U47648 (N_47648,N_31167,N_32819);
or U47649 (N_47649,N_38594,N_34218);
and U47650 (N_47650,N_39098,N_39883);
and U47651 (N_47651,N_30264,N_32937);
nand U47652 (N_47652,N_32626,N_34868);
or U47653 (N_47653,N_32410,N_34816);
nand U47654 (N_47654,N_34784,N_38075);
or U47655 (N_47655,N_38854,N_38496);
or U47656 (N_47656,N_33909,N_38528);
and U47657 (N_47657,N_34991,N_35746);
or U47658 (N_47658,N_39779,N_31681);
nor U47659 (N_47659,N_32142,N_35478);
or U47660 (N_47660,N_33061,N_32106);
and U47661 (N_47661,N_38186,N_37409);
xor U47662 (N_47662,N_32239,N_36233);
or U47663 (N_47663,N_33200,N_32471);
and U47664 (N_47664,N_38020,N_36560);
nor U47665 (N_47665,N_33343,N_30602);
or U47666 (N_47666,N_37589,N_39906);
nand U47667 (N_47667,N_38641,N_36619);
xor U47668 (N_47668,N_38305,N_34640);
nand U47669 (N_47669,N_30505,N_34843);
nor U47670 (N_47670,N_38399,N_36714);
and U47671 (N_47671,N_37275,N_32142);
nand U47672 (N_47672,N_39314,N_39357);
or U47673 (N_47673,N_31817,N_36063);
nand U47674 (N_47674,N_39718,N_31911);
and U47675 (N_47675,N_30360,N_34825);
or U47676 (N_47676,N_33799,N_36106);
nand U47677 (N_47677,N_36380,N_31700);
and U47678 (N_47678,N_35701,N_34445);
or U47679 (N_47679,N_39797,N_35200);
nand U47680 (N_47680,N_38330,N_31940);
nand U47681 (N_47681,N_37384,N_38100);
nand U47682 (N_47682,N_32845,N_38296);
and U47683 (N_47683,N_32775,N_31931);
nand U47684 (N_47684,N_38413,N_39472);
and U47685 (N_47685,N_33649,N_33830);
nor U47686 (N_47686,N_31451,N_36575);
xor U47687 (N_47687,N_37985,N_30913);
xor U47688 (N_47688,N_38950,N_34100);
nor U47689 (N_47689,N_31186,N_37286);
xor U47690 (N_47690,N_39851,N_34839);
nand U47691 (N_47691,N_30841,N_34665);
nand U47692 (N_47692,N_32055,N_35382);
or U47693 (N_47693,N_32990,N_30817);
nand U47694 (N_47694,N_34888,N_32721);
xor U47695 (N_47695,N_36958,N_34671);
and U47696 (N_47696,N_34736,N_37625);
or U47697 (N_47697,N_33337,N_35999);
nand U47698 (N_47698,N_31519,N_33422);
nand U47699 (N_47699,N_33853,N_38926);
or U47700 (N_47700,N_32058,N_33824);
nor U47701 (N_47701,N_39987,N_34671);
nand U47702 (N_47702,N_38762,N_30586);
nor U47703 (N_47703,N_30824,N_32509);
or U47704 (N_47704,N_34892,N_34029);
and U47705 (N_47705,N_35347,N_37042);
and U47706 (N_47706,N_31140,N_36480);
nand U47707 (N_47707,N_35564,N_35973);
nand U47708 (N_47708,N_34238,N_37542);
or U47709 (N_47709,N_32957,N_30957);
or U47710 (N_47710,N_39208,N_38902);
nand U47711 (N_47711,N_38081,N_30990);
xnor U47712 (N_47712,N_31115,N_31629);
xnor U47713 (N_47713,N_36186,N_38796);
xnor U47714 (N_47714,N_33218,N_38383);
and U47715 (N_47715,N_36088,N_38590);
xor U47716 (N_47716,N_39792,N_36699);
or U47717 (N_47717,N_30773,N_37090);
or U47718 (N_47718,N_33708,N_38347);
and U47719 (N_47719,N_34636,N_38716);
nor U47720 (N_47720,N_36761,N_39136);
xor U47721 (N_47721,N_34006,N_31360);
xor U47722 (N_47722,N_31821,N_37345);
or U47723 (N_47723,N_31711,N_39421);
or U47724 (N_47724,N_35329,N_35880);
and U47725 (N_47725,N_38015,N_33108);
and U47726 (N_47726,N_30326,N_30579);
nand U47727 (N_47727,N_35588,N_39433);
and U47728 (N_47728,N_36188,N_35864);
and U47729 (N_47729,N_30503,N_31334);
xor U47730 (N_47730,N_34961,N_30144);
nor U47731 (N_47731,N_33527,N_39595);
nor U47732 (N_47732,N_35703,N_36087);
nand U47733 (N_47733,N_39319,N_39602);
nand U47734 (N_47734,N_30474,N_31103);
and U47735 (N_47735,N_39463,N_30718);
nor U47736 (N_47736,N_39741,N_35809);
nand U47737 (N_47737,N_32074,N_37080);
nand U47738 (N_47738,N_33858,N_35362);
or U47739 (N_47739,N_30222,N_31583);
and U47740 (N_47740,N_39333,N_39397);
and U47741 (N_47741,N_32724,N_38087);
or U47742 (N_47742,N_33727,N_31988);
or U47743 (N_47743,N_30014,N_33052);
nand U47744 (N_47744,N_36262,N_33338);
or U47745 (N_47745,N_33899,N_36971);
and U47746 (N_47746,N_36818,N_36543);
or U47747 (N_47747,N_33554,N_32425);
nor U47748 (N_47748,N_39779,N_35786);
and U47749 (N_47749,N_39436,N_30223);
nor U47750 (N_47750,N_34274,N_32243);
or U47751 (N_47751,N_31007,N_30636);
xnor U47752 (N_47752,N_31959,N_33904);
nand U47753 (N_47753,N_30083,N_36988);
or U47754 (N_47754,N_32106,N_33409);
nand U47755 (N_47755,N_36045,N_32028);
nand U47756 (N_47756,N_36145,N_31519);
and U47757 (N_47757,N_33888,N_37026);
nand U47758 (N_47758,N_33647,N_31128);
and U47759 (N_47759,N_34541,N_38160);
and U47760 (N_47760,N_33369,N_36453);
xor U47761 (N_47761,N_34091,N_32819);
and U47762 (N_47762,N_35412,N_39804);
or U47763 (N_47763,N_34301,N_35670);
or U47764 (N_47764,N_36752,N_33946);
and U47765 (N_47765,N_33108,N_36339);
nand U47766 (N_47766,N_33870,N_31576);
or U47767 (N_47767,N_30578,N_36040);
nand U47768 (N_47768,N_36919,N_32847);
or U47769 (N_47769,N_35659,N_38100);
or U47770 (N_47770,N_34052,N_34636);
nand U47771 (N_47771,N_38117,N_39669);
nand U47772 (N_47772,N_38825,N_34976);
and U47773 (N_47773,N_38717,N_39452);
nand U47774 (N_47774,N_36456,N_37251);
and U47775 (N_47775,N_35891,N_38179);
xor U47776 (N_47776,N_32834,N_39250);
nand U47777 (N_47777,N_30015,N_39763);
nand U47778 (N_47778,N_34935,N_31241);
nand U47779 (N_47779,N_39171,N_35526);
nand U47780 (N_47780,N_31943,N_34496);
nor U47781 (N_47781,N_36175,N_32032);
nor U47782 (N_47782,N_34454,N_36089);
or U47783 (N_47783,N_30683,N_38803);
xnor U47784 (N_47784,N_31353,N_30838);
nor U47785 (N_47785,N_38967,N_34327);
and U47786 (N_47786,N_31190,N_34282);
or U47787 (N_47787,N_32208,N_35504);
or U47788 (N_47788,N_31558,N_31576);
nand U47789 (N_47789,N_33285,N_32863);
and U47790 (N_47790,N_34732,N_31135);
nand U47791 (N_47791,N_39079,N_31155);
or U47792 (N_47792,N_39646,N_30367);
nor U47793 (N_47793,N_37028,N_34388);
nand U47794 (N_47794,N_34031,N_37443);
nand U47795 (N_47795,N_37445,N_39015);
nor U47796 (N_47796,N_38155,N_37634);
or U47797 (N_47797,N_32772,N_36260);
nand U47798 (N_47798,N_37411,N_35702);
or U47799 (N_47799,N_38856,N_33820);
or U47800 (N_47800,N_33127,N_33728);
or U47801 (N_47801,N_32354,N_34373);
nor U47802 (N_47802,N_32259,N_31064);
and U47803 (N_47803,N_39578,N_39867);
or U47804 (N_47804,N_33838,N_39268);
nor U47805 (N_47805,N_30398,N_38087);
nor U47806 (N_47806,N_30883,N_36584);
nor U47807 (N_47807,N_35261,N_31488);
nor U47808 (N_47808,N_34256,N_34128);
and U47809 (N_47809,N_36583,N_35125);
nor U47810 (N_47810,N_37477,N_37925);
xnor U47811 (N_47811,N_36350,N_39113);
nor U47812 (N_47812,N_31186,N_32286);
and U47813 (N_47813,N_31102,N_36257);
nand U47814 (N_47814,N_34763,N_38677);
and U47815 (N_47815,N_36841,N_30966);
xor U47816 (N_47816,N_35484,N_32491);
nand U47817 (N_47817,N_37277,N_31668);
and U47818 (N_47818,N_32853,N_39966);
or U47819 (N_47819,N_39799,N_39481);
or U47820 (N_47820,N_37074,N_35700);
nor U47821 (N_47821,N_37435,N_37536);
or U47822 (N_47822,N_31466,N_32276);
nor U47823 (N_47823,N_30001,N_32973);
nor U47824 (N_47824,N_34176,N_33986);
nor U47825 (N_47825,N_31059,N_33886);
nor U47826 (N_47826,N_38930,N_37422);
nand U47827 (N_47827,N_35462,N_33060);
and U47828 (N_47828,N_30149,N_31903);
or U47829 (N_47829,N_39272,N_36251);
and U47830 (N_47830,N_37286,N_37669);
and U47831 (N_47831,N_32705,N_33888);
nor U47832 (N_47832,N_34475,N_38075);
and U47833 (N_47833,N_34448,N_38980);
and U47834 (N_47834,N_37959,N_31897);
and U47835 (N_47835,N_32658,N_39220);
or U47836 (N_47836,N_38578,N_34064);
nor U47837 (N_47837,N_36108,N_32671);
nor U47838 (N_47838,N_33310,N_35158);
nand U47839 (N_47839,N_39101,N_36289);
nor U47840 (N_47840,N_39810,N_32103);
nand U47841 (N_47841,N_31015,N_34101);
and U47842 (N_47842,N_35849,N_34895);
nor U47843 (N_47843,N_38949,N_30489);
nand U47844 (N_47844,N_30141,N_33983);
nor U47845 (N_47845,N_38697,N_38249);
nand U47846 (N_47846,N_38059,N_33418);
nor U47847 (N_47847,N_38843,N_35132);
and U47848 (N_47848,N_38873,N_34227);
xor U47849 (N_47849,N_38780,N_30057);
nor U47850 (N_47850,N_33918,N_35375);
and U47851 (N_47851,N_38833,N_34072);
or U47852 (N_47852,N_31955,N_37565);
nor U47853 (N_47853,N_31341,N_32639);
and U47854 (N_47854,N_38101,N_35520);
nand U47855 (N_47855,N_30177,N_34871);
nand U47856 (N_47856,N_32255,N_37145);
or U47857 (N_47857,N_36883,N_39477);
nor U47858 (N_47858,N_39305,N_37000);
and U47859 (N_47859,N_33815,N_30359);
and U47860 (N_47860,N_37446,N_32425);
nor U47861 (N_47861,N_38482,N_36709);
nand U47862 (N_47862,N_33933,N_39149);
nand U47863 (N_47863,N_34886,N_35589);
and U47864 (N_47864,N_31294,N_35492);
or U47865 (N_47865,N_32929,N_37039);
and U47866 (N_47866,N_36128,N_37495);
and U47867 (N_47867,N_30574,N_30450);
nand U47868 (N_47868,N_33473,N_34282);
nor U47869 (N_47869,N_36648,N_37270);
nor U47870 (N_47870,N_30814,N_36472);
and U47871 (N_47871,N_32992,N_34270);
nor U47872 (N_47872,N_36415,N_36276);
nor U47873 (N_47873,N_39226,N_38006);
or U47874 (N_47874,N_39363,N_37715);
nand U47875 (N_47875,N_31096,N_35967);
and U47876 (N_47876,N_37006,N_31670);
nor U47877 (N_47877,N_36471,N_32625);
or U47878 (N_47878,N_37340,N_32207);
or U47879 (N_47879,N_38586,N_37304);
xor U47880 (N_47880,N_37979,N_39933);
xor U47881 (N_47881,N_35017,N_39377);
nor U47882 (N_47882,N_38684,N_32687);
nor U47883 (N_47883,N_37540,N_38988);
xnor U47884 (N_47884,N_36435,N_35482);
nor U47885 (N_47885,N_32713,N_30096);
nand U47886 (N_47886,N_32284,N_32626);
nand U47887 (N_47887,N_32583,N_33712);
xnor U47888 (N_47888,N_36899,N_39652);
and U47889 (N_47889,N_35019,N_39967);
or U47890 (N_47890,N_33521,N_34778);
nand U47891 (N_47891,N_37703,N_33517);
or U47892 (N_47892,N_37210,N_33384);
or U47893 (N_47893,N_39165,N_34181);
and U47894 (N_47894,N_36028,N_32365);
and U47895 (N_47895,N_38312,N_35559);
or U47896 (N_47896,N_38517,N_30846);
or U47897 (N_47897,N_39685,N_31583);
and U47898 (N_47898,N_33549,N_31243);
nand U47899 (N_47899,N_32312,N_38462);
nor U47900 (N_47900,N_32947,N_35240);
nor U47901 (N_47901,N_37854,N_37291);
and U47902 (N_47902,N_38108,N_35385);
nor U47903 (N_47903,N_30509,N_31608);
nand U47904 (N_47904,N_36961,N_39055);
and U47905 (N_47905,N_30109,N_32633);
xnor U47906 (N_47906,N_32558,N_36730);
nand U47907 (N_47907,N_30059,N_34519);
or U47908 (N_47908,N_39832,N_38120);
nor U47909 (N_47909,N_32846,N_35028);
and U47910 (N_47910,N_36374,N_38604);
nand U47911 (N_47911,N_38405,N_34663);
nand U47912 (N_47912,N_34128,N_34724);
nand U47913 (N_47913,N_30266,N_36822);
and U47914 (N_47914,N_39598,N_36645);
nand U47915 (N_47915,N_33663,N_37261);
nand U47916 (N_47916,N_33746,N_37672);
nand U47917 (N_47917,N_33684,N_38883);
and U47918 (N_47918,N_38479,N_33726);
or U47919 (N_47919,N_31203,N_36590);
or U47920 (N_47920,N_30180,N_30073);
nand U47921 (N_47921,N_31020,N_32590);
nor U47922 (N_47922,N_35781,N_34324);
nor U47923 (N_47923,N_35874,N_32511);
or U47924 (N_47924,N_37499,N_36587);
and U47925 (N_47925,N_35037,N_31050);
or U47926 (N_47926,N_33136,N_36485);
nor U47927 (N_47927,N_39969,N_33368);
nor U47928 (N_47928,N_36827,N_31384);
or U47929 (N_47929,N_30340,N_32578);
xor U47930 (N_47930,N_37237,N_37193);
nor U47931 (N_47931,N_33580,N_30086);
nor U47932 (N_47932,N_33905,N_31182);
xor U47933 (N_47933,N_38435,N_36183);
nor U47934 (N_47934,N_39496,N_35356);
xnor U47935 (N_47935,N_34792,N_33486);
nor U47936 (N_47936,N_34667,N_33734);
nor U47937 (N_47937,N_33269,N_39933);
nand U47938 (N_47938,N_34398,N_34361);
and U47939 (N_47939,N_37990,N_36019);
nor U47940 (N_47940,N_39899,N_31194);
and U47941 (N_47941,N_39849,N_37473);
nand U47942 (N_47942,N_35640,N_31605);
nor U47943 (N_47943,N_32267,N_37135);
or U47944 (N_47944,N_31003,N_30587);
nand U47945 (N_47945,N_38556,N_32626);
or U47946 (N_47946,N_32623,N_32492);
and U47947 (N_47947,N_38036,N_37619);
and U47948 (N_47948,N_37723,N_34287);
nand U47949 (N_47949,N_39794,N_30417);
nor U47950 (N_47950,N_35821,N_36967);
and U47951 (N_47951,N_35229,N_30814);
nor U47952 (N_47952,N_39643,N_38740);
or U47953 (N_47953,N_38507,N_35084);
xor U47954 (N_47954,N_38990,N_36883);
or U47955 (N_47955,N_33675,N_34143);
nand U47956 (N_47956,N_37233,N_34848);
nor U47957 (N_47957,N_30354,N_35970);
nor U47958 (N_47958,N_31398,N_34954);
and U47959 (N_47959,N_37713,N_39711);
nor U47960 (N_47960,N_39091,N_36973);
nand U47961 (N_47961,N_36719,N_31532);
and U47962 (N_47962,N_35656,N_37120);
nand U47963 (N_47963,N_38338,N_31797);
nor U47964 (N_47964,N_37472,N_37881);
and U47965 (N_47965,N_32537,N_34649);
and U47966 (N_47966,N_39123,N_32904);
nand U47967 (N_47967,N_37891,N_35522);
xor U47968 (N_47968,N_35569,N_37458);
and U47969 (N_47969,N_36106,N_34150);
nand U47970 (N_47970,N_35347,N_35942);
nand U47971 (N_47971,N_34105,N_39979);
or U47972 (N_47972,N_35713,N_39004);
nand U47973 (N_47973,N_39060,N_30307);
nand U47974 (N_47974,N_34566,N_31036);
and U47975 (N_47975,N_34516,N_32364);
nand U47976 (N_47976,N_39392,N_38036);
or U47977 (N_47977,N_32637,N_37774);
nor U47978 (N_47978,N_35042,N_37928);
or U47979 (N_47979,N_36195,N_34972);
nor U47980 (N_47980,N_30874,N_30900);
and U47981 (N_47981,N_39173,N_33237);
nor U47982 (N_47982,N_31266,N_32669);
or U47983 (N_47983,N_31982,N_38375);
nand U47984 (N_47984,N_34219,N_37392);
xnor U47985 (N_47985,N_36505,N_33113);
or U47986 (N_47986,N_30316,N_33862);
or U47987 (N_47987,N_31536,N_35498);
xor U47988 (N_47988,N_35089,N_31206);
nor U47989 (N_47989,N_36081,N_32443);
or U47990 (N_47990,N_32279,N_38483);
or U47991 (N_47991,N_31332,N_32167);
nand U47992 (N_47992,N_34246,N_31766);
and U47993 (N_47993,N_32069,N_37456);
or U47994 (N_47994,N_38925,N_36982);
and U47995 (N_47995,N_39888,N_31230);
nor U47996 (N_47996,N_33880,N_36392);
or U47997 (N_47997,N_32435,N_38527);
xnor U47998 (N_47998,N_31907,N_34361);
nor U47999 (N_47999,N_37688,N_32882);
nand U48000 (N_48000,N_31955,N_38045);
nand U48001 (N_48001,N_32067,N_36107);
and U48002 (N_48002,N_39159,N_37612);
nand U48003 (N_48003,N_32145,N_31238);
nand U48004 (N_48004,N_37380,N_38212);
and U48005 (N_48005,N_38608,N_34888);
nor U48006 (N_48006,N_33845,N_38252);
or U48007 (N_48007,N_32392,N_34022);
nor U48008 (N_48008,N_33349,N_32205);
nor U48009 (N_48009,N_34410,N_39492);
and U48010 (N_48010,N_37375,N_30763);
xor U48011 (N_48011,N_34586,N_37039);
and U48012 (N_48012,N_31894,N_32036);
or U48013 (N_48013,N_38297,N_32596);
nand U48014 (N_48014,N_38794,N_32419);
xor U48015 (N_48015,N_37558,N_36976);
or U48016 (N_48016,N_37488,N_30466);
nor U48017 (N_48017,N_35875,N_30978);
or U48018 (N_48018,N_37555,N_36275);
or U48019 (N_48019,N_37909,N_39522);
xnor U48020 (N_48020,N_39815,N_39256);
nand U48021 (N_48021,N_38865,N_33818);
nor U48022 (N_48022,N_38355,N_30297);
and U48023 (N_48023,N_39162,N_32257);
or U48024 (N_48024,N_36870,N_33205);
and U48025 (N_48025,N_32192,N_37026);
and U48026 (N_48026,N_30013,N_30611);
or U48027 (N_48027,N_31316,N_31825);
xnor U48028 (N_48028,N_37363,N_35431);
nand U48029 (N_48029,N_35689,N_32546);
or U48030 (N_48030,N_37489,N_32270);
nand U48031 (N_48031,N_34858,N_31093);
nor U48032 (N_48032,N_39634,N_35728);
or U48033 (N_48033,N_30779,N_36952);
and U48034 (N_48034,N_31472,N_30563);
or U48035 (N_48035,N_35966,N_35033);
nor U48036 (N_48036,N_39310,N_33060);
nand U48037 (N_48037,N_39440,N_33351);
nor U48038 (N_48038,N_34064,N_32978);
and U48039 (N_48039,N_33095,N_38380);
nor U48040 (N_48040,N_39483,N_39720);
and U48041 (N_48041,N_34911,N_38302);
or U48042 (N_48042,N_38796,N_31159);
or U48043 (N_48043,N_37141,N_33530);
and U48044 (N_48044,N_32527,N_37361);
nor U48045 (N_48045,N_38059,N_31769);
and U48046 (N_48046,N_36918,N_36767);
and U48047 (N_48047,N_31042,N_39086);
nor U48048 (N_48048,N_34840,N_37332);
and U48049 (N_48049,N_38755,N_38879);
nor U48050 (N_48050,N_33771,N_35371);
nor U48051 (N_48051,N_35060,N_30486);
or U48052 (N_48052,N_32854,N_30583);
or U48053 (N_48053,N_36524,N_35146);
or U48054 (N_48054,N_31000,N_33889);
nor U48055 (N_48055,N_37465,N_31526);
xor U48056 (N_48056,N_32760,N_31305);
nor U48057 (N_48057,N_39540,N_39269);
or U48058 (N_48058,N_36256,N_31918);
or U48059 (N_48059,N_31775,N_39671);
nand U48060 (N_48060,N_37059,N_34687);
nor U48061 (N_48061,N_35837,N_36835);
and U48062 (N_48062,N_37018,N_38635);
xnor U48063 (N_48063,N_30468,N_33958);
nor U48064 (N_48064,N_30924,N_31295);
and U48065 (N_48065,N_32006,N_30798);
and U48066 (N_48066,N_36583,N_36750);
nand U48067 (N_48067,N_30606,N_38011);
and U48068 (N_48068,N_36270,N_31618);
nor U48069 (N_48069,N_38546,N_31501);
nor U48070 (N_48070,N_36019,N_37838);
nand U48071 (N_48071,N_34887,N_34353);
nor U48072 (N_48072,N_33397,N_30913);
and U48073 (N_48073,N_33375,N_34096);
and U48074 (N_48074,N_33202,N_39625);
xor U48075 (N_48075,N_32669,N_31781);
xnor U48076 (N_48076,N_39490,N_39982);
nand U48077 (N_48077,N_30225,N_31475);
and U48078 (N_48078,N_34731,N_36651);
and U48079 (N_48079,N_32948,N_39346);
and U48080 (N_48080,N_36208,N_32518);
or U48081 (N_48081,N_30068,N_37300);
nor U48082 (N_48082,N_35904,N_31489);
or U48083 (N_48083,N_30000,N_38125);
nor U48084 (N_48084,N_39933,N_30598);
nor U48085 (N_48085,N_32142,N_31656);
or U48086 (N_48086,N_33271,N_32021);
and U48087 (N_48087,N_31361,N_31654);
and U48088 (N_48088,N_30723,N_35014);
or U48089 (N_48089,N_37430,N_37410);
xnor U48090 (N_48090,N_37943,N_32304);
and U48091 (N_48091,N_35422,N_35293);
or U48092 (N_48092,N_35194,N_35837);
nor U48093 (N_48093,N_36305,N_37349);
or U48094 (N_48094,N_35477,N_33650);
nand U48095 (N_48095,N_37464,N_32944);
or U48096 (N_48096,N_35013,N_39524);
and U48097 (N_48097,N_37639,N_38604);
or U48098 (N_48098,N_36834,N_30523);
nand U48099 (N_48099,N_39553,N_34047);
xnor U48100 (N_48100,N_30852,N_35322);
xor U48101 (N_48101,N_33963,N_37624);
nor U48102 (N_48102,N_37538,N_30648);
nand U48103 (N_48103,N_38138,N_39254);
and U48104 (N_48104,N_31995,N_33686);
and U48105 (N_48105,N_35786,N_33314);
xor U48106 (N_48106,N_33706,N_38724);
nor U48107 (N_48107,N_33469,N_31759);
nor U48108 (N_48108,N_36167,N_31725);
nand U48109 (N_48109,N_33701,N_32164);
nor U48110 (N_48110,N_35040,N_37098);
and U48111 (N_48111,N_30620,N_33788);
xor U48112 (N_48112,N_37014,N_32707);
or U48113 (N_48113,N_35322,N_36677);
nand U48114 (N_48114,N_37849,N_33909);
xor U48115 (N_48115,N_35698,N_34245);
and U48116 (N_48116,N_38274,N_34008);
or U48117 (N_48117,N_37100,N_37013);
xor U48118 (N_48118,N_39354,N_31952);
or U48119 (N_48119,N_39004,N_32577);
nand U48120 (N_48120,N_35769,N_33097);
and U48121 (N_48121,N_38673,N_39526);
and U48122 (N_48122,N_39449,N_30087);
or U48123 (N_48123,N_39908,N_38820);
nand U48124 (N_48124,N_32951,N_35860);
and U48125 (N_48125,N_30830,N_31494);
or U48126 (N_48126,N_38633,N_37142);
nor U48127 (N_48127,N_34362,N_30230);
or U48128 (N_48128,N_30494,N_30241);
nand U48129 (N_48129,N_36643,N_36605);
xnor U48130 (N_48130,N_30856,N_38876);
nor U48131 (N_48131,N_33495,N_38259);
and U48132 (N_48132,N_34255,N_30981);
and U48133 (N_48133,N_38030,N_32922);
and U48134 (N_48134,N_35957,N_30261);
or U48135 (N_48135,N_30916,N_33211);
xor U48136 (N_48136,N_31274,N_34372);
xnor U48137 (N_48137,N_37750,N_37122);
or U48138 (N_48138,N_39383,N_39032);
and U48139 (N_48139,N_31086,N_32295);
and U48140 (N_48140,N_38681,N_30512);
nand U48141 (N_48141,N_32077,N_39551);
xnor U48142 (N_48142,N_35775,N_38109);
nor U48143 (N_48143,N_31033,N_31371);
nand U48144 (N_48144,N_33688,N_32290);
or U48145 (N_48145,N_34895,N_30614);
nand U48146 (N_48146,N_39161,N_37045);
or U48147 (N_48147,N_38212,N_38507);
xor U48148 (N_48148,N_36930,N_37715);
nor U48149 (N_48149,N_33019,N_39304);
nor U48150 (N_48150,N_37687,N_31608);
and U48151 (N_48151,N_39467,N_39399);
nand U48152 (N_48152,N_39680,N_38244);
or U48153 (N_48153,N_30450,N_34286);
or U48154 (N_48154,N_32693,N_30077);
and U48155 (N_48155,N_34721,N_30441);
or U48156 (N_48156,N_39726,N_32712);
xor U48157 (N_48157,N_37368,N_35062);
nand U48158 (N_48158,N_34315,N_31391);
or U48159 (N_48159,N_37591,N_37468);
and U48160 (N_48160,N_33676,N_33326);
xor U48161 (N_48161,N_35561,N_30084);
nand U48162 (N_48162,N_37163,N_36947);
and U48163 (N_48163,N_31330,N_34564);
nand U48164 (N_48164,N_34272,N_38711);
nand U48165 (N_48165,N_37714,N_30442);
nand U48166 (N_48166,N_35666,N_36707);
nor U48167 (N_48167,N_30720,N_37789);
or U48168 (N_48168,N_32612,N_31225);
xnor U48169 (N_48169,N_32721,N_32644);
nor U48170 (N_48170,N_35563,N_31078);
nand U48171 (N_48171,N_37099,N_39035);
or U48172 (N_48172,N_35225,N_37663);
or U48173 (N_48173,N_33073,N_30075);
nand U48174 (N_48174,N_37794,N_39159);
nor U48175 (N_48175,N_31820,N_37619);
and U48176 (N_48176,N_31571,N_31779);
nand U48177 (N_48177,N_32705,N_35087);
nor U48178 (N_48178,N_38613,N_37145);
nor U48179 (N_48179,N_39848,N_39018);
xnor U48180 (N_48180,N_31874,N_38169);
and U48181 (N_48181,N_32287,N_37038);
nand U48182 (N_48182,N_36215,N_32552);
nand U48183 (N_48183,N_32947,N_37567);
xnor U48184 (N_48184,N_31553,N_31128);
or U48185 (N_48185,N_34246,N_38375);
and U48186 (N_48186,N_34463,N_35951);
nor U48187 (N_48187,N_30454,N_38766);
nor U48188 (N_48188,N_30086,N_37617);
and U48189 (N_48189,N_32139,N_31972);
and U48190 (N_48190,N_30594,N_30448);
and U48191 (N_48191,N_36246,N_39562);
nor U48192 (N_48192,N_35579,N_35240);
xor U48193 (N_48193,N_36164,N_30885);
xnor U48194 (N_48194,N_38250,N_37982);
and U48195 (N_48195,N_37961,N_37422);
or U48196 (N_48196,N_30355,N_37243);
or U48197 (N_48197,N_30555,N_39783);
or U48198 (N_48198,N_38504,N_32659);
or U48199 (N_48199,N_31487,N_30869);
nor U48200 (N_48200,N_34187,N_39618);
and U48201 (N_48201,N_33255,N_39315);
and U48202 (N_48202,N_33018,N_35107);
nor U48203 (N_48203,N_37042,N_33492);
nor U48204 (N_48204,N_35416,N_32142);
nand U48205 (N_48205,N_30435,N_35968);
xor U48206 (N_48206,N_34274,N_31703);
or U48207 (N_48207,N_38487,N_35211);
and U48208 (N_48208,N_32347,N_32836);
and U48209 (N_48209,N_31853,N_36462);
nor U48210 (N_48210,N_31182,N_34848);
or U48211 (N_48211,N_34481,N_31209);
or U48212 (N_48212,N_36812,N_35234);
nand U48213 (N_48213,N_36387,N_34810);
nand U48214 (N_48214,N_33763,N_30097);
and U48215 (N_48215,N_31566,N_30574);
nand U48216 (N_48216,N_32440,N_33706);
nand U48217 (N_48217,N_32959,N_38730);
or U48218 (N_48218,N_33448,N_39483);
and U48219 (N_48219,N_37022,N_33263);
xnor U48220 (N_48220,N_39575,N_34615);
nor U48221 (N_48221,N_35193,N_37937);
nand U48222 (N_48222,N_35480,N_30435);
or U48223 (N_48223,N_35722,N_33043);
and U48224 (N_48224,N_30438,N_33899);
or U48225 (N_48225,N_33175,N_35732);
and U48226 (N_48226,N_33359,N_33345);
xnor U48227 (N_48227,N_39625,N_34353);
and U48228 (N_48228,N_36941,N_30883);
or U48229 (N_48229,N_34565,N_32756);
or U48230 (N_48230,N_34590,N_34373);
nand U48231 (N_48231,N_37107,N_30560);
xnor U48232 (N_48232,N_39384,N_39304);
xor U48233 (N_48233,N_39511,N_34873);
or U48234 (N_48234,N_35048,N_35683);
nor U48235 (N_48235,N_38994,N_38581);
nand U48236 (N_48236,N_39275,N_34961);
or U48237 (N_48237,N_32347,N_33191);
xor U48238 (N_48238,N_31607,N_38067);
nor U48239 (N_48239,N_30744,N_30419);
or U48240 (N_48240,N_35613,N_35272);
nor U48241 (N_48241,N_39611,N_32196);
and U48242 (N_48242,N_39563,N_39343);
nand U48243 (N_48243,N_34809,N_39194);
xnor U48244 (N_48244,N_35607,N_35261);
nor U48245 (N_48245,N_32058,N_35445);
or U48246 (N_48246,N_34331,N_32087);
or U48247 (N_48247,N_31049,N_39769);
nand U48248 (N_48248,N_30716,N_36992);
nand U48249 (N_48249,N_30832,N_31665);
or U48250 (N_48250,N_36668,N_38931);
nor U48251 (N_48251,N_38938,N_34034);
or U48252 (N_48252,N_34661,N_39853);
nand U48253 (N_48253,N_31249,N_32583);
and U48254 (N_48254,N_33909,N_30064);
nor U48255 (N_48255,N_34505,N_36975);
xor U48256 (N_48256,N_36455,N_39159);
nor U48257 (N_48257,N_30023,N_31686);
and U48258 (N_48258,N_35205,N_30212);
nand U48259 (N_48259,N_36757,N_31142);
nand U48260 (N_48260,N_39739,N_30444);
nor U48261 (N_48261,N_30707,N_35102);
and U48262 (N_48262,N_35087,N_32567);
nand U48263 (N_48263,N_36953,N_37050);
nand U48264 (N_48264,N_36855,N_38298);
or U48265 (N_48265,N_39892,N_30415);
and U48266 (N_48266,N_32048,N_37272);
or U48267 (N_48267,N_35532,N_35492);
xnor U48268 (N_48268,N_36377,N_32450);
or U48269 (N_48269,N_39318,N_31732);
or U48270 (N_48270,N_33818,N_38526);
or U48271 (N_48271,N_33918,N_33295);
or U48272 (N_48272,N_38694,N_35903);
and U48273 (N_48273,N_35907,N_39041);
and U48274 (N_48274,N_39643,N_37884);
nand U48275 (N_48275,N_36138,N_35561);
nor U48276 (N_48276,N_30667,N_30551);
and U48277 (N_48277,N_36565,N_34683);
or U48278 (N_48278,N_33412,N_30889);
or U48279 (N_48279,N_30516,N_33612);
and U48280 (N_48280,N_39437,N_31983);
or U48281 (N_48281,N_30267,N_39169);
nand U48282 (N_48282,N_30382,N_39883);
nand U48283 (N_48283,N_31465,N_30676);
and U48284 (N_48284,N_35592,N_36994);
or U48285 (N_48285,N_35287,N_32591);
or U48286 (N_48286,N_30049,N_33875);
nor U48287 (N_48287,N_38517,N_33929);
nand U48288 (N_48288,N_33069,N_31248);
nor U48289 (N_48289,N_30101,N_39076);
nand U48290 (N_48290,N_37179,N_34645);
and U48291 (N_48291,N_30707,N_36908);
nand U48292 (N_48292,N_38932,N_38218);
nand U48293 (N_48293,N_30490,N_30018);
and U48294 (N_48294,N_34094,N_36146);
and U48295 (N_48295,N_36776,N_38967);
and U48296 (N_48296,N_38124,N_34545);
or U48297 (N_48297,N_33639,N_33404);
nor U48298 (N_48298,N_37106,N_36582);
nand U48299 (N_48299,N_32755,N_30389);
and U48300 (N_48300,N_32506,N_30951);
or U48301 (N_48301,N_38962,N_37205);
nand U48302 (N_48302,N_35157,N_31676);
nor U48303 (N_48303,N_32039,N_35314);
and U48304 (N_48304,N_39786,N_34616);
nor U48305 (N_48305,N_31429,N_38910);
xnor U48306 (N_48306,N_34204,N_33324);
and U48307 (N_48307,N_38283,N_31249);
nand U48308 (N_48308,N_30982,N_39685);
nor U48309 (N_48309,N_39485,N_37669);
nor U48310 (N_48310,N_35931,N_35590);
or U48311 (N_48311,N_37134,N_37035);
nor U48312 (N_48312,N_32368,N_37545);
or U48313 (N_48313,N_39561,N_39811);
and U48314 (N_48314,N_32343,N_31295);
nand U48315 (N_48315,N_35279,N_39275);
and U48316 (N_48316,N_30428,N_34521);
xnor U48317 (N_48317,N_35526,N_37643);
nand U48318 (N_48318,N_31822,N_35966);
or U48319 (N_48319,N_37139,N_31036);
and U48320 (N_48320,N_37447,N_35393);
nand U48321 (N_48321,N_33106,N_33935);
nor U48322 (N_48322,N_39909,N_37858);
nor U48323 (N_48323,N_31515,N_37973);
nand U48324 (N_48324,N_38363,N_36080);
and U48325 (N_48325,N_30315,N_34198);
nand U48326 (N_48326,N_34238,N_32754);
xnor U48327 (N_48327,N_34232,N_39323);
nor U48328 (N_48328,N_38149,N_35617);
nand U48329 (N_48329,N_39606,N_37760);
nand U48330 (N_48330,N_38815,N_36730);
nor U48331 (N_48331,N_38544,N_34615);
or U48332 (N_48332,N_37009,N_31532);
nor U48333 (N_48333,N_35600,N_32987);
or U48334 (N_48334,N_34173,N_35112);
or U48335 (N_48335,N_36277,N_34329);
nor U48336 (N_48336,N_38550,N_36081);
and U48337 (N_48337,N_30535,N_38302);
nor U48338 (N_48338,N_30082,N_35444);
and U48339 (N_48339,N_34666,N_38534);
or U48340 (N_48340,N_30221,N_39561);
nand U48341 (N_48341,N_33418,N_38203);
xnor U48342 (N_48342,N_31281,N_34602);
and U48343 (N_48343,N_35696,N_39486);
or U48344 (N_48344,N_30094,N_36689);
nand U48345 (N_48345,N_36647,N_37499);
nand U48346 (N_48346,N_39299,N_33202);
nand U48347 (N_48347,N_34273,N_34577);
or U48348 (N_48348,N_33730,N_36410);
nand U48349 (N_48349,N_30871,N_37777);
and U48350 (N_48350,N_34337,N_31265);
and U48351 (N_48351,N_36055,N_34684);
nor U48352 (N_48352,N_38912,N_35902);
nand U48353 (N_48353,N_32478,N_34467);
or U48354 (N_48354,N_33881,N_34941);
nor U48355 (N_48355,N_37205,N_33318);
nand U48356 (N_48356,N_37285,N_35364);
nor U48357 (N_48357,N_33045,N_33892);
xor U48358 (N_48358,N_34694,N_31303);
or U48359 (N_48359,N_31250,N_37622);
xor U48360 (N_48360,N_36901,N_37122);
nor U48361 (N_48361,N_34215,N_38262);
nand U48362 (N_48362,N_36287,N_39329);
or U48363 (N_48363,N_38352,N_36533);
nor U48364 (N_48364,N_36697,N_34353);
nor U48365 (N_48365,N_31290,N_30008);
nor U48366 (N_48366,N_32130,N_30263);
and U48367 (N_48367,N_33357,N_30912);
or U48368 (N_48368,N_34962,N_34354);
or U48369 (N_48369,N_33030,N_37983);
or U48370 (N_48370,N_37891,N_30014);
nand U48371 (N_48371,N_35320,N_39806);
and U48372 (N_48372,N_32336,N_37570);
nand U48373 (N_48373,N_37357,N_36012);
and U48374 (N_48374,N_38827,N_30573);
and U48375 (N_48375,N_30824,N_31258);
xor U48376 (N_48376,N_36432,N_33363);
and U48377 (N_48377,N_33458,N_37697);
nor U48378 (N_48378,N_31372,N_32051);
xnor U48379 (N_48379,N_37776,N_31328);
or U48380 (N_48380,N_32608,N_36715);
nand U48381 (N_48381,N_34928,N_39138);
and U48382 (N_48382,N_39856,N_33852);
nor U48383 (N_48383,N_33023,N_38582);
or U48384 (N_48384,N_30018,N_33577);
nand U48385 (N_48385,N_38785,N_38620);
xnor U48386 (N_48386,N_30349,N_39351);
xor U48387 (N_48387,N_35618,N_37265);
nor U48388 (N_48388,N_39253,N_33289);
nor U48389 (N_48389,N_33169,N_37121);
or U48390 (N_48390,N_37785,N_38278);
nor U48391 (N_48391,N_35184,N_38232);
nand U48392 (N_48392,N_30093,N_38867);
nor U48393 (N_48393,N_35947,N_35867);
or U48394 (N_48394,N_30921,N_33644);
xnor U48395 (N_48395,N_36775,N_30068);
nand U48396 (N_48396,N_34840,N_37766);
and U48397 (N_48397,N_34474,N_33186);
nor U48398 (N_48398,N_30144,N_33283);
or U48399 (N_48399,N_36151,N_32953);
nand U48400 (N_48400,N_39041,N_37948);
or U48401 (N_48401,N_31630,N_30632);
or U48402 (N_48402,N_34800,N_33115);
or U48403 (N_48403,N_36388,N_30341);
nand U48404 (N_48404,N_30195,N_30979);
xor U48405 (N_48405,N_30960,N_30989);
xnor U48406 (N_48406,N_31648,N_38449);
xor U48407 (N_48407,N_33477,N_38965);
xnor U48408 (N_48408,N_32084,N_36899);
nor U48409 (N_48409,N_33337,N_34007);
or U48410 (N_48410,N_31138,N_36959);
and U48411 (N_48411,N_31666,N_36524);
or U48412 (N_48412,N_30227,N_35317);
nand U48413 (N_48413,N_30195,N_35817);
nand U48414 (N_48414,N_34359,N_38618);
nor U48415 (N_48415,N_36841,N_32634);
nor U48416 (N_48416,N_30097,N_39457);
nor U48417 (N_48417,N_36479,N_35892);
nor U48418 (N_48418,N_30970,N_31114);
xor U48419 (N_48419,N_32081,N_33235);
xor U48420 (N_48420,N_30979,N_38271);
and U48421 (N_48421,N_35725,N_30292);
or U48422 (N_48422,N_32150,N_33862);
nand U48423 (N_48423,N_38119,N_35919);
nor U48424 (N_48424,N_32230,N_31255);
nand U48425 (N_48425,N_35665,N_38139);
or U48426 (N_48426,N_38254,N_38423);
nor U48427 (N_48427,N_35409,N_32723);
nand U48428 (N_48428,N_34525,N_39732);
xor U48429 (N_48429,N_38925,N_34352);
or U48430 (N_48430,N_34097,N_35312);
nor U48431 (N_48431,N_36275,N_36272);
or U48432 (N_48432,N_32343,N_30153);
nor U48433 (N_48433,N_37949,N_34828);
or U48434 (N_48434,N_36008,N_33084);
nand U48435 (N_48435,N_37525,N_30883);
xnor U48436 (N_48436,N_37299,N_37636);
and U48437 (N_48437,N_34083,N_32088);
or U48438 (N_48438,N_36078,N_32863);
or U48439 (N_48439,N_33288,N_38275);
nor U48440 (N_48440,N_37288,N_36603);
or U48441 (N_48441,N_30705,N_37685);
nand U48442 (N_48442,N_36765,N_36427);
or U48443 (N_48443,N_37037,N_35518);
nand U48444 (N_48444,N_37345,N_37923);
and U48445 (N_48445,N_35594,N_32074);
nor U48446 (N_48446,N_35222,N_39621);
nor U48447 (N_48447,N_31929,N_39622);
or U48448 (N_48448,N_34269,N_31651);
nand U48449 (N_48449,N_30823,N_37444);
or U48450 (N_48450,N_34796,N_32825);
nand U48451 (N_48451,N_30396,N_36003);
nand U48452 (N_48452,N_39289,N_32450);
or U48453 (N_48453,N_38939,N_31284);
nand U48454 (N_48454,N_34085,N_31407);
and U48455 (N_48455,N_38900,N_35000);
and U48456 (N_48456,N_32928,N_33737);
nand U48457 (N_48457,N_39253,N_33241);
and U48458 (N_48458,N_32298,N_36371);
or U48459 (N_48459,N_39649,N_30130);
or U48460 (N_48460,N_30896,N_39795);
nand U48461 (N_48461,N_39763,N_32078);
and U48462 (N_48462,N_39831,N_39636);
nor U48463 (N_48463,N_30781,N_33031);
or U48464 (N_48464,N_39213,N_30959);
and U48465 (N_48465,N_34466,N_38184);
nand U48466 (N_48466,N_34504,N_30110);
xor U48467 (N_48467,N_34072,N_30748);
or U48468 (N_48468,N_35833,N_30662);
and U48469 (N_48469,N_38590,N_38709);
xor U48470 (N_48470,N_38300,N_30831);
xor U48471 (N_48471,N_33781,N_37586);
xnor U48472 (N_48472,N_30411,N_31486);
nor U48473 (N_48473,N_34211,N_34098);
nand U48474 (N_48474,N_32637,N_31599);
or U48475 (N_48475,N_33928,N_32565);
or U48476 (N_48476,N_30384,N_33024);
and U48477 (N_48477,N_34038,N_31372);
or U48478 (N_48478,N_31671,N_39881);
nand U48479 (N_48479,N_36729,N_35190);
nor U48480 (N_48480,N_38207,N_39781);
nand U48481 (N_48481,N_31493,N_32670);
nand U48482 (N_48482,N_33750,N_30189);
nand U48483 (N_48483,N_34983,N_36700);
nor U48484 (N_48484,N_38642,N_32425);
nor U48485 (N_48485,N_33067,N_34917);
or U48486 (N_48486,N_39594,N_32800);
nand U48487 (N_48487,N_33472,N_34963);
xnor U48488 (N_48488,N_32259,N_35902);
nor U48489 (N_48489,N_39713,N_38791);
nor U48490 (N_48490,N_39091,N_32105);
and U48491 (N_48491,N_32843,N_32063);
nor U48492 (N_48492,N_32230,N_38533);
and U48493 (N_48493,N_34041,N_33799);
or U48494 (N_48494,N_35953,N_36469);
and U48495 (N_48495,N_31624,N_30848);
nand U48496 (N_48496,N_37371,N_37454);
and U48497 (N_48497,N_34184,N_34639);
nor U48498 (N_48498,N_37415,N_34075);
or U48499 (N_48499,N_38448,N_39403);
nor U48500 (N_48500,N_31384,N_36308);
xor U48501 (N_48501,N_30819,N_30981);
or U48502 (N_48502,N_36148,N_37545);
and U48503 (N_48503,N_35790,N_32337);
or U48504 (N_48504,N_32599,N_33260);
nand U48505 (N_48505,N_37029,N_38433);
nand U48506 (N_48506,N_36983,N_32339);
nor U48507 (N_48507,N_34066,N_37059);
or U48508 (N_48508,N_31643,N_35320);
or U48509 (N_48509,N_31894,N_38463);
xnor U48510 (N_48510,N_36178,N_34785);
nor U48511 (N_48511,N_38678,N_36103);
nor U48512 (N_48512,N_34287,N_30645);
nand U48513 (N_48513,N_34530,N_32566);
nor U48514 (N_48514,N_34059,N_39539);
nand U48515 (N_48515,N_32410,N_37674);
xnor U48516 (N_48516,N_36721,N_35589);
and U48517 (N_48517,N_39110,N_39894);
xor U48518 (N_48518,N_31665,N_33996);
or U48519 (N_48519,N_36750,N_38436);
nand U48520 (N_48520,N_35264,N_39702);
or U48521 (N_48521,N_32207,N_30328);
nand U48522 (N_48522,N_38855,N_30836);
nand U48523 (N_48523,N_32388,N_32101);
nor U48524 (N_48524,N_33603,N_37692);
or U48525 (N_48525,N_31153,N_32036);
or U48526 (N_48526,N_39437,N_39977);
xnor U48527 (N_48527,N_38071,N_38310);
and U48528 (N_48528,N_31254,N_35268);
or U48529 (N_48529,N_36617,N_31220);
nand U48530 (N_48530,N_33794,N_31713);
nand U48531 (N_48531,N_38003,N_30927);
xnor U48532 (N_48532,N_36510,N_34508);
or U48533 (N_48533,N_31410,N_31579);
nor U48534 (N_48534,N_37864,N_32684);
or U48535 (N_48535,N_30140,N_31362);
and U48536 (N_48536,N_30516,N_31972);
or U48537 (N_48537,N_39596,N_32478);
nand U48538 (N_48538,N_33908,N_34662);
or U48539 (N_48539,N_39279,N_39167);
nand U48540 (N_48540,N_34208,N_36198);
and U48541 (N_48541,N_36003,N_37042);
and U48542 (N_48542,N_35225,N_31511);
and U48543 (N_48543,N_39805,N_38315);
or U48544 (N_48544,N_34343,N_33618);
nand U48545 (N_48545,N_38224,N_33379);
and U48546 (N_48546,N_38267,N_36793);
and U48547 (N_48547,N_32730,N_34521);
or U48548 (N_48548,N_39491,N_37014);
nor U48549 (N_48549,N_34766,N_37589);
or U48550 (N_48550,N_38427,N_36821);
and U48551 (N_48551,N_39176,N_36063);
or U48552 (N_48552,N_31739,N_32655);
or U48553 (N_48553,N_39054,N_32979);
nor U48554 (N_48554,N_37250,N_32730);
nor U48555 (N_48555,N_30594,N_38580);
xor U48556 (N_48556,N_39305,N_35907);
and U48557 (N_48557,N_32093,N_38336);
and U48558 (N_48558,N_33339,N_34851);
and U48559 (N_48559,N_31858,N_36011);
xnor U48560 (N_48560,N_31205,N_36620);
and U48561 (N_48561,N_33651,N_37405);
or U48562 (N_48562,N_31848,N_33123);
nand U48563 (N_48563,N_32005,N_39779);
and U48564 (N_48564,N_38732,N_31641);
nor U48565 (N_48565,N_36076,N_36950);
or U48566 (N_48566,N_30507,N_37346);
nor U48567 (N_48567,N_30834,N_37118);
nor U48568 (N_48568,N_33037,N_38629);
or U48569 (N_48569,N_37985,N_38780);
nand U48570 (N_48570,N_33602,N_34951);
or U48571 (N_48571,N_36351,N_35480);
nor U48572 (N_48572,N_35262,N_38239);
and U48573 (N_48573,N_30597,N_36870);
and U48574 (N_48574,N_33842,N_30115);
and U48575 (N_48575,N_33390,N_38643);
nor U48576 (N_48576,N_34014,N_32552);
and U48577 (N_48577,N_36859,N_30697);
and U48578 (N_48578,N_30831,N_32404);
and U48579 (N_48579,N_35600,N_37875);
xor U48580 (N_48580,N_39076,N_37569);
nand U48581 (N_48581,N_38344,N_39300);
or U48582 (N_48582,N_39384,N_35453);
or U48583 (N_48583,N_34769,N_33107);
nor U48584 (N_48584,N_38705,N_36710);
or U48585 (N_48585,N_33620,N_39664);
or U48586 (N_48586,N_38199,N_31388);
nor U48587 (N_48587,N_38837,N_39545);
xor U48588 (N_48588,N_34706,N_31629);
nand U48589 (N_48589,N_31769,N_35278);
or U48590 (N_48590,N_31032,N_34237);
nor U48591 (N_48591,N_30433,N_31662);
and U48592 (N_48592,N_34141,N_36235);
or U48593 (N_48593,N_39598,N_30253);
or U48594 (N_48594,N_35466,N_33199);
xnor U48595 (N_48595,N_34592,N_37578);
and U48596 (N_48596,N_33263,N_35984);
and U48597 (N_48597,N_30524,N_31977);
or U48598 (N_48598,N_39083,N_33954);
nor U48599 (N_48599,N_32331,N_32597);
nand U48600 (N_48600,N_33401,N_39175);
and U48601 (N_48601,N_34965,N_30251);
nor U48602 (N_48602,N_31571,N_31583);
and U48603 (N_48603,N_35281,N_30912);
nor U48604 (N_48604,N_37879,N_32819);
and U48605 (N_48605,N_32538,N_33574);
or U48606 (N_48606,N_35255,N_31678);
xnor U48607 (N_48607,N_35357,N_39041);
xor U48608 (N_48608,N_34118,N_34029);
and U48609 (N_48609,N_31907,N_32024);
nor U48610 (N_48610,N_32930,N_36534);
nor U48611 (N_48611,N_31742,N_33479);
nor U48612 (N_48612,N_33534,N_30624);
nand U48613 (N_48613,N_34989,N_31902);
nand U48614 (N_48614,N_34242,N_38395);
nor U48615 (N_48615,N_38013,N_36906);
nor U48616 (N_48616,N_37281,N_36147);
nand U48617 (N_48617,N_33652,N_30271);
and U48618 (N_48618,N_38983,N_32207);
nand U48619 (N_48619,N_37536,N_37618);
nand U48620 (N_48620,N_37263,N_39685);
nor U48621 (N_48621,N_37138,N_31019);
or U48622 (N_48622,N_30253,N_39678);
and U48623 (N_48623,N_36093,N_32734);
nor U48624 (N_48624,N_30927,N_39119);
nor U48625 (N_48625,N_39451,N_36194);
nand U48626 (N_48626,N_39437,N_35828);
and U48627 (N_48627,N_37387,N_38361);
nand U48628 (N_48628,N_38418,N_37410);
or U48629 (N_48629,N_30119,N_39825);
xnor U48630 (N_48630,N_35138,N_34062);
xor U48631 (N_48631,N_37927,N_33370);
nor U48632 (N_48632,N_33065,N_39135);
nand U48633 (N_48633,N_34630,N_39389);
xor U48634 (N_48634,N_33725,N_30294);
nand U48635 (N_48635,N_33245,N_37877);
nand U48636 (N_48636,N_37200,N_30779);
or U48637 (N_48637,N_38337,N_36331);
or U48638 (N_48638,N_38906,N_39521);
nand U48639 (N_48639,N_34471,N_39343);
xor U48640 (N_48640,N_33396,N_34416);
xor U48641 (N_48641,N_34987,N_35404);
or U48642 (N_48642,N_39163,N_34549);
and U48643 (N_48643,N_39109,N_34756);
nor U48644 (N_48644,N_31738,N_38613);
or U48645 (N_48645,N_33618,N_37891);
or U48646 (N_48646,N_38460,N_35463);
nand U48647 (N_48647,N_35810,N_31003);
nor U48648 (N_48648,N_37901,N_34986);
nand U48649 (N_48649,N_35206,N_39280);
nand U48650 (N_48650,N_34424,N_31342);
nor U48651 (N_48651,N_33533,N_36325);
nand U48652 (N_48652,N_38729,N_34645);
and U48653 (N_48653,N_32710,N_39073);
nand U48654 (N_48654,N_38113,N_30434);
nor U48655 (N_48655,N_38142,N_34640);
nand U48656 (N_48656,N_31089,N_32067);
nand U48657 (N_48657,N_37280,N_32311);
nor U48658 (N_48658,N_32689,N_33620);
or U48659 (N_48659,N_39016,N_36437);
nand U48660 (N_48660,N_35986,N_34414);
nand U48661 (N_48661,N_35241,N_35088);
and U48662 (N_48662,N_32302,N_30798);
nor U48663 (N_48663,N_34593,N_37567);
or U48664 (N_48664,N_39036,N_35650);
or U48665 (N_48665,N_32417,N_30909);
nand U48666 (N_48666,N_32441,N_36051);
nand U48667 (N_48667,N_35444,N_30601);
or U48668 (N_48668,N_33399,N_30821);
nand U48669 (N_48669,N_31567,N_38397);
or U48670 (N_48670,N_30793,N_38208);
nand U48671 (N_48671,N_36775,N_31003);
nor U48672 (N_48672,N_38591,N_33875);
and U48673 (N_48673,N_39091,N_38411);
or U48674 (N_48674,N_34583,N_39682);
nor U48675 (N_48675,N_32112,N_32907);
nand U48676 (N_48676,N_36892,N_39871);
nor U48677 (N_48677,N_37177,N_37164);
or U48678 (N_48678,N_38476,N_32099);
nor U48679 (N_48679,N_33204,N_34961);
nand U48680 (N_48680,N_38241,N_32527);
nand U48681 (N_48681,N_37456,N_34718);
or U48682 (N_48682,N_34061,N_39398);
and U48683 (N_48683,N_35139,N_36448);
nand U48684 (N_48684,N_37725,N_32478);
nor U48685 (N_48685,N_30411,N_38738);
and U48686 (N_48686,N_33538,N_35353);
nand U48687 (N_48687,N_33760,N_31659);
nand U48688 (N_48688,N_39956,N_30383);
and U48689 (N_48689,N_36562,N_33107);
and U48690 (N_48690,N_34503,N_32270);
and U48691 (N_48691,N_34318,N_37656);
nor U48692 (N_48692,N_39848,N_36705);
or U48693 (N_48693,N_33420,N_38019);
or U48694 (N_48694,N_33010,N_34036);
xor U48695 (N_48695,N_35609,N_30243);
and U48696 (N_48696,N_34959,N_32375);
and U48697 (N_48697,N_33905,N_35615);
nor U48698 (N_48698,N_36039,N_36343);
xnor U48699 (N_48699,N_38152,N_33197);
and U48700 (N_48700,N_32904,N_35542);
and U48701 (N_48701,N_39841,N_35603);
and U48702 (N_48702,N_34635,N_33570);
or U48703 (N_48703,N_34085,N_36675);
or U48704 (N_48704,N_31308,N_35859);
and U48705 (N_48705,N_30619,N_38231);
nor U48706 (N_48706,N_35327,N_30334);
nor U48707 (N_48707,N_34233,N_39346);
and U48708 (N_48708,N_32139,N_37154);
nor U48709 (N_48709,N_35866,N_31604);
xor U48710 (N_48710,N_32396,N_39790);
and U48711 (N_48711,N_35851,N_38646);
nand U48712 (N_48712,N_39850,N_39332);
xnor U48713 (N_48713,N_35017,N_32293);
xor U48714 (N_48714,N_37790,N_33911);
xnor U48715 (N_48715,N_33048,N_38785);
nor U48716 (N_48716,N_32757,N_39875);
xnor U48717 (N_48717,N_39367,N_32615);
and U48718 (N_48718,N_34383,N_32763);
nor U48719 (N_48719,N_31970,N_30809);
or U48720 (N_48720,N_37960,N_35528);
and U48721 (N_48721,N_38927,N_37624);
or U48722 (N_48722,N_35818,N_36610);
nor U48723 (N_48723,N_35304,N_35324);
nor U48724 (N_48724,N_37129,N_34785);
nor U48725 (N_48725,N_31171,N_39052);
nor U48726 (N_48726,N_35684,N_38727);
nor U48727 (N_48727,N_34143,N_37844);
nor U48728 (N_48728,N_30920,N_33858);
nor U48729 (N_48729,N_33156,N_34811);
nand U48730 (N_48730,N_38381,N_32565);
nand U48731 (N_48731,N_34653,N_39752);
and U48732 (N_48732,N_38876,N_37697);
or U48733 (N_48733,N_38752,N_32713);
and U48734 (N_48734,N_30327,N_39931);
xor U48735 (N_48735,N_33450,N_37146);
and U48736 (N_48736,N_31129,N_32658);
or U48737 (N_48737,N_36663,N_35859);
or U48738 (N_48738,N_37962,N_39342);
xor U48739 (N_48739,N_39867,N_37740);
or U48740 (N_48740,N_39240,N_33836);
and U48741 (N_48741,N_38716,N_33992);
or U48742 (N_48742,N_34033,N_38818);
or U48743 (N_48743,N_30136,N_33192);
and U48744 (N_48744,N_36193,N_31464);
nor U48745 (N_48745,N_32039,N_34695);
nor U48746 (N_48746,N_31490,N_32293);
xnor U48747 (N_48747,N_33730,N_36607);
nor U48748 (N_48748,N_30336,N_31765);
or U48749 (N_48749,N_34139,N_38799);
and U48750 (N_48750,N_35101,N_38984);
and U48751 (N_48751,N_31267,N_32882);
nor U48752 (N_48752,N_33039,N_39878);
nand U48753 (N_48753,N_36562,N_31412);
or U48754 (N_48754,N_38083,N_37526);
or U48755 (N_48755,N_37933,N_39408);
and U48756 (N_48756,N_39966,N_39862);
nand U48757 (N_48757,N_39546,N_33657);
nor U48758 (N_48758,N_33818,N_39690);
nor U48759 (N_48759,N_34631,N_37649);
and U48760 (N_48760,N_38935,N_38973);
nand U48761 (N_48761,N_39816,N_39318);
nand U48762 (N_48762,N_31308,N_32658);
and U48763 (N_48763,N_34919,N_30533);
and U48764 (N_48764,N_39295,N_39858);
or U48765 (N_48765,N_38152,N_38265);
or U48766 (N_48766,N_36118,N_38017);
nand U48767 (N_48767,N_30529,N_33495);
or U48768 (N_48768,N_34073,N_34228);
nand U48769 (N_48769,N_33892,N_39641);
nand U48770 (N_48770,N_38746,N_32879);
nand U48771 (N_48771,N_39122,N_33173);
and U48772 (N_48772,N_37204,N_39085);
nor U48773 (N_48773,N_38183,N_34277);
nand U48774 (N_48774,N_38447,N_35736);
or U48775 (N_48775,N_32607,N_31301);
nand U48776 (N_48776,N_33688,N_32036);
and U48777 (N_48777,N_38764,N_32415);
nor U48778 (N_48778,N_38420,N_31151);
nor U48779 (N_48779,N_37057,N_37244);
or U48780 (N_48780,N_30602,N_32892);
and U48781 (N_48781,N_32848,N_30468);
nand U48782 (N_48782,N_35885,N_33943);
or U48783 (N_48783,N_33982,N_36687);
nand U48784 (N_48784,N_38063,N_34088);
and U48785 (N_48785,N_32792,N_31254);
nor U48786 (N_48786,N_38795,N_31943);
and U48787 (N_48787,N_31942,N_33827);
nand U48788 (N_48788,N_39125,N_35816);
or U48789 (N_48789,N_36072,N_35132);
or U48790 (N_48790,N_36494,N_35606);
nor U48791 (N_48791,N_31170,N_37902);
nand U48792 (N_48792,N_36068,N_32858);
and U48793 (N_48793,N_37546,N_32139);
nand U48794 (N_48794,N_33352,N_33041);
or U48795 (N_48795,N_34931,N_35808);
nand U48796 (N_48796,N_37190,N_37487);
xnor U48797 (N_48797,N_36117,N_39486);
or U48798 (N_48798,N_39257,N_37811);
xor U48799 (N_48799,N_34633,N_37491);
nor U48800 (N_48800,N_37019,N_30278);
nor U48801 (N_48801,N_36932,N_30510);
nand U48802 (N_48802,N_36047,N_38697);
xor U48803 (N_48803,N_33108,N_36142);
and U48804 (N_48804,N_34890,N_37213);
nand U48805 (N_48805,N_32053,N_39779);
nor U48806 (N_48806,N_39291,N_32318);
nor U48807 (N_48807,N_33677,N_32884);
or U48808 (N_48808,N_38136,N_32324);
nor U48809 (N_48809,N_39779,N_38086);
xnor U48810 (N_48810,N_38548,N_38024);
nor U48811 (N_48811,N_35740,N_32151);
or U48812 (N_48812,N_32392,N_35533);
or U48813 (N_48813,N_37708,N_31233);
nand U48814 (N_48814,N_38024,N_37118);
nor U48815 (N_48815,N_38087,N_39802);
or U48816 (N_48816,N_39452,N_30170);
nand U48817 (N_48817,N_38935,N_30458);
nor U48818 (N_48818,N_31118,N_31355);
nor U48819 (N_48819,N_31643,N_31839);
nor U48820 (N_48820,N_35064,N_32478);
nor U48821 (N_48821,N_39791,N_37425);
and U48822 (N_48822,N_31201,N_32506);
nand U48823 (N_48823,N_35206,N_35863);
nor U48824 (N_48824,N_33222,N_36380);
xor U48825 (N_48825,N_39625,N_32279);
nor U48826 (N_48826,N_32987,N_30437);
nor U48827 (N_48827,N_36513,N_36877);
nand U48828 (N_48828,N_32724,N_30171);
and U48829 (N_48829,N_35033,N_31584);
and U48830 (N_48830,N_38651,N_32614);
nor U48831 (N_48831,N_32102,N_33759);
nand U48832 (N_48832,N_39326,N_31429);
nand U48833 (N_48833,N_31197,N_33409);
and U48834 (N_48834,N_39312,N_31847);
xnor U48835 (N_48835,N_34302,N_36689);
nand U48836 (N_48836,N_35971,N_37072);
nor U48837 (N_48837,N_39233,N_37602);
nand U48838 (N_48838,N_34723,N_30623);
nand U48839 (N_48839,N_34243,N_35416);
nor U48840 (N_48840,N_35032,N_30636);
or U48841 (N_48841,N_31140,N_38607);
nand U48842 (N_48842,N_35233,N_31816);
and U48843 (N_48843,N_35431,N_37881);
xor U48844 (N_48844,N_30271,N_39654);
nor U48845 (N_48845,N_34338,N_33658);
and U48846 (N_48846,N_37048,N_37514);
xnor U48847 (N_48847,N_31863,N_32124);
and U48848 (N_48848,N_31575,N_38759);
or U48849 (N_48849,N_37163,N_32636);
or U48850 (N_48850,N_36173,N_39111);
nand U48851 (N_48851,N_37410,N_37270);
nand U48852 (N_48852,N_39323,N_35714);
nand U48853 (N_48853,N_35499,N_33228);
and U48854 (N_48854,N_32978,N_34768);
and U48855 (N_48855,N_35805,N_35281);
nand U48856 (N_48856,N_31905,N_32520);
nor U48857 (N_48857,N_39088,N_30412);
or U48858 (N_48858,N_39808,N_33667);
or U48859 (N_48859,N_32413,N_33874);
nand U48860 (N_48860,N_35159,N_38695);
nor U48861 (N_48861,N_39248,N_38341);
xor U48862 (N_48862,N_35572,N_30425);
or U48863 (N_48863,N_33765,N_35443);
and U48864 (N_48864,N_34717,N_31184);
nand U48865 (N_48865,N_37995,N_32067);
or U48866 (N_48866,N_36050,N_38599);
or U48867 (N_48867,N_38868,N_39946);
or U48868 (N_48868,N_39945,N_36462);
and U48869 (N_48869,N_32054,N_38462);
or U48870 (N_48870,N_39432,N_32497);
nor U48871 (N_48871,N_35217,N_39434);
or U48872 (N_48872,N_30602,N_39135);
xor U48873 (N_48873,N_30908,N_39954);
nand U48874 (N_48874,N_32572,N_30201);
nor U48875 (N_48875,N_31521,N_36607);
or U48876 (N_48876,N_39106,N_33234);
nor U48877 (N_48877,N_38892,N_37584);
nand U48878 (N_48878,N_30772,N_31139);
and U48879 (N_48879,N_36343,N_39180);
xor U48880 (N_48880,N_32146,N_30978);
or U48881 (N_48881,N_33410,N_34985);
and U48882 (N_48882,N_32102,N_32048);
or U48883 (N_48883,N_39364,N_31996);
nor U48884 (N_48884,N_31243,N_32523);
and U48885 (N_48885,N_39809,N_38225);
nor U48886 (N_48886,N_32134,N_38698);
and U48887 (N_48887,N_33295,N_38278);
nor U48888 (N_48888,N_30052,N_36056);
nor U48889 (N_48889,N_39860,N_38884);
nor U48890 (N_48890,N_34810,N_37476);
or U48891 (N_48891,N_33179,N_31764);
nand U48892 (N_48892,N_39639,N_37133);
nor U48893 (N_48893,N_35852,N_37332);
nand U48894 (N_48894,N_36221,N_30787);
or U48895 (N_48895,N_38176,N_32808);
and U48896 (N_48896,N_32991,N_32068);
or U48897 (N_48897,N_37458,N_31109);
nor U48898 (N_48898,N_39536,N_36865);
and U48899 (N_48899,N_33297,N_31870);
and U48900 (N_48900,N_37480,N_30627);
nor U48901 (N_48901,N_31899,N_39330);
nor U48902 (N_48902,N_33425,N_38281);
nor U48903 (N_48903,N_39816,N_31747);
nand U48904 (N_48904,N_34136,N_38392);
or U48905 (N_48905,N_35751,N_30748);
or U48906 (N_48906,N_34752,N_30835);
nor U48907 (N_48907,N_30979,N_39903);
or U48908 (N_48908,N_32612,N_30880);
xor U48909 (N_48909,N_34044,N_37441);
nand U48910 (N_48910,N_35860,N_33426);
xnor U48911 (N_48911,N_32246,N_39905);
and U48912 (N_48912,N_37903,N_36677);
nand U48913 (N_48913,N_34731,N_37560);
nor U48914 (N_48914,N_39192,N_39652);
and U48915 (N_48915,N_35637,N_30441);
xor U48916 (N_48916,N_34442,N_30752);
and U48917 (N_48917,N_32170,N_34157);
or U48918 (N_48918,N_36853,N_37683);
or U48919 (N_48919,N_39298,N_31317);
and U48920 (N_48920,N_34767,N_32941);
nor U48921 (N_48921,N_34490,N_39256);
nor U48922 (N_48922,N_32735,N_36738);
and U48923 (N_48923,N_33757,N_39399);
nor U48924 (N_48924,N_37378,N_39206);
nor U48925 (N_48925,N_35448,N_35094);
nand U48926 (N_48926,N_38357,N_37561);
nor U48927 (N_48927,N_30947,N_38002);
xnor U48928 (N_48928,N_38436,N_38402);
nor U48929 (N_48929,N_31742,N_36334);
or U48930 (N_48930,N_33820,N_39040);
nor U48931 (N_48931,N_36870,N_34374);
or U48932 (N_48932,N_35763,N_31138);
and U48933 (N_48933,N_32878,N_37799);
or U48934 (N_48934,N_32302,N_33295);
or U48935 (N_48935,N_38307,N_33561);
and U48936 (N_48936,N_37172,N_32185);
or U48937 (N_48937,N_32016,N_31982);
or U48938 (N_48938,N_31124,N_33768);
and U48939 (N_48939,N_31919,N_35491);
and U48940 (N_48940,N_38585,N_36737);
or U48941 (N_48941,N_37615,N_30054);
and U48942 (N_48942,N_37523,N_33072);
nand U48943 (N_48943,N_31052,N_35172);
nor U48944 (N_48944,N_34899,N_30171);
and U48945 (N_48945,N_37480,N_39440);
or U48946 (N_48946,N_38944,N_34216);
nor U48947 (N_48947,N_37888,N_39562);
xnor U48948 (N_48948,N_34156,N_32868);
or U48949 (N_48949,N_30398,N_36921);
nor U48950 (N_48950,N_33767,N_31203);
and U48951 (N_48951,N_39236,N_33890);
or U48952 (N_48952,N_30140,N_39716);
and U48953 (N_48953,N_38813,N_34192);
xnor U48954 (N_48954,N_32978,N_39072);
or U48955 (N_48955,N_34553,N_30807);
nor U48956 (N_48956,N_37234,N_38401);
nor U48957 (N_48957,N_33673,N_39264);
nor U48958 (N_48958,N_34862,N_30365);
and U48959 (N_48959,N_34412,N_31599);
or U48960 (N_48960,N_39002,N_34443);
or U48961 (N_48961,N_31331,N_39022);
and U48962 (N_48962,N_34414,N_38601);
or U48963 (N_48963,N_36046,N_36730);
nor U48964 (N_48964,N_37092,N_36413);
or U48965 (N_48965,N_37937,N_36765);
nor U48966 (N_48966,N_32154,N_37306);
nand U48967 (N_48967,N_34083,N_35462);
and U48968 (N_48968,N_31792,N_32716);
and U48969 (N_48969,N_30447,N_38114);
nor U48970 (N_48970,N_36516,N_39935);
nor U48971 (N_48971,N_34310,N_39709);
nor U48972 (N_48972,N_39291,N_34709);
and U48973 (N_48973,N_30808,N_35191);
nor U48974 (N_48974,N_35221,N_34565);
xnor U48975 (N_48975,N_36850,N_38185);
or U48976 (N_48976,N_30668,N_31628);
nor U48977 (N_48977,N_37454,N_32148);
and U48978 (N_48978,N_32829,N_38726);
nand U48979 (N_48979,N_36068,N_36434);
nor U48980 (N_48980,N_30459,N_32214);
nand U48981 (N_48981,N_38432,N_36638);
nor U48982 (N_48982,N_38348,N_33065);
or U48983 (N_48983,N_30430,N_36739);
or U48984 (N_48984,N_38513,N_34080);
or U48985 (N_48985,N_36988,N_37745);
nor U48986 (N_48986,N_34175,N_39932);
and U48987 (N_48987,N_39669,N_32890);
or U48988 (N_48988,N_35637,N_30049);
nand U48989 (N_48989,N_39454,N_38431);
nand U48990 (N_48990,N_34041,N_32357);
and U48991 (N_48991,N_30705,N_35308);
xor U48992 (N_48992,N_36183,N_38973);
or U48993 (N_48993,N_30969,N_37799);
nor U48994 (N_48994,N_36887,N_35460);
nand U48995 (N_48995,N_32087,N_39897);
nor U48996 (N_48996,N_31339,N_34024);
and U48997 (N_48997,N_35556,N_35645);
or U48998 (N_48998,N_38417,N_35518);
xnor U48999 (N_48999,N_39261,N_34288);
xnor U49000 (N_49000,N_30822,N_39744);
or U49001 (N_49001,N_38951,N_34405);
and U49002 (N_49002,N_31880,N_34482);
nor U49003 (N_49003,N_34608,N_34231);
nand U49004 (N_49004,N_31435,N_34911);
and U49005 (N_49005,N_33707,N_30293);
and U49006 (N_49006,N_37533,N_39372);
nand U49007 (N_49007,N_33528,N_32505);
nor U49008 (N_49008,N_38977,N_31866);
and U49009 (N_49009,N_38135,N_39154);
nor U49010 (N_49010,N_33848,N_37006);
and U49011 (N_49011,N_30820,N_31471);
xor U49012 (N_49012,N_30379,N_34693);
or U49013 (N_49013,N_32786,N_38840);
nand U49014 (N_49014,N_32997,N_30239);
xor U49015 (N_49015,N_30607,N_32110);
nor U49016 (N_49016,N_38281,N_32876);
nor U49017 (N_49017,N_38098,N_34575);
and U49018 (N_49018,N_30051,N_30655);
or U49019 (N_49019,N_33811,N_32410);
and U49020 (N_49020,N_37285,N_31706);
nor U49021 (N_49021,N_30200,N_30896);
nand U49022 (N_49022,N_30935,N_37233);
and U49023 (N_49023,N_39051,N_31242);
xor U49024 (N_49024,N_38976,N_37600);
nand U49025 (N_49025,N_32257,N_38404);
nor U49026 (N_49026,N_33382,N_35095);
nand U49027 (N_49027,N_30633,N_35928);
nand U49028 (N_49028,N_33239,N_34752);
or U49029 (N_49029,N_38752,N_35458);
and U49030 (N_49030,N_38710,N_36829);
or U49031 (N_49031,N_37779,N_38557);
and U49032 (N_49032,N_33315,N_35432);
nor U49033 (N_49033,N_33383,N_34441);
and U49034 (N_49034,N_36208,N_34361);
nand U49035 (N_49035,N_36596,N_37181);
and U49036 (N_49036,N_32488,N_39820);
nor U49037 (N_49037,N_31598,N_32756);
nand U49038 (N_49038,N_34601,N_31758);
or U49039 (N_49039,N_30404,N_37548);
xor U49040 (N_49040,N_32741,N_30661);
nand U49041 (N_49041,N_32906,N_31423);
and U49042 (N_49042,N_34150,N_32290);
xor U49043 (N_49043,N_32384,N_36952);
nor U49044 (N_49044,N_31340,N_33777);
xor U49045 (N_49045,N_33980,N_39448);
xnor U49046 (N_49046,N_32439,N_31679);
or U49047 (N_49047,N_34087,N_33496);
nand U49048 (N_49048,N_39767,N_33357);
and U49049 (N_49049,N_36827,N_33555);
xnor U49050 (N_49050,N_36997,N_30215);
nor U49051 (N_49051,N_39395,N_35195);
and U49052 (N_49052,N_33056,N_32545);
nor U49053 (N_49053,N_37747,N_35070);
and U49054 (N_49054,N_34318,N_31174);
nor U49055 (N_49055,N_37938,N_35105);
xor U49056 (N_49056,N_30895,N_30440);
and U49057 (N_49057,N_36792,N_34106);
and U49058 (N_49058,N_36621,N_37957);
or U49059 (N_49059,N_36906,N_36603);
nor U49060 (N_49060,N_35885,N_37635);
nand U49061 (N_49061,N_31578,N_34545);
nor U49062 (N_49062,N_33626,N_38391);
or U49063 (N_49063,N_33590,N_35735);
nor U49064 (N_49064,N_38351,N_37747);
nand U49065 (N_49065,N_33060,N_31350);
or U49066 (N_49066,N_32244,N_32441);
and U49067 (N_49067,N_34781,N_30064);
nand U49068 (N_49068,N_38533,N_33428);
nand U49069 (N_49069,N_35894,N_32876);
or U49070 (N_49070,N_34920,N_31713);
or U49071 (N_49071,N_37482,N_39956);
or U49072 (N_49072,N_31828,N_35645);
nor U49073 (N_49073,N_37553,N_37868);
xor U49074 (N_49074,N_37662,N_36838);
nor U49075 (N_49075,N_31725,N_32167);
or U49076 (N_49076,N_30193,N_30027);
and U49077 (N_49077,N_34623,N_34631);
nand U49078 (N_49078,N_37741,N_35092);
and U49079 (N_49079,N_39505,N_35809);
and U49080 (N_49080,N_39149,N_32346);
and U49081 (N_49081,N_34244,N_35053);
or U49082 (N_49082,N_31811,N_34694);
nor U49083 (N_49083,N_35044,N_36202);
and U49084 (N_49084,N_37408,N_32038);
xor U49085 (N_49085,N_33496,N_39600);
or U49086 (N_49086,N_34408,N_36502);
and U49087 (N_49087,N_36227,N_37884);
nor U49088 (N_49088,N_38328,N_36008);
nand U49089 (N_49089,N_32492,N_32504);
nor U49090 (N_49090,N_30180,N_32791);
or U49091 (N_49091,N_32481,N_30185);
and U49092 (N_49092,N_34012,N_31451);
xor U49093 (N_49093,N_35534,N_33633);
and U49094 (N_49094,N_31785,N_34188);
and U49095 (N_49095,N_35395,N_39756);
nor U49096 (N_49096,N_34932,N_30305);
xnor U49097 (N_49097,N_39719,N_34084);
nor U49098 (N_49098,N_38541,N_34098);
nor U49099 (N_49099,N_38688,N_39614);
nor U49100 (N_49100,N_39042,N_35985);
and U49101 (N_49101,N_32391,N_36781);
nand U49102 (N_49102,N_37820,N_35138);
and U49103 (N_49103,N_30061,N_37232);
and U49104 (N_49104,N_36229,N_34961);
nand U49105 (N_49105,N_30887,N_39476);
xor U49106 (N_49106,N_31603,N_37272);
xnor U49107 (N_49107,N_31794,N_37570);
nor U49108 (N_49108,N_35776,N_34615);
or U49109 (N_49109,N_38615,N_31056);
or U49110 (N_49110,N_31554,N_33136);
and U49111 (N_49111,N_38148,N_36997);
or U49112 (N_49112,N_30498,N_35077);
nor U49113 (N_49113,N_39912,N_32813);
nand U49114 (N_49114,N_39008,N_34135);
and U49115 (N_49115,N_35797,N_37727);
nand U49116 (N_49116,N_33221,N_36009);
or U49117 (N_49117,N_31448,N_34961);
and U49118 (N_49118,N_32663,N_30489);
xor U49119 (N_49119,N_34527,N_38594);
or U49120 (N_49120,N_34358,N_36196);
or U49121 (N_49121,N_36257,N_35774);
xnor U49122 (N_49122,N_30633,N_33641);
or U49123 (N_49123,N_30607,N_35500);
xnor U49124 (N_49124,N_39631,N_30266);
nor U49125 (N_49125,N_39255,N_34054);
xor U49126 (N_49126,N_34115,N_37021);
or U49127 (N_49127,N_31856,N_34928);
and U49128 (N_49128,N_33582,N_37144);
nor U49129 (N_49129,N_37023,N_34070);
and U49130 (N_49130,N_38218,N_35322);
nand U49131 (N_49131,N_30974,N_35602);
xnor U49132 (N_49132,N_35072,N_30049);
and U49133 (N_49133,N_37665,N_32300);
and U49134 (N_49134,N_33665,N_36659);
or U49135 (N_49135,N_37649,N_33591);
nand U49136 (N_49136,N_36883,N_35946);
xor U49137 (N_49137,N_32327,N_30453);
nand U49138 (N_49138,N_35194,N_30928);
nor U49139 (N_49139,N_30388,N_39050);
nor U49140 (N_49140,N_36836,N_38697);
nor U49141 (N_49141,N_37524,N_33016);
nand U49142 (N_49142,N_35372,N_34419);
or U49143 (N_49143,N_38477,N_39943);
xor U49144 (N_49144,N_36616,N_30980);
or U49145 (N_49145,N_39010,N_34798);
xor U49146 (N_49146,N_38681,N_32695);
nor U49147 (N_49147,N_34005,N_33773);
nor U49148 (N_49148,N_31180,N_35053);
or U49149 (N_49149,N_39657,N_38645);
nand U49150 (N_49150,N_34079,N_31146);
and U49151 (N_49151,N_35134,N_31683);
and U49152 (N_49152,N_31647,N_38646);
nor U49153 (N_49153,N_30003,N_33493);
and U49154 (N_49154,N_37178,N_39765);
nand U49155 (N_49155,N_36503,N_37654);
and U49156 (N_49156,N_35728,N_36905);
xor U49157 (N_49157,N_34565,N_37009);
and U49158 (N_49158,N_38555,N_37087);
or U49159 (N_49159,N_32222,N_38801);
or U49160 (N_49160,N_31361,N_33685);
nor U49161 (N_49161,N_35126,N_37147);
nand U49162 (N_49162,N_39561,N_38306);
nor U49163 (N_49163,N_39245,N_34747);
nor U49164 (N_49164,N_37240,N_34654);
or U49165 (N_49165,N_39690,N_36820);
nor U49166 (N_49166,N_34685,N_35056);
or U49167 (N_49167,N_36718,N_30098);
or U49168 (N_49168,N_36532,N_38820);
and U49169 (N_49169,N_35755,N_37902);
nor U49170 (N_49170,N_36473,N_30914);
nor U49171 (N_49171,N_39775,N_33163);
or U49172 (N_49172,N_37870,N_30603);
and U49173 (N_49173,N_37005,N_30453);
nor U49174 (N_49174,N_35090,N_39090);
nor U49175 (N_49175,N_33033,N_39298);
and U49176 (N_49176,N_35441,N_39046);
or U49177 (N_49177,N_30627,N_34065);
nand U49178 (N_49178,N_30043,N_32364);
nand U49179 (N_49179,N_35670,N_31672);
xnor U49180 (N_49180,N_32497,N_34925);
or U49181 (N_49181,N_36904,N_38682);
nand U49182 (N_49182,N_30218,N_38113);
and U49183 (N_49183,N_31286,N_38345);
xnor U49184 (N_49184,N_33221,N_32486);
or U49185 (N_49185,N_30631,N_38215);
nand U49186 (N_49186,N_37336,N_34862);
or U49187 (N_49187,N_31159,N_31748);
nor U49188 (N_49188,N_33715,N_37200);
xor U49189 (N_49189,N_31709,N_34777);
xnor U49190 (N_49190,N_37063,N_32612);
nor U49191 (N_49191,N_33652,N_31167);
or U49192 (N_49192,N_37602,N_36961);
and U49193 (N_49193,N_32309,N_30372);
or U49194 (N_49194,N_30731,N_33490);
or U49195 (N_49195,N_33690,N_37514);
or U49196 (N_49196,N_33396,N_31603);
xnor U49197 (N_49197,N_31611,N_31014);
nor U49198 (N_49198,N_38602,N_33009);
or U49199 (N_49199,N_34512,N_32270);
nor U49200 (N_49200,N_32355,N_37643);
nor U49201 (N_49201,N_34418,N_30870);
or U49202 (N_49202,N_35375,N_36728);
and U49203 (N_49203,N_35109,N_38612);
nand U49204 (N_49204,N_35506,N_33934);
or U49205 (N_49205,N_38580,N_35532);
xor U49206 (N_49206,N_33214,N_32039);
and U49207 (N_49207,N_39718,N_38850);
nor U49208 (N_49208,N_37422,N_38942);
nand U49209 (N_49209,N_33998,N_35211);
nand U49210 (N_49210,N_33466,N_39279);
nand U49211 (N_49211,N_37903,N_39029);
nand U49212 (N_49212,N_38411,N_36766);
or U49213 (N_49213,N_38148,N_37690);
nor U49214 (N_49214,N_36668,N_34899);
or U49215 (N_49215,N_39220,N_30712);
or U49216 (N_49216,N_39710,N_39401);
or U49217 (N_49217,N_35203,N_33188);
nor U49218 (N_49218,N_39865,N_34093);
nand U49219 (N_49219,N_34053,N_35987);
and U49220 (N_49220,N_38117,N_35416);
or U49221 (N_49221,N_30816,N_36358);
nand U49222 (N_49222,N_31810,N_39093);
nor U49223 (N_49223,N_34430,N_30210);
xnor U49224 (N_49224,N_37719,N_31372);
nor U49225 (N_49225,N_32450,N_38228);
nor U49226 (N_49226,N_39906,N_35508);
or U49227 (N_49227,N_34416,N_37068);
nand U49228 (N_49228,N_38760,N_38196);
xor U49229 (N_49229,N_34925,N_30423);
nor U49230 (N_49230,N_38085,N_35722);
and U49231 (N_49231,N_33218,N_36348);
nand U49232 (N_49232,N_34563,N_36709);
xnor U49233 (N_49233,N_34339,N_35820);
nor U49234 (N_49234,N_36457,N_37984);
xor U49235 (N_49235,N_33906,N_37539);
nor U49236 (N_49236,N_31464,N_37858);
or U49237 (N_49237,N_39162,N_37020);
or U49238 (N_49238,N_30305,N_37652);
nor U49239 (N_49239,N_38185,N_31873);
or U49240 (N_49240,N_35702,N_35020);
and U49241 (N_49241,N_33519,N_35494);
nor U49242 (N_49242,N_30972,N_37242);
nor U49243 (N_49243,N_37147,N_33730);
xnor U49244 (N_49244,N_31521,N_30270);
nor U49245 (N_49245,N_39107,N_35123);
nor U49246 (N_49246,N_32336,N_30241);
nor U49247 (N_49247,N_32188,N_31957);
nor U49248 (N_49248,N_35633,N_34460);
or U49249 (N_49249,N_30909,N_30602);
or U49250 (N_49250,N_34175,N_39880);
or U49251 (N_49251,N_39335,N_38046);
xor U49252 (N_49252,N_38816,N_37655);
nand U49253 (N_49253,N_30450,N_30842);
and U49254 (N_49254,N_35954,N_35352);
nor U49255 (N_49255,N_37687,N_38650);
nor U49256 (N_49256,N_32506,N_38912);
nor U49257 (N_49257,N_39348,N_33471);
and U49258 (N_49258,N_32946,N_32371);
or U49259 (N_49259,N_33377,N_39639);
xnor U49260 (N_49260,N_36716,N_32036);
nor U49261 (N_49261,N_30655,N_37049);
nand U49262 (N_49262,N_30798,N_34881);
and U49263 (N_49263,N_39741,N_32887);
and U49264 (N_49264,N_32851,N_33266);
nor U49265 (N_49265,N_32059,N_36079);
nand U49266 (N_49266,N_39328,N_34720);
nand U49267 (N_49267,N_38070,N_34431);
and U49268 (N_49268,N_37978,N_30348);
or U49269 (N_49269,N_37829,N_38133);
nand U49270 (N_49270,N_31978,N_37012);
nor U49271 (N_49271,N_39288,N_39856);
or U49272 (N_49272,N_30314,N_38641);
and U49273 (N_49273,N_36329,N_38553);
and U49274 (N_49274,N_38155,N_35391);
or U49275 (N_49275,N_34049,N_33354);
nor U49276 (N_49276,N_37806,N_31877);
and U49277 (N_49277,N_32322,N_30436);
or U49278 (N_49278,N_37852,N_31448);
xnor U49279 (N_49279,N_32444,N_30283);
nor U49280 (N_49280,N_38935,N_38906);
and U49281 (N_49281,N_36984,N_37977);
nor U49282 (N_49282,N_33804,N_33581);
nor U49283 (N_49283,N_35334,N_31620);
nor U49284 (N_49284,N_36582,N_33610);
or U49285 (N_49285,N_34050,N_35728);
nand U49286 (N_49286,N_38721,N_30221);
nor U49287 (N_49287,N_30554,N_34460);
nor U49288 (N_49288,N_36181,N_38094);
and U49289 (N_49289,N_34979,N_33309);
nand U49290 (N_49290,N_36986,N_38145);
nand U49291 (N_49291,N_35634,N_30140);
xor U49292 (N_49292,N_30170,N_33010);
nor U49293 (N_49293,N_36352,N_30123);
or U49294 (N_49294,N_35085,N_39701);
nor U49295 (N_49295,N_31053,N_37916);
nand U49296 (N_49296,N_38788,N_34062);
nand U49297 (N_49297,N_33991,N_39755);
and U49298 (N_49298,N_38819,N_39204);
xnor U49299 (N_49299,N_32980,N_31658);
or U49300 (N_49300,N_37904,N_37096);
nand U49301 (N_49301,N_30048,N_32543);
xnor U49302 (N_49302,N_30135,N_31335);
xnor U49303 (N_49303,N_38437,N_37620);
and U49304 (N_49304,N_32399,N_31143);
and U49305 (N_49305,N_39407,N_30915);
and U49306 (N_49306,N_36699,N_35500);
or U49307 (N_49307,N_33984,N_34405);
nor U49308 (N_49308,N_36133,N_35264);
or U49309 (N_49309,N_33661,N_36793);
or U49310 (N_49310,N_31531,N_39547);
and U49311 (N_49311,N_37442,N_30185);
or U49312 (N_49312,N_38460,N_34437);
nand U49313 (N_49313,N_37436,N_33946);
and U49314 (N_49314,N_31114,N_38805);
nor U49315 (N_49315,N_37781,N_33442);
and U49316 (N_49316,N_36194,N_39309);
or U49317 (N_49317,N_31437,N_34965);
and U49318 (N_49318,N_33341,N_30199);
nand U49319 (N_49319,N_36564,N_33702);
nand U49320 (N_49320,N_38321,N_35407);
nor U49321 (N_49321,N_32546,N_35536);
and U49322 (N_49322,N_30833,N_36308);
and U49323 (N_49323,N_33269,N_37381);
or U49324 (N_49324,N_36267,N_33524);
or U49325 (N_49325,N_35683,N_35002);
xor U49326 (N_49326,N_39029,N_36618);
nor U49327 (N_49327,N_31954,N_34172);
nand U49328 (N_49328,N_33566,N_36366);
and U49329 (N_49329,N_33441,N_33515);
or U49330 (N_49330,N_30925,N_35093);
or U49331 (N_49331,N_33971,N_38976);
and U49332 (N_49332,N_35694,N_34364);
and U49333 (N_49333,N_39846,N_35964);
and U49334 (N_49334,N_39537,N_34097);
nand U49335 (N_49335,N_34448,N_39966);
nand U49336 (N_49336,N_34108,N_38260);
or U49337 (N_49337,N_39857,N_35319);
and U49338 (N_49338,N_37179,N_35905);
or U49339 (N_49339,N_38896,N_36372);
and U49340 (N_49340,N_33723,N_38674);
xnor U49341 (N_49341,N_37925,N_30561);
and U49342 (N_49342,N_30507,N_37284);
or U49343 (N_49343,N_32883,N_32204);
xnor U49344 (N_49344,N_31140,N_32124);
nand U49345 (N_49345,N_35944,N_38188);
and U49346 (N_49346,N_38388,N_35664);
nor U49347 (N_49347,N_34472,N_35464);
nand U49348 (N_49348,N_32082,N_32132);
nand U49349 (N_49349,N_35609,N_33495);
or U49350 (N_49350,N_33012,N_30687);
or U49351 (N_49351,N_39582,N_35967);
or U49352 (N_49352,N_33276,N_35625);
or U49353 (N_49353,N_31823,N_38882);
nor U49354 (N_49354,N_39351,N_37644);
nand U49355 (N_49355,N_39478,N_38839);
nand U49356 (N_49356,N_34270,N_35915);
nor U49357 (N_49357,N_31941,N_35222);
nand U49358 (N_49358,N_33540,N_39334);
nand U49359 (N_49359,N_38791,N_37413);
or U49360 (N_49360,N_35766,N_30856);
xor U49361 (N_49361,N_32024,N_39148);
and U49362 (N_49362,N_35959,N_36763);
or U49363 (N_49363,N_38806,N_34313);
and U49364 (N_49364,N_30529,N_36614);
or U49365 (N_49365,N_32999,N_34576);
nor U49366 (N_49366,N_34888,N_35317);
nor U49367 (N_49367,N_30702,N_36685);
nand U49368 (N_49368,N_32054,N_31690);
and U49369 (N_49369,N_36026,N_38052);
nand U49370 (N_49370,N_37051,N_39511);
and U49371 (N_49371,N_33342,N_30208);
xor U49372 (N_49372,N_37100,N_30898);
nand U49373 (N_49373,N_32523,N_36185);
and U49374 (N_49374,N_35520,N_39675);
and U49375 (N_49375,N_36965,N_38842);
nand U49376 (N_49376,N_35841,N_39833);
nor U49377 (N_49377,N_34106,N_35994);
or U49378 (N_49378,N_38550,N_31150);
nand U49379 (N_49379,N_38315,N_38492);
nand U49380 (N_49380,N_37909,N_38661);
xor U49381 (N_49381,N_30522,N_32119);
nor U49382 (N_49382,N_39411,N_33241);
or U49383 (N_49383,N_32050,N_38101);
and U49384 (N_49384,N_36431,N_37467);
or U49385 (N_49385,N_38140,N_38490);
or U49386 (N_49386,N_38988,N_33128);
nor U49387 (N_49387,N_35611,N_38738);
and U49388 (N_49388,N_37006,N_39574);
xor U49389 (N_49389,N_32642,N_32344);
nor U49390 (N_49390,N_38390,N_38905);
and U49391 (N_49391,N_30014,N_36559);
nand U49392 (N_49392,N_32489,N_34795);
or U49393 (N_49393,N_32686,N_32013);
or U49394 (N_49394,N_32447,N_30177);
nand U49395 (N_49395,N_38248,N_39510);
nand U49396 (N_49396,N_35116,N_32430);
or U49397 (N_49397,N_34834,N_37923);
and U49398 (N_49398,N_32250,N_35668);
and U49399 (N_49399,N_34276,N_31288);
xor U49400 (N_49400,N_39521,N_36066);
nor U49401 (N_49401,N_37738,N_32197);
or U49402 (N_49402,N_35102,N_37823);
or U49403 (N_49403,N_33452,N_34506);
or U49404 (N_49404,N_33624,N_36941);
or U49405 (N_49405,N_34189,N_33327);
nor U49406 (N_49406,N_34637,N_37126);
nand U49407 (N_49407,N_30790,N_31183);
nor U49408 (N_49408,N_31855,N_31645);
and U49409 (N_49409,N_30870,N_39056);
xor U49410 (N_49410,N_33780,N_37499);
or U49411 (N_49411,N_32044,N_32143);
nand U49412 (N_49412,N_34240,N_36440);
nor U49413 (N_49413,N_38022,N_34658);
and U49414 (N_49414,N_33626,N_31764);
and U49415 (N_49415,N_31555,N_39189);
or U49416 (N_49416,N_35468,N_39073);
and U49417 (N_49417,N_36940,N_37308);
or U49418 (N_49418,N_30486,N_35404);
and U49419 (N_49419,N_33667,N_32384);
nand U49420 (N_49420,N_37479,N_39148);
nand U49421 (N_49421,N_38729,N_39677);
and U49422 (N_49422,N_39970,N_36087);
or U49423 (N_49423,N_39974,N_37612);
nand U49424 (N_49424,N_34536,N_33346);
or U49425 (N_49425,N_33494,N_32694);
nor U49426 (N_49426,N_39543,N_38784);
and U49427 (N_49427,N_36296,N_35736);
nor U49428 (N_49428,N_37352,N_33273);
and U49429 (N_49429,N_34870,N_39232);
or U49430 (N_49430,N_30250,N_38162);
and U49431 (N_49431,N_32628,N_38270);
nand U49432 (N_49432,N_34447,N_30496);
or U49433 (N_49433,N_37470,N_37540);
or U49434 (N_49434,N_33846,N_33283);
nor U49435 (N_49435,N_35422,N_32177);
nor U49436 (N_49436,N_33081,N_33277);
nand U49437 (N_49437,N_34298,N_34736);
and U49438 (N_49438,N_32152,N_37163);
or U49439 (N_49439,N_33364,N_30143);
or U49440 (N_49440,N_35137,N_30820);
nor U49441 (N_49441,N_30310,N_30648);
nor U49442 (N_49442,N_39829,N_37831);
and U49443 (N_49443,N_35466,N_31764);
nand U49444 (N_49444,N_38755,N_32201);
nor U49445 (N_49445,N_30542,N_33573);
or U49446 (N_49446,N_35019,N_38987);
xor U49447 (N_49447,N_39495,N_36651);
nor U49448 (N_49448,N_39181,N_33202);
nand U49449 (N_49449,N_36715,N_32611);
and U49450 (N_49450,N_38236,N_38529);
nand U49451 (N_49451,N_32056,N_39811);
xor U49452 (N_49452,N_30167,N_32101);
and U49453 (N_49453,N_38620,N_39439);
or U49454 (N_49454,N_39471,N_34618);
and U49455 (N_49455,N_37334,N_38221);
nand U49456 (N_49456,N_38113,N_30116);
xor U49457 (N_49457,N_31046,N_38665);
or U49458 (N_49458,N_39690,N_33862);
and U49459 (N_49459,N_32599,N_31979);
or U49460 (N_49460,N_33658,N_37115);
nand U49461 (N_49461,N_38444,N_33968);
and U49462 (N_49462,N_31178,N_38945);
and U49463 (N_49463,N_35896,N_31217);
nor U49464 (N_49464,N_39946,N_30377);
and U49465 (N_49465,N_35449,N_33453);
nor U49466 (N_49466,N_36946,N_34498);
and U49467 (N_49467,N_39435,N_31149);
or U49468 (N_49468,N_35851,N_38725);
nor U49469 (N_49469,N_30958,N_35970);
and U49470 (N_49470,N_33261,N_31833);
or U49471 (N_49471,N_33073,N_31804);
or U49472 (N_49472,N_30221,N_30166);
nor U49473 (N_49473,N_32367,N_34048);
nand U49474 (N_49474,N_35826,N_34096);
nand U49475 (N_49475,N_35110,N_33019);
or U49476 (N_49476,N_32863,N_34944);
and U49477 (N_49477,N_31934,N_31020);
nor U49478 (N_49478,N_38907,N_30500);
or U49479 (N_49479,N_38259,N_36761);
xnor U49480 (N_49480,N_36914,N_39392);
or U49481 (N_49481,N_30643,N_31374);
nand U49482 (N_49482,N_31303,N_39634);
nand U49483 (N_49483,N_31017,N_34591);
and U49484 (N_49484,N_32878,N_38587);
and U49485 (N_49485,N_36420,N_38843);
or U49486 (N_49486,N_35838,N_37718);
or U49487 (N_49487,N_31246,N_31790);
nand U49488 (N_49488,N_32751,N_35981);
nand U49489 (N_49489,N_32978,N_39115);
or U49490 (N_49490,N_31889,N_34335);
nand U49491 (N_49491,N_36706,N_33249);
nand U49492 (N_49492,N_33605,N_35274);
nor U49493 (N_49493,N_38188,N_39424);
nor U49494 (N_49494,N_38622,N_31406);
or U49495 (N_49495,N_32370,N_31496);
or U49496 (N_49496,N_34871,N_36694);
xor U49497 (N_49497,N_39489,N_37524);
xor U49498 (N_49498,N_37539,N_36633);
and U49499 (N_49499,N_34480,N_32921);
nor U49500 (N_49500,N_36243,N_38830);
or U49501 (N_49501,N_38913,N_32898);
nor U49502 (N_49502,N_33808,N_30122);
xor U49503 (N_49503,N_35817,N_33729);
and U49504 (N_49504,N_31840,N_35890);
and U49505 (N_49505,N_33956,N_35326);
nand U49506 (N_49506,N_39708,N_33515);
nor U49507 (N_49507,N_39536,N_32373);
nor U49508 (N_49508,N_38120,N_37802);
xnor U49509 (N_49509,N_30179,N_32360);
xnor U49510 (N_49510,N_38553,N_30704);
nor U49511 (N_49511,N_36695,N_34647);
nand U49512 (N_49512,N_32931,N_39733);
or U49513 (N_49513,N_30953,N_30399);
and U49514 (N_49514,N_32933,N_33250);
and U49515 (N_49515,N_33992,N_31165);
and U49516 (N_49516,N_31469,N_36027);
nand U49517 (N_49517,N_37849,N_32970);
and U49518 (N_49518,N_34541,N_34201);
nand U49519 (N_49519,N_37468,N_35496);
or U49520 (N_49520,N_31076,N_39473);
xnor U49521 (N_49521,N_31556,N_37007);
or U49522 (N_49522,N_31975,N_30979);
nor U49523 (N_49523,N_32263,N_30443);
or U49524 (N_49524,N_37486,N_30968);
nor U49525 (N_49525,N_37975,N_39630);
nor U49526 (N_49526,N_30596,N_31333);
nor U49527 (N_49527,N_39571,N_36277);
nor U49528 (N_49528,N_36978,N_39856);
or U49529 (N_49529,N_37213,N_30968);
and U49530 (N_49530,N_35045,N_37402);
nand U49531 (N_49531,N_37860,N_36421);
nand U49532 (N_49532,N_33022,N_31369);
or U49533 (N_49533,N_31958,N_30435);
nand U49534 (N_49534,N_39079,N_37921);
and U49535 (N_49535,N_37023,N_30841);
or U49536 (N_49536,N_36279,N_30339);
nand U49537 (N_49537,N_35076,N_37295);
nand U49538 (N_49538,N_37071,N_33628);
and U49539 (N_49539,N_38079,N_37552);
or U49540 (N_49540,N_38756,N_33712);
or U49541 (N_49541,N_30390,N_34726);
and U49542 (N_49542,N_34286,N_39738);
nor U49543 (N_49543,N_38633,N_34362);
nand U49544 (N_49544,N_31538,N_31026);
nand U49545 (N_49545,N_33923,N_35999);
or U49546 (N_49546,N_31335,N_32864);
or U49547 (N_49547,N_30388,N_33744);
nand U49548 (N_49548,N_39873,N_32433);
and U49549 (N_49549,N_35602,N_36832);
nor U49550 (N_49550,N_34434,N_37853);
nand U49551 (N_49551,N_35750,N_36739);
or U49552 (N_49552,N_30622,N_30085);
nor U49553 (N_49553,N_35001,N_36328);
or U49554 (N_49554,N_39836,N_37450);
nand U49555 (N_49555,N_37513,N_30820);
nor U49556 (N_49556,N_31044,N_33502);
nor U49557 (N_49557,N_31833,N_39003);
nand U49558 (N_49558,N_33330,N_33534);
nand U49559 (N_49559,N_33057,N_35883);
xnor U49560 (N_49560,N_36344,N_39138);
nor U49561 (N_49561,N_36046,N_31186);
and U49562 (N_49562,N_35437,N_35231);
nand U49563 (N_49563,N_37581,N_33141);
nor U49564 (N_49564,N_34701,N_38278);
or U49565 (N_49565,N_36162,N_33170);
or U49566 (N_49566,N_34075,N_35772);
or U49567 (N_49567,N_31179,N_33461);
and U49568 (N_49568,N_33738,N_33607);
nand U49569 (N_49569,N_39726,N_38739);
and U49570 (N_49570,N_38307,N_33512);
and U49571 (N_49571,N_38507,N_38721);
nand U49572 (N_49572,N_33894,N_33897);
and U49573 (N_49573,N_31001,N_33162);
and U49574 (N_49574,N_32423,N_35950);
and U49575 (N_49575,N_38740,N_31488);
and U49576 (N_49576,N_35955,N_39299);
nor U49577 (N_49577,N_32630,N_33703);
and U49578 (N_49578,N_38931,N_36946);
nor U49579 (N_49579,N_39905,N_39287);
nand U49580 (N_49580,N_35365,N_38277);
and U49581 (N_49581,N_39046,N_38164);
or U49582 (N_49582,N_34875,N_31820);
or U49583 (N_49583,N_37314,N_36555);
or U49584 (N_49584,N_30510,N_33965);
and U49585 (N_49585,N_33679,N_31353);
nand U49586 (N_49586,N_31102,N_38076);
and U49587 (N_49587,N_32740,N_33351);
nor U49588 (N_49588,N_37442,N_32825);
or U49589 (N_49589,N_31763,N_34470);
nor U49590 (N_49590,N_32858,N_36444);
and U49591 (N_49591,N_38199,N_35203);
nor U49592 (N_49592,N_31177,N_35324);
nand U49593 (N_49593,N_39128,N_34123);
and U49594 (N_49594,N_33206,N_32543);
nor U49595 (N_49595,N_32251,N_34531);
or U49596 (N_49596,N_39054,N_37327);
nand U49597 (N_49597,N_38130,N_34292);
nand U49598 (N_49598,N_37530,N_35004);
and U49599 (N_49599,N_36797,N_38449);
or U49600 (N_49600,N_37055,N_38552);
and U49601 (N_49601,N_36767,N_37130);
nor U49602 (N_49602,N_36516,N_35603);
or U49603 (N_49603,N_36455,N_37980);
nand U49604 (N_49604,N_38460,N_38233);
nor U49605 (N_49605,N_36264,N_38091);
xnor U49606 (N_49606,N_32438,N_39254);
xor U49607 (N_49607,N_39826,N_35057);
nand U49608 (N_49608,N_32552,N_38880);
and U49609 (N_49609,N_35028,N_37921);
or U49610 (N_49610,N_32998,N_32050);
or U49611 (N_49611,N_35810,N_38136);
and U49612 (N_49612,N_38166,N_30484);
or U49613 (N_49613,N_33974,N_31992);
or U49614 (N_49614,N_36813,N_36952);
nand U49615 (N_49615,N_39266,N_32042);
or U49616 (N_49616,N_30137,N_33364);
nand U49617 (N_49617,N_36388,N_33703);
nor U49618 (N_49618,N_37778,N_39235);
nor U49619 (N_49619,N_37199,N_36893);
nand U49620 (N_49620,N_34527,N_38232);
nor U49621 (N_49621,N_39396,N_39856);
or U49622 (N_49622,N_31020,N_37450);
nand U49623 (N_49623,N_35014,N_38985);
or U49624 (N_49624,N_39367,N_36130);
nand U49625 (N_49625,N_37531,N_33851);
nand U49626 (N_49626,N_34147,N_33884);
nand U49627 (N_49627,N_37265,N_31544);
nand U49628 (N_49628,N_38965,N_38302);
and U49629 (N_49629,N_34772,N_32395);
nor U49630 (N_49630,N_32014,N_32640);
xor U49631 (N_49631,N_32492,N_37464);
nor U49632 (N_49632,N_35201,N_31411);
or U49633 (N_49633,N_39547,N_37132);
nand U49634 (N_49634,N_39141,N_32238);
and U49635 (N_49635,N_30958,N_39367);
and U49636 (N_49636,N_30675,N_37082);
nor U49637 (N_49637,N_32628,N_32588);
nor U49638 (N_49638,N_34120,N_39700);
nand U49639 (N_49639,N_38416,N_32186);
nand U49640 (N_49640,N_34052,N_30417);
or U49641 (N_49641,N_38467,N_34955);
nor U49642 (N_49642,N_35148,N_31251);
nor U49643 (N_49643,N_33257,N_39861);
and U49644 (N_49644,N_38126,N_36748);
nand U49645 (N_49645,N_39325,N_30751);
and U49646 (N_49646,N_36451,N_34055);
and U49647 (N_49647,N_33384,N_36028);
nor U49648 (N_49648,N_34151,N_34244);
and U49649 (N_49649,N_38671,N_33170);
xnor U49650 (N_49650,N_38522,N_32844);
nand U49651 (N_49651,N_31519,N_37411);
nor U49652 (N_49652,N_38831,N_38770);
nor U49653 (N_49653,N_30252,N_31213);
and U49654 (N_49654,N_39429,N_38924);
xor U49655 (N_49655,N_33793,N_31305);
or U49656 (N_49656,N_35193,N_31671);
and U49657 (N_49657,N_30410,N_39808);
or U49658 (N_49658,N_30009,N_33415);
nand U49659 (N_49659,N_31210,N_30577);
xnor U49660 (N_49660,N_38004,N_39875);
nand U49661 (N_49661,N_37119,N_38851);
or U49662 (N_49662,N_35306,N_36164);
or U49663 (N_49663,N_37927,N_34522);
nor U49664 (N_49664,N_34301,N_33031);
nand U49665 (N_49665,N_31810,N_34413);
or U49666 (N_49666,N_35698,N_37817);
nand U49667 (N_49667,N_36676,N_34893);
and U49668 (N_49668,N_32510,N_39334);
nor U49669 (N_49669,N_37981,N_37560);
or U49670 (N_49670,N_33480,N_30326);
nor U49671 (N_49671,N_34080,N_38185);
or U49672 (N_49672,N_34350,N_33923);
or U49673 (N_49673,N_31904,N_31416);
nand U49674 (N_49674,N_32830,N_35471);
or U49675 (N_49675,N_30722,N_30859);
or U49676 (N_49676,N_37068,N_34535);
nor U49677 (N_49677,N_33541,N_38735);
nand U49678 (N_49678,N_37293,N_30101);
nand U49679 (N_49679,N_33997,N_30813);
nor U49680 (N_49680,N_37370,N_35869);
nor U49681 (N_49681,N_33512,N_35691);
nor U49682 (N_49682,N_34922,N_30219);
nand U49683 (N_49683,N_32159,N_37006);
or U49684 (N_49684,N_34511,N_38830);
xor U49685 (N_49685,N_33972,N_34113);
nor U49686 (N_49686,N_31961,N_38781);
and U49687 (N_49687,N_38720,N_37261);
and U49688 (N_49688,N_32867,N_33913);
nor U49689 (N_49689,N_34986,N_36953);
xnor U49690 (N_49690,N_37963,N_31046);
nand U49691 (N_49691,N_33365,N_36490);
nand U49692 (N_49692,N_38657,N_36019);
and U49693 (N_49693,N_32534,N_31779);
nand U49694 (N_49694,N_30762,N_30346);
nor U49695 (N_49695,N_37571,N_30528);
nand U49696 (N_49696,N_32527,N_36192);
nor U49697 (N_49697,N_35971,N_30361);
nand U49698 (N_49698,N_39517,N_32460);
and U49699 (N_49699,N_31383,N_35431);
and U49700 (N_49700,N_32415,N_34218);
nand U49701 (N_49701,N_36803,N_35396);
or U49702 (N_49702,N_36103,N_35937);
or U49703 (N_49703,N_32049,N_31140);
xnor U49704 (N_49704,N_37608,N_36544);
nor U49705 (N_49705,N_30185,N_32720);
or U49706 (N_49706,N_34336,N_33607);
nand U49707 (N_49707,N_39468,N_37756);
or U49708 (N_49708,N_35068,N_36510);
and U49709 (N_49709,N_39522,N_30741);
nand U49710 (N_49710,N_39841,N_32354);
nor U49711 (N_49711,N_39469,N_33066);
nor U49712 (N_49712,N_36292,N_39927);
nand U49713 (N_49713,N_39034,N_31803);
nor U49714 (N_49714,N_36234,N_30473);
nand U49715 (N_49715,N_34084,N_30268);
nor U49716 (N_49716,N_38890,N_35327);
nand U49717 (N_49717,N_38923,N_33095);
nor U49718 (N_49718,N_34312,N_39548);
or U49719 (N_49719,N_31258,N_35369);
nand U49720 (N_49720,N_38045,N_35752);
and U49721 (N_49721,N_36960,N_39890);
or U49722 (N_49722,N_34754,N_33823);
nand U49723 (N_49723,N_36984,N_36896);
nand U49724 (N_49724,N_36436,N_32111);
nor U49725 (N_49725,N_38992,N_31104);
and U49726 (N_49726,N_33752,N_33400);
or U49727 (N_49727,N_30248,N_33284);
nand U49728 (N_49728,N_38499,N_37251);
nor U49729 (N_49729,N_30366,N_33104);
and U49730 (N_49730,N_37997,N_34266);
nand U49731 (N_49731,N_33389,N_36173);
and U49732 (N_49732,N_39940,N_36365);
or U49733 (N_49733,N_34058,N_39757);
nor U49734 (N_49734,N_38032,N_37161);
xor U49735 (N_49735,N_39674,N_34795);
nor U49736 (N_49736,N_31220,N_39215);
or U49737 (N_49737,N_30331,N_39649);
or U49738 (N_49738,N_32451,N_39893);
or U49739 (N_49739,N_36346,N_32674);
nor U49740 (N_49740,N_33955,N_39814);
and U49741 (N_49741,N_34240,N_35645);
and U49742 (N_49742,N_34831,N_38977);
nor U49743 (N_49743,N_35394,N_31750);
xnor U49744 (N_49744,N_35189,N_36548);
and U49745 (N_49745,N_30360,N_39103);
nor U49746 (N_49746,N_35850,N_37174);
or U49747 (N_49747,N_35452,N_36813);
nor U49748 (N_49748,N_38527,N_32849);
or U49749 (N_49749,N_32333,N_33092);
or U49750 (N_49750,N_31922,N_35608);
nand U49751 (N_49751,N_39706,N_39014);
and U49752 (N_49752,N_30609,N_38813);
and U49753 (N_49753,N_33240,N_33908);
or U49754 (N_49754,N_35192,N_33249);
or U49755 (N_49755,N_34913,N_36593);
nor U49756 (N_49756,N_38575,N_37928);
nor U49757 (N_49757,N_33725,N_31771);
and U49758 (N_49758,N_34725,N_32557);
xor U49759 (N_49759,N_34989,N_38837);
nand U49760 (N_49760,N_31467,N_39441);
or U49761 (N_49761,N_37726,N_36026);
nand U49762 (N_49762,N_36937,N_32077);
xor U49763 (N_49763,N_39723,N_36592);
nor U49764 (N_49764,N_34471,N_30492);
nor U49765 (N_49765,N_32426,N_34861);
and U49766 (N_49766,N_32054,N_37196);
xnor U49767 (N_49767,N_31509,N_38907);
nand U49768 (N_49768,N_37620,N_32621);
and U49769 (N_49769,N_37412,N_32211);
nor U49770 (N_49770,N_35016,N_30012);
and U49771 (N_49771,N_31568,N_36734);
nor U49772 (N_49772,N_37014,N_31194);
or U49773 (N_49773,N_35250,N_33186);
nand U49774 (N_49774,N_33391,N_36994);
nand U49775 (N_49775,N_30213,N_39211);
and U49776 (N_49776,N_39711,N_38918);
nand U49777 (N_49777,N_39030,N_38966);
or U49778 (N_49778,N_32152,N_38977);
or U49779 (N_49779,N_30425,N_35374);
xor U49780 (N_49780,N_31178,N_30606);
nor U49781 (N_49781,N_31152,N_38006);
nand U49782 (N_49782,N_39230,N_33597);
xnor U49783 (N_49783,N_30997,N_30308);
nor U49784 (N_49784,N_37893,N_33812);
and U49785 (N_49785,N_39283,N_36091);
or U49786 (N_49786,N_30446,N_38864);
or U49787 (N_49787,N_30560,N_31126);
nand U49788 (N_49788,N_33554,N_34429);
nand U49789 (N_49789,N_34643,N_38263);
and U49790 (N_49790,N_32926,N_34303);
and U49791 (N_49791,N_37720,N_36690);
nand U49792 (N_49792,N_38017,N_39792);
nand U49793 (N_49793,N_34406,N_33991);
nor U49794 (N_49794,N_35881,N_37960);
nand U49795 (N_49795,N_39802,N_36542);
nand U49796 (N_49796,N_36081,N_39387);
nand U49797 (N_49797,N_37308,N_34087);
and U49798 (N_49798,N_32226,N_37180);
or U49799 (N_49799,N_34125,N_38453);
nand U49800 (N_49800,N_33165,N_32302);
nand U49801 (N_49801,N_35507,N_31499);
and U49802 (N_49802,N_35169,N_35014);
or U49803 (N_49803,N_30060,N_33320);
nand U49804 (N_49804,N_39021,N_31726);
or U49805 (N_49805,N_33402,N_34141);
or U49806 (N_49806,N_36556,N_37649);
xnor U49807 (N_49807,N_34482,N_39708);
nor U49808 (N_49808,N_38207,N_31313);
or U49809 (N_49809,N_31312,N_34874);
nor U49810 (N_49810,N_35908,N_35443);
or U49811 (N_49811,N_38716,N_34664);
nor U49812 (N_49812,N_32679,N_37025);
and U49813 (N_49813,N_32393,N_36221);
or U49814 (N_49814,N_36294,N_39297);
or U49815 (N_49815,N_34142,N_30385);
or U49816 (N_49816,N_39122,N_38666);
or U49817 (N_49817,N_39355,N_39215);
xnor U49818 (N_49818,N_34459,N_37719);
or U49819 (N_49819,N_37528,N_35563);
nand U49820 (N_49820,N_30506,N_39755);
nor U49821 (N_49821,N_33466,N_34605);
or U49822 (N_49822,N_31914,N_36516);
xnor U49823 (N_49823,N_31413,N_36352);
nand U49824 (N_49824,N_39541,N_34492);
and U49825 (N_49825,N_30817,N_34403);
nand U49826 (N_49826,N_38841,N_30329);
or U49827 (N_49827,N_37823,N_36327);
or U49828 (N_49828,N_31820,N_37281);
nand U49829 (N_49829,N_38536,N_33965);
or U49830 (N_49830,N_31052,N_39228);
nand U49831 (N_49831,N_35774,N_30027);
nand U49832 (N_49832,N_35347,N_35182);
and U49833 (N_49833,N_35306,N_33594);
and U49834 (N_49834,N_33345,N_37600);
nor U49835 (N_49835,N_39715,N_37930);
or U49836 (N_49836,N_32191,N_36136);
and U49837 (N_49837,N_31473,N_33635);
and U49838 (N_49838,N_30833,N_32780);
and U49839 (N_49839,N_31347,N_30517);
or U49840 (N_49840,N_30591,N_32908);
nand U49841 (N_49841,N_38506,N_30540);
or U49842 (N_49842,N_35220,N_30906);
or U49843 (N_49843,N_33033,N_32338);
and U49844 (N_49844,N_33581,N_37950);
nand U49845 (N_49845,N_35490,N_39471);
and U49846 (N_49846,N_39584,N_32001);
or U49847 (N_49847,N_37388,N_33580);
nor U49848 (N_49848,N_35180,N_38223);
nand U49849 (N_49849,N_34788,N_39377);
or U49850 (N_49850,N_32121,N_36557);
nand U49851 (N_49851,N_36199,N_33380);
or U49852 (N_49852,N_32508,N_34681);
or U49853 (N_49853,N_38669,N_31280);
and U49854 (N_49854,N_36426,N_31694);
or U49855 (N_49855,N_30410,N_35223);
or U49856 (N_49856,N_31273,N_37451);
nor U49857 (N_49857,N_31136,N_32855);
nor U49858 (N_49858,N_30350,N_35045);
xnor U49859 (N_49859,N_32345,N_30007);
nor U49860 (N_49860,N_39727,N_38534);
nand U49861 (N_49861,N_37057,N_33184);
xor U49862 (N_49862,N_32816,N_34081);
nor U49863 (N_49863,N_34159,N_33193);
and U49864 (N_49864,N_38699,N_36131);
or U49865 (N_49865,N_31516,N_37558);
or U49866 (N_49866,N_34842,N_38818);
and U49867 (N_49867,N_37769,N_36076);
nand U49868 (N_49868,N_31458,N_33708);
nand U49869 (N_49869,N_31201,N_36008);
and U49870 (N_49870,N_32803,N_33381);
nand U49871 (N_49871,N_33366,N_37503);
nand U49872 (N_49872,N_36146,N_33494);
nor U49873 (N_49873,N_31608,N_33968);
nand U49874 (N_49874,N_36716,N_31678);
or U49875 (N_49875,N_31878,N_32022);
nand U49876 (N_49876,N_34117,N_35402);
nand U49877 (N_49877,N_31506,N_35929);
nor U49878 (N_49878,N_37254,N_39128);
and U49879 (N_49879,N_37075,N_37373);
and U49880 (N_49880,N_35758,N_38933);
nor U49881 (N_49881,N_39354,N_33368);
nor U49882 (N_49882,N_38097,N_38027);
and U49883 (N_49883,N_37687,N_32321);
and U49884 (N_49884,N_34979,N_37891);
nand U49885 (N_49885,N_35691,N_31004);
nand U49886 (N_49886,N_32263,N_32327);
nand U49887 (N_49887,N_37163,N_36641);
nor U49888 (N_49888,N_34499,N_32998);
xnor U49889 (N_49889,N_34695,N_31065);
and U49890 (N_49890,N_34212,N_34825);
or U49891 (N_49891,N_39727,N_33274);
nand U49892 (N_49892,N_32359,N_33327);
xor U49893 (N_49893,N_31938,N_30699);
nor U49894 (N_49894,N_39355,N_33403);
nor U49895 (N_49895,N_33377,N_39128);
and U49896 (N_49896,N_36950,N_31647);
or U49897 (N_49897,N_31592,N_38558);
or U49898 (N_49898,N_30334,N_31720);
nand U49899 (N_49899,N_33252,N_33434);
nor U49900 (N_49900,N_31518,N_34096);
nand U49901 (N_49901,N_33373,N_35912);
nand U49902 (N_49902,N_39942,N_34978);
xor U49903 (N_49903,N_34148,N_31842);
and U49904 (N_49904,N_36345,N_35023);
nand U49905 (N_49905,N_38528,N_38805);
nand U49906 (N_49906,N_37156,N_39383);
nor U49907 (N_49907,N_31449,N_36644);
nand U49908 (N_49908,N_33607,N_32730);
nor U49909 (N_49909,N_31393,N_36651);
xor U49910 (N_49910,N_32477,N_37147);
nand U49911 (N_49911,N_30667,N_32372);
nor U49912 (N_49912,N_38792,N_32231);
nand U49913 (N_49913,N_39153,N_31856);
nor U49914 (N_49914,N_39472,N_37925);
xor U49915 (N_49915,N_31029,N_38963);
nor U49916 (N_49916,N_31054,N_39853);
or U49917 (N_49917,N_31445,N_39926);
and U49918 (N_49918,N_37644,N_34183);
nor U49919 (N_49919,N_30460,N_35863);
nand U49920 (N_49920,N_30626,N_34508);
and U49921 (N_49921,N_37626,N_30508);
or U49922 (N_49922,N_32069,N_32226);
and U49923 (N_49923,N_33601,N_30280);
nor U49924 (N_49924,N_35492,N_37140);
nor U49925 (N_49925,N_35936,N_36490);
nor U49926 (N_49926,N_38505,N_32200);
or U49927 (N_49927,N_33650,N_38103);
or U49928 (N_49928,N_39603,N_32785);
or U49929 (N_49929,N_37406,N_30100);
xor U49930 (N_49930,N_34936,N_38845);
and U49931 (N_49931,N_32314,N_33019);
and U49932 (N_49932,N_37727,N_39541);
nand U49933 (N_49933,N_32205,N_38675);
or U49934 (N_49934,N_33334,N_37173);
and U49935 (N_49935,N_33230,N_32354);
xnor U49936 (N_49936,N_35672,N_33161);
or U49937 (N_49937,N_36593,N_39318);
nand U49938 (N_49938,N_35268,N_30285);
or U49939 (N_49939,N_32134,N_32502);
nor U49940 (N_49940,N_38412,N_36648);
nand U49941 (N_49941,N_39340,N_38332);
or U49942 (N_49942,N_37392,N_38824);
nand U49943 (N_49943,N_35548,N_39581);
and U49944 (N_49944,N_35681,N_32551);
and U49945 (N_49945,N_35989,N_37609);
or U49946 (N_49946,N_36211,N_35513);
or U49947 (N_49947,N_39309,N_30263);
nor U49948 (N_49948,N_35993,N_31881);
or U49949 (N_49949,N_30282,N_30037);
nor U49950 (N_49950,N_37432,N_32344);
and U49951 (N_49951,N_36527,N_30940);
nand U49952 (N_49952,N_34015,N_38011);
or U49953 (N_49953,N_34158,N_32423);
or U49954 (N_49954,N_36374,N_32319);
nand U49955 (N_49955,N_36483,N_39194);
nand U49956 (N_49956,N_31732,N_36963);
nand U49957 (N_49957,N_36510,N_34462);
or U49958 (N_49958,N_37520,N_32423);
or U49959 (N_49959,N_37138,N_38529);
and U49960 (N_49960,N_31015,N_33344);
and U49961 (N_49961,N_38250,N_37043);
and U49962 (N_49962,N_38088,N_34126);
nor U49963 (N_49963,N_38244,N_30153);
and U49964 (N_49964,N_32038,N_36960);
or U49965 (N_49965,N_32382,N_30640);
nor U49966 (N_49966,N_33514,N_30405);
or U49967 (N_49967,N_37103,N_31481);
or U49968 (N_49968,N_31599,N_35937);
nor U49969 (N_49969,N_34683,N_38372);
nor U49970 (N_49970,N_37885,N_36953);
and U49971 (N_49971,N_39892,N_32682);
and U49972 (N_49972,N_30464,N_38937);
or U49973 (N_49973,N_31997,N_36526);
and U49974 (N_49974,N_32763,N_32244);
nand U49975 (N_49975,N_35827,N_31109);
nand U49976 (N_49976,N_34614,N_32257);
and U49977 (N_49977,N_39645,N_30355);
nor U49978 (N_49978,N_37908,N_31373);
xor U49979 (N_49979,N_30822,N_32235);
nor U49980 (N_49980,N_34052,N_31638);
and U49981 (N_49981,N_36998,N_31212);
nand U49982 (N_49982,N_33627,N_30036);
nand U49983 (N_49983,N_38496,N_35202);
nand U49984 (N_49984,N_34728,N_38220);
and U49985 (N_49985,N_32114,N_36815);
or U49986 (N_49986,N_33326,N_33737);
nand U49987 (N_49987,N_35018,N_30849);
or U49988 (N_49988,N_32409,N_34452);
nor U49989 (N_49989,N_36285,N_37197);
nor U49990 (N_49990,N_30557,N_34369);
or U49991 (N_49991,N_34105,N_36774);
nand U49992 (N_49992,N_34196,N_35477);
or U49993 (N_49993,N_33841,N_35823);
and U49994 (N_49994,N_31415,N_31235);
nand U49995 (N_49995,N_31260,N_30229);
and U49996 (N_49996,N_35352,N_30922);
or U49997 (N_49997,N_30418,N_33372);
nand U49998 (N_49998,N_31285,N_38052);
and U49999 (N_49999,N_38885,N_33952);
nand UO_0 (O_0,N_44784,N_46133);
xor UO_1 (O_1,N_49775,N_43740);
or UO_2 (O_2,N_48459,N_49232);
and UO_3 (O_3,N_40069,N_40198);
nand UO_4 (O_4,N_49418,N_49040);
and UO_5 (O_5,N_40982,N_48383);
nand UO_6 (O_6,N_41133,N_41292);
or UO_7 (O_7,N_42643,N_41387);
nor UO_8 (O_8,N_48400,N_43367);
or UO_9 (O_9,N_47912,N_40443);
nor UO_10 (O_10,N_41913,N_46740);
nor UO_11 (O_11,N_42721,N_40054);
and UO_12 (O_12,N_47890,N_41120);
or UO_13 (O_13,N_46874,N_42405);
and UO_14 (O_14,N_43561,N_48328);
and UO_15 (O_15,N_47291,N_46758);
nor UO_16 (O_16,N_49609,N_44161);
or UO_17 (O_17,N_46213,N_42006);
nor UO_18 (O_18,N_47586,N_41032);
xnor UO_19 (O_19,N_49660,N_40649);
nand UO_20 (O_20,N_48418,N_49422);
nor UO_21 (O_21,N_41670,N_42935);
xor UO_22 (O_22,N_43227,N_49490);
nand UO_23 (O_23,N_40251,N_47934);
or UO_24 (O_24,N_43691,N_41452);
and UO_25 (O_25,N_45004,N_41963);
nor UO_26 (O_26,N_47919,N_43764);
nor UO_27 (O_27,N_41145,N_46806);
xnor UO_28 (O_28,N_47008,N_40902);
xor UO_29 (O_29,N_45929,N_44779);
or UO_30 (O_30,N_47419,N_48208);
nor UO_31 (O_31,N_49534,N_40551);
nand UO_32 (O_32,N_41716,N_49596);
and UO_33 (O_33,N_46148,N_41192);
nor UO_34 (O_34,N_47676,N_43244);
xnor UO_35 (O_35,N_41212,N_45480);
nor UO_36 (O_36,N_42111,N_47028);
and UO_37 (O_37,N_43897,N_49894);
and UO_38 (O_38,N_43117,N_43278);
or UO_39 (O_39,N_40557,N_47661);
xnor UO_40 (O_40,N_40810,N_41178);
and UO_41 (O_41,N_43995,N_47053);
xnor UO_42 (O_42,N_40527,N_41807);
nor UO_43 (O_43,N_48781,N_48940);
xor UO_44 (O_44,N_45448,N_48372);
and UO_45 (O_45,N_44757,N_46277);
and UO_46 (O_46,N_40926,N_43493);
nor UO_47 (O_47,N_42093,N_43961);
and UO_48 (O_48,N_42477,N_40834);
or UO_49 (O_49,N_45858,N_45769);
nor UO_50 (O_50,N_48345,N_46916);
nor UO_51 (O_51,N_40466,N_42435);
or UO_52 (O_52,N_49706,N_47873);
or UO_53 (O_53,N_41326,N_40680);
nor UO_54 (O_54,N_48915,N_40892);
nor UO_55 (O_55,N_41013,N_47668);
or UO_56 (O_56,N_43424,N_45810);
or UO_57 (O_57,N_40389,N_47738);
nand UO_58 (O_58,N_43472,N_47737);
nor UO_59 (O_59,N_49523,N_44297);
and UO_60 (O_60,N_48513,N_42122);
xnor UO_61 (O_61,N_41533,N_48299);
or UO_62 (O_62,N_41660,N_49725);
nand UO_63 (O_63,N_46479,N_48179);
nand UO_64 (O_64,N_46754,N_45643);
nand UO_65 (O_65,N_43575,N_40667);
or UO_66 (O_66,N_45823,N_49058);
and UO_67 (O_67,N_40660,N_41612);
or UO_68 (O_68,N_42912,N_47946);
and UO_69 (O_69,N_44206,N_46250);
nor UO_70 (O_70,N_46574,N_45699);
or UO_71 (O_71,N_42551,N_49566);
nor UO_72 (O_72,N_48376,N_40151);
or UO_73 (O_73,N_44371,N_46303);
and UO_74 (O_74,N_41845,N_40613);
nor UO_75 (O_75,N_44592,N_46198);
nor UO_76 (O_76,N_47201,N_48844);
nand UO_77 (O_77,N_42178,N_47740);
xor UO_78 (O_78,N_41558,N_40003);
nand UO_79 (O_79,N_44519,N_40411);
nor UO_80 (O_80,N_40476,N_49528);
nand UO_81 (O_81,N_48286,N_49608);
or UO_82 (O_82,N_47980,N_44201);
xnor UO_83 (O_83,N_45595,N_47424);
or UO_84 (O_84,N_44692,N_43400);
and UO_85 (O_85,N_46189,N_40158);
nand UO_86 (O_86,N_42423,N_41490);
nand UO_87 (O_87,N_47877,N_40758);
nor UO_88 (O_88,N_40799,N_42390);
nor UO_89 (O_89,N_42656,N_41456);
or UO_90 (O_90,N_47322,N_46736);
or UO_91 (O_91,N_40364,N_42595);
nand UO_92 (O_92,N_47109,N_47075);
or UO_93 (O_93,N_46535,N_48920);
xor UO_94 (O_94,N_45801,N_41856);
nand UO_95 (O_95,N_43011,N_48892);
and UO_96 (O_96,N_45720,N_40923);
and UO_97 (O_97,N_43337,N_43536);
nor UO_98 (O_98,N_43248,N_49001);
nor UO_99 (O_99,N_41019,N_41423);
nor UO_100 (O_100,N_45877,N_45686);
nand UO_101 (O_101,N_44656,N_43962);
and UO_102 (O_102,N_48644,N_48718);
or UO_103 (O_103,N_47776,N_49306);
nand UO_104 (O_104,N_45715,N_46931);
nor UO_105 (O_105,N_43670,N_48744);
nor UO_106 (O_106,N_45684,N_48619);
nor UO_107 (O_107,N_41770,N_44368);
nand UO_108 (O_108,N_43946,N_48965);
or UO_109 (O_109,N_43102,N_48051);
nor UO_110 (O_110,N_45656,N_49617);
nand UO_111 (O_111,N_44044,N_43888);
nand UO_112 (O_112,N_48034,N_48214);
or UO_113 (O_113,N_46426,N_45774);
nand UO_114 (O_114,N_49696,N_47393);
nor UO_115 (O_115,N_40007,N_49974);
nand UO_116 (O_116,N_40307,N_44636);
nand UO_117 (O_117,N_47832,N_48284);
nor UO_118 (O_118,N_41459,N_46613);
or UO_119 (O_119,N_42707,N_47047);
nor UO_120 (O_120,N_46842,N_49999);
and UO_121 (O_121,N_44011,N_46324);
and UO_122 (O_122,N_42027,N_40394);
xnor UO_123 (O_123,N_41154,N_42412);
nor UO_124 (O_124,N_41455,N_44872);
nand UO_125 (O_125,N_42969,N_43019);
and UO_126 (O_126,N_40679,N_48038);
or UO_127 (O_127,N_49474,N_46489);
and UO_128 (O_128,N_41174,N_44577);
nand UO_129 (O_129,N_44103,N_47566);
or UO_130 (O_130,N_49263,N_44419);
nand UO_131 (O_131,N_44416,N_41277);
and UO_132 (O_132,N_49722,N_43195);
nand UO_133 (O_133,N_47722,N_43144);
nor UO_134 (O_134,N_49159,N_48006);
nor UO_135 (O_135,N_49331,N_40049);
xnor UO_136 (O_136,N_45447,N_40037);
and UO_137 (O_137,N_41240,N_42863);
and UO_138 (O_138,N_43720,N_43461);
and UO_139 (O_139,N_40938,N_48267);
nand UO_140 (O_140,N_48012,N_47148);
or UO_141 (O_141,N_46436,N_48721);
or UO_142 (O_142,N_40584,N_44585);
nor UO_143 (O_143,N_43941,N_40859);
nand UO_144 (O_144,N_49977,N_48845);
and UO_145 (O_145,N_43005,N_46938);
or UO_146 (O_146,N_48447,N_42533);
and UO_147 (O_147,N_49926,N_43214);
nand UO_148 (O_148,N_45961,N_44530);
and UO_149 (O_149,N_49979,N_47183);
nand UO_150 (O_150,N_49491,N_43146);
or UO_151 (O_151,N_41257,N_45300);
or UO_152 (O_152,N_44306,N_44686);
nand UO_153 (O_153,N_44436,N_41772);
or UO_154 (O_154,N_46995,N_41655);
nor UO_155 (O_155,N_45621,N_49768);
xor UO_156 (O_156,N_40609,N_40981);
xor UO_157 (O_157,N_40869,N_40590);
or UO_158 (O_158,N_46811,N_45217);
and UO_159 (O_159,N_47007,N_47213);
nand UO_160 (O_160,N_47346,N_45239);
and UO_161 (O_161,N_47150,N_45211);
xor UO_162 (O_162,N_41918,N_46819);
and UO_163 (O_163,N_45160,N_43680);
xor UO_164 (O_164,N_44843,N_41247);
nand UO_165 (O_165,N_43257,N_43107);
or UO_166 (O_166,N_43523,N_44605);
nor UO_167 (O_167,N_44698,N_47695);
nand UO_168 (O_168,N_40681,N_43016);
nor UO_169 (O_169,N_42026,N_48771);
or UO_170 (O_170,N_44753,N_48494);
nor UO_171 (O_171,N_47503,N_49809);
nand UO_172 (O_172,N_49000,N_45265);
nor UO_173 (O_173,N_42943,N_47196);
and UO_174 (O_174,N_42997,N_46569);
xor UO_175 (O_175,N_46525,N_48117);
nand UO_176 (O_176,N_49430,N_47617);
and UO_177 (O_177,N_42017,N_49420);
nand UO_178 (O_178,N_47172,N_40781);
nand UO_179 (O_179,N_44350,N_48484);
nor UO_180 (O_180,N_42849,N_42054);
or UO_181 (O_181,N_47870,N_43057);
nor UO_182 (O_182,N_47572,N_40606);
nand UO_183 (O_183,N_47210,N_47765);
and UO_184 (O_184,N_47499,N_40496);
or UO_185 (O_185,N_40754,N_45902);
and UO_186 (O_186,N_40184,N_44431);
nor UO_187 (O_187,N_46820,N_47513);
xnor UO_188 (O_188,N_44058,N_47454);
nor UO_189 (O_189,N_44279,N_40168);
and UO_190 (O_190,N_42385,N_44898);
and UO_191 (O_191,N_40817,N_46888);
or UO_192 (O_192,N_48489,N_49754);
nand UO_193 (O_193,N_46331,N_47052);
or UO_194 (O_194,N_42244,N_47504);
nor UO_195 (O_195,N_42657,N_49689);
and UO_196 (O_196,N_43823,N_48618);
nand UO_197 (O_197,N_40809,N_47037);
nand UO_198 (O_198,N_49764,N_43258);
nand UO_199 (O_199,N_46263,N_44819);
and UO_200 (O_200,N_44772,N_49055);
and UO_201 (O_201,N_44937,N_49469);
or UO_202 (O_202,N_40638,N_46009);
or UO_203 (O_203,N_42584,N_41251);
nand UO_204 (O_204,N_48926,N_46582);
or UO_205 (O_205,N_48368,N_47861);
nor UO_206 (O_206,N_43846,N_46719);
xnor UO_207 (O_207,N_49903,N_45534);
nand UO_208 (O_208,N_44521,N_49154);
nand UO_209 (O_209,N_49393,N_47214);
or UO_210 (O_210,N_44746,N_48062);
and UO_211 (O_211,N_40963,N_47239);
nand UO_212 (O_212,N_46567,N_48266);
or UO_213 (O_213,N_45151,N_46134);
or UO_214 (O_214,N_41090,N_46738);
nor UO_215 (O_215,N_46257,N_41434);
nand UO_216 (O_216,N_47490,N_47173);
or UO_217 (O_217,N_48808,N_43128);
nand UO_218 (O_218,N_43466,N_46169);
nand UO_219 (O_219,N_42072,N_49398);
or UO_220 (O_220,N_40222,N_48321);
xnor UO_221 (O_221,N_40941,N_45983);
nand UO_222 (O_222,N_44296,N_49313);
nor UO_223 (O_223,N_41208,N_44104);
or UO_224 (O_224,N_43857,N_46722);
xor UO_225 (O_225,N_44211,N_45374);
or UO_226 (O_226,N_46790,N_44556);
nor UO_227 (O_227,N_46514,N_46383);
nand UO_228 (O_228,N_48191,N_40341);
nor UO_229 (O_229,N_49543,N_49243);
nor UO_230 (O_230,N_46953,N_43338);
nor UO_231 (O_231,N_44921,N_49225);
nand UO_232 (O_232,N_43620,N_45269);
nor UO_233 (O_233,N_40857,N_49426);
and UO_234 (O_234,N_45369,N_47843);
xnor UO_235 (O_235,N_42920,N_43546);
and UO_236 (O_236,N_49610,N_44609);
or UO_237 (O_237,N_44796,N_44008);
nor UO_238 (O_238,N_44839,N_45698);
and UO_239 (O_239,N_49217,N_43763);
or UO_240 (O_240,N_49712,N_45427);
and UO_241 (O_241,N_43473,N_40072);
nand UO_242 (O_242,N_45325,N_45779);
nor UO_243 (O_243,N_45851,N_41926);
nand UO_244 (O_244,N_46638,N_46203);
and UO_245 (O_245,N_42200,N_41173);
or UO_246 (O_246,N_42520,N_44853);
or UO_247 (O_247,N_45816,N_47905);
nor UO_248 (O_248,N_43965,N_41440);
or UO_249 (O_249,N_46441,N_43126);
xnor UO_250 (O_250,N_49260,N_43065);
nor UO_251 (O_251,N_44244,N_42288);
or UO_252 (O_252,N_44905,N_46417);
or UO_253 (O_253,N_40685,N_45388);
and UO_254 (O_254,N_43528,N_43990);
nand UO_255 (O_255,N_45033,N_44579);
and UO_256 (O_256,N_43767,N_45657);
or UO_257 (O_257,N_45892,N_41383);
nand UO_258 (O_258,N_48579,N_40644);
nor UO_259 (O_259,N_48592,N_45919);
nor UO_260 (O_260,N_41569,N_48736);
or UO_261 (O_261,N_44122,N_47753);
nor UO_262 (O_262,N_43164,N_44029);
nand UO_263 (O_263,N_49019,N_43984);
or UO_264 (O_264,N_40813,N_40547);
nand UO_265 (O_265,N_46763,N_44986);
nand UO_266 (O_266,N_49025,N_44290);
or UO_267 (O_267,N_41372,N_40126);
or UO_268 (O_268,N_44895,N_40604);
xor UO_269 (O_269,N_43912,N_49740);
nor UO_270 (O_270,N_40176,N_44170);
and UO_271 (O_271,N_43176,N_49056);
nor UO_272 (O_272,N_40587,N_42933);
nand UO_273 (O_273,N_49668,N_44259);
nor UO_274 (O_274,N_49219,N_43571);
nor UO_275 (O_275,N_49106,N_49865);
nand UO_276 (O_276,N_46202,N_40346);
nor UO_277 (O_277,N_47975,N_41519);
and UO_278 (O_278,N_40253,N_44687);
and UO_279 (O_279,N_44677,N_42189);
and UO_280 (O_280,N_46379,N_43987);
nor UO_281 (O_281,N_47604,N_43417);
or UO_282 (O_282,N_48571,N_40447);
or UO_283 (O_283,N_41900,N_45071);
and UO_284 (O_284,N_42641,N_40138);
and UO_285 (O_285,N_47672,N_42771);
xnor UO_286 (O_286,N_46832,N_48991);
or UO_287 (O_287,N_40544,N_43947);
nand UO_288 (O_288,N_46472,N_46421);
nand UO_289 (O_289,N_44846,N_44671);
xor UO_290 (O_290,N_45986,N_43430);
or UO_291 (O_291,N_48391,N_43796);
nor UO_292 (O_292,N_49088,N_47349);
nand UO_293 (O_293,N_45159,N_42469);
nand UO_294 (O_294,N_43913,N_46595);
nand UO_295 (O_295,N_46116,N_42999);
or UO_296 (O_296,N_42406,N_46409);
nand UO_297 (O_297,N_45402,N_48800);
nand UO_298 (O_298,N_43208,N_47016);
or UO_299 (O_299,N_45597,N_40572);
nand UO_300 (O_300,N_43569,N_42958);
xor UO_301 (O_301,N_45027,N_48962);
xor UO_302 (O_302,N_46999,N_48701);
nand UO_303 (O_303,N_47571,N_43242);
nor UO_304 (O_304,N_44775,N_41227);
or UO_305 (O_305,N_41288,N_49882);
nand UO_306 (O_306,N_43998,N_46265);
or UO_307 (O_307,N_46290,N_41930);
or UO_308 (O_308,N_47402,N_41441);
and UO_309 (O_309,N_45354,N_40872);
nand UO_310 (O_310,N_44048,N_46284);
nor UO_311 (O_311,N_42395,N_49606);
xor UO_312 (O_312,N_40302,N_42246);
nand UO_313 (O_313,N_49210,N_47774);
nand UO_314 (O_314,N_45462,N_41636);
nand UO_315 (O_315,N_47560,N_47473);
or UO_316 (O_316,N_49682,N_49544);
nor UO_317 (O_317,N_41307,N_48975);
and UO_318 (O_318,N_44845,N_43909);
and UO_319 (O_319,N_40712,N_41699);
or UO_320 (O_320,N_48311,N_46346);
nand UO_321 (O_321,N_45938,N_49024);
or UO_322 (O_322,N_49761,N_42851);
nand UO_323 (O_323,N_40214,N_42558);
and UO_324 (O_324,N_47918,N_43722);
and UO_325 (O_325,N_40110,N_49828);
nor UO_326 (O_326,N_48942,N_41182);
nand UO_327 (O_327,N_46125,N_47688);
nor UO_328 (O_328,N_42120,N_44216);
or UO_329 (O_329,N_42692,N_43127);
or UO_330 (O_330,N_48919,N_45293);
or UO_331 (O_331,N_41457,N_46870);
nor UO_332 (O_332,N_42381,N_42891);
or UO_333 (O_333,N_42050,N_44486);
and UO_334 (O_334,N_48141,N_42623);
nor UO_335 (O_335,N_47225,N_41891);
or UO_336 (O_336,N_47943,N_42287);
xnor UO_337 (O_337,N_46070,N_41953);
nand UO_338 (O_338,N_46992,N_45917);
or UO_339 (O_339,N_40970,N_48510);
or UO_340 (O_340,N_48547,N_42554);
xnor UO_341 (O_341,N_49231,N_49659);
nor UO_342 (O_342,N_49450,N_48938);
nand UO_343 (O_343,N_42087,N_49978);
nand UO_344 (O_344,N_41461,N_44653);
and UO_345 (O_345,N_46403,N_41373);
nand UO_346 (O_346,N_46356,N_46630);
nand UO_347 (O_347,N_44813,N_41754);
nand UO_348 (O_348,N_40514,N_41489);
xnor UO_349 (O_349,N_45654,N_47155);
nor UO_350 (O_350,N_44217,N_47992);
and UO_351 (O_351,N_48332,N_47486);
nor UO_352 (O_352,N_43351,N_42566);
nand UO_353 (O_353,N_49718,N_41828);
nor UO_354 (O_354,N_43723,N_42251);
xnor UO_355 (O_355,N_46020,N_40260);
nand UO_356 (O_356,N_42042,N_47494);
nor UO_357 (O_357,N_40569,N_48411);
nand UO_358 (O_358,N_42857,N_44620);
nand UO_359 (O_359,N_42784,N_41657);
nor UO_360 (O_360,N_45425,N_41391);
nor UO_361 (O_361,N_48517,N_41969);
nor UO_362 (O_362,N_44016,N_42445);
and UO_363 (O_363,N_43170,N_41728);
and UO_364 (O_364,N_44780,N_42025);
nor UO_365 (O_365,N_41711,N_42702);
nand UO_366 (O_366,N_46121,N_41948);
nand UO_367 (O_367,N_44578,N_45722);
nand UO_368 (O_368,N_40267,N_45825);
nand UO_369 (O_369,N_43784,N_45006);
nand UO_370 (O_370,N_45629,N_44334);
and UO_371 (O_371,N_47257,N_42911);
nor UO_372 (O_372,N_45944,N_48720);
or UO_373 (O_373,N_47019,N_49026);
and UO_374 (O_374,N_41725,N_46761);
and UO_375 (O_375,N_48145,N_47270);
xor UO_376 (O_376,N_45645,N_44920);
nand UO_377 (O_377,N_44908,N_45508);
nor UO_378 (O_378,N_43886,N_44747);
nor UO_379 (O_379,N_45023,N_47124);
or UO_380 (O_380,N_42767,N_43535);
or UO_381 (O_381,N_43850,N_48807);
or UO_382 (O_382,N_41837,N_47308);
and UO_383 (O_383,N_45193,N_46321);
and UO_384 (O_384,N_49859,N_40837);
and UO_385 (O_385,N_48973,N_45514);
or UO_386 (O_386,N_49151,N_49269);
xnor UO_387 (O_387,N_49816,N_40786);
nor UO_388 (O_388,N_46958,N_44730);
or UO_389 (O_389,N_46960,N_40836);
and UO_390 (O_390,N_49481,N_47704);
and UO_391 (O_391,N_41914,N_41933);
or UO_392 (O_392,N_49570,N_42177);
nor UO_393 (O_393,N_47897,N_42173);
and UO_394 (O_394,N_44418,N_45451);
nor UO_395 (O_395,N_48222,N_40111);
or UO_396 (O_396,N_41738,N_49757);
and UO_397 (O_397,N_42846,N_45258);
nand UO_398 (O_398,N_49078,N_48971);
nor UO_399 (O_399,N_43437,N_48458);
xnor UO_400 (O_400,N_49739,N_44551);
nand UO_401 (O_401,N_41915,N_40973);
and UO_402 (O_402,N_43206,N_41675);
nand UO_403 (O_403,N_42015,N_47309);
and UO_404 (O_404,N_40100,N_45605);
nand UO_405 (O_405,N_45081,N_45639);
and UO_406 (O_406,N_41961,N_49297);
nor UO_407 (O_407,N_42065,N_49588);
xnor UO_408 (O_408,N_44061,N_43226);
nand UO_409 (O_409,N_40403,N_46195);
nor UO_410 (O_410,N_49475,N_43296);
or UO_411 (O_411,N_47373,N_42145);
or UO_412 (O_412,N_48924,N_46127);
nor UO_413 (O_413,N_45222,N_44384);
and UO_414 (O_414,N_43618,N_49513);
and UO_415 (O_415,N_47036,N_44101);
nor UO_416 (O_416,N_46711,N_45827);
nand UO_417 (O_417,N_43234,N_44922);
and UO_418 (O_418,N_41443,N_44721);
or UO_419 (O_419,N_40994,N_44187);
and UO_420 (O_420,N_46547,N_46800);
and UO_421 (O_421,N_47274,N_48847);
xor UO_422 (O_422,N_47282,N_45273);
and UO_423 (O_423,N_45521,N_48862);
and UO_424 (O_424,N_42052,N_47336);
nor UO_425 (O_425,N_44553,N_43204);
or UO_426 (O_426,N_40920,N_41894);
nand UO_427 (O_427,N_46824,N_43381);
nand UO_428 (O_428,N_46564,N_46966);
xor UO_429 (O_429,N_40676,N_40853);
or UO_430 (O_430,N_40435,N_49562);
nand UO_431 (O_431,N_40276,N_41258);
and UO_432 (O_432,N_46972,N_40162);
nor UO_433 (O_433,N_48318,N_44032);
xnor UO_434 (O_434,N_43270,N_42678);
nand UO_435 (O_435,N_44050,N_49940);
nor UO_436 (O_436,N_46273,N_42427);
or UO_437 (O_437,N_42340,N_41767);
nor UO_438 (O_438,N_49301,N_45833);
and UO_439 (O_439,N_44265,N_47637);
xor UO_440 (O_440,N_47743,N_42495);
and UO_441 (O_441,N_42549,N_47711);
and UO_442 (O_442,N_46807,N_41927);
or UO_443 (O_443,N_46082,N_49885);
or UO_444 (O_444,N_46053,N_43364);
and UO_445 (O_445,N_49525,N_45275);
nand UO_446 (O_446,N_48980,N_48796);
nand UO_447 (O_447,N_46956,N_46367);
xnor UO_448 (O_448,N_40956,N_45137);
nand UO_449 (O_449,N_49998,N_44938);
and UO_450 (O_450,N_49637,N_45455);
nor UO_451 (O_451,N_44989,N_46700);
and UO_452 (O_452,N_45400,N_41128);
or UO_453 (O_453,N_45280,N_46899);
nor UO_454 (O_454,N_47553,N_40132);
nand UO_455 (O_455,N_44369,N_48017);
or UO_456 (O_456,N_45942,N_47584);
and UO_457 (O_457,N_49679,N_44068);
and UO_458 (O_458,N_41967,N_40377);
and UO_459 (O_459,N_41338,N_47375);
nand UO_460 (O_460,N_43556,N_43916);
or UO_461 (O_461,N_49500,N_45196);
or UO_462 (O_462,N_46219,N_49063);
nand UO_463 (O_463,N_43570,N_46340);
nand UO_464 (O_464,N_46280,N_47469);
nand UO_465 (O_465,N_40216,N_46221);
or UO_466 (O_466,N_48557,N_44465);
nor UO_467 (O_467,N_43657,N_45335);
xnor UO_468 (O_468,N_40090,N_42074);
nor UO_469 (O_469,N_43286,N_44013);
nor UO_470 (O_470,N_42561,N_45352);
nand UO_471 (O_471,N_49714,N_40131);
or UO_472 (O_472,N_40980,N_46007);
or UO_473 (O_473,N_43026,N_40542);
or UO_474 (O_474,N_45504,N_46518);
or UO_475 (O_475,N_44200,N_48841);
nor UO_476 (O_476,N_45199,N_43271);
and UO_477 (O_477,N_43901,N_47682);
or UO_478 (O_478,N_40412,N_41829);
nand UO_479 (O_479,N_45407,N_45515);
xnor UO_480 (O_480,N_43550,N_43549);
nor UO_481 (O_481,N_47057,N_40273);
and UO_482 (O_482,N_47273,N_47041);
or UO_483 (O_483,N_40028,N_47121);
and UO_484 (O_484,N_40862,N_42741);
or UO_485 (O_485,N_44935,N_47167);
nor UO_486 (O_486,N_42364,N_41631);
nand UO_487 (O_487,N_42511,N_46110);
or UO_488 (O_488,N_46102,N_48907);
and UO_489 (O_489,N_42600,N_43994);
and UO_490 (O_490,N_47440,N_43861);
xnor UO_491 (O_491,N_48706,N_47421);
nand UO_492 (O_492,N_46928,N_47778);
and UO_493 (O_493,N_41365,N_42014);
and UO_494 (O_494,N_47658,N_49361);
or UO_495 (O_495,N_41471,N_45382);
and UO_496 (O_496,N_47967,N_44360);
or UO_497 (O_497,N_47837,N_43157);
and UO_498 (O_498,N_48624,N_41756);
xnor UO_499 (O_499,N_45110,N_42530);
nand UO_500 (O_500,N_44354,N_43591);
or UO_501 (O_501,N_41034,N_48477);
nor UO_502 (O_502,N_43477,N_40112);
or UO_503 (O_503,N_41483,N_44683);
nor UO_504 (O_504,N_40170,N_43446);
nand UO_505 (O_505,N_47514,N_48830);
nor UO_506 (O_506,N_48854,N_48987);
nand UO_507 (O_507,N_44489,N_40326);
xnor UO_508 (O_508,N_48946,N_41595);
nor UO_509 (O_509,N_46145,N_43140);
nor UO_510 (O_510,N_49315,N_44702);
nand UO_511 (O_511,N_49930,N_45314);
nor UO_512 (O_512,N_41082,N_41797);
or UO_513 (O_513,N_47498,N_49778);
or UO_514 (O_514,N_42081,N_42835);
nor UO_515 (O_515,N_44673,N_42217);
and UO_516 (O_516,N_41745,N_49318);
nand UO_517 (O_517,N_47050,N_46146);
and UO_518 (O_518,N_44581,N_41705);
nor UO_519 (O_519,N_45750,N_47973);
xor UO_520 (O_520,N_49464,N_43974);
or UO_521 (O_521,N_46553,N_41191);
xor UO_522 (O_522,N_42038,N_45454);
or UO_523 (O_523,N_40436,N_46676);
nor UO_524 (O_524,N_42130,N_45806);
nor UO_525 (O_525,N_46838,N_41194);
nor UO_526 (O_526,N_41924,N_47206);
and UO_527 (O_527,N_41555,N_46448);
nor UO_528 (O_528,N_40934,N_40023);
nand UO_529 (O_529,N_44531,N_48108);
nand UO_530 (O_530,N_43061,N_49342);
and UO_531 (O_531,N_42380,N_43373);
or UO_532 (O_532,N_40721,N_40530);
nor UO_533 (O_533,N_46579,N_49798);
and UO_534 (O_534,N_47055,N_46641);
nand UO_535 (O_535,N_49349,N_49879);
nand UO_536 (O_536,N_46052,N_45732);
and UO_537 (O_537,N_40342,N_42023);
and UO_538 (O_538,N_49259,N_47230);
or UO_539 (O_539,N_49053,N_40367);
and UO_540 (O_540,N_48908,N_43073);
nor UO_541 (O_541,N_40627,N_42024);
nor UO_542 (O_542,N_49294,N_44751);
and UO_543 (O_543,N_40405,N_40563);
xnor UO_544 (O_544,N_40742,N_49097);
and UO_545 (O_545,N_41123,N_47796);
and UO_546 (O_546,N_49877,N_47423);
and UO_547 (O_547,N_40475,N_40718);
nand UO_548 (O_548,N_48539,N_43826);
nand UO_549 (O_549,N_47763,N_42097);
nor UO_550 (O_550,N_48264,N_48069);
nor UO_551 (O_551,N_44996,N_43819);
nand UO_552 (O_552,N_48478,N_43035);
nand UO_553 (O_553,N_40586,N_42576);
xor UO_554 (O_554,N_48795,N_49345);
nor UO_555 (O_555,N_42751,N_40525);
nor UO_556 (O_556,N_43565,N_47095);
or UO_557 (O_557,N_44950,N_45174);
and UO_558 (O_558,N_47930,N_49770);
nor UO_559 (O_559,N_43207,N_45237);
nand UO_560 (O_560,N_41607,N_41505);
xnor UO_561 (O_561,N_47482,N_40376);
and UO_562 (O_562,N_47447,N_43791);
nor UO_563 (O_563,N_45904,N_45486);
or UO_564 (O_564,N_41196,N_47714);
nor UO_565 (O_565,N_44624,N_44102);
nand UO_566 (O_566,N_41100,N_47234);
or UO_567 (O_567,N_43683,N_43112);
nand UO_568 (O_568,N_41633,N_46486);
and UO_569 (O_569,N_42160,N_47413);
nor UO_570 (O_570,N_43917,N_45311);
nor UO_571 (O_571,N_42646,N_44440);
nand UO_572 (O_572,N_40353,N_44595);
and UO_573 (O_573,N_45351,N_46358);
xnor UO_574 (O_574,N_44261,N_43532);
nor UO_575 (O_575,N_45638,N_49194);
nand UO_576 (O_576,N_41364,N_47247);
nor UO_577 (O_577,N_44240,N_49359);
or UO_578 (O_578,N_48759,N_48364);
and UO_579 (O_579,N_41768,N_44572);
or UO_580 (O_580,N_46698,N_48750);
and UO_581 (O_581,N_45468,N_46496);
nor UO_582 (O_582,N_49428,N_48464);
nor UO_583 (O_583,N_41722,N_45445);
nand UO_584 (O_584,N_47671,N_43890);
nand UO_585 (O_585,N_47358,N_42512);
nor UO_586 (O_586,N_41382,N_41375);
nand UO_587 (O_587,N_48455,N_48730);
nor UO_588 (O_588,N_42396,N_43671);
xnor UO_589 (O_589,N_46161,N_45709);
nor UO_590 (O_590,N_49631,N_48952);
nor UO_591 (O_591,N_46030,N_46848);
or UO_592 (O_592,N_46276,N_47591);
or UO_593 (O_593,N_47960,N_44195);
and UO_594 (O_594,N_42051,N_41743);
and UO_595 (O_595,N_49849,N_42972);
or UO_596 (O_596,N_47484,N_41177);
nor UO_597 (O_597,N_43508,N_48228);
nor UO_598 (O_598,N_43896,N_40724);
nand UO_599 (O_599,N_45726,N_43479);
nor UO_600 (O_600,N_46086,N_46287);
xor UO_601 (O_601,N_43782,N_48998);
and UO_602 (O_602,N_49196,N_48483);
nor UO_603 (O_603,N_43966,N_45843);
or UO_604 (O_604,N_40700,N_49901);
and UO_605 (O_605,N_42193,N_46435);
or UO_606 (O_606,N_42289,N_41587);
nand UO_607 (O_607,N_42163,N_45158);
or UO_608 (O_608,N_45546,N_41155);
and UO_609 (O_609,N_45106,N_44148);
and UO_610 (O_610,N_48535,N_41973);
and UO_611 (O_611,N_44662,N_45128);
nor UO_612 (O_612,N_41650,N_49869);
or UO_613 (O_613,N_43520,N_47558);
xor UO_614 (O_614,N_41340,N_41937);
nor UO_615 (O_615,N_44064,N_44181);
nor UO_616 (O_616,N_43390,N_49996);
and UO_617 (O_617,N_45090,N_49881);
or UO_618 (O_618,N_48532,N_48181);
and UO_619 (O_619,N_43469,N_41197);
or UO_620 (O_620,N_42858,N_43717);
and UO_621 (O_621,N_43854,N_40321);
or UO_622 (O_622,N_40549,N_44364);
nor UO_623 (O_623,N_47345,N_41988);
xor UO_624 (O_624,N_43274,N_44499);
nor UO_625 (O_625,N_48855,N_43243);
nand UO_626 (O_626,N_44470,N_42564);
or UO_627 (O_627,N_41496,N_43252);
and UO_628 (O_628,N_44688,N_41406);
or UO_629 (O_629,N_48569,N_44848);
nor UO_630 (O_630,N_41592,N_48438);
or UO_631 (O_631,N_43262,N_45376);
and UO_632 (O_632,N_41072,N_41517);
or UO_633 (O_633,N_41614,N_47638);
nand UO_634 (O_634,N_43696,N_48401);
or UO_635 (O_635,N_46345,N_49829);
or UO_636 (O_636,N_47384,N_48279);
nor UO_637 (O_637,N_40698,N_48212);
or UO_638 (O_638,N_46762,N_41295);
and UO_639 (O_639,N_45368,N_49845);
xnor UO_640 (O_640,N_40780,N_44990);
nand UO_641 (O_641,N_41502,N_45811);
or UO_642 (O_642,N_44451,N_48142);
or UO_643 (O_643,N_42803,N_45383);
nor UO_644 (O_644,N_40716,N_46948);
nand UO_645 (O_645,N_47697,N_46015);
and UO_646 (O_646,N_44821,N_46174);
nand UO_647 (O_647,N_48560,N_42485);
nor UO_648 (O_648,N_45792,N_43726);
nand UO_649 (O_649,N_43832,N_42281);
xnor UO_650 (O_650,N_41111,N_48377);
nor UO_651 (O_651,N_45016,N_40670);
or UO_652 (O_652,N_49130,N_44319);
and UO_653 (O_653,N_49512,N_47953);
nor UO_654 (O_654,N_48111,N_43042);
or UO_655 (O_655,N_46725,N_42926);
or UO_656 (O_656,N_42207,N_49399);
nor UO_657 (O_657,N_48794,N_47356);
nor UO_658 (O_658,N_48099,N_45242);
or UO_659 (O_659,N_40312,N_40993);
nand UO_660 (O_660,N_43602,N_42360);
or UO_661 (O_661,N_46809,N_48351);
and UO_662 (O_662,N_49455,N_47491);
or UO_663 (O_663,N_45933,N_43358);
and UO_664 (O_664,N_46295,N_45052);
nand UO_665 (O_665,N_47803,N_45591);
or UO_666 (O_666,N_49391,N_45039);
nand UO_667 (O_667,N_40319,N_40804);
xor UO_668 (O_668,N_48550,N_48308);
nand UO_669 (O_669,N_43745,N_45157);
nand UO_670 (O_670,N_48075,N_40951);
xor UO_671 (O_671,N_46418,N_47240);
xor UO_672 (O_672,N_45644,N_49466);
or UO_673 (O_673,N_40286,N_46746);
or UO_674 (O_674,N_45135,N_48549);
or UO_675 (O_675,N_48199,N_40630);
or UO_676 (O_676,N_44365,N_41949);
nand UO_677 (O_677,N_40348,N_43327);
and UO_678 (O_678,N_42482,N_44666);
nand UO_679 (O_679,N_49109,N_45077);
nand UO_680 (O_680,N_47030,N_49997);
and UO_681 (O_681,N_46344,N_40479);
and UO_682 (O_682,N_42816,N_48323);
nand UO_683 (O_683,N_40297,N_44389);
or UO_684 (O_684,N_45984,N_44243);
nand UO_685 (O_685,N_45846,N_49472);
or UO_686 (O_686,N_40199,N_46343);
and UO_687 (O_687,N_48474,N_49827);
nor UO_688 (O_688,N_48512,N_44902);
and UO_689 (O_689,N_49431,N_47287);
nand UO_690 (O_690,N_48409,N_43919);
or UO_691 (O_691,N_40815,N_49889);
or UO_692 (O_692,N_45510,N_45381);
xnor UO_693 (O_693,N_41507,N_44380);
xor UO_694 (O_694,N_45277,N_43736);
or UO_695 (O_695,N_48881,N_45328);
nor UO_696 (O_696,N_41048,N_46396);
or UO_697 (O_697,N_49462,N_42370);
nand UO_698 (O_698,N_49883,N_40891);
nor UO_699 (O_699,N_46036,N_41465);
xnor UO_700 (O_700,N_49192,N_42900);
or UO_701 (O_701,N_48522,N_41322);
xor UO_702 (O_702,N_48632,N_45875);
xnor UO_703 (O_703,N_40218,N_47092);
and UO_704 (O_704,N_42303,N_45423);
or UO_705 (O_705,N_42510,N_47522);
xnor UO_706 (O_706,N_43812,N_41074);
nand UO_707 (O_707,N_41397,N_44067);
or UO_708 (O_708,N_47628,N_42084);
nor UO_709 (O_709,N_47777,N_40831);
and UO_710 (O_710,N_44356,N_43012);
or UO_711 (O_711,N_42814,N_46028);
or UO_712 (O_712,N_43770,N_40277);
or UO_713 (O_713,N_43464,N_42250);
or UO_714 (O_714,N_40763,N_49152);
nor UO_715 (O_715,N_44967,N_43955);
and UO_716 (O_716,N_48711,N_41571);
nor UO_717 (O_717,N_45926,N_46118);
nor UO_718 (O_718,N_43078,N_42722);
and UO_719 (O_719,N_46191,N_45809);
xnor UO_720 (O_720,N_48576,N_48900);
nand UO_721 (O_721,N_42740,N_40483);
and UO_722 (O_722,N_42559,N_41600);
or UO_723 (O_723,N_40228,N_43223);
and UO_724 (O_724,N_40338,N_46180);
nor UO_725 (O_725,N_46467,N_47251);
and UO_726 (O_726,N_41874,N_47937);
nor UO_727 (O_727,N_41701,N_41125);
and UO_728 (O_728,N_45553,N_48913);
xor UO_729 (O_729,N_40081,N_49167);
or UO_730 (O_730,N_46115,N_44660);
and UO_731 (O_731,N_42085,N_43945);
nor UO_732 (O_732,N_48566,N_42436);
and UO_733 (O_733,N_49321,N_48083);
nor UO_734 (O_734,N_45582,N_43558);
nor UO_735 (O_735,N_44543,N_46322);
and UO_736 (O_736,N_47512,N_43820);
or UO_737 (O_737,N_49802,N_44051);
and UO_738 (O_738,N_42957,N_40196);
and UO_739 (O_739,N_46749,N_48454);
xnor UO_740 (O_740,N_48134,N_45754);
nand UO_741 (O_741,N_40143,N_40555);
nor UO_742 (O_742,N_40684,N_42548);
nand UO_743 (O_743,N_41649,N_48726);
or UO_744 (O_744,N_41064,N_46352);
or UO_745 (O_745,N_47332,N_46568);
or UO_746 (O_746,N_48331,N_46545);
and UO_747 (O_747,N_46329,N_45142);
and UO_748 (O_748,N_43335,N_40289);
nand UO_749 (O_749,N_46774,N_42515);
nor UO_750 (O_750,N_49895,N_42099);
or UO_751 (O_751,N_42708,N_44806);
or UO_752 (O_752,N_42563,N_44153);
and UO_753 (O_753,N_45393,N_44435);
nand UO_754 (O_754,N_48982,N_44434);
nor UO_755 (O_755,N_42152,N_46949);
nand UO_756 (O_756,N_48035,N_48206);
nand UO_757 (O_757,N_48103,N_43105);
nor UO_758 (O_758,N_49419,N_43789);
and UO_759 (O_759,N_45449,N_43729);
nor UO_760 (O_760,N_42155,N_49229);
xor UO_761 (O_761,N_48488,N_49021);
nor UO_762 (O_762,N_45696,N_49187);
and UO_763 (O_763,N_42421,N_46378);
and UO_764 (O_764,N_44039,N_41116);
nor UO_765 (O_765,N_48634,N_49680);
nand UO_766 (O_766,N_47675,N_49445);
and UO_767 (O_767,N_45814,N_42106);
xor UO_768 (O_768,N_44415,N_44915);
and UO_769 (O_769,N_41945,N_49069);
and UO_770 (O_770,N_47300,N_45741);
nand UO_771 (O_771,N_46469,N_43399);
xnor UO_772 (O_772,N_43272,N_46139);
nor UO_773 (O_773,N_43781,N_43395);
or UO_774 (O_774,N_43859,N_40449);
nor UO_775 (O_775,N_48085,N_45253);
nand UO_776 (O_776,N_40744,N_47457);
nor UO_777 (O_777,N_42267,N_42236);
nand UO_778 (O_778,N_42213,N_42527);
nand UO_779 (O_779,N_46833,N_46783);
and UO_780 (O_780,N_44351,N_45308);
or UO_781 (O_781,N_48250,N_47903);
xor UO_782 (O_782,N_49800,N_43332);
nand UO_783 (O_783,N_49618,N_41629);
or UO_784 (O_784,N_48865,N_40771);
nand UO_785 (O_785,N_40972,N_43963);
xor UO_786 (O_786,N_48198,N_48905);
nand UO_787 (O_787,N_47808,N_49356);
xor UO_788 (O_788,N_45405,N_46849);
nand UO_789 (O_789,N_42443,N_48352);
and UO_790 (O_790,N_42371,N_43744);
and UO_791 (O_791,N_41485,N_40705);
nor UO_792 (O_792,N_48020,N_49447);
and UO_793 (O_793,N_41950,N_49208);
nor UO_794 (O_794,N_41336,N_48140);
and UO_795 (O_795,N_47327,N_45494);
nor UO_796 (O_796,N_41033,N_43454);
or UO_797 (O_797,N_40696,N_46955);
and UO_798 (O_798,N_45865,N_48909);
or UO_799 (O_799,N_49344,N_45444);
nor UO_800 (O_800,N_48050,N_46389);
nand UO_801 (O_801,N_49101,N_46256);
nand UO_802 (O_802,N_48173,N_48049);
and UO_803 (O_803,N_45894,N_42815);
nor UO_804 (O_804,N_42039,N_49134);
or UO_805 (O_805,N_44094,N_41358);
nor UO_806 (O_806,N_49216,N_43590);
nor UO_807 (O_807,N_41712,N_49699);
and UO_808 (O_808,N_41374,N_43077);
xor UO_809 (O_809,N_45249,N_48147);
xor UO_810 (O_810,N_43707,N_49806);
xnor UO_811 (O_811,N_43283,N_49367);
nor UO_812 (O_812,N_43290,N_48660);
nor UO_813 (O_813,N_47097,N_40650);
xnor UO_814 (O_814,N_45872,N_42605);
or UO_815 (O_815,N_41942,N_43652);
and UO_816 (O_816,N_46816,N_42311);
or UO_817 (O_817,N_49482,N_43762);
or UO_818 (O_818,N_47412,N_48840);
xnor UO_819 (O_819,N_47253,N_49644);
nor UO_820 (O_820,N_46307,N_48087);
or UO_821 (O_821,N_41966,N_48702);
nand UO_822 (O_822,N_47664,N_47307);
or UO_823 (O_823,N_41117,N_44262);
and UO_824 (O_824,N_49371,N_41882);
nor UO_825 (O_825,N_42921,N_44007);
or UO_826 (O_826,N_47733,N_44483);
nor UO_827 (O_827,N_45438,N_41410);
nand UO_828 (O_828,N_40172,N_41096);
and UO_829 (O_829,N_40144,N_41218);
or UO_830 (O_830,N_41325,N_46957);
xnor UO_831 (O_831,N_42487,N_44631);
or UO_832 (O_832,N_45075,N_46494);
nand UO_833 (O_833,N_45370,N_43457);
nor UO_834 (O_834,N_49170,N_46501);
or UO_835 (O_835,N_48417,N_46546);
nand UO_836 (O_836,N_44566,N_45262);
xor UO_837 (O_837,N_48609,N_47441);
xor UO_838 (O_838,N_48540,N_41911);
xnor UO_839 (O_839,N_47269,N_48246);
nor UO_840 (O_840,N_48745,N_45074);
nand UO_841 (O_841,N_49769,N_40773);
nor UO_842 (O_842,N_42293,N_49337);
or UO_843 (O_843,N_40635,N_47146);
and UO_844 (O_844,N_45416,N_46645);
nand UO_845 (O_845,N_45973,N_48556);
and UO_846 (O_846,N_45954,N_49886);
nor UO_847 (O_847,N_48253,N_44946);
and UO_848 (O_848,N_49205,N_44053);
nand UO_849 (O_849,N_49076,N_41700);
nor UO_850 (O_850,N_41078,N_46988);
or UO_851 (O_851,N_41800,N_43111);
nor UO_852 (O_852,N_42773,N_45357);
or UO_853 (O_853,N_47177,N_40078);
nor UO_854 (O_854,N_46323,N_41784);
or UO_855 (O_855,N_47754,N_44568);
or UO_856 (O_856,N_41437,N_46293);
nor UO_857 (O_857,N_43485,N_45710);
nor UO_858 (O_858,N_40053,N_41870);
nor UO_859 (O_859,N_40636,N_44638);
and UO_860 (O_860,N_43099,N_41287);
or UO_861 (O_861,N_45527,N_42239);
nor UO_862 (O_862,N_46043,N_48880);
xnor UO_863 (O_863,N_41589,N_49727);
nand UO_864 (O_864,N_46969,N_48200);
and UO_865 (O_865,N_49786,N_41467);
or UO_866 (O_866,N_40757,N_40560);
nor UO_867 (O_867,N_48394,N_46571);
nor UO_868 (O_868,N_49228,N_40511);
nand UO_869 (O_869,N_40315,N_46088);
and UO_870 (O_870,N_49518,N_42242);
nor UO_871 (O_871,N_49514,N_49923);
or UO_872 (O_872,N_44079,N_47741);
and UO_873 (O_873,N_47147,N_40545);
nor UO_874 (O_874,N_40104,N_42066);
nor UO_875 (O_875,N_48806,N_40503);
nand UO_876 (O_876,N_46639,N_40608);
nand UO_877 (O_877,N_48594,N_47407);
nor UO_878 (O_878,N_41887,N_47058);
nand UO_879 (O_879,N_42971,N_40565);
or UO_880 (O_880,N_45168,N_41414);
nand UO_881 (O_881,N_40008,N_44883);
nor UO_882 (O_882,N_46947,N_48425);
nor UO_883 (O_883,N_47351,N_43504);
nor UO_884 (O_884,N_40135,N_44501);
and UO_885 (O_885,N_43774,N_44010);
and UO_886 (O_886,N_44330,N_45509);
nor UO_887 (O_887,N_47330,N_47132);
nand UO_888 (O_888,N_47849,N_42190);
xor UO_889 (O_889,N_45492,N_48722);
nor UO_890 (O_890,N_43254,N_40554);
nor UO_891 (O_891,N_47800,N_47784);
nor UO_892 (O_892,N_49920,N_49049);
nand UO_893 (O_893,N_42028,N_49086);
nand UO_894 (O_894,N_40453,N_48462);
nand UO_895 (O_895,N_47859,N_44340);
or UO_896 (O_896,N_43482,N_42729);
and UO_897 (O_897,N_42129,N_40388);
nand UO_898 (O_898,N_41110,N_44317);
nor UO_899 (O_899,N_41347,N_49252);
nand UO_900 (O_900,N_49148,N_46158);
xor UO_901 (O_901,N_42444,N_49890);
and UO_902 (O_902,N_41147,N_42092);
and UO_903 (O_903,N_41696,N_48370);
or UO_904 (O_904,N_46632,N_46927);
or UO_905 (O_905,N_45420,N_46918);
nand UO_906 (O_906,N_49034,N_46743);
or UO_907 (O_907,N_46537,N_46274);
nand UO_908 (O_908,N_42821,N_48994);
nand UO_909 (O_909,N_43392,N_48252);
nand UO_910 (O_910,N_48898,N_48499);
nor UO_911 (O_911,N_40770,N_46914);
xnor UO_912 (O_912,N_49015,N_45712);
and UO_913 (O_913,N_44035,N_40607);
or UO_914 (O_914,N_40802,N_44854);
nor UO_915 (O_915,N_46059,N_43097);
or UO_916 (O_916,N_49404,N_45120);
and UO_917 (O_917,N_47756,N_48010);
or UO_918 (O_918,N_42481,N_44378);
xor UO_919 (O_919,N_43356,N_40208);
nor UO_920 (O_920,N_45259,N_44237);
nor UO_921 (O_921,N_42930,N_41501);
nor UO_922 (O_922,N_43992,N_43768);
or UO_923 (O_923,N_43689,N_41639);
nor UO_924 (O_924,N_42433,N_43090);
nor UO_925 (O_925,N_47631,N_49368);
nand UO_926 (O_926,N_41736,N_40992);
nand UO_927 (O_927,N_45994,N_46945);
or UO_928 (O_928,N_40671,N_41820);
and UO_929 (O_929,N_44315,N_40661);
and UO_930 (O_930,N_49429,N_46596);
nor UO_931 (O_931,N_46650,N_44477);
and UO_932 (O_932,N_42504,N_47436);
nand UO_933 (O_933,N_42219,N_44246);
nand UO_934 (O_934,N_42961,N_49394);
or UO_935 (O_935,N_48468,N_42599);
nand UO_936 (O_936,N_41810,N_46420);
or UO_937 (O_937,N_42007,N_48014);
or UO_938 (O_938,N_49870,N_44108);
and UO_939 (O_939,N_45022,N_40485);
nor UO_940 (O_940,N_48521,N_47416);
nand UO_941 (O_941,N_41112,N_40068);
or UO_942 (O_942,N_49390,N_45676);
nor UO_943 (O_943,N_48154,N_47847);
or UO_944 (O_944,N_45278,N_40969);
nor UO_945 (O_945,N_40561,N_47382);
xor UO_946 (O_946,N_45791,N_42671);
nand UO_947 (O_947,N_47174,N_46505);
xor UO_948 (O_948,N_46044,N_46772);
nor UO_949 (O_949,N_47694,N_48211);
nor UO_950 (O_950,N_46349,N_44311);
nand UO_951 (O_951,N_46884,N_44866);
nand UO_952 (O_952,N_46453,N_41690);
nor UO_953 (O_953,N_44264,N_41735);
and UO_954 (O_954,N_43611,N_47089);
nand UO_955 (O_955,N_44532,N_45176);
nor UO_956 (O_956,N_45296,N_44594);
or UO_957 (O_957,N_49833,N_40728);
or UO_958 (O_958,N_43210,N_41693);
and UO_959 (O_959,N_48021,N_45751);
nor UO_960 (O_960,N_42414,N_49861);
or UO_961 (O_961,N_48680,N_40454);
or UO_962 (O_962,N_43365,N_44820);
nor UO_963 (O_963,N_44471,N_45963);
nand UO_964 (O_964,N_42491,N_41249);
and UO_965 (O_965,N_44943,N_45945);
xor UO_966 (O_966,N_44439,N_40964);
nor UO_967 (O_967,N_49959,N_42864);
nand UO_968 (O_968,N_45331,N_48864);
nand UO_969 (O_969,N_41300,N_40169);
nor UO_970 (O_970,N_48727,N_47067);
or UO_971 (O_971,N_43705,N_45067);
and UO_972 (O_972,N_40430,N_40562);
or UO_973 (O_973,N_47311,N_45611);
and UO_974 (O_974,N_47133,N_46907);
or UO_975 (O_975,N_45589,N_49169);
xnor UO_976 (O_976,N_46165,N_49146);
nor UO_977 (O_977,N_43926,N_45488);
and UO_978 (O_978,N_45216,N_40687);
nand UO_979 (O_979,N_41936,N_46341);
or UO_980 (O_980,N_49556,N_49120);
nand UO_981 (O_981,N_42666,N_47746);
nand UO_982 (O_982,N_47357,N_41863);
nor UO_983 (O_983,N_44835,N_42974);
nor UO_984 (O_984,N_40335,N_43879);
xnor UO_985 (O_985,N_45282,N_48631);
nor UO_986 (O_986,N_48408,N_44370);
and UO_987 (O_987,N_49144,N_42727);
or UO_988 (O_988,N_45068,N_45519);
and UO_989 (O_989,N_41470,N_48541);
nand UO_990 (O_990,N_42540,N_46720);
nand UO_991 (O_991,N_44145,N_44668);
or UO_992 (O_992,N_44685,N_42199);
xor UO_993 (O_993,N_41920,N_42261);
and UO_994 (O_994,N_40155,N_40400);
and UO_995 (O_995,N_42946,N_42775);
nand UO_996 (O_996,N_44644,N_46119);
and UO_997 (O_997,N_47315,N_43163);
and UO_998 (O_998,N_41527,N_40480);
nand UO_999 (O_999,N_40304,N_44127);
nand UO_1000 (O_1000,N_43658,N_46861);
nand UO_1001 (O_1001,N_45524,N_47561);
nor UO_1002 (O_1002,N_40825,N_41104);
nand UO_1003 (O_1003,N_48857,N_40789);
nand UO_1004 (O_1004,N_44442,N_49776);
and UO_1005 (O_1005,N_46799,N_42076);
nor UO_1006 (O_1006,N_49763,N_41190);
or UO_1007 (O_1007,N_43814,N_42966);
or UO_1008 (O_1008,N_45482,N_48395);
and UO_1009 (O_1009,N_48586,N_43694);
and UO_1010 (O_1010,N_49787,N_41698);
nor UO_1011 (O_1011,N_42459,N_48822);
or UO_1012 (O_1012,N_49108,N_46905);
and UO_1013 (O_1013,N_41952,N_49212);
or UO_1014 (O_1014,N_44105,N_49524);
nor UO_1015 (O_1015,N_45733,N_48307);
nand UO_1016 (O_1016,N_47517,N_46271);
nor UO_1017 (O_1017,N_41368,N_45635);
xor UO_1018 (O_1018,N_44612,N_41666);
nand UO_1019 (O_1019,N_49758,N_44390);
nor UO_1020 (O_1020,N_44918,N_41794);
nand UO_1021 (O_1021,N_41439,N_43153);
xor UO_1022 (O_1022,N_47304,N_44591);
or UO_1023 (O_1023,N_45024,N_41363);
and UO_1024 (O_1024,N_41839,N_41430);
xnor UO_1025 (O_1025,N_48995,N_47866);
nor UO_1026 (O_1026,N_45162,N_48452);
and UO_1027 (O_1027,N_41737,N_42766);
or UO_1028 (O_1028,N_44379,N_47853);
and UO_1029 (O_1029,N_44023,N_40459);
nand UO_1030 (O_1030,N_43434,N_46210);
nor UO_1031 (O_1031,N_42779,N_43018);
or UO_1032 (O_1032,N_45943,N_44728);
or UO_1033 (O_1033,N_43211,N_44174);
xnor UO_1034 (O_1034,N_40381,N_41580);
and UO_1035 (O_1035,N_47744,N_42285);
nand UO_1036 (O_1036,N_41760,N_46380);
and UO_1037 (O_1037,N_43187,N_47961);
xor UO_1038 (O_1038,N_49446,N_49378);
nand UO_1039 (O_1039,N_41426,N_45062);
or UO_1040 (O_1040,N_40779,N_44628);
nand UO_1041 (O_1041,N_47312,N_48313);
xnor UO_1042 (O_1042,N_42931,N_40298);
nor UO_1043 (O_1043,N_43491,N_45202);
and UO_1044 (O_1044,N_42776,N_46634);
or UO_1045 (O_1045,N_41301,N_42417);
nor UO_1046 (O_1046,N_47901,N_42252);
nand UO_1047 (O_1047,N_42376,N_41385);
nor UO_1048 (O_1048,N_47171,N_42300);
nand UO_1049 (O_1049,N_41842,N_48471);
nand UO_1050 (O_1050,N_47117,N_48066);
nor UO_1051 (O_1051,N_44941,N_49911);
or UO_1052 (O_1052,N_45736,N_45525);
or UO_1053 (O_1053,N_40269,N_40387);
nand UO_1054 (O_1054,N_49573,N_49181);
nand UO_1055 (O_1055,N_49582,N_42278);
xor UO_1056 (O_1056,N_44504,N_45417);
nor UO_1057 (O_1057,N_41010,N_43247);
xor UO_1058 (O_1058,N_44763,N_40535);
nor UO_1059 (O_1059,N_40861,N_46100);
nand UO_1060 (O_1060,N_42790,N_46530);
and UO_1061 (O_1061,N_45547,N_40187);
nor UO_1062 (O_1062,N_42356,N_47259);
or UO_1063 (O_1063,N_44749,N_49589);
or UO_1064 (O_1064,N_41400,N_46612);
xnor UO_1065 (O_1065,N_41267,N_45867);
nor UO_1066 (O_1066,N_46408,N_46410);
nor UO_1067 (O_1067,N_44815,N_42362);
nor UO_1068 (O_1068,N_44191,N_44190);
and UO_1069 (O_1069,N_40077,N_44700);
nand UO_1070 (O_1070,N_47712,N_45573);
nor UO_1071 (O_1071,N_41098,N_43141);
nor UO_1072 (O_1072,N_43559,N_41509);
nor UO_1073 (O_1073,N_47986,N_45231);
and UO_1074 (O_1074,N_44560,N_45979);
or UO_1075 (O_1075,N_49379,N_44175);
nor UO_1076 (O_1076,N_41270,N_45651);
nor UO_1077 (O_1077,N_47467,N_48319);
or UO_1078 (O_1078,N_45181,N_40739);
nand UO_1079 (O_1079,N_45272,N_45336);
and UO_1080 (O_1080,N_40116,N_45578);
nand UO_1081 (O_1081,N_49178,N_44057);
or UO_1082 (O_1082,N_48627,N_43906);
xnor UO_1083 (O_1083,N_47768,N_45091);
and UO_1084 (O_1084,N_44114,N_48416);
and UO_1085 (O_1085,N_48508,N_43780);
and UO_1086 (O_1086,N_47231,N_40866);
nand UO_1087 (O_1087,N_45784,N_45215);
xor UO_1088 (O_1088,N_46240,N_48263);
nand UO_1089 (O_1089,N_40611,N_41747);
nor UO_1090 (O_1090,N_44028,N_47091);
nand UO_1091 (O_1091,N_46597,N_41298);
nand UO_1092 (O_1092,N_46671,N_41153);
nor UO_1093 (O_1093,N_47855,N_42031);
xor UO_1094 (O_1094,N_49480,N_45538);
and UO_1095 (O_1095,N_49454,N_46714);
xnor UO_1096 (O_1096,N_47218,N_49489);
or UO_1097 (O_1097,N_48733,N_45443);
nand UO_1098 (O_1098,N_45797,N_45666);
and UO_1099 (O_1099,N_46536,N_43545);
and UO_1100 (O_1100,N_46864,N_43288);
nand UO_1101 (O_1101,N_45042,N_43401);
nor UO_1102 (O_1102,N_45285,N_47488);
and UO_1103 (O_1103,N_49941,N_49314);
nor UO_1104 (O_1104,N_49329,N_40145);
xor UO_1105 (O_1105,N_44610,N_41575);
and UO_1106 (O_1106,N_41304,N_42150);
or UO_1107 (O_1107,N_48879,N_49597);
nor UO_1108 (O_1108,N_40224,N_47180);
nand UO_1109 (O_1109,N_46973,N_44387);
nor UO_1110 (O_1110,N_47344,N_45257);
and UO_1111 (O_1111,N_42041,N_46524);
nand UO_1112 (O_1112,N_42290,N_44215);
nor UO_1113 (O_1113,N_43133,N_45145);
nor UO_1114 (O_1114,N_48244,N_41898);
nand UO_1115 (O_1115,N_40995,N_44277);
and UO_1116 (O_1116,N_49405,N_41922);
or UO_1117 (O_1117,N_49738,N_47822);
nand UO_1118 (O_1118,N_42916,N_40089);
and UO_1119 (O_1119,N_40191,N_41256);
and UO_1120 (O_1120,N_41324,N_46076);
nor UO_1121 (O_1121,N_46157,N_46667);
nand UO_1122 (O_1122,N_44476,N_45831);
and UO_1123 (O_1123,N_42368,N_40013);
nand UO_1124 (O_1124,N_48558,N_46306);
nand UO_1125 (O_1125,N_47154,N_49666);
and UO_1126 (O_1126,N_40878,N_46635);
or UO_1127 (O_1127,N_44140,N_44523);
nand UO_1128 (O_1128,N_46261,N_44944);
or UO_1129 (O_1129,N_47570,N_40881);
nand UO_1130 (O_1130,N_49463,N_42739);
nand UO_1131 (O_1131,N_41462,N_41982);
and UO_1132 (O_1132,N_42082,N_41020);
and UO_1133 (O_1133,N_40351,N_40356);
or UO_1134 (O_1134,N_45853,N_49760);
nand UO_1135 (O_1135,N_44087,N_49884);
and UO_1136 (O_1136,N_48148,N_49840);
or UO_1137 (O_1137,N_44622,N_42892);
or UO_1138 (O_1138,N_44221,N_45500);
nor UO_1139 (O_1139,N_46715,N_45321);
nor UO_1140 (O_1140,N_41415,N_43730);
nand UO_1141 (O_1141,N_49843,N_47707);
xnor UO_1142 (O_1142,N_40614,N_41004);
and UO_1143 (O_1143,N_48350,N_40212);
nor UO_1144 (O_1144,N_42868,N_46078);
nand UO_1145 (O_1145,N_47289,N_46744);
nor UO_1146 (O_1146,N_47446,N_49658);
nor UO_1147 (O_1147,N_49090,N_46980);
nor UO_1148 (O_1148,N_48931,N_46019);
xor UO_1149 (O_1149,N_42040,N_43197);
nand UO_1150 (O_1150,N_49479,N_48662);
and UO_1151 (O_1151,N_45115,N_41672);
nand UO_1152 (O_1152,N_46492,N_41543);
xnor UO_1153 (O_1153,N_49590,N_41740);
nor UO_1154 (O_1154,N_40807,N_43261);
or UO_1155 (O_1155,N_47128,N_49295);
nand UO_1156 (O_1156,N_43150,N_46561);
nor UO_1157 (O_1157,N_40769,N_41658);
and UO_1158 (O_1158,N_48801,N_45640);
and UO_1159 (O_1159,N_49547,N_46892);
or UO_1160 (O_1160,N_48078,N_45185);
or UO_1161 (O_1161,N_49312,N_44827);
nand UO_1162 (O_1162,N_41627,N_48232);
nand UO_1163 (O_1163,N_40233,N_40727);
nand UO_1164 (O_1164,N_45620,N_40841);
xor UO_1165 (O_1165,N_40413,N_45001);
or UO_1166 (O_1166,N_46476,N_43725);
nor UO_1167 (O_1167,N_47923,N_42716);
nand UO_1168 (O_1168,N_43869,N_43060);
or UO_1169 (O_1169,N_48741,N_43114);
xnor UO_1170 (O_1170,N_49860,N_49442);
xor UO_1171 (O_1171,N_48432,N_47835);
nor UO_1172 (O_1172,N_47523,N_45281);
nor UO_1173 (O_1173,N_41931,N_43511);
nand UO_1174 (O_1174,N_45602,N_48993);
or UO_1175 (O_1175,N_47303,N_42893);
or UO_1176 (O_1176,N_48763,N_45063);
or UO_1177 (O_1177,N_42582,N_47108);
nor UO_1178 (O_1178,N_44227,N_46887);
xor UO_1179 (O_1179,N_49052,N_40785);
nor UO_1180 (O_1180,N_49546,N_44424);
nor UO_1181 (O_1181,N_48381,N_49790);
or UO_1182 (O_1182,N_40153,N_45690);
or UO_1183 (O_1183,N_49133,N_43741);
nor UO_1184 (O_1184,N_43667,N_45248);
and UO_1185 (O_1185,N_49938,N_41908);
nor UO_1186 (O_1186,N_47650,N_45467);
nor UO_1187 (O_1187,N_48436,N_47942);
nand UO_1188 (O_1188,N_47787,N_43606);
nor UO_1189 (O_1189,N_45923,N_47188);
nand UO_1190 (O_1190,N_48874,N_42440);
nand UO_1191 (O_1191,N_47987,N_42430);
nor UO_1192 (O_1192,N_44086,N_49719);
nor UO_1193 (O_1193,N_46013,N_45665);
or UO_1194 (O_1194,N_41179,N_42113);
or UO_1195 (O_1195,N_42295,N_40264);
and UO_1196 (O_1196,N_41195,N_46051);
or UO_1197 (O_1197,N_46845,N_43104);
and UO_1198 (O_1198,N_49855,N_46282);
nor UO_1199 (O_1199,N_49586,N_48363);
and UO_1200 (O_1200,N_47971,N_41824);
nor UO_1201 (O_1201,N_45895,N_45126);
xor UO_1202 (O_1202,N_40564,N_46643);
or UO_1203 (O_1203,N_49811,N_42567);
or UO_1204 (O_1204,N_41965,N_48773);
or UO_1205 (O_1205,N_44881,N_40027);
and UO_1206 (O_1206,N_48245,N_48567);
nor UO_1207 (O_1207,N_42102,N_40029);
nor UO_1208 (O_1208,N_49240,N_42237);
and UO_1209 (O_1209,N_41283,N_49199);
nor UO_1210 (O_1210,N_44173,N_44366);
nand UO_1211 (O_1211,N_49932,N_42143);
nor UO_1212 (O_1212,N_44268,N_42407);
and UO_1213 (O_1213,N_42297,N_44210);
nor UO_1214 (O_1214,N_46882,N_46796);
xor UO_1215 (O_1215,N_40271,N_42953);
nor UO_1216 (O_1216,N_47149,N_41551);
or UO_1217 (O_1217,N_43579,N_49799);
and UO_1218 (O_1218,N_42182,N_42826);
or UO_1219 (O_1219,N_42901,N_45992);
nor UO_1220 (O_1220,N_49862,N_43716);
nor UO_1221 (O_1221,N_49504,N_47005);
nand UO_1222 (O_1222,N_41808,N_42463);
or UO_1223 (O_1223,N_49561,N_44756);
nand UO_1224 (O_1224,N_49826,N_42951);
xor UO_1225 (O_1225,N_44643,N_47825);
nand UO_1226 (O_1226,N_42655,N_40229);
nor UO_1227 (O_1227,N_43816,N_40977);
xnor UO_1228 (O_1228,N_41957,N_49365);
and UO_1229 (O_1229,N_41061,N_46222);
or UO_1230 (O_1230,N_44995,N_46818);
xnor UO_1231 (O_1231,N_48106,N_41318);
or UO_1232 (O_1232,N_45883,N_41261);
and UO_1233 (O_1233,N_48190,N_46771);
and UO_1234 (O_1234,N_45540,N_46626);
or UO_1235 (O_1235,N_49537,N_45526);
nand UO_1236 (O_1236,N_44025,N_47911);
nand UO_1237 (O_1237,N_45725,N_47639);
nand UO_1238 (O_1238,N_42804,N_44176);
or UO_1239 (O_1239,N_43238,N_42664);
nand UO_1240 (O_1240,N_41925,N_41974);
nand UO_1241 (O_1241,N_43425,N_47209);
nand UO_1242 (O_1242,N_48677,N_48772);
or UO_1243 (O_1243,N_42709,N_43034);
nand UO_1244 (O_1244,N_42735,N_46869);
and UO_1245 (O_1245,N_40175,N_48983);
or UO_1246 (O_1246,N_49452,N_44474);
xor UO_1247 (O_1247,N_44759,N_40034);
and UO_1248 (O_1248,N_45399,N_42660);
nor UO_1249 (O_1249,N_41958,N_40438);
and UO_1250 (O_1250,N_48461,N_41339);
nand UO_1251 (O_1251,N_41822,N_44805);
nand UO_1252 (O_1252,N_42327,N_43958);
xor UO_1253 (O_1253,N_42056,N_44506);
nor UO_1254 (O_1254,N_40301,N_47420);
and UO_1255 (O_1255,N_47526,N_46266);
and UO_1256 (O_1256,N_48355,N_43615);
nand UO_1257 (O_1257,N_48170,N_41697);
nor UO_1258 (O_1258,N_44649,N_48046);
xnor UO_1259 (O_1259,N_47350,N_48189);
nand UO_1260 (O_1260,N_47082,N_41495);
nor UO_1261 (O_1261,N_48182,N_41849);
nor UO_1262 (O_1262,N_49226,N_45375);
and UO_1263 (O_1263,N_49303,N_48872);
xnor UO_1264 (O_1264,N_43137,N_40818);
or UO_1265 (O_1265,N_48128,N_48875);
or UO_1266 (O_1266,N_43201,N_41099);
xnor UO_1267 (O_1267,N_44665,N_47511);
and UO_1268 (O_1268,N_40652,N_49782);
and UO_1269 (O_1269,N_40292,N_41224);
nor UO_1270 (O_1270,N_47263,N_47192);
or UO_1271 (O_1271,N_45220,N_41590);
nand UO_1272 (O_1272,N_43589,N_48422);
nor UO_1273 (O_1273,N_45224,N_41688);
and UO_1274 (O_1274,N_41630,N_42094);
nor UO_1275 (O_1275,N_40149,N_45485);
or UO_1276 (O_1276,N_48129,N_49741);
and UO_1277 (O_1277,N_46961,N_47074);
nor UO_1278 (O_1278,N_45433,N_42348);
nand UO_1279 (O_1279,N_40283,N_48607);
and UO_1280 (O_1280,N_49511,N_45108);
nand UO_1281 (O_1281,N_46588,N_45190);
nor UO_1282 (O_1282,N_47143,N_44133);
nand UO_1283 (O_1283,N_45002,N_43976);
nand UO_1284 (O_1284,N_43651,N_45749);
nor UO_1285 (O_1285,N_49348,N_43024);
nor UO_1286 (O_1286,N_40912,N_41054);
nor UO_1287 (O_1287,N_46813,N_48379);
xnor UO_1288 (O_1288,N_48876,N_44359);
xnor UO_1289 (O_1289,N_47550,N_46141);
nor UO_1290 (O_1290,N_46912,N_40533);
and UO_1291 (O_1291,N_49985,N_46862);
or UO_1292 (O_1292,N_43732,N_45554);
or UO_1293 (O_1293,N_45152,N_44252);
nor UO_1294 (O_1294,N_40656,N_41259);
xor UO_1295 (O_1295,N_42534,N_40819);
nand UO_1296 (O_1296,N_48925,N_47465);
nor UO_1297 (O_1297,N_45820,N_46328);
and UO_1298 (O_1298,N_49010,N_43250);
nor UO_1299 (O_1299,N_40986,N_41909);
nor UO_1300 (O_1300,N_48042,N_46193);
and UO_1301 (O_1301,N_45250,N_41273);
and UO_1302 (O_1302,N_42227,N_40898);
nand UO_1303 (O_1303,N_40402,N_49114);
nand UO_1304 (O_1304,N_49675,N_47319);
and UO_1305 (O_1305,N_49522,N_46583);
or UO_1306 (O_1306,N_44147,N_46936);
and UO_1307 (O_1307,N_47977,N_47186);
and UO_1308 (O_1308,N_44582,N_43884);
nor UO_1309 (O_1309,N_41367,N_47509);
or UO_1310 (O_1310,N_43253,N_40219);
nand UO_1311 (O_1311,N_42746,N_42358);
nand UO_1312 (O_1312,N_48843,N_45544);
nand UO_1313 (O_1313,N_45936,N_42373);
or UO_1314 (O_1314,N_43899,N_44333);
or UO_1315 (O_1315,N_41221,N_40842);
nor UO_1316 (O_1316,N_44496,N_47260);
and UO_1317 (O_1317,N_40431,N_49781);
nand UO_1318 (O_1318,N_48338,N_45922);
nor UO_1319 (O_1319,N_42114,N_42086);
nand UO_1320 (O_1320,N_48039,N_47485);
and UO_1321 (O_1321,N_43314,N_48317);
nor UO_1322 (O_1322,N_46310,N_47602);
nor UO_1323 (O_1323,N_47607,N_42480);
or UO_1324 (O_1324,N_44701,N_41085);
and UO_1325 (O_1325,N_49341,N_40708);
or UO_1326 (O_1326,N_41890,N_42596);
and UO_1327 (O_1327,N_46104,N_44570);
nor UO_1328 (O_1328,N_46320,N_46330);
or UO_1329 (O_1329,N_40830,N_40967);
nand UO_1330 (O_1330,N_46611,N_43971);
or UO_1331 (O_1331,N_45119,N_40055);
xnor UO_1332 (O_1332,N_45018,N_43010);
nor UO_1333 (O_1333,N_45678,N_42503);
nor UO_1334 (O_1334,N_45319,N_40765);
nor UO_1335 (O_1335,N_40678,N_46258);
or UO_1336 (O_1336,N_44851,N_45869);
nor UO_1337 (O_1337,N_46752,N_42895);
nand UO_1338 (O_1338,N_45094,N_43541);
nor UO_1339 (O_1339,N_43465,N_48060);
xor UO_1340 (O_1340,N_42620,N_47990);
nand UO_1341 (O_1341,N_46785,N_48639);
nor UO_1342 (O_1342,N_40579,N_44137);
or UO_1343 (O_1343,N_45737,N_43481);
and UO_1344 (O_1344,N_45430,N_42501);
nand UO_1345 (O_1345,N_46455,N_43510);
nand UO_1346 (O_1346,N_43172,N_48183);
xor UO_1347 (O_1347,N_42446,N_43580);
or UO_1348 (O_1348,N_45209,N_44283);
and UO_1349 (O_1349,N_49957,N_47736);
nor UO_1350 (O_1350,N_45288,N_47836);
nor UO_1351 (O_1351,N_44238,N_48450);
nand UO_1352 (O_1352,N_47817,N_46313);
nor UO_1353 (O_1353,N_49661,N_43810);
or UO_1354 (O_1354,N_40706,N_41167);
and UO_1355 (O_1355,N_49980,N_43876);
nor UO_1356 (O_1356,N_45636,N_42203);
nand UO_1357 (O_1357,N_48026,N_43384);
or UO_1358 (O_1358,N_42976,N_46919);
nand UO_1359 (O_1359,N_47046,N_40360);
or UO_1360 (O_1360,N_48235,N_44625);
or UO_1361 (O_1361,N_45503,N_43075);
nor UO_1362 (O_1362,N_44469,N_45461);
or UO_1363 (O_1363,N_48888,N_41578);
nor UO_1364 (O_1364,N_46620,N_41231);
nor UO_1365 (O_1365,N_49868,N_45506);
nor UO_1366 (O_1366,N_44955,N_46560);
nand UO_1367 (O_1367,N_46642,N_48739);
nand UO_1368 (O_1368,N_42461,N_43938);
nor UO_1369 (O_1369,N_41763,N_40146);
xnor UO_1370 (O_1370,N_45320,N_45909);
xnor UO_1371 (O_1371,N_41185,N_43988);
nand UO_1372 (O_1372,N_44722,N_47914);
nand UO_1373 (O_1373,N_46422,N_46181);
nor UO_1374 (O_1374,N_41567,N_42118);
xnor UO_1375 (O_1375,N_47025,N_41334);
nor UO_1376 (O_1376,N_40484,N_47073);
nor UO_1377 (O_1377,N_40491,N_47086);
or UO_1378 (O_1378,N_48769,N_40692);
xnor UO_1379 (O_1379,N_42088,N_49565);
or UO_1380 (O_1380,N_40888,N_47780);
nand UO_1381 (O_1381,N_45752,N_40422);
nor UO_1382 (O_1382,N_49916,N_47161);
xor UO_1383 (O_1383,N_49707,N_41867);
nor UO_1384 (O_1384,N_47298,N_47759);
or UO_1385 (O_1385,N_45403,N_41436);
nand UO_1386 (O_1386,N_48695,N_43525);
and UO_1387 (O_1387,N_49629,N_40643);
and UO_1388 (O_1388,N_48233,N_43116);
nor UO_1389 (O_1389,N_41836,N_46648);
or UO_1390 (O_1390,N_48287,N_46173);
or UO_1391 (O_1391,N_42521,N_41651);
and UO_1392 (O_1392,N_48775,N_42372);
or UO_1393 (O_1393,N_40128,N_44192);
and UO_1394 (O_1394,N_43865,N_44065);
nand UO_1395 (O_1395,N_40916,N_46251);
and UO_1396 (O_1396,N_48340,N_42876);
or UO_1397 (O_1397,N_40539,N_48268);
nor UO_1398 (O_1398,N_49568,N_43285);
or UO_1399 (O_1399,N_42782,N_40694);
xor UO_1400 (O_1400,N_44812,N_48063);
or UO_1401 (O_1401,N_43677,N_47220);
and UO_1402 (O_1402,N_49388,N_43766);
or UO_1403 (O_1403,N_49087,N_43870);
or UO_1404 (O_1404,N_41620,N_46211);
nor UO_1405 (O_1405,N_40846,N_40573);
nor UO_1406 (O_1406,N_48878,N_48492);
nor UO_1407 (O_1407,N_44571,N_43013);
and UO_1408 (O_1408,N_45876,N_43623);
xnor UO_1409 (O_1409,N_46732,N_40421);
and UO_1410 (O_1410,N_46996,N_44321);
or UO_1411 (O_1411,N_46991,N_43058);
or UO_1412 (O_1412,N_41466,N_41206);
nand UO_1413 (O_1413,N_45916,N_48916);
nor UO_1414 (O_1414,N_49135,N_48703);
nand UO_1415 (O_1415,N_42555,N_44139);
nand UO_1416 (O_1416,N_46254,N_45955);
nor UO_1417 (O_1417,N_48760,N_41812);
and UO_1418 (O_1418,N_40634,N_46940);
nor UO_1419 (O_1419,N_44587,N_44931);
nand UO_1420 (O_1420,N_47994,N_43000);
or UO_1421 (O_1421,N_41021,N_44083);
nor UO_1422 (O_1422,N_42389,N_42673);
nor UO_1423 (O_1423,N_46382,N_43378);
and UO_1424 (O_1424,N_43968,N_44755);
nand UO_1425 (O_1425,N_43943,N_45245);
or UO_1426 (O_1426,N_43713,N_49438);
xnor UO_1427 (O_1427,N_43937,N_42125);
nor UO_1428 (O_1428,N_43750,N_40895);
nand UO_1429 (O_1429,N_48276,N_41331);
or UO_1430 (O_1430,N_47189,N_46788);
or UO_1431 (O_1431,N_45304,N_41411);
and UO_1432 (O_1432,N_46246,N_44550);
nand UO_1433 (O_1433,N_49910,N_45395);
nand UO_1434 (O_1434,N_46490,N_43845);
xnor UO_1435 (O_1435,N_43230,N_46464);
nand UO_1436 (O_1436,N_43977,N_45140);
or UO_1437 (O_1437,N_49046,N_44443);
nand UO_1438 (O_1438,N_48853,N_49245);
nand UO_1439 (O_1439,N_41833,N_42853);
and UO_1440 (O_1440,N_46278,N_48999);
and UO_1441 (O_1441,N_47812,N_42854);
and UO_1442 (O_1442,N_45845,N_44493);
nor UO_1443 (O_1443,N_43302,N_42812);
or UO_1444 (O_1444,N_45100,N_47339);
or UO_1445 (O_1445,N_45874,N_46249);
and UO_1446 (O_1446,N_42787,N_42856);
and UO_1447 (O_1447,N_41741,N_44589);
and UO_1448 (O_1448,N_40948,N_43006);
or UO_1449 (O_1449,N_41653,N_44284);
xnor UO_1450 (O_1450,N_45824,N_44774);
and UO_1451 (O_1451,N_40379,N_44534);
nor UO_1452 (O_1452,N_41219,N_40546);
and UO_1453 (O_1453,N_48169,N_41635);
or UO_1454 (O_1454,N_40944,N_47439);
or UO_1455 (O_1455,N_46929,N_44111);
or UO_1456 (O_1456,N_46804,N_45627);
nor UO_1457 (O_1457,N_41713,N_41761);
nor UO_1458 (O_1458,N_41449,N_47113);
nor UO_1459 (O_1459,N_46227,N_41305);
and UO_1460 (O_1460,N_48115,N_40048);
nand UO_1461 (O_1461,N_40743,N_49083);
nand UO_1462 (O_1462,N_46817,N_47015);
and UO_1463 (O_1463,N_47492,N_44275);
or UO_1464 (O_1464,N_44164,N_48672);
nand UO_1465 (O_1465,N_43300,N_42744);
nand UO_1466 (O_1466,N_42522,N_44299);
or UO_1467 (O_1467,N_40275,N_49569);
or UO_1468 (O_1468,N_47951,N_44562);
nand UO_1469 (O_1469,N_40666,N_42750);
nor UO_1470 (O_1470,N_42323,N_41661);
nor UO_1471 (O_1471,N_41659,N_44600);
nand UO_1472 (O_1472,N_46814,N_48633);
nand UO_1473 (O_1473,N_49155,N_46402);
nand UO_1474 (O_1474,N_42745,N_48842);
and UO_1475 (O_1475,N_45703,N_46944);
or UO_1476 (O_1476,N_45793,N_41398);
or UO_1477 (O_1477,N_45340,N_43025);
or UO_1478 (O_1478,N_49954,N_40336);
and UO_1479 (O_1479,N_47116,N_43842);
nor UO_1480 (O_1480,N_41148,N_44430);
or UO_1481 (O_1481,N_47692,N_46779);
nand UO_1482 (O_1482,N_40540,N_44916);
xor UO_1483 (O_1483,N_48312,N_43260);
and UO_1484 (O_1484,N_46079,N_45826);
or UO_1485 (O_1485,N_47865,N_41885);
or UO_1486 (O_1486,N_42719,N_41991);
nor UO_1487 (O_1487,N_40618,N_42653);
nor UO_1488 (O_1488,N_42221,N_43323);
nor UO_1489 (O_1489,N_42764,N_41731);
or UO_1490 (O_1490,N_42309,N_41790);
nor UO_1491 (O_1491,N_48767,N_46304);
xnor UO_1492 (O_1492,N_48884,N_47551);
xnor UO_1493 (O_1493,N_43232,N_42101);
or UO_1494 (O_1494,N_46614,N_45014);
and UO_1495 (O_1495,N_45758,N_40150);
or UO_1496 (O_1496,N_41238,N_41044);
and UO_1497 (O_1497,N_47033,N_42774);
xor UO_1498 (O_1498,N_44002,N_42016);
or UO_1499 (O_1499,N_42195,N_45175);
or UO_1500 (O_1500,N_41748,N_42550);
nand UO_1501 (O_1501,N_43233,N_45536);
and UO_1502 (O_1502,N_44458,N_49640);
nand UO_1503 (O_1503,N_47101,N_42060);
nand UO_1504 (O_1504,N_45072,N_41835);
xnor UO_1505 (O_1505,N_47398,N_46674);
xor UO_1506 (O_1506,N_46523,N_40762);
nor UO_1507 (O_1507,N_48585,N_45655);
and UO_1508 (O_1508,N_44623,N_44152);
nor UO_1509 (O_1509,N_40623,N_42592);
nor UO_1510 (O_1510,N_48867,N_43863);
or UO_1511 (O_1511,N_40211,N_42785);
nor UO_1512 (O_1512,N_42057,N_46565);
and UO_1513 (O_1513,N_42255,N_40848);
or UO_1514 (O_1514,N_41040,N_44329);
or UO_1515 (O_1515,N_42544,N_40063);
or UO_1516 (O_1516,N_48052,N_40913);
nand UO_1517 (O_1517,N_44708,N_40215);
xor UO_1518 (O_1518,N_49943,N_48008);
nand UO_1519 (O_1519,N_42712,N_46708);
nand UO_1520 (O_1520,N_49671,N_48136);
and UO_1521 (O_1521,N_41841,N_47689);
or UO_1522 (O_1522,N_46716,N_49176);
nand UO_1523 (O_1523,N_46239,N_45134);
nor UO_1524 (O_1524,N_42590,N_47396);
and UO_1525 (O_1525,N_48316,N_40299);
and UO_1526 (O_1526,N_40704,N_41222);
nand UO_1527 (O_1527,N_48667,N_41819);
nor UO_1528 (O_1528,N_48518,N_41780);
or UO_1529 (O_1529,N_48045,N_48737);
xor UO_1530 (O_1530,N_45965,N_41799);
nor UO_1531 (O_1531,N_40473,N_46499);
or UO_1532 (O_1532,N_44205,N_46495);
nor UO_1533 (O_1533,N_49981,N_45695);
nor UO_1534 (O_1534,N_43455,N_49268);
nor UO_1535 (O_1535,N_43239,N_45144);
or UO_1536 (O_1536,N_48685,N_44402);
and UO_1537 (O_1537,N_49465,N_41214);
and UO_1538 (O_1538,N_40429,N_41769);
and UO_1539 (O_1539,N_47397,N_41895);
nor UO_1540 (O_1540,N_44958,N_42233);
nand UO_1541 (O_1541,N_48177,N_44172);
xor UO_1542 (O_1542,N_49698,N_48893);
nand UO_1543 (O_1543,N_45424,N_45830);
or UO_1544 (O_1544,N_48957,N_43307);
or UO_1545 (O_1545,N_46021,N_48162);
or UO_1546 (O_1546,N_47017,N_46335);
xnor UO_1547 (O_1547,N_48724,N_47453);
or UO_1548 (O_1548,N_49654,N_43329);
or UO_1549 (O_1549,N_47437,N_40152);
nand UO_1550 (O_1550,N_49847,N_44166);
or UO_1551 (O_1551,N_48265,N_47003);
or UO_1552 (O_1552,N_49937,N_44841);
nand UO_1553 (O_1553,N_46113,N_44059);
nand UO_1554 (O_1554,N_44982,N_46171);
nand UO_1555 (O_1555,N_46392,N_42831);
nor UO_1556 (O_1556,N_48638,N_42115);
and UO_1557 (O_1557,N_41750,N_47466);
nor UO_1558 (O_1558,N_42867,N_43495);
or UO_1559 (O_1559,N_45297,N_42850);
nor UO_1560 (O_1560,N_49363,N_43184);
and UO_1561 (O_1561,N_43551,N_42792);
nor UO_1562 (O_1562,N_41405,N_40120);
nand UO_1563 (O_1563,N_44952,N_45474);
nand UO_1564 (O_1564,N_43142,N_49287);
nand UO_1565 (O_1565,N_42598,N_40648);
or UO_1566 (O_1566,N_42829,N_47616);
and UO_1567 (O_1567,N_41641,N_43647);
nand UO_1568 (O_1568,N_47077,N_45036);
nor UO_1569 (O_1569,N_44316,N_47156);
or UO_1570 (O_1570,N_47622,N_48131);
xor UO_1571 (O_1571,N_43478,N_40330);
nand UO_1572 (O_1572,N_41851,N_47474);
and UO_1573 (O_1573,N_45708,N_45878);
nor UO_1574 (O_1574,N_40097,N_45082);
nand UO_1575 (O_1575,N_41561,N_44406);
and UO_1576 (O_1576,N_40067,N_44936);
or UO_1577 (O_1577,N_41418,N_47363);
or UO_1578 (O_1578,N_45531,N_47797);
and UO_1579 (O_1579,N_46072,N_40745);
or UO_1580 (O_1580,N_48533,N_46234);
or UO_1581 (O_1581,N_47199,N_43269);
nor UO_1582 (O_1582,N_41403,N_45702);
or UO_1583 (O_1583,N_43162,N_41513);
nor UO_1584 (O_1584,N_42243,N_45968);
and UO_1585 (O_1585,N_44393,N_46701);
nor UO_1586 (O_1586,N_40538,N_48496);
and UO_1587 (O_1587,N_42889,N_44729);
and UO_1588 (O_1588,N_44962,N_46515);
xnor UO_1589 (O_1589,N_46516,N_49519);
nand UO_1590 (O_1590,N_49912,N_49753);
or UO_1591 (O_1591,N_44278,N_48816);
nand UO_1592 (O_1592,N_44868,N_41528);
and UO_1593 (O_1593,N_42449,N_44225);
nor UO_1594 (O_1594,N_49585,N_40674);
and UO_1595 (O_1595,N_47048,N_47131);
and UO_1596 (O_1596,N_47701,N_45911);
and UO_1597 (O_1597,N_49441,N_44197);
and UO_1598 (O_1598,N_44537,N_45155);
nor UO_1599 (O_1599,N_46846,N_43598);
and UO_1600 (O_1600,N_48172,N_48951);
nor UO_1601 (O_1601,N_49516,N_40882);
and UO_1602 (O_1602,N_40209,N_46077);
or UO_1603 (O_1603,N_41482,N_41023);
nor UO_1604 (O_1604,N_44012,N_46965);
or UO_1605 (O_1605,N_44428,N_44449);
nand UO_1606 (O_1606,N_44336,N_45789);
xor UO_1607 (O_1607,N_48161,N_49035);
and UO_1608 (O_1608,N_40510,N_45234);
or UO_1609 (O_1609,N_45804,N_45309);
nand UO_1610 (O_1610,N_41573,N_40599);
and UO_1611 (O_1611,N_48573,N_48501);
or UO_1612 (O_1612,N_42205,N_44131);
or UO_1613 (O_1613,N_43851,N_41714);
nor UO_1614 (O_1614,N_48195,N_40824);
or UO_1615 (O_1615,N_44045,N_44720);
and UO_1616 (O_1616,N_44917,N_46777);
or UO_1617 (O_1617,N_43161,N_49433);
or UO_1618 (O_1618,N_43803,N_49250);
nor UO_1619 (O_1619,N_47630,N_44482);
or UO_1620 (O_1620,N_42507,N_44909);
nor UO_1621 (O_1621,N_44919,N_42478);
nand UO_1622 (O_1622,N_42684,N_46633);
and UO_1623 (O_1623,N_44177,N_46531);
xor UO_1624 (O_1624,N_46318,N_40262);
nand UO_1625 (O_1625,N_45410,N_49952);
xnor UO_1626 (O_1626,N_43056,N_44198);
nand UO_1627 (O_1627,N_46729,N_46830);
nor UO_1628 (O_1628,N_46430,N_42668);
nand UO_1629 (O_1629,N_41943,N_43411);
xnor UO_1630 (O_1630,N_48654,N_43818);
or UO_1631 (O_1631,N_47624,N_45812);
nor UO_1632 (O_1632,N_47022,N_48514);
or UO_1633 (O_1633,N_49968,N_45003);
or UO_1634 (O_1634,N_48341,N_46150);
and UO_1635 (O_1635,N_41785,N_46450);
nor UO_1636 (O_1636,N_45274,N_49351);
or UO_1637 (O_1637,N_45574,N_47645);
nor UO_1638 (O_1638,N_48259,N_47318);
nand UO_1639 (O_1639,N_42793,N_45458);
or UO_1640 (O_1640,N_42960,N_47828);
and UO_1641 (O_1641,N_45947,N_42457);
or UO_1642 (O_1642,N_41046,N_47976);
or UO_1643 (O_1643,N_49509,N_49499);
nor UO_1644 (O_1644,N_46825,N_41782);
nor UO_1645 (O_1645,N_47115,N_41500);
xnor UO_1646 (O_1646,N_49435,N_47227);
nor UO_1647 (O_1647,N_46279,N_49612);
or UO_1648 (O_1648,N_45848,N_41665);
nand UO_1649 (O_1649,N_44392,N_47893);
nor UO_1650 (O_1650,N_47038,N_45017);
and UO_1651 (O_1651,N_41409,N_44548);
or UO_1652 (O_1652,N_47941,N_45971);
nor UO_1653 (O_1653,N_42069,N_42711);
or UO_1654 (O_1654,N_46231,N_49197);
or UO_1655 (O_1655,N_41647,N_44460);
or UO_1656 (O_1656,N_46835,N_47719);
xor UO_1657 (O_1657,N_44834,N_43664);
and UO_1658 (O_1658,N_48296,N_45603);
nor UO_1659 (O_1659,N_48421,N_43304);
or UO_1660 (O_1660,N_43957,N_41559);
nor UO_1661 (O_1661,N_44983,N_43053);
nand UO_1662 (O_1662,N_47010,N_49383);
nand UO_1663 (O_1663,N_44089,N_42488);
or UO_1664 (O_1664,N_43530,N_44689);
or UO_1665 (O_1665,N_45799,N_44690);
and UO_1666 (O_1666,N_43369,N_47203);
nor UO_1667 (O_1667,N_40962,N_43241);
or UO_1668 (O_1668,N_41092,N_45359);
and UO_1669 (O_1669,N_46756,N_43216);
or UO_1670 (O_1670,N_46092,N_43975);
and UO_1671 (O_1671,N_46361,N_44768);
xnor UO_1672 (O_1672,N_42532,N_46228);
or UO_1673 (O_1673,N_46793,N_40406);
or UO_1674 (O_1674,N_47197,N_40843);
nor UO_1675 (O_1675,N_48500,N_45463);
nand UO_1676 (O_1676,N_44485,N_44157);
nand UO_1677 (O_1677,N_43155,N_49838);
nor UO_1678 (O_1678,N_49125,N_45386);
xnor UO_1679 (O_1679,N_44754,N_44642);
nand UO_1680 (O_1680,N_45711,N_47964);
nor UO_1681 (O_1681,N_46863,N_49600);
nor UO_1682 (O_1682,N_42637,N_43666);
xnor UO_1683 (O_1683,N_42944,N_46177);
and UO_1684 (O_1684,N_49414,N_46012);
nand UO_1685 (O_1685,N_40646,N_49871);
nand UO_1686 (O_1686,N_43471,N_46275);
nor UO_1687 (O_1687,N_43218,N_49595);
and UO_1688 (O_1688,N_45633,N_40633);
and UO_1689 (O_1689,N_43610,N_43786);
nand UO_1690 (O_1690,N_48714,N_45906);
and UO_1691 (O_1691,N_41791,N_45866);
nor UO_1692 (O_1692,N_40553,N_41557);
nand UO_1693 (O_1693,N_45829,N_43123);
nand UO_1694 (O_1694,N_47580,N_45472);
and UO_1695 (O_1695,N_40349,N_40354);
or UO_1696 (O_1696,N_46074,N_49487);
and UO_1697 (O_1697,N_48580,N_43772);
nand UO_1698 (O_1698,N_40243,N_49067);
or UO_1699 (O_1699,N_43470,N_48030);
nor UO_1700 (O_1700,N_41556,N_43970);
xnor UO_1701 (O_1701,N_42514,N_43719);
and UO_1702 (O_1702,N_43553,N_45777);
and UO_1703 (O_1703,N_45015,N_43191);
and UO_1704 (O_1704,N_45679,N_44658);
or UO_1705 (O_1705,N_42319,N_40798);
xor UO_1706 (O_1706,N_40827,N_42796);
nand UO_1707 (O_1707,N_49756,N_43552);
nand UO_1708 (O_1708,N_40070,N_49535);
xor UO_1709 (O_1709,N_45771,N_41548);
and UO_1710 (O_1710,N_47233,N_49635);
nand UO_1711 (O_1711,N_43492,N_44716);
nand UO_1712 (O_1712,N_40787,N_43412);
xor UO_1713 (O_1713,N_46458,N_43174);
nand UO_1714 (O_1714,N_44891,N_43049);
or UO_1715 (O_1715,N_45982,N_41369);
nor UO_1716 (O_1716,N_46901,N_47411);
or UO_1717 (O_1717,N_41230,N_44250);
nor UO_1718 (O_1718,N_48226,N_43334);
and UO_1719 (O_1719,N_49234,N_43687);
nand UO_1720 (O_1720,N_43326,N_46201);
or UO_1721 (O_1721,N_44875,N_42095);
xor UO_1722 (O_1722,N_40239,N_44017);
or UO_1723 (O_1723,N_49887,N_48783);
nor UO_1724 (O_1724,N_45687,N_48729);
xnor UO_1725 (O_1725,N_48373,N_45223);
or UO_1726 (O_1726,N_46401,N_43621);
and UO_1727 (O_1727,N_40493,N_42810);
xnor UO_1728 (O_1728,N_42208,N_43856);
nor UO_1729 (O_1729,N_48282,N_42923);
nand UO_1730 (O_1730,N_42231,N_46114);
nand UO_1731 (O_1731,N_45089,N_47651);
nor UO_1732 (O_1732,N_46192,N_47085);
and UO_1733 (O_1733,N_41323,N_48793);
nor UO_1734 (O_1734,N_45096,N_46637);
and UO_1735 (O_1735,N_42860,N_47313);
or UO_1736 (O_1736,N_47381,N_47892);
nor UO_1737 (O_1737,N_44529,N_44664);
or UO_1738 (O_1738,N_45267,N_40361);
and UO_1739 (O_1739,N_49242,N_44030);
or UO_1740 (O_1740,N_40729,N_45849);
nor UO_1741 (O_1741,N_49267,N_43212);
nand UO_1742 (O_1742,N_44472,N_45088);
nand UO_1743 (O_1743,N_48996,N_47811);
nor UO_1744 (O_1744,N_41715,N_46471);
xor UO_1745 (O_1745,N_43405,N_47406);
nor UO_1746 (O_1746,N_42304,N_44527);
and UO_1747 (O_1747,N_42049,N_47364);
and UO_1748 (O_1748,N_48110,N_47785);
nand UO_1749 (O_1749,N_47641,N_41009);
nor UO_1750 (O_1750,N_41417,N_45341);
nor UO_1751 (O_1751,N_46085,N_43778);
or UO_1752 (O_1752,N_45079,N_40752);
nor UO_1753 (O_1753,N_49935,N_44129);
nand UO_1754 (O_1754,N_40223,N_42934);
and UO_1755 (O_1755,N_41547,N_45493);
nor UO_1756 (O_1756,N_46298,N_44136);
nor UO_1757 (O_1757,N_48334,N_43452);
xnor UO_1758 (O_1758,N_40257,N_49338);
nor UO_1759 (O_1759,N_43458,N_46457);
nand UO_1760 (O_1760,N_40282,N_45575);
nor UO_1761 (O_1761,N_41097,N_49139);
and UO_1762 (O_1762,N_44288,N_48568);
or UO_1763 (O_1763,N_42560,N_46592);
nand UO_1764 (O_1764,N_43066,N_46462);
nor UO_1765 (O_1765,N_46528,N_44558);
xnor UO_1766 (O_1766,N_44447,N_43368);
nor UO_1767 (O_1767,N_43263,N_43497);
nor UO_1768 (O_1768,N_42538,N_45746);
and UO_1769 (O_1769,N_43564,N_41071);
or UO_1770 (O_1770,N_49102,N_43336);
nor UO_1771 (O_1771,N_40751,N_48774);
and UO_1772 (O_1772,N_41568,N_44769);
and UO_1773 (O_1773,N_42247,N_44849);
nand UO_1774 (O_1774,N_46555,N_43978);
nand UO_1775 (O_1775,N_43921,N_44948);
or UO_1776 (O_1776,N_44052,N_44966);
nand UO_1777 (O_1777,N_48036,N_47816);
or UO_1778 (O_1778,N_48663,N_45379);
nor UO_1779 (O_1779,N_41868,N_46011);
nand UO_1780 (O_1780,N_42575,N_42986);
nand UO_1781 (O_1781,N_42761,N_42736);
and UO_1782 (O_1782,N_40965,N_42100);
and UO_1783 (O_1783,N_41431,N_41095);
nor UO_1784 (O_1784,N_47938,N_47537);
or UO_1785 (O_1785,N_49803,N_47889);
and UO_1786 (O_1786,N_46197,N_49732);
nor UO_1787 (O_1787,N_42394,N_46188);
nor UO_1788 (O_1788,N_46934,N_46731);
nor UO_1789 (O_1789,N_47799,N_44003);
and UO_1790 (O_1790,N_45692,N_41972);
nand UO_1791 (O_1791,N_47690,N_43215);
nand UO_1792 (O_1792,N_45628,N_44542);
and UO_1793 (O_1793,N_47081,N_49172);
or UO_1794 (O_1794,N_49437,N_40331);
nand UO_1795 (O_1795,N_48033,N_40167);
and UO_1796 (O_1796,N_43771,N_45183);
nor UO_1797 (O_1797,N_48166,N_43346);
and UO_1798 (O_1798,N_45738,N_46018);
or UO_1799 (O_1799,N_43370,N_47072);
nor UO_1800 (O_1800,N_42805,N_44536);
xnor UO_1801 (O_1801,N_43840,N_47329);
or UO_1802 (O_1802,N_46218,N_43387);
nor UO_1803 (O_1803,N_46035,N_40946);
nor UO_1804 (O_1804,N_47278,N_47385);
nand UO_1805 (O_1805,N_45284,N_40512);
nand UO_1806 (O_1806,N_45757,N_44584);
nor UO_1807 (O_1807,N_41217,N_48326);
nand UO_1808 (O_1808,N_43605,N_46878);
and UO_1809 (O_1809,N_46398,N_47673);
nor UO_1810 (O_1810,N_43410,N_45899);
and UO_1811 (O_1811,N_47475,N_47824);
nor UO_1812 (O_1812,N_48684,N_40125);
nand UO_1813 (O_1813,N_44223,N_43151);
or UO_1814 (O_1814,N_46391,N_44830);
nand UO_1815 (O_1815,N_46602,N_49100);
nor UO_1816 (O_1816,N_44229,N_43783);
and UO_1817 (O_1817,N_45498,N_43480);
nor UO_1818 (O_1818,N_41638,N_46194);
nand UO_1819 (O_1819,N_42506,N_47533);
nand UO_1820 (O_1820,N_44155,N_41520);
and UO_1821 (O_1821,N_41976,N_43240);
and UO_1822 (O_1822,N_45030,N_45301);
nand UO_1823 (O_1823,N_43418,N_49839);
nand UO_1824 (O_1824,N_42517,N_49677);
nor UO_1825 (O_1825,N_48734,N_49532);
nand UO_1826 (O_1826,N_43106,N_47895);
nand UO_1827 (O_1827,N_41591,N_43074);
nand UO_1828 (O_1828,N_42928,N_45373);
or UO_1829 (O_1829,N_40140,N_46730);
and UO_1830 (O_1830,N_49486,N_45770);
xnor UO_1831 (O_1831,N_44425,N_46976);
and UO_1832 (O_1832,N_40740,N_45783);
xor UO_1833 (O_1833,N_49496,N_42078);
and UO_1834 (O_1834,N_41243,N_41644);
nor UO_1835 (O_1835,N_49248,N_45905);
or UO_1836 (O_1836,N_49856,N_41234);
nor UO_1837 (O_1837,N_43159,N_44816);
nor UO_1838 (O_1838,N_41656,N_42585);
xor UO_1839 (O_1839,N_47772,N_42606);
or UO_1840 (O_1840,N_40207,N_46727);
and UO_1841 (O_1841,N_45408,N_40025);
nor UO_1842 (O_1842,N_46580,N_43316);
or UO_1843 (O_1843,N_47496,N_47589);
nand UO_1844 (O_1844,N_45005,N_46176);
nand UO_1845 (O_1845,N_49817,N_44287);
nand UO_1846 (O_1846,N_42869,N_45165);
or UO_1847 (O_1847,N_43032,N_41873);
and UO_1848 (O_1848,N_47208,N_42141);
nand UO_1849 (O_1849,N_45729,N_40147);
or UO_1850 (O_1850,N_44006,N_47982);
nor UO_1851 (O_1851,N_44867,N_41971);
and UO_1852 (O_1852,N_47862,N_47328);
nor UO_1853 (O_1853,N_43833,N_41309);
and UO_1854 (O_1854,N_42927,N_41211);
nand UO_1855 (O_1855,N_41538,N_49506);
and UO_1856 (O_1856,N_41588,N_41282);
xnor UO_1857 (O_1857,N_46484,N_40548);
or UO_1858 (O_1858,N_42083,N_44188);
and UO_1859 (O_1859,N_47606,N_45680);
nor UO_1860 (O_1860,N_42698,N_48589);
nor UO_1861 (O_1861,N_40746,N_41135);
nand UO_1862 (O_1862,N_46091,N_46200);
or UO_1863 (O_1863,N_43076,N_40737);
nand UO_1864 (O_1864,N_49724,N_47403);
and UO_1865 (O_1865,N_41205,N_41934);
or UO_1866 (O_1866,N_44347,N_44773);
nand UO_1867 (O_1867,N_49149,N_44535);
and UO_1868 (O_1868,N_42675,N_40528);
and UO_1869 (O_1869,N_48692,N_40631);
or UO_1870 (O_1870,N_45479,N_44559);
nor UO_1871 (O_1871,N_43221,N_49291);
and UO_1872 (O_1872,N_42556,N_43622);
nand UO_1873 (O_1873,N_41454,N_48275);
and UO_1874 (O_1874,N_40507,N_40050);
nor UO_1875 (O_1875,N_40621,N_41109);
nand UO_1876 (O_1876,N_47751,N_40617);
and UO_1877 (O_1877,N_47838,N_49762);
nor UO_1878 (O_1878,N_48950,N_40509);
and UO_1879 (O_1879,N_40603,N_42448);
and UO_1880 (O_1880,N_41601,N_44888);
and UO_1881 (O_1881,N_46482,N_44627);
nand UO_1882 (O_1882,N_43062,N_47264);
or UO_1883 (O_1883,N_48077,N_46735);
and UO_1884 (O_1884,N_42691,N_46554);
or UO_1885 (O_1885,N_44876,N_47119);
nor UO_1886 (O_1886,N_47788,N_41776);
nand UO_1887 (O_1887,N_40333,N_42266);
and UO_1888 (O_1888,N_42670,N_48899);
nor UO_1889 (O_1889,N_46061,N_42845);
nand UO_1890 (O_1890,N_44134,N_46164);
and UO_1891 (O_1891,N_48151,N_46080);
and UO_1892 (O_1892,N_43306,N_43182);
and UO_1893 (O_1893,N_43877,N_42594);
and UO_1894 (O_1894,N_45707,N_49726);
or UO_1895 (O_1895,N_46987,N_47342);
xor UO_1896 (O_1896,N_42292,N_42685);
nor UO_1897 (O_1897,N_49241,N_49129);
or UO_1898 (O_1898,N_48604,N_41719);
nor UO_1899 (O_1899,N_46599,N_49443);
or UO_1900 (O_1900,N_47275,N_41706);
nand UO_1901 (O_1901,N_47433,N_43408);
nor UO_1902 (O_1902,N_41685,N_48770);
and UO_1903 (O_1903,N_48367,N_43196);
and UO_1904 (O_1904,N_40749,N_47229);
nand UO_1905 (O_1905,N_44826,N_44865);
or UO_1906 (O_1906,N_46658,N_41826);
xor UO_1907 (O_1907,N_48610,N_46058);
nand UO_1908 (O_1908,N_41932,N_45404);
nor UO_1909 (O_1909,N_48217,N_42183);
nand UO_1910 (O_1910,N_44991,N_49701);
or UO_1911 (O_1911,N_47354,N_43790);
xor UO_1912 (O_1912,N_45466,N_46207);
or UO_1913 (O_1913,N_45460,N_49962);
xor UO_1914 (O_1914,N_49971,N_45387);
nor UO_1915 (O_1915,N_41875,N_49678);
nor UO_1916 (O_1916,N_47996,N_47969);
xor UO_1917 (O_1917,N_47026,N_44092);
nor UO_1918 (O_1918,N_43445,N_47418);
nand UO_1919 (O_1919,N_47600,N_46659);
or UO_1920 (O_1920,N_40390,N_43281);
or UO_1921 (O_1921,N_43518,N_44969);
or UO_1922 (O_1922,N_42738,N_44597);
or UO_1923 (O_1923,N_48152,N_48949);
or UO_1924 (O_1924,N_44254,N_48937);
or UO_1925 (O_1925,N_43217,N_47065);
nand UO_1926 (O_1926,N_42791,N_47827);
xor UO_1927 (O_1927,N_46267,N_49070);
nand UO_1928 (O_1928,N_45593,N_48159);
and UO_1929 (O_1929,N_42524,N_49747);
or UO_1930 (O_1930,N_49456,N_42258);
nand UO_1931 (O_1931,N_48835,N_45315);
and UO_1932 (O_1932,N_48270,N_43699);
or UO_1933 (O_1933,N_44399,N_46347);
nand UO_1934 (O_1934,N_42222,N_49574);
and UO_1935 (O_1935,N_47487,N_41796);
nor UO_1936 (O_1936,N_41269,N_41378);
or UO_1937 (O_1937,N_45203,N_40663);
nand UO_1938 (O_1938,N_43908,N_40005);
xnor UO_1939 (O_1939,N_49702,N_41118);
xnor UO_1940 (O_1940,N_40612,N_40417);
or UO_1941 (O_1941,N_49902,N_49392);
nor UO_1942 (O_1942,N_41463,N_45775);
or UO_1943 (O_1943,N_40662,N_43625);
or UO_1944 (O_1944,N_44593,N_49737);
or UO_1945 (O_1945,N_45260,N_41460);
nor UO_1946 (O_1946,N_42367,N_42035);
nand UO_1947 (O_1947,N_46662,N_41626);
xor UO_1948 (O_1948,N_47235,N_44567);
and UO_1949 (O_1949,N_44771,N_43927);
or UO_1950 (O_1950,N_47294,N_49164);
and UO_1951 (O_1951,N_43376,N_45860);
xor UO_1952 (O_1952,N_47024,N_46244);
nor UO_1953 (O_1953,N_44245,N_45520);
nor UO_1954 (O_1954,N_46967,N_45256);
nor UO_1955 (O_1955,N_43008,N_47157);
xnor UO_1956 (O_1956,N_47663,N_40256);
nor UO_1957 (O_1957,N_47730,N_40917);
xnor UO_1958 (O_1958,N_42572,N_46190);
or UO_1959 (O_1959,N_49745,N_48339);
or UO_1960 (O_1960,N_47062,N_42742);
nand UO_1961 (O_1961,N_41739,N_45046);
nor UO_1962 (O_1962,N_46605,N_43256);
nand UO_1963 (O_1963,N_45714,N_42352);
nand UO_1964 (O_1964,N_46954,N_41425);
or UO_1965 (O_1965,N_45361,N_47217);
or UO_1966 (O_1966,N_47916,N_46627);
and UO_1967 (O_1967,N_49247,N_40179);
or UO_1968 (O_1968,N_42003,N_44037);
xor UO_1969 (O_1969,N_46326,N_43882);
nor UO_1970 (O_1970,N_46742,N_42119);
nand UO_1971 (O_1971,N_46444,N_43289);
and UO_1972 (O_1972,N_40852,N_43317);
xor UO_1973 (O_1973,N_48242,N_46172);
or UO_1974 (O_1974,N_40099,N_47660);
nor UO_1975 (O_1975,N_44088,N_45753);
xnor UO_1976 (O_1976,N_42611,N_44792);
nand UO_1977 (O_1977,N_48165,N_49307);
nor UO_1978 (O_1978,N_44459,N_40788);
and UO_1979 (O_1979,N_42844,N_45631);
xnor UO_1980 (O_1980,N_41297,N_41280);
nand UO_1981 (O_1981,N_49526,N_47470);
and UO_1982 (O_1982,N_41314,N_42615);
xnor UO_1983 (O_1983,N_41579,N_40311);
nand UO_1984 (O_1984,N_40796,N_49221);
nand UO_1985 (O_1985,N_44409,N_43737);
nand UO_1986 (O_1986,N_42331,N_41786);
nor UO_1987 (O_1987,N_43194,N_47540);
and UO_1988 (O_1988,N_41083,N_42635);
xor UO_1989 (O_1989,N_48877,N_46649);
nand UO_1990 (O_1990,N_45491,N_49408);
or UO_1991 (O_1991,N_48933,N_43222);
nor UO_1992 (O_1992,N_46776,N_40640);
nor UO_1993 (O_1993,N_43692,N_49147);
or UO_1994 (O_1994,N_45020,N_45236);
nor UO_1995 (O_1995,N_43685,N_42045);
nand UO_1996 (O_1996,N_41350,N_43712);
nand UO_1997 (O_1997,N_45561,N_48445);
or UO_1998 (O_1998,N_40279,N_47236);
xor UO_1999 (O_1999,N_45246,N_48428);
and UO_2000 (O_2000,N_47165,N_45208);
nand UO_2001 (O_2001,N_40163,N_43601);
and UO_2002 (O_2002,N_41027,N_48613);
xnor UO_2003 (O_2003,N_49866,N_47755);
nor UO_2004 (O_2004,N_41237,N_47926);
or UO_2005 (O_2005,N_47370,N_45932);
and UO_2006 (O_2006,N_41080,N_40955);
nand UO_2007 (O_2007,N_41726,N_41989);
or UO_2008 (O_2008,N_47340,N_48234);
or UO_2009 (O_2009,N_45344,N_45305);
or UO_2010 (O_2010,N_47372,N_47151);
or UO_2011 (O_2011,N_44913,N_49717);
xor UO_2012 (O_2012,N_49003,N_43079);
xor UO_2013 (O_2013,N_43148,N_44836);
nor UO_2014 (O_2014,N_47922,N_48676);
or UO_2015 (O_2015,N_41162,N_43490);
and UO_2016 (O_2016,N_43086,N_42220);
nor UO_2017 (O_2017,N_43733,N_43795);
nand UO_2018 (O_2018,N_46538,N_44879);
and UO_2019 (O_2019,N_42151,N_47789);
or UO_2020 (O_2020,N_47842,N_40767);
nor UO_2021 (O_2021,N_49016,N_46562);
nand UO_2022 (O_2022,N_41226,N_49614);
and UO_2023 (O_2023,N_46950,N_43597);
and UO_2024 (O_2024,N_44410,N_48004);
xnor UO_2025 (O_2025,N_48283,N_42171);
nand UO_2026 (O_2026,N_41062,N_48440);
or UO_2027 (O_2027,N_49611,N_41771);
or UO_2028 (O_2028,N_44987,N_46026);
or UO_2029 (O_2029,N_43936,N_46601);
xor UO_2030 (O_2030,N_49508,N_45532);
and UO_2031 (O_2031,N_47869,N_45045);
nand UO_2032 (O_2032,N_42728,N_42749);
and UO_2033 (O_2033,N_40122,N_41215);
or UO_2034 (O_2034,N_48743,N_49386);
and UO_2035 (O_2035,N_42268,N_44169);
or UO_2036 (O_2036,N_40441,N_40308);
nor UO_2037 (O_2037,N_40764,N_44121);
nor UO_2038 (O_2038,N_42833,N_48707);
nand UO_2039 (O_2039,N_41030,N_45080);
nor UO_2040 (O_2040,N_45390,N_40323);
and UO_2041 (O_2041,N_48261,N_42378);
nand UO_2042 (O_2042,N_48405,N_44078);
xnor UO_2043 (O_2043,N_47924,N_40531);
and UO_2044 (O_2044,N_49440,N_41815);
or UO_2045 (O_2045,N_49674,N_49094);
and UO_2046 (O_2046,N_48504,N_46926);
and UO_2047 (O_2047,N_43669,N_45078);
nor UO_2048 (O_2048,N_49400,N_48248);
nand UO_2049 (O_2049,N_46456,N_40395);
or UO_2050 (O_2050,N_41232,N_41613);
nand UO_2051 (O_2051,N_46040,N_44632);
xnor UO_2052 (O_2052,N_49615,N_43844);
and UO_2053 (O_2053,N_44717,N_42135);
or UO_2054 (O_2054,N_45291,N_43537);
nand UO_2055 (O_2055,N_46572,N_47501);
nand UO_2056 (O_2056,N_41146,N_40826);
nand UO_2057 (O_2057,N_45206,N_49755);
and UO_2058 (O_2058,N_41980,N_41412);
nand UO_2059 (O_2059,N_42676,N_46432);
nor UO_2060 (O_2060,N_44253,N_47001);
nand UO_2061 (O_2061,N_49089,N_48100);
nor UO_2062 (O_2062,N_48669,N_43064);
nor UO_2063 (O_2063,N_43681,N_41275);
xor UO_2064 (O_2064,N_48959,N_41204);
and UO_2065 (O_2065,N_48858,N_40550);
nor UO_2066 (O_2066,N_40463,N_42565);
nor UO_2067 (O_2067,N_46068,N_44549);
nor UO_2068 (O_2068,N_40205,N_42915);
nor UO_2069 (O_2069,N_49961,N_47310);
and UO_2070 (O_2070,N_48836,N_47034);
or UO_2071 (O_2071,N_44267,N_42777);
nand UO_2072 (O_2072,N_40747,N_40655);
nor UO_2073 (O_2073,N_44341,N_47846);
or UO_2074 (O_2074,N_40559,N_44125);
nand UO_2075 (O_2075,N_48687,N_43264);
or UO_2076 (O_2076,N_48120,N_40082);
nor UO_2077 (O_2077,N_45563,N_46459);
and UO_2078 (O_2078,N_45489,N_43362);
and UO_2079 (O_2079,N_49396,N_45343);
nand UO_2080 (O_2080,N_43805,N_41550);
nand UO_2081 (O_2081,N_49578,N_48406);
nor UO_2082 (O_2082,N_49820,N_48542);
or UO_2083 (O_2083,N_45131,N_46355);
xor UO_2084 (O_2084,N_45766,N_42000);
nor UO_2085 (O_2085,N_42962,N_47039);
nor UO_2086 (O_2086,N_49274,N_47422);
nand UO_2087 (O_2087,N_41175,N_40945);
nor UO_2088 (O_2088,N_42374,N_45173);
or UO_2089 (O_2089,N_40107,N_44042);
and UO_2090 (O_2090,N_45076,N_49593);
nand UO_2091 (O_2091,N_44408,N_45421);
nand UO_2092 (O_2092,N_47211,N_48935);
nand UO_2093 (O_2093,N_49381,N_44022);
or UO_2094 (O_2094,N_49370,N_47122);
nor UO_2095 (O_2095,N_42648,N_42144);
or UO_2096 (O_2096,N_48041,N_49022);
or UO_2097 (O_2097,N_40221,N_42715);
nor UO_2098 (O_2098,N_48443,N_44248);
and UO_2099 (O_2099,N_41065,N_46792);
xnor UO_2100 (O_2100,N_40433,N_43089);
or UO_2101 (O_2101,N_46064,N_40541);
and UO_2102 (O_2102,N_40074,N_47581);
nand UO_2103 (O_2103,N_47995,N_46797);
nor UO_2104 (O_2104,N_47626,N_46270);
nor UO_2105 (O_2105,N_42320,N_47066);
xor UO_2106 (O_2106,N_42754,N_48487);
nor UO_2107 (O_2107,N_43643,N_49960);
or UO_2108 (O_2108,N_49691,N_42388);
nor UO_2109 (O_2109,N_45232,N_40974);
nand UO_2110 (O_2110,N_48382,N_41294);
nand UO_2111 (O_2111,N_43701,N_44744);
nand UO_2112 (O_2112,N_40123,N_48197);
nor UO_2113 (O_2113,N_43029,N_46447);
or UO_2114 (O_2114,N_49864,N_49346);
nand UO_2115 (O_2115,N_46478,N_40343);
xnor UO_2116 (O_2116,N_48883,N_41718);
nor UO_2117 (O_2117,N_41671,N_46963);
nor UO_2118 (O_2118,N_47769,N_47534);
nor UO_2119 (O_2119,N_40592,N_42107);
nand UO_2120 (O_2120,N_48441,N_48310);
or UO_2121 (O_2121,N_43298,N_41199);
nand UO_2122 (O_2122,N_41052,N_40782);
xnor UO_2123 (O_2123,N_42379,N_46712);
nor UO_2124 (O_2124,N_44349,N_44808);
xnor UO_2125 (O_2125,N_41266,N_48555);
nand UO_2126 (O_2126,N_41401,N_44054);
or UO_2127 (O_2127,N_48964,N_43829);
nor UO_2128 (O_2128,N_40399,N_46032);
and UO_2129 (O_2129,N_42164,N_46784);
nand UO_2130 (O_2130,N_41859,N_47002);
and UO_2131 (O_2131,N_48815,N_49061);
nor UO_2132 (O_2132,N_48710,N_41137);
nand UO_2133 (O_2133,N_44512,N_45459);
or UO_2134 (O_2134,N_44213,N_41516);
xor UO_2135 (O_2135,N_42271,N_41492);
nor UO_2136 (O_2136,N_43526,N_40087);
nor UO_2137 (O_2137,N_47921,N_41545);
and UO_2138 (O_2138,N_45161,N_45674);
nor UO_2139 (O_2139,N_41921,N_40801);
nor UO_2140 (O_2140,N_42197,N_42603);
or UO_2141 (O_2141,N_41978,N_41103);
nor UO_2142 (O_2142,N_44663,N_49662);
xor UO_2143 (O_2143,N_47705,N_44323);
and UO_2144 (O_2144,N_41063,N_46757);
nand UO_2145 (O_2145,N_45583,N_42848);
xnor UO_2146 (O_2146,N_41854,N_40247);
or UO_2147 (O_2147,N_49583,N_42877);
or UO_2148 (O_2148,N_46707,N_47032);
xor UO_2149 (O_2149,N_41962,N_48548);
or UO_2150 (O_2150,N_46504,N_44159);
and UO_2151 (O_2151,N_42397,N_40041);
nor UO_2152 (O_2152,N_44062,N_45862);
and UO_2153 (O_2153,N_46581,N_40109);
nand UO_2154 (O_2154,N_48116,N_45084);
nand UO_2155 (O_2155,N_47681,N_40756);
and UO_2156 (O_2156,N_42133,N_47552);
or UO_2157 (O_2157,N_43594,N_42262);
or UO_2158 (O_2158,N_49209,N_42839);
nand UO_2159 (O_2159,N_43954,N_43091);
nand UO_2160 (O_2160,N_40935,N_47958);
nor UO_2161 (O_2161,N_42451,N_42731);
nor UO_2162 (O_2162,N_46770,N_42334);
nor UO_2163 (O_2163,N_43313,N_42187);
nand UO_2164 (O_2164,N_46291,N_42437);
nor UO_2165 (O_2165,N_47815,N_42058);
nor UO_2166 (O_2166,N_41445,N_42489);
and UO_2167 (O_2167,N_49946,N_46913);
nand UO_2168 (O_2168,N_42500,N_46010);
nand UO_2169 (O_2169,N_43642,N_42496);
nand UO_2170 (O_2170,N_42339,N_46510);
nor UO_2171 (O_2171,N_42954,N_46855);
and UO_2172 (O_2172,N_48274,N_44817);
and UO_2173 (O_2173,N_44063,N_42618);
nand UO_2174 (O_2174,N_42142,N_47576);
and UO_2175 (O_2175,N_40996,N_45289);
nor UO_2176 (O_2176,N_49458,N_47547);
nand UO_2177 (O_2177,N_42212,N_43438);
nand UO_2178 (O_2178,N_43540,N_41498);
nand UO_2179 (O_2179,N_41152,N_40066);
and UO_2180 (O_2180,N_49876,N_47460);
and UO_2181 (O_2181,N_44992,N_41362);
nand UO_2182 (O_2182,N_45871,N_47554);
nand UO_2183 (O_2183,N_48649,N_44455);
nor UO_2184 (O_2184,N_41136,N_44993);
nand UO_2185 (O_2185,N_41537,N_43291);
nand UO_2186 (O_2186,N_47793,N_44797);
nand UO_2187 (O_2187,N_41058,N_42663);
nor UO_2188 (O_2188,N_49376,N_47623);
or UO_2189 (O_2189,N_46230,N_40669);
nor UO_2190 (O_2190,N_47480,N_48713);
or UO_2191 (O_2191,N_41632,N_46606);
or UO_2192 (O_2192,N_41386,N_49238);
nor UO_2193 (O_2193,N_45238,N_46217);
or UO_2194 (O_2194,N_43366,N_44310);
xor UO_2195 (O_2195,N_49746,N_42310);
and UO_2196 (O_2196,N_42622,N_44682);
and UO_2197 (O_2197,N_44844,N_44743);
or UO_2198 (O_2198,N_44305,N_40329);
xnor UO_2199 (O_2199,N_40874,N_46549);
or UO_2200 (O_2200,N_46986,N_46751);
xnor UO_2201 (O_2201,N_47394,N_44652);
nor UO_2202 (O_2202,N_40080,N_43268);
nor UO_2203 (O_2203,N_40822,N_48068);
and UO_2204 (O_2204,N_45817,N_40736);
or UO_2205 (O_2205,N_45147,N_46903);
or UO_2206 (O_2206,N_40854,N_45856);
and UO_2207 (O_2207,N_43185,N_48679);
xnor UO_2208 (O_2208,N_48528,N_40092);
nor UO_2209 (O_2209,N_41354,N_48366);
and UO_2210 (O_2210,N_47102,N_43860);
nor UO_2211 (O_2211,N_43665,N_46646);
xnor UO_2212 (O_2212,N_48674,N_40121);
nand UO_2213 (O_2213,N_48961,N_48784);
nand UO_2214 (O_2214,N_45098,N_47126);
xor UO_2215 (O_2215,N_44400,N_49332);
and UO_2216 (O_2216,N_48562,N_46755);
and UO_2217 (O_2217,N_48859,N_42780);
and UO_2218 (O_2218,N_41413,N_46049);
nor UO_2219 (O_2219,N_41844,N_46908);
nor UO_2220 (O_2220,N_43475,N_47302);
or UO_2221 (O_2221,N_42338,N_43724);
nor UO_2222 (O_2222,N_42965,N_47461);
and UO_2223 (O_2223,N_44608,N_41384);
and UO_2224 (O_2224,N_47891,N_49409);
and UO_2225 (O_2225,N_41596,N_47408);
nor UO_2226 (O_2226,N_48595,N_43030);
and UO_2227 (O_2227,N_44639,N_48977);
and UO_2228 (O_2228,N_43402,N_47652);
and UO_2229 (O_2229,N_49048,N_45418);
and UO_2230 (O_2230,N_49220,N_45179);
or UO_2231 (O_2231,N_48911,N_40489);
or UO_2232 (O_2232,N_42471,N_47856);
nor UO_2233 (O_2233,N_46353,N_44178);
or UO_2234 (O_2234,N_40983,N_42280);
and UO_2235 (O_2235,N_40313,N_43404);
xnor UO_2236 (O_2236,N_43265,N_40691);
or UO_2237 (O_2237,N_45649,N_40226);
nor UO_2238 (O_2238,N_42633,N_40114);
xnor UO_2239 (O_2239,N_45731,N_47583);
nor UO_2240 (O_2240,N_43533,N_40889);
and UO_2241 (O_2241,N_49137,N_47527);
xnor UO_2242 (O_2242,N_46615,N_46551);
nand UO_2243 (O_2243,N_43835,N_40270);
nor UO_2244 (O_2244,N_42613,N_48302);
and UO_2245 (O_2245,N_45230,N_49340);
nor UO_2246 (O_2246,N_40186,N_40598);
xnor UO_2247 (O_2247,N_41042,N_44650);
nor UO_2248 (O_2248,N_41521,N_49030);
and UO_2249 (O_2249,N_43654,N_44069);
and UO_2250 (O_2250,N_45188,N_47338);
nor UO_2251 (O_2251,N_41707,N_49494);
and UO_2252 (O_2252,N_41070,N_41343);
and UO_2253 (O_2253,N_40073,N_44635);
nor UO_2254 (O_2254,N_41264,N_43567);
and UO_2255 (O_2255,N_43656,N_43361);
nand UO_2256 (O_2256,N_41534,N_45342);
and UO_2257 (O_2257,N_42147,N_40794);
or UO_2258 (O_2258,N_44116,N_46690);
nand UO_2259 (O_2259,N_45396,N_49710);
nand UO_2260 (O_2260,N_46689,N_48424);
or UO_2261 (O_2261,N_49360,N_47864);
and UO_2262 (O_2262,N_49140,N_45995);
nor UO_2263 (O_2263,N_40344,N_41542);
nand UO_2264 (O_2264,N_43588,N_43044);
nand UO_2265 (O_2265,N_44218,N_41821);
and UO_2266 (O_2266,N_48423,N_49118);
xor UO_2267 (O_2267,N_42185,N_40472);
and UO_2268 (O_2268,N_40642,N_43045);
xnor UO_2269 (O_2269,N_43939,N_45252);
nor UO_2270 (O_2270,N_48536,N_41929);
nand UO_2271 (O_2271,N_46802,N_40285);
nand UO_2272 (O_2272,N_41910,N_47648);
nand UO_2273 (O_2273,N_47449,N_45555);
xnor UO_2274 (O_2274,N_45535,N_45261);
nor UO_2275 (O_2275,N_44230,N_42531);
or UO_2276 (O_2276,N_47355,N_41396);
nor UO_2277 (O_2277,N_40113,N_40030);
nand UO_2278 (O_2278,N_44274,N_43002);
nor UO_2279 (O_2279,N_48970,N_40457);
nor UO_2280 (O_2280,N_46902,N_43752);
nor UO_2281 (O_2281,N_45347,N_43280);
or UO_2282 (O_2282,N_48032,N_44249);
or UO_2283 (O_2283,N_46837,N_43456);
or UO_2284 (O_2284,N_41917,N_48968);
or UO_2285 (O_2285,N_48603,N_49581);
nand UO_2286 (O_2286,N_48762,N_45377);
xor UO_2287 (O_2287,N_46688,N_46339);
xor UO_2288 (O_2288,N_49282,N_46096);
nor UO_2289 (O_2289,N_40396,N_41683);
xor UO_2290 (O_2290,N_46399,N_46468);
nand UO_2291 (O_2291,N_43229,N_46859);
and UO_2292 (O_2292,N_42121,N_43808);
nor UO_2293 (O_2293,N_48346,N_46625);
nand UO_2294 (O_2294,N_49387,N_49096);
or UO_2295 (O_2295,N_41239,N_47450);
nor UO_2296 (O_2296,N_46672,N_43499);
nand UO_2297 (O_2297,N_46132,N_43342);
nor UO_2298 (O_2298,N_40238,N_44997);
or UO_2299 (O_2299,N_40488,N_46069);
nand UO_2300 (O_2300,N_41268,N_48643);
xnor UO_2301 (O_2301,N_43862,N_43529);
nand UO_2302 (O_2302,N_49193,N_47807);
and UO_2303 (O_2303,N_41091,N_48939);
nand UO_2304 (O_2304,N_43738,N_41553);
nor UO_2305 (O_2305,N_45329,N_46001);
nand UO_2306 (O_2306,N_46167,N_43684);
and UO_2307 (O_2307,N_44547,N_45577);
nand UO_2308 (O_2308,N_47713,N_43113);
xnor UO_2309 (O_2309,N_44877,N_41002);
and UO_2310 (O_2310,N_42914,N_49976);
nor UO_2311 (O_2311,N_42137,N_49112);
nor UO_2312 (O_2312,N_43636,N_49449);
and UO_2313 (O_2313,N_45363,N_41491);
or UO_2314 (O_2314,N_41884,N_46678);
nand UO_2315 (O_2315,N_43502,N_49198);
and UO_2316 (O_2316,N_44828,N_45154);
nand UO_2317 (O_2317,N_46286,N_40793);
or UO_2318 (O_2318,N_40424,N_44954);
xor UO_2319 (O_2319,N_43432,N_44515);
and UO_2320 (O_2320,N_43996,N_46414);
and UO_2321 (O_2321,N_45641,N_45927);
or UO_2322 (O_2322,N_49189,N_41674);
nand UO_2323 (O_2323,N_44412,N_46433);
nor UO_2324 (O_2324,N_43439,N_47884);
nand UO_2325 (O_2325,N_47100,N_43839);
nand UO_2326 (O_2326,N_44395,N_48118);
or UO_2327 (O_2327,N_48114,N_40884);
or UO_2328 (O_2328,N_41242,N_46027);
or UO_2329 (O_2329,N_41877,N_48002);
xnor UO_2330 (O_2330,N_44599,N_45153);
nor UO_2331 (O_2331,N_41379,N_49550);
nor UO_2332 (O_2332,N_49988,N_43797);
and UO_2333 (O_2333,N_46575,N_45881);
xor UO_2334 (O_2334,N_45169,N_42772);
and UO_2335 (O_2335,N_43175,N_47438);
and UO_2336 (O_2336,N_42827,N_40863);
and UO_2337 (O_2337,N_41532,N_43521);
and UO_2338 (O_2338,N_42472,N_44871);
or UO_2339 (O_2339,N_41843,N_42230);
or UO_2340 (O_2340,N_47761,N_45481);
and UO_2341 (O_2341,N_46815,N_47767);
nand UO_2342 (O_2342,N_48333,N_44945);
nor UO_2343 (O_2343,N_45177,N_46138);
nor UO_2344 (O_2344,N_49041,N_48834);
nand UO_2345 (O_2345,N_44735,N_44186);
nor UO_2346 (O_2346,N_48954,N_46224);
and UO_2347 (O_2347,N_47896,N_44725);
nor UO_2348 (O_2348,N_48185,N_41615);
xnor UO_2349 (O_2349,N_43583,N_42186);
nand UO_2350 (O_2350,N_44505,N_47563);
nor UO_2351 (O_2351,N_44892,N_43769);
nand UO_2352 (O_2352,N_48832,N_47578);
and UO_2353 (O_2353,N_43668,N_49488);
nand UO_2354 (O_2354,N_46989,N_44429);
nor UO_2355 (O_2355,N_41676,N_43219);
nand UO_2356 (O_2356,N_44714,N_41536);
or UO_2357 (O_2357,N_47858,N_42062);
nor UO_2358 (O_2358,N_47538,N_46557);
or UO_2359 (O_2359,N_44964,N_48054);
nor UO_2360 (O_2360,N_42013,N_49931);
or UO_2361 (O_2361,N_45764,N_47595);
nand UO_2362 (O_2362,N_49785,N_47945);
nor UO_2363 (O_2363,N_44320,N_44781);
and UO_2364 (O_2364,N_48764,N_47483);
nor UO_2365 (O_2365,N_41296,N_48479);
nand UO_2366 (O_2366,N_40500,N_41059);
nor UO_2367 (O_2367,N_41156,N_40897);
nor UO_2368 (O_2368,N_48388,N_49616);
and UO_2369 (O_2369,N_42852,N_43675);
nor UO_2370 (O_2370,N_40622,N_47120);
or UO_2371 (O_2371,N_41346,N_46526);
nor UO_2372 (O_2372,N_43538,N_49014);
nand UO_2373 (O_2373,N_40296,N_40014);
and UO_2374 (O_2374,N_41724,N_45164);
and UO_2375 (O_2375,N_41395,N_42351);
nor UO_2376 (O_2376,N_49681,N_45456);
nand UO_2377 (O_2377,N_41990,N_49751);
and UO_2378 (O_2378,N_45637,N_44684);
or UO_2379 (O_2379,N_42798,N_45634);
and UO_2380 (O_2380,N_48018,N_42825);
nor UO_2381 (O_2381,N_46721,N_48163);
and UO_2382 (O_2382,N_49439,N_40141);
and UO_2383 (O_2383,N_43742,N_48277);
and UO_2384 (O_2384,N_41552,N_44182);
nand UO_2385 (O_2385,N_41008,N_43635);
nand UO_2386 (O_2386,N_43802,N_47974);
xnor UO_2387 (O_2387,N_40266,N_47592);
or UO_2388 (O_2388,N_43386,N_49899);
nor UO_2389 (O_2389,N_48765,N_45143);
nand UO_2390 (O_2390,N_44024,N_48009);
nand UO_2391 (O_2391,N_40026,N_45839);
or UO_2392 (O_2392,N_48851,N_41360);
or UO_2393 (O_2393,N_41026,N_43442);
and UO_2394 (O_2394,N_44870,N_41681);
xor UO_2395 (O_2395,N_46922,N_47464);
or UO_2396 (O_2396,N_43200,N_47103);
xnor UO_2397 (O_2397,N_48591,N_46135);
nand UO_2398 (O_2398,N_46823,N_45219);
or UO_2399 (O_2399,N_47141,N_41605);
nor UO_2400 (O_2400,N_46915,N_49695);
xor UO_2401 (O_2401,N_46185,N_46502);
or UO_2402 (O_2402,N_48694,N_45103);
nand UO_2403 (O_2403,N_44910,N_45167);
xor UO_2404 (O_2404,N_43022,N_40695);
xnor UO_2405 (O_2405,N_46098,N_42942);
nor UO_2406 (O_2406,N_47823,N_45704);
and UO_2407 (O_2407,N_47497,N_46233);
nand UO_2408 (O_2408,N_48171,N_40629);
or UO_2409 (O_2409,N_46522,N_48738);
nand UO_2410 (O_2410,N_49958,N_48249);
or UO_2411 (O_2411,N_45487,N_44374);
and UO_2412 (O_2412,N_42165,N_43991);
nor UO_2413 (O_2413,N_46301,N_44130);
nor UO_2414 (O_2414,N_48524,N_40281);
and UO_2415 (O_2415,N_40105,N_49896);
or UO_2416 (O_2416,N_45362,N_47568);
and UO_2417 (O_2417,N_43041,N_45619);
nor UO_2418 (O_2418,N_40062,N_49650);
or UO_2419 (O_2419,N_43088,N_45380);
nand UO_2420 (O_2420,N_45200,N_40518);
or UO_2421 (O_2421,N_42988,N_48057);
nor UO_2422 (O_2422,N_42828,N_49898);
and UO_2423 (O_2423,N_48180,N_41416);
nor UO_2424 (O_2424,N_48229,N_49451);
xor UO_2425 (O_2425,N_40192,N_43158);
nor UO_2426 (O_2426,N_44696,N_47848);
nand UO_2427 (O_2427,N_41076,N_44156);
nand UO_2428 (O_2428,N_43321,N_47931);
or UO_2429 (O_2429,N_48204,N_44980);
nand UO_2430 (O_2430,N_43199,N_49995);
or UO_2431 (O_2431,N_44361,N_41598);
and UO_2432 (O_2432,N_45870,N_42529);
nand UO_2433 (O_2433,N_47316,N_41709);
nor UO_2434 (O_2434,N_42453,N_43527);
nor UO_2435 (O_2435,N_44138,N_42359);
nand UO_2436 (O_2436,N_41947,N_43422);
nor UO_2437 (O_2437,N_42589,N_40709);
or UO_2438 (O_2438,N_41813,N_47585);
and UO_2439 (O_2439,N_46315,N_45852);
nor UO_2440 (O_2440,N_48393,N_47352);
nand UO_2441 (O_2441,N_42996,N_48225);
and UO_2442 (O_2442,N_40445,N_45671);
and UO_2443 (O_2443,N_41210,N_45987);
nand UO_2444 (O_2444,N_46325,N_43534);
nand UO_2445 (O_2445,N_43942,N_44882);
or UO_2446 (O_2446,N_49498,N_46877);
or UO_2447 (O_2447,N_48507,N_47764);
nor UO_2448 (O_2448,N_43135,N_49057);
nor UO_2449 (O_2449,N_43039,N_46405);
or UO_2450 (O_2450,N_43959,N_42341);
or UO_2451 (O_2451,N_41564,N_48792);
xnor UO_2452 (O_2452,N_42659,N_44189);
or UO_2453 (O_2453,N_40886,N_45609);
nor UO_2454 (O_2454,N_44831,N_44324);
nor UO_2455 (O_2455,N_40124,N_43374);
xor UO_2456 (O_2456,N_47125,N_43500);
xor UO_2457 (O_2457,N_42392,N_42329);
nor UO_2458 (O_2458,N_42523,N_49621);
and UO_2459 (O_2459,N_48658,N_41399);
nor UO_2460 (O_2460,N_49460,N_42952);
or UO_2461 (O_2461,N_41803,N_48716);
xor UO_2462 (O_2462,N_42765,N_42918);
nand UO_2463 (O_2463,N_40513,N_49939);
nor UO_2464 (O_2464,N_48918,N_49497);
nand UO_2465 (O_2465,N_45501,N_47272);
or UO_2466 (O_2466,N_40470,N_42153);
nand UO_2467 (O_2467,N_43967,N_41778);
nand UO_2468 (O_2468,N_48623,N_44634);
or UO_2469 (O_2469,N_46031,N_42568);
and UO_2470 (O_2470,N_46108,N_48791);
or UO_2471 (O_2471,N_49131,N_48593);
xor UO_2472 (O_2472,N_49266,N_45844);
nor UO_2473 (O_2473,N_42593,N_47959);
nor UO_2474 (O_2474,N_47399,N_41351);
nor UO_2475 (O_2475,N_42884,N_40904);
xnor UO_2476 (O_2476,N_40654,N_42464);
and UO_2477 (O_2477,N_45998,N_45105);
nor UO_2478 (O_2478,N_44313,N_42542);
and UO_2479 (O_2479,N_43852,N_44081);
nor UO_2480 (O_2480,N_42438,N_40000);
nor UO_2481 (O_2481,N_44438,N_43661);
xnor UO_2482 (O_2482,N_45432,N_46316);
nor UO_2483 (O_2483,N_49548,N_46163);
xnor UO_2484 (O_2484,N_46393,N_41951);
nor UO_2485 (O_2485,N_43979,N_46970);
and UO_2486 (O_2486,N_42286,N_40714);
xnor UO_2487 (O_2487,N_44291,N_41765);
or UO_2488 (O_2488,N_42030,N_43997);
and UO_2489 (O_2489,N_43935,N_40868);
or UO_2490 (O_2490,N_46844,N_49603);
and UO_2491 (O_2491,N_46766,N_45675);
or UO_2492 (O_2492,N_48251,N_42859);
or UO_2493 (O_2493,N_47182,N_48047);
or UO_2494 (O_2494,N_48174,N_47191);
nand UO_2495 (O_2495,N_43322,N_45044);
nand UO_2496 (O_2496,N_46187,N_45646);
nand UO_2497 (O_2497,N_44777,N_45192);
and UO_2498 (O_2498,N_49095,N_49880);
xnor UO_2499 (O_2499,N_40478,N_44074);
nor UO_2500 (O_2500,N_43355,N_47727);
nor UO_2501 (O_2501,N_48551,N_40200);
nor UO_2502 (O_2502,N_48601,N_49468);
or UO_2503 (O_2503,N_48641,N_43710);
or UO_2504 (O_2504,N_49283,N_45914);
nand UO_2505 (O_2505,N_46506,N_49339);
nand UO_2506 (O_2506,N_44862,N_47326);
nand UO_2507 (O_2507,N_43798,N_45422);
and UO_2508 (O_2508,N_40182,N_41997);
xnor UO_2509 (O_2509,N_48231,N_46503);
or UO_2510 (O_2510,N_45584,N_43173);
xnor UO_2511 (O_2511,N_48403,N_40268);
nand UO_2512 (O_2512,N_42224,N_40957);
nand UO_2513 (O_2513,N_49018,N_48850);
or UO_2514 (O_2514,N_43038,N_40393);
xor UO_2515 (O_2515,N_42090,N_45021);
xor UO_2516 (O_2516,N_40177,N_46782);
xnor UO_2517 (O_2517,N_42466,N_49715);
and UO_2518 (O_2518,N_43555,N_47749);
nand UO_2519 (O_2519,N_40657,N_47878);
or UO_2520 (O_2520,N_42713,N_42301);
nand UO_2521 (O_2521,N_48813,N_47135);
xor UO_2522 (O_2522,N_47775,N_41029);
and UO_2523 (O_2523,N_44697,N_49502);
nor UO_2524 (O_2524,N_47401,N_47685);
nor UO_2525 (O_2525,N_49290,N_44897);
or UO_2526 (O_2526,N_49075,N_40851);
nand UO_2527 (O_2527,N_43297,N_48025);
and UO_2528 (O_2528,N_40021,N_47548);
nor UO_2529 (O_2529,N_43037,N_43330);
nand UO_2530 (O_2530,N_42059,N_48673);
and UO_2531 (O_2531,N_44075,N_46262);
nand UO_2532 (O_2532,N_44214,N_45007);
and UO_2533 (O_2533,N_43989,N_45618);
and UO_2534 (O_2534,N_46067,N_44607);
xnor UO_2535 (O_2535,N_40171,N_48271);
or UO_2536 (O_2536,N_45834,N_41565);
nand UO_2537 (O_2537,N_48071,N_40458);
nor UO_2538 (O_2538,N_41752,N_44414);
and UO_2539 (O_2539,N_44971,N_41159);
or UO_2540 (O_2540,N_43169,N_43441);
and UO_2541 (O_2541,N_47852,N_46935);
nor UO_2542 (O_2542,N_45415,N_40915);
and UO_2543 (O_2543,N_46474,N_44445);
nand UO_2544 (O_2544,N_46373,N_41554);
nand UO_2545 (O_2545,N_46791,N_46669);
xor UO_2546 (O_2546,N_48000,N_47250);
and UO_2547 (O_2547,N_46822,N_48902);
nand UO_2548 (O_2548,N_47325,N_42046);
xnor UO_2549 (O_2549,N_46886,N_48384);
nor UO_2550 (O_2550,N_44331,N_45558);
and UO_2551 (O_2551,N_46519,N_41689);
or UO_2552 (O_2552,N_46371,N_44788);
nand UO_2553 (O_2553,N_42139,N_46112);
nor UO_2554 (O_2554,N_40689,N_48630);
nor UO_2555 (O_2555,N_44713,N_42408);
nor UO_2556 (O_2556,N_44100,N_48158);
or UO_2557 (O_2557,N_44107,N_47949);
and UO_2558 (O_2558,N_47998,N_40451);
or UO_2559 (O_2559,N_48475,N_46827);
or UO_2560 (O_2560,N_47079,N_46665);
or UO_2561 (O_2561,N_46419,N_41729);
and UO_2562 (O_2562,N_46411,N_44031);
or UO_2563 (O_2563,N_42866,N_40940);
and UO_2564 (O_2564,N_46048,N_46624);
nand UO_2565 (O_2565,N_49642,N_46685);
and UO_2566 (O_2566,N_47587,N_46726);
and UO_2567 (O_2567,N_49320,N_43864);
nand UO_2568 (O_2568,N_40230,N_48546);
nor UO_2569 (O_2569,N_41229,N_41530);
nand UO_2570 (O_2570,N_43501,N_48349);
nor UO_2571 (O_2571,N_46795,N_46808);
nand UO_2572 (O_2572,N_41678,N_49878);
nand UO_2573 (O_2573,N_48670,N_46533);
and UO_2574 (O_2574,N_48828,N_45873);
nor UO_2575 (O_2575,N_48281,N_46424);
xnor UO_2576 (O_2576,N_45484,N_49950);
nor UO_2577 (O_2577,N_48956,N_47435);
nand UO_2578 (O_2578,N_44464,N_42283);
nand UO_2579 (O_2579,N_40383,N_46439);
nor UO_2580 (O_2580,N_47611,N_44726);
xnor UO_2581 (O_2581,N_48976,N_48696);
xnor UO_2582 (O_2582,N_43409,N_40249);
and UO_2583 (O_2583,N_41168,N_49795);
and UO_2584 (O_2584,N_43951,N_43371);
nand UO_2585 (O_2585,N_43662,N_42813);
and UO_2586 (O_2586,N_41477,N_40959);
nor UO_2587 (O_2587,N_44208,N_40805);
nor UO_2588 (O_2588,N_44694,N_43397);
nand UO_2589 (O_2589,N_49575,N_47619);
nand UO_2590 (O_2590,N_43001,N_40726);
or UO_2591 (O_2591,N_47968,N_45967);
nor UO_2592 (O_2592,N_43277,N_42588);
nor UO_2593 (O_2593,N_47854,N_49857);
xor UO_2594 (O_2594,N_45473,N_44695);
nor UO_2595 (O_2595,N_40772,N_43708);
xnor UO_2596 (O_2596,N_42124,N_42467);
or UO_2597 (O_2597,N_48084,N_49374);
nand UO_2598 (O_2598,N_44766,N_48590);
nand UO_2599 (O_2599,N_46748,N_44555);
and UO_2600 (O_2600,N_45429,N_42508);
and UO_2601 (O_2601,N_49375,N_40303);
xor UO_2602 (O_2602,N_42316,N_41744);
nor UO_2603 (O_2603,N_40032,N_42597);
or UO_2604 (O_2604,N_43083,N_42176);
and UO_2605 (O_2605,N_46865,N_49919);
and UO_2606 (O_2606,N_41779,N_48126);
nor UO_2607 (O_2607,N_43747,N_45125);
and UO_2608 (O_2608,N_43416,N_49789);
nor UO_2609 (O_2609,N_45065,N_45993);
xor UO_2610 (O_2610,N_43815,N_41024);
and UO_2611 (O_2611,N_45988,N_43031);
nor UO_2612 (O_2612,N_49576,N_49270);
xor UO_2613 (O_2613,N_44678,N_40958);
nor UO_2614 (O_2614,N_43213,N_48691);
nand UO_2615 (O_2615,N_46370,N_49357);
or UO_2616 (O_2616,N_43413,N_46137);
nand UO_2617 (O_2617,N_46532,N_47368);
nand UO_2618 (O_2618,N_47898,N_49093);
or UO_2619 (O_2619,N_49195,N_46488);
xnor UO_2620 (O_2620,N_42270,N_40157);
nor UO_2621 (O_2621,N_49538,N_44810);
or UO_2622 (O_2622,N_48187,N_45697);
xor UO_2623 (O_2623,N_49571,N_42875);
nand UO_2624 (O_2624,N_43584,N_45840);
nor UO_2625 (O_2625,N_48221,N_44798);
xnor UO_2626 (O_2626,N_42703,N_48704);
nand UO_2627 (O_2627,N_49507,N_45537);
xor UO_2628 (O_2628,N_47442,N_42586);
nand UO_2629 (O_2629,N_41998,N_40325);
nand UO_2630 (O_2630,N_46364,N_42795);
nor UO_2631 (O_2631,N_42470,N_49207);
or UO_2632 (O_2632,N_43294,N_42649);
nand UO_2633 (O_2633,N_48719,N_42269);
and UO_2634 (O_2634,N_46769,N_44345);
or UO_2635 (O_2635,N_47093,N_42880);
or UO_2636 (O_2636,N_43700,N_48777);
xnor UO_2637 (O_2637,N_40821,N_48269);
nand UO_2638 (O_2638,N_43866,N_45610);
or UO_2639 (O_2639,N_48064,N_43585);
xnor UO_2640 (O_2640,N_48053,N_49663);
xnor UO_2641 (O_2641,N_47925,N_40287);
and UO_2642 (O_2642,N_46056,N_49459);
or UO_2643 (O_2643,N_43910,N_40085);
nor UO_2644 (O_2644,N_49249,N_48175);
or UO_2645 (O_2645,N_44615,N_41003);
nor UO_2646 (O_2646,N_49891,N_44077);
or UO_2647 (O_2647,N_42398,N_41225);
or UO_2648 (O_2648,N_49353,N_49645);
and UO_2649 (O_2649,N_44256,N_49577);
or UO_2650 (O_2650,N_43577,N_47605);
or UO_2651 (O_2651,N_44143,N_47252);
or UO_2652 (O_2652,N_46840,N_49970);
nor UO_2653 (O_2653,N_48387,N_49186);
or UO_2654 (O_2654,N_42737,N_45034);
xnor UO_2655 (O_2655,N_49520,N_43189);
and UO_2656 (O_2656,N_42021,N_44736);
and UO_2657 (O_2657,N_46365,N_42447);
nor UO_2658 (O_2658,N_45579,N_40462);
nor UO_2659 (O_2659,N_43398,N_40991);
nand UO_2660 (O_2660,N_44672,N_45907);
nor UO_2661 (O_2661,N_46312,N_42747);
and UO_2662 (O_2662,N_40467,N_47387);
and UO_2663 (O_2663,N_48511,N_43357);
or UO_2664 (O_2664,N_41686,N_49206);
or UO_2665 (O_2665,N_44513,N_44968);
nor UO_2666 (O_2666,N_48457,N_46906);
nor UO_2667 (O_2667,N_41825,N_46212);
and UO_2668 (O_2668,N_49145,N_45681);
nand UO_2669 (O_2669,N_44889,N_46431);
and UO_2670 (O_2670,N_46724,N_44500);
and UO_2671 (O_2671,N_48871,N_46220);
nor UO_2672 (O_2672,N_41602,N_47929);
nor UO_2673 (O_2673,N_42547,N_41646);
and UO_2674 (O_2674,N_42369,N_40213);
nand UO_2675 (O_2675,N_43503,N_42170);
xnor UO_2676 (O_2676,N_49412,N_49044);
and UO_2677 (O_2677,N_44977,N_45759);
nand UO_2678 (O_2678,N_43349,N_45397);
nor UO_2679 (O_2679,N_45832,N_46985);
nor UO_2680 (O_2680,N_41793,N_48325);
nand UO_2681 (O_2681,N_43688,N_46385);
or UO_2682 (O_2682,N_46951,N_42841);
or UO_2683 (O_2683,N_41254,N_46452);
and UO_2684 (O_2684,N_44000,N_47567);
xor UO_2685 (O_2685,N_41424,N_42234);
or UO_2686 (O_2686,N_42890,N_46475);
and UO_2687 (O_2687,N_46943,N_49648);
or UO_2688 (O_2688,N_49579,N_47006);
xor UO_2689 (O_2689,N_45928,N_49793);
and UO_2690 (O_2690,N_44270,N_48081);
nand UO_2691 (O_2691,N_40602,N_43871);
nor UO_2692 (O_2692,N_43494,N_45307);
or UO_2693 (O_2693,N_45312,N_47887);
or UO_2694 (O_2694,N_49716,N_43948);
nand UO_2695 (O_2695,N_42919,N_45888);
and UO_2696 (O_2696,N_44034,N_41968);
or UO_2697 (O_2697,N_49141,N_42284);
nor UO_2698 (O_2698,N_47353,N_45204);
and UO_2699 (O_2699,N_42018,N_45700);
xor UO_2700 (O_2700,N_48886,N_45765);
or UO_2701 (O_2701,N_49625,N_45442);
and UO_2702 (O_2702,N_45951,N_47367);
nor UO_2703 (O_2703,N_49382,N_47725);
nor UO_2704 (O_2704,N_46741,N_47425);
nor UO_2705 (O_2705,N_44251,N_41827);
and UO_2706 (O_2706,N_46705,N_45330);
nor UO_2707 (O_2707,N_41345,N_43582);
nand UO_2708 (O_2708,N_45608,N_47721);
nor UO_2709 (O_2709,N_43758,N_41801);
or UO_2710 (O_2710,N_43612,N_43599);
or UO_2711 (O_2711,N_43604,N_42647);
xnor UO_2712 (O_2712,N_44304,N_44019);
and UO_2713 (O_2713,N_47452,N_47819);
or UO_2714 (O_2714,N_41617,N_43644);
and UO_2715 (O_2715,N_42801,N_45350);
nand UO_2716 (O_2716,N_40879,N_45727);
nand UO_2717 (O_2717,N_41272,N_42621);
nand UO_2718 (O_2718,N_43563,N_42387);
nor UO_2719 (O_2719,N_49774,N_44046);
nor UO_2720 (O_2720,N_43054,N_44109);
and UO_2721 (O_2721,N_49549,N_48929);
nand UO_2722 (O_2722,N_45058,N_45941);
and UO_2723 (O_2723,N_48756,N_48255);
or UO_2724 (O_2724,N_49688,N_42196);
nor UO_2725 (O_2725,N_41108,N_47655);
or UO_2726 (O_2726,N_47137,N_45552);
nor UO_2727 (O_2727,N_44385,N_41278);
or UO_2728 (O_2728,N_48890,N_45170);
or UO_2729 (O_2729,N_48526,N_48124);
and UO_2730 (O_2730,N_45092,N_49622);
nor UO_2731 (O_2731,N_43237,N_44670);
nor UO_2732 (O_2732,N_49969,N_40071);
nor UO_2733 (O_2733,N_48426,N_40871);
nor UO_2734 (O_2734,N_47642,N_46223);
nor UO_2735 (O_2735,N_47770,N_40347);
and UO_2736 (O_2736,N_46160,N_42783);
nand UO_2737 (O_2737,N_48359,N_44234);
or UO_2738 (O_2738,N_46682,N_45290);
and UO_2739 (O_2739,N_45251,N_40091);
and UO_2740 (O_2740,N_46253,N_46697);
nand UO_2741 (O_2741,N_41144,N_42291);
nand UO_2742 (O_2742,N_49110,N_43303);
or UO_2743 (O_2743,N_42484,N_41447);
and UO_2744 (O_2744,N_45585,N_40136);
nor UO_2745 (O_2745,N_48753,N_43315);
and UO_2746 (O_2746,N_48698,N_43340);
and UO_2747 (O_2747,N_44241,N_46860);
or UO_2748 (O_2748,N_45530,N_42978);
xor UO_2749 (O_2749,N_43120,N_47659);
nor UO_2750 (O_2750,N_49665,N_41679);
and UO_2751 (O_2751,N_45212,N_45149);
and UO_2752 (O_2752,N_47134,N_48559);
and UO_2753 (O_2753,N_44574,N_42409);
and UO_2754 (O_2754,N_45958,N_44357);
nor UO_2755 (O_2755,N_48309,N_49858);
and UO_2756 (O_2756,N_45890,N_41427);
and UO_2757 (O_2757,N_45171,N_40639);
xor UO_2758 (O_2758,N_48449,N_48213);
and UO_2759 (O_2759,N_42820,N_45496);
xnor UO_2760 (O_2760,N_47679,N_48746);
or UO_2761 (O_2761,N_43415,N_43617);
or UO_2762 (O_2762,N_49822,N_46311);
xor UO_2763 (O_2763,N_42645,N_46709);
or UO_2764 (O_2764,N_44199,N_49204);
nand UO_2765 (O_2765,N_42272,N_43487);
or UO_2766 (O_2766,N_44124,N_40188);
nand UO_2767 (O_2767,N_40481,N_41983);
and UO_2768 (O_2768,N_45658,N_49539);
nand UO_2769 (O_2769,N_46272,N_40720);
nor UO_2770 (O_2770,N_40811,N_45452);
nor UO_2771 (O_2771,N_44712,N_45898);
or UO_2772 (O_2772,N_45378,N_46109);
or UO_2773 (O_2773,N_41905,N_44707);
nor UO_2774 (O_2774,N_47981,N_49117);
nor UO_2775 (O_2775,N_49922,N_49071);
nand UO_2776 (O_2776,N_46843,N_41628);
nor UO_2777 (O_2777,N_45721,N_45761);
and UO_2778 (O_2778,N_48602,N_44894);
nand UO_2779 (O_2779,N_49664,N_47809);
nor UO_2780 (O_2780,N_42781,N_40783);
nor UO_2781 (O_2781,N_47939,N_46000);
or UO_2782 (O_2782,N_40426,N_43581);
or UO_2783 (O_2783,N_43149,N_48011);
xor UO_2784 (O_2784,N_48797,N_47194);
nand UO_2785 (O_2785,N_46047,N_44144);
or UO_2786 (O_2786,N_41446,N_48646);
and UO_2787 (O_2787,N_47445,N_40921);
nor UO_2788 (O_2788,N_45730,N_42752);
and UO_2789 (O_2789,N_48666,N_49163);
nor UO_2790 (O_2790,N_43794,N_49279);
and UO_2791 (O_2791,N_43177,N_46209);
and UO_2792 (O_2792,N_46268,N_42518);
or UO_2793 (O_2793,N_46930,N_44884);
nand UO_2794 (O_2794,N_44076,N_45901);
or UO_2795 (O_2795,N_40468,N_46975);
nand UO_2796 (O_2796,N_47615,N_49552);
or UO_2797 (O_2797,N_40452,N_40201);
and UO_2798 (O_2798,N_46152,N_46810);
xor UO_2799 (O_2799,N_42363,N_47647);
nand UO_2800 (O_2800,N_49647,N_45802);
xor UO_2801 (O_2801,N_46964,N_48742);
nand UO_2802 (O_2802,N_47562,N_42932);
or UO_2803 (O_2803,N_48895,N_42486);
nor UO_2804 (O_2804,N_43015,N_45453);
or UO_2805 (O_2805,N_49214,N_48757);
nand UO_2806 (O_2806,N_40594,N_47216);
nor UO_2807 (O_2807,N_48374,N_48616);
xor UO_2808 (O_2808,N_40532,N_44391);
and UO_2809 (O_2809,N_47256,N_44294);
nor UO_2810 (O_2810,N_45776,N_47669);
nand UO_2811 (O_2811,N_41984,N_47489);
nand UO_2812 (O_2812,N_42343,N_43092);
or UO_2813 (O_2813,N_47341,N_42519);
nand UO_2814 (O_2814,N_40305,N_49646);
nand UO_2815 (O_2815,N_46993,N_41150);
nor UO_2816 (O_2816,N_40543,N_42899);
or UO_2817 (O_2817,N_46653,N_47305);
or UO_2818 (O_2818,N_49064,N_41333);
nor UO_2819 (O_2819,N_48029,N_49784);
nor UO_2820 (O_2820,N_40022,N_43902);
nand UO_2821 (O_2821,N_49236,N_43450);
nor UO_2822 (O_2822,N_47107,N_47226);
and UO_2823 (O_2823,N_45669,N_49983);
nor UO_2824 (O_2824,N_44293,N_48280);
nand UO_2825 (O_2825,N_41366,N_46247);
nand UO_2826 (O_2826,N_44014,N_43659);
nor UO_2827 (O_2827,N_42681,N_48891);
nand UO_2828 (O_2828,N_47254,N_45592);
and UO_2829 (O_2829,N_44953,N_49636);
or UO_2830 (O_2830,N_49284,N_49492);
and UO_2831 (O_2831,N_44657,N_49244);
nand UO_2832 (O_2832,N_41959,N_41852);
and UO_2833 (O_2833,N_44541,N_44071);
nand UO_2834 (O_2834,N_46651,N_46300);
and UO_2835 (O_2835,N_47677,N_44448);
and UO_2836 (O_2836,N_46904,N_47674);
nor UO_2837 (O_2837,N_44300,N_46369);
nand UO_2838 (O_2838,N_48928,N_41727);
or UO_2839 (O_2839,N_48543,N_41043);
and UO_2840 (O_2840,N_44842,N_42998);
nand UO_2841 (O_2841,N_49293,N_40455);
or UO_2842 (O_2842,N_43428,N_43592);
nand UO_2843 (O_2843,N_42188,N_42146);
and UO_2844 (O_2844,N_46151,N_45270);
and UO_2845 (O_2845,N_42047,N_42248);
nor UO_2846 (O_2846,N_40597,N_49503);
or UO_2847 (O_2847,N_42581,N_41129);
nand UO_2848 (O_2848,N_44149,N_41236);
nand UO_2849 (O_2849,N_49461,N_41535);
nand UO_2850 (O_2850,N_42887,N_47710);
nand UO_2851 (O_2851,N_43923,N_49963);
or UO_2852 (O_2852,N_42473,N_40368);
or UO_2853 (O_2853,N_41066,N_44565);
nand UO_2854 (O_2854,N_40086,N_42640);
nor UO_2855 (O_2855,N_41640,N_47703);
and UO_2856 (O_2856,N_40628,N_42696);
nor UO_2857 (O_2857,N_40664,N_42807);
nor UO_2858 (O_2858,N_49792,N_46852);
xnor UO_2859 (O_2859,N_43831,N_42462);
and UO_2860 (O_2860,N_43702,N_45475);
nand UO_2861 (O_2861,N_47978,N_46828);
xnor UO_2862 (O_2862,N_46130,N_44927);
nor UO_2863 (O_2863,N_45748,N_43573);
and UO_2864 (O_2864,N_47380,N_43440);
nor UO_2865 (O_2865,N_48930,N_42718);
nand UO_2866 (O_2866,N_41733,N_45590);
nor UO_2867 (O_2867,N_41101,N_41606);
or UO_2868 (O_2868,N_42132,N_44637);
nand UO_2869 (O_2869,N_48731,N_46765);
and UO_2870 (O_2870,N_47083,N_47549);
nor UO_2871 (O_2871,N_49853,N_45760);
nor UO_2872 (O_2872,N_40768,N_49271);
nand UO_2873 (O_2873,N_49115,N_48096);
nand UO_2874 (O_2874,N_48811,N_47088);
and UO_2875 (O_2875,N_41170,N_47829);
nand UO_2876 (O_2876,N_46745,N_41134);
or UO_2877 (O_2877,N_43637,N_48019);
and UO_2878 (O_2878,N_46511,N_49453);
nand UO_2879 (O_2879,N_45271,N_43190);
nor UO_2880 (O_2880,N_45642,N_40820);
or UO_2881 (O_2881,N_42349,N_48978);
and UO_2882 (O_2882,N_40733,N_45935);
xor UO_2883 (O_2883,N_42131,N_43040);
nor UO_2884 (O_2884,N_43775,N_47261);
and UO_2885 (O_2885,N_48209,N_43047);
nand UO_2886 (O_2886,N_43305,N_42167);
or UO_2887 (O_2887,N_45691,N_40943);
or UO_2888 (O_2888,N_43980,N_48563);
or UO_2889 (O_2889,N_48947,N_47948);
and UO_2890 (O_2890,N_41271,N_44912);
nor UO_2891 (O_2891,N_47594,N_44710);
xnor UO_2892 (O_2892,N_46144,N_44709);
nor UO_2893 (O_2893,N_43560,N_49530);
xnor UO_2894 (O_2894,N_43868,N_40876);
or UO_2895 (O_2895,N_46853,N_41540);
or UO_2896 (O_2896,N_40860,N_46368);
and UO_2897 (O_2897,N_47245,N_42116);
nor UO_2898 (O_2898,N_44396,N_48080);
or UO_2899 (O_2899,N_43950,N_48070);
and UO_2900 (O_2900,N_45887,N_43486);
and UO_2901 (O_2901,N_41157,N_46775);
and UO_2902 (O_2902,N_44285,N_47049);
xnor UO_2903 (O_2903,N_44838,N_48827);
xor UO_2904 (O_2904,N_43043,N_45497);
and UO_2905 (O_2905,N_45931,N_49092);
nand UO_2906 (O_2906,N_42695,N_48104);
and UO_2907 (O_2907,N_43363,N_48485);
and UO_2908 (O_2908,N_43914,N_46338);
nor UO_2909 (O_2909,N_41899,N_40502);
nor UO_2910 (O_2910,N_40658,N_47285);
and UO_2911 (O_2911,N_48365,N_42984);
nand UO_2912 (O_2912,N_43608,N_40240);
nand UO_2913 (O_2913,N_43513,N_40061);
nand UO_2914 (O_2914,N_48621,N_48442);
xor UO_2915 (O_2915,N_40697,N_42689);
and UO_2916 (O_2916,N_42260,N_49915);
and UO_2917 (O_2917,N_47054,N_43462);
nand UO_2918 (O_2918,N_41954,N_42968);
nand UO_2919 (O_2919,N_44544,N_46465);
nand UO_2920 (O_2920,N_42904,N_43383);
nor UO_2921 (O_2921,N_44539,N_48427);
or UO_2922 (O_2922,N_49265,N_48498);
xnor UO_2923 (O_2923,N_47463,N_49554);
nor UO_2924 (O_2924,N_47164,N_47629);
or UO_2925 (O_2925,N_42948,N_43421);
or UO_2926 (O_2926,N_48067,N_42768);
and UO_2927 (O_2927,N_40352,N_44601);
xor UO_2928 (O_2928,N_44573,N_40919);
nor UO_2929 (O_2929,N_48537,N_41216);
or UO_2930 (O_2930,N_47362,N_43489);
and UO_2931 (O_2931,N_40001,N_43419);
or UO_2932 (O_2932,N_44480,N_44026);
and UO_2933 (O_2933,N_49047,N_47212);
or UO_2934 (O_2934,N_48780,N_44282);
nor UO_2935 (O_2935,N_45566,N_40906);
nand UO_2936 (O_2936,N_47000,N_43052);
and UO_2937 (O_2937,N_47042,N_40576);
nor UO_2938 (O_2938,N_41245,N_43444);
and UO_2939 (O_2939,N_44375,N_42907);
nand UO_2940 (O_2940,N_48058,N_46407);
or UO_2941 (O_2941,N_46925,N_40359);
nand UO_2942 (O_2942,N_43676,N_40010);
and UO_2943 (O_2943,N_47111,N_44761);
and UO_2944 (O_2944,N_42426,N_43809);
or UO_2945 (O_2945,N_44160,N_47874);
nand UO_2946 (O_2946,N_40011,N_45925);
xnor UO_2947 (O_2947,N_42112,N_43255);
and UO_2948 (O_2948,N_45490,N_48122);
nand UO_2949 (O_2949,N_43813,N_43964);
nor UO_2950 (O_2950,N_45435,N_44093);
and UO_2951 (O_2951,N_41886,N_40918);
nor UO_2952 (O_2952,N_41113,N_47390);
or UO_2953 (O_2953,N_49834,N_45441);
and UO_2954 (O_2954,N_45828,N_48399);
and UO_2955 (O_2955,N_48936,N_45172);
nand UO_2956 (O_2956,N_43385,N_46087);
nor UO_2957 (O_2957,N_47288,N_44273);
or UO_2958 (O_2958,N_47900,N_45019);
nand UO_2959 (O_2959,N_41881,N_41356);
nor UO_2960 (O_2960,N_41075,N_42730);
nand UO_2961 (O_2961,N_44128,N_47323);
nand UO_2962 (O_2962,N_40855,N_40300);
or UO_2963 (O_2963,N_40750,N_40375);
nand UO_2964 (O_2964,N_48413,N_41668);
and UO_2965 (O_2965,N_43103,N_45705);
or UO_2966 (O_2966,N_42879,N_42987);
nor UO_2967 (O_2967,N_44358,N_43603);
nand UO_2968 (O_2968,N_40370,N_45962);
or UO_2969 (O_2969,N_42992,N_43429);
nand UO_2970 (O_2970,N_40966,N_40404);
or UO_2971 (O_2971,N_47715,N_42259);
or UO_2972 (O_2972,N_46412,N_49545);
nand UO_2973 (O_2973,N_45083,N_44005);
nor UO_2974 (O_2974,N_47477,N_43225);
nand UO_2975 (O_2975,N_45121,N_48348);
and UO_2976 (O_2976,N_49444,N_47004);
xor UO_2977 (O_2977,N_47386,N_48133);
nor UO_2978 (O_2978,N_49652,N_47609);
nor UO_2979 (O_2979,N_44733,N_46552);
or UO_2980 (O_2980,N_49121,N_48708);
nor UO_2981 (O_2981,N_42509,N_43714);
nand UO_2982 (O_2982,N_40699,N_47084);
and UO_2983 (O_2983,N_40306,N_49334);
xnor UO_2984 (O_2984,N_49619,N_41680);
nor UO_2985 (O_2985,N_48491,N_44461);
nand UO_2986 (O_2986,N_42096,N_42256);
and UO_2987 (O_2987,N_40651,N_47027);
nor UO_2988 (O_2988,N_49326,N_48882);
xor UO_2989 (O_2989,N_43109,N_45313);
nand UO_2990 (O_2990,N_41695,N_49011);
and UO_2991 (O_2991,N_47556,N_49653);
nor UO_2992 (O_2992,N_43098,N_42963);
xor UO_2993 (O_2993,N_41860,N_43547);
nor UO_2994 (O_2994,N_48396,N_46184);
or UO_2995 (O_2995,N_41624,N_42366);
xnor UO_2996 (O_2996,N_43180,N_49191);
nand UO_2997 (O_2997,N_42717,N_45337);
and UO_2998 (O_2998,N_49563,N_47105);
and UO_2999 (O_2999,N_41664,N_41608);
nand UO_3000 (O_3000,N_47599,N_41049);
and UO_3001 (O_3001,N_43167,N_42587);
nand UO_3002 (O_3002,N_43483,N_45323);
or UO_3003 (O_3003,N_40242,N_45529);
nor UO_3004 (O_3004,N_49605,N_48523);
nor UO_3005 (O_3005,N_42240,N_42830);
and UO_3006 (O_3006,N_40309,N_42682);
xor UO_3007 (O_3007,N_49185,N_46594);
nor UO_3008 (O_3008,N_43245,N_43484);
nand UO_3009 (O_3009,N_44869,N_48967);
xor UO_3010 (O_3010,N_49233,N_43093);
xnor UO_3011 (O_3011,N_40334,N_40051);
or UO_3012 (O_3012,N_47404,N_41577);
nand UO_3013 (O_3013,N_41667,N_48596);
and UO_3014 (O_3014,N_48344,N_40803);
or UO_3015 (O_3015,N_40039,N_46932);
nand UO_3016 (O_3016,N_47806,N_47944);
xor UO_3017 (O_3017,N_45884,N_41012);
and UO_3018 (O_3018,N_48894,N_42985);
or UO_3019 (O_3019,N_43220,N_40766);
nor UO_3020 (O_3020,N_44741,N_44491);
or UO_3021 (O_3021,N_46695,N_42838);
nor UO_3022 (O_3022,N_43898,N_40210);
nand UO_3023 (O_3023,N_40903,N_45111);
nand UO_3024 (O_3024,N_48671,N_43275);
nand UO_3025 (O_3025,N_45879,N_48090);
nor UO_3026 (O_3026,N_49697,N_43828);
xnor UO_3027 (O_3027,N_46982,N_45221);
nor UO_3028 (O_3028,N_49772,N_48988);
nand UO_3029 (O_3029,N_46025,N_45893);
xor UO_3030 (O_3030,N_44731,N_47909);
or UO_3031 (O_3031,N_42861,N_45356);
nand UO_3032 (O_3032,N_41081,N_48502);
and UO_3033 (O_3033,N_40366,N_49875);
nand UO_3034 (O_3034,N_49651,N_43145);
or UO_3035 (O_3035,N_45997,N_49037);
and UO_3036 (O_3036,N_49744,N_49068);
or UO_3037 (O_3037,N_46034,N_41809);
nor UO_3038 (O_3038,N_43068,N_45718);
xor UO_3039 (O_3039,N_44118,N_40314);
nor UO_3040 (O_3040,N_44423,N_49700);
nand UO_3041 (O_3041,N_40976,N_42103);
nor UO_3042 (O_3042,N_40139,N_44325);
or UO_3043 (O_3043,N_47248,N_42123);
nor UO_3044 (O_3044,N_41610,N_43596);
and UO_3045 (O_3045,N_42809,N_40936);
xnor UO_3046 (O_3046,N_49081,N_44466);
or UO_3047 (O_3047,N_44603,N_41308);
or UO_3048 (O_3048,N_43087,N_42929);
or UO_3049 (O_3049,N_47195,N_48470);
nand UO_3050 (O_3050,N_45073,N_45054);
xor UO_3051 (O_3051,N_40363,N_41376);
nor UO_3052 (O_3052,N_40494,N_40583);
nor UO_3053 (O_3053,N_44099,N_41985);
nand UO_3054 (O_3054,N_43325,N_48927);
or UO_3055 (O_3055,N_46858,N_44421);
or UO_3056 (O_3056,N_42326,N_41453);
nand UO_3057 (O_3057,N_44276,N_42552);
nand UO_3058 (O_3058,N_46681,N_41140);
or UO_3059 (O_3059,N_41450,N_41499);
and UO_3060 (O_3060,N_44171,N_43476);
nand UO_3061 (O_3061,N_45788,N_41126);
nand UO_3062 (O_3062,N_46037,N_42897);
nor UO_3063 (O_3063,N_41176,N_42679);
or UO_3064 (O_3064,N_45950,N_48958);
and UO_3065 (O_3065,N_40231,N_41392);
xor UO_3066 (O_3066,N_41119,N_41022);
or UO_3067 (O_3067,N_48072,N_45622);
nor UO_3068 (O_3068,N_42325,N_46055);
nand UO_3069 (O_3069,N_45744,N_48606);
nor UO_3070 (O_3070,N_49917,N_40774);
or UO_3071 (O_3071,N_44162,N_48439);
nand UO_3072 (O_3072,N_41508,N_49316);
nand UO_3073 (O_3073,N_48168,N_45773);
nor UO_3074 (O_3074,N_41349,N_44723);
nand UO_3075 (O_3075,N_46252,N_46046);
xor UO_3076 (O_3076,N_48529,N_44860);
or UO_3077 (O_3077,N_47720,N_49824);
and UO_3078 (O_3078,N_46962,N_45086);
xnor UO_3079 (O_3079,N_44782,N_45795);
nor UO_3080 (O_3080,N_41260,N_41151);
xor UO_3081 (O_3081,N_40931,N_49966);
and UO_3082 (O_3082,N_47528,N_43609);
or UO_3083 (O_3083,N_49470,N_46500);
and UO_3084 (O_3084,N_45719,N_47324);
and UO_3085 (O_3085,N_45580,N_49693);
nor UO_3086 (O_3086,N_47374,N_41774);
and UO_3087 (O_3087,N_44949,N_49807);
nor UO_3088 (O_3088,N_44576,N_41634);
nand UO_3089 (O_3089,N_45706,N_41964);
nand UO_3090 (O_3090,N_40952,N_46175);
nor UO_3091 (O_3091,N_45685,N_44060);
nand UO_3092 (O_3092,N_40142,N_44974);
and UO_3093 (O_3093,N_49473,N_49029);
and UO_3094 (O_3094,N_49008,N_44167);
nand UO_3095 (O_3095,N_43519,N_47657);
or UO_3096 (O_3096,N_44580,N_40924);
nand UO_3097 (O_3097,N_42263,N_45426);
or UO_3098 (O_3098,N_45668,N_46550);
or UO_3099 (O_3099,N_42843,N_44335);
nand UO_3100 (O_3100,N_40887,N_42661);
nor UO_3101 (O_3101,N_48584,N_49317);
xnor UO_3102 (O_3102,N_41622,N_49863);
nand UO_3103 (O_3103,N_45037,N_43875);
nor UO_3104 (O_3104,N_41036,N_47955);
and UO_3105 (O_3105,N_42543,N_43139);
or UO_3106 (O_3106,N_47863,N_46416);
nor UO_3107 (O_3107,N_46587,N_49815);
nand UO_3108 (O_3108,N_49673,N_44426);
nor UO_3109 (O_3109,N_48402,N_41992);
xnor UO_3110 (O_3110,N_44629,N_43463);
nand UO_3111 (O_3111,N_48914,N_45939);
nor UO_3112 (O_3112,N_42651,N_45306);
and UO_3113 (O_3113,N_41139,N_47296);
or UO_3114 (O_3114,N_44616,N_42546);
and UO_3115 (O_3115,N_43080,N_44289);
nor UO_3116 (O_3116,N_44583,N_47223);
nor UO_3117 (O_3117,N_46998,N_47021);
nand UO_3118 (O_3118,N_47555,N_44233);
and UO_3119 (O_3119,N_43436,N_42734);
nand UO_3120 (O_3120,N_42452,N_40593);
or UO_3121 (O_3121,N_47510,N_41302);
or UO_3122 (O_3122,N_48570,N_46868);
nand UO_3123 (O_3123,N_48577,N_41584);
nor UO_3124 (O_3124,N_44932,N_48665);
and UO_3125 (O_3125,N_46750,N_47292);
or UO_3126 (O_3126,N_40386,N_46831);
nor UO_3127 (O_3127,N_48787,N_40490);
and UO_3128 (O_3128,N_40784,N_44960);
and UO_3129 (O_3129,N_40380,N_42842);
and UO_3130 (O_3130,N_49711,N_44802);
or UO_3131 (O_3131,N_42577,N_40759);
nand UO_3132 (O_3132,N_45562,N_41893);
or UO_3133 (O_3133,N_47262,N_43807);
or UO_3134 (O_3134,N_42169,N_44433);
nor UO_3135 (O_3135,N_40060,N_46205);
nor UO_3136 (O_3136,N_47850,N_40374);
or UO_3137 (O_3137,N_42824,N_45533);
and UO_3138 (O_3138,N_45095,N_46016);
nor UO_3139 (O_3139,N_40345,N_46566);
nor UO_3140 (O_3140,N_41604,N_49223);
and UO_3141 (O_3141,N_40272,N_42386);
and UO_3142 (O_3142,N_45060,N_43650);
nand UO_3143 (O_3143,N_42732,N_42117);
nor UO_3144 (O_3144,N_47614,N_45255);
nand UO_3145 (O_3145,N_46994,N_40317);
nand UO_3146 (O_3146,N_48941,N_40730);
nand UO_3147 (O_3147,N_48717,N_42245);
nand UO_3148 (O_3148,N_44929,N_46829);
nand UO_3149 (O_3149,N_40520,N_40722);
nor UO_3150 (O_3150,N_40717,N_44219);
xnor UO_3151 (O_3151,N_40295,N_42902);
nor UO_3152 (O_3152,N_43023,N_43628);
and UO_3153 (O_3153,N_47451,N_45339);
or UO_3154 (O_3154,N_49945,N_49175);
xor UO_3155 (O_3155,N_44655,N_48768);
and UO_3156 (O_3156,N_45953,N_48243);
xor UO_3157 (O_3157,N_45949,N_47625);
and UO_3158 (O_3158,N_44073,N_46153);
and UO_3159 (O_3159,N_45166,N_40710);
or UO_3160 (O_3160,N_41834,N_42886);
xnor UO_3161 (O_3161,N_46348,N_40290);
nand UO_3162 (O_3162,N_42226,N_48917);
nor UO_3163 (O_3163,N_47999,N_44711);
nand UO_3164 (O_3164,N_47043,N_49927);
and UO_3165 (O_3165,N_48202,N_45803);
nor UO_3166 (O_3166,N_46655,N_40760);
nand UO_3167 (O_3167,N_45913,N_49991);
or UO_3168 (O_3168,N_44413,N_48848);
nand UO_3169 (O_3169,N_45355,N_46073);
nand UO_3170 (O_3170,N_48239,N_49672);
xor UO_3171 (O_3171,N_43889,N_44207);
nand UO_3172 (O_3172,N_49336,N_43903);
nand UO_3173 (O_3173,N_44348,N_42265);
and UO_3174 (O_3174,N_44015,N_43834);
xor UO_3175 (O_3175,N_43203,N_47613);
and UO_3176 (O_3176,N_46071,N_48073);
nand UO_3177 (O_3177,N_45513,N_42945);
or UO_3178 (O_3178,N_48473,N_40118);
nor UO_3179 (O_3179,N_43731,N_47443);
and UO_3180 (O_3180,N_45507,N_49074);
nand UO_3181 (O_3181,N_47290,N_43394);
nand UO_3182 (O_3182,N_45038,N_42539);
nor UO_3183 (O_3183,N_48790,N_44586);
nand UO_3184 (O_3184,N_45835,N_45360);
or UO_3185 (O_3185,N_40526,N_44959);
nand UO_3186 (O_3186,N_45978,N_42981);
nand UO_3187 (O_3187,N_44896,N_46617);
and UO_3188 (O_3188,N_45880,N_49380);
or UO_3189 (O_3189,N_41094,N_40506);
xor UO_3190 (O_3190,N_46237,N_43543);
and UO_3191 (O_3191,N_46920,N_49909);
or UO_3192 (O_3192,N_40419,N_46260);
xor UO_3193 (O_3193,N_43739,N_49780);
xnor UO_3194 (O_3194,N_49555,N_49467);
or UO_3195 (O_3195,N_48480,N_49099);
nand UO_3196 (O_3196,N_41897,N_40909);
nor UO_3197 (O_3197,N_40791,N_46120);
nor UO_3198 (O_3198,N_40930,N_42756);
nor UO_3199 (O_3199,N_41503,N_46292);
nand UO_3200 (O_3200,N_40234,N_48953);
or UO_3201 (O_3201,N_42697,N_42763);
xnor UO_3202 (O_3202,N_44520,N_49324);
xnor UO_3203 (O_3203,N_48683,N_44850);
nor UO_3204 (O_3204,N_41038,N_46660);
or UO_3205 (O_3205,N_48184,N_43420);
nand UO_3206 (O_3206,N_45859,N_40469);
nand UO_3207 (O_3207,N_48415,N_48640);
xor UO_3208 (O_3208,N_47795,N_45133);
nand UO_3209 (O_3209,N_41901,N_42964);
nand UO_3210 (O_3210,N_45059,N_49421);
nor UO_3211 (O_3211,N_46429,N_48608);
nor UO_3212 (O_3212,N_43426,N_46126);
nand UO_3213 (O_3213,N_49993,N_46060);
and UO_3214 (O_3214,N_46534,N_44488);
xor UO_3215 (O_3215,N_44914,N_44117);
xnor UO_3216 (O_3216,N_46008,N_46696);
and UO_3217 (O_3217,N_43674,N_42535);
xor UO_3218 (O_3218,N_44115,N_47426);
nor UO_3219 (O_3219,N_48709,N_44452);
and UO_3220 (O_3220,N_45102,N_42257);
nand UO_3221 (O_3221,N_41599,N_45518);
or UO_3222 (O_3222,N_40096,N_42192);
or UO_3223 (O_3223,N_45055,N_40937);
or UO_3224 (O_3224,N_48809,N_40927);
nand UO_3225 (O_3225,N_46154,N_43028);
nand UO_3226 (O_3226,N_41903,N_45201);
or UO_3227 (O_3227,N_45129,N_43101);
nand UO_3228 (O_3228,N_48657,N_44680);
xnor UO_3229 (O_3229,N_46850,N_41663);
xnor UO_3230 (O_3230,N_49825,N_47724);
and UO_3231 (O_3231,N_46875,N_43179);
and UO_3232 (O_3232,N_43887,N_49831);
or UO_3233 (O_3233,N_47683,N_40154);
nand UO_3234 (O_3234,N_43765,N_44080);
and UO_3235 (O_3235,N_43129,N_48298);
and UO_3236 (O_3236,N_44900,N_48149);
or UO_3237 (O_3237,N_45855,N_48167);
nor UO_3238 (O_3238,N_40701,N_42570);
nor UO_3239 (O_3239,N_48963,N_45745);
and UO_3240 (O_3240,N_42694,N_45150);
nor UO_3241 (O_3241,N_42898,N_47136);
nand UO_3242 (O_3242,N_48782,N_44923);
and UO_3243 (O_3243,N_48121,N_45069);
or UO_3244 (O_3244,N_40327,N_48960);
xnor UO_3245 (O_3245,N_41402,N_46942);
or UO_3246 (O_3246,N_49292,N_46984);
nor UO_3247 (O_3247,N_40378,N_40407);
nand UO_3248 (O_3248,N_44928,N_45235);
and UO_3249 (O_3249,N_43496,N_49628);
or UO_3250 (O_3250,N_48305,N_41846);
and UO_3251 (O_3251,N_48829,N_47782);
nor UO_3252 (O_3252,N_47104,N_43125);
nor UO_3253 (O_3253,N_40601,N_42525);
xnor UO_3254 (O_3254,N_43855,N_40245);
nor UO_3255 (O_3255,N_48588,N_43885);
nand UO_3256 (O_3256,N_45385,N_47588);
and UO_3257 (O_3257,N_40094,N_42967);
or UO_3258 (O_3258,N_47640,N_45818);
or UO_3259 (O_3259,N_40133,N_48904);
nor UO_3260 (O_3260,N_49914,N_46981);
nor UO_3261 (O_3261,N_43460,N_46946);
nor UO_3262 (O_3262,N_47635,N_44893);
and UO_3263 (O_3263,N_47577,N_44463);
nand UO_3264 (O_3264,N_46142,N_48831);
or UO_3265 (O_3265,N_48354,N_48490);
and UO_3266 (O_3266,N_47915,N_42513);
nor UO_3267 (O_3267,N_44861,N_43156);
xnor UO_3268 (O_3268,N_41124,N_41515);
and UO_3269 (O_3269,N_49730,N_41570);
xnor UO_3270 (O_3270,N_46739,N_45093);
or UO_3271 (O_3271,N_44072,N_41420);
nand UO_3272 (O_3272,N_43576,N_44353);
nor UO_3273 (O_3273,N_46099,N_43119);
nor UO_3274 (O_3274,N_47620,N_49032);
and UO_3275 (O_3275,N_45813,N_41193);
xnor UO_3276 (O_3276,N_49743,N_45009);
nor UO_3277 (O_3277,N_44715,N_43686);
and UO_3278 (O_3278,N_43776,N_40610);
and UO_3279 (O_3279,N_48901,N_48505);
and UO_3280 (O_3280,N_46351,N_45970);
nand UO_3281 (O_3281,N_49947,N_45545);
xnor UO_3282 (O_3282,N_48272,N_40591);
and UO_3283 (O_3283,N_41203,N_44271);
nor UO_3284 (O_3284,N_42336,N_41691);
nor UO_3285 (O_3285,N_44070,N_43515);
or UO_3286 (O_3286,N_49705,N_46647);
nor UO_3287 (O_3287,N_42204,N_48839);
xor UO_3288 (O_3288,N_48022,N_45345);
nand UO_3289 (O_3289,N_46687,N_47726);
and UO_3290 (O_3290,N_49531,N_48675);
nand UO_3291 (O_3291,N_49051,N_42465);
and UO_3292 (O_3292,N_49536,N_43972);
or UO_3293 (O_3293,N_45310,N_49669);
xor UO_3294 (O_3294,N_48699,N_46216);
xnor UO_3295 (O_3295,N_47175,N_49773);
or UO_3296 (O_3296,N_47502,N_40600);
and UO_3297 (O_3297,N_47279,N_48433);
nor UO_3298 (O_3298,N_42557,N_41603);
and UO_3299 (O_3299,N_44232,N_48682);
and UO_3300 (O_3300,N_40465,N_48320);
or UO_3301 (O_3301,N_47841,N_40998);
nand UO_3302 (O_3302,N_42619,N_49158);
xnor UO_3303 (O_3303,N_44606,N_44528);
and UO_3304 (O_3304,N_42888,N_45969);
nor UO_3305 (O_3305,N_47636,N_45101);
nand UO_3306 (O_3306,N_41202,N_43122);
or UO_3307 (O_3307,N_49485,N_44090);
nand UO_3308 (O_3308,N_49160,N_42161);
or UO_3309 (O_3309,N_46041,N_49328);
nand UO_3310 (O_3310,N_44794,N_42723);
or UO_3311 (O_3311,N_43453,N_46487);
nor UO_3312 (O_3312,N_45682,N_40084);
and UO_3313 (O_3313,N_41263,N_42483);
and UO_3314 (O_3314,N_48095,N_44383);
and UO_3315 (O_3315,N_48414,N_42669);
and UO_3316 (O_3316,N_42571,N_49505);
xor UO_3317 (O_3317,N_44204,N_43328);
nand UO_3318 (O_3318,N_48446,N_42494);
nor UO_3319 (O_3319,N_48329,N_48923);
nor UO_3320 (O_3320,N_47415,N_42905);
nor UO_3321 (O_3321,N_41562,N_42317);
or UO_3322 (O_3322,N_45908,N_43800);
and UO_3323 (O_3323,N_43613,N_46983);
and UO_3324 (O_3324,N_45299,N_49066);
or UO_3325 (O_3325,N_46229,N_46734);
or UO_3326 (O_3326,N_43715,N_47306);
nor UO_3327 (O_3327,N_49529,N_45366);
nor UO_3328 (O_3328,N_40020,N_47798);
nand UO_3329 (O_3329,N_45568,N_48031);
and UO_3330 (O_3330,N_42680,N_48814);
and UO_3331 (O_3331,N_40665,N_44507);
nand UO_3332 (O_3332,N_40004,N_49986);
xnor UO_3333 (O_3333,N_49072,N_44762);
nor UO_3334 (O_3334,N_42762,N_48088);
nor UO_3335 (O_3335,N_41390,N_41015);
nor UO_3336 (O_3336,N_48826,N_41993);
nor UO_3337 (O_3337,N_42012,N_44021);
and UO_3338 (O_3338,N_42029,N_46269);
nor UO_3339 (O_3339,N_48481,N_42569);
nand UO_3340 (O_3340,N_49656,N_45064);
xor UO_3341 (O_3341,N_48655,N_40065);
nor UO_3342 (O_3342,N_43517,N_47546);
or UO_3343 (O_3343,N_45915,N_46375);
nor UO_3344 (O_3344,N_45523,N_46781);
or UO_3345 (O_3345,N_44132,N_41276);
and UO_3346 (O_3346,N_49273,N_45191);
nand UO_3347 (O_3347,N_45615,N_45047);
or UO_3348 (O_3348,N_40504,N_47876);
nand UO_3349 (O_3349,N_48237,N_47902);
or UO_3350 (O_3350,N_43205,N_45886);
xor UO_3351 (O_3351,N_41014,N_41045);
nor UO_3352 (O_3352,N_40574,N_46851);
and UO_3353 (O_3353,N_40508,N_49256);
xnor UO_3354 (O_3354,N_41028,N_45302);
and UO_3355 (O_3355,N_41648,N_42071);
nor UO_3356 (O_3356,N_47400,N_43063);
or UO_3357 (O_3357,N_40619,N_48210);
nand UO_3358 (O_3358,N_45588,N_45097);
and UO_3359 (O_3359,N_42458,N_48611);
nor UO_3360 (O_3360,N_49045,N_46854);
nor UO_3361 (O_3361,N_40035,N_40515);
nand UO_3362 (O_3362,N_43382,N_47747);
nor UO_3363 (O_3363,N_42724,N_44212);
or UO_3364 (O_3364,N_48754,N_43703);
or UO_3365 (O_3365,N_40517,N_43734);
nand UO_3366 (O_3366,N_46924,N_43881);
nand UO_3367 (O_3367,N_43801,N_49084);
or UO_3368 (O_3368,N_46155,N_44874);
or UO_3369 (O_3369,N_47680,N_44367);
or UO_3370 (O_3370,N_47693,N_48289);
or UO_3371 (O_3371,N_44588,N_47820);
nor UO_3372 (O_3372,N_44703,N_43312);
or UO_3373 (O_3373,N_47579,N_45924);
and UO_3374 (O_3374,N_41919,N_49202);
nand UO_3375 (O_3375,N_49713,N_40434);
or UO_3376 (O_3376,N_43673,N_40156);
xnor UO_3377 (O_3377,N_49812,N_46692);
or UO_3378 (O_3378,N_46299,N_43853);
nor UO_3379 (O_3379,N_40350,N_42683);
nand UO_3380 (O_3380,N_47597,N_45782);
nand UO_3381 (O_3381,N_40865,N_44110);
nor UO_3382 (O_3382,N_42404,N_45647);
or UO_3383 (O_3383,N_42136,N_41549);
or UO_3384 (O_3384,N_43353,N_42616);
nor UO_3385 (O_3385,N_46789,N_43121);
or UO_3386 (O_3386,N_40534,N_41444);
nor UO_3387 (O_3387,N_41188,N_41582);
and UO_3388 (O_3388,N_42229,N_44823);
xor UO_3389 (O_3389,N_44258,N_40795);
or UO_3390 (O_3390,N_40844,N_46801);
nor UO_3391 (O_3391,N_48207,N_45197);
or UO_3392 (O_3392,N_47320,N_41805);
or UO_3393 (O_3393,N_41084,N_47932);
nand UO_3394 (O_3394,N_46075,N_44097);
nor UO_3395 (O_3395,N_47991,N_45392);
nand UO_3396 (O_3396,N_48125,N_48689);
nor UO_3397 (O_3397,N_49905,N_42786);
xnor UO_3398 (O_3398,N_49643,N_48779);
nor UO_3399 (O_3399,N_40856,N_49592);
nand UO_3400 (O_3400,N_42991,N_49188);
nor UO_3401 (O_3401,N_41291,N_44611);
and UO_3402 (O_3402,N_41160,N_46542);
xnor UO_3403 (O_3403,N_49607,N_42382);
and UO_3404 (O_3404,N_46283,N_40761);
or UO_3405 (O_3405,N_44453,N_47090);
nand UO_3406 (O_3406,N_49079,N_42490);
and UO_3407 (O_3407,N_41290,N_40497);
nor UO_3408 (O_3408,N_42353,N_44228);
or UO_3409 (O_3409,N_47532,N_46006);
or UO_3410 (O_3410,N_49630,N_40914);
nand UO_3411 (O_3411,N_47644,N_43633);
nor UO_3412 (O_3412,N_48335,N_47879);
and UO_3413 (O_3413,N_47377,N_46764);
nor UO_3414 (O_3414,N_41293,N_47653);
or UO_3415 (O_3415,N_46123,N_48109);
nor UO_3416 (O_3416,N_44679,N_45623);
or UO_3417 (O_3417,N_43646,N_46971);
xor UO_3418 (O_3418,N_40845,N_47575);
nand UO_3419 (O_3419,N_45959,N_45398);
xnor UO_3420 (O_3420,N_40372,N_42454);
xor UO_3421 (O_3421,N_40487,N_45808);
or UO_3422 (O_3422,N_41005,N_47662);
nand UO_3423 (O_3423,N_43619,N_46680);
nand UO_3424 (O_3424,N_49009,N_42720);
and UO_3425 (O_3425,N_40339,N_40165);
nor UO_3426 (O_3426,N_47045,N_47170);
nor UO_3427 (O_3427,N_47472,N_41370);
nor UO_3428 (O_3428,N_46585,N_43787);
or UO_3429 (O_3429,N_45673,N_49721);
nand UO_3430 (O_3430,N_46977,N_40161);
nor UO_3431 (O_3431,N_44502,N_49964);
xor UO_3432 (O_3432,N_41847,N_40471);
and UO_3433 (O_3433,N_49122,N_42211);
or UO_3434 (O_3434,N_40715,N_45550);
and UO_3435 (O_3435,N_44659,N_49580);
and UO_3436 (O_3436,N_43108,N_43759);
nand UO_3437 (O_3437,N_48048,N_43350);
nor UO_3438 (O_3438,N_40932,N_47935);
nand UO_3439 (O_3439,N_42063,N_45539);
nand UO_3440 (O_3440,N_46140,N_48866);
and UO_3441 (O_3441,N_46577,N_45981);
nand UO_3442 (O_3442,N_45436,N_45511);
and UO_3443 (O_3443,N_42180,N_48188);
xnor UO_3444 (O_3444,N_43825,N_43838);
or UO_3445 (O_3445,N_45972,N_45112);
and UO_3446 (O_3446,N_45990,N_43718);
xnor UO_3447 (O_3447,N_41879,N_41189);
nand UO_3448 (O_3448,N_45241,N_43542);
nand UO_3449 (O_3449,N_42312,N_45464);
or UO_3450 (O_3450,N_42004,N_48292);
nor UO_3451 (O_3451,N_42553,N_49779);
and UO_3452 (O_3452,N_47621,N_48327);
nand UO_3453 (O_3453,N_44903,N_43375);
or UO_3454 (O_3454,N_45512,N_49602);
nand UO_3455 (O_3455,N_40103,N_41093);
xor UO_3456 (O_3456,N_43389,N_43663);
or UO_3457 (O_3457,N_47762,N_49355);
and UO_3458 (O_3458,N_47271,N_45348);
nor UO_3459 (O_3459,N_40332,N_46162);
xor UO_3460 (O_3460,N_45617,N_42885);
nor UO_3461 (O_3461,N_49126,N_41916);
and UO_3462 (O_3462,N_45934,N_42862);
and UO_3463 (O_3463,N_48581,N_47804);
nand UO_3464 (O_3464,N_45996,N_48870);
nor UO_3465 (O_3465,N_47610,N_41361);
and UO_3466 (O_3466,N_47894,N_43793);
and UO_3467 (O_3467,N_44508,N_40686);
and UO_3468 (O_3468,N_44314,N_49427);
nor UO_3469 (O_3469,N_49156,N_45053);
nor UO_3470 (O_3470,N_41316,N_41171);
nor UO_3471 (O_3471,N_44098,N_45136);
xor UO_3472 (O_3472,N_40949,N_40521);
nand UO_3473 (O_3473,N_46897,N_40748);
nand UO_3474 (O_3474,N_43110,N_48802);
nand UO_3475 (O_3475,N_47432,N_41102);
or UO_3476 (O_3476,N_49832,N_45772);
or UO_3477 (O_3477,N_45182,N_40180);
and UO_3478 (O_3478,N_47557,N_46702);
xor UO_3479 (O_3479,N_48989,N_42910);
nor UO_3480 (O_3480,N_40195,N_42138);
nand UO_3481 (O_3481,N_40703,N_42439);
nor UO_3482 (O_3482,N_49992,N_40707);
xnor UO_3483 (O_3483,N_46374,N_45495);
and UO_3484 (O_3484,N_45279,N_42940);
nor UO_3485 (O_3485,N_45032,N_44119);
xnor UO_3486 (O_3486,N_42416,N_45040);
or UO_3487 (O_3487,N_45316,N_49771);
nand UO_3488 (O_3488,N_49967,N_49091);
or UO_3489 (O_3489,N_49425,N_41623);
or UO_3490 (O_3490,N_45148,N_41088);
or UO_3491 (O_3491,N_44646,N_41464);
or UO_3492 (O_3492,N_48132,N_47293);
and UO_3493 (O_3493,N_43228,N_44307);
nand UO_3494 (O_3494,N_40075,N_47508);
xor UO_3495 (O_3495,N_44557,N_47429);
nand UO_3496 (O_3496,N_49908,N_48430);
nand UO_3497 (O_3497,N_41279,N_48637);
nand UO_3498 (O_3498,N_44614,N_42008);
or UO_3499 (O_3499,N_42475,N_40616);
and UO_3500 (O_3500,N_44904,N_41488);
nand UO_3501 (O_3501,N_42909,N_46759);
and UO_3502 (O_3502,N_49676,N_49300);
xor UO_3503 (O_3503,N_49116,N_43193);
and UO_3504 (O_3504,N_43867,N_48404);
or UO_3505 (O_3505,N_44422,N_41007);
or UO_3506 (O_3506,N_49023,N_46893);
or UO_3507 (O_3507,N_49515,N_42706);
xnor UO_3508 (O_3508,N_47280,N_44972);
nor UO_3509 (O_3509,N_47029,N_42837);
or UO_3510 (O_3510,N_44598,N_49258);
and UO_3511 (O_3511,N_45189,N_45821);
xnor UO_3512 (O_3512,N_46900,N_48375);
nand UO_3513 (O_3513,N_43562,N_47813);
or UO_3514 (O_3514,N_45505,N_41652);
and UO_3515 (O_3515,N_49564,N_42476);
and UO_3516 (O_3516,N_42499,N_47181);
and UO_3517 (O_3517,N_40079,N_47242);
or UO_3518 (O_3518,N_40595,N_49457);
nor UO_3519 (O_3519,N_49020,N_44926);
nand UO_3520 (O_3520,N_49728,N_47478);
or UO_3521 (O_3521,N_47880,N_49982);
nand UO_3522 (O_3522,N_46281,N_49343);
and UO_3523 (O_3523,N_46090,N_44193);
xor UO_3524 (O_3524,N_45000,N_48463);
nor UO_3525 (O_3525,N_49655,N_43756);
xor UO_3526 (O_3526,N_44878,N_44981);
or UO_3527 (O_3527,N_46029,N_42383);
nor UO_3528 (O_3528,N_45569,N_48460);
and UO_3529 (O_3529,N_42498,N_42140);
nor UO_3530 (O_3530,N_44150,N_47543);
nor UO_3531 (O_3531,N_45365,N_48688);
or UO_3532 (O_3532,N_49873,N_42528);
and UO_3533 (O_3533,N_48597,N_41213);
or UO_3534 (O_3534,N_44095,N_45805);
nor UO_3535 (O_3535,N_46618,N_46657);
or UO_3536 (O_3536,N_44750,N_44654);
or UO_3537 (O_3537,N_47063,N_48013);
nand UO_3538 (O_3538,N_48278,N_48291);
nor UO_3539 (O_3539,N_40777,N_46038);
or UO_3540 (O_3540,N_47505,N_44705);
and UO_3541 (O_3541,N_41335,N_42415);
and UO_3542 (O_3542,N_44203,N_41673);
nor UO_3543 (O_3543,N_46675,N_40725);
or UO_3544 (O_3544,N_44444,N_41576);
nand UO_3545 (O_3545,N_44247,N_47794);
nor UO_3546 (O_3546,N_44640,N_43743);
and UO_3547 (O_3547,N_47612,N_46302);
nand UO_3548 (O_3548,N_40088,N_40558);
or UO_3549 (O_3549,N_47529,N_44933);
and UO_3550 (O_3550,N_47632,N_41979);
or UO_3551 (O_3551,N_41669,N_45099);
and UO_3552 (O_3552,N_47536,N_47051);
nor UO_3553 (O_3553,N_41814,N_40057);
nor UO_3554 (O_3554,N_48986,N_47507);
or UO_3555 (O_3555,N_41816,N_43072);
or UO_3556 (O_3556,N_42053,N_42610);
nor UO_3557 (O_3557,N_49373,N_47962);
nor UO_3558 (O_3558,N_46826,N_40864);
or UO_3559 (O_3559,N_41016,N_44142);
nor UO_3560 (O_3560,N_47495,N_42043);
or UO_3561 (O_3561,N_48258,N_40637);
nand UO_3562 (O_3562,N_48290,N_46097);
and UO_3563 (O_3563,N_49759,N_48160);
nand UO_3564 (O_3564,N_41106,N_41107);
and UO_3565 (O_3565,N_45980,N_49765);
or UO_3566 (O_3566,N_49362,N_41975);
and UO_3567 (O_3567,N_40127,N_47185);
xnor UO_3568 (O_3568,N_42896,N_41862);
nor UO_3569 (O_3569,N_41753,N_41566);
nand UO_3570 (O_3570,N_48486,N_48256);
nand UO_3571 (O_3571,N_49723,N_40901);
nor UO_3572 (O_3572,N_43341,N_40456);
or UO_3573 (O_3573,N_48645,N_44799);
nor UO_3574 (O_3574,N_40423,N_41421);
nor UO_3575 (O_3575,N_48065,N_47950);
or UO_3576 (O_3576,N_40427,N_44475);
or UO_3577 (O_3577,N_42956,N_43880);
nand UO_3578 (O_3578,N_47506,N_45882);
nand UO_3579 (O_3579,N_43918,N_48431);
nand UO_3580 (O_3580,N_47389,N_41734);
nand UO_3581 (O_3581,N_49867,N_47193);
and UO_3582 (O_3582,N_41994,N_47265);
nand UO_3583 (O_3583,N_42393,N_47821);
and UO_3584 (O_3584,N_44617,N_47745);
or UO_3585 (O_3585,N_40324,N_42994);
or UO_3586 (O_3586,N_40947,N_49483);
xor UO_3587 (O_3587,N_41394,N_47952);
or UO_3588 (O_3588,N_40408,N_46206);
or UO_3589 (O_3589,N_41086,N_48818);
or UO_3590 (O_3590,N_45477,N_49389);
or UO_3591 (O_3591,N_47383,N_42979);
nand UO_3592 (O_3592,N_48497,N_43837);
and UO_3593 (O_3593,N_40910,N_46885);
and UO_3594 (O_3594,N_43539,N_46628);
nand UO_3595 (O_3595,N_44179,N_45976);
nand UO_3596 (O_3596,N_45431,N_47731);
or UO_3597 (O_3597,N_42434,N_41327);
and UO_3598 (O_3598,N_44800,N_42322);
xor UO_3599 (O_3599,N_46480,N_41255);
nor UO_3600 (O_3600,N_49904,N_42748);
nand UO_3601 (O_3601,N_49542,N_40647);
nand UO_3602 (O_3602,N_45918,N_44168);
nand UO_3603 (O_3603,N_45450,N_40019);
and UO_3604 (O_3604,N_45483,N_46094);
and UO_3605 (O_3605,N_43554,N_49033);
nor UO_3606 (O_3606,N_41654,N_46921);
and UO_3607 (O_3607,N_49436,N_48861);
nor UO_3608 (O_3608,N_48493,N_44704);
xor UO_3609 (O_3609,N_46512,N_49366);
nand UO_3610 (O_3610,N_42010,N_45857);
nor UO_3611 (O_3611,N_44309,N_48617);
nor UO_3612 (O_3612,N_48863,N_44457);
xor UO_3613 (O_3613,N_48992,N_40953);
xor UO_3614 (O_3614,N_42913,N_41352);
and UO_3615 (O_3615,N_49142,N_42215);
nor UO_3616 (O_3616,N_43324,N_43749);
or UO_3617 (O_3617,N_42628,N_46891);
nand UO_3618 (O_3618,N_44604,N_48979);
nor UO_3619 (O_3619,N_49846,N_48059);
nand UO_3620 (O_3620,N_42206,N_48040);
and UO_3621 (O_3621,N_41892,N_46387);
and UO_3622 (O_3622,N_42333,N_44807);
xor UO_3623 (O_3623,N_49942,N_45560);
nand UO_3624 (O_3624,N_44363,N_41616);
and UO_3625 (O_3625,N_45565,N_46723);
xnor UO_3626 (O_3626,N_45861,N_45755);
nand UO_3627 (O_3627,N_40102,N_40316);
xnor UO_3628 (O_3628,N_46466,N_42789);
xor UO_3629 (O_3629,N_47244,N_40641);
nand UO_3630 (O_3630,N_44951,N_41469);
nor UO_3631 (O_3631,N_41493,N_45672);
nand UO_3632 (O_3632,N_43014,N_43407);
or UO_3633 (O_3633,N_45587,N_44804);
nor UO_3634 (O_3634,N_41313,N_41621);
and UO_3635 (O_3635,N_46319,N_40416);
or UO_3636 (O_3636,N_44151,N_48007);
nor UO_3637 (O_3637,N_46677,N_47335);
or UO_3638 (O_3638,N_47871,N_41073);
xnor UO_3639 (O_3639,N_46679,N_43682);
nor UO_3640 (O_3640,N_47481,N_46917);
or UO_3641 (O_3641,N_41546,N_47739);
or UO_3642 (O_3642,N_49333,N_41510);
or UO_3643 (O_3643,N_48112,N_45178);
and UO_3644 (O_3644,N_45141,N_46317);
and UO_3645 (O_3645,N_43414,N_49777);
nand UO_3646 (O_3646,N_46890,N_46896);
xor UO_3647 (O_3647,N_48943,N_45338);
nand UO_3648 (O_3648,N_45985,N_47471);
or UO_3649 (O_3649,N_42420,N_41506);
nor UO_3650 (O_3650,N_42105,N_46623);
or UO_3651 (O_3651,N_46425,N_46388);
and UO_3652 (O_3652,N_42305,N_47826);
or UO_3653 (O_3653,N_46978,N_42166);
or UO_3654 (O_3654,N_41764,N_45287);
and UO_3655 (O_3655,N_40925,N_42665);
nand UO_3656 (O_3656,N_48825,N_44004);
and UO_3657 (O_3657,N_46363,N_48812);
or UO_3658 (O_3658,N_40792,N_43933);
nand UO_3659 (O_3659,N_49471,N_48016);
and UO_3660 (O_3660,N_45439,N_41476);
and UO_3661 (O_3661,N_41348,N_47993);
nand UO_3662 (O_3662,N_48294,N_40529);
nand UO_3663 (O_3663,N_47068,N_46168);
or UO_3664 (O_3664,N_48482,N_44942);
or UO_3665 (O_3665,N_40877,N_40978);
nand UO_3666 (O_3666,N_49239,N_46491);
nand UO_3667 (O_3667,N_44514,N_44437);
nor UO_3668 (O_3668,N_42579,N_48300);
or UO_3669 (O_3669,N_44344,N_45070);
or UO_3670 (O_3670,N_49852,N_49310);
and UO_3671 (O_3671,N_44790,N_43360);
or UO_3672 (O_3672,N_42157,N_40401);
or UO_3673 (O_3673,N_40185,N_43507);
nor UO_3674 (O_3674,N_45977,N_40442);
xnor UO_3675 (O_3675,N_41645,N_48778);
nor UO_3676 (O_3676,N_43009,N_48503);
or UO_3677 (O_3677,N_49541,N_44040);
xor UO_3678 (O_3678,N_40961,N_43693);
nor UO_3679 (O_3679,N_47840,N_45785);
nand UO_3680 (O_3680,N_40258,N_46423);
nor UO_3681 (O_3681,N_41746,N_43094);
or UO_3682 (O_3682,N_41321,N_47831);
or UO_3683 (O_3683,N_46684,N_42479);
or UO_3684 (O_3684,N_44822,N_43393);
and UO_3685 (O_3685,N_42686,N_40672);
and UO_3686 (O_3686,N_41995,N_45841);
xnor UO_3687 (O_3687,N_40362,N_43284);
nor UO_3688 (O_3688,N_41380,N_48023);
and UO_3689 (O_3689,N_45227,N_40738);
xnor UO_3690 (O_3690,N_41585,N_47493);
xnor UO_3691 (O_3691,N_47521,N_43344);
and UO_3692 (O_3692,N_48378,N_43443);
nor UO_3693 (O_3693,N_46544,N_43843);
or UO_3694 (O_3694,N_47904,N_47818);
nor UO_3695 (O_3695,N_48113,N_49928);
or UO_3696 (O_3696,N_43183,N_48362);
and UO_3697 (O_3697,N_45557,N_45353);
nor UO_3698 (O_3698,N_43435,N_44786);
or UO_3699 (O_3699,N_44727,N_46327);
xnor UO_3700 (O_3700,N_49411,N_41262);
and UO_3701 (O_3701,N_47060,N_47700);
and UO_3702 (O_3702,N_46483,N_46856);
or UO_3703 (O_3703,N_49634,N_42361);
and UO_3704 (O_3704,N_40690,N_48219);
and UO_3705 (O_3705,N_44494,N_46563);
nand UO_3706 (O_3706,N_48094,N_41200);
and UO_3707 (O_3707,N_43377,N_46305);
nor UO_3708 (O_3708,N_44403,N_45767);
nand UO_3709 (O_3709,N_45989,N_48205);
or UO_3710 (O_3710,N_42650,N_40890);
nand UO_3711 (O_3711,N_48119,N_45087);
or UO_3712 (O_3712,N_45384,N_46170);
or UO_3713 (O_3713,N_42324,N_40254);
nor UO_3714 (O_3714,N_40589,N_41889);
and UO_3715 (O_3715,N_46131,N_42526);
nor UO_3716 (O_3716,N_41855,N_46235);
and UO_3717 (O_3717,N_40414,N_47643);
and UO_3718 (O_3718,N_46622,N_42873);
or UO_3719 (O_3719,N_44106,N_41896);
nand UO_3720 (O_3720,N_42418,N_45187);
nand UO_3721 (O_3721,N_42690,N_46065);
nor UO_3722 (O_3722,N_49403,N_43544);
nor UO_3723 (O_3723,N_49254,N_40880);
and UO_3724 (O_3724,N_44675,N_41475);
nor UO_3725 (O_3725,N_48295,N_47956);
nand UO_3726 (O_3726,N_41442,N_47972);
nand UO_3727 (O_3727,N_48824,N_44492);
nor UO_3728 (O_3728,N_42652,N_44706);
nand UO_3729 (O_3729,N_46381,N_49553);
nand UO_3730 (O_3730,N_44963,N_41703);
and UO_3731 (O_3731,N_45132,N_48273);
or UO_3732 (O_3732,N_45406,N_46798);
and UO_3733 (O_3733,N_47297,N_43273);
and UO_3734 (O_3734,N_42536,N_49476);
or UO_3735 (O_3735,N_42693,N_48314);
and UO_3736 (O_3736,N_45358,N_49956);
nand UO_3737 (O_3737,N_40552,N_44648);
nor UO_3738 (O_3738,N_43178,N_45960);
or UO_3739 (O_3739,N_46111,N_47771);
and UO_3740 (O_3740,N_40577,N_40237);
nor UO_3741 (O_3741,N_41865,N_47801);
nand UO_3742 (O_3742,N_47130,N_42034);
xor UO_3743 (O_3743,N_43706,N_40984);
nand UO_3744 (O_3744,N_44647,N_43055);
nor UO_3745 (O_3745,N_45606,N_40250);
xnor UO_3746 (O_3746,N_49261,N_44758);
or UO_3747 (O_3747,N_42625,N_44880);
and UO_3748 (O_3748,N_43391,N_46941);
nand UO_3749 (O_3749,N_49085,N_44907);
or UO_3750 (O_3750,N_49190,N_45394);
and UO_3751 (O_3751,N_46873,N_42537);
or UO_3752 (O_3752,N_42401,N_42428);
xor UO_3753 (O_3753,N_43587,N_44540);
nand UO_3754 (O_3754,N_42959,N_40486);
nand UO_3755 (O_3755,N_41381,N_41310);
and UO_3756 (O_3756,N_45225,N_42127);
or UO_3757 (O_3757,N_42908,N_40385);
nor UO_3758 (O_3758,N_43505,N_41286);
nand UO_3759 (O_3759,N_47076,N_42468);
and UO_3760 (O_3760,N_40990,N_42541);
and UO_3761 (O_3761,N_43548,N_42032);
nand UO_3762 (O_3762,N_48419,N_45264);
nand UO_3763 (O_3763,N_46106,N_46199);
nand UO_3764 (O_3764,N_41518,N_44911);
and UO_3765 (O_3765,N_49138,N_48093);
nand UO_3766 (O_3766,N_44226,N_42332);
nand UO_3767 (O_3767,N_44718,N_48240);
nand UO_3768 (O_3768,N_45607,N_42626);
nand UO_3769 (O_3769,N_46909,N_42573);
and UO_3770 (O_3770,N_40056,N_41006);
nand UO_3771 (O_3771,N_43893,N_40046);
nand UO_3772 (O_3772,N_45326,N_43607);
xnor UO_3773 (O_3773,N_44852,N_48337);
or UO_3774 (O_3774,N_42019,N_40850);
or UO_3775 (O_3775,N_47886,N_41047);
nand UO_3776 (O_3776,N_43777,N_42591);
nor UO_3777 (O_3777,N_46004,N_49161);
and UO_3778 (O_3778,N_47608,N_40166);
and UO_3779 (O_3779,N_46226,N_41878);
and UO_3780 (O_3780,N_42104,N_40398);
nand UO_3781 (O_3781,N_44154,N_45747);
or UO_3782 (O_3782,N_48247,N_41299);
nand UO_3783 (O_3783,N_45057,N_43915);
or UO_3784 (O_3784,N_42425,N_47168);
or UO_3785 (O_3785,N_41037,N_48985);
and UO_3786 (O_3786,N_49322,N_43704);
and UO_3787 (O_3787,N_46232,N_43427);
nor UO_3788 (O_3788,N_44554,N_42949);
xnor UO_3789 (O_3789,N_44901,N_49028);
nand UO_3790 (O_3790,N_43632,N_47476);
or UO_3791 (O_3791,N_43403,N_42627);
nor UO_3792 (O_3792,N_43136,N_42995);
nand UO_3793 (O_3793,N_42769,N_48215);
nand UO_3794 (O_3794,N_40045,N_47544);
and UO_3795 (O_3795,N_41594,N_41572);
or UO_3796 (O_3796,N_46737,N_40183);
nor UO_3797 (O_3797,N_48353,N_41522);
nor UO_3798 (O_3798,N_40979,N_41311);
and UO_3799 (O_3799,N_47525,N_43878);
nand UO_3800 (O_3800,N_49557,N_42840);
and UO_3801 (O_3801,N_42687,N_45516);
nor UO_3802 (O_3802,N_42174,N_47020);
or UO_3803 (O_3803,N_49039,N_43406);
xor UO_3804 (O_3804,N_42924,N_42758);
or UO_3805 (O_3805,N_42941,N_44441);
nand UO_3806 (O_3806,N_42241,N_40355);
xnor UO_3807 (O_3807,N_41832,N_44257);
or UO_3808 (O_3808,N_41053,N_42313);
nor UO_3809 (O_3809,N_43920,N_40516);
nor UO_3810 (O_3810,N_44975,N_40076);
and UO_3811 (O_3811,N_47590,N_47791);
nor UO_3812 (O_3812,N_43259,N_43343);
nor UO_3813 (O_3813,N_48015,N_48740);
nor UO_3814 (O_3814,N_44824,N_48137);
xnor UO_3815 (O_3815,N_49477,N_45050);
nor UO_3816 (O_3816,N_43310,N_47691);
or UO_3817 (O_3817,N_46664,N_45117);
nand UO_3818 (O_3818,N_43973,N_43999);
or UO_3819 (O_3819,N_40248,N_49235);
nand UO_3820 (O_3820,N_40536,N_46149);
nand UO_3821 (O_3821,N_46603,N_44479);
and UO_3822 (O_3822,N_48153,N_45616);
and UO_3823 (O_3823,N_47735,N_49620);
xnor UO_3824 (O_3824,N_43388,N_43348);
xnor UO_3825 (O_3825,N_48906,N_43872);
xnor UO_3826 (O_3826,N_46461,N_41581);
nor UO_3827 (O_3827,N_48819,N_44978);
nor UO_3828 (O_3828,N_46243,N_45207);
xor UO_3829 (O_3829,N_46357,N_46610);
nand UO_3830 (O_3830,N_42636,N_45499);
or UO_3831 (O_3831,N_45948,N_45522);
nor UO_3832 (O_3832,N_43301,N_42198);
nor UO_3833 (O_3833,N_49690,N_46778);
nand UO_3834 (O_3834,N_48690,N_42079);
nand UO_3835 (O_3835,N_47748,N_44801);
and UO_3836 (O_3836,N_49604,N_47979);
and UO_3837 (O_3837,N_42817,N_45205);
and UO_3838 (O_3838,N_48330,N_46062);
xnor UO_3839 (O_3839,N_49013,N_46105);
nand UO_3840 (O_3840,N_47190,N_45837);
nand UO_3841 (O_3841,N_49384,N_48371);
nor UO_3842 (O_3842,N_43295,N_45891);
nand UO_3843 (O_3843,N_44135,N_42330);
nor UO_3844 (O_3844,N_48123,N_40371);
nand UO_3845 (O_3845,N_43799,N_44411);
and UO_3846 (O_3846,N_44141,N_45854);
nor UO_3847 (O_3847,N_49289,N_43354);
nand UO_3848 (O_3848,N_49703,N_47142);
xor UO_3849 (O_3849,N_40734,N_47699);
or UO_3850 (O_3850,N_47702,N_44401);
or UO_3851 (O_3851,N_47378,N_45717);
xnor UO_3852 (O_3852,N_41788,N_41143);
or UO_3853 (O_3853,N_45409,N_41574);
or UO_3854 (O_3854,N_44934,N_49128);
and UO_3855 (O_3855,N_41751,N_47009);
or UO_3856 (O_3856,N_44041,N_47070);
nand UO_3857 (O_3857,N_45724,N_46460);
xor UO_3858 (O_3858,N_41432,N_44049);
nor UO_3859 (O_3859,N_48652,N_41928);
or UO_3860 (O_3860,N_48974,N_49042);
and UO_3861 (O_3861,N_40373,N_45734);
or UO_3862 (O_3862,N_42701,N_49407);
and UO_3863 (O_3863,N_48260,N_46259);
nor UO_3864 (O_3864,N_48910,N_42308);
nor UO_3865 (O_3865,N_40997,N_47098);
or UO_3866 (O_3866,N_45122,N_40907);
and UO_3867 (O_3867,N_45008,N_48224);
nand UO_3868 (O_3868,N_42410,N_48227);
nand UO_3869 (O_3869,N_44906,N_40835);
or UO_3870 (O_3870,N_40134,N_48990);
nand UO_3871 (O_3871,N_49327,N_46543);
and UO_3872 (O_3872,N_49323,N_48196);
or UO_3873 (O_3873,N_45303,N_48525);
or UO_3874 (O_3874,N_45401,N_45559);
and UO_3875 (O_3875,N_45701,N_40731);
nand UO_3876 (O_3876,N_45567,N_45683);
or UO_3877 (O_3877,N_49872,N_46083);
nor UO_3878 (O_3878,N_43631,N_45626);
nand UO_3879 (O_3879,N_42181,N_42422);
and UO_3880 (O_3880,N_41404,N_42402);
nand UO_3881 (O_3881,N_44855,N_44669);
or UO_3882 (O_3882,N_45885,N_49308);
or UO_3883 (O_3883,N_48735,N_43188);
or UO_3884 (O_3884,N_49623,N_44661);
and UO_3885 (O_3885,N_44970,N_46404);
or UO_3886 (O_3886,N_44382,N_48626);
nand UO_3887 (O_3887,N_43761,N_42108);
xnor UO_3888 (O_3888,N_41428,N_46124);
nor UO_3889 (O_3889,N_48697,N_40673);
xnor UO_3890 (O_3890,N_41161,N_48143);
or UO_3891 (O_3891,N_42755,N_47627);
nor UO_3892 (O_3892,N_41317,N_49929);
nand UO_3893 (O_3893,N_47276,N_49921);
and UO_3894 (O_3894,N_48293,N_41923);
nand UO_3895 (O_3895,N_46539,N_43171);
and UO_3896 (O_3896,N_48798,N_44495);
and UO_3897 (O_3897,N_41759,N_48257);
nand UO_3898 (O_3898,N_44454,N_41831);
nand UO_3899 (O_3899,N_47200,N_41789);
and UO_3900 (O_3900,N_48467,N_48969);
nand UO_3901 (O_3901,N_42516,N_41723);
and UO_3902 (O_3902,N_41996,N_44338);
and UO_3903 (O_3903,N_44123,N_48412);
or UO_3904 (O_3904,N_41039,N_43266);
or UO_3905 (O_3905,N_43568,N_44809);
nand UO_3906 (O_3906,N_46394,N_42302);
nor UO_3907 (O_3907,N_47732,N_45780);
or UO_3908 (O_3908,N_48530,N_46242);
or UO_3909 (O_3909,N_48921,N_41732);
nor UO_3910 (O_3910,N_47545,N_48656);
nor UO_3911 (O_3911,N_42700,N_41858);
nand UO_3912 (O_3912,N_45011,N_43817);
or UO_3913 (O_3913,N_49237,N_45214);
xor UO_3914 (O_3914,N_49082,N_43081);
or UO_3915 (O_3915,N_40461,N_46103);
nor UO_3916 (O_3916,N_42001,N_42264);
nand UO_3917 (O_3917,N_49797,N_40038);
nand UO_3918 (O_3918,N_46107,N_42872);
nor UO_3919 (O_3919,N_41241,N_41625);
xor UO_3920 (O_3920,N_44517,N_44832);
xor UO_3921 (O_3921,N_42128,N_47573);
and UO_3922 (O_3922,N_47559,N_40905);
nand UO_3923 (O_3923,N_41474,N_42631);
nor UO_3924 (O_3924,N_49749,N_40217);
nor UO_3925 (O_3925,N_43931,N_47152);
nor UO_3926 (O_3926,N_46128,N_48912);
nand UO_3927 (O_3927,N_46493,N_44450);
or UO_3928 (O_3928,N_42002,N_43379);
nand UO_3929 (O_3929,N_43033,N_43396);
nand UO_3930 (O_3930,N_43050,N_40939);
nand UO_3931 (O_3931,N_45910,N_41857);
nor UO_3932 (O_3932,N_42832,N_43858);
and UO_3933 (O_3933,N_44260,N_46451);
and UO_3934 (O_3934,N_46179,N_43928);
nor UO_3935 (O_3935,N_49369,N_40012);
xnor UO_3936 (O_3936,N_48024,N_48700);
nand UO_3937 (O_3937,N_47888,N_40293);
nand UO_3938 (O_3938,N_45367,N_47331);
and UO_3939 (O_3939,N_42209,N_42365);
and UO_3940 (O_3940,N_47284,N_46438);
nand UO_3941 (O_3941,N_42064,N_44417);
nor UO_3942 (O_3942,N_43593,N_41438);
and UO_3943 (O_3943,N_49893,N_41955);
nor UO_3944 (O_3944,N_46857,N_43932);
or UO_3945 (O_3945,N_40775,N_46760);
nand UO_3946 (O_3946,N_40225,N_41389);
or UO_3947 (O_3947,N_49157,N_49004);
or UO_3948 (O_3948,N_45937,N_42254);
nor UO_3949 (O_3949,N_48838,N_43757);
xnor UO_3950 (O_3950,N_41804,N_48833);
xor UO_3951 (O_3951,N_41035,N_49854);
nor UO_3952 (O_3952,N_46498,N_47667);
nand UO_3953 (O_3953,N_43639,N_44864);
nand UO_3954 (O_3954,N_41758,N_40235);
or UO_3955 (O_3955,N_41209,N_44651);
nor UO_3956 (O_3956,N_40883,N_46434);
or UO_3957 (O_3957,N_43004,N_45061);
nor UO_3958 (O_3958,N_43727,N_49347);
nand UO_3959 (O_3959,N_46333,N_42347);
or UO_3960 (O_3960,N_44490,N_46024);
nand UO_3961 (O_3961,N_46485,N_40675);
xnor UO_3962 (O_3962,N_47750,N_47301);
and UO_3963 (O_3963,N_48218,N_43655);
nand UO_3964 (O_3964,N_42667,N_44890);
and UO_3965 (O_3965,N_40130,N_47456);
and UO_3966 (O_3966,N_46366,N_48076);
and UO_3967 (O_3967,N_49330,N_44056);
and UO_3968 (O_3968,N_44332,N_49766);
nor UO_3969 (O_3969,N_49933,N_45085);
nand UO_3970 (O_3970,N_45346,N_46670);
nand UO_3971 (O_3971,N_43246,N_43118);
nand UO_3972 (O_3972,N_46129,N_47883);
or UO_3973 (O_3973,N_45229,N_45794);
and UO_3974 (O_3974,N_46122,N_47875);
and UO_3975 (O_3975,N_40093,N_41164);
and UO_3976 (O_3976,N_44352,N_41017);
and UO_3977 (O_3977,N_41127,N_49527);
or UO_3978 (O_3978,N_40492,N_41069);
or UO_3979 (O_3979,N_49372,N_46045);
nand UO_3980 (O_3980,N_45903,N_40252);
nand UO_3981 (O_3981,N_42639,N_43048);
xor UO_3982 (O_3982,N_48531,N_47947);
or UO_3983 (O_3983,N_49251,N_46898);
or UO_3984 (O_3984,N_41122,N_43506);
nand UO_3985 (O_3985,N_40009,N_41051);
nand UO_3986 (O_3986,N_45768,N_45975);
or UO_3987 (O_3987,N_44263,N_49821);
and UO_3988 (O_3988,N_47654,N_44269);
nand UO_3989 (O_3989,N_47910,N_41848);
nor UO_3990 (O_3990,N_41525,N_40971);
nor UO_3991 (O_3991,N_42346,N_49272);
and UO_3992 (O_3992,N_47833,N_47539);
or UO_3993 (O_3993,N_44863,N_41597);
nand UO_3994 (O_3994,N_45889,N_48693);
nor UO_3995 (O_3995,N_45543,N_40450);
nand UO_3996 (O_3996,N_40129,N_44740);
or UO_3997 (O_3997,N_45263,N_44120);
or UO_3998 (O_3998,N_47716,N_44575);
or UO_3999 (O_3999,N_46910,N_42450);
nand UO_4000 (O_4000,N_48747,N_49594);
or UO_4001 (O_4001,N_47814,N_43124);
nor UO_4002 (O_4002,N_47646,N_41757);
nor UO_4003 (O_4003,N_46990,N_40015);
nand UO_4004 (O_4004,N_47706,N_44163);
or UO_4005 (O_4005,N_44292,N_41494);
nor UO_4006 (O_4006,N_43753,N_43905);
nor UO_4007 (O_4007,N_40702,N_49162);
nand UO_4008 (O_4008,N_46166,N_49262);
nand UO_4009 (O_4009,N_46143,N_41235);
nand UO_4010 (O_4010,N_46413,N_49253);
nor UO_4011 (O_4011,N_42214,N_47906);
and UO_4012 (O_4012,N_40885,N_41250);
xor UO_4013 (O_4013,N_41207,N_49735);
and UO_4014 (O_4014,N_45124,N_40083);
and UO_4015 (O_4015,N_42688,N_41344);
or UO_4016 (O_4016,N_48628,N_44516);
or UO_4017 (O_4017,N_41619,N_42939);
nand UO_4018 (O_4018,N_40823,N_48572);
xnor UO_4019 (O_4019,N_46136,N_46033);
nand UO_4020 (O_4020,N_47202,N_44033);
or UO_4021 (O_4021,N_47388,N_49601);
or UO_4022 (O_4022,N_48635,N_44590);
nand UO_4023 (O_4023,N_44681,N_46241);
and UO_4024 (O_4024,N_46607,N_42162);
or UO_4025 (O_4025,N_41448,N_46668);
or UO_4026 (O_4026,N_46666,N_41166);
nor UO_4027 (O_4027,N_41944,N_43447);
nor UO_4028 (O_4028,N_48981,N_49521);
or UO_4029 (O_4029,N_40870,N_46661);
nor UO_4030 (O_4030,N_41977,N_42080);
and UO_4031 (O_4031,N_45465,N_45184);
nand UO_4032 (O_4032,N_47179,N_42460);
or UO_4033 (O_4033,N_47198,N_40816);
or UO_4034 (O_4034,N_43806,N_49801);
xnor UO_4035 (O_4035,N_47140,N_40278);
and UO_4036 (O_4036,N_41523,N_42950);
nand UO_4037 (O_4037,N_44641,N_48061);
nand UO_4038 (O_4038,N_43132,N_41512);
or UO_4039 (O_4039,N_44924,N_40284);
nor UO_4040 (O_4040,N_40753,N_45446);
xor UO_4041 (O_4041,N_47255,N_49281);
nand UO_4042 (O_4042,N_44397,N_42089);
or UO_4043 (O_4043,N_45457,N_43788);
or UO_4044 (O_4044,N_45723,N_47266);
and UO_4045 (O_4045,N_47603,N_41866);
nand UO_4046 (O_4046,N_45614,N_47427);
xnor UO_4047 (O_4047,N_43331,N_43380);
nor UO_4048 (O_4048,N_41677,N_41018);
nor UO_4049 (O_4049,N_46591,N_49031);
xnor UO_4050 (O_4050,N_41131,N_47989);
nand UO_4051 (O_4051,N_49948,N_46390);
and UO_4052 (O_4052,N_45756,N_43082);
nor UO_4053 (O_4053,N_48538,N_49257);
nand UO_4054 (O_4054,N_47601,N_46586);
nor UO_4055 (O_4055,N_43892,N_41130);
nand UO_4056 (O_4056,N_44887,N_45476);
nand UO_4057 (O_4057,N_49836,N_43811);
xor UO_4058 (O_4058,N_47519,N_46773);
or UO_4059 (O_4059,N_42328,N_42502);
nor UO_4060 (O_4060,N_49808,N_41315);
and UO_4061 (O_4061,N_42011,N_41407);
or UO_4062 (O_4062,N_47868,N_40808);
xnor UO_4063 (O_4063,N_49975,N_44674);
nor UO_4064 (O_4064,N_44764,N_49627);
and UO_4065 (O_4065,N_45661,N_48776);
and UO_4066 (O_4066,N_42344,N_47376);
or UO_4067 (O_4067,N_40006,N_42753);
and UO_4068 (O_4068,N_42159,N_45863);
and UO_4069 (O_4069,N_43929,N_46710);
or UO_4070 (O_4070,N_43695,N_41987);
nor UO_4071 (O_4071,N_47723,N_43751);
nor UO_4072 (O_4072,N_47802,N_40755);
nand UO_4073 (O_4073,N_45318,N_48545);
nand UO_4074 (O_4074,N_48037,N_47936);
or UO_4075 (O_4075,N_40975,N_42883);
nand UO_4076 (O_4076,N_44027,N_41149);
and UO_4077 (O_4077,N_44619,N_42674);
or UO_4078 (O_4078,N_47448,N_44857);
and UO_4079 (O_4079,N_47118,N_42733);
nand UO_4080 (O_4080,N_42277,N_43130);
and UO_4081 (O_4081,N_45624,N_45470);
xor UO_4082 (O_4082,N_49729,N_45123);
nand UO_4083 (O_4083,N_48107,N_44691);
and UO_4084 (O_4084,N_40432,N_42770);
or UO_4085 (O_4085,N_40190,N_43468);
and UO_4086 (O_4086,N_49913,N_47114);
xnor UO_4087 (O_4087,N_48561,N_48156);
nor UO_4088 (O_4088,N_41504,N_46717);
nor UO_4089 (O_4089,N_47757,N_44613);
or UO_4090 (O_4090,N_48749,N_45198);
nand UO_4091 (O_4091,N_46517,N_45604);
and UO_4092 (O_4092,N_43512,N_46497);
nor UO_4093 (O_4093,N_47317,N_47760);
nor UO_4094 (O_4094,N_46867,N_49182);
and UO_4095 (O_4095,N_49027,N_49994);
nor UO_4096 (O_4096,N_46631,N_49667);
and UO_4097 (O_4097,N_40322,N_47634);
nor UO_4098 (O_4098,N_41662,N_48803);
nor UO_4099 (O_4099,N_48429,N_44420);
nand UO_4100 (O_4100,N_45107,N_46636);
and UO_4101 (O_4101,N_48789,N_46362);
nand UO_4102 (O_4102,N_44239,N_43251);
nor UO_4103 (O_4103,N_40832,N_48230);
xnor UO_4104 (O_4104,N_49907,N_43922);
and UO_4105 (O_4105,N_46608,N_41880);
or UO_4106 (O_4106,N_42642,N_46397);
nand UO_4107 (O_4107,N_43944,N_48642);
nand UO_4108 (O_4108,N_41643,N_45266);
and UO_4109 (O_4109,N_48448,N_48241);
nand UO_4110 (O_4110,N_45240,N_48821);
xor UO_4111 (O_4111,N_40194,N_45163);
or UO_4112 (O_4112,N_48598,N_41940);
or UO_4113 (O_4113,N_44224,N_49709);
or UO_4114 (O_4114,N_46937,N_43433);
nor UO_4115 (O_4115,N_44312,N_40677);
and UO_4116 (O_4116,N_49830,N_48466);
and UO_4117 (O_4117,N_49406,N_40181);
nand UO_4118 (O_4118,N_46952,N_43467);
or UO_4119 (O_4119,N_43614,N_49277);
nand UO_4120 (O_4120,N_49900,N_49385);
or UO_4121 (O_4121,N_44318,N_47997);
or UO_4122 (O_4122,N_49413,N_48098);
xnor UO_4123 (O_4123,N_46933,N_45528);
or UO_4124 (O_4124,N_49848,N_46974);
nand UO_4125 (O_4125,N_45576,N_45012);
nand UO_4126 (O_4126,N_48138,N_47963);
nand UO_4127 (O_4127,N_45790,N_44676);
and UO_4128 (O_4128,N_49559,N_43311);
and UO_4129 (O_4129,N_41357,N_41458);
nor UO_4130 (O_4130,N_45630,N_48236);
nand UO_4131 (O_4131,N_48288,N_41332);
and UO_4132 (O_4132,N_43069,N_44602);
or UO_4133 (O_4133,N_40437,N_43711);
nor UO_4134 (O_4134,N_43983,N_49495);
or UO_4135 (O_4135,N_41031,N_45572);
and UO_4136 (O_4136,N_45109,N_45807);
or UO_4137 (O_4137,N_41050,N_40024);
or UO_4138 (O_4138,N_47907,N_48686);
or UO_4139 (O_4139,N_49587,N_47881);
nand UO_4140 (O_4140,N_42980,N_48304);
and UO_4141 (O_4141,N_49255,N_43638);
xor UO_4142 (O_4142,N_45517,N_44509);
nand UO_4143 (O_4143,N_41935,N_45596);
xor UO_4144 (O_4144,N_42878,N_49850);
nand UO_4145 (O_4145,N_49686,N_49275);
and UO_4146 (O_4146,N_46386,N_48636);
nor UO_4147 (O_4147,N_49708,N_48786);
xnor UO_4148 (O_4148,N_40280,N_43841);
nor UO_4149 (O_4149,N_44220,N_48091);
or UO_4150 (O_4150,N_42077,N_43007);
or UO_4151 (O_4151,N_42274,N_46541);
nor UO_4152 (O_4152,N_47985,N_42725);
and UO_4153 (O_4153,N_46520,N_45847);
or UO_4154 (O_4154,N_40002,N_44984);
or UO_4155 (O_4155,N_41055,N_40988);
nand UO_4156 (O_4156,N_47268,N_40320);
or UO_4157 (O_4157,N_41337,N_42811);
or UO_4158 (O_4158,N_41692,N_45013);
nor UO_4159 (O_4159,N_47023,N_40896);
or UO_4160 (O_4160,N_42061,N_42989);
nand UO_4161 (O_4161,N_48515,N_46428);
or UO_4162 (O_4162,N_41163,N_44752);
or UO_4163 (O_4163,N_48889,N_46881);
or UO_4164 (O_4164,N_43070,N_43952);
xor UO_4165 (O_4165,N_41201,N_49584);
and UO_4166 (O_4166,N_45440,N_45051);
and UO_4167 (O_4167,N_44394,N_42148);
xnor UO_4168 (O_4168,N_48520,N_42442);
nand UO_4169 (O_4169,N_42797,N_49298);
xor UO_4170 (O_4170,N_48324,N_49350);
or UO_4171 (O_4171,N_47129,N_46002);
and UO_4172 (O_4172,N_41181,N_42882);
nand UO_4173 (O_4173,N_40719,N_49054);
or UO_4174 (O_4174,N_49286,N_43672);
nor UO_4175 (O_4175,N_44767,N_40052);
or UO_4176 (O_4176,N_48027,N_40137);
or UO_4177 (O_4177,N_42179,N_41132);
and UO_4178 (O_4178,N_48997,N_41541);
or UO_4179 (O_4179,N_49633,N_40498);
or UO_4180 (O_4180,N_43347,N_43953);
nor UO_4181 (O_4181,N_40193,N_46208);
and UO_4182 (O_4182,N_43021,N_47087);
xnor UO_4183 (O_4183,N_49736,N_46057);
and UO_4184 (O_4184,N_47687,N_42168);
and UO_4185 (O_4185,N_48472,N_42906);
and UO_4186 (O_4186,N_43653,N_46437);
or UO_4187 (O_4187,N_48044,N_41115);
and UO_4188 (O_4188,N_45632,N_49888);
and UO_4189 (O_4189,N_42822,N_46654);
or UO_4190 (O_4190,N_46182,N_48723);
nor UO_4191 (O_4191,N_42201,N_44645);
nor UO_4192 (O_4192,N_49720,N_49007);
and UO_4193 (O_4193,N_43320,N_44194);
nand UO_4194 (O_4194,N_44776,N_47928);
or UO_4195 (O_4195,N_48223,N_49641);
nor UO_4196 (O_4196,N_46629,N_42672);
nor UO_4197 (O_4197,N_42937,N_45564);
xor UO_4198 (O_4198,N_43267,N_41479);
nor UO_4199 (O_4199,N_40632,N_46440);
or UO_4200 (O_4200,N_43981,N_43827);
or UO_4201 (O_4201,N_41067,N_47742);
and UO_4202 (O_4202,N_48135,N_48653);
xnor UO_4203 (O_4203,N_40033,N_40567);
or UO_4204 (O_4204,N_48984,N_41105);
nand UO_4205 (O_4205,N_43181,N_44018);
and UO_4206 (O_4206,N_46509,N_41087);
or UO_4207 (O_4207,N_42037,N_47698);
and UO_4208 (O_4208,N_47281,N_49002);
nand UO_4209 (O_4209,N_47267,N_46604);
xnor UO_4210 (O_4210,N_46923,N_48357);
nor UO_4211 (O_4211,N_46508,N_46556);
and UO_4212 (O_4212,N_44473,N_47044);
or UO_4213 (O_4213,N_44825,N_42808);
nand UO_4214 (O_4214,N_44343,N_48758);
or UO_4215 (O_4215,N_41025,N_45713);
nor UO_4216 (O_4216,N_48817,N_45104);
nor UO_4217 (O_4217,N_48614,N_42634);
nand UO_4218 (O_4218,N_48527,N_40790);
nand UO_4219 (O_4219,N_49174,N_41708);
nor UO_4220 (O_4220,N_42249,N_45146);
nor UO_4221 (O_4221,N_44082,N_45127);
and UO_4222 (O_4222,N_42608,N_47224);
nand UO_4223 (O_4223,N_48849,N_40178);
nand UO_4224 (O_4224,N_45742,N_40197);
and UO_4225 (O_4225,N_45478,N_46042);
nand UO_4226 (O_4226,N_48092,N_42294);
or UO_4227 (O_4227,N_48089,N_42432);
or UO_4228 (O_4228,N_49364,N_47670);
and UO_4229 (O_4229,N_44724,N_49841);
or UO_4230 (O_4230,N_40797,N_42172);
nand UO_4231 (O_4231,N_49302,N_42806);
nand UO_4232 (O_4232,N_48420,N_40688);
nand UO_4233 (O_4233,N_48804,N_43557);
nor UO_4234 (O_4234,N_49059,N_40840);
nand UO_4235 (O_4235,N_45413,N_44985);
nand UO_4236 (O_4236,N_48150,N_46812);
or UO_4237 (O_4237,N_40806,N_44280);
and UO_4238 (O_4238,N_42894,N_41902);
nor UO_4239 (O_4239,N_47040,N_47014);
or UO_4240 (O_4240,N_41312,N_48176);
nor UO_4241 (O_4241,N_46005,N_48873);
and UO_4242 (O_4242,N_44180,N_47966);
and UO_4243 (O_4243,N_46699,N_44184);
nor UO_4244 (O_4244,N_43224,N_49936);
and UO_4245 (O_4245,N_49955,N_46081);
or UO_4246 (O_4246,N_41223,N_41583);
or UO_4247 (O_4247,N_41792,N_40693);
or UO_4248 (O_4248,N_40409,N_41811);
or UO_4249 (O_4249,N_44231,N_48146);
or UO_4250 (O_4250,N_42337,N_44342);
nor UO_4251 (O_4251,N_40232,N_49987);
or UO_4252 (O_4252,N_41941,N_43046);
and UO_4253 (O_4253,N_41869,N_42424);
nand UO_4254 (O_4254,N_43847,N_49203);
and UO_4255 (O_4255,N_42847,N_47369);
nor UO_4256 (O_4256,N_45778,N_46794);
xnor UO_4257 (O_4257,N_49230,N_41904);
nor UO_4258 (O_4258,N_41041,N_41749);
or UO_4259 (O_4259,N_44446,N_42225);
nor UO_4260 (O_4260,N_47988,N_47365);
xor UO_4261 (O_4261,N_42399,N_44295);
or UO_4262 (O_4262,N_45570,N_43431);
nand UO_4263 (O_4263,N_47258,N_49837);
and UO_4264 (O_4264,N_40942,N_42067);
and UO_4265 (O_4265,N_43925,N_43309);
and UO_4266 (O_4266,N_41906,N_48451);
nand UO_4267 (O_4267,N_44719,N_41960);
or UO_4268 (O_4268,N_46839,N_40174);
and UO_4269 (O_4269,N_43824,N_45025);
xnor UO_4270 (O_4270,N_41939,N_41817);
xnor UO_4271 (O_4271,N_43848,N_44308);
nor UO_4272 (O_4272,N_45130,N_49448);
nor UO_4273 (O_4273,N_45815,N_46895);
or UO_4274 (O_4274,N_48732,N_40357);
and UO_4275 (O_4275,N_40568,N_43821);
nand UO_4276 (O_4276,N_41472,N_44998);
or UO_4277 (O_4277,N_42022,N_47455);
or UO_4278 (O_4278,N_41970,N_42881);
nor UO_4279 (O_4279,N_41755,N_45469);
nor UO_4280 (O_4280,N_48343,N_49692);
or UO_4281 (O_4281,N_48615,N_42411);
nand UO_4282 (O_4282,N_42377,N_47123);
or UO_4283 (O_4283,N_41702,N_44859);
nand UO_4284 (O_4284,N_48315,N_47127);
or UO_4285 (O_4285,N_43282,N_46911);
xor UO_4286 (O_4286,N_48681,N_47459);
or UO_4287 (O_4287,N_46415,N_46050);
and UO_4288 (O_4288,N_46548,N_40043);
or UO_4289 (O_4289,N_47106,N_41244);
nand UO_4290 (O_4290,N_45031,N_48509);
nand UO_4291 (O_4291,N_44036,N_43095);
and UO_4292 (O_4292,N_43891,N_40523);
nand UO_4293 (O_4293,N_48216,N_45688);
and UO_4294 (O_4294,N_44266,N_47752);
or UO_4295 (O_4295,N_44947,N_41342);
and UO_4296 (O_4296,N_47984,N_40382);
and UO_4297 (O_4297,N_45247,N_40814);
or UO_4298 (O_4298,N_49818,N_49132);
or UO_4299 (O_4299,N_44956,N_41609);
and UO_4300 (O_4300,N_43600,N_40522);
or UO_4301 (O_4301,N_47011,N_44783);
and UO_4302 (O_4302,N_47518,N_47708);
nor UO_4303 (O_4303,N_42156,N_46644);
xnor UO_4304 (O_4304,N_42384,N_47414);
and UO_4305 (O_4305,N_46054,N_46214);
nand UO_4306 (O_4306,N_46704,N_49788);
or UO_4307 (O_4307,N_45798,N_41435);
nand UO_4308 (O_4308,N_40732,N_42275);
and UO_4309 (O_4309,N_40929,N_44112);
nor UO_4310 (O_4310,N_46879,N_40847);
nand UO_4311 (O_4311,N_45735,N_45372);
nor UO_4312 (O_4312,N_46309,N_46570);
nand UO_4313 (O_4313,N_41138,N_44183);
nor UO_4314 (O_4314,N_45957,N_48469);
and UO_4315 (O_4315,N_48600,N_47792);
nor UO_4316 (O_4316,N_49694,N_47805);
and UO_4317 (O_4317,N_41539,N_45056);
nor UO_4318 (O_4318,N_48164,N_47686);
or UO_4319 (O_4319,N_42743,N_42870);
nand UO_4320 (O_4320,N_44281,N_43498);
nand UO_4321 (O_4321,N_46883,N_42917);
and UO_4322 (O_4322,N_49098,N_44091);
nand UO_4323 (O_4323,N_40524,N_45660);
nand UO_4324 (O_4324,N_49264,N_45966);
nand UO_4325 (O_4325,N_41274,N_43059);
and UO_4326 (O_4326,N_42228,N_40397);
and UO_4327 (O_4327,N_46621,N_40246);
or UO_4328 (O_4328,N_46780,N_46821);
nand UO_4329 (O_4329,N_43319,N_44961);
or UO_4330 (O_4330,N_44837,N_48194);
nand UO_4331 (O_4331,N_41529,N_45195);
or UO_4332 (O_4332,N_45389,N_43202);
nor UO_4333 (O_4333,N_40263,N_49077);
xnor UO_4334 (O_4334,N_40310,N_49657);
nor UO_4335 (O_4335,N_43036,N_43616);
or UO_4336 (O_4336,N_46872,N_44742);
nor UO_4337 (O_4337,N_48186,N_46372);
nor UO_4338 (O_4338,N_49103,N_46527);
and UO_4339 (O_4339,N_45650,N_43873);
nand UO_4340 (O_4340,N_47222,N_48945);
or UO_4341 (O_4341,N_40384,N_40410);
and UO_4342 (O_4342,N_41341,N_40337);
nor UO_4343 (O_4343,N_44432,N_40653);
and UO_4344 (O_4344,N_49484,N_42778);
nor UO_4345 (O_4345,N_49874,N_42134);
and UO_4346 (O_4346,N_40227,N_46703);
nor UO_4347 (O_4347,N_42235,N_45243);
and UO_4348 (O_4348,N_46183,N_48130);
or UO_4349 (O_4349,N_41720,N_49123);
nor UO_4350 (O_4350,N_48837,N_43067);
nor UO_4351 (O_4351,N_48748,N_48620);
xor UO_4352 (O_4352,N_47160,N_44467);
nor UO_4353 (O_4353,N_48575,N_40873);
or UO_4354 (O_4354,N_43459,N_42609);
and UO_4355 (O_4355,N_48565,N_44618);
nand UO_4356 (O_4356,N_49119,N_41320);
nor UO_4357 (O_4357,N_47428,N_49309);
and UO_4358 (O_4358,N_45836,N_46089);
xor UO_4359 (O_4359,N_46590,N_42705);
and UO_4360 (O_4360,N_46871,N_40899);
nor UO_4361 (O_4361,N_41956,N_42048);
nand UO_4362 (O_4362,N_45974,N_42505);
and UO_4363 (O_4363,N_46578,N_42216);
or UO_4364 (O_4364,N_47249,N_40474);
nor UO_4365 (O_4365,N_41802,N_41329);
nor UO_4366 (O_4366,N_40047,N_45667);
nor UO_4367 (O_4367,N_42044,N_47138);
nor UO_4368 (O_4368,N_46443,N_46204);
and UO_4369 (O_4369,N_40446,N_46619);
nand UO_4370 (O_4370,N_43911,N_45286);
nor UO_4371 (O_4371,N_42279,N_47094);
nor UO_4372 (O_4372,N_40900,N_49177);
nand UO_4373 (O_4373,N_44272,N_47228);
or UO_4374 (O_4374,N_41433,N_46156);
nor UO_4375 (O_4375,N_40723,N_46017);
xnor UO_4376 (O_4376,N_49934,N_45556);
nor UO_4377 (O_4377,N_42073,N_45317);
nor UO_4378 (O_4378,N_49222,N_48647);
nor UO_4379 (O_4379,N_44322,N_44158);
nand UO_4380 (O_4380,N_40626,N_45586);
nand UO_4381 (O_4381,N_46084,N_42818);
nand UO_4382 (O_4382,N_48648,N_44404);
nor UO_4383 (O_4383,N_44630,N_47099);
nand UO_4384 (O_4384,N_42658,N_48444);
and UO_4385 (O_4385,N_49136,N_48003);
nor UO_4386 (O_4386,N_48437,N_43115);
nor UO_4387 (O_4387,N_47860,N_43678);
nand UO_4388 (O_4388,N_42345,N_46427);
and UO_4389 (O_4389,N_49783,N_48788);
nand UO_4390 (O_4390,N_45625,N_49990);
xnor UO_4391 (O_4391,N_42865,N_42202);
nor UO_4392 (O_4392,N_43449,N_48389);
or UO_4393 (O_4393,N_49006,N_48434);
nand UO_4394 (O_4394,N_40776,N_44925);
nand UO_4395 (O_4395,N_41883,N_42456);
nand UO_4396 (O_4396,N_48629,N_49276);
and UO_4397 (O_4397,N_49105,N_40645);
or UO_4398 (O_4398,N_44526,N_41907);
and UO_4399 (O_4399,N_42903,N_46693);
nand UO_4400 (O_4400,N_48519,N_43698);
and UO_4401 (O_4401,N_47162,N_49124);
nor UO_4402 (O_4402,N_48972,N_43634);
nor UO_4403 (O_4403,N_45581,N_49533);
nand UO_4404 (O_4404,N_45716,N_47717);
or UO_4405 (O_4405,N_43160,N_48001);
or UO_4406 (O_4406,N_47582,N_49731);
and UO_4407 (O_4407,N_44043,N_47444);
or UO_4408 (O_4408,N_42947,N_44765);
and UO_4409 (O_4409,N_45542,N_41169);
xor UO_4410 (O_4410,N_48678,N_41289);
and UO_4411 (O_4411,N_40922,N_49805);
and UO_4412 (O_4412,N_48516,N_43649);
nor UO_4413 (O_4413,N_45659,N_42710);
or UO_4414 (O_4414,N_43760,N_40018);
or UO_4415 (O_4415,N_44242,N_42644);
and UO_4416 (O_4416,N_46101,N_47709);
nor UO_4417 (O_4417,N_41158,N_43276);
nor UO_4418 (O_4418,N_49733,N_43524);
or UO_4419 (O_4419,N_43152,N_42662);
and UO_4420 (O_4420,N_48144,N_44355);
nor UO_4421 (O_4421,N_44373,N_48810);
and UO_4422 (O_4422,N_47535,N_40615);
and UO_4423 (O_4423,N_43640,N_42184);
or UO_4424 (O_4424,N_46733,N_44165);
nand UO_4425 (O_4425,N_40893,N_49989);
and UO_4426 (O_4426,N_46297,N_43930);
and UO_4427 (O_4427,N_42276,N_40340);
xor UO_4428 (O_4428,N_42654,N_47064);
or UO_4429 (O_4429,N_43085,N_47839);
or UO_4430 (O_4430,N_45740,N_40894);
xor UO_4431 (O_4431,N_49752,N_47031);
nor UO_4432 (O_4432,N_46093,N_49501);
nand UO_4433 (O_4433,N_45324,N_42091);
or UO_4434 (O_4434,N_47153,N_49352);
nand UO_4435 (O_4435,N_44328,N_48254);
and UO_4436 (O_4436,N_47834,N_42296);
or UO_4437 (O_4437,N_40908,N_44699);
xnor UO_4438 (O_4438,N_44793,N_40987);
or UO_4439 (O_4439,N_43755,N_49143);
nand UO_4440 (O_4440,N_44126,N_41637);
nor UO_4441 (O_4441,N_44748,N_42604);
or UO_4442 (O_4442,N_44522,N_40148);
nand UO_4443 (O_4443,N_46576,N_43934);
and UO_4444 (O_4444,N_41830,N_41840);
nor UO_4445 (O_4445,N_49296,N_48322);
nor UO_4446 (O_4446,N_41220,N_45419);
and UO_4447 (O_4447,N_40477,N_47851);
nand UO_4448 (O_4448,N_46473,N_45728);
nand UO_4449 (O_4449,N_44847,N_43960);
xor UO_4450 (O_4450,N_40867,N_45662);
nor UO_4451 (O_4451,N_48955,N_48082);
nor UO_4452 (O_4452,N_47333,N_43339);
nand UO_4453 (O_4453,N_44202,N_47056);
nor UO_4454 (O_4454,N_49280,N_44973);
nor UO_4455 (O_4455,N_45276,N_48476);
or UO_4456 (O_4456,N_44339,N_42126);
or UO_4457 (O_4457,N_43192,N_44407);
nor UO_4458 (O_4458,N_45322,N_45412);
or UO_4459 (O_4459,N_47069,N_45138);
nor UO_4460 (O_4460,N_42342,N_42545);
or UO_4461 (O_4461,N_49285,N_40036);
nand UO_4462 (O_4462,N_43372,N_43522);
nor UO_4463 (O_4463,N_40778,N_41057);
nor UO_4464 (O_4464,N_47035,N_48705);
or UO_4465 (O_4465,N_42925,N_41353);
nand UO_4466 (O_4466,N_44546,N_47430);
nand UO_4467 (O_4467,N_42759,N_42794);
nand UO_4468 (O_4468,N_47205,N_44497);
and UO_4469 (O_4469,N_48564,N_46713);
or UO_4470 (O_4470,N_44957,N_41077);
and UO_4471 (O_4471,N_46600,N_42098);
nor UO_4472 (O_4472,N_47080,N_46264);
nand UO_4473 (O_4473,N_41682,N_41938);
and UO_4474 (O_4474,N_44737,N_45612);
nor UO_4475 (O_4475,N_42955,N_41285);
xor UO_4476 (O_4476,N_46289,N_41060);
or UO_4477 (O_4477,N_46747,N_42318);
nand UO_4478 (O_4478,N_48178,N_41068);
xor UO_4479 (O_4479,N_44626,N_41248);
nand UO_4480 (O_4480,N_45677,N_44833);
nand UO_4481 (O_4481,N_43100,N_40101);
or UO_4482 (O_4482,N_40160,N_44778);
or UO_4483 (O_4483,N_49613,N_45226);
or UO_4484 (O_4484,N_49288,N_47366);
or UO_4485 (O_4485,N_47360,N_43051);
and UO_4486 (O_4486,N_40596,N_44481);
nand UO_4487 (O_4487,N_41359,N_42403);
nor UO_4488 (O_4488,N_41563,N_46939);
or UO_4489 (O_4489,N_49687,N_49558);
and UO_4490 (O_4490,N_43168,N_41544);
and UO_4491 (O_4491,N_41246,N_42977);
and UO_4492 (O_4492,N_43165,N_48948);
or UO_4493 (O_4493,N_47343,N_43578);
nor UO_4494 (O_4494,N_44940,N_46609);
nand UO_4495 (O_4495,N_48157,N_47096);
nor UO_4496 (O_4496,N_48005,N_49823);
and UO_4497 (O_4497,N_44346,N_41429);
and UO_4498 (O_4498,N_45428,N_44518);
or UO_4499 (O_4499,N_40581,N_40585);
and UO_4500 (O_4500,N_48386,N_47569);
and UO_4501 (O_4501,N_47970,N_41328);
nor UO_4502 (O_4502,N_40620,N_49510);
xor UO_4503 (O_4503,N_44301,N_44994);
and UO_4504 (O_4504,N_40428,N_49246);
nor UO_4505 (O_4505,N_43626,N_46248);
xor UO_4506 (O_4506,N_48380,N_49704);
nor UO_4507 (O_4507,N_44667,N_45049);
nand UO_4508 (O_4508,N_41642,N_46866);
nand UO_4509 (O_4509,N_40265,N_43586);
nand UO_4510 (O_4510,N_44760,N_40683);
and UO_4511 (O_4511,N_45194,N_46186);
nand UO_4512 (O_4512,N_43785,N_42607);
and UO_4513 (O_4513,N_44236,N_46787);
or UO_4514 (O_4514,N_40588,N_49844);
and UO_4515 (O_4515,N_42677,N_45594);
xor UO_4516 (O_4516,N_41142,N_43318);
or UO_4517 (O_4517,N_49670,N_43754);
nand UO_4518 (O_4518,N_46255,N_47379);
or UO_4519 (O_4519,N_47773,N_48301);
xnor UO_4520 (O_4520,N_48102,N_49626);
or UO_4521 (O_4521,N_47882,N_44478);
and UO_4522 (O_4522,N_48799,N_48262);
and UO_4523 (O_4523,N_40420,N_42617);
or UO_4524 (O_4524,N_49111,N_40164);
or UO_4525 (O_4525,N_43308,N_44873);
and UO_4526 (O_4526,N_46117,N_49638);
nor UO_4527 (O_4527,N_48712,N_41478);
nand UO_4528 (O_4528,N_49168,N_47061);
or UO_4529 (O_4529,N_46513,N_40117);
and UO_4530 (O_4530,N_45028,N_47965);
nor UO_4531 (O_4531,N_44302,N_40106);
or UO_4532 (O_4532,N_48932,N_47783);
nor UO_4533 (O_4533,N_40291,N_43690);
nand UO_4534 (O_4534,N_48922,N_41233);
nand UO_4535 (O_4535,N_41704,N_46841);
and UO_4536 (O_4536,N_46215,N_47596);
nor UO_4537 (O_4537,N_48751,N_48766);
xor UO_4538 (O_4538,N_48306,N_47479);
nor UO_4539 (O_4539,N_49540,N_40119);
and UO_4540 (O_4540,N_43020,N_40365);
nor UO_4541 (O_4541,N_48358,N_49551);
nor UO_4542 (O_4542,N_43084,N_49748);
nor UO_4543 (O_4543,N_41773,N_46308);
xor UO_4544 (O_4544,N_42429,N_47405);
nor UO_4545 (O_4545,N_42799,N_49319);
xnor UO_4546 (O_4546,N_43293,N_42474);
xnor UO_4547 (O_4547,N_49183,N_41319);
or UO_4548 (O_4548,N_45113,N_49796);
or UO_4549 (O_4549,N_40833,N_41710);
nand UO_4550 (O_4550,N_44745,N_40031);
nand UO_4551 (O_4551,N_45391,N_49224);
and UO_4552 (O_4552,N_41079,N_46663);
xor UO_4553 (O_4553,N_46521,N_48856);
nand UO_4554 (O_4554,N_44405,N_43956);
nor UO_4555 (O_4555,N_46288,N_45502);
nor UO_4556 (O_4556,N_42493,N_41480);
or UO_4557 (O_4557,N_45912,N_42109);
or UO_4558 (O_4558,N_48552,N_48752);
or UO_4559 (O_4559,N_49560,N_44113);
nor UO_4560 (O_4560,N_45819,N_46559);
and UO_4561 (O_4561,N_47516,N_47500);
nand UO_4562 (O_4562,N_44020,N_49417);
nor UO_4563 (O_4563,N_44545,N_41228);
and UO_4564 (O_4564,N_48820,N_40968);
nand UO_4565 (O_4565,N_40580,N_46294);
or UO_4566 (O_4566,N_44976,N_46336);
nor UO_4567 (O_4567,N_46063,N_49639);
nand UO_4568 (O_4568,N_42802,N_49984);
nor UO_4569 (O_4569,N_40537,N_40911);
or UO_4570 (O_4570,N_44235,N_45599);
nand UO_4571 (O_4571,N_48303,N_47238);
nand UO_4572 (O_4572,N_43231,N_45244);
or UO_4573 (O_4573,N_47810,N_41486);
and UO_4574 (O_4574,N_41783,N_40858);
xnor UO_4575 (O_4575,N_40950,N_47957);
nor UO_4576 (O_4576,N_48903,N_49944);
or UO_4577 (O_4577,N_41487,N_48369);
or UO_4578 (O_4578,N_40989,N_40659);
nor UO_4579 (O_4579,N_42068,N_41818);
xor UO_4580 (O_4580,N_44858,N_46376);
nor UO_4581 (O_4581,N_49113,N_47187);
xnor UO_4582 (O_4582,N_47277,N_40220);
nand UO_4583 (O_4583,N_40244,N_42299);
nand UO_4584 (O_4584,N_43993,N_44885);
nor UO_4585 (O_4585,N_48043,N_43904);
or UO_4586 (O_4586,N_44185,N_43574);
or UO_4587 (O_4587,N_42306,N_49304);
and UO_4588 (O_4588,N_46694,N_48155);
nor UO_4589 (O_4589,N_49153,N_47321);
or UO_4590 (O_4590,N_40741,N_46573);
nand UO_4591 (O_4591,N_40875,N_49299);
nand UO_4592 (O_4592,N_41864,N_41687);
xnor UO_4593 (O_4593,N_48201,N_46786);
nand UO_4594 (O_4594,N_40204,N_41419);
nor UO_4595 (O_4595,N_45838,N_49424);
nor UO_4596 (O_4596,N_49107,N_47908);
or UO_4597 (O_4597,N_48885,N_41306);
nor UO_4598 (O_4598,N_44362,N_41141);
and UO_4599 (O_4599,N_49050,N_46753);
nor UO_4600 (O_4600,N_43830,N_44939);
nor UO_4601 (O_4601,N_48869,N_47564);
or UO_4602 (O_4602,N_48554,N_47221);
xor UO_4603 (O_4603,N_42819,N_42419);
and UO_4604 (O_4604,N_43359,N_42232);
nand UO_4605 (O_4605,N_45952,N_48336);
and UO_4606 (O_4606,N_47458,N_43003);
nand UO_4607 (O_4607,N_41183,N_42970);
nand UO_4608 (O_4608,N_47779,N_42036);
nor UO_4609 (O_4609,N_44524,N_48725);
or UO_4610 (O_4610,N_44377,N_47684);
nand UO_4611 (O_4611,N_48342,N_47299);
nand UO_4612 (O_4612,N_43894,N_43186);
and UO_4613 (O_4613,N_49354,N_49227);
and UO_4614 (O_4614,N_44066,N_42983);
or UO_4615 (O_4615,N_44999,N_42699);
or UO_4616 (O_4616,N_45029,N_40571);
nor UO_4617 (O_4617,N_44484,N_49906);
or UO_4618 (O_4618,N_40259,N_42070);
nor UO_4619 (O_4619,N_46225,N_44829);
and UO_4620 (O_4620,N_47110,N_49567);
nand UO_4621 (O_4621,N_49397,N_46095);
nor UO_4622 (O_4622,N_43627,N_41393);
nor UO_4623 (O_4623,N_42973,N_40519);
or UO_4624 (O_4624,N_44327,N_46406);
and UO_4625 (O_4625,N_41253,N_49835);
and UO_4626 (O_4626,N_40566,N_41781);
and UO_4627 (O_4627,N_41001,N_40828);
nor UO_4628 (O_4628,N_48055,N_42175);
nand UO_4629 (O_4629,N_41473,N_46979);
or UO_4630 (O_4630,N_41511,N_41056);
nand UO_4631 (O_4631,N_42110,N_47410);
or UO_4632 (O_4632,N_44596,N_40288);
nor UO_4633 (O_4633,N_46847,N_43849);
or UO_4634 (O_4634,N_43630,N_41284);
or UO_4635 (O_4635,N_44533,N_45762);
nand UO_4636 (O_4636,N_47541,N_41377);
and UO_4637 (O_4637,N_44388,N_47359);
and UO_4638 (O_4638,N_46880,N_40985);
or UO_4639 (O_4639,N_43249,N_43071);
nand UO_4640 (O_4640,N_46507,N_42210);
nand UO_4641 (O_4641,N_49804,N_46481);
nor UO_4642 (O_4642,N_47246,N_48664);
and UO_4643 (O_4643,N_49423,N_42273);
nor UO_4644 (O_4644,N_41946,N_46003);
or UO_4645 (O_4645,N_40713,N_47295);
nor UO_4646 (O_4646,N_45796,N_47790);
nand UO_4647 (O_4647,N_47018,N_40928);
or UO_4648 (O_4648,N_41795,N_40017);
nand UO_4649 (O_4649,N_40369,N_41999);
xnor UO_4650 (O_4650,N_48506,N_47178);
and UO_4651 (O_4651,N_49179,N_47392);
nand UO_4652 (O_4652,N_49150,N_46767);
or UO_4653 (O_4653,N_42922,N_41717);
nor UO_4654 (O_4654,N_44055,N_46196);
nand UO_4655 (O_4655,N_41252,N_48297);
nand UO_4656 (O_4656,N_44498,N_43292);
nand UO_4657 (O_4657,N_43624,N_45781);
nand UO_4658 (O_4658,N_47163,N_49325);
and UO_4659 (O_4659,N_48097,N_47857);
xor UO_4660 (O_4660,N_44222,N_43154);
nor UO_4661 (O_4661,N_44787,N_46593);
and UO_4662 (O_4662,N_49415,N_42612);
xor UO_4663 (O_4663,N_42354,N_46449);
or UO_4664 (O_4664,N_42788,N_41180);
and UO_4665 (O_4665,N_48356,N_44739);
nor UO_4666 (O_4666,N_47933,N_45228);
nor UO_4667 (O_4667,N_45850,N_41388);
or UO_4668 (O_4668,N_41721,N_41872);
or UO_4669 (O_4669,N_43595,N_48220);
nor UO_4670 (O_4670,N_48823,N_45739);
and UO_4671 (O_4671,N_43709,N_44814);
or UO_4672 (O_4672,N_48755,N_46805);
nand UO_4673 (O_4673,N_40849,N_49572);
or UO_4674 (O_4674,N_42307,N_45332);
or UO_4675 (O_4675,N_43982,N_44738);
and UO_4676 (O_4676,N_46454,N_44811);
nand UO_4677 (O_4677,N_45652,N_46598);
or UO_4678 (O_4678,N_49005,N_40999);
and UO_4679 (O_4679,N_43969,N_42055);
xnor UO_4680 (O_4680,N_42413,N_48553);
nand UO_4681 (O_4681,N_40668,N_49036);
nor UO_4682 (O_4682,N_46360,N_45991);
or UO_4683 (O_4683,N_49358,N_45035);
nor UO_4684 (O_4684,N_43874,N_41422);
or UO_4685 (O_4685,N_46354,N_49734);
xnor UO_4686 (O_4686,N_46445,N_40095);
and UO_4687 (O_4687,N_46014,N_41611);
nand UO_4688 (O_4688,N_49517,N_47361);
nand UO_4689 (O_4689,N_45434,N_46470);
nor UO_4690 (O_4690,N_40954,N_46876);
nor UO_4691 (O_4691,N_40241,N_42630);
nor UO_4692 (O_4692,N_49311,N_47241);
and UO_4693 (O_4693,N_41777,N_49104);
xnor UO_4694 (O_4694,N_49434,N_48397);
or UO_4695 (O_4695,N_45327,N_47334);
or UO_4696 (O_4696,N_45864,N_46673);
xor UO_4697 (O_4697,N_43735,N_46616);
or UO_4698 (O_4698,N_48193,N_44818);
nand UO_4699 (O_4699,N_49624,N_47314);
or UO_4700 (O_4700,N_41888,N_46377);
and UO_4701 (O_4701,N_44255,N_42871);
nand UO_4702 (O_4702,N_41766,N_43804);
nand UO_4703 (O_4703,N_44789,N_46894);
nor UO_4704 (O_4704,N_43648,N_40682);
and UO_4705 (O_4705,N_47718,N_45653);
nand UO_4706 (O_4706,N_42602,N_46314);
nor UO_4707 (O_4707,N_40800,N_48659);
nor UO_4708 (O_4708,N_47542,N_42194);
nor UO_4709 (O_4709,N_42033,N_47112);
nor UO_4710 (O_4710,N_49742,N_47593);
or UO_4711 (O_4711,N_49410,N_46023);
or UO_4712 (O_4712,N_47059,N_47176);
or UO_4713 (O_4713,N_48661,N_45551);
nor UO_4714 (O_4714,N_48390,N_41011);
nand UO_4715 (O_4715,N_45414,N_45218);
and UO_4716 (O_4716,N_42757,N_40575);
and UO_4717 (O_4717,N_43143,N_44001);
or UO_4718 (O_4718,N_40464,N_46442);
or UO_4719 (O_4719,N_46159,N_49127);
nand UO_4720 (O_4720,N_49767,N_45041);
nand UO_4721 (O_4721,N_40556,N_45116);
and UO_4722 (O_4722,N_49973,N_40255);
or UO_4723 (O_4723,N_42335,N_40501);
xor UO_4724 (O_4724,N_49591,N_49402);
nand UO_4725 (O_4725,N_44988,N_42315);
or UO_4726 (O_4726,N_49598,N_45471);
nand UO_4727 (O_4727,N_49171,N_43423);
nor UO_4728 (O_4728,N_49416,N_45371);
and UO_4729 (O_4729,N_40933,N_49377);
nand UO_4730 (O_4730,N_41876,N_46706);
nor UO_4731 (O_4731,N_43895,N_49892);
and UO_4732 (O_4732,N_41861,N_48347);
nor UO_4733 (O_4733,N_46039,N_48410);
xor UO_4734 (O_4734,N_45930,N_43333);
nand UO_4735 (O_4735,N_43940,N_40624);
and UO_4736 (O_4736,N_40838,N_42253);
and UO_4737 (O_4737,N_41787,N_42583);
xor UO_4738 (O_4738,N_44538,N_48715);
xnor UO_4739 (O_4739,N_47395,N_48852);
nor UO_4740 (O_4740,N_45292,N_42574);
nand UO_4741 (O_4741,N_47781,N_47885);
and UO_4742 (O_4742,N_49897,N_43514);
and UO_4743 (O_4743,N_46334,N_42149);
and UO_4744 (O_4744,N_49278,N_43027);
nor UO_4745 (O_4745,N_43287,N_48139);
nor UO_4746 (O_4746,N_47184,N_44372);
or UO_4747 (O_4747,N_49649,N_43509);
and UO_4748 (O_4748,N_41981,N_46446);
nand UO_4749 (O_4749,N_40274,N_48534);
or UO_4750 (O_4750,N_41481,N_42580);
and UO_4751 (O_4751,N_41593,N_48582);
nand UO_4752 (O_4752,N_47867,N_46656);
nand UO_4753 (O_4753,N_41408,N_44376);
and UO_4754 (O_4754,N_42431,N_43779);
nand UO_4755 (O_4755,N_44337,N_48761);
nand UO_4756 (O_4756,N_48127,N_45786);
nand UO_4757 (O_4757,N_49791,N_47524);
nor UO_4758 (O_4758,N_46558,N_45601);
nand UO_4759 (O_4759,N_49065,N_41986);
nor UO_4760 (O_4760,N_44734,N_43488);
nand UO_4761 (O_4761,N_44511,N_44298);
xnor UO_4762 (O_4762,N_44563,N_42400);
nor UO_4763 (O_4763,N_49166,N_44569);
xor UO_4764 (O_4764,N_47729,N_42005);
nand UO_4765 (O_4765,N_42629,N_42990);
nand UO_4766 (O_4766,N_47666,N_40044);
and UO_4767 (O_4767,N_49819,N_45541);
nand UO_4768 (O_4768,N_41265,N_48668);
nand UO_4769 (O_4769,N_42321,N_44899);
nor UO_4770 (O_4770,N_49951,N_48079);
nor UO_4771 (O_4771,N_41798,N_45254);
or UO_4772 (O_4772,N_44326,N_40460);
or UO_4773 (O_4773,N_49012,N_40203);
or UO_4774 (O_4774,N_43645,N_43451);
nor UO_4775 (O_4775,N_45571,N_49060);
nor UO_4776 (O_4776,N_47696,N_41694);
or UO_4777 (O_4777,N_43924,N_49632);
or UO_4778 (O_4778,N_47013,N_49949);
nor UO_4779 (O_4779,N_45964,N_40605);
nand UO_4780 (O_4780,N_42314,N_45689);
or UO_4781 (O_4781,N_46997,N_49211);
and UO_4782 (O_4782,N_40294,N_41531);
nand UO_4783 (O_4783,N_46529,N_43660);
nor UO_4784 (O_4784,N_43883,N_49305);
xnor UO_4785 (O_4785,N_48203,N_45114);
or UO_4786 (O_4786,N_48385,N_40059);
and UO_4787 (O_4787,N_48785,N_43773);
nor UO_4788 (O_4788,N_40318,N_47530);
or UO_4789 (O_4789,N_45956,N_47169);
nor UO_4790 (O_4790,N_42993,N_45921);
nand UO_4791 (O_4791,N_47434,N_44468);
nor UO_4792 (O_4792,N_49213,N_43792);
or UO_4793 (O_4793,N_48578,N_44503);
nand UO_4794 (O_4794,N_42938,N_41762);
and UO_4795 (O_4795,N_49972,N_43198);
nand UO_4796 (O_4796,N_44633,N_41775);
nor UO_4797 (O_4797,N_40495,N_47927);
or UO_4798 (O_4798,N_48056,N_41172);
or UO_4799 (O_4799,N_42726,N_49924);
nor UO_4800 (O_4800,N_42009,N_47204);
and UO_4801 (O_4801,N_40328,N_48605);
and UO_4802 (O_4802,N_48612,N_41468);
nand UO_4803 (O_4803,N_41871,N_49599);
nand UO_4804 (O_4804,N_48465,N_44930);
nor UO_4805 (O_4805,N_47656,N_40960);
nand UO_4806 (O_4806,N_43721,N_47899);
nand UO_4807 (O_4807,N_42800,N_40444);
nor UO_4808 (O_4808,N_42441,N_46959);
nand UO_4809 (O_4809,N_42624,N_45549);
nand UO_4810 (O_4810,N_47159,N_46395);
xor UO_4811 (O_4811,N_48897,N_43134);
nand UO_4812 (O_4812,N_45437,N_48074);
nor UO_4813 (O_4813,N_48285,N_47219);
nor UO_4814 (O_4814,N_46968,N_42375);
nor UO_4815 (O_4815,N_44462,N_45598);
xnor UO_4816 (O_4816,N_40448,N_44886);
nand UO_4817 (O_4817,N_49165,N_40173);
nor UO_4818 (O_4818,N_45411,N_41514);
nand UO_4819 (O_4819,N_48435,N_43949);
and UO_4820 (O_4820,N_42982,N_49180);
xor UO_4821 (O_4821,N_43138,N_43748);
nand UO_4822 (O_4822,N_40261,N_41806);
nor UO_4823 (O_4823,N_43822,N_48625);
or UO_4824 (O_4824,N_45298,N_45648);
nor UO_4825 (O_4825,N_46022,N_40159);
or UO_4826 (O_4826,N_49794,N_43907);
nor UO_4827 (O_4827,N_46889,N_49918);
or UO_4828 (O_4828,N_44487,N_40839);
or UO_4829 (O_4829,N_40206,N_45822);
and UO_4830 (O_4830,N_48086,N_45010);
nand UO_4831 (O_4831,N_49814,N_45026);
or UO_4832 (O_4832,N_41121,N_47348);
and UO_4833 (O_4833,N_46728,N_46066);
xor UO_4834 (O_4834,N_49683,N_44209);
xor UO_4835 (O_4835,N_41184,N_44386);
or UO_4836 (O_4836,N_47078,N_41730);
xnor UO_4837 (O_4837,N_40735,N_45800);
nand UO_4838 (O_4838,N_46589,N_46652);
nand UO_4839 (O_4839,N_47337,N_42836);
nor UO_4840 (O_4840,N_48392,N_47243);
and UO_4841 (O_4841,N_47158,N_45233);
and UO_4842 (O_4842,N_47144,N_43572);
xor UO_4843 (O_4843,N_42191,N_47215);
or UO_4844 (O_4844,N_42714,N_44096);
nor UO_4845 (O_4845,N_42874,N_45842);
or UO_4846 (O_4846,N_47139,N_47565);
and UO_4847 (O_4847,N_40440,N_45999);
and UO_4848 (O_4848,N_47347,N_48846);
nand UO_4849 (O_4849,N_41850,N_44840);
xnor UO_4850 (O_4850,N_45743,N_46463);
or UO_4851 (O_4851,N_46178,N_45600);
or UO_4852 (O_4852,N_43641,N_47830);
xor UO_4853 (O_4853,N_46400,N_40499);
nand UO_4854 (O_4854,N_47845,N_44856);
nor UO_4855 (O_4855,N_44398,N_49851);
nor UO_4856 (O_4856,N_41684,N_43516);
and UO_4857 (O_4857,N_45066,N_46640);
nor UO_4858 (O_4858,N_42238,N_42282);
or UO_4859 (O_4859,N_48495,N_49173);
nor UO_4860 (O_4860,N_48728,N_46834);
or UO_4861 (O_4861,N_42357,N_49684);
xor UO_4862 (O_4862,N_48934,N_41330);
nand UO_4863 (O_4863,N_43017,N_49201);
or UO_4864 (O_4864,N_49395,N_43474);
and UO_4865 (O_4865,N_41371,N_40625);
nor UO_4866 (O_4866,N_42492,N_48101);
nand UO_4867 (O_4867,N_44009,N_44621);
xnor UO_4868 (O_4868,N_45364,N_42298);
nor UO_4869 (O_4869,N_47872,N_48944);
and UO_4870 (O_4870,N_44286,N_40711);
nor UO_4871 (O_4871,N_49478,N_49080);
or UO_4872 (O_4872,N_43209,N_47431);
and UO_4873 (O_4873,N_40418,N_41187);
nor UO_4874 (O_4874,N_42704,N_42223);
or UO_4875 (O_4875,N_44196,N_46147);
or UO_4876 (O_4876,N_46359,N_44381);
nor UO_4877 (O_4877,N_45946,N_42020);
and UO_4878 (O_4878,N_48650,N_42614);
and UO_4879 (O_4879,N_44803,N_47371);
xnor UO_4880 (O_4880,N_42601,N_47954);
xnor UO_4881 (O_4881,N_41000,N_41560);
and UO_4882 (O_4882,N_49184,N_45349);
and UO_4883 (O_4883,N_48887,N_40582);
nor UO_4884 (O_4884,N_42497,N_48360);
or UO_4885 (O_4885,N_48583,N_49493);
nor UO_4886 (O_4886,N_49842,N_42975);
nand UO_4887 (O_4887,N_46691,N_47758);
nand UO_4888 (O_4888,N_43448,N_47207);
nand UO_4889 (O_4889,N_46342,N_44770);
nand UO_4890 (O_4890,N_43679,N_43235);
or UO_4891 (O_4891,N_43697,N_45139);
xnor UO_4892 (O_4892,N_41912,N_48456);
or UO_4893 (O_4893,N_49017,N_43629);
xnor UO_4894 (O_4894,N_47520,N_43096);
nand UO_4895 (O_4895,N_42158,N_40098);
nor UO_4896 (O_4896,N_45283,N_47012);
nor UO_4897 (O_4897,N_47678,N_47913);
and UO_4898 (O_4898,N_41303,N_49925);
nand UO_4899 (O_4899,N_45333,N_49062);
nand UO_4900 (O_4900,N_45210,N_42455);
xor UO_4901 (O_4901,N_41823,N_45693);
or UO_4902 (O_4902,N_49953,N_46718);
xnor UO_4903 (O_4903,N_41114,N_46337);
or UO_4904 (O_4904,N_48587,N_46285);
nand UO_4905 (O_4905,N_43352,N_47633);
nand UO_4906 (O_4906,N_47983,N_43299);
nand UO_4907 (O_4907,N_45663,N_46238);
or UO_4908 (O_4908,N_47237,N_47531);
and UO_4909 (O_4909,N_49401,N_49432);
xnor UO_4910 (O_4910,N_46332,N_48599);
nor UO_4911 (O_4911,N_49685,N_45268);
nor UO_4912 (O_4912,N_48407,N_45186);
and UO_4913 (O_4913,N_45180,N_40064);
nor UO_4914 (O_4914,N_41355,N_46477);
and UO_4915 (O_4915,N_44525,N_49043);
nand UO_4916 (O_4916,N_44561,N_40425);
xor UO_4917 (O_4917,N_49038,N_43166);
xor UO_4918 (O_4918,N_41497,N_48966);
or UO_4919 (O_4919,N_40392,N_44456);
or UO_4920 (O_4920,N_47071,N_43728);
nor UO_4921 (O_4921,N_41526,N_40202);
nand UO_4922 (O_4922,N_48860,N_40570);
xor UO_4923 (O_4923,N_47618,N_41586);
or UO_4924 (O_4924,N_40058,N_41524);
and UO_4925 (O_4925,N_42638,N_44564);
nand UO_4926 (O_4926,N_47286,N_44047);
or UO_4927 (O_4927,N_45048,N_40415);
or UO_4928 (O_4928,N_46540,N_40115);
xnor UO_4929 (O_4929,N_44085,N_48105);
nand UO_4930 (O_4930,N_45334,N_40482);
nor UO_4931 (O_4931,N_49073,N_43147);
nor UO_4932 (O_4932,N_46768,N_45940);
nand UO_4933 (O_4933,N_42562,N_47166);
nand UO_4934 (O_4934,N_47462,N_49335);
and UO_4935 (O_4935,N_40439,N_44084);
nor UO_4936 (O_4936,N_48192,N_47409);
and UO_4937 (O_4937,N_47574,N_48868);
nand UO_4938 (O_4938,N_48574,N_43236);
nand UO_4939 (O_4939,N_41853,N_41281);
or UO_4940 (O_4940,N_49965,N_46683);
xor UO_4941 (O_4941,N_40189,N_40108);
nor UO_4942 (O_4942,N_42823,N_42075);
or UO_4943 (O_4943,N_45213,N_45548);
nand UO_4944 (O_4944,N_48622,N_47665);
nand UO_4945 (O_4945,N_46584,N_47940);
and UO_4946 (O_4946,N_44732,N_41198);
nand UO_4947 (O_4947,N_45295,N_47283);
and UO_4948 (O_4948,N_48544,N_42855);
nand UO_4949 (O_4949,N_41186,N_45920);
and UO_4950 (O_4950,N_44795,N_48028);
or UO_4951 (O_4951,N_45156,N_45613);
nand UO_4952 (O_4952,N_46803,N_49218);
nand UO_4953 (O_4953,N_48805,N_47844);
or UO_4954 (O_4954,N_43985,N_43836);
or UO_4955 (O_4955,N_43345,N_41838);
nand UO_4956 (O_4956,N_47728,N_46686);
nor UO_4957 (O_4957,N_47391,N_45118);
xor UO_4958 (O_4958,N_46836,N_40016);
xnor UO_4959 (O_4959,N_49215,N_45868);
or UO_4960 (O_4960,N_42760,N_45694);
and UO_4961 (O_4961,N_48896,N_43279);
nor UO_4962 (O_4962,N_40391,N_48361);
and UO_4963 (O_4963,N_40829,N_45043);
and UO_4964 (O_4964,N_40358,N_40040);
or UO_4965 (O_4965,N_49750,N_45763);
nand UO_4966 (O_4966,N_44693,N_42391);
nor UO_4967 (O_4967,N_44965,N_41484);
and UO_4968 (O_4968,N_47766,N_48398);
nand UO_4969 (O_4969,N_44552,N_44303);
and UO_4970 (O_4970,N_46384,N_42218);
nor UO_4971 (O_4971,N_43531,N_45897);
or UO_4972 (O_4972,N_44791,N_44146);
or UO_4973 (O_4973,N_42632,N_43131);
or UO_4974 (O_4974,N_46296,N_41742);
and UO_4975 (O_4975,N_41451,N_41165);
nand UO_4976 (O_4976,N_47786,N_40042);
xor UO_4977 (O_4977,N_43566,N_42834);
nand UO_4978 (O_4978,N_42355,N_47920);
or UO_4979 (O_4979,N_49810,N_40236);
or UO_4980 (O_4980,N_44785,N_46245);
xor UO_4981 (O_4981,N_40578,N_49200);
xor UO_4982 (O_4982,N_48238,N_44038);
and UO_4983 (O_4983,N_45294,N_44979);
nor UO_4984 (O_4984,N_48453,N_40505);
or UO_4985 (O_4985,N_41089,N_45900);
and UO_4986 (O_4986,N_45787,N_47917);
nor UO_4987 (O_4987,N_45664,N_47417);
and UO_4988 (O_4988,N_43900,N_46236);
and UO_4989 (O_4989,N_43746,N_41618);
or UO_4990 (O_4990,N_47649,N_44510);
and UO_4991 (O_4991,N_42578,N_47468);
nand UO_4992 (O_4992,N_48651,N_42936);
nor UO_4993 (O_4993,N_47232,N_46350);
or UO_4994 (O_4994,N_47598,N_43986);
and UO_4995 (O_4995,N_40812,N_47734);
and UO_4996 (O_4996,N_47515,N_45896);
nor UO_4997 (O_4997,N_42350,N_42154);
nor UO_4998 (O_4998,N_45670,N_47145);
nor UO_4999 (O_4999,N_49813,N_44427);
endmodule