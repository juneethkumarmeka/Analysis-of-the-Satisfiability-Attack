module basic_2000_20000_2500_20_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_690,In_1592);
xor U1 (N_1,In_1980,In_1133);
nor U2 (N_2,In_1295,In_524);
or U3 (N_3,In_1613,In_1899);
xor U4 (N_4,In_499,In_644);
xor U5 (N_5,In_312,In_1563);
and U6 (N_6,In_1139,In_1169);
and U7 (N_7,In_1817,In_1081);
xnor U8 (N_8,In_1180,In_1161);
or U9 (N_9,In_1176,In_1950);
xor U10 (N_10,In_981,In_859);
or U11 (N_11,In_62,In_1994);
nor U12 (N_12,In_1825,In_982);
nor U13 (N_13,In_422,In_1603);
xor U14 (N_14,In_270,In_344);
or U15 (N_15,In_161,In_653);
and U16 (N_16,In_667,In_1101);
nand U17 (N_17,In_1668,In_1845);
or U18 (N_18,In_1400,In_49);
nand U19 (N_19,In_57,In_1061);
xor U20 (N_20,In_553,In_1401);
nand U21 (N_21,In_319,In_254);
or U22 (N_22,In_894,In_1475);
nand U23 (N_23,In_1941,In_624);
and U24 (N_24,In_103,In_4);
xnor U25 (N_25,In_188,In_1364);
xnor U26 (N_26,In_1215,In_990);
or U27 (N_27,In_154,In_750);
xnor U28 (N_28,In_1968,In_120);
nor U29 (N_29,In_515,In_1699);
nand U30 (N_30,In_144,In_955);
nor U31 (N_31,In_1499,In_500);
or U32 (N_32,In_480,In_1884);
xor U33 (N_33,In_852,In_522);
and U34 (N_34,In_386,In_761);
xnor U35 (N_35,In_431,In_1284);
nand U36 (N_36,In_964,In_1883);
or U37 (N_37,In_822,In_862);
nor U38 (N_38,In_1121,In_96);
nor U39 (N_39,In_591,In_1643);
or U40 (N_40,In_1595,In_655);
and U41 (N_41,In_742,In_730);
nor U42 (N_42,In_148,In_1085);
or U43 (N_43,In_1765,In_658);
and U44 (N_44,In_1137,In_132);
and U45 (N_45,In_130,In_1008);
and U46 (N_46,In_393,In_1182);
nor U47 (N_47,In_752,In_1484);
nand U48 (N_48,In_1443,In_537);
nor U49 (N_49,In_569,In_1472);
and U50 (N_50,In_809,In_347);
nand U51 (N_51,In_107,In_1524);
and U52 (N_52,In_1311,In_861);
or U53 (N_53,In_1453,In_71);
nor U54 (N_54,In_1653,In_1394);
xnor U55 (N_55,In_532,In_1103);
and U56 (N_56,In_1261,In_1220);
nand U57 (N_57,In_1018,In_1332);
nand U58 (N_58,In_455,In_1546);
nand U59 (N_59,In_1576,In_1266);
and U60 (N_60,In_1894,In_58);
and U61 (N_61,In_1494,In_1992);
or U62 (N_62,In_484,In_266);
or U63 (N_63,In_244,In_211);
nand U64 (N_64,In_1775,In_1226);
xnor U65 (N_65,In_1709,In_1673);
and U66 (N_66,In_164,In_1767);
xnor U67 (N_67,In_612,In_453);
and U68 (N_68,In_382,In_926);
and U69 (N_69,In_885,In_1834);
or U70 (N_70,In_1896,In_1536);
or U71 (N_71,In_596,In_378);
nor U72 (N_72,In_660,In_1143);
xnor U73 (N_73,In_390,In_592);
xnor U74 (N_74,In_1307,In_814);
xor U75 (N_75,In_479,In_415);
and U76 (N_76,In_1642,In_664);
xnor U77 (N_77,In_235,In_157);
nand U78 (N_78,In_406,In_588);
or U79 (N_79,In_1624,In_1551);
or U80 (N_80,In_1124,In_1744);
xnor U81 (N_81,In_1793,In_67);
nor U82 (N_82,In_1958,In_1373);
xor U83 (N_83,In_1265,In_452);
and U84 (N_84,In_1031,In_1891);
or U85 (N_85,In_1144,In_68);
and U86 (N_86,In_1518,In_940);
or U87 (N_87,In_679,In_192);
and U88 (N_88,In_368,In_463);
xnor U89 (N_89,In_520,In_1108);
xor U90 (N_90,In_392,In_478);
or U91 (N_91,In_1727,In_1131);
nand U92 (N_92,In_1325,In_1488);
nor U93 (N_93,In_1390,In_284);
nand U94 (N_94,In_40,In_399);
nor U95 (N_95,In_430,In_123);
nor U96 (N_96,In_1395,In_376);
and U97 (N_97,In_1384,In_714);
xnor U98 (N_98,In_195,In_1357);
xnor U99 (N_99,In_1809,In_137);
xnor U100 (N_100,In_208,In_202);
and U101 (N_101,In_1051,In_1663);
and U102 (N_102,In_259,In_1969);
xor U103 (N_103,In_1520,In_1508);
and U104 (N_104,In_1013,In_1150);
and U105 (N_105,In_1612,In_807);
and U106 (N_106,In_1882,In_1286);
nor U107 (N_107,In_1289,In_307);
nor U108 (N_108,In_700,In_1356);
nand U109 (N_109,In_1088,In_1294);
xnor U110 (N_110,In_1147,In_22);
nor U111 (N_111,In_1922,In_1846);
nor U112 (N_112,In_1399,In_385);
nor U113 (N_113,In_207,In_12);
nand U114 (N_114,In_554,In_863);
and U115 (N_115,In_1376,In_950);
and U116 (N_116,In_1723,In_1900);
nor U117 (N_117,In_369,In_1111);
xor U118 (N_118,In_48,In_1116);
nor U119 (N_119,In_912,In_389);
nand U120 (N_120,In_379,In_1585);
or U121 (N_121,In_1389,In_1632);
or U122 (N_122,In_1194,In_39);
or U123 (N_123,In_705,In_1577);
or U124 (N_124,In_840,In_535);
nand U125 (N_125,In_362,In_1388);
nor U126 (N_126,In_1532,In_1438);
or U127 (N_127,In_1635,In_634);
nand U128 (N_128,In_1828,In_829);
xor U129 (N_129,In_165,In_986);
nor U130 (N_130,In_1513,In_720);
nor U131 (N_131,In_1756,In_1029);
and U132 (N_132,In_676,In_1944);
nand U133 (N_133,In_1718,In_1140);
xnor U134 (N_134,In_474,In_909);
or U135 (N_135,In_127,In_1857);
xnor U136 (N_136,In_1670,In_567);
or U137 (N_137,In_963,In_666);
nor U138 (N_138,In_1501,In_1048);
and U139 (N_139,In_1757,In_907);
and U140 (N_140,In_1849,In_134);
and U141 (N_141,In_1319,In_823);
nor U142 (N_142,In_197,In_849);
nand U143 (N_143,In_1171,In_1231);
nand U144 (N_144,In_1737,In_1354);
nor U145 (N_145,In_1596,In_199);
xnor U146 (N_146,In_543,In_1213);
or U147 (N_147,In_928,In_1210);
or U148 (N_148,In_301,In_383);
xnor U149 (N_149,In_736,In_693);
and U150 (N_150,In_1032,In_1919);
and U151 (N_151,In_1745,In_23);
xnor U152 (N_152,In_349,In_366);
nand U153 (N_153,In_1788,In_1517);
nand U154 (N_154,In_317,In_182);
and U155 (N_155,In_518,In_30);
nor U156 (N_156,In_293,In_267);
nor U157 (N_157,In_684,In_771);
xor U158 (N_158,In_291,In_1437);
nor U159 (N_159,In_1128,In_1540);
and U160 (N_160,In_490,In_1254);
xnor U161 (N_161,In_1089,In_297);
nor U162 (N_162,In_348,In_1504);
and U163 (N_163,In_827,In_359);
or U164 (N_164,In_1905,In_1803);
or U165 (N_165,In_1,In_832);
nor U166 (N_166,In_943,In_1114);
nand U167 (N_167,In_1710,In_264);
or U168 (N_168,In_1850,In_1134);
nor U169 (N_169,In_1346,In_63);
xnor U170 (N_170,In_606,In_810);
nor U171 (N_171,In_1310,In_582);
and U172 (N_172,In_458,In_128);
or U173 (N_173,In_296,In_1255);
or U174 (N_174,In_64,In_657);
or U175 (N_175,In_28,In_1448);
nand U176 (N_176,In_1503,In_557);
nand U177 (N_177,In_1872,In_1976);
nand U178 (N_178,In_1010,In_129);
or U179 (N_179,In_1561,In_670);
nand U180 (N_180,In_513,In_1716);
or U181 (N_181,In_895,In_1371);
nor U182 (N_182,In_650,In_1921);
nand U183 (N_183,In_962,In_131);
nand U184 (N_184,In_1059,In_1330);
nand U185 (N_185,In_1746,In_139);
and U186 (N_186,In_918,In_1587);
nor U187 (N_187,In_1962,In_1074);
and U188 (N_188,In_1351,In_1338);
xor U189 (N_189,In_1270,In_751);
or U190 (N_190,In_1822,In_914);
nor U191 (N_191,In_294,In_1100);
xnor U192 (N_192,In_1211,In_1043);
nand U193 (N_193,In_1440,In_1873);
or U194 (N_194,In_1446,In_61);
nor U195 (N_195,In_1467,In_1071);
or U196 (N_196,In_642,In_1852);
nand U197 (N_197,In_1300,In_159);
nand U198 (N_198,In_475,In_1120);
or U199 (N_199,In_538,In_1249);
or U200 (N_200,In_184,In_1041);
and U201 (N_201,In_1073,In_1275);
xor U202 (N_202,In_571,In_1918);
nand U203 (N_203,In_258,In_231);
nor U204 (N_204,In_930,In_1479);
and U205 (N_205,In_602,In_101);
or U206 (N_206,In_864,In_1303);
xor U207 (N_207,In_168,In_1908);
nor U208 (N_208,In_476,In_597);
nand U209 (N_209,In_1471,In_1527);
or U210 (N_210,In_420,In_1207);
and U211 (N_211,In_257,In_276);
nor U212 (N_212,In_710,In_1413);
or U213 (N_213,In_1327,In_35);
xnor U214 (N_214,In_425,In_1362);
nand U215 (N_215,In_1023,In_821);
or U216 (N_216,In_1953,In_1618);
xor U217 (N_217,In_502,In_1189);
nand U218 (N_218,In_1195,In_1700);
nand U219 (N_219,In_1515,In_1667);
nor U220 (N_220,In_1753,In_1854);
nor U221 (N_221,In_1014,In_1072);
nor U222 (N_222,In_1291,In_1886);
nand U223 (N_223,In_577,In_1251);
and U224 (N_224,In_1246,In_726);
nand U225 (N_225,In_1223,In_1069);
and U226 (N_226,In_1611,In_247);
xor U227 (N_227,In_958,In_1414);
and U228 (N_228,In_1687,In_245);
nor U229 (N_229,In_1320,In_1661);
and U230 (N_230,In_782,In_1412);
nor U231 (N_231,In_566,In_551);
xor U232 (N_232,In_1110,In_135);
nor U233 (N_233,In_1135,In_1447);
nand U234 (N_234,In_473,In_1481);
and U235 (N_235,In_629,In_1786);
nor U236 (N_236,In_1118,In_1880);
nor U237 (N_237,In_1863,In_1277);
or U238 (N_238,In_1993,In_367);
and U239 (N_239,In_1916,In_1094);
nor U240 (N_240,In_394,In_739);
nand U241 (N_241,In_808,In_433);
or U242 (N_242,In_1923,In_1168);
or U243 (N_243,In_768,In_590);
or U244 (N_244,In_371,In_239);
nand U245 (N_245,In_281,In_898);
nor U246 (N_246,In_1904,In_1201);
xor U247 (N_247,In_806,In_681);
nand U248 (N_248,In_892,In_1827);
nor U249 (N_249,In_1491,In_1256);
nor U250 (N_250,In_1847,In_1198);
xor U251 (N_251,In_1998,In_753);
or U252 (N_252,In_1728,In_1044);
nand U253 (N_253,In_398,In_1910);
nand U254 (N_254,In_1681,In_1777);
nand U255 (N_255,In_260,In_1196);
and U256 (N_256,In_114,In_97);
nand U257 (N_257,In_610,In_1529);
xnor U258 (N_258,In_1463,In_1773);
or U259 (N_259,In_793,In_384);
nor U260 (N_260,In_977,In_1404);
and U261 (N_261,In_1224,In_1935);
or U262 (N_262,In_1977,In_662);
nand U263 (N_263,In_865,In_1877);
and U264 (N_264,In_796,In_18);
and U265 (N_265,In_1819,In_727);
nor U266 (N_266,In_1222,In_1634);
and U267 (N_267,In_1557,In_1898);
nor U268 (N_268,In_36,In_27);
and U269 (N_269,In_632,In_1490);
and U270 (N_270,In_1741,In_1622);
or U271 (N_271,In_613,In_1554);
nand U272 (N_272,In_1640,In_1917);
and U273 (N_273,In_1715,In_1017);
nor U274 (N_274,In_1441,In_873);
and U275 (N_275,In_1566,In_363);
xnor U276 (N_276,In_925,In_1739);
xnor U277 (N_277,In_1027,In_204);
or U278 (N_278,In_1648,In_1263);
xor U279 (N_279,In_1934,In_1016);
xnor U280 (N_280,In_1380,In_9);
and U281 (N_281,In_150,In_449);
or U282 (N_282,In_1138,In_501);
xnor U283 (N_283,In_418,In_1903);
and U284 (N_284,In_747,In_675);
xor U285 (N_285,In_643,In_1057);
and U286 (N_286,In_286,In_1348);
nor U287 (N_287,In_84,In_915);
nor U288 (N_288,In_929,In_1333);
xor U289 (N_289,In_1841,In_21);
nor U290 (N_290,In_991,In_731);
nand U291 (N_291,In_481,In_460);
and U292 (N_292,In_292,In_265);
or U293 (N_293,In_1456,In_1843);
or U294 (N_294,In_1290,In_1530);
nand U295 (N_295,In_1459,In_1269);
nor U296 (N_296,In_375,In_702);
or U297 (N_297,In_81,In_724);
nor U298 (N_298,In_1403,In_1274);
xor U299 (N_299,In_279,In_1418);
xnor U300 (N_300,In_1287,In_403);
nand U301 (N_301,In_74,In_373);
nand U302 (N_302,In_1646,In_54);
and U303 (N_303,In_549,In_1734);
nand U304 (N_304,In_489,In_1783);
nand U305 (N_305,In_11,In_1855);
nand U306 (N_306,In_850,In_948);
or U307 (N_307,In_315,In_1034);
and U308 (N_308,In_716,In_1974);
nor U309 (N_309,In_787,In_66);
xnor U310 (N_310,In_1507,In_471);
nor U311 (N_311,In_608,In_1153);
and U312 (N_312,In_1967,In_570);
and U313 (N_313,In_172,In_1415);
nor U314 (N_314,In_138,In_778);
xor U315 (N_315,In_125,In_1858);
or U316 (N_316,In_1558,In_145);
nand U317 (N_317,In_584,In_1689);
nor U318 (N_318,In_212,In_116);
and U319 (N_319,In_409,In_1343);
nor U320 (N_320,In_10,In_1302);
xnor U321 (N_321,In_1408,In_1945);
nor U322 (N_322,In_1060,In_253);
nand U323 (N_323,In_618,In_1505);
or U324 (N_324,In_1946,In_777);
xor U325 (N_325,In_842,In_1590);
and U326 (N_326,In_167,In_337);
nand U327 (N_327,In_1797,In_1717);
xor U328 (N_328,In_13,In_1659);
nor U329 (N_329,In_1848,In_941);
nor U330 (N_330,In_938,In_1936);
or U331 (N_331,In_1575,In_889);
xor U332 (N_332,In_1091,In_556);
or U333 (N_333,In_820,In_530);
or U334 (N_334,In_246,In_1282);
nand U335 (N_335,In_741,In_527);
nand U336 (N_336,In_769,In_1141);
xor U337 (N_337,In_1461,In_121);
nand U338 (N_338,In_652,In_365);
nor U339 (N_339,In_1426,In_42);
nor U340 (N_340,In_1301,In_124);
and U341 (N_341,In_218,In_1204);
or U342 (N_342,In_934,In_1729);
or U343 (N_343,In_1627,In_446);
nand U344 (N_344,In_198,In_1604);
nor U345 (N_345,In_352,In_1097);
nand U346 (N_346,In_1760,In_1245);
and U347 (N_347,In_1015,In_1542);
or U348 (N_348,In_555,In_927);
or U349 (N_349,In_1241,In_615);
and U350 (N_350,In_193,In_723);
xnor U351 (N_351,In_1402,In_1104);
xor U352 (N_352,In_1234,In_1784);
nor U353 (N_353,In_1068,In_133);
nor U354 (N_354,In_573,In_303);
or U355 (N_355,In_1159,In_316);
or U356 (N_356,In_1424,In_654);
nand U357 (N_357,In_1063,In_942);
nor U358 (N_358,In_900,In_637);
and U359 (N_359,In_100,In_1541);
or U360 (N_360,In_853,In_638);
xnor U361 (N_361,In_931,In_1377);
nor U362 (N_362,In_510,In_249);
xor U363 (N_363,In_1844,In_1242);
nand U364 (N_364,In_1191,In_507);
or U365 (N_365,In_1209,In_630);
and U366 (N_366,In_1615,In_1620);
or U367 (N_367,In_1427,In_412);
and U368 (N_368,In_1257,In_289);
xor U369 (N_369,In_1173,In_1656);
and U370 (N_370,In_440,In_1129);
nand U371 (N_371,In_1605,In_1123);
nor U372 (N_372,In_1470,In_997);
nand U373 (N_373,In_661,In_799);
nor U374 (N_374,In_1981,In_1954);
xnor U375 (N_375,In_1239,In_1761);
and U376 (N_376,In_250,In_448);
nor U377 (N_377,In_432,In_342);
nor U378 (N_378,In_1019,In_243);
and U379 (N_379,In_206,In_1562);
xor U380 (N_380,In_579,In_228);
nand U381 (N_381,In_72,In_287);
nor U382 (N_382,In_434,In_1056);
nor U383 (N_383,In_795,In_665);
nor U384 (N_384,In_1956,In_1132);
nand U385 (N_385,In_883,In_44);
nor U386 (N_386,In_1458,In_1691);
xnor U387 (N_387,In_1658,In_746);
nor U388 (N_388,In_881,In_1392);
and U389 (N_389,In_171,In_1747);
nand U390 (N_390,In_1293,In_830);
nand U391 (N_391,In_837,In_1047);
xnor U392 (N_392,In_516,In_1385);
nor U393 (N_393,In_322,In_16);
nand U394 (N_394,In_687,In_1077);
or U395 (N_395,In_308,In_488);
nor U396 (N_396,In_76,In_785);
xor U397 (N_397,In_457,In_1359);
and U398 (N_398,In_1525,In_1457);
nand U399 (N_399,In_1625,In_1684);
nor U400 (N_400,In_1644,In_1943);
xnor U401 (N_401,In_1477,In_1205);
or U402 (N_402,In_784,In_1581);
nor U403 (N_403,In_512,In_1701);
or U404 (N_404,In_1225,In_946);
nor U405 (N_405,In_1267,In_222);
nor U406 (N_406,In_1712,In_701);
or U407 (N_407,In_214,In_646);
or U408 (N_408,In_1548,In_696);
or U409 (N_409,In_65,In_178);
and U410 (N_410,In_428,In_450);
nor U411 (N_411,In_486,In_572);
and U412 (N_412,In_1965,In_419);
nand U413 (N_413,In_268,In_32);
or U414 (N_414,In_1959,In_185);
nor U415 (N_415,In_151,In_232);
or U416 (N_416,In_789,In_920);
xor U417 (N_417,In_774,In_1009);
xor U418 (N_418,In_326,In_583);
or U419 (N_419,In_1315,In_1028);
nand U420 (N_420,In_1680,In_1192);
or U421 (N_421,In_1406,In_217);
or U422 (N_422,In_974,In_98);
nand U423 (N_423,In_858,In_999);
or U424 (N_424,In_1478,In_715);
nor U425 (N_425,In_1573,In_1154);
nand U426 (N_426,In_1156,In_411);
or U427 (N_427,In_798,In_1454);
xnor U428 (N_428,In_519,In_1678);
and U429 (N_429,In_1174,In_1940);
nand U430 (N_430,In_323,In_1358);
and U431 (N_431,In_695,In_1162);
xnor U432 (N_432,In_770,In_1907);
and U433 (N_433,In_1719,In_1724);
and U434 (N_434,In_825,In_117);
and U435 (N_435,In_5,In_1951);
nand U436 (N_436,In_495,In_321);
xor U437 (N_437,In_1510,In_1531);
or U438 (N_438,In_1878,In_1928);
or U439 (N_439,In_973,In_1004);
nor U440 (N_440,In_1722,In_1771);
or U441 (N_441,In_680,In_1949);
xnor U442 (N_442,In_1617,In_1422);
or U443 (N_443,In_1007,In_1421);
and U444 (N_444,In_1042,In_1961);
or U445 (N_445,In_536,In_1862);
nor U446 (N_446,In_1353,In_1334);
and U447 (N_447,In_589,In_1219);
nand U448 (N_448,In_1258,In_86);
nor U449 (N_449,In_1374,In_1083);
xnor U450 (N_450,In_913,In_1690);
xnor U451 (N_451,In_1344,In_174);
nand U452 (N_452,In_968,In_1608);
or U453 (N_453,In_698,In_1197);
and U454 (N_454,In_438,In_240);
nand U455 (N_455,In_1519,In_560);
and U456 (N_456,In_1732,In_764);
nor U457 (N_457,In_1299,In_1052);
nor U458 (N_458,In_550,In_357);
xor U459 (N_459,In_1306,In_1764);
and U460 (N_460,In_332,In_581);
nor U461 (N_461,In_1157,In_783);
or U462 (N_462,In_1349,In_1466);
xor U463 (N_463,In_558,In_1802);
and U464 (N_464,In_1645,In_372);
xor U465 (N_465,In_952,In_1790);
or U466 (N_466,In_755,In_1890);
nand U467 (N_467,In_605,In_491);
nor U468 (N_468,In_180,In_1297);
nor U469 (N_469,In_749,In_181);
and U470 (N_470,In_890,In_1526);
nand U471 (N_471,In_108,In_984);
nor U472 (N_472,In_1831,In_370);
and U473 (N_473,In_1200,In_1978);
nand U474 (N_474,In_1247,In_544);
or U475 (N_475,In_1423,In_1093);
nor U476 (N_476,In_1360,In_106);
or U477 (N_477,In_1864,In_227);
and U478 (N_478,In_1473,In_713);
nand U479 (N_479,In_305,In_1833);
nor U480 (N_480,In_1988,In_737);
nand U481 (N_481,In_1033,In_1758);
or U482 (N_482,In_1050,In_1990);
or U483 (N_483,In_547,In_966);
and U484 (N_484,In_1160,In_1657);
or U485 (N_485,In_645,In_1593);
nor U486 (N_486,In_1808,In_1233);
xor U487 (N_487,In_53,In_1816);
nand U488 (N_488,In_59,In_158);
or U489 (N_489,In_1496,In_1971);
xnor U490 (N_490,In_528,In_122);
nor U491 (N_491,In_600,In_1675);
or U492 (N_492,In_3,In_1000);
and U493 (N_493,In_1555,In_1708);
nor U494 (N_494,In_169,In_1102);
nand U495 (N_495,In_754,In_563);
and U496 (N_496,In_1407,In_334);
and U497 (N_497,In_856,In_1942);
or U498 (N_498,In_1149,In_324);
nor U499 (N_499,In_762,In_498);
nor U500 (N_500,In_1572,In_1537);
xor U501 (N_501,In_792,In_380);
and U502 (N_502,In_923,In_735);
xor U503 (N_503,In_1750,In_190);
nand U504 (N_504,In_1410,In_1539);
or U505 (N_505,In_1972,In_1054);
or U506 (N_506,In_1146,In_1323);
nor U507 (N_507,In_953,In_295);
or U508 (N_508,In_1707,In_874);
nand U509 (N_509,In_1804,In_722);
nor U510 (N_510,In_1740,In_976);
nor U511 (N_511,In_1080,In_83);
and U512 (N_512,In_1851,In_766);
or U513 (N_513,In_1511,In_1130);
or U514 (N_514,In_1142,In_1316);
nor U515 (N_515,In_587,In_320);
and U516 (N_516,In_995,In_603);
and U517 (N_517,In_1250,In_1262);
xnor U518 (N_518,In_870,In_176);
and U519 (N_519,In_1126,In_1957);
nor U520 (N_520,In_704,In_975);
nor U521 (N_521,In_1748,In_1682);
and U522 (N_522,In_104,In_1973);
nand U523 (N_523,In_402,In_811);
and U524 (N_524,In_1328,In_1070);
nor U525 (N_525,In_1567,In_1937);
nand U526 (N_526,In_236,In_1688);
and U527 (N_527,In_336,In_465);
nand U528 (N_528,In_313,In_1914);
and U529 (N_529,In_8,In_1498);
xor U530 (N_530,In_1711,In_1175);
and U531 (N_531,In_93,In_780);
xnor U532 (N_532,In_1202,In_1125);
xor U533 (N_533,In_1769,In_1897);
nand U534 (N_534,In_1317,In_262);
or U535 (N_535,In_1782,In_309);
xor U536 (N_536,In_1181,In_1964);
xor U537 (N_537,In_1002,In_179);
or U538 (N_538,In_744,In_1464);
xnor U539 (N_539,In_1662,In_304);
and U540 (N_540,In_980,In_73);
xnor U541 (N_541,In_1650,In_1610);
xor U542 (N_542,In_1483,In_1288);
or U543 (N_543,In_126,In_1594);
xor U544 (N_544,In_341,In_1006);
xnor U545 (N_545,In_1005,In_947);
nand U546 (N_546,In_678,In_351);
nand U547 (N_547,In_1151,In_1696);
nand U548 (N_548,In_229,In_1868);
nand U549 (N_549,In_280,In_1279);
nand U550 (N_550,In_1697,In_1814);
and U551 (N_551,In_836,In_585);
or U552 (N_552,In_921,In_496);
and U553 (N_553,In_355,In_466);
and U554 (N_554,In_441,In_1218);
and U555 (N_555,In_1516,In_1870);
or U556 (N_556,In_1136,In_738);
nand U557 (N_557,In_56,In_364);
nor U558 (N_558,In_1975,In_1654);
nor U559 (N_559,In_905,In_887);
nor U560 (N_560,In_788,In_707);
nand U561 (N_561,In_436,In_879);
xnor U562 (N_562,In_649,In_1902);
xnor U563 (N_563,In_1875,In_781);
nand U564 (N_564,In_1296,In_377);
or U565 (N_565,In_1228,In_1393);
nor U566 (N_566,In_1666,In_672);
and U567 (N_567,In_94,In_1731);
and U568 (N_568,In_884,In_916);
xor U569 (N_569,In_1281,In_1442);
nor U570 (N_570,In_1705,In_343);
nor U571 (N_571,In_1035,In_237);
nand U572 (N_572,In_423,In_269);
nand U573 (N_573,In_311,In_1553);
and U574 (N_574,In_191,In_1861);
or U575 (N_575,In_1036,In_1738);
xor U576 (N_576,In_1253,In_1906);
xnor U577 (N_577,In_1217,In_1468);
nand U578 (N_578,In_105,In_508);
nand U579 (N_579,In_580,In_1079);
or U580 (N_580,In_802,In_1801);
nor U581 (N_581,In_972,In_1584);
nand U582 (N_582,In_330,In_187);
xnor U583 (N_583,In_1309,In_860);
and U584 (N_584,In_1859,In_663);
nand U585 (N_585,In_998,In_954);
xor U586 (N_586,In_1337,In_1651);
xor U587 (N_587,In_1509,In_772);
or U588 (N_588,In_899,In_1779);
and U589 (N_589,In_1113,In_1240);
nor U590 (N_590,In_1347,In_1331);
nand U591 (N_591,In_414,In_338);
or U592 (N_592,In_1649,In_686);
xor U593 (N_593,In_1931,In_47);
xor U594 (N_594,In_1742,In_290);
or U595 (N_595,In_483,In_539);
xnor U596 (N_596,In_867,In_1836);
or U597 (N_597,In_639,In_328);
nand U598 (N_598,In_405,In_743);
nor U599 (N_599,In_85,In_1227);
and U600 (N_600,In_1735,In_1638);
nand U601 (N_601,In_194,In_1669);
nand U602 (N_602,In_813,In_1927);
or U603 (N_603,In_41,In_1476);
nand U604 (N_604,In_1796,In_728);
nand U605 (N_605,In_937,In_92);
or U606 (N_606,In_1046,In_611);
nand U607 (N_607,In_1730,In_456);
or U608 (N_608,In_880,In_801);
or U609 (N_609,In_115,In_339);
nand U610 (N_610,In_1785,In_404);
and U611 (N_611,In_69,In_1789);
and U612 (N_612,In_1329,In_435);
or U613 (N_613,In_1571,In_1552);
and U614 (N_614,In_1772,In_1926);
xor U615 (N_615,In_1702,In_318);
nor U616 (N_616,In_1107,In_37);
nand U617 (N_617,In_327,In_1938);
and U618 (N_618,In_1469,In_1623);
nor U619 (N_619,In_882,In_1445);
nor U620 (N_620,In_445,In_621);
xnor U621 (N_621,In_443,In_1419);
or U622 (N_622,In_1574,In_908);
nand U623 (N_623,In_1292,In_1930);
xnor U624 (N_624,In_1893,In_1806);
and U625 (N_625,In_1318,In_1811);
or U626 (N_626,In_220,In_381);
nand U627 (N_627,In_302,In_1183);
xnor U628 (N_628,In_223,In_815);
or U629 (N_629,In_1874,In_1815);
xor U630 (N_630,In_356,In_1020);
nor U631 (N_631,In_1455,In_1158);
xnor U632 (N_632,In_1591,In_299);
xor U633 (N_633,In_521,In_361);
xnor U634 (N_634,In_300,In_1355);
and U635 (N_635,In_617,In_1480);
xor U636 (N_636,In_1433,In_1214);
nand U637 (N_637,In_397,In_844);
or U638 (N_638,In_838,In_252);
nand U639 (N_639,In_1986,In_523);
xor U640 (N_640,In_1314,In_1145);
or U641 (N_641,In_396,In_1820);
and U642 (N_642,In_80,In_1979);
xnor U643 (N_643,In_1055,In_1985);
nor U644 (N_644,In_400,In_360);
nor U645 (N_645,In_857,In_1733);
and U646 (N_646,In_1067,In_1547);
and U647 (N_647,In_824,In_1078);
nand U648 (N_648,In_358,In_854);
nor U649 (N_649,In_797,In_1500);
or U650 (N_650,In_595,In_1621);
or U651 (N_651,In_209,In_775);
nand U652 (N_652,In_442,In_1165);
and U653 (N_653,In_1752,In_1003);
or U654 (N_654,In_1989,In_733);
xnor U655 (N_655,In_689,In_936);
and U656 (N_656,In_878,In_1628);
nor U657 (N_657,In_1172,In_1339);
or U658 (N_658,In_278,In_1759);
nand U659 (N_659,In_1075,In_626);
nor U660 (N_660,In_285,In_1298);
nor U661 (N_661,In_1342,In_871);
nor U662 (N_662,In_46,In_485);
xor U663 (N_663,In_1177,In_1235);
nor U664 (N_664,In_111,In_170);
and U665 (N_665,In_1304,In_29);
and U666 (N_666,In_1794,In_469);
xor U667 (N_667,In_1924,In_1800);
nor U668 (N_668,In_851,In_1853);
nor U669 (N_669,In_848,In_288);
nor U670 (N_670,In_633,In_1867);
or U671 (N_671,In_1583,In_186);
and U672 (N_672,In_841,In_1535);
and U673 (N_673,In_1382,In_1939);
and U674 (N_674,In_1308,In_956);
xnor U675 (N_675,In_897,In_779);
nor U676 (N_676,In_1580,In_345);
and U677 (N_677,In_1065,In_1086);
or U678 (N_678,In_740,In_1221);
nand U679 (N_679,In_835,In_271);
or U680 (N_680,In_467,In_1092);
or U681 (N_681,In_1889,In_886);
nand U682 (N_682,In_647,In_1664);
xor U683 (N_683,In_719,In_1322);
xor U684 (N_684,In_1276,In_1285);
nand U685 (N_685,In_599,In_1026);
xor U686 (N_686,In_505,In_1933);
or U687 (N_687,In_979,In_1340);
nor U688 (N_688,In_99,In_1929);
nor U689 (N_689,In_996,In_1112);
xnor U690 (N_690,In_153,In_1411);
or U691 (N_691,In_1109,In_1324);
or U692 (N_692,In_641,In_960);
and U693 (N_693,In_1805,In_2);
nand U694 (N_694,In_607,In_1025);
nand U695 (N_695,In_685,In_1881);
and U696 (N_696,In_224,In_1391);
nand U697 (N_697,In_298,In_353);
nand U698 (N_698,In_620,In_776);
nor U699 (N_699,In_951,In_1465);
and U700 (N_700,In_1090,In_1082);
xnor U701 (N_701,In_1429,In_1148);
xnor U702 (N_702,In_1647,In_1960);
nand U703 (N_703,In_156,In_911);
and U704 (N_704,In_493,In_598);
nor U705 (N_705,In_651,In_1367);
xor U706 (N_706,In_1770,In_335);
nor U707 (N_707,In_1244,In_877);
and U708 (N_708,In_272,In_1589);
nor U709 (N_709,In_1533,In_763);
nand U710 (N_710,In_804,In_718);
nor U711 (N_711,In_526,In_1982);
and U712 (N_712,In_511,In_1030);
xnor U713 (N_713,In_868,In_514);
xnor U714 (N_714,In_1341,In_1486);
nor U715 (N_715,In_1602,In_869);
nand U716 (N_716,In_160,In_791);
and U717 (N_717,In_1720,In_576);
xor U718 (N_718,In_1117,In_711);
xnor U719 (N_719,In_669,In_628);
nand U720 (N_720,In_906,In_162);
and U721 (N_721,In_1865,In_1170);
or U722 (N_722,In_1766,In_1378);
nand U723 (N_723,In_1749,In_1326);
nor U724 (N_724,In_454,In_812);
and U725 (N_725,In_1600,In_1345);
nand U726 (N_726,In_401,In_1430);
or U727 (N_727,In_506,In_374);
nand U728 (N_728,In_1076,In_1879);
nand U729 (N_729,In_201,In_1698);
xnor U730 (N_730,In_1066,In_1636);
or U731 (N_731,In_470,In_91);
and U732 (N_732,In_767,In_1305);
xor U733 (N_733,In_855,In_1095);
nand U734 (N_734,In_1842,In_866);
or U735 (N_735,In_816,In_1963);
xor U736 (N_736,In_329,In_1606);
or U737 (N_737,In_1631,In_1167);
or U738 (N_738,In_1776,In_1064);
or U739 (N_739,In_1920,In_668);
or U740 (N_740,In_504,In_1996);
nand U741 (N_741,In_333,In_346);
and U742 (N_742,In_1186,In_1671);
and U743 (N_743,In_847,In_143);
nor U744 (N_744,In_1570,In_45);
and U745 (N_745,In_1460,In_1686);
nor U746 (N_746,In_1660,In_902);
xor U747 (N_747,In_759,In_472);
and U748 (N_748,In_26,In_70);
or U749 (N_749,In_609,In_1703);
nor U750 (N_750,In_1559,In_985);
or U751 (N_751,In_1966,In_310);
or U752 (N_752,In_118,In_325);
and U753 (N_753,In_1049,In_552);
or U754 (N_754,In_1449,In_1368);
xnor U755 (N_755,In_1363,In_983);
nor U756 (N_756,In_1237,In_1932);
or U757 (N_757,In_993,In_119);
nand U758 (N_758,In_1040,In_461);
nor U759 (N_759,In_1768,In_203);
nor U760 (N_760,In_213,In_568);
nand U761 (N_761,In_238,In_1260);
and U762 (N_762,In_1283,In_1272);
and U763 (N_763,In_756,In_875);
and U764 (N_764,In_659,In_216);
or U765 (N_765,In_147,In_1892);
nor U766 (N_766,In_87,In_477);
and U767 (N_767,In_24,In_1361);
or U768 (N_768,In_708,In_944);
xnor U769 (N_769,In_627,In_1674);
and U770 (N_770,In_1398,In_712);
nor U771 (N_771,In_932,In_1432);
and U772 (N_772,In_541,In_1278);
and U773 (N_773,In_1692,In_1821);
xnor U774 (N_774,In_1826,In_1350);
and U775 (N_775,In_1835,In_1512);
nand U776 (N_776,In_1912,In_989);
or U777 (N_777,In_413,In_1616);
and U778 (N_778,In_533,In_1236);
nor U779 (N_779,In_1672,In_15);
xnor U780 (N_780,In_1199,In_1683);
or U781 (N_781,In_1037,In_800);
and U782 (N_782,In_614,In_845);
or U783 (N_783,In_509,In_1987);
nor U784 (N_784,In_1544,In_1983);
and U785 (N_785,In_683,In_17);
or U786 (N_786,In_1369,In_671);
or U787 (N_787,In_1238,In_487);
or U788 (N_788,In_1633,In_1451);
xnor U789 (N_789,In_1780,In_439);
xor U790 (N_790,In_545,In_1736);
xnor U791 (N_791,In_1754,In_1439);
xnor U792 (N_792,In_1474,In_559);
nor U793 (N_793,In_60,In_1655);
nand U794 (N_794,In_95,In_1155);
nand U795 (N_795,In_1273,In_1127);
and U796 (N_796,In_922,In_1492);
or U797 (N_797,In_540,In_1970);
nand U798 (N_798,In_757,In_31);
nor U799 (N_799,In_1417,In_1084);
nor U800 (N_800,In_833,In_1321);
and U801 (N_801,In_1991,In_673);
nand U802 (N_802,In_1396,In_1452);
nor U803 (N_803,In_1058,In_1586);
nand U804 (N_804,In_1096,In_1352);
and U805 (N_805,In_1915,In_760);
nor U806 (N_806,In_1495,In_462);
nor U807 (N_807,In_149,In_575);
xnor U808 (N_808,In_1428,In_970);
xor U809 (N_809,In_706,In_388);
nor U810 (N_810,In_803,In_1832);
and U811 (N_811,In_640,In_919);
nor U812 (N_812,In_843,In_1335);
xnor U813 (N_813,In_531,In_173);
xor U814 (N_814,In_282,In_1545);
nand U815 (N_815,In_1838,In_142);
nand U816 (N_816,In_1206,In_904);
and U817 (N_817,In_1774,In_444);
or U818 (N_818,In_656,In_1743);
nand U819 (N_819,In_113,In_1506);
nor U820 (N_820,In_1641,In_574);
and U821 (N_821,In_1614,In_1652);
and U822 (N_822,In_786,In_758);
xnor U823 (N_823,In_1839,In_1212);
or U824 (N_824,In_586,In_140);
nor U825 (N_825,In_725,In_748);
nand U826 (N_826,In_1871,In_699);
nor U827 (N_827,In_410,In_525);
or U828 (N_828,In_421,In_1522);
nor U829 (N_829,In_263,In_408);
and U830 (N_830,In_1259,In_1038);
or U831 (N_831,In_75,In_1053);
nor U832 (N_832,In_189,In_677);
or U833 (N_833,In_429,In_562);
xnor U834 (N_834,In_251,In_497);
and U835 (N_835,In_1781,In_1630);
xnor U836 (N_836,In_939,In_1909);
and U837 (N_837,In_1012,In_965);
and U838 (N_838,In_565,In_82);
or U839 (N_839,In_274,In_1493);
or U840 (N_840,In_831,In_447);
or U841 (N_841,In_839,In_1232);
and U842 (N_842,In_51,In_709);
xnor U843 (N_843,In_1436,In_935);
nor U844 (N_844,In_622,In_492);
xnor U845 (N_845,In_534,In_945);
and U846 (N_846,In_200,In_241);
or U847 (N_847,In_225,In_988);
or U848 (N_848,In_994,In_33);
and U849 (N_849,In_1997,In_1087);
nor U850 (N_850,In_1725,In_1565);
xnor U851 (N_851,In_1045,In_1830);
or U852 (N_852,In_205,In_917);
or U853 (N_853,In_1714,In_1755);
xnor U854 (N_854,In_697,In_6);
and U855 (N_855,In_1869,In_790);
nor U856 (N_856,In_1829,In_1948);
xnor U857 (N_857,In_1425,In_1243);
xnor U858 (N_858,In_1866,In_1556);
nor U859 (N_859,In_102,In_275);
or U860 (N_860,In_903,In_78);
or U861 (N_861,In_1485,In_427);
or U862 (N_862,In_90,In_1695);
or U863 (N_863,In_1911,In_25);
or U864 (N_864,In_1538,In_52);
and U865 (N_865,In_1375,In_1840);
nand U866 (N_866,In_1601,In_688);
xor U867 (N_867,In_593,In_542);
or U868 (N_868,In_1597,In_175);
nand U869 (N_869,In_273,In_1679);
nor U870 (N_870,In_89,In_872);
nor U871 (N_871,In_256,In_152);
nor U872 (N_872,In_1021,In_1435);
and U873 (N_873,In_1185,In_691);
xor U874 (N_874,In_1887,In_1810);
and U875 (N_875,In_635,In_1431);
or U876 (N_876,In_1895,In_340);
and U877 (N_877,In_1164,In_391);
or U878 (N_878,In_1179,In_1313);
and U879 (N_879,In_1381,In_177);
nand U880 (N_880,In_1860,In_1885);
nor U881 (N_881,In_459,In_1203);
or U882 (N_882,In_1952,In_166);
or U883 (N_883,In_1216,In_529);
xor U884 (N_884,In_146,In_7);
nand U885 (N_885,In_1818,In_546);
or U886 (N_886,In_1489,In_717);
and U887 (N_887,In_1588,In_1178);
nor U888 (N_888,In_636,In_1534);
nand U889 (N_889,In_20,In_1995);
nor U890 (N_890,In_1823,In_306);
or U891 (N_891,In_616,In_1416);
xnor U892 (N_892,In_14,In_1629);
and U893 (N_893,In_1578,In_196);
nor U894 (N_894,In_426,In_805);
and U895 (N_895,In_248,In_648);
or U896 (N_896,In_1497,In_1799);
or U897 (N_897,In_19,In_732);
nand U898 (N_898,In_910,In_234);
xnor U899 (N_899,In_1444,In_692);
nor U900 (N_900,In_183,In_1502);
nand U901 (N_901,In_1568,In_1564);
or U902 (N_902,In_1187,In_221);
and U903 (N_903,In_682,In_1876);
xnor U904 (N_904,In_1947,In_826);
or U905 (N_905,In_283,In_1550);
or U906 (N_906,In_387,In_978);
xor U907 (N_907,In_1370,In_1762);
nand U908 (N_908,In_1271,In_1252);
or U909 (N_909,In_1379,In_1386);
nand U910 (N_910,In_1665,In_1813);
xnor U911 (N_911,In_1397,In_314);
nand U912 (N_912,In_846,In_1778);
and U913 (N_913,In_1264,In_210);
and U914 (N_914,In_1685,In_959);
xor U915 (N_915,In_619,In_933);
xor U916 (N_916,In_1280,In_773);
nand U917 (N_917,In_1856,In_703);
or U918 (N_918,In_1011,In_1152);
and U919 (N_919,In_1268,In_242);
nand U920 (N_920,In_961,In_110);
or U921 (N_921,In_1409,In_494);
nor U922 (N_922,In_354,In_1122);
nand U923 (N_923,In_1795,In_1763);
nor U924 (N_924,In_1798,In_1365);
or U925 (N_925,In_1713,In_424);
xor U926 (N_926,In_1106,In_1514);
nor U927 (N_927,In_987,In_1190);
nand U928 (N_928,In_451,In_55);
and U929 (N_929,In_1582,In_623);
nand U930 (N_930,In_604,In_155);
and U931 (N_931,In_1560,In_261);
or U932 (N_932,In_564,In_1677);
nor U933 (N_933,In_765,In_876);
and U934 (N_934,In_464,In_819);
or U935 (N_935,In_1405,In_1024);
nand U936 (N_936,In_1807,In_417);
or U937 (N_937,In_548,In_1676);
and U938 (N_938,In_1721,In_1482);
nand U939 (N_939,In_350,In_1098);
and U940 (N_940,In_901,In_1726);
or U941 (N_941,In_1119,In_1487);
nor U942 (N_942,In_1901,In_1105);
nand U943 (N_943,In_1039,In_215);
nand U944 (N_944,In_1184,In_77);
nor U945 (N_945,In_888,In_1248);
nand U946 (N_946,In_1888,In_828);
nand U947 (N_947,In_1569,In_43);
nor U948 (N_948,In_578,In_1837);
nand U949 (N_949,In_992,In_1366);
nor U950 (N_950,In_1824,In_1229);
nor U951 (N_951,In_1434,In_1607);
xor U952 (N_952,In_1599,In_631);
or U953 (N_953,In_109,In_1099);
nand U954 (N_954,In_625,In_34);
or U955 (N_955,In_817,In_1420);
and U956 (N_956,In_594,In_1022);
or U957 (N_957,In_1913,In_834);
xnor U958 (N_958,In_331,In_1706);
or U959 (N_959,In_219,In_1383);
nand U960 (N_960,In_1693,In_924);
xor U961 (N_961,In_1751,In_971);
nand U962 (N_962,In_1619,In_1462);
and U963 (N_963,In_967,In_79);
nor U964 (N_964,In_601,In_1543);
and U965 (N_965,In_1062,In_88);
nand U966 (N_966,In_1694,In_1450);
or U967 (N_967,In_794,In_255);
nand U968 (N_968,In_437,In_1230);
xnor U969 (N_969,In_1115,In_1001);
nand U970 (N_970,In_949,In_1812);
nor U971 (N_971,In_1792,In_1208);
nor U972 (N_972,In_395,In_136);
and U973 (N_973,In_1637,In_694);
nand U974 (N_974,In_1387,In_1955);
and U975 (N_975,In_416,In_818);
nor U976 (N_976,In_1163,In_230);
nand U977 (N_977,In_141,In_891);
and U978 (N_978,In_50,In_1188);
or U979 (N_979,In_38,In_674);
and U980 (N_980,In_957,In_1528);
and U981 (N_981,In_517,In_729);
nand U982 (N_982,In_0,In_1372);
or U983 (N_983,In_893,In_1579);
or U984 (N_984,In_1999,In_503);
nor U985 (N_985,In_896,In_1639);
and U986 (N_986,In_277,In_734);
nor U987 (N_987,In_468,In_1166);
and U988 (N_988,In_1336,In_1521);
nand U989 (N_989,In_1626,In_482);
or U990 (N_990,In_407,In_721);
and U991 (N_991,In_1984,In_233);
and U992 (N_992,In_1925,In_1787);
nor U993 (N_993,In_1523,In_1704);
and U994 (N_994,In_1791,In_1312);
nand U995 (N_995,In_226,In_163);
or U996 (N_996,In_969,In_1598);
nand U997 (N_997,In_745,In_1549);
and U998 (N_998,In_1193,In_1609);
nor U999 (N_999,In_561,In_112);
nand U1000 (N_1000,N_68,N_57);
and U1001 (N_1001,N_534,N_742);
or U1002 (N_1002,N_42,N_712);
nand U1003 (N_1003,N_190,N_448);
and U1004 (N_1004,N_917,N_199);
or U1005 (N_1005,N_375,N_855);
nand U1006 (N_1006,N_601,N_37);
and U1007 (N_1007,N_876,N_619);
or U1008 (N_1008,N_966,N_890);
and U1009 (N_1009,N_850,N_512);
and U1010 (N_1010,N_571,N_660);
and U1011 (N_1011,N_752,N_803);
or U1012 (N_1012,N_854,N_10);
and U1013 (N_1013,N_411,N_615);
or U1014 (N_1014,N_973,N_170);
nand U1015 (N_1015,N_406,N_428);
nand U1016 (N_1016,N_441,N_185);
nand U1017 (N_1017,N_487,N_54);
and U1018 (N_1018,N_419,N_169);
and U1019 (N_1019,N_272,N_904);
nor U1020 (N_1020,N_330,N_447);
or U1021 (N_1021,N_520,N_50);
and U1022 (N_1022,N_969,N_596);
xnor U1023 (N_1023,N_344,N_664);
nand U1024 (N_1024,N_47,N_777);
xnor U1025 (N_1025,N_8,N_795);
nand U1026 (N_1026,N_705,N_907);
or U1027 (N_1027,N_390,N_912);
xor U1028 (N_1028,N_178,N_3);
xnor U1029 (N_1029,N_131,N_298);
or U1030 (N_1030,N_933,N_519);
or U1031 (N_1031,N_654,N_55);
and U1032 (N_1032,N_453,N_893);
nand U1033 (N_1033,N_176,N_704);
nand U1034 (N_1034,N_460,N_463);
and U1035 (N_1035,N_840,N_322);
nor U1036 (N_1036,N_783,N_767);
nand U1037 (N_1037,N_565,N_835);
xor U1038 (N_1038,N_799,N_814);
and U1039 (N_1039,N_155,N_276);
and U1040 (N_1040,N_680,N_924);
xor U1041 (N_1041,N_147,N_386);
xor U1042 (N_1042,N_96,N_584);
nand U1043 (N_1043,N_314,N_834);
nor U1044 (N_1044,N_58,N_655);
or U1045 (N_1045,N_533,N_246);
and U1046 (N_1046,N_343,N_241);
nand U1047 (N_1047,N_837,N_122);
xnor U1048 (N_1048,N_184,N_320);
or U1049 (N_1049,N_726,N_354);
nand U1050 (N_1050,N_616,N_825);
and U1051 (N_1051,N_93,N_938);
and U1052 (N_1052,N_336,N_380);
nand U1053 (N_1053,N_543,N_427);
and U1054 (N_1054,N_388,N_225);
nor U1055 (N_1055,N_323,N_807);
and U1056 (N_1056,N_724,N_468);
nand U1057 (N_1057,N_217,N_686);
or U1058 (N_1058,N_983,N_20);
nand U1059 (N_1059,N_793,N_670);
nor U1060 (N_1060,N_366,N_668);
xor U1061 (N_1061,N_171,N_945);
nor U1062 (N_1062,N_236,N_667);
nand U1063 (N_1063,N_977,N_243);
xnor U1064 (N_1064,N_549,N_501);
nand U1065 (N_1065,N_963,N_905);
nand U1066 (N_1066,N_162,N_770);
nor U1067 (N_1067,N_639,N_101);
and U1068 (N_1068,N_226,N_317);
nand U1069 (N_1069,N_237,N_947);
nand U1070 (N_1070,N_315,N_651);
or U1071 (N_1071,N_551,N_598);
and U1072 (N_1072,N_249,N_385);
and U1073 (N_1073,N_9,N_896);
nor U1074 (N_1074,N_577,N_284);
nand U1075 (N_1075,N_245,N_14);
or U1076 (N_1076,N_949,N_987);
and U1077 (N_1077,N_262,N_497);
and U1078 (N_1078,N_177,N_698);
nand U1079 (N_1079,N_785,N_479);
or U1080 (N_1080,N_418,N_197);
or U1081 (N_1081,N_701,N_989);
and U1082 (N_1082,N_346,N_73);
and U1083 (N_1083,N_493,N_283);
nand U1084 (N_1084,N_721,N_400);
nand U1085 (N_1085,N_474,N_306);
xor U1086 (N_1086,N_557,N_454);
and U1087 (N_1087,N_863,N_558);
xor U1088 (N_1088,N_473,N_700);
and U1089 (N_1089,N_786,N_656);
nor U1090 (N_1090,N_791,N_163);
nor U1091 (N_1091,N_848,N_653);
nand U1092 (N_1092,N_796,N_477);
xor U1093 (N_1093,N_142,N_729);
and U1094 (N_1094,N_23,N_426);
nor U1095 (N_1095,N_342,N_117);
nor U1096 (N_1096,N_504,N_674);
xor U1097 (N_1097,N_295,N_164);
and U1098 (N_1098,N_393,N_148);
or U1099 (N_1099,N_864,N_90);
or U1100 (N_1100,N_188,N_451);
and U1101 (N_1101,N_383,N_125);
nor U1102 (N_1102,N_608,N_260);
and U1103 (N_1103,N_970,N_561);
and U1104 (N_1104,N_467,N_110);
nor U1105 (N_1105,N_693,N_285);
xnor U1106 (N_1106,N_340,N_156);
xnor U1107 (N_1107,N_205,N_351);
nand U1108 (N_1108,N_921,N_114);
and U1109 (N_1109,N_648,N_416);
or U1110 (N_1110,N_939,N_613);
xor U1111 (N_1111,N_990,N_361);
xnor U1112 (N_1112,N_529,N_830);
or U1113 (N_1113,N_89,N_845);
xnor U1114 (N_1114,N_51,N_684);
nand U1115 (N_1115,N_46,N_365);
nand U1116 (N_1116,N_919,N_564);
and U1117 (N_1117,N_646,N_822);
xnor U1118 (N_1118,N_301,N_682);
or U1119 (N_1119,N_918,N_76);
xnor U1120 (N_1120,N_768,N_310);
nand U1121 (N_1121,N_761,N_254);
or U1122 (N_1122,N_95,N_161);
or U1123 (N_1123,N_847,N_82);
nor U1124 (N_1124,N_488,N_815);
nor U1125 (N_1125,N_457,N_494);
nand U1126 (N_1126,N_778,N_997);
nand U1127 (N_1127,N_934,N_797);
nand U1128 (N_1128,N_103,N_112);
or U1129 (N_1129,N_787,N_157);
nor U1130 (N_1130,N_431,N_857);
and U1131 (N_1131,N_79,N_720);
nand U1132 (N_1132,N_6,N_374);
and U1133 (N_1133,N_688,N_287);
and U1134 (N_1134,N_52,N_935);
and U1135 (N_1135,N_749,N_600);
xnor U1136 (N_1136,N_137,N_308);
nor U1137 (N_1137,N_300,N_327);
and U1138 (N_1138,N_874,N_376);
and U1139 (N_1139,N_649,N_925);
nand U1140 (N_1140,N_647,N_193);
xor U1141 (N_1141,N_542,N_572);
nor U1142 (N_1142,N_620,N_811);
nand U1143 (N_1143,N_610,N_221);
xor U1144 (N_1144,N_207,N_747);
nand U1145 (N_1145,N_339,N_717);
and U1146 (N_1146,N_806,N_515);
and U1147 (N_1147,N_633,N_115);
xor U1148 (N_1148,N_422,N_63);
or U1149 (N_1149,N_192,N_500);
xnor U1150 (N_1150,N_402,N_818);
nor U1151 (N_1151,N_303,N_823);
and U1152 (N_1152,N_508,N_470);
and U1153 (N_1153,N_434,N_191);
xnor U1154 (N_1154,N_420,N_444);
or U1155 (N_1155,N_930,N_991);
nor U1156 (N_1156,N_370,N_862);
xnor U1157 (N_1157,N_92,N_695);
or U1158 (N_1158,N_59,N_491);
nor U1159 (N_1159,N_732,N_663);
or U1160 (N_1160,N_84,N_524);
and U1161 (N_1161,N_410,N_461);
nor U1162 (N_1162,N_526,N_265);
or U1163 (N_1163,N_395,N_34);
xor U1164 (N_1164,N_439,N_540);
and U1165 (N_1165,N_291,N_134);
nor U1166 (N_1166,N_946,N_979);
and U1167 (N_1167,N_809,N_452);
nand U1168 (N_1168,N_1,N_556);
nor U1169 (N_1169,N_538,N_774);
nand U1170 (N_1170,N_928,N_546);
and U1171 (N_1171,N_999,N_319);
xor U1172 (N_1172,N_903,N_658);
and U1173 (N_1173,N_296,N_527);
nand U1174 (N_1174,N_897,N_634);
nand U1175 (N_1175,N_861,N_288);
nor U1176 (N_1176,N_708,N_865);
xor U1177 (N_1177,N_817,N_87);
nor U1178 (N_1178,N_91,N_455);
or U1179 (N_1179,N_898,N_77);
nor U1180 (N_1180,N_438,N_880);
or U1181 (N_1181,N_628,N_988);
xor U1182 (N_1182,N_443,N_618);
nand U1183 (N_1183,N_743,N_360);
nor U1184 (N_1184,N_25,N_635);
nor U1185 (N_1185,N_105,N_790);
nor U1186 (N_1186,N_675,N_820);
and U1187 (N_1187,N_812,N_72);
nor U1188 (N_1188,N_212,N_513);
or U1189 (N_1189,N_804,N_703);
and U1190 (N_1190,N_173,N_640);
or U1191 (N_1191,N_259,N_99);
nor U1192 (N_1192,N_17,N_728);
nand U1193 (N_1193,N_216,N_960);
nor U1194 (N_1194,N_588,N_813);
xnor U1195 (N_1195,N_582,N_409);
nor U1196 (N_1196,N_130,N_309);
nor U1197 (N_1197,N_779,N_396);
xnor U1198 (N_1198,N_38,N_430);
or U1199 (N_1199,N_916,N_962);
and U1200 (N_1200,N_40,N_146);
xor U1201 (N_1201,N_127,N_280);
or U1202 (N_1202,N_794,N_614);
xnor U1203 (N_1203,N_44,N_433);
and U1204 (N_1204,N_141,N_516);
nand U1205 (N_1205,N_858,N_875);
nor U1206 (N_1206,N_484,N_626);
or U1207 (N_1207,N_362,N_523);
xor U1208 (N_1208,N_950,N_21);
xor U1209 (N_1209,N_329,N_382);
xor U1210 (N_1210,N_891,N_920);
xnor U1211 (N_1211,N_915,N_328);
nor U1212 (N_1212,N_53,N_222);
nand U1213 (N_1213,N_959,N_716);
or U1214 (N_1214,N_948,N_469);
xnor U1215 (N_1215,N_581,N_78);
nand U1216 (N_1216,N_702,N_100);
nand U1217 (N_1217,N_650,N_405);
nand U1218 (N_1218,N_839,N_61);
and U1219 (N_1219,N_802,N_555);
xnor U1220 (N_1220,N_578,N_19);
nand U1221 (N_1221,N_771,N_56);
xnor U1222 (N_1222,N_364,N_605);
or U1223 (N_1223,N_906,N_776);
xnor U1224 (N_1224,N_294,N_261);
nor U1225 (N_1225,N_681,N_709);
nor U1226 (N_1226,N_311,N_595);
and U1227 (N_1227,N_210,N_168);
and U1228 (N_1228,N_860,N_851);
or U1229 (N_1229,N_894,N_781);
nand U1230 (N_1230,N_394,N_70);
nor U1231 (N_1231,N_609,N_83);
nor U1232 (N_1232,N_580,N_195);
and U1233 (N_1233,N_149,N_174);
and U1234 (N_1234,N_269,N_154);
or U1235 (N_1235,N_186,N_943);
nor U1236 (N_1236,N_982,N_313);
and U1237 (N_1237,N_35,N_60);
xor U1238 (N_1238,N_412,N_741);
nand U1239 (N_1239,N_801,N_631);
or U1240 (N_1240,N_235,N_810);
nor U1241 (N_1241,N_737,N_109);
xor U1242 (N_1242,N_937,N_659);
nor U1243 (N_1243,N_877,N_586);
and U1244 (N_1244,N_363,N_525);
nor U1245 (N_1245,N_445,N_334);
xor U1246 (N_1246,N_119,N_151);
xnor U1247 (N_1247,N_305,N_927);
nor U1248 (N_1248,N_277,N_118);
xnor U1249 (N_1249,N_722,N_4);
and U1250 (N_1250,N_152,N_13);
and U1251 (N_1251,N_872,N_417);
nor U1252 (N_1252,N_45,N_643);
and U1253 (N_1253,N_180,N_392);
or U1254 (N_1254,N_889,N_942);
or U1255 (N_1255,N_532,N_331);
nor U1256 (N_1256,N_81,N_636);
or U1257 (N_1257,N_97,N_414);
xnor U1258 (N_1258,N_788,N_121);
or U1259 (N_1259,N_506,N_356);
nand U1260 (N_1260,N_275,N_604);
nand U1261 (N_1261,N_559,N_359);
xnor U1262 (N_1262,N_878,N_337);
nand U1263 (N_1263,N_766,N_248);
nor U1264 (N_1264,N_691,N_353);
nor U1265 (N_1265,N_745,N_568);
and U1266 (N_1266,N_744,N_486);
and U1267 (N_1267,N_998,N_748);
and U1268 (N_1268,N_446,N_387);
nand U1269 (N_1269,N_931,N_282);
nand U1270 (N_1270,N_685,N_575);
nor U1271 (N_1271,N_593,N_268);
and U1272 (N_1272,N_391,N_531);
or U1273 (N_1273,N_499,N_31);
xor U1274 (N_1274,N_914,N_539);
or U1275 (N_1275,N_821,N_954);
nand U1276 (N_1276,N_378,N_733);
or U1277 (N_1277,N_763,N_699);
nor U1278 (N_1278,N_683,N_886);
nor U1279 (N_1279,N_437,N_238);
and U1280 (N_1280,N_852,N_381);
nor U1281 (N_1281,N_489,N_348);
and U1282 (N_1282,N_570,N_407);
xnor U1283 (N_1283,N_624,N_43);
or U1284 (N_1284,N_754,N_567);
nand U1285 (N_1285,N_838,N_591);
or U1286 (N_1286,N_302,N_866);
xnor U1287 (N_1287,N_267,N_228);
nor U1288 (N_1288,N_910,N_24);
or U1289 (N_1289,N_389,N_573);
xor U1290 (N_1290,N_321,N_106);
xnor U1291 (N_1291,N_718,N_832);
xnor U1292 (N_1292,N_765,N_849);
and U1293 (N_1293,N_579,N_630);
nand U1294 (N_1294,N_369,N_373);
and U1295 (N_1295,N_677,N_574);
or U1296 (N_1296,N_711,N_951);
xor U1297 (N_1297,N_66,N_165);
or U1298 (N_1298,N_279,N_111);
or U1299 (N_1299,N_867,N_629);
xnor U1300 (N_1300,N_341,N_908);
nor U1301 (N_1301,N_88,N_873);
xor U1302 (N_1302,N_883,N_828);
or U1303 (N_1303,N_278,N_968);
nor U1304 (N_1304,N_459,N_41);
xnor U1305 (N_1305,N_972,N_856);
nor U1306 (N_1306,N_144,N_773);
or U1307 (N_1307,N_661,N_853);
xor U1308 (N_1308,N_672,N_671);
nor U1309 (N_1309,N_252,N_625);
xnor U1310 (N_1310,N_492,N_882);
and U1311 (N_1311,N_885,N_338);
and U1312 (N_1312,N_956,N_597);
or U1313 (N_1313,N_318,N_870);
nand U1314 (N_1314,N_941,N_759);
and U1315 (N_1315,N_297,N_255);
nor U1316 (N_1316,N_425,N_827);
nor U1317 (N_1317,N_290,N_64);
and U1318 (N_1318,N_498,N_18);
xor U1319 (N_1319,N_316,N_644);
or U1320 (N_1320,N_984,N_350);
nand U1321 (N_1321,N_900,N_775);
and U1322 (N_1322,N_136,N_541);
xnor U1323 (N_1323,N_569,N_550);
or U1324 (N_1324,N_731,N_976);
nand U1325 (N_1325,N_462,N_611);
and U1326 (N_1326,N_456,N_368);
nand U1327 (N_1327,N_562,N_760);
or U1328 (N_1328,N_859,N_736);
nand U1329 (N_1329,N_332,N_798);
nor U1330 (N_1330,N_150,N_730);
xor U1331 (N_1331,N_922,N_995);
or U1332 (N_1332,N_535,N_490);
and U1333 (N_1333,N_971,N_12);
nor U1334 (N_1334,N_869,N_432);
xnor U1335 (N_1335,N_780,N_563);
and U1336 (N_1336,N_377,N_957);
or U1337 (N_1337,N_404,N_401);
xor U1338 (N_1338,N_29,N_179);
nand U1339 (N_1339,N_167,N_22);
nand U1340 (N_1340,N_113,N_482);
nand U1341 (N_1341,N_511,N_274);
or U1342 (N_1342,N_622,N_621);
nor U1343 (N_1343,N_208,N_518);
and U1344 (N_1344,N_175,N_218);
or U1345 (N_1345,N_710,N_138);
xor U1346 (N_1346,N_266,N_399);
and U1347 (N_1347,N_958,N_413);
nor U1348 (N_1348,N_139,N_892);
and U1349 (N_1349,N_836,N_902);
nand U1350 (N_1350,N_784,N_230);
and U1351 (N_1351,N_442,N_547);
xnor U1352 (N_1352,N_756,N_33);
nand U1353 (N_1353,N_762,N_120);
nor U1354 (N_1354,N_974,N_215);
xnor U1355 (N_1355,N_270,N_201);
and U1356 (N_1356,N_792,N_738);
and U1357 (N_1357,N_209,N_145);
xor U1358 (N_1358,N_657,N_476);
nand U1359 (N_1359,N_772,N_424);
or U1360 (N_1360,N_507,N_471);
nor U1361 (N_1361,N_62,N_183);
nor U1362 (N_1362,N_537,N_49);
nand U1363 (N_1363,N_612,N_955);
nor U1364 (N_1364,N_423,N_253);
and U1365 (N_1365,N_819,N_231);
xor U1366 (N_1366,N_355,N_627);
and U1367 (N_1367,N_307,N_98);
and U1368 (N_1368,N_623,N_367);
or U1369 (N_1369,N_757,N_204);
nor U1370 (N_1370,N_715,N_980);
xnor U1371 (N_1371,N_669,N_379);
nor U1372 (N_1372,N_816,N_953);
and U1373 (N_1373,N_913,N_713);
nand U1374 (N_1374,N_528,N_881);
nand U1375 (N_1375,N_645,N_961);
and U1376 (N_1376,N_753,N_831);
or U1377 (N_1377,N_239,N_326);
nand U1378 (N_1378,N_871,N_517);
xnor U1379 (N_1379,N_843,N_472);
or U1380 (N_1380,N_530,N_251);
nand U1381 (N_1381,N_271,N_94);
and U1382 (N_1382,N_696,N_992);
and U1383 (N_1383,N_879,N_652);
and U1384 (N_1384,N_244,N_135);
or U1385 (N_1385,N_219,N_104);
and U1386 (N_1386,N_159,N_641);
nand U1387 (N_1387,N_264,N_65);
nor U1388 (N_1388,N_27,N_223);
or U1389 (N_1389,N_545,N_449);
nor U1390 (N_1390,N_143,N_755);
or U1391 (N_1391,N_16,N_676);
nand U1392 (N_1392,N_258,N_7);
or U1393 (N_1393,N_544,N_71);
and U1394 (N_1394,N_229,N_687);
and U1395 (N_1395,N_214,N_576);
or U1396 (N_1396,N_750,N_429);
nand U1397 (N_1397,N_929,N_560);
and U1398 (N_1398,N_189,N_769);
nor U1399 (N_1399,N_74,N_679);
or U1400 (N_1400,N_458,N_981);
or U1401 (N_1401,N_403,N_899);
or U1402 (N_1402,N_944,N_440);
and U1403 (N_1403,N_521,N_509);
nor U1404 (N_1404,N_589,N_232);
or U1405 (N_1405,N_714,N_345);
and U1406 (N_1406,N_846,N_800);
nor U1407 (N_1407,N_289,N_751);
or U1408 (N_1408,N_335,N_996);
and U1409 (N_1409,N_30,N_187);
nand U1410 (N_1410,N_602,N_107);
xor U1411 (N_1411,N_102,N_952);
nor U1412 (N_1412,N_782,N_789);
nor U1413 (N_1413,N_554,N_352);
xor U1414 (N_1414,N_478,N_75);
nand U1415 (N_1415,N_86,N_690);
nand U1416 (N_1416,N_481,N_80);
nor U1417 (N_1417,N_123,N_133);
or U1418 (N_1418,N_116,N_833);
nor U1419 (N_1419,N_510,N_536);
nor U1420 (N_1420,N_994,N_740);
xor U1421 (N_1421,N_895,N_202);
nand U1422 (N_1422,N_247,N_964);
xnor U1423 (N_1423,N_421,N_888);
and U1424 (N_1424,N_39,N_415);
or U1425 (N_1425,N_764,N_932);
and U1426 (N_1426,N_985,N_692);
or U1427 (N_1427,N_592,N_140);
and U1428 (N_1428,N_673,N_108);
nand U1429 (N_1429,N_240,N_503);
and U1430 (N_1430,N_993,N_485);
and U1431 (N_1431,N_436,N_590);
xnor U1432 (N_1432,N_926,N_32);
xnor U1433 (N_1433,N_256,N_706);
nor U1434 (N_1434,N_181,N_496);
nor U1435 (N_1435,N_132,N_665);
nor U1436 (N_1436,N_126,N_213);
xor U1437 (N_1437,N_372,N_450);
or U1438 (N_1438,N_464,N_28);
or U1439 (N_1439,N_678,N_397);
or U1440 (N_1440,N_465,N_617);
or U1441 (N_1441,N_642,N_233);
nor U1442 (N_1442,N_0,N_408);
and U1443 (N_1443,N_583,N_224);
or U1444 (N_1444,N_203,N_257);
nand U1445 (N_1445,N_735,N_182);
or U1446 (N_1446,N_967,N_694);
nor U1447 (N_1447,N_844,N_868);
or U1448 (N_1448,N_5,N_67);
nand U1449 (N_1449,N_293,N_603);
nand U1450 (N_1450,N_196,N_250);
nand U1451 (N_1451,N_505,N_2);
nand U1452 (N_1452,N_398,N_841);
xnor U1453 (N_1453,N_211,N_194);
or U1454 (N_1454,N_829,N_986);
xnor U1455 (N_1455,N_124,N_566);
nand U1456 (N_1456,N_166,N_689);
nand U1457 (N_1457,N_585,N_325);
xnor U1458 (N_1458,N_502,N_808);
nand U1459 (N_1459,N_637,N_299);
or U1460 (N_1460,N_826,N_36);
nand U1461 (N_1461,N_936,N_522);
nor U1462 (N_1462,N_723,N_198);
or U1463 (N_1463,N_69,N_739);
and U1464 (N_1464,N_281,N_304);
and U1465 (N_1465,N_884,N_153);
or U1466 (N_1466,N_349,N_324);
xnor U1467 (N_1467,N_662,N_587);
xor U1468 (N_1468,N_358,N_172);
nor U1469 (N_1469,N_234,N_357);
and U1470 (N_1470,N_200,N_160);
nand U1471 (N_1471,N_707,N_128);
nor U1472 (N_1472,N_746,N_466);
or U1473 (N_1473,N_11,N_887);
and U1474 (N_1474,N_697,N_548);
and U1475 (N_1475,N_824,N_371);
xor U1476 (N_1476,N_158,N_475);
and U1477 (N_1477,N_965,N_206);
nand U1478 (N_1478,N_552,N_129);
or U1479 (N_1479,N_758,N_594);
or U1480 (N_1480,N_15,N_599);
nand U1481 (N_1481,N_638,N_435);
and U1482 (N_1482,N_312,N_495);
and U1483 (N_1483,N_292,N_480);
nand U1484 (N_1484,N_719,N_805);
xnor U1485 (N_1485,N_940,N_909);
nor U1486 (N_1486,N_333,N_553);
nand U1487 (N_1487,N_923,N_978);
or U1488 (N_1488,N_842,N_26);
nand U1489 (N_1489,N_48,N_727);
xnor U1490 (N_1490,N_384,N_514);
or U1491 (N_1491,N_220,N_606);
xnor U1492 (N_1492,N_286,N_347);
or U1493 (N_1493,N_263,N_975);
nor U1494 (N_1494,N_607,N_725);
or U1495 (N_1495,N_85,N_242);
or U1496 (N_1496,N_911,N_901);
xnor U1497 (N_1497,N_734,N_227);
or U1498 (N_1498,N_273,N_632);
and U1499 (N_1499,N_666,N_483);
or U1500 (N_1500,N_933,N_251);
nand U1501 (N_1501,N_244,N_360);
nand U1502 (N_1502,N_825,N_511);
or U1503 (N_1503,N_314,N_493);
nor U1504 (N_1504,N_465,N_932);
nor U1505 (N_1505,N_412,N_710);
nand U1506 (N_1506,N_327,N_606);
or U1507 (N_1507,N_339,N_74);
nand U1508 (N_1508,N_94,N_940);
nor U1509 (N_1509,N_80,N_400);
or U1510 (N_1510,N_705,N_786);
and U1511 (N_1511,N_263,N_467);
nand U1512 (N_1512,N_450,N_83);
nor U1513 (N_1513,N_57,N_280);
nor U1514 (N_1514,N_674,N_960);
nand U1515 (N_1515,N_831,N_376);
and U1516 (N_1516,N_91,N_356);
nor U1517 (N_1517,N_800,N_586);
nand U1518 (N_1518,N_249,N_459);
and U1519 (N_1519,N_223,N_58);
and U1520 (N_1520,N_27,N_91);
nand U1521 (N_1521,N_11,N_332);
xor U1522 (N_1522,N_220,N_247);
and U1523 (N_1523,N_678,N_104);
nand U1524 (N_1524,N_564,N_951);
nor U1525 (N_1525,N_955,N_441);
nand U1526 (N_1526,N_206,N_99);
or U1527 (N_1527,N_466,N_677);
xnor U1528 (N_1528,N_42,N_965);
and U1529 (N_1529,N_650,N_112);
nor U1530 (N_1530,N_795,N_783);
and U1531 (N_1531,N_607,N_731);
or U1532 (N_1532,N_594,N_354);
nor U1533 (N_1533,N_51,N_364);
nand U1534 (N_1534,N_341,N_420);
or U1535 (N_1535,N_706,N_961);
nor U1536 (N_1536,N_338,N_639);
nor U1537 (N_1537,N_488,N_298);
or U1538 (N_1538,N_157,N_671);
xnor U1539 (N_1539,N_483,N_971);
xor U1540 (N_1540,N_740,N_28);
nor U1541 (N_1541,N_384,N_670);
nand U1542 (N_1542,N_992,N_584);
nand U1543 (N_1543,N_850,N_522);
nor U1544 (N_1544,N_558,N_603);
xor U1545 (N_1545,N_999,N_112);
nor U1546 (N_1546,N_932,N_3);
nand U1547 (N_1547,N_819,N_693);
nand U1548 (N_1548,N_879,N_162);
xor U1549 (N_1549,N_318,N_575);
and U1550 (N_1550,N_624,N_847);
nor U1551 (N_1551,N_509,N_823);
nand U1552 (N_1552,N_604,N_241);
nand U1553 (N_1553,N_481,N_726);
xnor U1554 (N_1554,N_302,N_409);
nand U1555 (N_1555,N_142,N_250);
or U1556 (N_1556,N_477,N_978);
xnor U1557 (N_1557,N_864,N_93);
or U1558 (N_1558,N_571,N_467);
nand U1559 (N_1559,N_755,N_425);
nand U1560 (N_1560,N_432,N_529);
and U1561 (N_1561,N_869,N_583);
xor U1562 (N_1562,N_959,N_641);
nor U1563 (N_1563,N_143,N_280);
xor U1564 (N_1564,N_410,N_959);
xnor U1565 (N_1565,N_231,N_637);
nand U1566 (N_1566,N_824,N_906);
or U1567 (N_1567,N_533,N_921);
nand U1568 (N_1568,N_475,N_812);
nand U1569 (N_1569,N_226,N_692);
nand U1570 (N_1570,N_56,N_241);
xor U1571 (N_1571,N_529,N_596);
xor U1572 (N_1572,N_153,N_923);
nor U1573 (N_1573,N_549,N_249);
or U1574 (N_1574,N_153,N_779);
nand U1575 (N_1575,N_906,N_32);
nor U1576 (N_1576,N_886,N_951);
or U1577 (N_1577,N_255,N_553);
nand U1578 (N_1578,N_506,N_76);
and U1579 (N_1579,N_936,N_669);
nor U1580 (N_1580,N_262,N_199);
xnor U1581 (N_1581,N_28,N_250);
nand U1582 (N_1582,N_69,N_283);
nand U1583 (N_1583,N_306,N_480);
nor U1584 (N_1584,N_307,N_473);
xor U1585 (N_1585,N_746,N_295);
or U1586 (N_1586,N_971,N_81);
nor U1587 (N_1587,N_78,N_664);
and U1588 (N_1588,N_804,N_933);
and U1589 (N_1589,N_990,N_578);
nand U1590 (N_1590,N_298,N_717);
nand U1591 (N_1591,N_280,N_894);
or U1592 (N_1592,N_411,N_107);
or U1593 (N_1593,N_920,N_542);
nor U1594 (N_1594,N_726,N_872);
xnor U1595 (N_1595,N_120,N_279);
xnor U1596 (N_1596,N_874,N_610);
nor U1597 (N_1597,N_415,N_239);
and U1598 (N_1598,N_559,N_521);
xor U1599 (N_1599,N_433,N_879);
or U1600 (N_1600,N_788,N_857);
xnor U1601 (N_1601,N_593,N_45);
nand U1602 (N_1602,N_721,N_617);
nand U1603 (N_1603,N_276,N_600);
or U1604 (N_1604,N_636,N_226);
or U1605 (N_1605,N_279,N_688);
nand U1606 (N_1606,N_963,N_420);
and U1607 (N_1607,N_665,N_675);
xor U1608 (N_1608,N_952,N_30);
xnor U1609 (N_1609,N_359,N_378);
or U1610 (N_1610,N_873,N_618);
nor U1611 (N_1611,N_430,N_601);
and U1612 (N_1612,N_426,N_183);
nand U1613 (N_1613,N_23,N_886);
nor U1614 (N_1614,N_194,N_487);
and U1615 (N_1615,N_620,N_15);
and U1616 (N_1616,N_961,N_578);
or U1617 (N_1617,N_60,N_259);
nor U1618 (N_1618,N_754,N_61);
and U1619 (N_1619,N_552,N_701);
and U1620 (N_1620,N_600,N_312);
or U1621 (N_1621,N_56,N_406);
nand U1622 (N_1622,N_462,N_616);
and U1623 (N_1623,N_835,N_602);
or U1624 (N_1624,N_310,N_455);
nand U1625 (N_1625,N_866,N_677);
or U1626 (N_1626,N_620,N_107);
nor U1627 (N_1627,N_569,N_926);
xnor U1628 (N_1628,N_569,N_198);
or U1629 (N_1629,N_657,N_411);
or U1630 (N_1630,N_425,N_621);
nand U1631 (N_1631,N_268,N_876);
nor U1632 (N_1632,N_510,N_487);
or U1633 (N_1633,N_722,N_264);
xor U1634 (N_1634,N_653,N_100);
nand U1635 (N_1635,N_595,N_399);
nor U1636 (N_1636,N_369,N_228);
and U1637 (N_1637,N_580,N_498);
nor U1638 (N_1638,N_501,N_106);
and U1639 (N_1639,N_506,N_278);
and U1640 (N_1640,N_511,N_815);
nand U1641 (N_1641,N_521,N_819);
and U1642 (N_1642,N_76,N_377);
nand U1643 (N_1643,N_416,N_311);
or U1644 (N_1644,N_603,N_186);
or U1645 (N_1645,N_482,N_831);
and U1646 (N_1646,N_357,N_691);
nand U1647 (N_1647,N_437,N_313);
xnor U1648 (N_1648,N_504,N_856);
or U1649 (N_1649,N_469,N_853);
or U1650 (N_1650,N_225,N_903);
xnor U1651 (N_1651,N_735,N_653);
and U1652 (N_1652,N_497,N_263);
and U1653 (N_1653,N_100,N_13);
or U1654 (N_1654,N_977,N_571);
or U1655 (N_1655,N_89,N_767);
and U1656 (N_1656,N_5,N_160);
nor U1657 (N_1657,N_407,N_266);
nor U1658 (N_1658,N_858,N_695);
nor U1659 (N_1659,N_565,N_485);
or U1660 (N_1660,N_672,N_799);
xnor U1661 (N_1661,N_705,N_366);
nand U1662 (N_1662,N_927,N_842);
nor U1663 (N_1663,N_633,N_577);
nor U1664 (N_1664,N_33,N_280);
or U1665 (N_1665,N_908,N_124);
nor U1666 (N_1666,N_624,N_877);
xor U1667 (N_1667,N_272,N_648);
nand U1668 (N_1668,N_240,N_753);
nor U1669 (N_1669,N_110,N_363);
or U1670 (N_1670,N_644,N_786);
xnor U1671 (N_1671,N_911,N_840);
nand U1672 (N_1672,N_885,N_153);
and U1673 (N_1673,N_279,N_686);
xnor U1674 (N_1674,N_129,N_733);
and U1675 (N_1675,N_101,N_103);
nand U1676 (N_1676,N_514,N_492);
and U1677 (N_1677,N_135,N_509);
nand U1678 (N_1678,N_746,N_456);
xnor U1679 (N_1679,N_893,N_408);
xnor U1680 (N_1680,N_131,N_358);
xnor U1681 (N_1681,N_801,N_605);
xnor U1682 (N_1682,N_219,N_291);
nand U1683 (N_1683,N_241,N_558);
nand U1684 (N_1684,N_219,N_870);
xnor U1685 (N_1685,N_291,N_944);
nor U1686 (N_1686,N_881,N_827);
or U1687 (N_1687,N_836,N_172);
nand U1688 (N_1688,N_942,N_388);
or U1689 (N_1689,N_440,N_460);
nor U1690 (N_1690,N_691,N_91);
xnor U1691 (N_1691,N_959,N_966);
or U1692 (N_1692,N_227,N_154);
or U1693 (N_1693,N_306,N_501);
xnor U1694 (N_1694,N_861,N_274);
xor U1695 (N_1695,N_762,N_340);
or U1696 (N_1696,N_761,N_983);
xnor U1697 (N_1697,N_222,N_410);
nand U1698 (N_1698,N_256,N_903);
and U1699 (N_1699,N_414,N_265);
or U1700 (N_1700,N_84,N_282);
or U1701 (N_1701,N_127,N_309);
nor U1702 (N_1702,N_291,N_153);
nor U1703 (N_1703,N_727,N_450);
and U1704 (N_1704,N_729,N_337);
and U1705 (N_1705,N_74,N_941);
nor U1706 (N_1706,N_531,N_595);
xor U1707 (N_1707,N_999,N_511);
nand U1708 (N_1708,N_126,N_184);
nand U1709 (N_1709,N_638,N_883);
nand U1710 (N_1710,N_538,N_17);
and U1711 (N_1711,N_538,N_152);
or U1712 (N_1712,N_405,N_710);
nand U1713 (N_1713,N_457,N_963);
nor U1714 (N_1714,N_366,N_358);
nor U1715 (N_1715,N_521,N_575);
nor U1716 (N_1716,N_831,N_679);
or U1717 (N_1717,N_218,N_731);
and U1718 (N_1718,N_142,N_675);
nor U1719 (N_1719,N_922,N_678);
and U1720 (N_1720,N_796,N_230);
nor U1721 (N_1721,N_79,N_857);
nor U1722 (N_1722,N_129,N_948);
and U1723 (N_1723,N_199,N_569);
nand U1724 (N_1724,N_161,N_284);
and U1725 (N_1725,N_331,N_647);
and U1726 (N_1726,N_124,N_317);
nor U1727 (N_1727,N_696,N_59);
or U1728 (N_1728,N_234,N_979);
and U1729 (N_1729,N_483,N_56);
nand U1730 (N_1730,N_78,N_475);
nand U1731 (N_1731,N_407,N_561);
nor U1732 (N_1732,N_719,N_369);
and U1733 (N_1733,N_25,N_984);
and U1734 (N_1734,N_330,N_31);
and U1735 (N_1735,N_497,N_381);
nand U1736 (N_1736,N_391,N_183);
or U1737 (N_1737,N_556,N_978);
nor U1738 (N_1738,N_145,N_884);
or U1739 (N_1739,N_422,N_637);
nor U1740 (N_1740,N_721,N_333);
xor U1741 (N_1741,N_460,N_768);
or U1742 (N_1742,N_86,N_493);
nand U1743 (N_1743,N_729,N_203);
nand U1744 (N_1744,N_30,N_90);
or U1745 (N_1745,N_675,N_611);
and U1746 (N_1746,N_328,N_402);
or U1747 (N_1747,N_160,N_266);
xor U1748 (N_1748,N_523,N_455);
xor U1749 (N_1749,N_914,N_392);
xor U1750 (N_1750,N_658,N_74);
or U1751 (N_1751,N_51,N_524);
and U1752 (N_1752,N_133,N_19);
nor U1753 (N_1753,N_87,N_932);
or U1754 (N_1754,N_908,N_491);
and U1755 (N_1755,N_804,N_394);
nand U1756 (N_1756,N_779,N_86);
and U1757 (N_1757,N_167,N_807);
nor U1758 (N_1758,N_990,N_404);
and U1759 (N_1759,N_110,N_595);
xnor U1760 (N_1760,N_192,N_611);
nand U1761 (N_1761,N_533,N_456);
nand U1762 (N_1762,N_247,N_824);
nor U1763 (N_1763,N_981,N_910);
or U1764 (N_1764,N_655,N_957);
and U1765 (N_1765,N_729,N_597);
nand U1766 (N_1766,N_934,N_20);
xor U1767 (N_1767,N_23,N_403);
nand U1768 (N_1768,N_412,N_983);
or U1769 (N_1769,N_931,N_239);
xor U1770 (N_1770,N_930,N_600);
nand U1771 (N_1771,N_743,N_911);
xnor U1772 (N_1772,N_100,N_528);
nand U1773 (N_1773,N_35,N_635);
xor U1774 (N_1774,N_335,N_255);
and U1775 (N_1775,N_611,N_912);
or U1776 (N_1776,N_808,N_568);
xnor U1777 (N_1777,N_892,N_697);
nand U1778 (N_1778,N_980,N_939);
or U1779 (N_1779,N_394,N_101);
nand U1780 (N_1780,N_2,N_970);
xor U1781 (N_1781,N_766,N_238);
nand U1782 (N_1782,N_358,N_164);
nor U1783 (N_1783,N_181,N_245);
nor U1784 (N_1784,N_76,N_691);
nand U1785 (N_1785,N_535,N_45);
nand U1786 (N_1786,N_839,N_690);
nor U1787 (N_1787,N_499,N_869);
or U1788 (N_1788,N_585,N_878);
xor U1789 (N_1789,N_635,N_679);
nand U1790 (N_1790,N_147,N_493);
and U1791 (N_1791,N_398,N_847);
or U1792 (N_1792,N_550,N_763);
and U1793 (N_1793,N_299,N_157);
or U1794 (N_1794,N_514,N_336);
and U1795 (N_1795,N_254,N_628);
nand U1796 (N_1796,N_983,N_154);
nor U1797 (N_1797,N_126,N_262);
or U1798 (N_1798,N_215,N_444);
xnor U1799 (N_1799,N_785,N_132);
and U1800 (N_1800,N_751,N_293);
nor U1801 (N_1801,N_105,N_179);
nand U1802 (N_1802,N_590,N_400);
nor U1803 (N_1803,N_739,N_96);
nand U1804 (N_1804,N_67,N_645);
nand U1805 (N_1805,N_315,N_25);
and U1806 (N_1806,N_494,N_260);
nand U1807 (N_1807,N_637,N_647);
nand U1808 (N_1808,N_841,N_139);
nand U1809 (N_1809,N_121,N_503);
nor U1810 (N_1810,N_599,N_816);
nand U1811 (N_1811,N_971,N_440);
or U1812 (N_1812,N_798,N_867);
xnor U1813 (N_1813,N_457,N_184);
nand U1814 (N_1814,N_148,N_655);
nand U1815 (N_1815,N_899,N_238);
or U1816 (N_1816,N_782,N_557);
nor U1817 (N_1817,N_786,N_815);
nor U1818 (N_1818,N_647,N_852);
or U1819 (N_1819,N_187,N_572);
xor U1820 (N_1820,N_468,N_959);
or U1821 (N_1821,N_574,N_714);
nor U1822 (N_1822,N_240,N_862);
nor U1823 (N_1823,N_706,N_113);
xor U1824 (N_1824,N_267,N_405);
nor U1825 (N_1825,N_299,N_948);
or U1826 (N_1826,N_344,N_337);
nor U1827 (N_1827,N_802,N_782);
nor U1828 (N_1828,N_574,N_605);
and U1829 (N_1829,N_673,N_373);
nand U1830 (N_1830,N_591,N_623);
or U1831 (N_1831,N_525,N_626);
nor U1832 (N_1832,N_371,N_402);
xor U1833 (N_1833,N_373,N_322);
nor U1834 (N_1834,N_879,N_909);
xnor U1835 (N_1835,N_160,N_436);
nand U1836 (N_1836,N_119,N_685);
xor U1837 (N_1837,N_23,N_913);
or U1838 (N_1838,N_951,N_183);
xnor U1839 (N_1839,N_103,N_720);
or U1840 (N_1840,N_47,N_203);
nor U1841 (N_1841,N_211,N_896);
nor U1842 (N_1842,N_845,N_653);
and U1843 (N_1843,N_321,N_13);
and U1844 (N_1844,N_352,N_385);
nor U1845 (N_1845,N_561,N_592);
nor U1846 (N_1846,N_256,N_749);
or U1847 (N_1847,N_340,N_604);
nor U1848 (N_1848,N_296,N_973);
and U1849 (N_1849,N_160,N_879);
nor U1850 (N_1850,N_586,N_447);
nand U1851 (N_1851,N_972,N_707);
or U1852 (N_1852,N_706,N_332);
nand U1853 (N_1853,N_265,N_439);
xor U1854 (N_1854,N_191,N_52);
and U1855 (N_1855,N_400,N_303);
nor U1856 (N_1856,N_817,N_895);
nor U1857 (N_1857,N_769,N_695);
nand U1858 (N_1858,N_506,N_533);
nor U1859 (N_1859,N_111,N_235);
xor U1860 (N_1860,N_839,N_854);
xor U1861 (N_1861,N_726,N_755);
nor U1862 (N_1862,N_435,N_741);
nand U1863 (N_1863,N_539,N_853);
nand U1864 (N_1864,N_495,N_492);
nand U1865 (N_1865,N_552,N_108);
nor U1866 (N_1866,N_159,N_545);
nand U1867 (N_1867,N_942,N_4);
nand U1868 (N_1868,N_571,N_193);
and U1869 (N_1869,N_693,N_250);
xor U1870 (N_1870,N_530,N_243);
and U1871 (N_1871,N_44,N_459);
and U1872 (N_1872,N_419,N_352);
nor U1873 (N_1873,N_931,N_789);
and U1874 (N_1874,N_138,N_966);
nand U1875 (N_1875,N_423,N_556);
nand U1876 (N_1876,N_927,N_811);
nand U1877 (N_1877,N_746,N_780);
nand U1878 (N_1878,N_869,N_867);
xor U1879 (N_1879,N_515,N_360);
and U1880 (N_1880,N_913,N_31);
nor U1881 (N_1881,N_71,N_54);
or U1882 (N_1882,N_201,N_764);
xnor U1883 (N_1883,N_629,N_603);
and U1884 (N_1884,N_67,N_618);
or U1885 (N_1885,N_487,N_449);
xor U1886 (N_1886,N_253,N_84);
nand U1887 (N_1887,N_679,N_260);
xor U1888 (N_1888,N_646,N_344);
and U1889 (N_1889,N_269,N_613);
and U1890 (N_1890,N_341,N_738);
xnor U1891 (N_1891,N_34,N_937);
and U1892 (N_1892,N_490,N_688);
and U1893 (N_1893,N_357,N_427);
nor U1894 (N_1894,N_7,N_132);
nand U1895 (N_1895,N_716,N_40);
nor U1896 (N_1896,N_419,N_485);
nor U1897 (N_1897,N_37,N_139);
nor U1898 (N_1898,N_792,N_902);
xor U1899 (N_1899,N_741,N_918);
or U1900 (N_1900,N_796,N_270);
xnor U1901 (N_1901,N_343,N_201);
xor U1902 (N_1902,N_433,N_962);
nor U1903 (N_1903,N_623,N_409);
nand U1904 (N_1904,N_129,N_54);
nand U1905 (N_1905,N_701,N_208);
or U1906 (N_1906,N_574,N_812);
nand U1907 (N_1907,N_524,N_655);
and U1908 (N_1908,N_715,N_788);
nor U1909 (N_1909,N_373,N_623);
or U1910 (N_1910,N_378,N_780);
nand U1911 (N_1911,N_74,N_483);
nor U1912 (N_1912,N_432,N_821);
xnor U1913 (N_1913,N_796,N_875);
or U1914 (N_1914,N_162,N_245);
nor U1915 (N_1915,N_811,N_978);
nand U1916 (N_1916,N_507,N_730);
and U1917 (N_1917,N_715,N_124);
nor U1918 (N_1918,N_354,N_307);
nor U1919 (N_1919,N_177,N_113);
nand U1920 (N_1920,N_752,N_724);
and U1921 (N_1921,N_255,N_68);
and U1922 (N_1922,N_211,N_599);
nor U1923 (N_1923,N_191,N_38);
nand U1924 (N_1924,N_184,N_202);
xor U1925 (N_1925,N_125,N_324);
nand U1926 (N_1926,N_953,N_597);
and U1927 (N_1927,N_39,N_613);
nor U1928 (N_1928,N_910,N_134);
nand U1929 (N_1929,N_231,N_461);
nand U1930 (N_1930,N_184,N_381);
and U1931 (N_1931,N_79,N_220);
or U1932 (N_1932,N_643,N_901);
xor U1933 (N_1933,N_418,N_217);
xor U1934 (N_1934,N_1,N_433);
xor U1935 (N_1935,N_326,N_547);
nor U1936 (N_1936,N_849,N_863);
and U1937 (N_1937,N_829,N_285);
or U1938 (N_1938,N_616,N_86);
nand U1939 (N_1939,N_80,N_292);
xnor U1940 (N_1940,N_29,N_499);
and U1941 (N_1941,N_383,N_500);
or U1942 (N_1942,N_858,N_893);
nor U1943 (N_1943,N_973,N_69);
xor U1944 (N_1944,N_316,N_641);
and U1945 (N_1945,N_148,N_661);
or U1946 (N_1946,N_2,N_812);
and U1947 (N_1947,N_738,N_291);
xnor U1948 (N_1948,N_840,N_522);
and U1949 (N_1949,N_834,N_814);
and U1950 (N_1950,N_189,N_843);
or U1951 (N_1951,N_41,N_396);
nand U1952 (N_1952,N_15,N_240);
nor U1953 (N_1953,N_54,N_695);
and U1954 (N_1954,N_418,N_598);
xor U1955 (N_1955,N_161,N_221);
and U1956 (N_1956,N_691,N_93);
nand U1957 (N_1957,N_12,N_330);
and U1958 (N_1958,N_896,N_7);
and U1959 (N_1959,N_16,N_702);
and U1960 (N_1960,N_822,N_249);
or U1961 (N_1961,N_467,N_670);
nand U1962 (N_1962,N_257,N_273);
or U1963 (N_1963,N_218,N_600);
nor U1964 (N_1964,N_470,N_597);
nand U1965 (N_1965,N_854,N_950);
nand U1966 (N_1966,N_75,N_835);
or U1967 (N_1967,N_180,N_46);
and U1968 (N_1968,N_118,N_599);
xor U1969 (N_1969,N_438,N_75);
nand U1970 (N_1970,N_16,N_913);
xnor U1971 (N_1971,N_116,N_259);
xnor U1972 (N_1972,N_383,N_321);
or U1973 (N_1973,N_92,N_819);
nor U1974 (N_1974,N_387,N_645);
and U1975 (N_1975,N_965,N_223);
nor U1976 (N_1976,N_766,N_521);
xnor U1977 (N_1977,N_392,N_133);
nor U1978 (N_1978,N_714,N_857);
nand U1979 (N_1979,N_393,N_362);
nand U1980 (N_1980,N_427,N_522);
xnor U1981 (N_1981,N_629,N_320);
or U1982 (N_1982,N_821,N_276);
xnor U1983 (N_1983,N_482,N_478);
nor U1984 (N_1984,N_686,N_917);
nor U1985 (N_1985,N_388,N_12);
nor U1986 (N_1986,N_542,N_333);
nand U1987 (N_1987,N_299,N_459);
nor U1988 (N_1988,N_217,N_241);
nor U1989 (N_1989,N_191,N_258);
and U1990 (N_1990,N_742,N_888);
nand U1991 (N_1991,N_515,N_328);
or U1992 (N_1992,N_33,N_739);
xor U1993 (N_1993,N_779,N_404);
nand U1994 (N_1994,N_915,N_565);
nand U1995 (N_1995,N_568,N_207);
nor U1996 (N_1996,N_5,N_286);
xor U1997 (N_1997,N_715,N_817);
nor U1998 (N_1998,N_931,N_174);
and U1999 (N_1999,N_255,N_950);
nand U2000 (N_2000,N_1354,N_1046);
and U2001 (N_2001,N_1775,N_1386);
nand U2002 (N_2002,N_1207,N_1611);
or U2003 (N_2003,N_1944,N_1906);
nand U2004 (N_2004,N_1209,N_1844);
and U2005 (N_2005,N_1073,N_1296);
and U2006 (N_2006,N_1187,N_1005);
xor U2007 (N_2007,N_1016,N_1934);
nand U2008 (N_2008,N_1822,N_1013);
or U2009 (N_2009,N_1765,N_1315);
or U2010 (N_2010,N_1426,N_1247);
nand U2011 (N_2011,N_1782,N_1672);
xnor U2012 (N_2012,N_1523,N_1175);
nand U2013 (N_2013,N_1729,N_1221);
and U2014 (N_2014,N_1358,N_1986);
xnor U2015 (N_2015,N_1253,N_1940);
and U2016 (N_2016,N_1798,N_1548);
and U2017 (N_2017,N_1955,N_1120);
or U2018 (N_2018,N_1361,N_1741);
nand U2019 (N_2019,N_1463,N_1905);
nor U2020 (N_2020,N_1242,N_1731);
xnor U2021 (N_2021,N_1717,N_1928);
xor U2022 (N_2022,N_1500,N_1884);
nor U2023 (N_2023,N_1943,N_1017);
xor U2024 (N_2024,N_1843,N_1606);
nor U2025 (N_2025,N_1563,N_1237);
xor U2026 (N_2026,N_1302,N_1541);
and U2027 (N_2027,N_1544,N_1430);
and U2028 (N_2028,N_1234,N_1058);
or U2029 (N_2029,N_1012,N_1599);
or U2030 (N_2030,N_1888,N_1461);
and U2031 (N_2031,N_1300,N_1041);
nor U2032 (N_2032,N_1492,N_1057);
nand U2033 (N_2033,N_1042,N_1538);
or U2034 (N_2034,N_1923,N_1200);
xor U2035 (N_2035,N_1483,N_1681);
xor U2036 (N_2036,N_1124,N_1524);
nor U2037 (N_2037,N_1521,N_1048);
nand U2038 (N_2038,N_1738,N_1661);
nor U2039 (N_2039,N_1146,N_1640);
or U2040 (N_2040,N_1091,N_1632);
or U2041 (N_2041,N_1010,N_1197);
or U2042 (N_2042,N_1753,N_1388);
xnor U2043 (N_2043,N_1812,N_1589);
and U2044 (N_2044,N_1994,N_1869);
or U2045 (N_2045,N_1066,N_1825);
or U2046 (N_2046,N_1759,N_1078);
and U2047 (N_2047,N_1920,N_1101);
nand U2048 (N_2048,N_1852,N_1348);
and U2049 (N_2049,N_1049,N_1513);
and U2050 (N_2050,N_1192,N_1368);
xor U2051 (N_2051,N_1227,N_1180);
nor U2052 (N_2052,N_1097,N_1927);
nand U2053 (N_2053,N_1686,N_1113);
xnor U2054 (N_2054,N_1896,N_1429);
nor U2055 (N_2055,N_1325,N_1576);
nor U2056 (N_2056,N_1445,N_1470);
nand U2057 (N_2057,N_1229,N_1918);
and U2058 (N_2058,N_1722,N_1022);
nor U2059 (N_2059,N_1841,N_1208);
and U2060 (N_2060,N_1441,N_1107);
or U2061 (N_2061,N_1614,N_1402);
nand U2062 (N_2062,N_1342,N_1625);
nor U2063 (N_2063,N_1117,N_1960);
or U2064 (N_2064,N_1181,N_1322);
xnor U2065 (N_2065,N_1901,N_1559);
and U2066 (N_2066,N_1875,N_1929);
nand U2067 (N_2067,N_1275,N_1536);
nor U2068 (N_2068,N_1155,N_1919);
nand U2069 (N_2069,N_1420,N_1836);
xnor U2070 (N_2070,N_1450,N_1027);
nor U2071 (N_2071,N_1469,N_1511);
xor U2072 (N_2072,N_1479,N_1439);
nand U2073 (N_2073,N_1055,N_1396);
nor U2074 (N_2074,N_1863,N_1937);
and U2075 (N_2075,N_1405,N_1615);
nor U2076 (N_2076,N_1635,N_1881);
or U2077 (N_2077,N_1594,N_1842);
or U2078 (N_2078,N_1164,N_1975);
xnor U2079 (N_2079,N_1032,N_1566);
xor U2080 (N_2080,N_1643,N_1845);
and U2081 (N_2081,N_1561,N_1867);
and U2082 (N_2082,N_1831,N_1504);
xnor U2083 (N_2083,N_1848,N_1334);
nand U2084 (N_2084,N_1721,N_1428);
nor U2085 (N_2085,N_1535,N_1703);
xnor U2086 (N_2086,N_1318,N_1104);
or U2087 (N_2087,N_1416,N_1704);
nand U2088 (N_2088,N_1166,N_1959);
or U2089 (N_2089,N_1945,N_1894);
xor U2090 (N_2090,N_1382,N_1593);
nor U2091 (N_2091,N_1758,N_1417);
nand U2092 (N_2092,N_1760,N_1198);
or U2093 (N_2093,N_1186,N_1067);
xnor U2094 (N_2094,N_1433,N_1040);
or U2095 (N_2095,N_1321,N_1021);
and U2096 (N_2096,N_1886,N_1231);
xnor U2097 (N_2097,N_1774,N_1803);
nor U2098 (N_2098,N_1303,N_1965);
and U2099 (N_2099,N_1832,N_1462);
xor U2100 (N_2100,N_1385,N_1381);
and U2101 (N_2101,N_1512,N_1281);
and U2102 (N_2102,N_1217,N_1719);
nor U2103 (N_2103,N_1079,N_1408);
xor U2104 (N_2104,N_1478,N_1711);
nand U2105 (N_2105,N_1948,N_1103);
or U2106 (N_2106,N_1284,N_1367);
xnor U2107 (N_2107,N_1194,N_1584);
or U2108 (N_2108,N_1476,N_1618);
nand U2109 (N_2109,N_1880,N_1043);
nand U2110 (N_2110,N_1678,N_1609);
and U2111 (N_2111,N_1258,N_1581);
and U2112 (N_2112,N_1437,N_1074);
or U2113 (N_2113,N_1977,N_1460);
xnor U2114 (N_2114,N_1018,N_1213);
nor U2115 (N_2115,N_1784,N_1464);
xor U2116 (N_2116,N_1723,N_1634);
nand U2117 (N_2117,N_1442,N_1510);
and U2118 (N_2118,N_1333,N_1817);
xnor U2119 (N_2119,N_1708,N_1082);
nor U2120 (N_2120,N_1826,N_1954);
nor U2121 (N_2121,N_1345,N_1885);
xnor U2122 (N_2122,N_1392,N_1298);
nor U2123 (N_2123,N_1569,N_1664);
or U2124 (N_2124,N_1801,N_1114);
xor U2125 (N_2125,N_1056,N_1412);
xnor U2126 (N_2126,N_1639,N_1020);
or U2127 (N_2127,N_1421,N_1667);
nand U2128 (N_2128,N_1932,N_1550);
or U2129 (N_2129,N_1794,N_1659);
xor U2130 (N_2130,N_1178,N_1185);
nor U2131 (N_2131,N_1063,N_1150);
nand U2132 (N_2132,N_1356,N_1481);
and U2133 (N_2133,N_1369,N_1821);
nand U2134 (N_2134,N_1655,N_1520);
or U2135 (N_2135,N_1309,N_1813);
and U2136 (N_2136,N_1262,N_1330);
nand U2137 (N_2137,N_1182,N_1740);
and U2138 (N_2138,N_1828,N_1980);
or U2139 (N_2139,N_1274,N_1856);
nand U2140 (N_2140,N_1733,N_1952);
and U2141 (N_2141,N_1264,N_1866);
and U2142 (N_2142,N_1053,N_1241);
and U2143 (N_2143,N_1037,N_1574);
or U2144 (N_2144,N_1993,N_1077);
and U2145 (N_2145,N_1080,N_1174);
and U2146 (N_2146,N_1793,N_1202);
xor U2147 (N_2147,N_1691,N_1316);
or U2148 (N_2148,N_1707,N_1489);
nand U2149 (N_2149,N_1438,N_1709);
and U2150 (N_2150,N_1344,N_1914);
nor U2151 (N_2151,N_1145,N_1604);
nand U2152 (N_2152,N_1839,N_1362);
nor U2153 (N_2153,N_1061,N_1773);
xor U2154 (N_2154,N_1143,N_1751);
nand U2155 (N_2155,N_1534,N_1697);
and U2156 (N_2156,N_1950,N_1799);
xor U2157 (N_2157,N_1583,N_1849);
and U2158 (N_2158,N_1169,N_1311);
nand U2159 (N_2159,N_1682,N_1338);
or U2160 (N_2160,N_1240,N_1642);
xor U2161 (N_2161,N_1163,N_1516);
and U2162 (N_2162,N_1997,N_1151);
nor U2163 (N_2163,N_1230,N_1468);
or U2164 (N_2164,N_1808,N_1910);
and U2165 (N_2165,N_1289,N_1352);
nand U2166 (N_2166,N_1728,N_1419);
or U2167 (N_2167,N_1525,N_1501);
nand U2168 (N_2168,N_1855,N_1715);
nand U2169 (N_2169,N_1677,N_1554);
nand U2170 (N_2170,N_1130,N_1327);
and U2171 (N_2171,N_1689,N_1968);
nand U2172 (N_2172,N_1071,N_1065);
nor U2173 (N_2173,N_1670,N_1467);
and U2174 (N_2174,N_1788,N_1602);
nand U2175 (N_2175,N_1936,N_1783);
or U2176 (N_2176,N_1573,N_1393);
xor U2177 (N_2177,N_1269,N_1792);
xnor U2178 (N_2178,N_1093,N_1015);
and U2179 (N_2179,N_1714,N_1118);
nor U2180 (N_2180,N_1373,N_1949);
nand U2181 (N_2181,N_1546,N_1451);
nand U2182 (N_2182,N_1394,N_1626);
xnor U2183 (N_2183,N_1448,N_1777);
nand U2184 (N_2184,N_1768,N_1487);
xor U2185 (N_2185,N_1283,N_1038);
nor U2186 (N_2186,N_1987,N_1854);
or U2187 (N_2187,N_1624,N_1789);
xor U2188 (N_2188,N_1216,N_1658);
nor U2189 (N_2189,N_1045,N_1355);
or U2190 (N_2190,N_1688,N_1224);
xor U2191 (N_2191,N_1853,N_1176);
xnor U2192 (N_2192,N_1374,N_1805);
or U2193 (N_2193,N_1830,N_1075);
xnor U2194 (N_2194,N_1877,N_1098);
and U2195 (N_2195,N_1299,N_1449);
or U2196 (N_2196,N_1956,N_1070);
and U2197 (N_2197,N_1736,N_1526);
nand U2198 (N_2198,N_1482,N_1495);
xor U2199 (N_2199,N_1455,N_1909);
nand U2200 (N_2200,N_1440,N_1263);
nand U2201 (N_2201,N_1564,N_1819);
nor U2202 (N_2202,N_1656,N_1543);
nor U2203 (N_2203,N_1484,N_1857);
nand U2204 (N_2204,N_1490,N_1111);
nand U2205 (N_2205,N_1779,N_1982);
nand U2206 (N_2206,N_1054,N_1557);
xor U2207 (N_2207,N_1239,N_1232);
xnor U2208 (N_2208,N_1245,N_1129);
and U2209 (N_2209,N_1925,N_1149);
nor U2210 (N_2210,N_1999,N_1941);
nand U2211 (N_2211,N_1148,N_1834);
nand U2212 (N_2212,N_1305,N_1273);
or U2213 (N_2213,N_1648,N_1962);
or U2214 (N_2214,N_1776,N_1366);
xnor U2215 (N_2215,N_1364,N_1961);
nor U2216 (N_2216,N_1924,N_1814);
xor U2217 (N_2217,N_1218,N_1638);
or U2218 (N_2218,N_1457,N_1858);
and U2219 (N_2219,N_1882,N_1008);
or U2220 (N_2220,N_1860,N_1319);
nor U2221 (N_2221,N_1903,N_1404);
nand U2222 (N_2222,N_1147,N_1797);
nor U2223 (N_2223,N_1400,N_1372);
nand U2224 (N_2224,N_1921,N_1807);
or U2225 (N_2225,N_1996,N_1096);
and U2226 (N_2226,N_1219,N_1555);
or U2227 (N_2227,N_1293,N_1974);
nand U2228 (N_2228,N_1754,N_1418);
and U2229 (N_2229,N_1683,N_1039);
nor U2230 (N_2230,N_1387,N_1621);
nor U2231 (N_2231,N_1970,N_1837);
nand U2232 (N_2232,N_1761,N_1818);
and U2233 (N_2233,N_1631,N_1846);
nor U2234 (N_2234,N_1767,N_1654);
or U2235 (N_2235,N_1126,N_1502);
and U2236 (N_2236,N_1726,N_1081);
or U2237 (N_2237,N_1616,N_1095);
xor U2238 (N_2238,N_1899,N_1350);
nor U2239 (N_2239,N_1306,N_1553);
nor U2240 (N_2240,N_1290,N_1623);
nand U2241 (N_2241,N_1183,N_1904);
nand U2242 (N_2242,N_1585,N_1529);
xor U2243 (N_2243,N_1637,N_1424);
or U2244 (N_2244,N_1244,N_1674);
xor U2245 (N_2245,N_1001,N_1475);
xnor U2246 (N_2246,N_1864,N_1131);
nor U2247 (N_2247,N_1106,N_1873);
or U2248 (N_2248,N_1435,N_1279);
and U2249 (N_2249,N_1514,N_1699);
and U2250 (N_2250,N_1379,N_1427);
and U2251 (N_2251,N_1991,N_1389);
xor U2252 (N_2252,N_1320,N_1436);
nand U2253 (N_2253,N_1608,N_1735);
or U2254 (N_2254,N_1749,N_1161);
or U2255 (N_2255,N_1995,N_1907);
nor U2256 (N_2256,N_1170,N_1014);
xor U2257 (N_2257,N_1233,N_1254);
or U2258 (N_2258,N_1718,N_1085);
nand U2259 (N_2259,N_1981,N_1339);
nand U2260 (N_2260,N_1630,N_1720);
nor U2261 (N_2261,N_1734,N_1809);
or U2262 (N_2262,N_1669,N_1212);
nor U2263 (N_2263,N_1157,N_1598);
or U2264 (N_2264,N_1990,N_1930);
xor U2265 (N_2265,N_1102,N_1190);
xor U2266 (N_2266,N_1786,N_1908);
xor U2267 (N_2267,N_1862,N_1052);
or U2268 (N_2268,N_1973,N_1824);
xnor U2269 (N_2269,N_1280,N_1804);
nor U2270 (N_2270,N_1033,N_1547);
or U2271 (N_2271,N_1665,N_1755);
nand U2272 (N_2272,N_1727,N_1532);
or U2273 (N_2273,N_1653,N_1222);
nand U2274 (N_2274,N_1375,N_1971);
xnor U2275 (N_2275,N_1282,N_1456);
or U2276 (N_2276,N_1023,N_1189);
nor U2277 (N_2277,N_1570,N_1984);
nor U2278 (N_2278,N_1823,N_1485);
and U2279 (N_2279,N_1795,N_1173);
and U2280 (N_2280,N_1086,N_1215);
and U2281 (N_2281,N_1307,N_1029);
xnor U2282 (N_2282,N_1006,N_1693);
and U2283 (N_2283,N_1992,N_1480);
and U2284 (N_2284,N_1756,N_1335);
or U2285 (N_2285,N_1211,N_1380);
xor U2286 (N_2286,N_1769,N_1138);
xnor U2287 (N_2287,N_1730,N_1351);
nand U2288 (N_2288,N_1158,N_1474);
or U2289 (N_2289,N_1494,N_1540);
and U2290 (N_2290,N_1410,N_1477);
nor U2291 (N_2291,N_1287,N_1542);
xor U2292 (N_2292,N_1411,N_1633);
nand U2293 (N_2293,N_1515,N_1601);
xnor U2294 (N_2294,N_1278,N_1261);
or U2295 (N_2295,N_1499,N_1815);
nand U2296 (N_2296,N_1787,N_1887);
nand U2297 (N_2297,N_1266,N_1458);
and U2298 (N_2298,N_1235,N_1329);
nand U2299 (N_2299,N_1099,N_1324);
or U2300 (N_2300,N_1331,N_1859);
nand U2301 (N_2301,N_1226,N_1911);
or U2302 (N_2302,N_1011,N_1926);
xnor U2303 (N_2303,N_1549,N_1090);
and U2304 (N_2304,N_1705,N_1087);
nor U2305 (N_2305,N_1252,N_1644);
and U2306 (N_2306,N_1946,N_1084);
nand U2307 (N_2307,N_1024,N_1916);
nand U2308 (N_2308,N_1127,N_1370);
or U2309 (N_2309,N_1204,N_1142);
and U2310 (N_2310,N_1108,N_1236);
or U2311 (N_2311,N_1912,N_1139);
nand U2312 (N_2312,N_1133,N_1184);
nor U2313 (N_2313,N_1568,N_1377);
nor U2314 (N_2314,N_1026,N_1636);
or U2315 (N_2315,N_1663,N_1214);
xnor U2316 (N_2316,N_1137,N_1503);
nand U2317 (N_2317,N_1953,N_1466);
or U2318 (N_2318,N_1687,N_1778);
nand U2319 (N_2319,N_1592,N_1036);
xnor U2320 (N_2320,N_1443,N_1942);
nand U2321 (N_2321,N_1810,N_1878);
xor U2322 (N_2322,N_1872,N_1452);
and U2323 (N_2323,N_1519,N_1575);
xnor U2324 (N_2324,N_1128,N_1545);
xor U2325 (N_2325,N_1668,N_1619);
nand U2326 (N_2326,N_1816,N_1179);
nand U2327 (N_2327,N_1265,N_1250);
or U2328 (N_2328,N_1931,N_1694);
nor U2329 (N_2329,N_1763,N_1431);
and U2330 (N_2330,N_1747,N_1917);
nand U2331 (N_2331,N_1288,N_1414);
or U2332 (N_2332,N_1228,N_1317);
or U2333 (N_2333,N_1893,N_1360);
xor U2334 (N_2334,N_1695,N_1507);
xor U2335 (N_2335,N_1115,N_1371);
xor U2336 (N_2336,N_1383,N_1835);
or U2337 (N_2337,N_1092,N_1268);
or U2338 (N_2338,N_1193,N_1110);
nand U2339 (N_2339,N_1238,N_1764);
and U2340 (N_2340,N_1684,N_1702);
or U2341 (N_2341,N_1031,N_1790);
nor U2342 (N_2342,N_1225,N_1685);
nor U2343 (N_2343,N_1444,N_1802);
nand U2344 (N_2344,N_1791,N_1301);
or U2345 (N_2345,N_1064,N_1785);
nand U2346 (N_2346,N_1201,N_1246);
nand U2347 (N_2347,N_1454,N_1652);
nor U2348 (N_2348,N_1447,N_1935);
nand U2349 (N_2349,N_1223,N_1340);
or U2350 (N_2350,N_1595,N_1255);
and U2351 (N_2351,N_1676,N_1353);
nor U2352 (N_2352,N_1493,N_1833);
xor U2353 (N_2353,N_1121,N_1028);
or U2354 (N_2354,N_1059,N_1646);
nor U2355 (N_2355,N_1591,N_1989);
nand U2356 (N_2356,N_1210,N_1167);
nor U2357 (N_2357,N_1517,N_1083);
xnor U2358 (N_2358,N_1947,N_1409);
nand U2359 (N_2359,N_1617,N_1336);
nand U2360 (N_2360,N_1294,N_1257);
xnor U2361 (N_2361,N_1295,N_1313);
or U2362 (N_2362,N_1969,N_1528);
nor U2363 (N_2363,N_1551,N_1587);
xnor U2364 (N_2364,N_1248,N_1607);
and U2365 (N_2365,N_1889,N_1508);
and U2366 (N_2366,N_1978,N_1800);
xnor U2367 (N_2367,N_1406,N_1939);
nor U2368 (N_2368,N_1742,N_1610);
nor U2369 (N_2369,N_1871,N_1270);
nand U2370 (N_2370,N_1004,N_1983);
nand U2371 (N_2371,N_1578,N_1243);
xor U2372 (N_2372,N_1671,N_1365);
and U2373 (N_2373,N_1675,N_1622);
xnor U2374 (N_2374,N_1891,N_1701);
xor U2375 (N_2375,N_1915,N_1567);
and U2376 (N_2376,N_1162,N_1895);
or U2377 (N_2377,N_1132,N_1260);
nor U2378 (N_2378,N_1870,N_1657);
nand U2379 (N_2379,N_1732,N_1666);
xor U2380 (N_2380,N_1744,N_1002);
nand U2381 (N_2381,N_1141,N_1390);
nand U2382 (N_2382,N_1620,N_1647);
or U2383 (N_2383,N_1752,N_1820);
and U2384 (N_2384,N_1259,N_1471);
and U2385 (N_2385,N_1172,N_1159);
nand U2386 (N_2386,N_1898,N_1902);
or U2387 (N_2387,N_1425,N_1518);
nand U2388 (N_2388,N_1527,N_1883);
xnor U2389 (N_2389,N_1432,N_1152);
or U2390 (N_2390,N_1838,N_1491);
and U2391 (N_2391,N_1326,N_1109);
nand U2392 (N_2392,N_1119,N_1035);
nand U2393 (N_2393,N_1153,N_1310);
xnor U2394 (N_2394,N_1144,N_1879);
nand U2395 (N_2395,N_1706,N_1922);
and U2396 (N_2396,N_1397,N_1533);
nand U2397 (N_2397,N_1698,N_1572);
nand U2398 (N_2398,N_1913,N_1068);
or U2399 (N_2399,N_1465,N_1044);
xnor U2400 (N_2400,N_1505,N_1972);
and U2401 (N_2401,N_1136,N_1892);
or U2402 (N_2402,N_1413,N_1154);
or U2403 (N_2403,N_1395,N_1384);
or U2404 (N_2404,N_1496,N_1649);
nand U2405 (N_2405,N_1558,N_1700);
and U2406 (N_2406,N_1865,N_1556);
xnor U2407 (N_2407,N_1771,N_1051);
xnor U2408 (N_2408,N_1047,N_1453);
or U2409 (N_2409,N_1531,N_1285);
or U2410 (N_2410,N_1597,N_1267);
or U2411 (N_2411,N_1600,N_1089);
nor U2412 (N_2412,N_1314,N_1488);
xor U2413 (N_2413,N_1772,N_1840);
or U2414 (N_2414,N_1613,N_1007);
nor U2415 (N_2415,N_1750,N_1034);
and U2416 (N_2416,N_1874,N_1188);
xnor U2417 (N_2417,N_1271,N_1349);
xnor U2418 (N_2418,N_1580,N_1156);
nor U2419 (N_2419,N_1000,N_1276);
xnor U2420 (N_2420,N_1586,N_1199);
nand U2421 (N_2421,N_1168,N_1486);
nand U2422 (N_2422,N_1423,N_1003);
or U2423 (N_2423,N_1897,N_1641);
xor U2424 (N_2424,N_1088,N_1737);
nand U2425 (N_2425,N_1019,N_1562);
nand U2426 (N_2426,N_1125,N_1337);
nand U2427 (N_2427,N_1692,N_1745);
nand U2428 (N_2428,N_1757,N_1291);
and U2429 (N_2429,N_1506,N_1957);
xor U2430 (N_2430,N_1123,N_1762);
and U2431 (N_2431,N_1900,N_1713);
nand U2432 (N_2432,N_1712,N_1645);
xor U2433 (N_2433,N_1780,N_1629);
or U2434 (N_2434,N_1509,N_1680);
nand U2435 (N_2435,N_1341,N_1596);
or U2436 (N_2436,N_1347,N_1766);
and U2437 (N_2437,N_1025,N_1249);
nand U2438 (N_2438,N_1662,N_1679);
nor U2439 (N_2439,N_1100,N_1277);
or U2440 (N_2440,N_1459,N_1297);
nor U2441 (N_2441,N_1312,N_1069);
or U2442 (N_2442,N_1868,N_1963);
or U2443 (N_2443,N_1292,N_1748);
and U2444 (N_2444,N_1256,N_1196);
nand U2445 (N_2445,N_1399,N_1378);
xor U2446 (N_2446,N_1498,N_1134);
xnor U2447 (N_2447,N_1203,N_1979);
nor U2448 (N_2448,N_1391,N_1951);
or U2449 (N_2449,N_1605,N_1851);
nor U2450 (N_2450,N_1272,N_1195);
or U2451 (N_2451,N_1122,N_1050);
xor U2452 (N_2452,N_1690,N_1220);
xnor U2453 (N_2453,N_1560,N_1135);
xor U2454 (N_2454,N_1473,N_1627);
nor U2455 (N_2455,N_1363,N_1829);
and U2456 (N_2456,N_1407,N_1850);
nor U2457 (N_2457,N_1743,N_1191);
and U2458 (N_2458,N_1062,N_1890);
nand U2459 (N_2459,N_1612,N_1781);
xnor U2460 (N_2460,N_1522,N_1796);
nor U2461 (N_2461,N_1552,N_1072);
xor U2462 (N_2462,N_1628,N_1827);
xor U2463 (N_2463,N_1725,N_1060);
nand U2464 (N_2464,N_1415,N_1094);
xor U2465 (N_2465,N_1346,N_1976);
nand U2466 (N_2466,N_1206,N_1177);
nor U2467 (N_2467,N_1171,N_1603);
xnor U2468 (N_2468,N_1998,N_1847);
xnor U2469 (N_2469,N_1582,N_1251);
or U2470 (N_2470,N_1539,N_1076);
nor U2471 (N_2471,N_1588,N_1116);
nor U2472 (N_2472,N_1357,N_1590);
nor U2473 (N_2473,N_1571,N_1497);
xnor U2474 (N_2474,N_1530,N_1650);
and U2475 (N_2475,N_1308,N_1112);
nand U2476 (N_2476,N_1716,N_1140);
xor U2477 (N_2477,N_1673,N_1286);
xnor U2478 (N_2478,N_1710,N_1323);
xor U2479 (N_2479,N_1105,N_1160);
nor U2480 (N_2480,N_1359,N_1403);
and U2481 (N_2481,N_1434,N_1205);
nand U2482 (N_2482,N_1938,N_1739);
nor U2483 (N_2483,N_1565,N_1958);
or U2484 (N_2484,N_1811,N_1966);
nand U2485 (N_2485,N_1964,N_1579);
nand U2486 (N_2486,N_1985,N_1696);
or U2487 (N_2487,N_1401,N_1343);
xnor U2488 (N_2488,N_1724,N_1746);
and U2489 (N_2489,N_1030,N_1537);
or U2490 (N_2490,N_1651,N_1009);
nand U2491 (N_2491,N_1328,N_1165);
nand U2492 (N_2492,N_1422,N_1933);
or U2493 (N_2493,N_1861,N_1376);
nor U2494 (N_2494,N_1304,N_1660);
or U2495 (N_2495,N_1577,N_1806);
xnor U2496 (N_2496,N_1988,N_1446);
nor U2497 (N_2497,N_1472,N_1398);
and U2498 (N_2498,N_1770,N_1876);
xnor U2499 (N_2499,N_1967,N_1332);
nor U2500 (N_2500,N_1335,N_1204);
xor U2501 (N_2501,N_1087,N_1735);
and U2502 (N_2502,N_1352,N_1649);
nand U2503 (N_2503,N_1236,N_1692);
xnor U2504 (N_2504,N_1756,N_1691);
nor U2505 (N_2505,N_1283,N_1082);
xor U2506 (N_2506,N_1315,N_1137);
nand U2507 (N_2507,N_1529,N_1393);
nand U2508 (N_2508,N_1392,N_1317);
and U2509 (N_2509,N_1395,N_1359);
xnor U2510 (N_2510,N_1795,N_1625);
nor U2511 (N_2511,N_1950,N_1093);
and U2512 (N_2512,N_1697,N_1117);
nand U2513 (N_2513,N_1794,N_1221);
nor U2514 (N_2514,N_1610,N_1334);
nor U2515 (N_2515,N_1226,N_1197);
nand U2516 (N_2516,N_1403,N_1505);
or U2517 (N_2517,N_1419,N_1551);
xor U2518 (N_2518,N_1382,N_1988);
nand U2519 (N_2519,N_1785,N_1619);
or U2520 (N_2520,N_1274,N_1989);
and U2521 (N_2521,N_1962,N_1862);
or U2522 (N_2522,N_1274,N_1172);
or U2523 (N_2523,N_1378,N_1736);
xnor U2524 (N_2524,N_1554,N_1846);
nor U2525 (N_2525,N_1970,N_1550);
nor U2526 (N_2526,N_1454,N_1964);
and U2527 (N_2527,N_1135,N_1498);
xor U2528 (N_2528,N_1444,N_1591);
and U2529 (N_2529,N_1747,N_1545);
or U2530 (N_2530,N_1031,N_1532);
nor U2531 (N_2531,N_1737,N_1672);
or U2532 (N_2532,N_1472,N_1124);
nor U2533 (N_2533,N_1526,N_1757);
or U2534 (N_2534,N_1368,N_1055);
or U2535 (N_2535,N_1236,N_1398);
and U2536 (N_2536,N_1540,N_1705);
nand U2537 (N_2537,N_1175,N_1498);
xnor U2538 (N_2538,N_1602,N_1446);
nor U2539 (N_2539,N_1754,N_1307);
nand U2540 (N_2540,N_1553,N_1480);
nor U2541 (N_2541,N_1149,N_1497);
nor U2542 (N_2542,N_1785,N_1598);
or U2543 (N_2543,N_1673,N_1811);
and U2544 (N_2544,N_1465,N_1383);
nor U2545 (N_2545,N_1576,N_1852);
nand U2546 (N_2546,N_1374,N_1945);
nand U2547 (N_2547,N_1217,N_1947);
nor U2548 (N_2548,N_1925,N_1346);
or U2549 (N_2549,N_1451,N_1955);
xnor U2550 (N_2550,N_1489,N_1806);
or U2551 (N_2551,N_1534,N_1366);
or U2552 (N_2552,N_1080,N_1622);
nor U2553 (N_2553,N_1027,N_1017);
nand U2554 (N_2554,N_1925,N_1083);
and U2555 (N_2555,N_1233,N_1829);
and U2556 (N_2556,N_1882,N_1310);
and U2557 (N_2557,N_1152,N_1398);
and U2558 (N_2558,N_1497,N_1043);
and U2559 (N_2559,N_1099,N_1949);
xnor U2560 (N_2560,N_1531,N_1845);
nor U2561 (N_2561,N_1065,N_1483);
and U2562 (N_2562,N_1658,N_1835);
xnor U2563 (N_2563,N_1223,N_1291);
xor U2564 (N_2564,N_1892,N_1032);
nand U2565 (N_2565,N_1750,N_1328);
nor U2566 (N_2566,N_1891,N_1297);
and U2567 (N_2567,N_1836,N_1656);
nand U2568 (N_2568,N_1876,N_1403);
and U2569 (N_2569,N_1267,N_1657);
or U2570 (N_2570,N_1345,N_1278);
nand U2571 (N_2571,N_1402,N_1130);
xnor U2572 (N_2572,N_1061,N_1672);
and U2573 (N_2573,N_1394,N_1902);
nand U2574 (N_2574,N_1592,N_1354);
and U2575 (N_2575,N_1240,N_1576);
nand U2576 (N_2576,N_1723,N_1833);
nor U2577 (N_2577,N_1469,N_1087);
nor U2578 (N_2578,N_1105,N_1427);
and U2579 (N_2579,N_1167,N_1126);
nand U2580 (N_2580,N_1306,N_1739);
xnor U2581 (N_2581,N_1854,N_1527);
xnor U2582 (N_2582,N_1975,N_1518);
nand U2583 (N_2583,N_1067,N_1504);
nand U2584 (N_2584,N_1049,N_1571);
and U2585 (N_2585,N_1051,N_1758);
nand U2586 (N_2586,N_1765,N_1858);
and U2587 (N_2587,N_1391,N_1690);
nor U2588 (N_2588,N_1230,N_1777);
nand U2589 (N_2589,N_1381,N_1451);
nand U2590 (N_2590,N_1433,N_1927);
xor U2591 (N_2591,N_1090,N_1952);
and U2592 (N_2592,N_1719,N_1291);
nand U2593 (N_2593,N_1275,N_1413);
nand U2594 (N_2594,N_1012,N_1188);
xor U2595 (N_2595,N_1044,N_1958);
and U2596 (N_2596,N_1976,N_1494);
or U2597 (N_2597,N_1658,N_1252);
or U2598 (N_2598,N_1875,N_1955);
xnor U2599 (N_2599,N_1270,N_1925);
and U2600 (N_2600,N_1775,N_1783);
and U2601 (N_2601,N_1772,N_1836);
xor U2602 (N_2602,N_1704,N_1806);
or U2603 (N_2603,N_1482,N_1642);
or U2604 (N_2604,N_1507,N_1995);
nand U2605 (N_2605,N_1135,N_1918);
and U2606 (N_2606,N_1599,N_1200);
xor U2607 (N_2607,N_1949,N_1333);
or U2608 (N_2608,N_1857,N_1125);
xnor U2609 (N_2609,N_1302,N_1279);
or U2610 (N_2610,N_1229,N_1177);
or U2611 (N_2611,N_1543,N_1121);
and U2612 (N_2612,N_1303,N_1098);
and U2613 (N_2613,N_1374,N_1188);
nand U2614 (N_2614,N_1631,N_1948);
and U2615 (N_2615,N_1058,N_1880);
or U2616 (N_2616,N_1856,N_1313);
nand U2617 (N_2617,N_1447,N_1974);
xor U2618 (N_2618,N_1002,N_1969);
nor U2619 (N_2619,N_1419,N_1933);
nor U2620 (N_2620,N_1682,N_1818);
or U2621 (N_2621,N_1307,N_1710);
nand U2622 (N_2622,N_1408,N_1966);
nor U2623 (N_2623,N_1046,N_1865);
xor U2624 (N_2624,N_1893,N_1400);
and U2625 (N_2625,N_1764,N_1662);
or U2626 (N_2626,N_1948,N_1193);
xor U2627 (N_2627,N_1427,N_1674);
nand U2628 (N_2628,N_1306,N_1851);
and U2629 (N_2629,N_1069,N_1390);
xor U2630 (N_2630,N_1423,N_1481);
and U2631 (N_2631,N_1638,N_1564);
xnor U2632 (N_2632,N_1715,N_1499);
nor U2633 (N_2633,N_1927,N_1761);
nand U2634 (N_2634,N_1365,N_1900);
or U2635 (N_2635,N_1353,N_1485);
and U2636 (N_2636,N_1046,N_1496);
and U2637 (N_2637,N_1043,N_1256);
nor U2638 (N_2638,N_1186,N_1783);
nand U2639 (N_2639,N_1109,N_1713);
nand U2640 (N_2640,N_1753,N_1982);
and U2641 (N_2641,N_1327,N_1783);
nand U2642 (N_2642,N_1026,N_1273);
nand U2643 (N_2643,N_1355,N_1658);
nand U2644 (N_2644,N_1038,N_1644);
and U2645 (N_2645,N_1928,N_1562);
nand U2646 (N_2646,N_1651,N_1336);
nor U2647 (N_2647,N_1214,N_1296);
nor U2648 (N_2648,N_1664,N_1136);
and U2649 (N_2649,N_1824,N_1202);
xnor U2650 (N_2650,N_1375,N_1042);
xor U2651 (N_2651,N_1364,N_1208);
nor U2652 (N_2652,N_1690,N_1958);
and U2653 (N_2653,N_1088,N_1561);
and U2654 (N_2654,N_1940,N_1198);
nand U2655 (N_2655,N_1678,N_1116);
nor U2656 (N_2656,N_1761,N_1303);
and U2657 (N_2657,N_1698,N_1740);
nor U2658 (N_2658,N_1286,N_1145);
and U2659 (N_2659,N_1312,N_1762);
or U2660 (N_2660,N_1827,N_1684);
xnor U2661 (N_2661,N_1161,N_1390);
xor U2662 (N_2662,N_1732,N_1243);
xnor U2663 (N_2663,N_1037,N_1058);
nor U2664 (N_2664,N_1347,N_1647);
xor U2665 (N_2665,N_1411,N_1074);
xor U2666 (N_2666,N_1428,N_1595);
nand U2667 (N_2667,N_1845,N_1992);
or U2668 (N_2668,N_1209,N_1258);
and U2669 (N_2669,N_1976,N_1044);
nor U2670 (N_2670,N_1710,N_1750);
and U2671 (N_2671,N_1702,N_1969);
or U2672 (N_2672,N_1173,N_1352);
or U2673 (N_2673,N_1230,N_1143);
or U2674 (N_2674,N_1810,N_1405);
and U2675 (N_2675,N_1599,N_1489);
xor U2676 (N_2676,N_1877,N_1841);
nor U2677 (N_2677,N_1809,N_1588);
or U2678 (N_2678,N_1085,N_1797);
and U2679 (N_2679,N_1760,N_1017);
nand U2680 (N_2680,N_1381,N_1255);
and U2681 (N_2681,N_1027,N_1161);
xor U2682 (N_2682,N_1693,N_1130);
or U2683 (N_2683,N_1256,N_1399);
nor U2684 (N_2684,N_1555,N_1829);
nor U2685 (N_2685,N_1695,N_1824);
xor U2686 (N_2686,N_1870,N_1857);
xor U2687 (N_2687,N_1202,N_1847);
xnor U2688 (N_2688,N_1624,N_1069);
nor U2689 (N_2689,N_1515,N_1129);
nand U2690 (N_2690,N_1750,N_1187);
xnor U2691 (N_2691,N_1318,N_1416);
or U2692 (N_2692,N_1971,N_1209);
xor U2693 (N_2693,N_1802,N_1663);
or U2694 (N_2694,N_1767,N_1923);
nand U2695 (N_2695,N_1490,N_1441);
nand U2696 (N_2696,N_1739,N_1722);
xor U2697 (N_2697,N_1124,N_1018);
xor U2698 (N_2698,N_1547,N_1320);
or U2699 (N_2699,N_1833,N_1000);
or U2700 (N_2700,N_1998,N_1325);
nand U2701 (N_2701,N_1801,N_1844);
xnor U2702 (N_2702,N_1992,N_1002);
xor U2703 (N_2703,N_1448,N_1861);
or U2704 (N_2704,N_1364,N_1529);
nand U2705 (N_2705,N_1408,N_1021);
nand U2706 (N_2706,N_1791,N_1781);
xor U2707 (N_2707,N_1427,N_1495);
nor U2708 (N_2708,N_1705,N_1454);
nand U2709 (N_2709,N_1342,N_1774);
or U2710 (N_2710,N_1387,N_1287);
or U2711 (N_2711,N_1934,N_1399);
and U2712 (N_2712,N_1281,N_1144);
and U2713 (N_2713,N_1390,N_1197);
or U2714 (N_2714,N_1837,N_1194);
nand U2715 (N_2715,N_1589,N_1555);
nand U2716 (N_2716,N_1015,N_1121);
xor U2717 (N_2717,N_1812,N_1347);
nand U2718 (N_2718,N_1484,N_1564);
and U2719 (N_2719,N_1493,N_1852);
nor U2720 (N_2720,N_1832,N_1670);
and U2721 (N_2721,N_1504,N_1996);
nor U2722 (N_2722,N_1913,N_1954);
nand U2723 (N_2723,N_1861,N_1876);
or U2724 (N_2724,N_1283,N_1594);
and U2725 (N_2725,N_1380,N_1916);
and U2726 (N_2726,N_1639,N_1377);
xnor U2727 (N_2727,N_1400,N_1820);
and U2728 (N_2728,N_1508,N_1053);
xnor U2729 (N_2729,N_1501,N_1537);
xnor U2730 (N_2730,N_1242,N_1903);
or U2731 (N_2731,N_1176,N_1018);
and U2732 (N_2732,N_1291,N_1261);
xor U2733 (N_2733,N_1572,N_1670);
nor U2734 (N_2734,N_1499,N_1014);
xnor U2735 (N_2735,N_1704,N_1895);
nand U2736 (N_2736,N_1638,N_1516);
nor U2737 (N_2737,N_1244,N_1742);
nand U2738 (N_2738,N_1409,N_1546);
xor U2739 (N_2739,N_1734,N_1316);
nor U2740 (N_2740,N_1207,N_1062);
xor U2741 (N_2741,N_1720,N_1896);
nor U2742 (N_2742,N_1002,N_1161);
nand U2743 (N_2743,N_1934,N_1266);
nand U2744 (N_2744,N_1161,N_1765);
xnor U2745 (N_2745,N_1176,N_1543);
nand U2746 (N_2746,N_1746,N_1365);
nor U2747 (N_2747,N_1947,N_1904);
xor U2748 (N_2748,N_1811,N_1573);
nor U2749 (N_2749,N_1722,N_1638);
nand U2750 (N_2750,N_1000,N_1112);
nor U2751 (N_2751,N_1957,N_1381);
xnor U2752 (N_2752,N_1505,N_1882);
xnor U2753 (N_2753,N_1829,N_1658);
nand U2754 (N_2754,N_1266,N_1702);
nor U2755 (N_2755,N_1595,N_1241);
xor U2756 (N_2756,N_1298,N_1718);
nor U2757 (N_2757,N_1066,N_1674);
nor U2758 (N_2758,N_1020,N_1164);
xnor U2759 (N_2759,N_1600,N_1883);
or U2760 (N_2760,N_1738,N_1397);
xor U2761 (N_2761,N_1778,N_1992);
and U2762 (N_2762,N_1671,N_1085);
nor U2763 (N_2763,N_1884,N_1032);
xor U2764 (N_2764,N_1298,N_1796);
nor U2765 (N_2765,N_1280,N_1410);
nor U2766 (N_2766,N_1618,N_1755);
nand U2767 (N_2767,N_1153,N_1268);
or U2768 (N_2768,N_1817,N_1574);
nand U2769 (N_2769,N_1267,N_1842);
xor U2770 (N_2770,N_1497,N_1010);
and U2771 (N_2771,N_1303,N_1790);
nand U2772 (N_2772,N_1686,N_1683);
xnor U2773 (N_2773,N_1069,N_1197);
or U2774 (N_2774,N_1927,N_1721);
and U2775 (N_2775,N_1392,N_1718);
nand U2776 (N_2776,N_1351,N_1196);
or U2777 (N_2777,N_1890,N_1639);
or U2778 (N_2778,N_1206,N_1249);
xor U2779 (N_2779,N_1367,N_1761);
and U2780 (N_2780,N_1283,N_1032);
or U2781 (N_2781,N_1402,N_1443);
or U2782 (N_2782,N_1175,N_1698);
nand U2783 (N_2783,N_1440,N_1035);
and U2784 (N_2784,N_1219,N_1901);
xnor U2785 (N_2785,N_1589,N_1069);
xor U2786 (N_2786,N_1264,N_1992);
and U2787 (N_2787,N_1269,N_1914);
xor U2788 (N_2788,N_1858,N_1399);
and U2789 (N_2789,N_1738,N_1960);
and U2790 (N_2790,N_1428,N_1609);
or U2791 (N_2791,N_1079,N_1788);
or U2792 (N_2792,N_1115,N_1751);
nand U2793 (N_2793,N_1522,N_1275);
xnor U2794 (N_2794,N_1831,N_1446);
or U2795 (N_2795,N_1561,N_1380);
nor U2796 (N_2796,N_1252,N_1997);
xor U2797 (N_2797,N_1573,N_1922);
nand U2798 (N_2798,N_1197,N_1217);
nor U2799 (N_2799,N_1015,N_1476);
and U2800 (N_2800,N_1965,N_1202);
or U2801 (N_2801,N_1933,N_1198);
nor U2802 (N_2802,N_1925,N_1483);
or U2803 (N_2803,N_1119,N_1725);
or U2804 (N_2804,N_1041,N_1063);
or U2805 (N_2805,N_1448,N_1692);
nand U2806 (N_2806,N_1499,N_1771);
nand U2807 (N_2807,N_1555,N_1695);
and U2808 (N_2808,N_1970,N_1998);
or U2809 (N_2809,N_1364,N_1710);
nor U2810 (N_2810,N_1517,N_1978);
and U2811 (N_2811,N_1129,N_1355);
nor U2812 (N_2812,N_1307,N_1711);
or U2813 (N_2813,N_1526,N_1864);
nor U2814 (N_2814,N_1590,N_1702);
xnor U2815 (N_2815,N_1833,N_1420);
xor U2816 (N_2816,N_1170,N_1609);
nand U2817 (N_2817,N_1584,N_1745);
nor U2818 (N_2818,N_1077,N_1514);
nor U2819 (N_2819,N_1772,N_1050);
nand U2820 (N_2820,N_1064,N_1521);
xor U2821 (N_2821,N_1502,N_1518);
and U2822 (N_2822,N_1798,N_1927);
or U2823 (N_2823,N_1564,N_1589);
or U2824 (N_2824,N_1510,N_1046);
nor U2825 (N_2825,N_1887,N_1346);
or U2826 (N_2826,N_1256,N_1946);
or U2827 (N_2827,N_1925,N_1956);
xor U2828 (N_2828,N_1469,N_1450);
or U2829 (N_2829,N_1638,N_1873);
nand U2830 (N_2830,N_1063,N_1752);
and U2831 (N_2831,N_1643,N_1885);
or U2832 (N_2832,N_1726,N_1578);
and U2833 (N_2833,N_1623,N_1074);
and U2834 (N_2834,N_1266,N_1070);
nand U2835 (N_2835,N_1813,N_1597);
nand U2836 (N_2836,N_1140,N_1248);
xor U2837 (N_2837,N_1851,N_1184);
xor U2838 (N_2838,N_1168,N_1733);
xnor U2839 (N_2839,N_1314,N_1103);
xor U2840 (N_2840,N_1289,N_1652);
xnor U2841 (N_2841,N_1800,N_1121);
and U2842 (N_2842,N_1979,N_1131);
nand U2843 (N_2843,N_1563,N_1198);
or U2844 (N_2844,N_1327,N_1186);
or U2845 (N_2845,N_1915,N_1269);
xnor U2846 (N_2846,N_1145,N_1639);
nor U2847 (N_2847,N_1940,N_1145);
and U2848 (N_2848,N_1067,N_1697);
xnor U2849 (N_2849,N_1499,N_1802);
or U2850 (N_2850,N_1123,N_1274);
nand U2851 (N_2851,N_1776,N_1686);
or U2852 (N_2852,N_1433,N_1607);
or U2853 (N_2853,N_1382,N_1843);
nor U2854 (N_2854,N_1581,N_1904);
or U2855 (N_2855,N_1734,N_1968);
or U2856 (N_2856,N_1078,N_1587);
and U2857 (N_2857,N_1216,N_1253);
and U2858 (N_2858,N_1524,N_1399);
and U2859 (N_2859,N_1986,N_1038);
or U2860 (N_2860,N_1851,N_1507);
xnor U2861 (N_2861,N_1494,N_1952);
nand U2862 (N_2862,N_1662,N_1485);
or U2863 (N_2863,N_1972,N_1324);
xor U2864 (N_2864,N_1889,N_1464);
nor U2865 (N_2865,N_1731,N_1929);
and U2866 (N_2866,N_1388,N_1094);
or U2867 (N_2867,N_1674,N_1538);
or U2868 (N_2868,N_1667,N_1687);
and U2869 (N_2869,N_1457,N_1275);
xnor U2870 (N_2870,N_1642,N_1361);
and U2871 (N_2871,N_1399,N_1899);
and U2872 (N_2872,N_1590,N_1715);
or U2873 (N_2873,N_1787,N_1340);
nand U2874 (N_2874,N_1368,N_1826);
and U2875 (N_2875,N_1051,N_1227);
and U2876 (N_2876,N_1683,N_1728);
xor U2877 (N_2877,N_1123,N_1137);
nand U2878 (N_2878,N_1899,N_1657);
nor U2879 (N_2879,N_1155,N_1285);
or U2880 (N_2880,N_1655,N_1029);
nand U2881 (N_2881,N_1105,N_1410);
nor U2882 (N_2882,N_1242,N_1410);
and U2883 (N_2883,N_1625,N_1747);
xnor U2884 (N_2884,N_1694,N_1276);
nand U2885 (N_2885,N_1817,N_1785);
xnor U2886 (N_2886,N_1850,N_1598);
nor U2887 (N_2887,N_1487,N_1610);
nand U2888 (N_2888,N_1129,N_1720);
nor U2889 (N_2889,N_1614,N_1059);
or U2890 (N_2890,N_1509,N_1180);
and U2891 (N_2891,N_1422,N_1877);
xnor U2892 (N_2892,N_1781,N_1629);
nor U2893 (N_2893,N_1988,N_1595);
or U2894 (N_2894,N_1449,N_1571);
nand U2895 (N_2895,N_1661,N_1864);
nand U2896 (N_2896,N_1301,N_1103);
or U2897 (N_2897,N_1007,N_1165);
nor U2898 (N_2898,N_1039,N_1438);
and U2899 (N_2899,N_1968,N_1797);
and U2900 (N_2900,N_1025,N_1683);
nand U2901 (N_2901,N_1045,N_1545);
and U2902 (N_2902,N_1489,N_1476);
nor U2903 (N_2903,N_1429,N_1424);
xor U2904 (N_2904,N_1587,N_1362);
nand U2905 (N_2905,N_1383,N_1378);
or U2906 (N_2906,N_1150,N_1947);
nor U2907 (N_2907,N_1626,N_1415);
or U2908 (N_2908,N_1892,N_1825);
nor U2909 (N_2909,N_1917,N_1347);
or U2910 (N_2910,N_1189,N_1969);
xor U2911 (N_2911,N_1123,N_1867);
nor U2912 (N_2912,N_1241,N_1060);
or U2913 (N_2913,N_1087,N_1433);
nand U2914 (N_2914,N_1884,N_1131);
xor U2915 (N_2915,N_1591,N_1883);
nor U2916 (N_2916,N_1755,N_1843);
or U2917 (N_2917,N_1459,N_1438);
xor U2918 (N_2918,N_1614,N_1097);
or U2919 (N_2919,N_1894,N_1639);
or U2920 (N_2920,N_1063,N_1620);
or U2921 (N_2921,N_1817,N_1206);
and U2922 (N_2922,N_1267,N_1209);
and U2923 (N_2923,N_1533,N_1065);
nor U2924 (N_2924,N_1212,N_1197);
and U2925 (N_2925,N_1217,N_1269);
or U2926 (N_2926,N_1121,N_1584);
and U2927 (N_2927,N_1819,N_1084);
nand U2928 (N_2928,N_1365,N_1213);
nor U2929 (N_2929,N_1129,N_1034);
nand U2930 (N_2930,N_1561,N_1905);
and U2931 (N_2931,N_1550,N_1538);
or U2932 (N_2932,N_1273,N_1085);
and U2933 (N_2933,N_1142,N_1371);
or U2934 (N_2934,N_1596,N_1940);
nor U2935 (N_2935,N_1624,N_1694);
xor U2936 (N_2936,N_1676,N_1359);
nand U2937 (N_2937,N_1676,N_1957);
xnor U2938 (N_2938,N_1386,N_1989);
nor U2939 (N_2939,N_1184,N_1268);
nand U2940 (N_2940,N_1452,N_1136);
nand U2941 (N_2941,N_1846,N_1806);
nor U2942 (N_2942,N_1679,N_1128);
or U2943 (N_2943,N_1965,N_1677);
nor U2944 (N_2944,N_1232,N_1797);
or U2945 (N_2945,N_1231,N_1300);
nor U2946 (N_2946,N_1833,N_1656);
nor U2947 (N_2947,N_1751,N_1459);
and U2948 (N_2948,N_1879,N_1649);
xor U2949 (N_2949,N_1600,N_1791);
and U2950 (N_2950,N_1959,N_1818);
nand U2951 (N_2951,N_1499,N_1904);
and U2952 (N_2952,N_1909,N_1928);
or U2953 (N_2953,N_1466,N_1270);
and U2954 (N_2954,N_1085,N_1044);
nor U2955 (N_2955,N_1454,N_1069);
nand U2956 (N_2956,N_1890,N_1833);
or U2957 (N_2957,N_1776,N_1861);
nor U2958 (N_2958,N_1441,N_1904);
nor U2959 (N_2959,N_1700,N_1083);
nor U2960 (N_2960,N_1012,N_1944);
and U2961 (N_2961,N_1352,N_1176);
nand U2962 (N_2962,N_1771,N_1385);
nand U2963 (N_2963,N_1714,N_1021);
or U2964 (N_2964,N_1342,N_1704);
and U2965 (N_2965,N_1199,N_1811);
or U2966 (N_2966,N_1842,N_1606);
xnor U2967 (N_2967,N_1926,N_1680);
or U2968 (N_2968,N_1487,N_1594);
nor U2969 (N_2969,N_1958,N_1319);
or U2970 (N_2970,N_1535,N_1600);
nand U2971 (N_2971,N_1943,N_1197);
nor U2972 (N_2972,N_1192,N_1999);
and U2973 (N_2973,N_1769,N_1678);
or U2974 (N_2974,N_1756,N_1409);
or U2975 (N_2975,N_1550,N_1284);
and U2976 (N_2976,N_1313,N_1930);
nand U2977 (N_2977,N_1314,N_1576);
nor U2978 (N_2978,N_1568,N_1355);
nand U2979 (N_2979,N_1946,N_1448);
and U2980 (N_2980,N_1559,N_1868);
or U2981 (N_2981,N_1986,N_1567);
or U2982 (N_2982,N_1902,N_1351);
nor U2983 (N_2983,N_1692,N_1335);
xor U2984 (N_2984,N_1248,N_1216);
and U2985 (N_2985,N_1612,N_1117);
nand U2986 (N_2986,N_1357,N_1097);
or U2987 (N_2987,N_1590,N_1594);
nor U2988 (N_2988,N_1700,N_1119);
and U2989 (N_2989,N_1192,N_1840);
xor U2990 (N_2990,N_1905,N_1593);
and U2991 (N_2991,N_1628,N_1449);
and U2992 (N_2992,N_1686,N_1073);
nor U2993 (N_2993,N_1543,N_1364);
and U2994 (N_2994,N_1057,N_1465);
or U2995 (N_2995,N_1710,N_1206);
xor U2996 (N_2996,N_1074,N_1892);
nand U2997 (N_2997,N_1401,N_1968);
and U2998 (N_2998,N_1799,N_1021);
nand U2999 (N_2999,N_1276,N_1731);
xor U3000 (N_3000,N_2973,N_2049);
xnor U3001 (N_3001,N_2608,N_2750);
or U3002 (N_3002,N_2508,N_2219);
or U3003 (N_3003,N_2194,N_2812);
nand U3004 (N_3004,N_2776,N_2343);
and U3005 (N_3005,N_2994,N_2493);
nand U3006 (N_3006,N_2753,N_2984);
nand U3007 (N_3007,N_2141,N_2490);
or U3008 (N_3008,N_2624,N_2284);
or U3009 (N_3009,N_2247,N_2023);
or U3010 (N_3010,N_2839,N_2547);
nor U3011 (N_3011,N_2091,N_2925);
nor U3012 (N_3012,N_2859,N_2110);
and U3013 (N_3013,N_2788,N_2897);
and U3014 (N_3014,N_2068,N_2342);
nand U3015 (N_3015,N_2852,N_2965);
and U3016 (N_3016,N_2726,N_2321);
nand U3017 (N_3017,N_2885,N_2456);
xor U3018 (N_3018,N_2792,N_2677);
and U3019 (N_3019,N_2798,N_2265);
or U3020 (N_3020,N_2675,N_2283);
nor U3021 (N_3021,N_2511,N_2730);
or U3022 (N_3022,N_2097,N_2768);
nand U3023 (N_3023,N_2656,N_2356);
and U3024 (N_3024,N_2276,N_2101);
and U3025 (N_3025,N_2992,N_2563);
or U3026 (N_3026,N_2825,N_2209);
nand U3027 (N_3027,N_2880,N_2519);
xnor U3028 (N_3028,N_2902,N_2290);
nand U3029 (N_3029,N_2771,N_2257);
or U3030 (N_3030,N_2549,N_2597);
xnor U3031 (N_3031,N_2454,N_2757);
nand U3032 (N_3032,N_2630,N_2680);
nor U3033 (N_3033,N_2400,N_2186);
xnor U3034 (N_3034,N_2772,N_2015);
xor U3035 (N_3035,N_2893,N_2020);
nor U3036 (N_3036,N_2762,N_2940);
xor U3037 (N_3037,N_2409,N_2153);
or U3038 (N_3038,N_2924,N_2410);
or U3039 (N_3039,N_2561,N_2138);
or U3040 (N_3040,N_2007,N_2044);
nand U3041 (N_3041,N_2710,N_2124);
and U3042 (N_3042,N_2297,N_2235);
or U3043 (N_3043,N_2039,N_2244);
nand U3044 (N_3044,N_2018,N_2424);
nand U3045 (N_3045,N_2657,N_2942);
nor U3046 (N_3046,N_2134,N_2793);
nand U3047 (N_3047,N_2129,N_2104);
nor U3048 (N_3048,N_2031,N_2197);
nor U3049 (N_3049,N_2051,N_2906);
nor U3050 (N_3050,N_2160,N_2874);
or U3051 (N_3051,N_2105,N_2215);
xor U3052 (N_3052,N_2899,N_2483);
xnor U3053 (N_3053,N_2616,N_2352);
nor U3054 (N_3054,N_2972,N_2954);
or U3055 (N_3055,N_2045,N_2208);
and U3056 (N_3056,N_2056,N_2399);
or U3057 (N_3057,N_2698,N_2350);
xor U3058 (N_3058,N_2095,N_2347);
and U3059 (N_3059,N_2038,N_2166);
xnor U3060 (N_3060,N_2791,N_2365);
and U3061 (N_3061,N_2345,N_2494);
nor U3062 (N_3062,N_2133,N_2724);
and U3063 (N_3063,N_2152,N_2576);
nand U3064 (N_3064,N_2654,N_2921);
nand U3065 (N_3065,N_2504,N_2575);
or U3066 (N_3066,N_2505,N_2195);
nand U3067 (N_3067,N_2452,N_2571);
or U3068 (N_3068,N_2125,N_2836);
xor U3069 (N_3069,N_2484,N_2869);
nand U3070 (N_3070,N_2299,N_2453);
or U3071 (N_3071,N_2474,N_2282);
and U3072 (N_3072,N_2557,N_2733);
or U3073 (N_3073,N_2327,N_2055);
nand U3074 (N_3074,N_2446,N_2043);
or U3075 (N_3075,N_2574,N_2736);
nor U3076 (N_3076,N_2064,N_2976);
nand U3077 (N_3077,N_2422,N_2932);
and U3078 (N_3078,N_2222,N_2722);
nor U3079 (N_3079,N_2469,N_2503);
nor U3080 (N_3080,N_2185,N_2671);
or U3081 (N_3081,N_2151,N_2473);
xor U3082 (N_3082,N_2599,N_2059);
xnor U3083 (N_3083,N_2876,N_2635);
xor U3084 (N_3084,N_2079,N_2866);
nor U3085 (N_3085,N_2602,N_2956);
nand U3086 (N_3086,N_2568,N_2263);
xnor U3087 (N_3087,N_2041,N_2692);
xnor U3088 (N_3088,N_2864,N_2584);
nand U3089 (N_3089,N_2022,N_2298);
nand U3090 (N_3090,N_2790,N_2457);
nor U3091 (N_3091,N_2117,N_2950);
nand U3092 (N_3092,N_2036,N_2867);
nand U3093 (N_3093,N_2759,N_2200);
nand U3094 (N_3094,N_2914,N_2649);
or U3095 (N_3095,N_2471,N_2379);
nand U3096 (N_3096,N_2711,N_2781);
xor U3097 (N_3097,N_2851,N_2006);
and U3098 (N_3098,N_2936,N_2818);
nand U3099 (N_3099,N_2248,N_2307);
or U3100 (N_3100,N_2386,N_2164);
and U3101 (N_3101,N_2898,N_2233);
nor U3102 (N_3102,N_2854,N_2609);
and U3103 (N_3103,N_2188,N_2312);
nor U3104 (N_3104,N_2580,N_2011);
or U3105 (N_3105,N_2252,N_2319);
xor U3106 (N_3106,N_2841,N_2001);
or U3107 (N_3107,N_2491,N_2534);
nor U3108 (N_3108,N_2989,N_2699);
xnor U3109 (N_3109,N_2767,N_2966);
nor U3110 (N_3110,N_2857,N_2934);
or U3111 (N_3111,N_2032,N_2081);
and U3112 (N_3112,N_2017,N_2288);
or U3113 (N_3113,N_2048,N_2178);
and U3114 (N_3114,N_2529,N_2458);
nor U3115 (N_3115,N_2427,N_2074);
or U3116 (N_3116,N_2909,N_2196);
or U3117 (N_3117,N_2643,N_2465);
or U3118 (N_3118,N_2951,N_2660);
and U3119 (N_3119,N_2860,N_2943);
or U3120 (N_3120,N_2702,N_2187);
and U3121 (N_3121,N_2294,N_2640);
nor U3122 (N_3122,N_2224,N_2856);
xor U3123 (N_3123,N_2392,N_2106);
nand U3124 (N_3124,N_2535,N_2611);
or U3125 (N_3125,N_2337,N_2167);
nand U3126 (N_3126,N_2203,N_2947);
nand U3127 (N_3127,N_2567,N_2175);
nand U3128 (N_3128,N_2112,N_2644);
nand U3129 (N_3129,N_2232,N_2277);
and U3130 (N_3130,N_2174,N_2501);
xnor U3131 (N_3131,N_2542,N_2132);
or U3132 (N_3132,N_2681,N_2123);
nand U3133 (N_3133,N_2614,N_2182);
xnor U3134 (N_3134,N_2538,N_2517);
nor U3135 (N_3135,N_2676,N_2751);
or U3136 (N_3136,N_2945,N_2543);
nand U3137 (N_3137,N_2046,N_2809);
nor U3138 (N_3138,N_2027,N_2369);
or U3139 (N_3139,N_2553,N_2340);
and U3140 (N_3140,N_2601,N_2536);
nor U3141 (N_3141,N_2506,N_2009);
and U3142 (N_3142,N_2663,N_2833);
and U3143 (N_3143,N_2295,N_2326);
xnor U3144 (N_3144,N_2354,N_2374);
nand U3145 (N_3145,N_2367,N_2202);
xnor U3146 (N_3146,N_2192,N_2764);
or U3147 (N_3147,N_2709,N_2338);
nand U3148 (N_3148,N_2548,N_2376);
nand U3149 (N_3149,N_2468,N_2708);
or U3150 (N_3150,N_2755,N_2849);
nand U3151 (N_3151,N_2887,N_2334);
xnor U3152 (N_3152,N_2441,N_2370);
nand U3153 (N_3153,N_2066,N_2477);
xor U3154 (N_3154,N_2440,N_2245);
or U3155 (N_3155,N_2403,N_2844);
nand U3156 (N_3156,N_2689,N_2974);
and U3157 (N_3157,N_2894,N_2627);
nand U3158 (N_3158,N_2946,N_2981);
and U3159 (N_3159,N_2439,N_2638);
xnor U3160 (N_3160,N_2390,N_2804);
and U3161 (N_3161,N_2889,N_2479);
xor U3162 (N_3162,N_2811,N_2274);
nor U3163 (N_3163,N_2432,N_2131);
or U3164 (N_3164,N_2513,N_2729);
or U3165 (N_3165,N_2908,N_2805);
and U3166 (N_3166,N_2230,N_2193);
nand U3167 (N_3167,N_2189,N_2030);
nand U3168 (N_3168,N_2959,N_2114);
xor U3169 (N_3169,N_2533,N_2314);
and U3170 (N_3170,N_2637,N_2096);
or U3171 (N_3171,N_2107,N_2785);
or U3172 (N_3172,N_2619,N_2537);
nand U3173 (N_3173,N_2148,N_2080);
xnor U3174 (N_3174,N_2691,N_2273);
or U3175 (N_3175,N_2564,N_2871);
and U3176 (N_3176,N_2429,N_2728);
xor U3177 (N_3177,N_2413,N_2615);
nor U3178 (N_3178,N_2891,N_2156);
xnor U3179 (N_3179,N_2489,N_2863);
xor U3180 (N_3180,N_2645,N_2987);
and U3181 (N_3181,N_2977,N_2870);
and U3182 (N_3182,N_2855,N_2569);
or U3183 (N_3183,N_2396,N_2648);
xor U3184 (N_3184,N_2888,N_2366);
nand U3185 (N_3185,N_2301,N_2378);
xor U3186 (N_3186,N_2651,N_2398);
nor U3187 (N_3187,N_2831,N_2344);
nor U3188 (N_3188,N_2258,N_2165);
or U3189 (N_3189,N_2500,N_2223);
xor U3190 (N_3190,N_2596,N_2389);
xnor U3191 (N_3191,N_2442,N_2103);
or U3192 (N_3192,N_2975,N_2652);
and U3193 (N_3193,N_2917,N_2169);
and U3194 (N_3194,N_2406,N_2672);
nand U3195 (N_3195,N_2475,N_2270);
nand U3196 (N_3196,N_2998,N_2142);
nor U3197 (N_3197,N_2929,N_2029);
nor U3198 (N_3198,N_2361,N_2428);
or U3199 (N_3199,N_2019,N_2911);
and U3200 (N_3200,N_2100,N_2521);
and U3201 (N_3201,N_2430,N_2184);
and U3202 (N_3202,N_2901,N_2589);
or U3203 (N_3203,N_2254,N_2734);
xnor U3204 (N_3204,N_2316,N_2618);
nand U3205 (N_3205,N_2878,N_2421);
nor U3206 (N_3206,N_2317,N_2359);
nor U3207 (N_3207,N_2154,N_2122);
or U3208 (N_3208,N_2808,N_2799);
or U3209 (N_3209,N_2118,N_2664);
nand U3210 (N_3210,N_2279,N_2000);
and U3211 (N_3211,N_2752,N_2843);
xor U3212 (N_3212,N_2250,N_2229);
nor U3213 (N_3213,N_2336,N_2748);
or U3214 (N_3214,N_2806,N_2935);
or U3215 (N_3215,N_2613,N_2948);
or U3216 (N_3216,N_2666,N_2587);
nand U3217 (N_3217,N_2732,N_2016);
or U3218 (N_3218,N_2621,N_2173);
and U3219 (N_3219,N_2402,N_2737);
nor U3220 (N_3220,N_2585,N_2783);
nor U3221 (N_3221,N_2289,N_2706);
nand U3222 (N_3222,N_2071,N_2008);
or U3223 (N_3223,N_2249,N_2719);
xor U3224 (N_3224,N_2397,N_2552);
xnor U3225 (N_3225,N_2139,N_2647);
or U3226 (N_3226,N_2979,N_2447);
nand U3227 (N_3227,N_2784,N_2915);
nor U3228 (N_3228,N_2920,N_2723);
nor U3229 (N_3229,N_2941,N_2499);
and U3230 (N_3230,N_2582,N_2577);
or U3231 (N_3231,N_2172,N_2181);
or U3232 (N_3232,N_2829,N_2050);
and U3233 (N_3233,N_2617,N_2512);
or U3234 (N_3234,N_2612,N_2769);
nand U3235 (N_3235,N_2639,N_2416);
nand U3236 (N_3236,N_2971,N_2158);
or U3237 (N_3237,N_2659,N_2267);
or U3238 (N_3238,N_2655,N_2522);
or U3239 (N_3239,N_2291,N_2381);
nand U3240 (N_3240,N_2143,N_2296);
or U3241 (N_3241,N_2873,N_2982);
or U3242 (N_3242,N_2024,N_2339);
and U3243 (N_3243,N_2275,N_2944);
or U3244 (N_3244,N_2451,N_2961);
nand U3245 (N_3245,N_2685,N_2445);
xor U3246 (N_3246,N_2845,N_2418);
and U3247 (N_3247,N_2625,N_2094);
nor U3248 (N_3248,N_2905,N_2955);
xnor U3249 (N_3249,N_2037,N_2077);
nor U3250 (N_3250,N_2882,N_2305);
nor U3251 (N_3251,N_2003,N_2720);
xor U3252 (N_3252,N_2526,N_2658);
nor U3253 (N_3253,N_2532,N_2434);
xnor U3254 (N_3254,N_2260,N_2555);
xor U3255 (N_3255,N_2687,N_2444);
xor U3256 (N_3256,N_2251,N_2813);
xor U3257 (N_3257,N_2650,N_2419);
or U3258 (N_3258,N_2240,N_2395);
nand U3259 (N_3259,N_2821,N_2383);
nand U3260 (N_3260,N_2060,N_2155);
or U3261 (N_3261,N_2488,N_2286);
or U3262 (N_3262,N_2388,N_2877);
or U3263 (N_3263,N_2357,N_2999);
xnor U3264 (N_3264,N_2329,N_2147);
nand U3265 (N_3265,N_2405,N_2372);
and U3266 (N_3266,N_2495,N_2042);
and U3267 (N_3267,N_2626,N_2377);
xnor U3268 (N_3268,N_2157,N_2448);
or U3269 (N_3269,N_2610,N_2727);
nor U3270 (N_3270,N_2819,N_2515);
nor U3271 (N_3271,N_2697,N_2211);
xnor U3272 (N_3272,N_2603,N_2803);
nor U3273 (N_3273,N_2335,N_2120);
nand U3274 (N_3274,N_2756,N_2606);
or U3275 (N_3275,N_2330,N_2144);
and U3276 (N_3276,N_2628,N_2775);
xnor U3277 (N_3277,N_2594,N_2514);
or U3278 (N_3278,N_2665,N_2591);
nand U3279 (N_3279,N_2472,N_2140);
and U3280 (N_3280,N_2426,N_2331);
nand U3281 (N_3281,N_2486,N_2528);
or U3282 (N_3282,N_2743,N_2896);
or U3283 (N_3283,N_2206,N_2739);
and U3284 (N_3284,N_2242,N_2588);
nor U3285 (N_3285,N_2358,N_2904);
xnor U3286 (N_3286,N_2082,N_2363);
xor U3287 (N_3287,N_2810,N_2180);
and U3288 (N_3288,N_2320,N_2835);
xor U3289 (N_3289,N_2725,N_2765);
xor U3290 (N_3290,N_2108,N_2669);
nor U3291 (N_3291,N_2963,N_2065);
or U3292 (N_3292,N_2470,N_2923);
or U3293 (N_3293,N_2559,N_2098);
nor U3294 (N_3294,N_2927,N_2881);
or U3295 (N_3295,N_2969,N_2115);
nand U3296 (N_3296,N_2570,N_2579);
nand U3297 (N_3297,N_2498,N_2145);
nor U3298 (N_3298,N_2128,N_2231);
or U3299 (N_3299,N_2773,N_2130);
nor U3300 (N_3300,N_2436,N_2938);
nand U3301 (N_3301,N_2707,N_2323);
nor U3302 (N_3302,N_2482,N_2527);
and U3303 (N_3303,N_2986,N_2238);
nand U3304 (N_3304,N_2745,N_2464);
and U3305 (N_3305,N_2126,N_2341);
or U3306 (N_3306,N_2777,N_2673);
nand U3307 (N_3307,N_2268,N_2102);
nor U3308 (N_3308,N_2520,N_2467);
xnor U3309 (N_3309,N_2928,N_2086);
or U3310 (N_3310,N_2304,N_2485);
and U3311 (N_3311,N_2246,N_2414);
nand U3312 (N_3312,N_2420,N_2269);
or U3313 (N_3313,N_2415,N_2237);
nand U3314 (N_3314,N_2822,N_2324);
nor U3315 (N_3315,N_2315,N_2820);
nand U3316 (N_3316,N_2113,N_2502);
and U3317 (N_3317,N_2243,N_2682);
xor U3318 (N_3318,N_2510,N_2539);
and U3319 (N_3319,N_2070,N_2480);
xnor U3320 (N_3320,N_2900,N_2620);
nand U3321 (N_3321,N_2583,N_2278);
nor U3322 (N_3322,N_2700,N_2631);
xor U3323 (N_3323,N_2010,N_2487);
or U3324 (N_3324,N_2742,N_2088);
nor U3325 (N_3325,N_2013,N_2253);
and U3326 (N_3326,N_2207,N_2837);
or U3327 (N_3327,N_2668,N_2912);
xnor U3328 (N_3328,N_2595,N_2199);
xnor U3329 (N_3329,N_2816,N_2721);
nand U3330 (N_3330,N_2558,N_2696);
nand U3331 (N_3331,N_2364,N_2228);
nor U3332 (N_3332,N_2481,N_2057);
or U3333 (N_3333,N_2496,N_2546);
xor U3334 (N_3334,N_2217,N_2629);
and U3335 (N_3335,N_2308,N_2411);
and U3336 (N_3336,N_2531,N_2201);
or U3337 (N_3337,N_2162,N_2449);
xor U3338 (N_3338,N_2779,N_2394);
nand U3339 (N_3339,N_2313,N_2566);
nand U3340 (N_3340,N_2221,N_2256);
or U3341 (N_3341,N_2084,N_2530);
xor U3342 (N_3342,N_2592,N_2600);
or U3343 (N_3343,N_2333,N_2853);
and U3344 (N_3344,N_2826,N_2425);
nor U3345 (N_3345,N_2089,N_2695);
nand U3346 (N_3346,N_2264,N_2712);
xnor U3347 (N_3347,N_2868,N_2438);
nor U3348 (N_3348,N_2052,N_2949);
and U3349 (N_3349,N_2646,N_2581);
and U3350 (N_3350,N_2259,N_2507);
nand U3351 (N_3351,N_2679,N_2962);
xor U3352 (N_3352,N_2814,N_2827);
or U3353 (N_3353,N_2910,N_2300);
xnor U3354 (N_3354,N_2832,N_2271);
and U3355 (N_3355,N_2346,N_2541);
nand U3356 (N_3356,N_2433,N_2562);
nand U3357 (N_3357,N_2287,N_2879);
xor U3358 (N_3358,N_2703,N_2353);
xnor U3359 (N_3359,N_2239,N_2028);
nand U3360 (N_3360,N_2075,N_2328);
nand U3361 (N_3361,N_2968,N_2450);
nor U3362 (N_3362,N_2492,N_2062);
and U3363 (N_3363,N_2761,N_2760);
and U3364 (N_3364,N_2985,N_2701);
or U3365 (N_3365,N_2593,N_2926);
or U3366 (N_3366,N_2774,N_2861);
nand U3367 (N_3367,N_2033,N_2318);
and U3368 (N_3368,N_2572,N_2800);
and U3369 (N_3369,N_2190,N_2306);
and U3370 (N_3370,N_2713,N_2466);
and U3371 (N_3371,N_2476,N_2807);
or U3372 (N_3372,N_2407,N_2127);
xor U3373 (N_3373,N_2842,N_2636);
nor U3374 (N_3374,N_2053,N_2838);
nand U3375 (N_3375,N_2463,N_2633);
nor U3376 (N_3376,N_2005,N_2325);
or U3377 (N_3377,N_2205,N_2198);
and U3378 (N_3378,N_2653,N_2021);
nor U3379 (N_3379,N_2303,N_2933);
nor U3380 (N_3380,N_2795,N_2310);
and U3381 (N_3381,N_2778,N_2092);
and U3382 (N_3382,N_2311,N_2964);
xor U3383 (N_3383,N_2280,N_2754);
nor U3384 (N_3384,N_2996,N_2216);
nand U3385 (N_3385,N_2550,N_2740);
xnor U3386 (N_3386,N_2136,N_2116);
nand U3387 (N_3387,N_2978,N_2437);
xor U3388 (N_3388,N_2161,N_2302);
nand U3389 (N_3389,N_2758,N_2266);
nand U3390 (N_3390,N_2360,N_2509);
nand U3391 (N_3391,N_2622,N_2850);
or U3392 (N_3392,N_2401,N_2741);
xor U3393 (N_3393,N_2847,N_2980);
nor U3394 (N_3394,N_2385,N_2191);
or U3395 (N_3395,N_2830,N_2632);
and U3396 (N_3396,N_2525,N_2524);
nor U3397 (N_3397,N_2738,N_2078);
xnor U3398 (N_3398,N_2380,N_2607);
or U3399 (N_3399,N_2796,N_2460);
or U3400 (N_3400,N_2309,N_2014);
xor U3401 (N_3401,N_2705,N_2214);
nor U3402 (N_3402,N_2993,N_2391);
nand U3403 (N_3403,N_2349,N_2171);
nand U3404 (N_3404,N_2693,N_2293);
xnor U3405 (N_3405,N_2261,N_2953);
xnor U3406 (N_3406,N_2351,N_2149);
nand U3407 (N_3407,N_2642,N_2137);
nor U3408 (N_3408,N_2997,N_2907);
or U3409 (N_3409,N_2034,N_2236);
and U3410 (N_3410,N_2002,N_2227);
nor U3411 (N_3411,N_2012,N_2952);
or U3412 (N_3412,N_2431,N_2858);
xnor U3413 (N_3413,N_2717,N_2272);
nor U3414 (N_3414,N_2170,N_2087);
and U3415 (N_3415,N_2076,N_2970);
nand U3416 (N_3416,N_2694,N_2573);
or U3417 (N_3417,N_2213,N_2801);
nor U3418 (N_3418,N_2744,N_2786);
xor U3419 (N_3419,N_2135,N_2047);
nor U3420 (N_3420,N_2718,N_2478);
or U3421 (N_3421,N_2085,N_2332);
xnor U3422 (N_3422,N_2382,N_2459);
or U3423 (N_3423,N_2794,N_2348);
or U3424 (N_3424,N_2417,N_2119);
and U3425 (N_3425,N_2824,N_2040);
nand U3426 (N_3426,N_2111,N_2072);
nor U3427 (N_3427,N_2674,N_2281);
nand U3428 (N_3428,N_2913,N_2605);
and U3429 (N_3429,N_2886,N_2890);
or U3430 (N_3430,N_2735,N_2225);
or U3431 (N_3431,N_2146,N_2983);
and U3432 (N_3432,N_2523,N_2285);
or U3433 (N_3433,N_2516,N_2789);
nor U3434 (N_3434,N_2556,N_2061);
nor U3435 (N_3435,N_2919,N_2026);
xor U3436 (N_3436,N_2183,N_2883);
and U3437 (N_3437,N_2895,N_2497);
xnor U3438 (N_3438,N_2404,N_2766);
nor U3439 (N_3439,N_2960,N_2641);
and U3440 (N_3440,N_2875,N_2518);
or U3441 (N_3441,N_2545,N_2939);
or U3442 (N_3442,N_2931,N_2565);
and U3443 (N_3443,N_2846,N_2025);
nand U3444 (N_3444,N_2544,N_2930);
or U3445 (N_3445,N_2226,N_2443);
and U3446 (N_3446,N_2937,N_2678);
or U3447 (N_3447,N_2035,N_2918);
xnor U3448 (N_3448,N_2922,N_2780);
nand U3449 (N_3449,N_2865,N_2099);
or U3450 (N_3450,N_2560,N_2770);
nor U3451 (N_3451,N_2054,N_2892);
or U3452 (N_3452,N_2872,N_2373);
and U3453 (N_3453,N_2848,N_2991);
or U3454 (N_3454,N_2393,N_2958);
nand U3455 (N_3455,N_2179,N_2990);
or U3456 (N_3456,N_2554,N_2540);
or U3457 (N_3457,N_2234,N_2995);
and U3458 (N_3458,N_2662,N_2903);
nand U3459 (N_3459,N_2371,N_2815);
and U3460 (N_3460,N_2797,N_2731);
xor U3461 (N_3461,N_2746,N_2322);
or U3462 (N_3462,N_2093,N_2763);
nor U3463 (N_3463,N_2090,N_2578);
nand U3464 (N_3464,N_2834,N_2704);
and U3465 (N_3465,N_2715,N_2455);
nor U3466 (N_3466,N_2067,N_2461);
and U3467 (N_3467,N_2159,N_2817);
or U3468 (N_3468,N_2716,N_2967);
nor U3469 (N_3469,N_2828,N_2121);
and U3470 (N_3470,N_2686,N_2177);
nand U3471 (N_3471,N_2204,N_2069);
nor U3472 (N_3472,N_2598,N_2862);
nand U3473 (N_3473,N_2241,N_2747);
and U3474 (N_3474,N_2661,N_2109);
xnor U3475 (N_3475,N_2150,N_2262);
and U3476 (N_3476,N_2212,N_2688);
nor U3477 (N_3477,N_2684,N_2787);
xor U3478 (N_3478,N_2802,N_2218);
or U3479 (N_3479,N_2163,N_2435);
nand U3480 (N_3480,N_2957,N_2368);
nand U3481 (N_3481,N_2670,N_2412);
nand U3482 (N_3482,N_2220,N_2604);
nand U3483 (N_3483,N_2840,N_2255);
and U3484 (N_3484,N_2083,N_2210);
nand U3485 (N_3485,N_2375,N_2634);
and U3486 (N_3486,N_2004,N_2063);
nand U3487 (N_3487,N_2749,N_2823);
or U3488 (N_3488,N_2590,N_2884);
nor U3489 (N_3489,N_2551,N_2292);
nor U3490 (N_3490,N_2683,N_2690);
and U3491 (N_3491,N_2423,N_2408);
nand U3492 (N_3492,N_2714,N_2355);
and U3493 (N_3493,N_2384,N_2988);
or U3494 (N_3494,N_2362,N_2667);
or U3495 (N_3495,N_2073,N_2623);
and U3496 (N_3496,N_2058,N_2916);
and U3497 (N_3497,N_2387,N_2782);
nand U3498 (N_3498,N_2586,N_2462);
nor U3499 (N_3499,N_2176,N_2168);
nand U3500 (N_3500,N_2607,N_2657);
nor U3501 (N_3501,N_2899,N_2348);
nor U3502 (N_3502,N_2762,N_2102);
nand U3503 (N_3503,N_2249,N_2624);
and U3504 (N_3504,N_2111,N_2696);
nand U3505 (N_3505,N_2674,N_2434);
xnor U3506 (N_3506,N_2748,N_2435);
or U3507 (N_3507,N_2885,N_2853);
nor U3508 (N_3508,N_2436,N_2144);
nand U3509 (N_3509,N_2410,N_2901);
and U3510 (N_3510,N_2737,N_2373);
xor U3511 (N_3511,N_2246,N_2138);
and U3512 (N_3512,N_2865,N_2150);
or U3513 (N_3513,N_2278,N_2735);
nand U3514 (N_3514,N_2311,N_2587);
and U3515 (N_3515,N_2569,N_2502);
nand U3516 (N_3516,N_2510,N_2899);
or U3517 (N_3517,N_2133,N_2514);
xnor U3518 (N_3518,N_2809,N_2400);
and U3519 (N_3519,N_2496,N_2244);
xnor U3520 (N_3520,N_2865,N_2700);
xor U3521 (N_3521,N_2795,N_2611);
and U3522 (N_3522,N_2781,N_2879);
nand U3523 (N_3523,N_2304,N_2214);
xnor U3524 (N_3524,N_2707,N_2606);
or U3525 (N_3525,N_2642,N_2862);
and U3526 (N_3526,N_2003,N_2747);
and U3527 (N_3527,N_2976,N_2537);
xor U3528 (N_3528,N_2736,N_2938);
or U3529 (N_3529,N_2570,N_2480);
nor U3530 (N_3530,N_2527,N_2522);
nor U3531 (N_3531,N_2823,N_2760);
xnor U3532 (N_3532,N_2821,N_2999);
nand U3533 (N_3533,N_2302,N_2151);
nor U3534 (N_3534,N_2735,N_2763);
or U3535 (N_3535,N_2735,N_2217);
and U3536 (N_3536,N_2336,N_2508);
and U3537 (N_3537,N_2506,N_2402);
nand U3538 (N_3538,N_2929,N_2524);
or U3539 (N_3539,N_2619,N_2640);
and U3540 (N_3540,N_2344,N_2377);
and U3541 (N_3541,N_2214,N_2828);
nand U3542 (N_3542,N_2390,N_2063);
nor U3543 (N_3543,N_2262,N_2325);
and U3544 (N_3544,N_2249,N_2270);
or U3545 (N_3545,N_2980,N_2929);
nand U3546 (N_3546,N_2626,N_2359);
xnor U3547 (N_3547,N_2671,N_2279);
xnor U3548 (N_3548,N_2684,N_2566);
nor U3549 (N_3549,N_2053,N_2023);
or U3550 (N_3550,N_2362,N_2843);
nor U3551 (N_3551,N_2116,N_2342);
or U3552 (N_3552,N_2037,N_2779);
nor U3553 (N_3553,N_2310,N_2313);
xnor U3554 (N_3554,N_2094,N_2434);
and U3555 (N_3555,N_2477,N_2078);
or U3556 (N_3556,N_2320,N_2008);
nor U3557 (N_3557,N_2189,N_2775);
nand U3558 (N_3558,N_2821,N_2170);
nand U3559 (N_3559,N_2273,N_2976);
or U3560 (N_3560,N_2212,N_2281);
xnor U3561 (N_3561,N_2805,N_2171);
and U3562 (N_3562,N_2324,N_2472);
and U3563 (N_3563,N_2265,N_2943);
and U3564 (N_3564,N_2175,N_2627);
or U3565 (N_3565,N_2775,N_2535);
or U3566 (N_3566,N_2370,N_2399);
and U3567 (N_3567,N_2773,N_2355);
nand U3568 (N_3568,N_2905,N_2240);
or U3569 (N_3569,N_2010,N_2114);
and U3570 (N_3570,N_2541,N_2492);
nand U3571 (N_3571,N_2877,N_2080);
nor U3572 (N_3572,N_2626,N_2341);
or U3573 (N_3573,N_2182,N_2086);
nand U3574 (N_3574,N_2624,N_2453);
and U3575 (N_3575,N_2540,N_2927);
or U3576 (N_3576,N_2817,N_2363);
and U3577 (N_3577,N_2013,N_2051);
or U3578 (N_3578,N_2829,N_2329);
and U3579 (N_3579,N_2123,N_2147);
nand U3580 (N_3580,N_2342,N_2899);
xor U3581 (N_3581,N_2472,N_2868);
nor U3582 (N_3582,N_2081,N_2331);
or U3583 (N_3583,N_2895,N_2332);
nand U3584 (N_3584,N_2503,N_2854);
and U3585 (N_3585,N_2754,N_2189);
xnor U3586 (N_3586,N_2688,N_2980);
or U3587 (N_3587,N_2996,N_2230);
xor U3588 (N_3588,N_2970,N_2596);
nand U3589 (N_3589,N_2363,N_2879);
and U3590 (N_3590,N_2582,N_2552);
and U3591 (N_3591,N_2591,N_2275);
or U3592 (N_3592,N_2351,N_2502);
and U3593 (N_3593,N_2927,N_2130);
or U3594 (N_3594,N_2748,N_2541);
and U3595 (N_3595,N_2741,N_2813);
nor U3596 (N_3596,N_2148,N_2099);
and U3597 (N_3597,N_2940,N_2504);
nor U3598 (N_3598,N_2384,N_2100);
and U3599 (N_3599,N_2655,N_2581);
and U3600 (N_3600,N_2956,N_2226);
and U3601 (N_3601,N_2544,N_2413);
and U3602 (N_3602,N_2607,N_2955);
xnor U3603 (N_3603,N_2417,N_2442);
or U3604 (N_3604,N_2954,N_2649);
or U3605 (N_3605,N_2568,N_2972);
nand U3606 (N_3606,N_2155,N_2663);
xnor U3607 (N_3607,N_2212,N_2980);
or U3608 (N_3608,N_2324,N_2576);
nor U3609 (N_3609,N_2332,N_2811);
xnor U3610 (N_3610,N_2798,N_2591);
nand U3611 (N_3611,N_2140,N_2856);
or U3612 (N_3612,N_2774,N_2077);
xor U3613 (N_3613,N_2156,N_2451);
or U3614 (N_3614,N_2596,N_2775);
nand U3615 (N_3615,N_2391,N_2717);
or U3616 (N_3616,N_2730,N_2721);
nor U3617 (N_3617,N_2825,N_2394);
nand U3618 (N_3618,N_2301,N_2327);
nand U3619 (N_3619,N_2132,N_2799);
and U3620 (N_3620,N_2102,N_2786);
and U3621 (N_3621,N_2945,N_2400);
and U3622 (N_3622,N_2436,N_2161);
nor U3623 (N_3623,N_2577,N_2657);
nand U3624 (N_3624,N_2359,N_2286);
xor U3625 (N_3625,N_2992,N_2893);
and U3626 (N_3626,N_2607,N_2833);
nor U3627 (N_3627,N_2623,N_2218);
and U3628 (N_3628,N_2335,N_2728);
or U3629 (N_3629,N_2734,N_2915);
nor U3630 (N_3630,N_2016,N_2609);
and U3631 (N_3631,N_2936,N_2900);
and U3632 (N_3632,N_2718,N_2606);
nor U3633 (N_3633,N_2780,N_2195);
and U3634 (N_3634,N_2590,N_2307);
nand U3635 (N_3635,N_2217,N_2159);
and U3636 (N_3636,N_2420,N_2402);
nor U3637 (N_3637,N_2757,N_2284);
or U3638 (N_3638,N_2361,N_2447);
and U3639 (N_3639,N_2107,N_2058);
or U3640 (N_3640,N_2288,N_2528);
nand U3641 (N_3641,N_2953,N_2862);
and U3642 (N_3642,N_2927,N_2442);
and U3643 (N_3643,N_2374,N_2475);
nand U3644 (N_3644,N_2604,N_2031);
nor U3645 (N_3645,N_2966,N_2980);
and U3646 (N_3646,N_2176,N_2608);
or U3647 (N_3647,N_2892,N_2086);
nor U3648 (N_3648,N_2042,N_2408);
nand U3649 (N_3649,N_2169,N_2869);
nand U3650 (N_3650,N_2867,N_2950);
xor U3651 (N_3651,N_2037,N_2409);
nand U3652 (N_3652,N_2575,N_2610);
or U3653 (N_3653,N_2555,N_2999);
and U3654 (N_3654,N_2764,N_2430);
xnor U3655 (N_3655,N_2325,N_2724);
and U3656 (N_3656,N_2317,N_2449);
xnor U3657 (N_3657,N_2444,N_2320);
nand U3658 (N_3658,N_2490,N_2410);
or U3659 (N_3659,N_2070,N_2160);
or U3660 (N_3660,N_2018,N_2107);
and U3661 (N_3661,N_2873,N_2809);
and U3662 (N_3662,N_2741,N_2355);
xor U3663 (N_3663,N_2618,N_2814);
nor U3664 (N_3664,N_2619,N_2905);
nand U3665 (N_3665,N_2435,N_2235);
nand U3666 (N_3666,N_2100,N_2952);
and U3667 (N_3667,N_2251,N_2442);
nand U3668 (N_3668,N_2055,N_2348);
nor U3669 (N_3669,N_2411,N_2963);
xor U3670 (N_3670,N_2901,N_2969);
or U3671 (N_3671,N_2917,N_2374);
xnor U3672 (N_3672,N_2801,N_2282);
nor U3673 (N_3673,N_2887,N_2722);
nor U3674 (N_3674,N_2304,N_2425);
nor U3675 (N_3675,N_2977,N_2735);
or U3676 (N_3676,N_2213,N_2523);
and U3677 (N_3677,N_2985,N_2619);
or U3678 (N_3678,N_2699,N_2740);
nor U3679 (N_3679,N_2004,N_2937);
nor U3680 (N_3680,N_2129,N_2014);
nand U3681 (N_3681,N_2322,N_2953);
xor U3682 (N_3682,N_2065,N_2993);
nor U3683 (N_3683,N_2015,N_2633);
nand U3684 (N_3684,N_2758,N_2726);
xor U3685 (N_3685,N_2830,N_2714);
xnor U3686 (N_3686,N_2920,N_2225);
nand U3687 (N_3687,N_2927,N_2431);
or U3688 (N_3688,N_2450,N_2677);
xnor U3689 (N_3689,N_2691,N_2229);
nor U3690 (N_3690,N_2923,N_2655);
nor U3691 (N_3691,N_2682,N_2639);
nand U3692 (N_3692,N_2015,N_2332);
xor U3693 (N_3693,N_2683,N_2085);
nand U3694 (N_3694,N_2588,N_2651);
or U3695 (N_3695,N_2142,N_2310);
nor U3696 (N_3696,N_2433,N_2424);
nand U3697 (N_3697,N_2444,N_2673);
xor U3698 (N_3698,N_2496,N_2160);
nand U3699 (N_3699,N_2281,N_2992);
nor U3700 (N_3700,N_2823,N_2104);
and U3701 (N_3701,N_2367,N_2253);
nor U3702 (N_3702,N_2312,N_2515);
xnor U3703 (N_3703,N_2267,N_2643);
or U3704 (N_3704,N_2010,N_2432);
nor U3705 (N_3705,N_2320,N_2254);
nand U3706 (N_3706,N_2837,N_2570);
or U3707 (N_3707,N_2465,N_2194);
nor U3708 (N_3708,N_2697,N_2274);
xor U3709 (N_3709,N_2554,N_2545);
nor U3710 (N_3710,N_2478,N_2398);
nand U3711 (N_3711,N_2075,N_2107);
nor U3712 (N_3712,N_2097,N_2713);
and U3713 (N_3713,N_2730,N_2193);
and U3714 (N_3714,N_2856,N_2696);
nor U3715 (N_3715,N_2895,N_2208);
and U3716 (N_3716,N_2002,N_2705);
and U3717 (N_3717,N_2086,N_2256);
nand U3718 (N_3718,N_2762,N_2673);
nand U3719 (N_3719,N_2429,N_2158);
or U3720 (N_3720,N_2810,N_2133);
or U3721 (N_3721,N_2095,N_2569);
nand U3722 (N_3722,N_2463,N_2267);
or U3723 (N_3723,N_2957,N_2589);
nand U3724 (N_3724,N_2028,N_2180);
nor U3725 (N_3725,N_2755,N_2711);
and U3726 (N_3726,N_2938,N_2303);
nand U3727 (N_3727,N_2666,N_2607);
nor U3728 (N_3728,N_2312,N_2215);
xnor U3729 (N_3729,N_2144,N_2485);
or U3730 (N_3730,N_2465,N_2778);
or U3731 (N_3731,N_2623,N_2291);
xor U3732 (N_3732,N_2749,N_2860);
and U3733 (N_3733,N_2857,N_2265);
or U3734 (N_3734,N_2106,N_2776);
or U3735 (N_3735,N_2739,N_2111);
and U3736 (N_3736,N_2244,N_2749);
and U3737 (N_3737,N_2682,N_2865);
nand U3738 (N_3738,N_2195,N_2366);
or U3739 (N_3739,N_2668,N_2334);
or U3740 (N_3740,N_2630,N_2752);
xnor U3741 (N_3741,N_2125,N_2046);
and U3742 (N_3742,N_2657,N_2323);
nor U3743 (N_3743,N_2694,N_2900);
and U3744 (N_3744,N_2830,N_2083);
xor U3745 (N_3745,N_2023,N_2890);
or U3746 (N_3746,N_2250,N_2797);
xor U3747 (N_3747,N_2349,N_2756);
xnor U3748 (N_3748,N_2835,N_2343);
and U3749 (N_3749,N_2444,N_2931);
xnor U3750 (N_3750,N_2426,N_2701);
and U3751 (N_3751,N_2673,N_2747);
or U3752 (N_3752,N_2153,N_2711);
nand U3753 (N_3753,N_2131,N_2874);
xor U3754 (N_3754,N_2006,N_2040);
or U3755 (N_3755,N_2018,N_2000);
xnor U3756 (N_3756,N_2036,N_2792);
xor U3757 (N_3757,N_2267,N_2665);
xor U3758 (N_3758,N_2531,N_2030);
nand U3759 (N_3759,N_2176,N_2528);
and U3760 (N_3760,N_2716,N_2423);
nand U3761 (N_3761,N_2431,N_2985);
xor U3762 (N_3762,N_2318,N_2189);
or U3763 (N_3763,N_2189,N_2869);
nand U3764 (N_3764,N_2772,N_2077);
and U3765 (N_3765,N_2778,N_2820);
xor U3766 (N_3766,N_2334,N_2292);
nor U3767 (N_3767,N_2895,N_2619);
xnor U3768 (N_3768,N_2109,N_2320);
and U3769 (N_3769,N_2930,N_2901);
and U3770 (N_3770,N_2961,N_2730);
nand U3771 (N_3771,N_2128,N_2285);
and U3772 (N_3772,N_2211,N_2397);
xnor U3773 (N_3773,N_2012,N_2909);
xor U3774 (N_3774,N_2826,N_2657);
or U3775 (N_3775,N_2860,N_2611);
xnor U3776 (N_3776,N_2721,N_2589);
or U3777 (N_3777,N_2391,N_2958);
xnor U3778 (N_3778,N_2660,N_2554);
or U3779 (N_3779,N_2343,N_2083);
xnor U3780 (N_3780,N_2491,N_2636);
and U3781 (N_3781,N_2471,N_2747);
or U3782 (N_3782,N_2720,N_2153);
nor U3783 (N_3783,N_2186,N_2626);
xor U3784 (N_3784,N_2510,N_2654);
nand U3785 (N_3785,N_2450,N_2543);
and U3786 (N_3786,N_2597,N_2798);
nand U3787 (N_3787,N_2328,N_2887);
xnor U3788 (N_3788,N_2316,N_2329);
xnor U3789 (N_3789,N_2516,N_2715);
xnor U3790 (N_3790,N_2014,N_2158);
nand U3791 (N_3791,N_2403,N_2754);
nor U3792 (N_3792,N_2808,N_2174);
xnor U3793 (N_3793,N_2986,N_2384);
xnor U3794 (N_3794,N_2023,N_2060);
or U3795 (N_3795,N_2060,N_2624);
nand U3796 (N_3796,N_2117,N_2495);
xor U3797 (N_3797,N_2645,N_2283);
xor U3798 (N_3798,N_2898,N_2106);
or U3799 (N_3799,N_2598,N_2079);
xor U3800 (N_3800,N_2989,N_2634);
or U3801 (N_3801,N_2972,N_2322);
nor U3802 (N_3802,N_2939,N_2675);
nand U3803 (N_3803,N_2718,N_2342);
xnor U3804 (N_3804,N_2861,N_2686);
and U3805 (N_3805,N_2461,N_2317);
xnor U3806 (N_3806,N_2469,N_2826);
or U3807 (N_3807,N_2374,N_2550);
nor U3808 (N_3808,N_2474,N_2583);
and U3809 (N_3809,N_2165,N_2536);
and U3810 (N_3810,N_2665,N_2125);
nand U3811 (N_3811,N_2811,N_2177);
nand U3812 (N_3812,N_2728,N_2030);
or U3813 (N_3813,N_2695,N_2324);
xnor U3814 (N_3814,N_2449,N_2528);
nor U3815 (N_3815,N_2362,N_2280);
or U3816 (N_3816,N_2751,N_2734);
and U3817 (N_3817,N_2062,N_2293);
and U3818 (N_3818,N_2088,N_2601);
or U3819 (N_3819,N_2323,N_2257);
nor U3820 (N_3820,N_2383,N_2432);
xor U3821 (N_3821,N_2145,N_2087);
nand U3822 (N_3822,N_2228,N_2478);
or U3823 (N_3823,N_2036,N_2576);
xnor U3824 (N_3824,N_2677,N_2915);
nor U3825 (N_3825,N_2847,N_2610);
nor U3826 (N_3826,N_2068,N_2320);
nor U3827 (N_3827,N_2052,N_2828);
xnor U3828 (N_3828,N_2554,N_2736);
nor U3829 (N_3829,N_2077,N_2092);
or U3830 (N_3830,N_2716,N_2410);
nor U3831 (N_3831,N_2254,N_2515);
xnor U3832 (N_3832,N_2738,N_2353);
and U3833 (N_3833,N_2471,N_2792);
and U3834 (N_3834,N_2001,N_2730);
xnor U3835 (N_3835,N_2707,N_2098);
nor U3836 (N_3836,N_2009,N_2598);
nor U3837 (N_3837,N_2451,N_2953);
xnor U3838 (N_3838,N_2594,N_2104);
xnor U3839 (N_3839,N_2782,N_2228);
nand U3840 (N_3840,N_2022,N_2355);
nand U3841 (N_3841,N_2268,N_2948);
nor U3842 (N_3842,N_2850,N_2574);
xnor U3843 (N_3843,N_2242,N_2181);
nor U3844 (N_3844,N_2292,N_2688);
nand U3845 (N_3845,N_2440,N_2176);
nand U3846 (N_3846,N_2232,N_2246);
xnor U3847 (N_3847,N_2036,N_2276);
nand U3848 (N_3848,N_2827,N_2562);
or U3849 (N_3849,N_2593,N_2087);
nor U3850 (N_3850,N_2526,N_2643);
and U3851 (N_3851,N_2978,N_2764);
nor U3852 (N_3852,N_2253,N_2049);
and U3853 (N_3853,N_2832,N_2999);
nor U3854 (N_3854,N_2313,N_2233);
and U3855 (N_3855,N_2626,N_2207);
and U3856 (N_3856,N_2666,N_2274);
and U3857 (N_3857,N_2727,N_2396);
xnor U3858 (N_3858,N_2324,N_2105);
nand U3859 (N_3859,N_2882,N_2405);
or U3860 (N_3860,N_2835,N_2762);
nand U3861 (N_3861,N_2632,N_2500);
nand U3862 (N_3862,N_2953,N_2745);
xor U3863 (N_3863,N_2902,N_2986);
nand U3864 (N_3864,N_2961,N_2855);
nand U3865 (N_3865,N_2392,N_2236);
xnor U3866 (N_3866,N_2367,N_2879);
nor U3867 (N_3867,N_2090,N_2595);
and U3868 (N_3868,N_2299,N_2692);
nand U3869 (N_3869,N_2817,N_2970);
or U3870 (N_3870,N_2388,N_2309);
and U3871 (N_3871,N_2741,N_2801);
or U3872 (N_3872,N_2220,N_2122);
nand U3873 (N_3873,N_2045,N_2110);
xnor U3874 (N_3874,N_2012,N_2791);
and U3875 (N_3875,N_2262,N_2290);
nand U3876 (N_3876,N_2080,N_2374);
nor U3877 (N_3877,N_2152,N_2543);
nand U3878 (N_3878,N_2410,N_2872);
xor U3879 (N_3879,N_2785,N_2332);
nor U3880 (N_3880,N_2282,N_2455);
and U3881 (N_3881,N_2160,N_2058);
nor U3882 (N_3882,N_2899,N_2993);
nor U3883 (N_3883,N_2655,N_2806);
xor U3884 (N_3884,N_2020,N_2141);
nand U3885 (N_3885,N_2196,N_2544);
nand U3886 (N_3886,N_2475,N_2880);
nor U3887 (N_3887,N_2314,N_2358);
nor U3888 (N_3888,N_2750,N_2232);
nand U3889 (N_3889,N_2987,N_2354);
or U3890 (N_3890,N_2609,N_2041);
or U3891 (N_3891,N_2087,N_2692);
nand U3892 (N_3892,N_2836,N_2847);
and U3893 (N_3893,N_2371,N_2293);
and U3894 (N_3894,N_2613,N_2757);
nor U3895 (N_3895,N_2482,N_2586);
or U3896 (N_3896,N_2108,N_2962);
xnor U3897 (N_3897,N_2508,N_2120);
xnor U3898 (N_3898,N_2771,N_2384);
or U3899 (N_3899,N_2099,N_2132);
nor U3900 (N_3900,N_2891,N_2511);
or U3901 (N_3901,N_2860,N_2926);
nor U3902 (N_3902,N_2888,N_2660);
nor U3903 (N_3903,N_2324,N_2997);
and U3904 (N_3904,N_2288,N_2664);
nand U3905 (N_3905,N_2181,N_2280);
xnor U3906 (N_3906,N_2640,N_2139);
and U3907 (N_3907,N_2600,N_2830);
xor U3908 (N_3908,N_2207,N_2362);
and U3909 (N_3909,N_2929,N_2052);
nor U3910 (N_3910,N_2234,N_2339);
xor U3911 (N_3911,N_2289,N_2470);
xor U3912 (N_3912,N_2228,N_2373);
nor U3913 (N_3913,N_2690,N_2313);
and U3914 (N_3914,N_2046,N_2059);
or U3915 (N_3915,N_2502,N_2833);
nor U3916 (N_3916,N_2863,N_2909);
xor U3917 (N_3917,N_2418,N_2778);
nand U3918 (N_3918,N_2294,N_2552);
or U3919 (N_3919,N_2026,N_2653);
and U3920 (N_3920,N_2057,N_2875);
xnor U3921 (N_3921,N_2873,N_2606);
xnor U3922 (N_3922,N_2912,N_2330);
nor U3923 (N_3923,N_2276,N_2040);
nand U3924 (N_3924,N_2232,N_2553);
and U3925 (N_3925,N_2487,N_2536);
or U3926 (N_3926,N_2690,N_2804);
or U3927 (N_3927,N_2524,N_2347);
xnor U3928 (N_3928,N_2795,N_2178);
or U3929 (N_3929,N_2913,N_2895);
or U3930 (N_3930,N_2486,N_2000);
xnor U3931 (N_3931,N_2459,N_2650);
xnor U3932 (N_3932,N_2051,N_2795);
or U3933 (N_3933,N_2802,N_2144);
or U3934 (N_3934,N_2099,N_2691);
nand U3935 (N_3935,N_2990,N_2942);
nor U3936 (N_3936,N_2223,N_2147);
and U3937 (N_3937,N_2427,N_2103);
nor U3938 (N_3938,N_2541,N_2081);
and U3939 (N_3939,N_2104,N_2793);
nand U3940 (N_3940,N_2156,N_2989);
nor U3941 (N_3941,N_2880,N_2274);
or U3942 (N_3942,N_2029,N_2803);
or U3943 (N_3943,N_2931,N_2402);
and U3944 (N_3944,N_2818,N_2379);
nand U3945 (N_3945,N_2517,N_2625);
nand U3946 (N_3946,N_2932,N_2675);
nand U3947 (N_3947,N_2177,N_2774);
nand U3948 (N_3948,N_2975,N_2412);
nand U3949 (N_3949,N_2147,N_2600);
nand U3950 (N_3950,N_2090,N_2113);
and U3951 (N_3951,N_2758,N_2713);
nor U3952 (N_3952,N_2932,N_2996);
nor U3953 (N_3953,N_2361,N_2325);
xnor U3954 (N_3954,N_2741,N_2420);
nor U3955 (N_3955,N_2900,N_2636);
nand U3956 (N_3956,N_2883,N_2922);
or U3957 (N_3957,N_2148,N_2604);
xor U3958 (N_3958,N_2661,N_2972);
or U3959 (N_3959,N_2687,N_2078);
nor U3960 (N_3960,N_2585,N_2462);
or U3961 (N_3961,N_2330,N_2960);
and U3962 (N_3962,N_2970,N_2043);
xnor U3963 (N_3963,N_2627,N_2829);
and U3964 (N_3964,N_2768,N_2606);
xnor U3965 (N_3965,N_2803,N_2054);
nand U3966 (N_3966,N_2829,N_2387);
or U3967 (N_3967,N_2737,N_2708);
nor U3968 (N_3968,N_2973,N_2269);
xnor U3969 (N_3969,N_2763,N_2912);
nor U3970 (N_3970,N_2595,N_2883);
and U3971 (N_3971,N_2206,N_2510);
or U3972 (N_3972,N_2614,N_2127);
and U3973 (N_3973,N_2910,N_2712);
nor U3974 (N_3974,N_2763,N_2677);
xor U3975 (N_3975,N_2956,N_2954);
nand U3976 (N_3976,N_2902,N_2278);
nand U3977 (N_3977,N_2319,N_2181);
nor U3978 (N_3978,N_2996,N_2386);
nand U3979 (N_3979,N_2880,N_2843);
xor U3980 (N_3980,N_2963,N_2425);
and U3981 (N_3981,N_2623,N_2062);
nand U3982 (N_3982,N_2822,N_2742);
xor U3983 (N_3983,N_2431,N_2298);
nor U3984 (N_3984,N_2105,N_2259);
nand U3985 (N_3985,N_2465,N_2222);
or U3986 (N_3986,N_2924,N_2732);
and U3987 (N_3987,N_2180,N_2834);
or U3988 (N_3988,N_2734,N_2266);
nand U3989 (N_3989,N_2902,N_2469);
nor U3990 (N_3990,N_2698,N_2111);
xnor U3991 (N_3991,N_2197,N_2573);
and U3992 (N_3992,N_2488,N_2984);
nand U3993 (N_3993,N_2220,N_2019);
and U3994 (N_3994,N_2473,N_2981);
xnor U3995 (N_3995,N_2007,N_2122);
nor U3996 (N_3996,N_2379,N_2233);
nor U3997 (N_3997,N_2567,N_2357);
and U3998 (N_3998,N_2075,N_2884);
nand U3999 (N_3999,N_2734,N_2168);
xnor U4000 (N_4000,N_3088,N_3113);
and U4001 (N_4001,N_3900,N_3241);
nand U4002 (N_4002,N_3595,N_3896);
nand U4003 (N_4003,N_3265,N_3050);
or U4004 (N_4004,N_3234,N_3583);
or U4005 (N_4005,N_3806,N_3476);
and U4006 (N_4006,N_3567,N_3540);
or U4007 (N_4007,N_3230,N_3755);
nand U4008 (N_4008,N_3040,N_3168);
nor U4009 (N_4009,N_3329,N_3115);
or U4010 (N_4010,N_3042,N_3535);
or U4011 (N_4011,N_3193,N_3488);
nand U4012 (N_4012,N_3859,N_3381);
nand U4013 (N_4013,N_3988,N_3290);
xnor U4014 (N_4014,N_3256,N_3940);
or U4015 (N_4015,N_3893,N_3098);
xnor U4016 (N_4016,N_3428,N_3450);
and U4017 (N_4017,N_3471,N_3282);
nor U4018 (N_4018,N_3120,N_3456);
nor U4019 (N_4019,N_3196,N_3674);
and U4020 (N_4020,N_3106,N_3031);
nand U4021 (N_4021,N_3043,N_3739);
nor U4022 (N_4022,N_3372,N_3746);
xnor U4023 (N_4023,N_3716,N_3506);
nor U4024 (N_4024,N_3610,N_3200);
nand U4025 (N_4025,N_3046,N_3968);
and U4026 (N_4026,N_3872,N_3284);
and U4027 (N_4027,N_3552,N_3620);
nor U4028 (N_4028,N_3886,N_3976);
and U4029 (N_4029,N_3248,N_3820);
or U4030 (N_4030,N_3192,N_3667);
nor U4031 (N_4031,N_3159,N_3440);
and U4032 (N_4032,N_3487,N_3484);
xnor U4033 (N_4033,N_3842,N_3005);
xor U4034 (N_4034,N_3094,N_3796);
and U4035 (N_4035,N_3383,N_3330);
xnor U4036 (N_4036,N_3603,N_3235);
nand U4037 (N_4037,N_3604,N_3978);
xnor U4038 (N_4038,N_3062,N_3399);
nand U4039 (N_4039,N_3589,N_3435);
or U4040 (N_4040,N_3298,N_3243);
nor U4041 (N_4041,N_3108,N_3026);
or U4042 (N_4042,N_3994,N_3149);
xnor U4043 (N_4043,N_3948,N_3029);
or U4044 (N_4044,N_3051,N_3384);
nor U4045 (N_4045,N_3002,N_3360);
nor U4046 (N_4046,N_3732,N_3331);
or U4047 (N_4047,N_3786,N_3371);
nor U4048 (N_4048,N_3854,N_3165);
and U4049 (N_4049,N_3414,N_3791);
and U4050 (N_4050,N_3466,N_3780);
and U4051 (N_4051,N_3255,N_3459);
xnor U4052 (N_4052,N_3016,N_3673);
and U4053 (N_4053,N_3364,N_3368);
or U4054 (N_4054,N_3246,N_3028);
and U4055 (N_4055,N_3418,N_3267);
nand U4056 (N_4056,N_3578,N_3299);
and U4057 (N_4057,N_3332,N_3410);
or U4058 (N_4058,N_3056,N_3308);
xnor U4059 (N_4059,N_3542,N_3928);
or U4060 (N_4060,N_3180,N_3478);
nand U4061 (N_4061,N_3217,N_3382);
or U4062 (N_4062,N_3742,N_3228);
nor U4063 (N_4063,N_3153,N_3346);
xnor U4064 (N_4064,N_3812,N_3519);
xnor U4065 (N_4065,N_3628,N_3075);
xnor U4066 (N_4066,N_3293,N_3232);
or U4067 (N_4067,N_3751,N_3426);
nor U4068 (N_4068,N_3808,N_3609);
and U4069 (N_4069,N_3563,N_3491);
and U4070 (N_4070,N_3635,N_3183);
nand U4071 (N_4071,N_3433,N_3670);
xor U4072 (N_4072,N_3825,N_3336);
nand U4073 (N_4073,N_3866,N_3084);
nor U4074 (N_4074,N_3137,N_3104);
xnor U4075 (N_4075,N_3935,N_3145);
or U4076 (N_4076,N_3672,N_3849);
and U4077 (N_4077,N_3760,N_3434);
or U4078 (N_4078,N_3320,N_3961);
and U4079 (N_4079,N_3807,N_3868);
xor U4080 (N_4080,N_3163,N_3500);
and U4081 (N_4081,N_3348,N_3489);
and U4082 (N_4082,N_3924,N_3733);
xnor U4083 (N_4083,N_3641,N_3162);
nand U4084 (N_4084,N_3878,N_3663);
or U4085 (N_4085,N_3054,N_3593);
and U4086 (N_4086,N_3653,N_3432);
nand U4087 (N_4087,N_3199,N_3444);
or U4088 (N_4088,N_3511,N_3779);
nand U4089 (N_4089,N_3136,N_3592);
and U4090 (N_4090,N_3123,N_3474);
or U4091 (N_4091,N_3438,N_3274);
or U4092 (N_4092,N_3852,N_3768);
nor U4093 (N_4093,N_3985,N_3864);
xor U4094 (N_4094,N_3577,N_3917);
xor U4095 (N_4095,N_3294,N_3020);
and U4096 (N_4096,N_3622,N_3950);
xnor U4097 (N_4097,N_3208,N_3226);
xnor U4098 (N_4098,N_3752,N_3572);
xor U4099 (N_4099,N_3288,N_3262);
and U4100 (N_4100,N_3831,N_3300);
xor U4101 (N_4101,N_3482,N_3549);
nand U4102 (N_4102,N_3377,N_3649);
and U4103 (N_4103,N_3957,N_3130);
and U4104 (N_4104,N_3206,N_3677);
and U4105 (N_4105,N_3212,N_3838);
or U4106 (N_4106,N_3443,N_3380);
nand U4107 (N_4107,N_3470,N_3556);
or U4108 (N_4108,N_3997,N_3057);
xor U4109 (N_4109,N_3337,N_3654);
nor U4110 (N_4110,N_3023,N_3615);
or U4111 (N_4111,N_3581,N_3605);
nor U4112 (N_4112,N_3499,N_3127);
nand U4113 (N_4113,N_3365,N_3087);
nor U4114 (N_4114,N_3458,N_3036);
nor U4115 (N_4115,N_3078,N_3931);
and U4116 (N_4116,N_3638,N_3338);
or U4117 (N_4117,N_3110,N_3204);
nand U4118 (N_4118,N_3770,N_3277);
xor U4119 (N_4119,N_3353,N_3698);
nor U4120 (N_4120,N_3363,N_3264);
nand U4121 (N_4121,N_3452,N_3731);
or U4122 (N_4122,N_3251,N_3824);
or U4123 (N_4123,N_3086,N_3930);
nor U4124 (N_4124,N_3063,N_3323);
and U4125 (N_4125,N_3850,N_3403);
xor U4126 (N_4126,N_3446,N_3469);
or U4127 (N_4127,N_3793,N_3205);
nor U4128 (N_4128,N_3125,N_3409);
nand U4129 (N_4129,N_3652,N_3743);
nand U4130 (N_4130,N_3555,N_3766);
and U4131 (N_4131,N_3269,N_3468);
and U4132 (N_4132,N_3493,N_3547);
and U4133 (N_4133,N_3520,N_3981);
or U4134 (N_4134,N_3953,N_3013);
nand U4135 (N_4135,N_3613,N_3802);
xnor U4136 (N_4136,N_3441,N_3437);
nand U4137 (N_4137,N_3625,N_3436);
nand U4138 (N_4138,N_3310,N_3503);
or U4139 (N_4139,N_3415,N_3883);
nor U4140 (N_4140,N_3929,N_3092);
or U4141 (N_4141,N_3461,N_3322);
and U4142 (N_4142,N_3958,N_3970);
and U4143 (N_4143,N_3987,N_3447);
and U4144 (N_4144,N_3210,N_3637);
and U4145 (N_4145,N_3758,N_3140);
xnor U4146 (N_4146,N_3767,N_3933);
xnor U4147 (N_4147,N_3512,N_3903);
nand U4148 (N_4148,N_3753,N_3498);
or U4149 (N_4149,N_3376,N_3799);
or U4150 (N_4150,N_3216,N_3128);
or U4151 (N_4151,N_3618,N_3782);
nand U4152 (N_4152,N_3501,N_3533);
xnor U4153 (N_4153,N_3263,N_3867);
and U4154 (N_4154,N_3964,N_3923);
xor U4155 (N_4155,N_3892,N_3223);
and U4156 (N_4156,N_3211,N_3669);
or U4157 (N_4157,N_3366,N_3938);
nor U4158 (N_4158,N_3502,N_3295);
nor U4159 (N_4159,N_3354,N_3551);
and U4160 (N_4160,N_3642,N_3664);
nor U4161 (N_4161,N_3811,N_3693);
and U4162 (N_4162,N_3843,N_3774);
xnor U4163 (N_4163,N_3147,N_3144);
nor U4164 (N_4164,N_3352,N_3229);
nand U4165 (N_4165,N_3496,N_3068);
and U4166 (N_4166,N_3829,N_3202);
and U4167 (N_4167,N_3719,N_3008);
nand U4168 (N_4168,N_3562,N_3992);
or U4169 (N_4169,N_3252,N_3772);
or U4170 (N_4170,N_3207,N_3853);
and U4171 (N_4171,N_3021,N_3738);
and U4172 (N_4172,N_3543,N_3579);
or U4173 (N_4173,N_3754,N_3907);
nand U4174 (N_4174,N_3465,N_3334);
xor U4175 (N_4175,N_3534,N_3550);
nand U4176 (N_4176,N_3764,N_3836);
nand U4177 (N_4177,N_3761,N_3236);
xnor U4178 (N_4178,N_3497,N_3848);
or U4179 (N_4179,N_3333,N_3946);
and U4180 (N_4180,N_3715,N_3397);
xor U4181 (N_4181,N_3213,N_3630);
and U4182 (N_4182,N_3973,N_3982);
nand U4183 (N_4183,N_3600,N_3906);
or U4184 (N_4184,N_3061,N_3312);
nor U4185 (N_4185,N_3922,N_3190);
or U4186 (N_4186,N_3387,N_3189);
nor U4187 (N_4187,N_3690,N_3797);
nor U4188 (N_4188,N_3015,N_3851);
and U4189 (N_4189,N_3995,N_3894);
or U4190 (N_4190,N_3845,N_3584);
nand U4191 (N_4191,N_3143,N_3239);
nand U4192 (N_4192,N_3350,N_3072);
or U4193 (N_4193,N_3448,N_3275);
xor U4194 (N_4194,N_3833,N_3166);
xor U4195 (N_4195,N_3794,N_3568);
and U4196 (N_4196,N_3640,N_3627);
nand U4197 (N_4197,N_3671,N_3518);
nor U4198 (N_4198,N_3626,N_3530);
xnor U4199 (N_4199,N_3475,N_3385);
nand U4200 (N_4200,N_3749,N_3773);
nor U4201 (N_4201,N_3517,N_3045);
or U4202 (N_4202,N_3081,N_3430);
and U4203 (N_4203,N_3736,N_3596);
or U4204 (N_4204,N_3951,N_3585);
xor U4205 (N_4205,N_3138,N_3846);
nor U4206 (N_4206,N_3662,N_3035);
nand U4207 (N_4207,N_3188,N_3142);
and U4208 (N_4208,N_3326,N_3058);
xor U4209 (N_4209,N_3943,N_3569);
nor U4210 (N_4210,N_3740,N_3784);
and U4211 (N_4211,N_3184,N_3744);
and U4212 (N_4212,N_3340,N_3717);
nand U4213 (N_4213,N_3522,N_3071);
xor U4214 (N_4214,N_3356,N_3097);
xor U4215 (N_4215,N_3112,N_3510);
nor U4216 (N_4216,N_3913,N_3093);
or U4217 (N_4217,N_3521,N_3473);
nor U4218 (N_4218,N_3492,N_3697);
and U4219 (N_4219,N_3801,N_3965);
and U4220 (N_4220,N_3890,N_3453);
nand U4221 (N_4221,N_3860,N_3704);
xnor U4222 (N_4222,N_3100,N_3271);
nor U4223 (N_4223,N_3575,N_3897);
xor U4224 (N_4224,N_3116,N_3686);
xor U4225 (N_4225,N_3775,N_3374);
nor U4226 (N_4226,N_3823,N_3266);
and U4227 (N_4227,N_3816,N_3813);
and U4228 (N_4228,N_3479,N_3590);
nand U4229 (N_4229,N_3735,N_3911);
xor U4230 (N_4230,N_3616,N_3421);
xnor U4231 (N_4231,N_3546,N_3974);
xor U4232 (N_4232,N_3401,N_3526);
xnor U4233 (N_4233,N_3442,N_3975);
nor U4234 (N_4234,N_3727,N_3185);
xnor U4235 (N_4235,N_3278,N_3598);
nor U4236 (N_4236,N_3395,N_3027);
nand U4237 (N_4237,N_3316,N_3632);
and U4238 (N_4238,N_3971,N_3821);
or U4239 (N_4239,N_3524,N_3073);
nor U4240 (N_4240,N_3012,N_3762);
or U4241 (N_4241,N_3955,N_3827);
xnor U4242 (N_4242,N_3619,N_3194);
nor U4243 (N_4243,N_3857,N_3835);
or U4244 (N_4244,N_3949,N_3601);
xor U4245 (N_4245,N_3963,N_3822);
and U4246 (N_4246,N_3238,N_3203);
xnor U4247 (N_4247,N_3684,N_3999);
or U4248 (N_4248,N_3480,N_3926);
xnor U4249 (N_4249,N_3341,N_3388);
or U4250 (N_4250,N_3879,N_3612);
nor U4251 (N_4251,N_3392,N_3874);
xor U4252 (N_4252,N_3309,N_3621);
xnor U4253 (N_4253,N_3571,N_3699);
nand U4254 (N_4254,N_3695,N_3582);
and U4255 (N_4255,N_3132,N_3010);
nor U4256 (N_4256,N_3431,N_3895);
nand U4257 (N_4257,N_3798,N_3167);
or U4258 (N_4258,N_3483,N_3525);
nand U4259 (N_4259,N_3661,N_3915);
nor U4260 (N_4260,N_3881,N_3862);
nor U4261 (N_4261,N_3317,N_3745);
nor U4262 (N_4262,N_3650,N_3729);
xor U4263 (N_4263,N_3422,N_3398);
or U4264 (N_4264,N_3599,N_3757);
or U4265 (N_4265,N_3841,N_3657);
or U4266 (N_4266,N_3700,N_3614);
xor U4267 (N_4267,N_3391,N_3351);
xnor U4268 (N_4268,N_3541,N_3509);
or U4269 (N_4269,N_3718,N_3665);
and U4270 (N_4270,N_3728,N_3324);
nor U4271 (N_4271,N_3030,N_3722);
nand U4272 (N_4272,N_3573,N_3880);
nor U4273 (N_4273,N_3787,N_3055);
nor U4274 (N_4274,N_3464,N_3462);
nor U4275 (N_4275,N_3747,N_3285);
and U4276 (N_4276,N_3118,N_3396);
or U4277 (N_4277,N_3227,N_3945);
or U4278 (N_4278,N_3668,N_3004);
xnor U4279 (N_4279,N_3545,N_3647);
and U4280 (N_4280,N_3678,N_3925);
xor U4281 (N_4281,N_3701,N_3910);
and U4282 (N_4282,N_3861,N_3400);
nand U4283 (N_4283,N_3457,N_3494);
nand U4284 (N_4284,N_3259,N_3869);
nor U4285 (N_4285,N_3083,N_3289);
and U4286 (N_4286,N_3696,N_3099);
or U4287 (N_4287,N_3721,N_3817);
nor U4288 (N_4288,N_3281,N_3169);
nand U4289 (N_4289,N_3276,N_3810);
nand U4290 (N_4290,N_3844,N_3656);
xor U4291 (N_4291,N_3863,N_3792);
nand U4292 (N_4292,N_3369,N_3122);
or U4293 (N_4293,N_3889,N_3176);
nor U4294 (N_4294,N_3225,N_3709);
nand U4295 (N_4295,N_3785,N_3018);
or U4296 (N_4296,N_3151,N_3565);
and U4297 (N_4297,N_3803,N_3998);
or U4298 (N_4298,N_3339,N_3914);
nor U4299 (N_4299,N_3408,N_3523);
xor U4300 (N_4300,N_3544,N_3685);
xor U4301 (N_4301,N_3150,N_3187);
nand U4302 (N_4302,N_3712,N_3916);
xor U4303 (N_4303,N_3379,N_3032);
or U4304 (N_4304,N_3148,N_3177);
nand U4305 (N_4305,N_3311,N_3074);
nor U4306 (N_4306,N_3920,N_3713);
xor U4307 (N_4307,N_3611,N_3305);
and U4308 (N_4308,N_3066,N_3837);
xor U4309 (N_4309,N_3114,N_3378);
and U4310 (N_4310,N_3195,N_3179);
xnor U4311 (N_4311,N_3576,N_3367);
or U4312 (N_4312,N_3539,N_3318);
nor U4313 (N_4313,N_3633,N_3531);
nor U4314 (N_4314,N_3485,N_3080);
nor U4315 (N_4315,N_3319,N_3706);
nor U4316 (N_4316,N_3557,N_3887);
and U4317 (N_4317,N_3901,N_3847);
nand U4318 (N_4318,N_3591,N_3876);
xor U4319 (N_4319,N_3375,N_3636);
xor U4320 (N_4320,N_3313,N_3904);
and U4321 (N_4321,N_3424,N_3011);
nor U4322 (N_4322,N_3197,N_3245);
nand U4323 (N_4323,N_3991,N_3307);
xor U4324 (N_4324,N_3201,N_3805);
nand U4325 (N_4325,N_3077,N_3157);
or U4326 (N_4326,N_3172,N_3680);
nor U4327 (N_4327,N_3101,N_3048);
xor U4328 (N_4328,N_3932,N_3454);
xnor U4329 (N_4329,N_3306,N_3191);
nand U4330 (N_4330,N_3419,N_3304);
nor U4331 (N_4331,N_3089,N_3175);
and U4332 (N_4332,N_3606,N_3898);
xnor U4333 (N_4333,N_3538,N_3007);
and U4334 (N_4334,N_3830,N_3607);
or U4335 (N_4335,N_3537,N_3209);
nand U4336 (N_4336,N_3242,N_3160);
and U4337 (N_4337,N_3634,N_3560);
nor U4338 (N_4338,N_3070,N_3679);
and U4339 (N_4339,N_3629,N_3257);
xor U4340 (N_4340,N_3643,N_3888);
or U4341 (N_4341,N_3956,N_3182);
or U4342 (N_4342,N_3102,N_3960);
nor U4343 (N_4343,N_3111,N_3834);
nor U4344 (N_4344,N_3303,N_3608);
nor U4345 (N_4345,N_3065,N_3186);
xor U4346 (N_4346,N_3855,N_3809);
nor U4347 (N_4347,N_3297,N_3639);
or U4348 (N_4348,N_3840,N_3344);
and U4349 (N_4349,N_3617,N_3273);
nand U4350 (N_4350,N_3646,N_3778);
xnor U4351 (N_4351,N_3158,N_3393);
nor U4352 (N_4352,N_3689,N_3763);
xnor U4353 (N_4353,N_3258,N_3570);
or U4354 (N_4354,N_3707,N_3472);
xor U4355 (N_4355,N_3079,N_3765);
nand U4356 (N_4356,N_3909,N_3181);
xor U4357 (N_4357,N_3342,N_3423);
xor U4358 (N_4358,N_3224,N_3268);
or U4359 (N_4359,N_3060,N_3359);
nand U4360 (N_4360,N_3873,N_3449);
or U4361 (N_4361,N_3495,N_3119);
nor U4362 (N_4362,N_3952,N_3548);
or U4363 (N_4363,N_3871,N_3631);
xor U4364 (N_4364,N_3655,N_3725);
xnor U4365 (N_4365,N_3327,N_3566);
nand U4366 (N_4366,N_3741,N_3373);
nand U4367 (N_4367,N_3301,N_3771);
nand U4368 (N_4368,N_3105,N_3781);
and U4369 (N_4369,N_3139,N_3355);
xor U4370 (N_4370,N_3681,N_3934);
and U4371 (N_4371,N_3135,N_3404);
nand U4372 (N_4372,N_3455,N_3003);
nor U4373 (N_4373,N_3984,N_3759);
or U4374 (N_4374,N_3460,N_3708);
xnor U4375 (N_4375,N_3756,N_3828);
xnor U4376 (N_4376,N_3882,N_3411);
nor U4377 (N_4377,N_3215,N_3052);
xor U4378 (N_4378,N_3554,N_3532);
nand U4379 (N_4379,N_3407,N_3624);
xnor U4380 (N_4380,N_3173,N_3644);
and U4381 (N_4381,N_3034,N_3986);
or U4382 (N_4382,N_3218,N_3033);
nand U4383 (N_4383,N_3865,N_3133);
nand U4384 (N_4384,N_3164,N_3941);
nand U4385 (N_4385,N_3726,N_3559);
nand U4386 (N_4386,N_3345,N_3047);
or U4387 (N_4387,N_3505,N_3270);
nor U4388 (N_4388,N_3966,N_3737);
nand U4389 (N_4389,N_3000,N_3939);
and U4390 (N_4390,N_3870,N_3979);
xor U4391 (N_4391,N_3103,N_3788);
and U4392 (N_4392,N_3921,N_3683);
or U4393 (N_4393,N_3390,N_3445);
nor U4394 (N_4394,N_3908,N_3343);
nor U4395 (N_4395,N_3420,N_3789);
or U4396 (N_4396,N_3049,N_3315);
nor U4397 (N_4397,N_3959,N_3291);
or U4398 (N_4398,N_3937,N_3280);
nand U4399 (N_4399,N_3253,N_3272);
and U4400 (N_4400,N_3134,N_3902);
nor U4401 (N_4401,N_3705,N_3286);
xnor U4402 (N_4402,N_3425,N_3769);
and U4403 (N_4403,N_3154,N_3394);
or U4404 (N_4404,N_3124,N_3942);
nor U4405 (N_4405,N_3146,N_3856);
or U4406 (N_4406,N_3730,N_3085);
nand U4407 (N_4407,N_3832,N_3386);
or U4408 (N_4408,N_3858,N_3427);
and U4409 (N_4409,N_3954,N_3711);
xor U4410 (N_4410,N_3121,N_3839);
and U4411 (N_4411,N_3983,N_3260);
xnor U4412 (N_4412,N_3152,N_3587);
or U4413 (N_4413,N_3358,N_3927);
xnor U4414 (N_4414,N_3660,N_3648);
xor U4415 (N_4415,N_3481,N_3783);
nor U4416 (N_4416,N_3658,N_3117);
or U4417 (N_4417,N_3335,N_3439);
or U4418 (N_4418,N_3748,N_3347);
nor U4419 (N_4419,N_3357,N_3389);
or U4420 (N_4420,N_3349,N_3156);
and U4421 (N_4421,N_3006,N_3221);
nor U4422 (N_4422,N_3734,N_3815);
nor U4423 (N_4423,N_3795,N_3039);
nor U4424 (N_4424,N_3918,N_3328);
and U4425 (N_4425,N_3174,N_3059);
nand U4426 (N_4426,N_3090,N_3022);
nand U4427 (N_4427,N_3676,N_3413);
or U4428 (N_4428,N_3107,N_3877);
nand U4429 (N_4429,N_3899,N_3477);
or U4430 (N_4430,N_3109,N_3126);
xnor U4431 (N_4431,N_3416,N_3219);
and U4432 (N_4432,N_3980,N_3623);
nor U4433 (N_4433,N_3666,N_3944);
nor U4434 (N_4434,N_3091,N_3405);
nand U4435 (N_4435,N_3429,N_3804);
and U4436 (N_4436,N_3129,N_3515);
and U4437 (N_4437,N_3237,N_3412);
xnor U4438 (N_4438,N_3231,N_3076);
xnor U4439 (N_4439,N_3233,N_3659);
nand U4440 (N_4440,N_3588,N_3041);
and U4441 (N_4441,N_3038,N_3694);
xnor U4442 (N_4442,N_3250,N_3777);
nor U4443 (N_4443,N_3516,N_3161);
xor U4444 (N_4444,N_3170,N_3529);
nor U4445 (N_4445,N_3361,N_3536);
or U4446 (N_4446,N_3017,N_3936);
or U4447 (N_4447,N_3486,N_3586);
and U4448 (N_4448,N_3467,N_3597);
nor U4449 (N_4449,N_3082,N_3508);
or U4450 (N_4450,N_3687,N_3406);
or U4451 (N_4451,N_3025,N_3561);
nor U4452 (N_4452,N_3222,N_3024);
or U4453 (N_4453,N_3885,N_3451);
or U4454 (N_4454,N_3826,N_3989);
or U4455 (N_4455,N_3947,N_3279);
and U4456 (N_4456,N_3249,N_3513);
nor U4457 (N_4457,N_3723,N_3069);
nor U4458 (N_4458,N_3703,N_3247);
xor U4459 (N_4459,N_3990,N_3891);
and U4460 (N_4460,N_3504,N_3688);
nand U4461 (N_4461,N_3507,N_3096);
nand U4462 (N_4462,N_3064,N_3972);
nor U4463 (N_4463,N_3261,N_3014);
nand U4464 (N_4464,N_3321,N_3993);
xnor U4465 (N_4465,N_3296,N_3244);
nor U4466 (N_4466,N_3714,N_3818);
nor U4467 (N_4467,N_3651,N_3967);
and U4468 (N_4468,N_3302,N_3558);
and U4469 (N_4469,N_3996,N_3594);
and U4470 (N_4470,N_3977,N_3178);
or U4471 (N_4471,N_3724,N_3564);
nand U4472 (N_4472,N_3402,N_3240);
or U4473 (N_4473,N_3067,N_3155);
and U4474 (N_4474,N_3325,N_3417);
xnor U4475 (N_4475,N_3814,N_3528);
or U4476 (N_4476,N_3750,N_3710);
nor U4477 (N_4477,N_3287,N_3580);
and U4478 (N_4478,N_3905,N_3283);
nor U4479 (N_4479,N_3019,N_3490);
xor U4480 (N_4480,N_3884,N_3682);
nor U4481 (N_4481,N_3800,N_3514);
nand U4482 (N_4482,N_3692,N_3702);
xor U4483 (N_4483,N_3602,N_3969);
xor U4484 (N_4484,N_3691,N_3553);
nand U4485 (N_4485,N_3645,N_3001);
or U4486 (N_4486,N_3370,N_3009);
xnor U4487 (N_4487,N_3463,N_3198);
nor U4488 (N_4488,N_3095,N_3044);
or U4489 (N_4489,N_3875,N_3574);
or U4490 (N_4490,N_3254,N_3141);
and U4491 (N_4491,N_3790,N_3912);
nand U4492 (N_4492,N_3362,N_3314);
and U4493 (N_4493,N_3819,N_3919);
and U4494 (N_4494,N_3776,N_3214);
nor U4495 (N_4495,N_3053,N_3962);
or U4496 (N_4496,N_3037,N_3220);
nor U4497 (N_4497,N_3171,N_3675);
nand U4498 (N_4498,N_3720,N_3292);
nand U4499 (N_4499,N_3131,N_3527);
nand U4500 (N_4500,N_3588,N_3975);
nand U4501 (N_4501,N_3277,N_3689);
nand U4502 (N_4502,N_3198,N_3658);
nand U4503 (N_4503,N_3972,N_3517);
xor U4504 (N_4504,N_3473,N_3763);
nand U4505 (N_4505,N_3529,N_3191);
or U4506 (N_4506,N_3944,N_3155);
and U4507 (N_4507,N_3692,N_3901);
xnor U4508 (N_4508,N_3885,N_3287);
or U4509 (N_4509,N_3106,N_3789);
or U4510 (N_4510,N_3322,N_3611);
or U4511 (N_4511,N_3981,N_3499);
and U4512 (N_4512,N_3588,N_3125);
or U4513 (N_4513,N_3655,N_3593);
nor U4514 (N_4514,N_3833,N_3344);
xnor U4515 (N_4515,N_3135,N_3559);
xnor U4516 (N_4516,N_3516,N_3547);
xnor U4517 (N_4517,N_3329,N_3332);
nor U4518 (N_4518,N_3202,N_3866);
xnor U4519 (N_4519,N_3365,N_3067);
and U4520 (N_4520,N_3352,N_3203);
and U4521 (N_4521,N_3396,N_3293);
nor U4522 (N_4522,N_3453,N_3325);
nand U4523 (N_4523,N_3818,N_3404);
nor U4524 (N_4524,N_3878,N_3257);
or U4525 (N_4525,N_3870,N_3470);
and U4526 (N_4526,N_3114,N_3051);
nor U4527 (N_4527,N_3987,N_3957);
nand U4528 (N_4528,N_3453,N_3152);
or U4529 (N_4529,N_3613,N_3164);
nand U4530 (N_4530,N_3681,N_3870);
and U4531 (N_4531,N_3251,N_3229);
xnor U4532 (N_4532,N_3056,N_3142);
nand U4533 (N_4533,N_3437,N_3752);
xor U4534 (N_4534,N_3295,N_3282);
xor U4535 (N_4535,N_3542,N_3722);
and U4536 (N_4536,N_3245,N_3213);
nand U4537 (N_4537,N_3491,N_3932);
nor U4538 (N_4538,N_3562,N_3445);
nor U4539 (N_4539,N_3947,N_3362);
and U4540 (N_4540,N_3149,N_3077);
nor U4541 (N_4541,N_3443,N_3516);
or U4542 (N_4542,N_3870,N_3365);
and U4543 (N_4543,N_3308,N_3679);
xnor U4544 (N_4544,N_3542,N_3362);
or U4545 (N_4545,N_3935,N_3357);
xnor U4546 (N_4546,N_3407,N_3944);
nand U4547 (N_4547,N_3641,N_3468);
or U4548 (N_4548,N_3779,N_3657);
nand U4549 (N_4549,N_3321,N_3405);
nor U4550 (N_4550,N_3398,N_3697);
nor U4551 (N_4551,N_3601,N_3134);
nor U4552 (N_4552,N_3198,N_3066);
nor U4553 (N_4553,N_3046,N_3401);
or U4554 (N_4554,N_3739,N_3769);
nand U4555 (N_4555,N_3893,N_3533);
nand U4556 (N_4556,N_3335,N_3745);
and U4557 (N_4557,N_3501,N_3260);
or U4558 (N_4558,N_3587,N_3452);
and U4559 (N_4559,N_3149,N_3949);
or U4560 (N_4560,N_3625,N_3132);
xor U4561 (N_4561,N_3199,N_3016);
nor U4562 (N_4562,N_3258,N_3587);
and U4563 (N_4563,N_3323,N_3329);
and U4564 (N_4564,N_3744,N_3972);
and U4565 (N_4565,N_3112,N_3489);
nor U4566 (N_4566,N_3771,N_3428);
nand U4567 (N_4567,N_3254,N_3685);
nor U4568 (N_4568,N_3235,N_3958);
nor U4569 (N_4569,N_3804,N_3659);
xor U4570 (N_4570,N_3492,N_3581);
nor U4571 (N_4571,N_3271,N_3534);
nor U4572 (N_4572,N_3698,N_3726);
nand U4573 (N_4573,N_3054,N_3713);
xor U4574 (N_4574,N_3770,N_3383);
or U4575 (N_4575,N_3048,N_3036);
nand U4576 (N_4576,N_3471,N_3534);
or U4577 (N_4577,N_3917,N_3455);
and U4578 (N_4578,N_3370,N_3142);
or U4579 (N_4579,N_3601,N_3259);
nand U4580 (N_4580,N_3239,N_3667);
and U4581 (N_4581,N_3977,N_3713);
or U4582 (N_4582,N_3716,N_3577);
and U4583 (N_4583,N_3525,N_3865);
nor U4584 (N_4584,N_3238,N_3427);
and U4585 (N_4585,N_3325,N_3782);
nor U4586 (N_4586,N_3916,N_3134);
nor U4587 (N_4587,N_3572,N_3561);
nor U4588 (N_4588,N_3333,N_3098);
xnor U4589 (N_4589,N_3385,N_3300);
xnor U4590 (N_4590,N_3934,N_3706);
nand U4591 (N_4591,N_3329,N_3277);
nand U4592 (N_4592,N_3121,N_3057);
nand U4593 (N_4593,N_3304,N_3173);
nand U4594 (N_4594,N_3134,N_3926);
xor U4595 (N_4595,N_3014,N_3625);
xnor U4596 (N_4596,N_3241,N_3717);
nand U4597 (N_4597,N_3363,N_3314);
nor U4598 (N_4598,N_3203,N_3975);
and U4599 (N_4599,N_3135,N_3284);
or U4600 (N_4600,N_3551,N_3195);
and U4601 (N_4601,N_3799,N_3768);
nand U4602 (N_4602,N_3509,N_3629);
and U4603 (N_4603,N_3435,N_3854);
nand U4604 (N_4604,N_3177,N_3165);
xnor U4605 (N_4605,N_3265,N_3237);
nor U4606 (N_4606,N_3124,N_3969);
and U4607 (N_4607,N_3620,N_3901);
xor U4608 (N_4608,N_3700,N_3600);
nand U4609 (N_4609,N_3818,N_3458);
nor U4610 (N_4610,N_3083,N_3106);
nand U4611 (N_4611,N_3345,N_3708);
or U4612 (N_4612,N_3434,N_3698);
nor U4613 (N_4613,N_3419,N_3392);
nor U4614 (N_4614,N_3500,N_3295);
nor U4615 (N_4615,N_3361,N_3777);
xor U4616 (N_4616,N_3008,N_3125);
or U4617 (N_4617,N_3538,N_3305);
nand U4618 (N_4618,N_3083,N_3380);
nand U4619 (N_4619,N_3225,N_3427);
nor U4620 (N_4620,N_3596,N_3784);
and U4621 (N_4621,N_3526,N_3746);
nor U4622 (N_4622,N_3679,N_3941);
nand U4623 (N_4623,N_3956,N_3592);
xor U4624 (N_4624,N_3847,N_3180);
or U4625 (N_4625,N_3833,N_3513);
or U4626 (N_4626,N_3136,N_3585);
or U4627 (N_4627,N_3665,N_3164);
xor U4628 (N_4628,N_3252,N_3718);
and U4629 (N_4629,N_3807,N_3726);
and U4630 (N_4630,N_3951,N_3179);
or U4631 (N_4631,N_3770,N_3868);
nand U4632 (N_4632,N_3547,N_3134);
and U4633 (N_4633,N_3067,N_3559);
nor U4634 (N_4634,N_3209,N_3548);
nor U4635 (N_4635,N_3419,N_3172);
and U4636 (N_4636,N_3319,N_3236);
nand U4637 (N_4637,N_3930,N_3651);
or U4638 (N_4638,N_3041,N_3742);
xnor U4639 (N_4639,N_3665,N_3290);
and U4640 (N_4640,N_3033,N_3720);
and U4641 (N_4641,N_3867,N_3769);
and U4642 (N_4642,N_3822,N_3386);
nand U4643 (N_4643,N_3287,N_3751);
nand U4644 (N_4644,N_3051,N_3418);
or U4645 (N_4645,N_3859,N_3866);
xnor U4646 (N_4646,N_3296,N_3070);
nor U4647 (N_4647,N_3550,N_3545);
or U4648 (N_4648,N_3602,N_3869);
xor U4649 (N_4649,N_3367,N_3231);
xnor U4650 (N_4650,N_3503,N_3640);
nor U4651 (N_4651,N_3737,N_3540);
and U4652 (N_4652,N_3061,N_3235);
or U4653 (N_4653,N_3798,N_3087);
or U4654 (N_4654,N_3690,N_3416);
nor U4655 (N_4655,N_3547,N_3637);
nand U4656 (N_4656,N_3776,N_3743);
or U4657 (N_4657,N_3496,N_3650);
nor U4658 (N_4658,N_3405,N_3397);
and U4659 (N_4659,N_3126,N_3548);
xnor U4660 (N_4660,N_3161,N_3621);
or U4661 (N_4661,N_3755,N_3675);
and U4662 (N_4662,N_3369,N_3052);
and U4663 (N_4663,N_3810,N_3854);
nand U4664 (N_4664,N_3091,N_3331);
and U4665 (N_4665,N_3719,N_3605);
xnor U4666 (N_4666,N_3719,N_3971);
or U4667 (N_4667,N_3189,N_3166);
xnor U4668 (N_4668,N_3310,N_3234);
nor U4669 (N_4669,N_3026,N_3173);
nor U4670 (N_4670,N_3888,N_3649);
and U4671 (N_4671,N_3122,N_3505);
and U4672 (N_4672,N_3663,N_3795);
and U4673 (N_4673,N_3786,N_3138);
nor U4674 (N_4674,N_3935,N_3596);
or U4675 (N_4675,N_3012,N_3110);
or U4676 (N_4676,N_3697,N_3090);
and U4677 (N_4677,N_3929,N_3791);
nand U4678 (N_4678,N_3505,N_3942);
and U4679 (N_4679,N_3772,N_3300);
nand U4680 (N_4680,N_3619,N_3804);
xor U4681 (N_4681,N_3348,N_3331);
or U4682 (N_4682,N_3373,N_3029);
xnor U4683 (N_4683,N_3469,N_3691);
xnor U4684 (N_4684,N_3102,N_3830);
nor U4685 (N_4685,N_3528,N_3807);
nor U4686 (N_4686,N_3310,N_3086);
nand U4687 (N_4687,N_3242,N_3956);
or U4688 (N_4688,N_3335,N_3517);
xnor U4689 (N_4689,N_3783,N_3063);
or U4690 (N_4690,N_3814,N_3147);
xor U4691 (N_4691,N_3404,N_3323);
or U4692 (N_4692,N_3393,N_3011);
or U4693 (N_4693,N_3093,N_3440);
and U4694 (N_4694,N_3190,N_3132);
and U4695 (N_4695,N_3398,N_3051);
and U4696 (N_4696,N_3602,N_3608);
and U4697 (N_4697,N_3386,N_3688);
or U4698 (N_4698,N_3534,N_3632);
xor U4699 (N_4699,N_3863,N_3659);
and U4700 (N_4700,N_3853,N_3759);
or U4701 (N_4701,N_3978,N_3387);
nand U4702 (N_4702,N_3035,N_3341);
xor U4703 (N_4703,N_3703,N_3083);
or U4704 (N_4704,N_3540,N_3362);
nor U4705 (N_4705,N_3054,N_3288);
or U4706 (N_4706,N_3997,N_3656);
nor U4707 (N_4707,N_3332,N_3414);
nor U4708 (N_4708,N_3251,N_3728);
nand U4709 (N_4709,N_3629,N_3248);
xnor U4710 (N_4710,N_3857,N_3285);
or U4711 (N_4711,N_3060,N_3586);
and U4712 (N_4712,N_3847,N_3778);
nand U4713 (N_4713,N_3110,N_3386);
nand U4714 (N_4714,N_3569,N_3391);
nor U4715 (N_4715,N_3248,N_3188);
nor U4716 (N_4716,N_3483,N_3545);
nand U4717 (N_4717,N_3361,N_3078);
or U4718 (N_4718,N_3618,N_3892);
xnor U4719 (N_4719,N_3130,N_3122);
or U4720 (N_4720,N_3462,N_3259);
nand U4721 (N_4721,N_3638,N_3476);
xnor U4722 (N_4722,N_3459,N_3527);
xnor U4723 (N_4723,N_3511,N_3879);
and U4724 (N_4724,N_3031,N_3677);
nand U4725 (N_4725,N_3720,N_3118);
nor U4726 (N_4726,N_3805,N_3752);
or U4727 (N_4727,N_3619,N_3416);
and U4728 (N_4728,N_3847,N_3911);
nor U4729 (N_4729,N_3551,N_3624);
and U4730 (N_4730,N_3337,N_3128);
and U4731 (N_4731,N_3005,N_3317);
nor U4732 (N_4732,N_3441,N_3791);
nand U4733 (N_4733,N_3328,N_3365);
nor U4734 (N_4734,N_3163,N_3026);
nor U4735 (N_4735,N_3612,N_3515);
nor U4736 (N_4736,N_3126,N_3068);
nor U4737 (N_4737,N_3049,N_3488);
nand U4738 (N_4738,N_3735,N_3848);
nor U4739 (N_4739,N_3006,N_3907);
and U4740 (N_4740,N_3703,N_3061);
and U4741 (N_4741,N_3966,N_3338);
nand U4742 (N_4742,N_3813,N_3096);
xor U4743 (N_4743,N_3466,N_3230);
xor U4744 (N_4744,N_3931,N_3470);
nand U4745 (N_4745,N_3502,N_3960);
or U4746 (N_4746,N_3807,N_3034);
nand U4747 (N_4747,N_3526,N_3447);
or U4748 (N_4748,N_3639,N_3073);
nand U4749 (N_4749,N_3347,N_3722);
or U4750 (N_4750,N_3144,N_3879);
nand U4751 (N_4751,N_3818,N_3784);
nor U4752 (N_4752,N_3183,N_3285);
or U4753 (N_4753,N_3752,N_3417);
or U4754 (N_4754,N_3004,N_3105);
nand U4755 (N_4755,N_3408,N_3160);
nor U4756 (N_4756,N_3431,N_3550);
or U4757 (N_4757,N_3435,N_3390);
nand U4758 (N_4758,N_3597,N_3001);
and U4759 (N_4759,N_3589,N_3723);
or U4760 (N_4760,N_3853,N_3790);
nand U4761 (N_4761,N_3861,N_3298);
xnor U4762 (N_4762,N_3681,N_3155);
or U4763 (N_4763,N_3118,N_3116);
and U4764 (N_4764,N_3210,N_3310);
nor U4765 (N_4765,N_3817,N_3858);
nand U4766 (N_4766,N_3053,N_3461);
nor U4767 (N_4767,N_3060,N_3058);
nor U4768 (N_4768,N_3401,N_3482);
nand U4769 (N_4769,N_3552,N_3860);
and U4770 (N_4770,N_3789,N_3934);
and U4771 (N_4771,N_3225,N_3410);
xor U4772 (N_4772,N_3859,N_3936);
nand U4773 (N_4773,N_3070,N_3238);
xor U4774 (N_4774,N_3917,N_3218);
nand U4775 (N_4775,N_3137,N_3836);
and U4776 (N_4776,N_3216,N_3698);
xor U4777 (N_4777,N_3633,N_3789);
or U4778 (N_4778,N_3219,N_3499);
nor U4779 (N_4779,N_3550,N_3043);
or U4780 (N_4780,N_3404,N_3990);
or U4781 (N_4781,N_3893,N_3888);
nand U4782 (N_4782,N_3151,N_3731);
or U4783 (N_4783,N_3951,N_3879);
or U4784 (N_4784,N_3584,N_3144);
nor U4785 (N_4785,N_3416,N_3092);
nor U4786 (N_4786,N_3798,N_3640);
and U4787 (N_4787,N_3870,N_3327);
xor U4788 (N_4788,N_3519,N_3085);
and U4789 (N_4789,N_3957,N_3313);
and U4790 (N_4790,N_3131,N_3464);
or U4791 (N_4791,N_3419,N_3396);
nand U4792 (N_4792,N_3246,N_3145);
or U4793 (N_4793,N_3570,N_3569);
nor U4794 (N_4794,N_3043,N_3962);
or U4795 (N_4795,N_3125,N_3308);
and U4796 (N_4796,N_3262,N_3030);
and U4797 (N_4797,N_3895,N_3490);
or U4798 (N_4798,N_3009,N_3916);
and U4799 (N_4799,N_3275,N_3305);
and U4800 (N_4800,N_3219,N_3057);
xor U4801 (N_4801,N_3779,N_3003);
nor U4802 (N_4802,N_3964,N_3710);
and U4803 (N_4803,N_3230,N_3065);
or U4804 (N_4804,N_3249,N_3296);
nand U4805 (N_4805,N_3728,N_3356);
xor U4806 (N_4806,N_3394,N_3476);
or U4807 (N_4807,N_3779,N_3400);
nand U4808 (N_4808,N_3695,N_3848);
nand U4809 (N_4809,N_3289,N_3875);
and U4810 (N_4810,N_3675,N_3771);
xor U4811 (N_4811,N_3825,N_3934);
or U4812 (N_4812,N_3083,N_3902);
nand U4813 (N_4813,N_3469,N_3895);
or U4814 (N_4814,N_3143,N_3435);
nand U4815 (N_4815,N_3818,N_3767);
and U4816 (N_4816,N_3014,N_3054);
and U4817 (N_4817,N_3482,N_3185);
or U4818 (N_4818,N_3996,N_3300);
nand U4819 (N_4819,N_3505,N_3555);
nand U4820 (N_4820,N_3836,N_3082);
and U4821 (N_4821,N_3013,N_3545);
nand U4822 (N_4822,N_3090,N_3515);
and U4823 (N_4823,N_3093,N_3291);
xor U4824 (N_4824,N_3818,N_3377);
nand U4825 (N_4825,N_3538,N_3235);
nor U4826 (N_4826,N_3847,N_3890);
and U4827 (N_4827,N_3953,N_3014);
nor U4828 (N_4828,N_3961,N_3656);
xor U4829 (N_4829,N_3892,N_3087);
or U4830 (N_4830,N_3854,N_3382);
xnor U4831 (N_4831,N_3349,N_3926);
xnor U4832 (N_4832,N_3417,N_3915);
and U4833 (N_4833,N_3414,N_3379);
and U4834 (N_4834,N_3556,N_3120);
nor U4835 (N_4835,N_3267,N_3936);
xnor U4836 (N_4836,N_3753,N_3249);
or U4837 (N_4837,N_3837,N_3884);
nor U4838 (N_4838,N_3869,N_3532);
and U4839 (N_4839,N_3171,N_3601);
xnor U4840 (N_4840,N_3250,N_3345);
or U4841 (N_4841,N_3479,N_3802);
xor U4842 (N_4842,N_3209,N_3687);
nand U4843 (N_4843,N_3397,N_3157);
nor U4844 (N_4844,N_3005,N_3665);
nand U4845 (N_4845,N_3049,N_3166);
or U4846 (N_4846,N_3634,N_3963);
or U4847 (N_4847,N_3046,N_3788);
xor U4848 (N_4848,N_3773,N_3826);
xor U4849 (N_4849,N_3462,N_3648);
and U4850 (N_4850,N_3938,N_3343);
and U4851 (N_4851,N_3152,N_3952);
and U4852 (N_4852,N_3645,N_3182);
xor U4853 (N_4853,N_3506,N_3144);
or U4854 (N_4854,N_3380,N_3602);
or U4855 (N_4855,N_3243,N_3998);
or U4856 (N_4856,N_3662,N_3557);
nand U4857 (N_4857,N_3941,N_3127);
xnor U4858 (N_4858,N_3802,N_3744);
or U4859 (N_4859,N_3915,N_3460);
nor U4860 (N_4860,N_3734,N_3304);
and U4861 (N_4861,N_3176,N_3869);
nand U4862 (N_4862,N_3589,N_3389);
xor U4863 (N_4863,N_3075,N_3594);
nor U4864 (N_4864,N_3108,N_3209);
nand U4865 (N_4865,N_3992,N_3185);
and U4866 (N_4866,N_3358,N_3001);
nor U4867 (N_4867,N_3467,N_3190);
and U4868 (N_4868,N_3203,N_3868);
nor U4869 (N_4869,N_3220,N_3093);
and U4870 (N_4870,N_3623,N_3887);
or U4871 (N_4871,N_3593,N_3418);
and U4872 (N_4872,N_3017,N_3770);
and U4873 (N_4873,N_3475,N_3314);
and U4874 (N_4874,N_3691,N_3280);
and U4875 (N_4875,N_3187,N_3077);
nor U4876 (N_4876,N_3241,N_3249);
nand U4877 (N_4877,N_3939,N_3338);
nand U4878 (N_4878,N_3243,N_3520);
xor U4879 (N_4879,N_3331,N_3825);
and U4880 (N_4880,N_3447,N_3334);
nand U4881 (N_4881,N_3998,N_3578);
xor U4882 (N_4882,N_3571,N_3934);
and U4883 (N_4883,N_3193,N_3123);
or U4884 (N_4884,N_3119,N_3916);
or U4885 (N_4885,N_3302,N_3919);
nand U4886 (N_4886,N_3211,N_3629);
nor U4887 (N_4887,N_3382,N_3386);
xnor U4888 (N_4888,N_3934,N_3178);
nand U4889 (N_4889,N_3262,N_3512);
nor U4890 (N_4890,N_3516,N_3727);
nor U4891 (N_4891,N_3330,N_3855);
and U4892 (N_4892,N_3780,N_3064);
and U4893 (N_4893,N_3654,N_3803);
nor U4894 (N_4894,N_3278,N_3960);
nand U4895 (N_4895,N_3464,N_3085);
xnor U4896 (N_4896,N_3357,N_3581);
or U4897 (N_4897,N_3617,N_3796);
or U4898 (N_4898,N_3618,N_3112);
and U4899 (N_4899,N_3771,N_3523);
or U4900 (N_4900,N_3673,N_3717);
nor U4901 (N_4901,N_3987,N_3078);
xnor U4902 (N_4902,N_3002,N_3648);
xnor U4903 (N_4903,N_3641,N_3674);
or U4904 (N_4904,N_3580,N_3347);
nor U4905 (N_4905,N_3902,N_3118);
and U4906 (N_4906,N_3758,N_3822);
or U4907 (N_4907,N_3211,N_3480);
xor U4908 (N_4908,N_3844,N_3808);
xnor U4909 (N_4909,N_3560,N_3436);
or U4910 (N_4910,N_3922,N_3062);
and U4911 (N_4911,N_3842,N_3744);
nor U4912 (N_4912,N_3126,N_3130);
xnor U4913 (N_4913,N_3577,N_3956);
and U4914 (N_4914,N_3549,N_3737);
nand U4915 (N_4915,N_3824,N_3398);
nor U4916 (N_4916,N_3414,N_3403);
or U4917 (N_4917,N_3251,N_3249);
nand U4918 (N_4918,N_3830,N_3943);
nor U4919 (N_4919,N_3640,N_3117);
or U4920 (N_4920,N_3740,N_3456);
xnor U4921 (N_4921,N_3930,N_3371);
xnor U4922 (N_4922,N_3359,N_3416);
and U4923 (N_4923,N_3693,N_3159);
nand U4924 (N_4924,N_3092,N_3366);
or U4925 (N_4925,N_3705,N_3314);
and U4926 (N_4926,N_3811,N_3761);
or U4927 (N_4927,N_3765,N_3836);
and U4928 (N_4928,N_3201,N_3856);
and U4929 (N_4929,N_3738,N_3932);
xor U4930 (N_4930,N_3674,N_3473);
or U4931 (N_4931,N_3326,N_3039);
nor U4932 (N_4932,N_3820,N_3506);
or U4933 (N_4933,N_3936,N_3977);
or U4934 (N_4934,N_3691,N_3321);
xor U4935 (N_4935,N_3526,N_3036);
or U4936 (N_4936,N_3621,N_3409);
xor U4937 (N_4937,N_3130,N_3505);
or U4938 (N_4938,N_3651,N_3597);
xnor U4939 (N_4939,N_3800,N_3918);
nand U4940 (N_4940,N_3147,N_3107);
nand U4941 (N_4941,N_3560,N_3418);
nand U4942 (N_4942,N_3340,N_3612);
or U4943 (N_4943,N_3465,N_3887);
or U4944 (N_4944,N_3476,N_3872);
and U4945 (N_4945,N_3096,N_3649);
or U4946 (N_4946,N_3797,N_3907);
nor U4947 (N_4947,N_3615,N_3132);
or U4948 (N_4948,N_3157,N_3056);
and U4949 (N_4949,N_3973,N_3792);
or U4950 (N_4950,N_3612,N_3695);
xor U4951 (N_4951,N_3901,N_3000);
and U4952 (N_4952,N_3004,N_3580);
nor U4953 (N_4953,N_3498,N_3472);
or U4954 (N_4954,N_3883,N_3249);
nand U4955 (N_4955,N_3001,N_3949);
nor U4956 (N_4956,N_3257,N_3822);
nor U4957 (N_4957,N_3058,N_3722);
and U4958 (N_4958,N_3978,N_3820);
xnor U4959 (N_4959,N_3700,N_3310);
nor U4960 (N_4960,N_3378,N_3306);
nand U4961 (N_4961,N_3603,N_3875);
and U4962 (N_4962,N_3844,N_3148);
nor U4963 (N_4963,N_3530,N_3914);
and U4964 (N_4964,N_3857,N_3644);
xor U4965 (N_4965,N_3633,N_3791);
nand U4966 (N_4966,N_3227,N_3911);
xnor U4967 (N_4967,N_3880,N_3469);
nand U4968 (N_4968,N_3679,N_3726);
xnor U4969 (N_4969,N_3404,N_3289);
and U4970 (N_4970,N_3138,N_3965);
or U4971 (N_4971,N_3293,N_3683);
nor U4972 (N_4972,N_3429,N_3965);
xor U4973 (N_4973,N_3577,N_3690);
nor U4974 (N_4974,N_3931,N_3054);
xor U4975 (N_4975,N_3020,N_3115);
or U4976 (N_4976,N_3847,N_3965);
or U4977 (N_4977,N_3263,N_3865);
nand U4978 (N_4978,N_3644,N_3757);
nor U4979 (N_4979,N_3508,N_3042);
nor U4980 (N_4980,N_3900,N_3349);
and U4981 (N_4981,N_3230,N_3191);
xor U4982 (N_4982,N_3039,N_3960);
nor U4983 (N_4983,N_3058,N_3432);
and U4984 (N_4984,N_3918,N_3192);
nor U4985 (N_4985,N_3881,N_3696);
nand U4986 (N_4986,N_3129,N_3003);
nor U4987 (N_4987,N_3377,N_3399);
xor U4988 (N_4988,N_3794,N_3219);
xor U4989 (N_4989,N_3327,N_3938);
xnor U4990 (N_4990,N_3625,N_3442);
nand U4991 (N_4991,N_3145,N_3061);
and U4992 (N_4992,N_3898,N_3894);
nor U4993 (N_4993,N_3566,N_3902);
nor U4994 (N_4994,N_3682,N_3553);
xor U4995 (N_4995,N_3478,N_3715);
xor U4996 (N_4996,N_3101,N_3283);
nand U4997 (N_4997,N_3928,N_3157);
nor U4998 (N_4998,N_3426,N_3478);
nor U4999 (N_4999,N_3200,N_3638);
nand U5000 (N_5000,N_4245,N_4857);
nand U5001 (N_5001,N_4499,N_4617);
or U5002 (N_5002,N_4235,N_4162);
or U5003 (N_5003,N_4516,N_4152);
and U5004 (N_5004,N_4914,N_4785);
or U5005 (N_5005,N_4236,N_4514);
nand U5006 (N_5006,N_4479,N_4070);
nand U5007 (N_5007,N_4530,N_4438);
or U5008 (N_5008,N_4822,N_4435);
nor U5009 (N_5009,N_4296,N_4308);
nand U5010 (N_5010,N_4420,N_4050);
xnor U5011 (N_5011,N_4712,N_4574);
nor U5012 (N_5012,N_4706,N_4551);
nand U5013 (N_5013,N_4628,N_4796);
xnor U5014 (N_5014,N_4542,N_4772);
nand U5015 (N_5015,N_4798,N_4925);
nand U5016 (N_5016,N_4836,N_4404);
nand U5017 (N_5017,N_4111,N_4249);
nand U5018 (N_5018,N_4810,N_4428);
and U5019 (N_5019,N_4447,N_4646);
xnor U5020 (N_5020,N_4618,N_4139);
nor U5021 (N_5021,N_4960,N_4086);
xor U5022 (N_5022,N_4113,N_4945);
nand U5023 (N_5023,N_4425,N_4667);
or U5024 (N_5024,N_4434,N_4575);
or U5025 (N_5025,N_4637,N_4660);
and U5026 (N_5026,N_4862,N_4506);
and U5027 (N_5027,N_4768,N_4054);
and U5028 (N_5028,N_4399,N_4795);
and U5029 (N_5029,N_4647,N_4031);
xnor U5030 (N_5030,N_4163,N_4649);
nand U5031 (N_5031,N_4701,N_4352);
or U5032 (N_5032,N_4418,N_4902);
or U5033 (N_5033,N_4926,N_4720);
nand U5034 (N_5034,N_4200,N_4459);
and U5035 (N_5035,N_4354,N_4958);
or U5036 (N_5036,N_4167,N_4419);
and U5037 (N_5037,N_4762,N_4155);
xnor U5038 (N_5038,N_4266,N_4400);
nor U5039 (N_5039,N_4933,N_4893);
nand U5040 (N_5040,N_4251,N_4688);
and U5041 (N_5041,N_4461,N_4882);
nor U5042 (N_5042,N_4346,N_4788);
or U5043 (N_5043,N_4654,N_4085);
nand U5044 (N_5044,N_4759,N_4069);
and U5045 (N_5045,N_4002,N_4920);
or U5046 (N_5046,N_4967,N_4659);
and U5047 (N_5047,N_4600,N_4465);
nor U5048 (N_5048,N_4135,N_4755);
or U5049 (N_5049,N_4820,N_4790);
nand U5050 (N_5050,N_4067,N_4416);
xor U5051 (N_5051,N_4833,N_4169);
and U5052 (N_5052,N_4073,N_4782);
nor U5053 (N_5053,N_4319,N_4947);
nor U5054 (N_5054,N_4008,N_4809);
and U5055 (N_5055,N_4905,N_4766);
nor U5056 (N_5056,N_4781,N_4440);
and U5057 (N_5057,N_4627,N_4068);
or U5058 (N_5058,N_4610,N_4382);
nor U5059 (N_5059,N_4472,N_4823);
or U5060 (N_5060,N_4394,N_4669);
xnor U5061 (N_5061,N_4645,N_4448);
nor U5062 (N_5062,N_4477,N_4621);
xnor U5063 (N_5063,N_4579,N_4132);
nor U5064 (N_5064,N_4909,N_4577);
xnor U5065 (N_5065,N_4345,N_4136);
nor U5066 (N_5066,N_4769,N_4391);
xor U5067 (N_5067,N_4800,N_4183);
nand U5068 (N_5068,N_4306,N_4558);
xor U5069 (N_5069,N_4992,N_4032);
or U5070 (N_5070,N_4390,N_4268);
xor U5071 (N_5071,N_4223,N_4494);
nor U5072 (N_5072,N_4034,N_4110);
nor U5073 (N_5073,N_4778,N_4733);
xnor U5074 (N_5074,N_4289,N_4896);
nand U5075 (N_5075,N_4606,N_4535);
or U5076 (N_5076,N_4300,N_4238);
nand U5077 (N_5077,N_4738,N_4567);
or U5078 (N_5078,N_4279,N_4021);
nand U5079 (N_5079,N_4675,N_4184);
nor U5080 (N_5080,N_4464,N_4367);
nor U5081 (N_5081,N_4397,N_4969);
nor U5082 (N_5082,N_4554,N_4944);
and U5083 (N_5083,N_4817,N_4341);
and U5084 (N_5084,N_4087,N_4512);
or U5085 (N_5085,N_4732,N_4194);
or U5086 (N_5086,N_4583,N_4107);
and U5087 (N_5087,N_4897,N_4175);
nand U5088 (N_5088,N_4985,N_4791);
or U5089 (N_5089,N_4090,N_4919);
and U5090 (N_5090,N_4539,N_4414);
nor U5091 (N_5091,N_4240,N_4563);
nand U5092 (N_5092,N_4550,N_4062);
xor U5093 (N_5093,N_4195,N_4784);
and U5094 (N_5094,N_4994,N_4865);
xnor U5095 (N_5095,N_4060,N_4509);
xnor U5096 (N_5096,N_4389,N_4138);
xnor U5097 (N_5097,N_4177,N_4265);
nand U5098 (N_5098,N_4084,N_4151);
and U5099 (N_5099,N_4779,N_4642);
xnor U5100 (N_5100,N_4964,N_4189);
nor U5101 (N_5101,N_4248,N_4871);
and U5102 (N_5102,N_4777,N_4363);
or U5103 (N_5103,N_4039,N_4611);
nand U5104 (N_5104,N_4749,N_4752);
nor U5105 (N_5105,N_4388,N_4063);
nor U5106 (N_5106,N_4100,N_4475);
or U5107 (N_5107,N_4540,N_4044);
or U5108 (N_5108,N_4536,N_4644);
or U5109 (N_5109,N_4453,N_4584);
or U5110 (N_5110,N_4529,N_4601);
or U5111 (N_5111,N_4524,N_4874);
and U5112 (N_5112,N_4545,N_4984);
nor U5113 (N_5113,N_4292,N_4689);
nand U5114 (N_5114,N_4674,N_4504);
xnor U5115 (N_5115,N_4928,N_4305);
nor U5116 (N_5116,N_4557,N_4204);
and U5117 (N_5117,N_4685,N_4590);
nor U5118 (N_5118,N_4597,N_4185);
nand U5119 (N_5119,N_4114,N_4112);
nand U5120 (N_5120,N_4285,N_4402);
xnor U5121 (N_5121,N_4878,N_4742);
nand U5122 (N_5122,N_4199,N_4001);
or U5123 (N_5123,N_4312,N_4497);
nor U5124 (N_5124,N_4852,N_4144);
nand U5125 (N_5125,N_4255,N_4115);
and U5126 (N_5126,N_4526,N_4966);
or U5127 (N_5127,N_4356,N_4883);
or U5128 (N_5128,N_4188,N_4323);
or U5129 (N_5129,N_4716,N_4775);
and U5130 (N_5130,N_4117,N_4821);
nor U5131 (N_5131,N_4968,N_4517);
xor U5132 (N_5132,N_4409,N_4190);
nor U5133 (N_5133,N_4206,N_4377);
nor U5134 (N_5134,N_4916,N_4929);
or U5135 (N_5135,N_4875,N_4787);
nand U5136 (N_5136,N_4744,N_4614);
xnor U5137 (N_5137,N_4845,N_4398);
or U5138 (N_5138,N_4095,N_4217);
or U5139 (N_5139,N_4057,N_4080);
or U5140 (N_5140,N_4620,N_4375);
xor U5141 (N_5141,N_4757,N_4205);
xor U5142 (N_5142,N_4867,N_4172);
nand U5143 (N_5143,N_4089,N_4527);
nand U5144 (N_5144,N_4708,N_4005);
nand U5145 (N_5145,N_4840,N_4518);
nand U5146 (N_5146,N_4962,N_4892);
xor U5147 (N_5147,N_4898,N_4123);
xor U5148 (N_5148,N_4666,N_4049);
nand U5149 (N_5149,N_4260,N_4756);
or U5150 (N_5150,N_4181,N_4083);
and U5151 (N_5151,N_4835,N_4580);
nor U5152 (N_5152,N_4267,N_4048);
nand U5153 (N_5153,N_4912,N_4587);
nand U5154 (N_5154,N_4218,N_4652);
and U5155 (N_5155,N_4740,N_4826);
nor U5156 (N_5156,N_4664,N_4815);
or U5157 (N_5157,N_4168,N_4698);
xnor U5158 (N_5158,N_4573,N_4956);
xnor U5159 (N_5159,N_4941,N_4449);
or U5160 (N_5160,N_4564,N_4870);
or U5161 (N_5161,N_4816,N_4326);
nand U5162 (N_5162,N_4348,N_4244);
xor U5163 (N_5163,N_4441,N_4598);
and U5164 (N_5164,N_4156,N_4018);
or U5165 (N_5165,N_4490,N_4714);
nand U5166 (N_5166,N_4247,N_4886);
xnor U5167 (N_5167,N_4640,N_4071);
or U5168 (N_5168,N_4340,N_4496);
nand U5169 (N_5169,N_4844,N_4128);
xor U5170 (N_5170,N_4805,N_4252);
xnor U5171 (N_5171,N_4224,N_4794);
nand U5172 (N_5172,N_4328,N_4332);
nand U5173 (N_5173,N_4015,N_4361);
or U5174 (N_5174,N_4819,N_4212);
xor U5175 (N_5175,N_4572,N_4849);
or U5176 (N_5176,N_4722,N_4301);
nand U5177 (N_5177,N_4770,N_4040);
nor U5178 (N_5178,N_4066,N_4754);
xnor U5179 (N_5179,N_4847,N_4273);
or U5180 (N_5180,N_4746,N_4250);
nand U5181 (N_5181,N_4231,N_4006);
and U5182 (N_5182,N_4724,N_4170);
and U5183 (N_5183,N_4451,N_4274);
xor U5184 (N_5184,N_4313,N_4476);
nand U5185 (N_5185,N_4264,N_4661);
and U5186 (N_5186,N_4099,N_4201);
or U5187 (N_5187,N_4275,N_4478);
and U5188 (N_5188,N_4541,N_4663);
or U5189 (N_5189,N_4237,N_4693);
nor U5190 (N_5190,N_4403,N_4012);
xor U5191 (N_5191,N_4094,N_4159);
or U5192 (N_5192,N_4043,N_4373);
nor U5193 (N_5193,N_4780,N_4767);
nand U5194 (N_5194,N_4904,N_4894);
or U5195 (N_5195,N_4327,N_4207);
xnor U5196 (N_5196,N_4830,N_4225);
nor U5197 (N_5197,N_4405,N_4284);
xor U5198 (N_5198,N_4197,N_4142);
nand U5199 (N_5199,N_4764,N_4337);
and U5200 (N_5200,N_4407,N_4814);
and U5201 (N_5201,N_4466,N_4020);
and U5202 (N_5202,N_4276,N_4046);
or U5203 (N_5203,N_4091,N_4304);
xor U5204 (N_5204,N_4662,N_4711);
xor U5205 (N_5205,N_4609,N_4634);
xnor U5206 (N_5206,N_4565,N_4687);
or U5207 (N_5207,N_4379,N_4710);
and U5208 (N_5208,N_4707,N_4650);
and U5209 (N_5209,N_4220,N_4092);
nor U5210 (N_5210,N_4013,N_4677);
nand U5211 (N_5211,N_4473,N_4331);
nand U5212 (N_5212,N_4961,N_4741);
or U5213 (N_5213,N_4619,N_4522);
nand U5214 (N_5214,N_4360,N_4651);
nand U5215 (N_5215,N_4846,N_4730);
and U5216 (N_5216,N_4173,N_4854);
or U5217 (N_5217,N_4719,N_4934);
xor U5218 (N_5218,N_4624,N_4807);
and U5219 (N_5219,N_4818,N_4374);
nand U5220 (N_5220,N_4347,N_4198);
and U5221 (N_5221,N_4316,N_4510);
nor U5222 (N_5222,N_4813,N_4436);
or U5223 (N_5223,N_4042,N_4148);
or U5224 (N_5224,N_4072,N_4942);
xnor U5225 (N_5225,N_4576,N_4949);
and U5226 (N_5226,N_4271,N_4653);
nand U5227 (N_5227,N_4191,N_4676);
or U5228 (N_5228,N_4828,N_4310);
nor U5229 (N_5229,N_4922,N_4413);
and U5230 (N_5230,N_4444,N_4485);
and U5231 (N_5231,N_4839,N_4578);
and U5232 (N_5232,N_4480,N_4439);
nand U5233 (N_5233,N_4432,N_4082);
nand U5234 (N_5234,N_4804,N_4736);
or U5235 (N_5235,N_4989,N_4433);
nand U5236 (N_5236,N_4026,N_4950);
and U5237 (N_5237,N_4076,N_4307);
or U5238 (N_5238,N_4443,N_4290);
nor U5239 (N_5239,N_4125,N_4311);
or U5240 (N_5240,N_4513,N_4939);
nor U5241 (N_5241,N_4729,N_4981);
and U5242 (N_5242,N_4641,N_4555);
or U5243 (N_5243,N_4129,N_4164);
and U5244 (N_5244,N_4548,N_4131);
nand U5245 (N_5245,N_4531,N_4035);
xor U5246 (N_5246,N_4569,N_4500);
and U5247 (N_5247,N_4229,N_4078);
nand U5248 (N_5248,N_4421,N_4010);
or U5249 (N_5249,N_4126,N_4498);
nand U5250 (N_5250,N_4334,N_4027);
or U5251 (N_5251,N_4105,N_4869);
xnor U5252 (N_5252,N_4482,N_4723);
nor U5253 (N_5253,N_4806,N_4612);
nor U5254 (N_5254,N_4460,N_4365);
xor U5255 (N_5255,N_4931,N_4362);
nor U5256 (N_5256,N_4033,N_4519);
nor U5257 (N_5257,N_4014,N_4471);
or U5258 (N_5258,N_4387,N_4630);
and U5259 (N_5259,N_4045,N_4915);
and U5260 (N_5260,N_4431,N_4457);
xor U5261 (N_5261,N_4437,N_4302);
and U5262 (N_5262,N_4680,N_4684);
nand U5263 (N_5263,N_4446,N_4940);
nor U5264 (N_5264,N_4488,N_4463);
or U5265 (N_5265,N_4349,N_4074);
nand U5266 (N_5266,N_4607,N_4253);
xor U5267 (N_5267,N_4228,N_4280);
nor U5268 (N_5268,N_4291,N_4287);
and U5269 (N_5269,N_4843,N_4203);
or U5270 (N_5270,N_4986,N_4546);
nor U5271 (N_5271,N_4880,N_4511);
nand U5272 (N_5272,N_4995,N_4145);
nor U5273 (N_5273,N_4470,N_4242);
or U5274 (N_5274,N_4158,N_4016);
xor U5275 (N_5275,N_4562,N_4106);
or U5276 (N_5276,N_4282,N_4368);
xor U5277 (N_5277,N_4834,N_4081);
nand U5278 (N_5278,N_4118,N_4501);
xor U5279 (N_5279,N_4671,N_4560);
and U5280 (N_5280,N_4568,N_4879);
and U5281 (N_5281,N_4422,N_4978);
or U5282 (N_5282,N_4987,N_4004);
and U5283 (N_5283,N_4889,N_4691);
nand U5284 (N_5284,N_4241,N_4298);
nand U5285 (N_5285,N_4553,N_4802);
nor U5286 (N_5286,N_4797,N_4219);
nor U5287 (N_5287,N_4592,N_4455);
nor U5288 (N_5288,N_4952,N_4727);
or U5289 (N_5289,N_4096,N_4335);
and U5290 (N_5290,N_4765,N_4127);
nor U5291 (N_5291,N_4116,N_4980);
xnor U5292 (N_5292,N_4381,N_4976);
xor U5293 (N_5293,N_4186,N_4411);
nor U5294 (N_5294,N_4863,N_4261);
or U5295 (N_5295,N_4990,N_4364);
nand U5296 (N_5296,N_4988,N_4193);
nor U5297 (N_5297,N_4591,N_4695);
nor U5298 (N_5298,N_4380,N_4528);
nor U5299 (N_5299,N_4355,N_4700);
and U5300 (N_5300,N_4523,N_4595);
nor U5301 (N_5301,N_4841,N_4119);
and U5302 (N_5302,N_4903,N_4538);
xnor U5303 (N_5303,N_4864,N_4948);
nor U5304 (N_5304,N_4808,N_4632);
xnor U5305 (N_5305,N_4140,N_4344);
xnor U5306 (N_5306,N_4616,N_4288);
nor U5307 (N_5307,N_4629,N_4907);
nand U5308 (N_5308,N_4927,N_4101);
xor U5309 (N_5309,N_4581,N_4038);
nor U5310 (N_5310,N_4486,N_4481);
and U5311 (N_5311,N_4887,N_4406);
and U5312 (N_5312,N_4593,N_4051);
and U5313 (N_5313,N_4702,N_4429);
or U5314 (N_5314,N_4303,N_4508);
nand U5315 (N_5315,N_4622,N_4133);
and U5316 (N_5316,N_4801,N_4997);
or U5317 (N_5317,N_4525,N_4643);
and U5318 (N_5318,N_4491,N_4900);
and U5319 (N_5319,N_4343,N_4998);
nor U5320 (N_5320,N_4556,N_4254);
nor U5321 (N_5321,N_4187,N_4673);
xnor U5322 (N_5322,N_4951,N_4061);
and U5323 (N_5323,N_4369,N_4561);
and U5324 (N_5324,N_4342,N_4717);
xor U5325 (N_5325,N_4665,N_4633);
nor U5326 (N_5326,N_4921,N_4751);
or U5327 (N_5327,N_4594,N_4745);
and U5328 (N_5328,N_4150,N_4393);
nor U5329 (N_5329,N_4009,N_4851);
xnor U5330 (N_5330,N_4336,N_4631);
or U5331 (N_5331,N_4024,N_4454);
xor U5332 (N_5332,N_4829,N_4281);
or U5333 (N_5333,N_4211,N_4655);
nor U5334 (N_5334,N_4739,N_4868);
and U5335 (N_5335,N_4171,N_4837);
nand U5336 (N_5336,N_4353,N_4503);
nor U5337 (N_5337,N_4608,N_4648);
xor U5338 (N_5338,N_4325,N_4917);
nand U5339 (N_5339,N_4955,N_4410);
nor U5340 (N_5340,N_4657,N_4278);
nand U5341 (N_5341,N_4726,N_4263);
nand U5342 (N_5342,N_4605,N_4639);
and U5343 (N_5343,N_4321,N_4991);
and U5344 (N_5344,N_4370,N_4521);
and U5345 (N_5345,N_4737,N_4103);
and U5346 (N_5346,N_4697,N_4146);
and U5347 (N_5347,N_4971,N_4532);
or U5348 (N_5348,N_4309,N_4682);
xor U5349 (N_5349,N_4214,N_4121);
xor U5350 (N_5350,N_4339,N_4690);
nand U5351 (N_5351,N_4876,N_4623);
or U5352 (N_5352,N_4458,N_4256);
xor U5353 (N_5353,N_4913,N_4943);
and U5354 (N_5354,N_4147,N_4036);
or U5355 (N_5355,N_4104,N_4549);
nor U5356 (N_5356,N_4866,N_4141);
and U5357 (N_5357,N_4773,N_4566);
nand U5358 (N_5358,N_4963,N_4210);
and U5359 (N_5359,N_4753,N_4456);
nor U5360 (N_5360,N_4239,N_4371);
nand U5361 (N_5361,N_4993,N_4603);
xor U5362 (N_5362,N_4696,N_4075);
nand U5363 (N_5363,N_4208,N_4077);
nand U5364 (N_5364,N_4395,N_4350);
nor U5365 (N_5365,N_4378,N_4462);
nor U5366 (N_5366,N_4028,N_4196);
and U5367 (N_5367,N_4317,N_4970);
and U5368 (N_5368,N_4983,N_4924);
nand U5369 (N_5369,N_4445,N_4743);
or U5370 (N_5370,N_4295,N_4093);
nand U5371 (N_5371,N_4906,N_4856);
xnor U5372 (N_5372,N_4474,N_4493);
and U5373 (N_5373,N_4396,N_4636);
nor U5374 (N_5374,N_4789,N_4358);
xnor U5375 (N_5375,N_4615,N_4859);
or U5376 (N_5376,N_4489,N_4703);
nand U5377 (N_5377,N_4977,N_4423);
xor U5378 (N_5378,N_4771,N_4972);
xor U5379 (N_5379,N_4330,N_4811);
nand U5380 (N_5380,N_4022,N_4705);
and U5381 (N_5381,N_4827,N_4174);
xor U5382 (N_5382,N_4625,N_4495);
xor U5383 (N_5383,N_4315,N_4023);
xor U5384 (N_5384,N_4715,N_4386);
or U5385 (N_5385,N_4954,N_4761);
or U5386 (N_5386,N_4679,N_4333);
xnor U5387 (N_5387,N_4246,N_4234);
nor U5388 (N_5388,N_4812,N_4037);
nand U5389 (N_5389,N_4709,N_4544);
and U5390 (N_5390,N_4957,N_4401);
and U5391 (N_5391,N_4872,N_4672);
or U5392 (N_5392,N_4025,N_4946);
nand U5393 (N_5393,N_4824,N_4029);
nand U5394 (N_5394,N_4257,N_4272);
and U5395 (N_5395,N_4728,N_4873);
and U5396 (N_5396,N_4430,N_4047);
nand U5397 (N_5397,N_4881,N_4003);
nor U5398 (N_5398,N_4799,N_4585);
or U5399 (N_5399,N_4178,N_4681);
nand U5400 (N_5400,N_4936,N_4179);
xnor U5401 (N_5401,N_4877,N_4277);
xor U5402 (N_5402,N_4979,N_4861);
or U5403 (N_5403,N_4832,N_4792);
nand U5404 (N_5404,N_4232,N_4923);
xnor U5405 (N_5405,N_4314,N_4450);
and U5406 (N_5406,N_4901,N_4270);
and U5407 (N_5407,N_4226,N_4383);
xor U5408 (N_5408,N_4392,N_4570);
nand U5409 (N_5409,N_4176,N_4599);
nor U5410 (N_5410,N_4102,N_4124);
and U5411 (N_5411,N_4351,N_4259);
nor U5412 (N_5412,N_4357,N_4098);
and U5413 (N_5413,N_4937,N_4783);
or U5414 (N_5414,N_4318,N_4059);
xor U5415 (N_5415,N_4774,N_4758);
nor U5416 (N_5416,N_4216,N_4965);
nand U5417 (N_5417,N_4735,N_4065);
or U5418 (N_5418,N_4213,N_4613);
or U5419 (N_5419,N_4166,N_4384);
or U5420 (N_5420,N_4959,N_4019);
or U5421 (N_5421,N_4996,N_4515);
or U5422 (N_5422,N_4953,N_4017);
nor U5423 (N_5423,N_4858,N_4324);
xnor U5424 (N_5424,N_4547,N_4750);
or U5425 (N_5425,N_4297,N_4202);
nor U5426 (N_5426,N_4860,N_4683);
xor U5427 (N_5427,N_4134,N_4221);
or U5428 (N_5428,N_4895,N_4154);
nand U5429 (N_5429,N_4322,N_4492);
or U5430 (N_5430,N_4786,N_4932);
nand U5431 (N_5431,N_4699,N_4588);
xor U5432 (N_5432,N_4359,N_4692);
xnor U5433 (N_5433,N_4502,N_4122);
or U5434 (N_5434,N_4215,N_4533);
nor U5435 (N_5435,N_4670,N_4803);
and U5436 (N_5436,N_4999,N_4222);
and U5437 (N_5437,N_4372,N_4776);
nand U5438 (N_5438,N_4484,N_4678);
nor U5439 (N_5439,N_4537,N_4058);
nor U5440 (N_5440,N_4721,N_4731);
or U5441 (N_5441,N_4725,N_4329);
and U5442 (N_5442,N_4052,N_4890);
xnor U5443 (N_5443,N_4408,N_4097);
nor U5444 (N_5444,N_4793,N_4694);
xor U5445 (N_5445,N_4534,N_4262);
or U5446 (N_5446,N_4120,N_4658);
xor U5447 (N_5447,N_4505,N_4320);
and U5448 (N_5448,N_4734,N_4713);
xor U5449 (N_5449,N_4283,N_4899);
or U5450 (N_5450,N_4487,N_4938);
or U5451 (N_5451,N_4596,N_4974);
nor U5452 (N_5452,N_4041,N_4415);
xnor U5453 (N_5453,N_4638,N_4831);
or U5454 (N_5454,N_4853,N_4850);
and U5455 (N_5455,N_4842,N_4269);
and U5456 (N_5456,N_4559,N_4930);
xor U5457 (N_5457,N_4137,N_4884);
and U5458 (N_5458,N_4975,N_4299);
and U5459 (N_5459,N_4908,N_4626);
and U5460 (N_5460,N_4161,N_4376);
xnor U5461 (N_5461,N_4424,N_4589);
nand U5462 (N_5462,N_4088,N_4079);
nor U5463 (N_5463,N_4109,N_4855);
and U5464 (N_5464,N_4385,N_4412);
nand U5465 (N_5465,N_4825,N_4571);
nor U5466 (N_5466,N_4911,N_4192);
nand U5467 (N_5467,N_4007,N_4426);
nand U5468 (N_5468,N_4468,N_4130);
xor U5469 (N_5469,N_4602,N_4143);
nand U5470 (N_5470,N_4760,N_4552);
and U5471 (N_5471,N_4520,N_4582);
xor U5472 (N_5472,N_4230,N_4763);
or U5473 (N_5473,N_4293,N_4053);
nand U5474 (N_5474,N_4153,N_4483);
xnor U5475 (N_5475,N_4888,N_4182);
and U5476 (N_5476,N_4586,N_4011);
and U5477 (N_5477,N_4157,N_4180);
nand U5478 (N_5478,N_4030,N_4160);
xor U5479 (N_5479,N_4165,N_4469);
or U5480 (N_5480,N_4227,N_4910);
and U5481 (N_5481,N_4108,N_4848);
nand U5482 (N_5482,N_4243,N_4656);
or U5483 (N_5483,N_4452,N_4442);
xnor U5484 (N_5484,N_4507,N_4668);
xor U5485 (N_5485,N_4366,N_4718);
and U5486 (N_5486,N_4467,N_4543);
nand U5487 (N_5487,N_4338,N_4973);
nand U5488 (N_5488,N_4635,N_4747);
and U5489 (N_5489,N_4885,N_4233);
and U5490 (N_5490,N_4417,N_4427);
and U5491 (N_5491,N_4686,N_4918);
nor U5492 (N_5492,N_4294,N_4935);
or U5493 (N_5493,N_4064,N_4748);
or U5494 (N_5494,N_4838,N_4258);
xor U5495 (N_5495,N_4286,N_4149);
nor U5496 (N_5496,N_4056,N_4055);
nor U5497 (N_5497,N_4891,N_4604);
or U5498 (N_5498,N_4704,N_4000);
nor U5499 (N_5499,N_4982,N_4209);
and U5500 (N_5500,N_4615,N_4754);
nand U5501 (N_5501,N_4903,N_4183);
xnor U5502 (N_5502,N_4851,N_4265);
xor U5503 (N_5503,N_4932,N_4670);
xnor U5504 (N_5504,N_4448,N_4642);
nor U5505 (N_5505,N_4192,N_4213);
and U5506 (N_5506,N_4748,N_4379);
nor U5507 (N_5507,N_4393,N_4191);
nand U5508 (N_5508,N_4012,N_4595);
and U5509 (N_5509,N_4396,N_4427);
xor U5510 (N_5510,N_4227,N_4102);
xnor U5511 (N_5511,N_4325,N_4533);
xor U5512 (N_5512,N_4274,N_4320);
xnor U5513 (N_5513,N_4922,N_4347);
nor U5514 (N_5514,N_4653,N_4279);
nand U5515 (N_5515,N_4788,N_4867);
nor U5516 (N_5516,N_4957,N_4497);
and U5517 (N_5517,N_4984,N_4113);
nor U5518 (N_5518,N_4813,N_4419);
xnor U5519 (N_5519,N_4185,N_4207);
nand U5520 (N_5520,N_4723,N_4916);
or U5521 (N_5521,N_4949,N_4442);
nand U5522 (N_5522,N_4450,N_4661);
or U5523 (N_5523,N_4759,N_4387);
nand U5524 (N_5524,N_4125,N_4398);
and U5525 (N_5525,N_4517,N_4061);
or U5526 (N_5526,N_4143,N_4624);
nand U5527 (N_5527,N_4650,N_4909);
xnor U5528 (N_5528,N_4635,N_4055);
nand U5529 (N_5529,N_4669,N_4465);
or U5530 (N_5530,N_4170,N_4086);
nand U5531 (N_5531,N_4063,N_4506);
or U5532 (N_5532,N_4322,N_4351);
or U5533 (N_5533,N_4242,N_4180);
or U5534 (N_5534,N_4120,N_4427);
and U5535 (N_5535,N_4320,N_4479);
nand U5536 (N_5536,N_4102,N_4687);
xnor U5537 (N_5537,N_4869,N_4950);
nand U5538 (N_5538,N_4373,N_4746);
nand U5539 (N_5539,N_4200,N_4186);
nor U5540 (N_5540,N_4690,N_4501);
nor U5541 (N_5541,N_4573,N_4354);
nand U5542 (N_5542,N_4189,N_4038);
xnor U5543 (N_5543,N_4499,N_4329);
nor U5544 (N_5544,N_4728,N_4095);
nand U5545 (N_5545,N_4915,N_4210);
nor U5546 (N_5546,N_4591,N_4633);
xor U5547 (N_5547,N_4074,N_4893);
or U5548 (N_5548,N_4664,N_4045);
nand U5549 (N_5549,N_4873,N_4357);
nor U5550 (N_5550,N_4841,N_4054);
and U5551 (N_5551,N_4274,N_4510);
nand U5552 (N_5552,N_4934,N_4422);
xor U5553 (N_5553,N_4948,N_4374);
xor U5554 (N_5554,N_4094,N_4582);
or U5555 (N_5555,N_4655,N_4871);
nand U5556 (N_5556,N_4929,N_4934);
or U5557 (N_5557,N_4431,N_4116);
nor U5558 (N_5558,N_4998,N_4197);
xnor U5559 (N_5559,N_4745,N_4749);
nand U5560 (N_5560,N_4904,N_4003);
nor U5561 (N_5561,N_4794,N_4738);
nor U5562 (N_5562,N_4043,N_4685);
and U5563 (N_5563,N_4077,N_4281);
nand U5564 (N_5564,N_4804,N_4425);
or U5565 (N_5565,N_4691,N_4862);
nand U5566 (N_5566,N_4446,N_4526);
or U5567 (N_5567,N_4680,N_4612);
or U5568 (N_5568,N_4977,N_4117);
nor U5569 (N_5569,N_4314,N_4310);
nand U5570 (N_5570,N_4852,N_4153);
and U5571 (N_5571,N_4332,N_4861);
and U5572 (N_5572,N_4704,N_4372);
and U5573 (N_5573,N_4070,N_4533);
nor U5574 (N_5574,N_4874,N_4612);
or U5575 (N_5575,N_4651,N_4431);
nor U5576 (N_5576,N_4153,N_4428);
nor U5577 (N_5577,N_4392,N_4013);
and U5578 (N_5578,N_4119,N_4854);
xnor U5579 (N_5579,N_4023,N_4171);
nor U5580 (N_5580,N_4083,N_4172);
nand U5581 (N_5581,N_4204,N_4750);
and U5582 (N_5582,N_4993,N_4879);
nand U5583 (N_5583,N_4149,N_4577);
nor U5584 (N_5584,N_4149,N_4277);
nand U5585 (N_5585,N_4847,N_4550);
nor U5586 (N_5586,N_4969,N_4187);
nor U5587 (N_5587,N_4014,N_4347);
nand U5588 (N_5588,N_4083,N_4149);
xor U5589 (N_5589,N_4595,N_4915);
nand U5590 (N_5590,N_4564,N_4400);
or U5591 (N_5591,N_4776,N_4798);
or U5592 (N_5592,N_4272,N_4579);
xor U5593 (N_5593,N_4688,N_4320);
nand U5594 (N_5594,N_4676,N_4245);
xnor U5595 (N_5595,N_4556,N_4071);
nand U5596 (N_5596,N_4315,N_4620);
nor U5597 (N_5597,N_4669,N_4139);
xnor U5598 (N_5598,N_4973,N_4429);
xor U5599 (N_5599,N_4426,N_4292);
nor U5600 (N_5600,N_4696,N_4744);
and U5601 (N_5601,N_4336,N_4922);
and U5602 (N_5602,N_4547,N_4123);
and U5603 (N_5603,N_4337,N_4467);
or U5604 (N_5604,N_4907,N_4598);
or U5605 (N_5605,N_4346,N_4158);
xnor U5606 (N_5606,N_4257,N_4785);
xor U5607 (N_5607,N_4285,N_4978);
nand U5608 (N_5608,N_4400,N_4277);
nand U5609 (N_5609,N_4100,N_4566);
xnor U5610 (N_5610,N_4236,N_4114);
and U5611 (N_5611,N_4089,N_4665);
nor U5612 (N_5612,N_4390,N_4783);
nand U5613 (N_5613,N_4793,N_4764);
nand U5614 (N_5614,N_4507,N_4320);
nand U5615 (N_5615,N_4576,N_4501);
nand U5616 (N_5616,N_4627,N_4669);
or U5617 (N_5617,N_4631,N_4397);
nand U5618 (N_5618,N_4236,N_4153);
nand U5619 (N_5619,N_4780,N_4402);
nand U5620 (N_5620,N_4299,N_4468);
xor U5621 (N_5621,N_4925,N_4836);
nand U5622 (N_5622,N_4588,N_4923);
nand U5623 (N_5623,N_4027,N_4437);
nor U5624 (N_5624,N_4212,N_4853);
nand U5625 (N_5625,N_4545,N_4985);
xor U5626 (N_5626,N_4982,N_4343);
or U5627 (N_5627,N_4380,N_4987);
xor U5628 (N_5628,N_4846,N_4346);
and U5629 (N_5629,N_4424,N_4181);
xor U5630 (N_5630,N_4858,N_4874);
nand U5631 (N_5631,N_4567,N_4164);
nor U5632 (N_5632,N_4693,N_4612);
xnor U5633 (N_5633,N_4397,N_4896);
nand U5634 (N_5634,N_4907,N_4501);
nor U5635 (N_5635,N_4132,N_4327);
nor U5636 (N_5636,N_4299,N_4477);
xor U5637 (N_5637,N_4150,N_4140);
nand U5638 (N_5638,N_4237,N_4944);
or U5639 (N_5639,N_4636,N_4437);
nor U5640 (N_5640,N_4225,N_4388);
or U5641 (N_5641,N_4979,N_4095);
or U5642 (N_5642,N_4212,N_4614);
or U5643 (N_5643,N_4236,N_4641);
and U5644 (N_5644,N_4310,N_4791);
or U5645 (N_5645,N_4414,N_4330);
and U5646 (N_5646,N_4319,N_4808);
nand U5647 (N_5647,N_4936,N_4380);
nand U5648 (N_5648,N_4483,N_4721);
xor U5649 (N_5649,N_4728,N_4703);
xor U5650 (N_5650,N_4684,N_4791);
or U5651 (N_5651,N_4660,N_4055);
nor U5652 (N_5652,N_4356,N_4818);
nand U5653 (N_5653,N_4932,N_4095);
and U5654 (N_5654,N_4395,N_4548);
and U5655 (N_5655,N_4614,N_4967);
nand U5656 (N_5656,N_4040,N_4998);
xor U5657 (N_5657,N_4222,N_4364);
nor U5658 (N_5658,N_4079,N_4185);
xor U5659 (N_5659,N_4023,N_4468);
and U5660 (N_5660,N_4077,N_4740);
nand U5661 (N_5661,N_4138,N_4356);
xnor U5662 (N_5662,N_4096,N_4357);
and U5663 (N_5663,N_4469,N_4602);
xnor U5664 (N_5664,N_4150,N_4945);
nor U5665 (N_5665,N_4460,N_4542);
or U5666 (N_5666,N_4449,N_4248);
or U5667 (N_5667,N_4855,N_4788);
and U5668 (N_5668,N_4910,N_4132);
and U5669 (N_5669,N_4919,N_4228);
nand U5670 (N_5670,N_4996,N_4505);
xor U5671 (N_5671,N_4034,N_4113);
and U5672 (N_5672,N_4171,N_4677);
nor U5673 (N_5673,N_4542,N_4139);
or U5674 (N_5674,N_4216,N_4903);
and U5675 (N_5675,N_4612,N_4888);
xnor U5676 (N_5676,N_4614,N_4861);
nor U5677 (N_5677,N_4551,N_4637);
and U5678 (N_5678,N_4793,N_4543);
xnor U5679 (N_5679,N_4863,N_4974);
or U5680 (N_5680,N_4746,N_4570);
nor U5681 (N_5681,N_4396,N_4460);
and U5682 (N_5682,N_4836,N_4652);
and U5683 (N_5683,N_4613,N_4153);
nand U5684 (N_5684,N_4529,N_4758);
or U5685 (N_5685,N_4616,N_4595);
or U5686 (N_5686,N_4643,N_4664);
xor U5687 (N_5687,N_4770,N_4920);
and U5688 (N_5688,N_4261,N_4299);
or U5689 (N_5689,N_4419,N_4092);
and U5690 (N_5690,N_4753,N_4489);
xnor U5691 (N_5691,N_4718,N_4651);
and U5692 (N_5692,N_4457,N_4746);
and U5693 (N_5693,N_4452,N_4517);
or U5694 (N_5694,N_4825,N_4238);
and U5695 (N_5695,N_4636,N_4606);
nand U5696 (N_5696,N_4098,N_4674);
and U5697 (N_5697,N_4526,N_4750);
or U5698 (N_5698,N_4836,N_4728);
and U5699 (N_5699,N_4848,N_4539);
and U5700 (N_5700,N_4249,N_4421);
xor U5701 (N_5701,N_4690,N_4192);
nor U5702 (N_5702,N_4629,N_4536);
nand U5703 (N_5703,N_4719,N_4645);
nand U5704 (N_5704,N_4137,N_4208);
and U5705 (N_5705,N_4905,N_4154);
xnor U5706 (N_5706,N_4058,N_4263);
and U5707 (N_5707,N_4499,N_4415);
nand U5708 (N_5708,N_4902,N_4513);
nor U5709 (N_5709,N_4902,N_4674);
and U5710 (N_5710,N_4265,N_4982);
and U5711 (N_5711,N_4728,N_4989);
nand U5712 (N_5712,N_4004,N_4321);
and U5713 (N_5713,N_4528,N_4690);
and U5714 (N_5714,N_4625,N_4258);
or U5715 (N_5715,N_4081,N_4127);
nor U5716 (N_5716,N_4487,N_4936);
xnor U5717 (N_5717,N_4048,N_4799);
xnor U5718 (N_5718,N_4688,N_4345);
and U5719 (N_5719,N_4137,N_4729);
or U5720 (N_5720,N_4285,N_4825);
or U5721 (N_5721,N_4596,N_4903);
nand U5722 (N_5722,N_4180,N_4600);
nor U5723 (N_5723,N_4238,N_4419);
and U5724 (N_5724,N_4772,N_4199);
or U5725 (N_5725,N_4545,N_4050);
and U5726 (N_5726,N_4653,N_4801);
nand U5727 (N_5727,N_4991,N_4579);
nor U5728 (N_5728,N_4241,N_4018);
nor U5729 (N_5729,N_4076,N_4540);
xor U5730 (N_5730,N_4351,N_4716);
nand U5731 (N_5731,N_4170,N_4033);
xor U5732 (N_5732,N_4307,N_4453);
and U5733 (N_5733,N_4406,N_4728);
nand U5734 (N_5734,N_4511,N_4219);
and U5735 (N_5735,N_4369,N_4330);
or U5736 (N_5736,N_4996,N_4584);
and U5737 (N_5737,N_4049,N_4824);
xor U5738 (N_5738,N_4881,N_4514);
nand U5739 (N_5739,N_4716,N_4794);
nor U5740 (N_5740,N_4268,N_4178);
nor U5741 (N_5741,N_4683,N_4742);
nand U5742 (N_5742,N_4186,N_4397);
xor U5743 (N_5743,N_4557,N_4686);
xor U5744 (N_5744,N_4261,N_4861);
and U5745 (N_5745,N_4459,N_4657);
or U5746 (N_5746,N_4779,N_4572);
nand U5747 (N_5747,N_4076,N_4774);
or U5748 (N_5748,N_4146,N_4744);
nand U5749 (N_5749,N_4101,N_4169);
nand U5750 (N_5750,N_4274,N_4606);
nand U5751 (N_5751,N_4499,N_4925);
xor U5752 (N_5752,N_4514,N_4437);
nand U5753 (N_5753,N_4281,N_4548);
or U5754 (N_5754,N_4822,N_4631);
or U5755 (N_5755,N_4205,N_4500);
or U5756 (N_5756,N_4306,N_4082);
and U5757 (N_5757,N_4143,N_4832);
nand U5758 (N_5758,N_4193,N_4166);
nand U5759 (N_5759,N_4013,N_4330);
and U5760 (N_5760,N_4764,N_4445);
nor U5761 (N_5761,N_4576,N_4674);
nand U5762 (N_5762,N_4219,N_4607);
nor U5763 (N_5763,N_4681,N_4027);
and U5764 (N_5764,N_4849,N_4672);
xor U5765 (N_5765,N_4857,N_4152);
xnor U5766 (N_5766,N_4213,N_4669);
xnor U5767 (N_5767,N_4481,N_4234);
xnor U5768 (N_5768,N_4278,N_4220);
nor U5769 (N_5769,N_4240,N_4820);
nor U5770 (N_5770,N_4775,N_4801);
nor U5771 (N_5771,N_4152,N_4847);
and U5772 (N_5772,N_4699,N_4992);
nor U5773 (N_5773,N_4555,N_4833);
nor U5774 (N_5774,N_4982,N_4852);
nand U5775 (N_5775,N_4301,N_4900);
nand U5776 (N_5776,N_4653,N_4108);
or U5777 (N_5777,N_4308,N_4460);
xor U5778 (N_5778,N_4670,N_4787);
nand U5779 (N_5779,N_4998,N_4646);
xnor U5780 (N_5780,N_4834,N_4345);
or U5781 (N_5781,N_4495,N_4483);
nor U5782 (N_5782,N_4369,N_4922);
nand U5783 (N_5783,N_4869,N_4653);
or U5784 (N_5784,N_4705,N_4682);
and U5785 (N_5785,N_4929,N_4011);
and U5786 (N_5786,N_4602,N_4252);
xnor U5787 (N_5787,N_4679,N_4039);
or U5788 (N_5788,N_4771,N_4497);
nand U5789 (N_5789,N_4990,N_4575);
and U5790 (N_5790,N_4784,N_4172);
and U5791 (N_5791,N_4517,N_4822);
xor U5792 (N_5792,N_4781,N_4935);
and U5793 (N_5793,N_4945,N_4324);
xor U5794 (N_5794,N_4962,N_4111);
xor U5795 (N_5795,N_4100,N_4937);
nand U5796 (N_5796,N_4852,N_4135);
and U5797 (N_5797,N_4445,N_4536);
and U5798 (N_5798,N_4652,N_4997);
and U5799 (N_5799,N_4687,N_4717);
nor U5800 (N_5800,N_4589,N_4033);
xnor U5801 (N_5801,N_4090,N_4648);
xnor U5802 (N_5802,N_4424,N_4554);
nand U5803 (N_5803,N_4742,N_4854);
and U5804 (N_5804,N_4444,N_4677);
or U5805 (N_5805,N_4197,N_4070);
xnor U5806 (N_5806,N_4483,N_4443);
or U5807 (N_5807,N_4233,N_4568);
and U5808 (N_5808,N_4495,N_4656);
and U5809 (N_5809,N_4099,N_4748);
or U5810 (N_5810,N_4478,N_4522);
and U5811 (N_5811,N_4527,N_4813);
and U5812 (N_5812,N_4290,N_4649);
nand U5813 (N_5813,N_4637,N_4459);
and U5814 (N_5814,N_4317,N_4691);
nor U5815 (N_5815,N_4239,N_4812);
nand U5816 (N_5816,N_4995,N_4283);
xor U5817 (N_5817,N_4508,N_4869);
and U5818 (N_5818,N_4606,N_4228);
or U5819 (N_5819,N_4859,N_4941);
or U5820 (N_5820,N_4463,N_4769);
xnor U5821 (N_5821,N_4272,N_4895);
and U5822 (N_5822,N_4842,N_4568);
nand U5823 (N_5823,N_4910,N_4187);
xnor U5824 (N_5824,N_4927,N_4987);
and U5825 (N_5825,N_4504,N_4931);
or U5826 (N_5826,N_4198,N_4869);
or U5827 (N_5827,N_4078,N_4668);
xnor U5828 (N_5828,N_4869,N_4190);
nor U5829 (N_5829,N_4305,N_4584);
nor U5830 (N_5830,N_4703,N_4081);
nand U5831 (N_5831,N_4002,N_4520);
and U5832 (N_5832,N_4444,N_4224);
xor U5833 (N_5833,N_4886,N_4118);
or U5834 (N_5834,N_4567,N_4625);
nand U5835 (N_5835,N_4387,N_4463);
nor U5836 (N_5836,N_4599,N_4385);
nor U5837 (N_5837,N_4974,N_4144);
nand U5838 (N_5838,N_4604,N_4838);
nand U5839 (N_5839,N_4336,N_4929);
xnor U5840 (N_5840,N_4538,N_4464);
nor U5841 (N_5841,N_4222,N_4173);
nor U5842 (N_5842,N_4015,N_4475);
and U5843 (N_5843,N_4740,N_4397);
or U5844 (N_5844,N_4311,N_4474);
xor U5845 (N_5845,N_4830,N_4755);
nand U5846 (N_5846,N_4850,N_4954);
nor U5847 (N_5847,N_4901,N_4680);
nor U5848 (N_5848,N_4627,N_4969);
and U5849 (N_5849,N_4183,N_4731);
nor U5850 (N_5850,N_4105,N_4034);
nor U5851 (N_5851,N_4700,N_4068);
and U5852 (N_5852,N_4341,N_4767);
nor U5853 (N_5853,N_4144,N_4929);
nand U5854 (N_5854,N_4949,N_4505);
or U5855 (N_5855,N_4716,N_4918);
or U5856 (N_5856,N_4044,N_4246);
or U5857 (N_5857,N_4997,N_4380);
nor U5858 (N_5858,N_4456,N_4029);
nand U5859 (N_5859,N_4166,N_4606);
or U5860 (N_5860,N_4139,N_4038);
or U5861 (N_5861,N_4356,N_4013);
and U5862 (N_5862,N_4856,N_4317);
nor U5863 (N_5863,N_4731,N_4846);
nand U5864 (N_5864,N_4383,N_4611);
nand U5865 (N_5865,N_4979,N_4343);
nand U5866 (N_5866,N_4384,N_4447);
or U5867 (N_5867,N_4284,N_4092);
nor U5868 (N_5868,N_4127,N_4551);
nor U5869 (N_5869,N_4924,N_4025);
nor U5870 (N_5870,N_4127,N_4118);
nand U5871 (N_5871,N_4161,N_4929);
nand U5872 (N_5872,N_4420,N_4728);
nand U5873 (N_5873,N_4873,N_4339);
and U5874 (N_5874,N_4099,N_4242);
or U5875 (N_5875,N_4090,N_4943);
and U5876 (N_5876,N_4563,N_4645);
nand U5877 (N_5877,N_4241,N_4683);
nand U5878 (N_5878,N_4170,N_4566);
xor U5879 (N_5879,N_4553,N_4023);
nand U5880 (N_5880,N_4797,N_4120);
or U5881 (N_5881,N_4684,N_4472);
or U5882 (N_5882,N_4259,N_4056);
or U5883 (N_5883,N_4855,N_4524);
or U5884 (N_5884,N_4766,N_4894);
nand U5885 (N_5885,N_4321,N_4857);
and U5886 (N_5886,N_4614,N_4503);
or U5887 (N_5887,N_4817,N_4857);
nand U5888 (N_5888,N_4106,N_4908);
nand U5889 (N_5889,N_4374,N_4440);
xor U5890 (N_5890,N_4058,N_4522);
nor U5891 (N_5891,N_4681,N_4824);
nor U5892 (N_5892,N_4348,N_4362);
nor U5893 (N_5893,N_4785,N_4261);
or U5894 (N_5894,N_4306,N_4760);
or U5895 (N_5895,N_4682,N_4346);
and U5896 (N_5896,N_4505,N_4501);
nand U5897 (N_5897,N_4466,N_4100);
xor U5898 (N_5898,N_4423,N_4096);
nor U5899 (N_5899,N_4832,N_4921);
xnor U5900 (N_5900,N_4733,N_4504);
and U5901 (N_5901,N_4229,N_4533);
nor U5902 (N_5902,N_4605,N_4127);
nor U5903 (N_5903,N_4703,N_4540);
nand U5904 (N_5904,N_4938,N_4203);
nand U5905 (N_5905,N_4410,N_4678);
or U5906 (N_5906,N_4093,N_4426);
nand U5907 (N_5907,N_4345,N_4525);
and U5908 (N_5908,N_4320,N_4963);
and U5909 (N_5909,N_4801,N_4232);
and U5910 (N_5910,N_4627,N_4637);
nor U5911 (N_5911,N_4813,N_4193);
and U5912 (N_5912,N_4378,N_4836);
nand U5913 (N_5913,N_4353,N_4294);
or U5914 (N_5914,N_4950,N_4565);
or U5915 (N_5915,N_4806,N_4616);
xnor U5916 (N_5916,N_4490,N_4298);
nand U5917 (N_5917,N_4850,N_4338);
xnor U5918 (N_5918,N_4558,N_4893);
xnor U5919 (N_5919,N_4122,N_4409);
xnor U5920 (N_5920,N_4269,N_4552);
and U5921 (N_5921,N_4476,N_4154);
or U5922 (N_5922,N_4465,N_4446);
xnor U5923 (N_5923,N_4739,N_4122);
or U5924 (N_5924,N_4775,N_4243);
and U5925 (N_5925,N_4650,N_4559);
xor U5926 (N_5926,N_4002,N_4381);
xor U5927 (N_5927,N_4485,N_4125);
nor U5928 (N_5928,N_4040,N_4056);
or U5929 (N_5929,N_4247,N_4955);
and U5930 (N_5930,N_4360,N_4948);
xor U5931 (N_5931,N_4640,N_4306);
xor U5932 (N_5932,N_4703,N_4058);
nor U5933 (N_5933,N_4825,N_4435);
xor U5934 (N_5934,N_4039,N_4608);
and U5935 (N_5935,N_4242,N_4934);
and U5936 (N_5936,N_4958,N_4909);
or U5937 (N_5937,N_4422,N_4974);
or U5938 (N_5938,N_4240,N_4029);
and U5939 (N_5939,N_4339,N_4442);
and U5940 (N_5940,N_4357,N_4943);
and U5941 (N_5941,N_4083,N_4308);
nand U5942 (N_5942,N_4037,N_4056);
or U5943 (N_5943,N_4384,N_4340);
nor U5944 (N_5944,N_4201,N_4800);
and U5945 (N_5945,N_4048,N_4921);
and U5946 (N_5946,N_4304,N_4490);
xnor U5947 (N_5947,N_4399,N_4438);
or U5948 (N_5948,N_4258,N_4688);
nand U5949 (N_5949,N_4876,N_4057);
nor U5950 (N_5950,N_4263,N_4623);
nor U5951 (N_5951,N_4516,N_4551);
xor U5952 (N_5952,N_4372,N_4070);
nor U5953 (N_5953,N_4187,N_4519);
nand U5954 (N_5954,N_4275,N_4550);
nand U5955 (N_5955,N_4459,N_4297);
nor U5956 (N_5956,N_4889,N_4907);
nor U5957 (N_5957,N_4161,N_4663);
or U5958 (N_5958,N_4012,N_4343);
nor U5959 (N_5959,N_4258,N_4113);
nor U5960 (N_5960,N_4441,N_4536);
xnor U5961 (N_5961,N_4518,N_4998);
xnor U5962 (N_5962,N_4071,N_4130);
nand U5963 (N_5963,N_4031,N_4074);
and U5964 (N_5964,N_4308,N_4107);
nand U5965 (N_5965,N_4176,N_4750);
nand U5966 (N_5966,N_4328,N_4093);
nor U5967 (N_5967,N_4540,N_4094);
xor U5968 (N_5968,N_4625,N_4347);
nor U5969 (N_5969,N_4165,N_4792);
nor U5970 (N_5970,N_4406,N_4256);
or U5971 (N_5971,N_4276,N_4518);
or U5972 (N_5972,N_4949,N_4379);
or U5973 (N_5973,N_4342,N_4438);
nor U5974 (N_5974,N_4827,N_4778);
nand U5975 (N_5975,N_4035,N_4164);
xor U5976 (N_5976,N_4775,N_4560);
or U5977 (N_5977,N_4979,N_4945);
xor U5978 (N_5978,N_4153,N_4278);
or U5979 (N_5979,N_4714,N_4440);
or U5980 (N_5980,N_4786,N_4382);
xnor U5981 (N_5981,N_4862,N_4024);
xnor U5982 (N_5982,N_4726,N_4306);
nor U5983 (N_5983,N_4019,N_4569);
nand U5984 (N_5984,N_4186,N_4822);
or U5985 (N_5985,N_4104,N_4749);
or U5986 (N_5986,N_4125,N_4200);
or U5987 (N_5987,N_4141,N_4619);
xor U5988 (N_5988,N_4712,N_4490);
nor U5989 (N_5989,N_4695,N_4246);
or U5990 (N_5990,N_4721,N_4532);
nor U5991 (N_5991,N_4635,N_4309);
nand U5992 (N_5992,N_4970,N_4266);
and U5993 (N_5993,N_4825,N_4838);
nor U5994 (N_5994,N_4006,N_4554);
and U5995 (N_5995,N_4366,N_4558);
nor U5996 (N_5996,N_4018,N_4764);
and U5997 (N_5997,N_4382,N_4599);
or U5998 (N_5998,N_4845,N_4288);
nor U5999 (N_5999,N_4292,N_4224);
nand U6000 (N_6000,N_5921,N_5407);
nor U6001 (N_6001,N_5665,N_5278);
or U6002 (N_6002,N_5668,N_5513);
nand U6003 (N_6003,N_5899,N_5705);
xor U6004 (N_6004,N_5862,N_5515);
nor U6005 (N_6005,N_5678,N_5401);
and U6006 (N_6006,N_5071,N_5775);
or U6007 (N_6007,N_5386,N_5587);
nor U6008 (N_6008,N_5671,N_5545);
nor U6009 (N_6009,N_5510,N_5853);
nand U6010 (N_6010,N_5528,N_5752);
xor U6011 (N_6011,N_5082,N_5747);
xor U6012 (N_6012,N_5025,N_5114);
and U6013 (N_6013,N_5798,N_5660);
and U6014 (N_6014,N_5590,N_5479);
xor U6015 (N_6015,N_5631,N_5723);
nor U6016 (N_6016,N_5319,N_5315);
xor U6017 (N_6017,N_5121,N_5334);
nand U6018 (N_6018,N_5138,N_5179);
nand U6019 (N_6019,N_5928,N_5362);
xor U6020 (N_6020,N_5016,N_5229);
nor U6021 (N_6021,N_5603,N_5007);
nor U6022 (N_6022,N_5271,N_5172);
and U6023 (N_6023,N_5283,N_5640);
nand U6024 (N_6024,N_5583,N_5103);
xor U6025 (N_6025,N_5392,N_5126);
nor U6026 (N_6026,N_5904,N_5262);
xor U6027 (N_6027,N_5874,N_5889);
and U6028 (N_6028,N_5883,N_5284);
nand U6029 (N_6029,N_5553,N_5572);
or U6030 (N_6030,N_5318,N_5035);
or U6031 (N_6031,N_5717,N_5730);
nand U6032 (N_6032,N_5820,N_5537);
or U6033 (N_6033,N_5626,N_5501);
and U6034 (N_6034,N_5194,N_5463);
or U6035 (N_6035,N_5241,N_5586);
or U6036 (N_6036,N_5252,N_5803);
nor U6037 (N_6037,N_5566,N_5959);
or U6038 (N_6038,N_5967,N_5650);
nand U6039 (N_6039,N_5514,N_5689);
nand U6040 (N_6040,N_5378,N_5055);
nor U6041 (N_6041,N_5765,N_5111);
nand U6042 (N_6042,N_5424,N_5696);
and U6043 (N_6043,N_5520,N_5212);
nand U6044 (N_6044,N_5247,N_5502);
nand U6045 (N_6045,N_5589,N_5374);
nor U6046 (N_6046,N_5571,N_5535);
nor U6047 (N_6047,N_5702,N_5246);
or U6048 (N_6048,N_5742,N_5109);
xnor U6049 (N_6049,N_5833,N_5473);
nor U6050 (N_6050,N_5823,N_5302);
or U6051 (N_6051,N_5504,N_5677);
and U6052 (N_6052,N_5654,N_5758);
and U6053 (N_6053,N_5522,N_5734);
or U6054 (N_6054,N_5085,N_5128);
or U6055 (N_6055,N_5037,N_5259);
nand U6056 (N_6056,N_5680,N_5347);
or U6057 (N_6057,N_5153,N_5119);
and U6058 (N_6058,N_5503,N_5321);
or U6059 (N_6059,N_5715,N_5370);
xnor U6060 (N_6060,N_5968,N_5471);
or U6061 (N_6061,N_5089,N_5641);
and U6062 (N_6062,N_5763,N_5682);
nor U6063 (N_6063,N_5711,N_5648);
and U6064 (N_6064,N_5317,N_5215);
nor U6065 (N_6065,N_5716,N_5745);
xnor U6066 (N_6066,N_5203,N_5836);
and U6067 (N_6067,N_5004,N_5686);
and U6068 (N_6068,N_5125,N_5393);
nand U6069 (N_6069,N_5398,N_5530);
nand U6070 (N_6070,N_5040,N_5421);
or U6071 (N_6071,N_5186,N_5365);
nor U6072 (N_6072,N_5301,N_5584);
xor U6073 (N_6073,N_5270,N_5929);
xnor U6074 (N_6074,N_5466,N_5494);
xnor U6075 (N_6075,N_5828,N_5342);
nand U6076 (N_6076,N_5199,N_5244);
xor U6077 (N_6077,N_5253,N_5949);
nand U6078 (N_6078,N_5056,N_5779);
or U6079 (N_6079,N_5913,N_5737);
and U6080 (N_6080,N_5826,N_5307);
nor U6081 (N_6081,N_5916,N_5827);
and U6082 (N_6082,N_5957,N_5699);
and U6083 (N_6083,N_5210,N_5805);
or U6084 (N_6084,N_5002,N_5406);
xor U6085 (N_6085,N_5396,N_5303);
or U6086 (N_6086,N_5695,N_5867);
nand U6087 (N_6087,N_5355,N_5178);
nand U6088 (N_6088,N_5709,N_5546);
nand U6089 (N_6089,N_5997,N_5330);
or U6090 (N_6090,N_5163,N_5389);
and U6091 (N_6091,N_5608,N_5804);
nor U6092 (N_6092,N_5467,N_5456);
or U6093 (N_6093,N_5776,N_5934);
or U6094 (N_6094,N_5982,N_5093);
nor U6095 (N_6095,N_5525,N_5851);
and U6096 (N_6096,N_5847,N_5345);
and U6097 (N_6097,N_5558,N_5011);
nor U6098 (N_6098,N_5840,N_5611);
nand U6099 (N_6099,N_5106,N_5265);
nor U6100 (N_6100,N_5796,N_5969);
and U6101 (N_6101,N_5733,N_5293);
xor U6102 (N_6102,N_5079,N_5996);
and U6103 (N_6103,N_5769,N_5364);
nand U6104 (N_6104,N_5306,N_5003);
nor U6105 (N_6105,N_5906,N_5605);
nand U6106 (N_6106,N_5074,N_5475);
nor U6107 (N_6107,N_5839,N_5896);
nand U6108 (N_6108,N_5816,N_5001);
or U6109 (N_6109,N_5489,N_5991);
or U6110 (N_6110,N_5084,N_5581);
nand U6111 (N_6111,N_5376,N_5073);
and U6112 (N_6112,N_5622,N_5455);
xor U6113 (N_6113,N_5683,N_5846);
xnor U6114 (N_6114,N_5443,N_5653);
and U6115 (N_6115,N_5633,N_5655);
nor U6116 (N_6116,N_5395,N_5998);
and U6117 (N_6117,N_5162,N_5618);
nand U6118 (N_6118,N_5604,N_5094);
nor U6119 (N_6119,N_5459,N_5610);
nor U6120 (N_6120,N_5511,N_5277);
and U6121 (N_6121,N_5445,N_5434);
and U6122 (N_6122,N_5736,N_5615);
xor U6123 (N_6123,N_5329,N_5320);
and U6124 (N_6124,N_5635,N_5684);
or U6125 (N_6125,N_5720,N_5036);
and U6126 (N_6126,N_5010,N_5045);
xnor U6127 (N_6127,N_5166,N_5218);
nor U6128 (N_6128,N_5299,N_5592);
and U6129 (N_6129,N_5136,N_5426);
or U6130 (N_6130,N_5806,N_5978);
or U6131 (N_6131,N_5360,N_5794);
xor U6132 (N_6132,N_5557,N_5623);
nand U6133 (N_6133,N_5612,N_5534);
nor U6134 (N_6134,N_5131,N_5230);
nand U6135 (N_6135,N_5919,N_5613);
or U6136 (N_6136,N_5254,N_5432);
xnor U6137 (N_6137,N_5134,N_5710);
nand U6138 (N_6138,N_5296,N_5966);
nor U6139 (N_6139,N_5047,N_5105);
and U6140 (N_6140,N_5160,N_5243);
nor U6141 (N_6141,N_5273,N_5394);
nand U6142 (N_6142,N_5531,N_5951);
or U6143 (N_6143,N_5038,N_5454);
or U6144 (N_6144,N_5110,N_5795);
and U6145 (N_6145,N_5700,N_5063);
xnor U6146 (N_6146,N_5188,N_5550);
and U6147 (N_6147,N_5076,N_5800);
or U6148 (N_6148,N_5102,N_5529);
or U6149 (N_6149,N_5679,N_5240);
nand U6150 (N_6150,N_5607,N_5909);
nor U6151 (N_6151,N_5481,N_5606);
or U6152 (N_6152,N_5461,N_5880);
xnor U6153 (N_6153,N_5636,N_5390);
nand U6154 (N_6154,N_5656,N_5672);
and U6155 (N_6155,N_5219,N_5113);
xor U6156 (N_6156,N_5349,N_5685);
and U6157 (N_6157,N_5402,N_5280);
xnor U6158 (N_6158,N_5989,N_5182);
xnor U6159 (N_6159,N_5591,N_5044);
xnor U6160 (N_6160,N_5112,N_5888);
nand U6161 (N_6161,N_5895,N_5005);
nor U6162 (N_6162,N_5981,N_5621);
or U6163 (N_6163,N_5143,N_5924);
xnor U6164 (N_6164,N_5980,N_5670);
nand U6165 (N_6165,N_5496,N_5274);
or U6166 (N_6166,N_5070,N_5498);
nor U6167 (N_6167,N_5596,N_5228);
or U6168 (N_6168,N_5869,N_5799);
nor U6169 (N_6169,N_5123,N_5220);
nand U6170 (N_6170,N_5669,N_5115);
nor U6171 (N_6171,N_5863,N_5559);
nand U6172 (N_6172,N_5095,N_5643);
and U6173 (N_6173,N_5400,N_5485);
nand U6174 (N_6174,N_5767,N_5465);
and U6175 (N_6175,N_5645,N_5021);
and U6176 (N_6176,N_5064,N_5328);
nand U6177 (N_6177,N_5915,N_5287);
nand U6178 (N_6178,N_5950,N_5708);
and U6179 (N_6179,N_5420,N_5780);
or U6180 (N_6180,N_5351,N_5956);
nor U6181 (N_6181,N_5857,N_5236);
xor U6182 (N_6182,N_5771,N_5358);
xor U6183 (N_6183,N_5873,N_5910);
nand U6184 (N_6184,N_5474,N_5158);
nor U6185 (N_6185,N_5777,N_5937);
and U6186 (N_6186,N_5524,N_5773);
nor U6187 (N_6187,N_5339,N_5970);
xnor U6188 (N_6188,N_5714,N_5995);
nor U6189 (N_6189,N_5770,N_5092);
or U6190 (N_6190,N_5174,N_5107);
nand U6191 (N_6191,N_5460,N_5782);
nand U6192 (N_6192,N_5728,N_5878);
nor U6193 (N_6193,N_5807,N_5185);
or U6194 (N_6194,N_5974,N_5499);
and U6195 (N_6195,N_5431,N_5724);
xor U6196 (N_6196,N_5681,N_5565);
nand U6197 (N_6197,N_5088,N_5532);
or U6198 (N_6198,N_5411,N_5519);
nor U6199 (N_6199,N_5914,N_5135);
nor U6200 (N_6200,N_5762,N_5784);
nor U6201 (N_6201,N_5601,N_5006);
and U6202 (N_6202,N_5594,N_5316);
or U6203 (N_6203,N_5698,N_5286);
nand U6204 (N_6204,N_5170,N_5920);
nor U6205 (N_6205,N_5870,N_5642);
and U6206 (N_6206,N_5462,N_5427);
nand U6207 (N_6207,N_5740,N_5544);
nor U6208 (N_6208,N_5813,N_5161);
and U6209 (N_6209,N_5834,N_5907);
or U6210 (N_6210,N_5637,N_5054);
nand U6211 (N_6211,N_5041,N_5439);
and U6212 (N_6212,N_5187,N_5117);
nor U6213 (N_6213,N_5447,N_5225);
or U6214 (N_6214,N_5385,N_5688);
or U6215 (N_6215,N_5985,N_5887);
nand U6216 (N_6216,N_5436,N_5130);
xor U6217 (N_6217,N_5925,N_5760);
nor U6218 (N_6218,N_5205,N_5922);
nor U6219 (N_6219,N_5815,N_5190);
and U6220 (N_6220,N_5062,N_5704);
and U6221 (N_6221,N_5333,N_5304);
nand U6222 (N_6222,N_5597,N_5232);
nand U6223 (N_6223,N_5051,N_5894);
or U6224 (N_6224,N_5291,N_5526);
and U6225 (N_6225,N_5940,N_5579);
and U6226 (N_6226,N_5491,N_5375);
nand U6227 (N_6227,N_5211,N_5639);
and U6228 (N_6228,N_5438,N_5990);
or U6229 (N_6229,N_5031,N_5898);
xnor U6230 (N_6230,N_5311,N_5701);
nor U6231 (N_6231,N_5268,N_5100);
or U6232 (N_6232,N_5649,N_5832);
xnor U6233 (N_6233,N_5488,N_5359);
nor U6234 (N_6234,N_5741,N_5150);
nand U6235 (N_6235,N_5842,N_5647);
or U6236 (N_6236,N_5340,N_5790);
xor U6237 (N_6237,N_5221,N_5468);
xnor U6238 (N_6238,N_5120,N_5744);
nand U6239 (N_6239,N_5327,N_5573);
nand U6240 (N_6240,N_5337,N_5024);
xor U6241 (N_6241,N_5946,N_5013);
nor U6242 (N_6242,N_5091,N_5885);
nor U6243 (N_6243,N_5156,N_5541);
nand U6244 (N_6244,N_5059,N_5941);
xor U6245 (N_6245,N_5052,N_5876);
nor U6246 (N_6246,N_5289,N_5948);
and U6247 (N_6247,N_5201,N_5691);
nor U6248 (N_6248,N_5200,N_5387);
or U6249 (N_6249,N_5632,N_5808);
nor U6250 (N_6250,N_5818,N_5487);
xor U6251 (N_6251,N_5255,N_5464);
xor U6252 (N_6252,N_5204,N_5441);
nand U6253 (N_6253,N_5242,N_5954);
or U6254 (N_6254,N_5155,N_5449);
nor U6255 (N_6255,N_5743,N_5066);
nor U6256 (N_6256,N_5727,N_5324);
xnor U6257 (N_6257,N_5458,N_5297);
or U6258 (N_6258,N_5209,N_5585);
and U6259 (N_6259,N_5197,N_5947);
xnor U6260 (N_6260,N_5213,N_5739);
nand U6261 (N_6261,N_5470,N_5020);
nor U6262 (N_6262,N_5480,N_5176);
nor U6263 (N_6263,N_5731,N_5202);
and U6264 (N_6264,N_5933,N_5146);
nand U6265 (N_6265,N_5619,N_5657);
and U6266 (N_6266,N_5602,N_5457);
xnor U6267 (N_6267,N_5101,N_5017);
xnor U6268 (N_6268,N_5167,N_5028);
nor U6269 (N_6269,N_5482,N_5429);
xnor U6270 (N_6270,N_5772,N_5373);
nand U6271 (N_6271,N_5738,N_5858);
and U6272 (N_6272,N_5538,N_5567);
nand U6273 (N_6273,N_5713,N_5658);
nand U6274 (N_6274,N_5331,N_5938);
or U6275 (N_6275,N_5628,N_5835);
nor U6276 (N_6276,N_5415,N_5072);
xor U6277 (N_6277,N_5962,N_5256);
and U6278 (N_6278,N_5931,N_5484);
nor U6279 (N_6279,N_5061,N_5987);
nand U6280 (N_6280,N_5452,N_5509);
xor U6281 (N_6281,N_5893,N_5231);
xor U6282 (N_6282,N_5549,N_5164);
nand U6283 (N_6283,N_5552,N_5570);
or U6284 (N_6284,N_5266,N_5145);
nand U6285 (N_6285,N_5976,N_5450);
nor U6286 (N_6286,N_5152,N_5992);
xnor U6287 (N_6287,N_5226,N_5809);
xor U6288 (N_6288,N_5593,N_5697);
and U6289 (N_6289,N_5298,N_5490);
nor U6290 (N_6290,N_5175,N_5430);
or U6291 (N_6291,N_5646,N_5352);
or U6292 (N_6292,N_5476,N_5864);
or U6293 (N_6293,N_5972,N_5812);
xor U6294 (N_6294,N_5428,N_5718);
or U6295 (N_6295,N_5019,N_5600);
or U6296 (N_6296,N_5032,N_5448);
nor U6297 (N_6297,N_5108,N_5859);
nand U6298 (N_6298,N_5451,N_5217);
xor U6299 (N_6299,N_5446,N_5381);
xnor U6300 (N_6300,N_5801,N_5361);
nand U6301 (N_6301,N_5944,N_5905);
or U6302 (N_6302,N_5569,N_5129);
xnor U6303 (N_6303,N_5027,N_5346);
xor U6304 (N_6304,N_5249,N_5416);
nor U6305 (N_6305,N_5308,N_5932);
xor U6306 (N_6306,N_5159,N_5477);
nand U6307 (N_6307,N_5960,N_5860);
nand U6308 (N_6308,N_5292,N_5788);
nor U6309 (N_6309,N_5638,N_5575);
xnor U6310 (N_6310,N_5761,N_5486);
nand U6311 (N_6311,N_5844,N_5104);
and U6312 (N_6312,N_5667,N_5323);
nor U6313 (N_6313,N_5015,N_5825);
or U6314 (N_6314,N_5322,N_5380);
nor U6315 (N_6315,N_5872,N_5332);
nor U6316 (N_6316,N_5408,N_5759);
xnor U6317 (N_6317,N_5258,N_5263);
or U6318 (N_6318,N_5757,N_5539);
nor U6319 (N_6319,N_5042,N_5151);
or U6320 (N_6320,N_5118,N_5830);
or U6321 (N_6321,N_5177,N_5659);
nand U6322 (N_6322,N_5492,N_5797);
xor U6323 (N_6323,N_5141,N_5372);
xor U6324 (N_6324,N_5171,N_5754);
nand U6325 (N_6325,N_5912,N_5423);
xnor U6326 (N_6326,N_5852,N_5892);
or U6327 (N_6327,N_5096,N_5472);
nor U6328 (N_6328,N_5952,N_5814);
and U6329 (N_6329,N_5831,N_5382);
xnor U6330 (N_6330,N_5282,N_5617);
nand U6331 (N_6331,N_5856,N_5897);
nand U6332 (N_6332,N_5824,N_5943);
xor U6333 (N_6333,N_5314,N_5662);
nand U6334 (N_6334,N_5276,N_5057);
xnor U6335 (N_6335,N_5687,N_5012);
nand U6336 (N_6336,N_5050,N_5144);
and U6337 (N_6337,N_5692,N_5576);
xor U6338 (N_6338,N_5336,N_5865);
xnor U6339 (N_6339,N_5195,N_5994);
nor U6340 (N_6340,N_5674,N_5595);
and U6341 (N_6341,N_5269,N_5341);
nor U6342 (N_6342,N_5305,N_5518);
nand U6343 (N_6343,N_5309,N_5866);
or U6344 (N_6344,N_5453,N_5766);
nor U6345 (N_6345,N_5444,N_5988);
nand U6346 (N_6346,N_5366,N_5644);
xnor U6347 (N_6347,N_5580,N_5180);
and U6348 (N_6348,N_5787,N_5868);
nor U6349 (N_6349,N_5403,N_5192);
nand U6350 (N_6350,N_5900,N_5239);
xor U6351 (N_6351,N_5676,N_5440);
and U6352 (N_6352,N_5122,N_5543);
xnor U6353 (N_6353,N_5555,N_5540);
and U6354 (N_6354,N_5993,N_5902);
nor U6355 (N_6355,N_5384,N_5116);
and U6356 (N_6356,N_5694,N_5248);
and U6357 (N_6357,N_5578,N_5469);
and U6358 (N_6358,N_5478,N_5369);
or U6359 (N_6359,N_5556,N_5207);
or U6360 (N_6360,N_5206,N_5625);
nor U6361 (N_6361,N_5077,N_5942);
xor U6362 (N_6362,N_5986,N_5560);
xor U6363 (N_6363,N_5367,N_5018);
nor U6364 (N_6364,N_5811,N_5245);
xor U6365 (N_6365,N_5624,N_5792);
xor U6366 (N_6366,N_5582,N_5312);
or U6367 (N_6367,N_5058,N_5810);
nor U6368 (N_6368,N_5154,N_5264);
nor U6369 (N_6369,N_5785,N_5417);
nand U6370 (N_6370,N_5442,N_5357);
nor U6371 (N_6371,N_5127,N_5707);
nand U6372 (N_6372,N_5173,N_5999);
and U6373 (N_6373,N_5789,N_5690);
nand U6374 (N_6374,N_5973,N_5124);
or U6375 (N_6375,N_5132,N_5075);
or U6376 (N_6376,N_5497,N_5764);
or U6377 (N_6377,N_5425,N_5325);
xor U6378 (N_6378,N_5845,N_5412);
xnor U6379 (N_6379,N_5009,N_5030);
nand U6380 (N_6380,N_5958,N_5721);
nor U6381 (N_6381,N_5749,N_5008);
xnor U6382 (N_6382,N_5251,N_5848);
and U6383 (N_6383,N_5148,N_5547);
nor U6384 (N_6384,N_5768,N_5379);
nand U6385 (N_6385,N_5719,N_5574);
and U6386 (N_6386,N_5279,N_5261);
nand U6387 (N_6387,N_5078,N_5726);
nand U6388 (N_6388,N_5523,N_5599);
nand U6389 (N_6389,N_5397,N_5908);
xnor U6390 (N_6390,N_5911,N_5965);
nor U6391 (N_6391,N_5554,N_5854);
nand U6392 (N_6392,N_5133,N_5930);
or U6393 (N_6393,N_5879,N_5886);
xnor U6394 (N_6394,N_5551,N_5377);
nand U6395 (N_6395,N_5977,N_5272);
nor U6396 (N_6396,N_5838,N_5026);
nand U6397 (N_6397,N_5196,N_5029);
nor U6398 (N_6398,N_5663,N_5348);
and U6399 (N_6399,N_5413,N_5861);
nor U6400 (N_6400,N_5191,N_5140);
or U6401 (N_6401,N_5053,N_5536);
or U6402 (N_6402,N_5168,N_5495);
nand U6403 (N_6403,N_5043,N_5137);
and U6404 (N_6404,N_5542,N_5193);
xnor U6405 (N_6405,N_5087,N_5198);
nor U6406 (N_6406,N_5984,N_5774);
nor U6407 (N_6407,N_5527,N_5383);
or U6408 (N_6408,N_5802,N_5149);
and U6409 (N_6409,N_5099,N_5652);
and U6410 (N_6410,N_5926,N_5049);
or U6411 (N_6411,N_5285,N_5000);
nand U6412 (N_6412,N_5290,N_5756);
nor U6413 (N_6413,N_5781,N_5048);
or U6414 (N_6414,N_5927,N_5516);
and U6415 (N_6415,N_5791,N_5849);
or U6416 (N_6416,N_5953,N_5598);
nand U6417 (N_6417,N_5500,N_5363);
or U6418 (N_6418,N_5142,N_5353);
nand U6419 (N_6419,N_5275,N_5548);
xnor U6420 (N_6420,N_5616,N_5184);
or U6421 (N_6421,N_5065,N_5356);
nand U6422 (N_6422,N_5732,N_5081);
nand U6423 (N_6423,N_5562,N_5841);
nor U6424 (N_6424,N_5882,N_5399);
nor U6425 (N_6425,N_5183,N_5533);
xnor U6426 (N_6426,N_5961,N_5060);
nor U6427 (N_6427,N_5310,N_5778);
xnor U6428 (N_6428,N_5281,N_5693);
nor U6429 (N_6429,N_5850,N_5414);
or U6430 (N_6430,N_5181,N_5703);
and U6431 (N_6431,N_5368,N_5521);
xnor U6432 (N_6432,N_5344,N_5577);
nor U6433 (N_6433,N_5673,N_5023);
and U6434 (N_6434,N_5214,N_5257);
or U6435 (N_6435,N_5097,N_5409);
xnor U6436 (N_6436,N_5338,N_5661);
or U6437 (N_6437,N_5822,N_5651);
nor U6438 (N_6438,N_5568,N_5169);
xor U6439 (N_6439,N_5725,N_5975);
nand U6440 (N_6440,N_5067,N_5267);
and U6441 (N_6441,N_5493,N_5189);
or U6442 (N_6442,N_5260,N_5234);
and U6443 (N_6443,N_5033,N_5793);
nor U6444 (N_6444,N_5335,N_5294);
and U6445 (N_6445,N_5404,N_5923);
nand U6446 (N_6446,N_5422,N_5901);
or U6447 (N_6447,N_5945,N_5877);
or U6448 (N_6448,N_5080,N_5817);
nor U6449 (N_6449,N_5939,N_5964);
nand U6450 (N_6450,N_5343,N_5222);
or U6451 (N_6451,N_5216,N_5235);
and U6452 (N_6452,N_5620,N_5722);
xnor U6453 (N_6453,N_5371,N_5208);
and U6454 (N_6454,N_5069,N_5735);
or U6455 (N_6455,N_5614,N_5855);
nand U6456 (N_6456,N_5629,N_5391);
nand U6457 (N_6457,N_5675,N_5630);
or U6458 (N_6458,N_5068,N_5588);
and U6459 (N_6459,N_5435,N_5233);
or U6460 (N_6460,N_5890,N_5783);
xnor U6461 (N_6461,N_5300,N_5609);
nor U6462 (N_6462,N_5664,N_5751);
nor U6463 (N_6463,N_5936,N_5837);
xor U6464 (N_6464,N_5821,N_5753);
or U6465 (N_6465,N_5712,N_5437);
xor U6466 (N_6466,N_5634,N_5223);
and U6467 (N_6467,N_5963,N_5917);
xnor U6468 (N_6468,N_5508,N_5083);
nor U6469 (N_6469,N_5561,N_5517);
xor U6470 (N_6470,N_5871,N_5086);
and U6471 (N_6471,N_5729,N_5786);
nand U6472 (N_6472,N_5418,N_5139);
xnor U6473 (N_6473,N_5979,N_5295);
xnor U6474 (N_6474,N_5935,N_5022);
and U6475 (N_6475,N_5955,N_5227);
and U6476 (N_6476,N_5507,N_5090);
or U6477 (N_6477,N_5237,N_5563);
or U6478 (N_6478,N_5627,N_5039);
and U6479 (N_6479,N_5755,N_5238);
xor U6480 (N_6480,N_5881,N_5918);
xnor U6481 (N_6481,N_5748,N_5165);
xnor U6482 (N_6482,N_5875,N_5313);
nand U6483 (N_6483,N_5746,N_5157);
or U6484 (N_6484,N_5354,N_5147);
nand U6485 (N_6485,N_5666,N_5350);
nor U6486 (N_6486,N_5829,N_5505);
and U6487 (N_6487,N_5224,N_5250);
and U6488 (N_6488,N_5706,N_5405);
or U6489 (N_6489,N_5512,N_5971);
nand U6490 (N_6490,N_5388,N_5891);
or U6491 (N_6491,N_5098,N_5326);
nand U6492 (N_6492,N_5819,N_5288);
and U6493 (N_6493,N_5433,N_5843);
and U6494 (N_6494,N_5983,N_5046);
xor U6495 (N_6495,N_5903,N_5884);
or U6496 (N_6496,N_5419,N_5750);
or U6497 (N_6497,N_5014,N_5483);
xnor U6498 (N_6498,N_5034,N_5410);
or U6499 (N_6499,N_5506,N_5564);
and U6500 (N_6500,N_5298,N_5506);
or U6501 (N_6501,N_5823,N_5728);
xnor U6502 (N_6502,N_5544,N_5421);
or U6503 (N_6503,N_5365,N_5087);
xnor U6504 (N_6504,N_5316,N_5788);
xnor U6505 (N_6505,N_5377,N_5825);
nor U6506 (N_6506,N_5092,N_5907);
nand U6507 (N_6507,N_5488,N_5529);
nand U6508 (N_6508,N_5983,N_5151);
nand U6509 (N_6509,N_5226,N_5983);
xor U6510 (N_6510,N_5469,N_5474);
nor U6511 (N_6511,N_5680,N_5717);
or U6512 (N_6512,N_5523,N_5323);
and U6513 (N_6513,N_5574,N_5096);
nor U6514 (N_6514,N_5172,N_5744);
and U6515 (N_6515,N_5692,N_5412);
xor U6516 (N_6516,N_5277,N_5604);
or U6517 (N_6517,N_5866,N_5863);
and U6518 (N_6518,N_5765,N_5070);
xor U6519 (N_6519,N_5184,N_5719);
or U6520 (N_6520,N_5345,N_5553);
or U6521 (N_6521,N_5027,N_5042);
nor U6522 (N_6522,N_5954,N_5602);
or U6523 (N_6523,N_5753,N_5329);
and U6524 (N_6524,N_5870,N_5747);
nand U6525 (N_6525,N_5715,N_5603);
xnor U6526 (N_6526,N_5407,N_5118);
or U6527 (N_6527,N_5484,N_5717);
nand U6528 (N_6528,N_5854,N_5045);
xor U6529 (N_6529,N_5565,N_5268);
and U6530 (N_6530,N_5401,N_5428);
nand U6531 (N_6531,N_5570,N_5885);
or U6532 (N_6532,N_5009,N_5296);
nand U6533 (N_6533,N_5242,N_5422);
nor U6534 (N_6534,N_5633,N_5585);
xor U6535 (N_6535,N_5540,N_5410);
nor U6536 (N_6536,N_5417,N_5254);
xor U6537 (N_6537,N_5612,N_5010);
or U6538 (N_6538,N_5018,N_5345);
or U6539 (N_6539,N_5983,N_5826);
xor U6540 (N_6540,N_5316,N_5384);
nand U6541 (N_6541,N_5389,N_5208);
nor U6542 (N_6542,N_5167,N_5088);
or U6543 (N_6543,N_5177,N_5571);
nand U6544 (N_6544,N_5703,N_5826);
nor U6545 (N_6545,N_5177,N_5055);
xor U6546 (N_6546,N_5513,N_5457);
xnor U6547 (N_6547,N_5445,N_5973);
and U6548 (N_6548,N_5332,N_5478);
and U6549 (N_6549,N_5930,N_5044);
nor U6550 (N_6550,N_5486,N_5001);
and U6551 (N_6551,N_5717,N_5708);
nor U6552 (N_6552,N_5643,N_5088);
nand U6553 (N_6553,N_5245,N_5130);
nor U6554 (N_6554,N_5892,N_5508);
nor U6555 (N_6555,N_5584,N_5641);
and U6556 (N_6556,N_5590,N_5251);
and U6557 (N_6557,N_5654,N_5593);
xnor U6558 (N_6558,N_5114,N_5742);
nand U6559 (N_6559,N_5177,N_5387);
nor U6560 (N_6560,N_5510,N_5454);
or U6561 (N_6561,N_5144,N_5596);
and U6562 (N_6562,N_5007,N_5240);
and U6563 (N_6563,N_5658,N_5211);
nor U6564 (N_6564,N_5365,N_5073);
nand U6565 (N_6565,N_5018,N_5390);
nand U6566 (N_6566,N_5818,N_5595);
xor U6567 (N_6567,N_5093,N_5747);
and U6568 (N_6568,N_5302,N_5583);
and U6569 (N_6569,N_5069,N_5405);
and U6570 (N_6570,N_5578,N_5294);
nand U6571 (N_6571,N_5761,N_5169);
nor U6572 (N_6572,N_5479,N_5255);
nand U6573 (N_6573,N_5588,N_5263);
nor U6574 (N_6574,N_5233,N_5052);
or U6575 (N_6575,N_5763,N_5822);
nand U6576 (N_6576,N_5442,N_5980);
and U6577 (N_6577,N_5664,N_5762);
and U6578 (N_6578,N_5724,N_5335);
and U6579 (N_6579,N_5853,N_5569);
nand U6580 (N_6580,N_5203,N_5903);
or U6581 (N_6581,N_5504,N_5789);
nand U6582 (N_6582,N_5081,N_5860);
or U6583 (N_6583,N_5697,N_5692);
and U6584 (N_6584,N_5423,N_5950);
nand U6585 (N_6585,N_5862,N_5062);
and U6586 (N_6586,N_5610,N_5893);
nor U6587 (N_6587,N_5919,N_5609);
nor U6588 (N_6588,N_5916,N_5389);
nand U6589 (N_6589,N_5687,N_5485);
or U6590 (N_6590,N_5395,N_5343);
and U6591 (N_6591,N_5896,N_5502);
nand U6592 (N_6592,N_5277,N_5725);
xor U6593 (N_6593,N_5868,N_5532);
nand U6594 (N_6594,N_5041,N_5435);
xnor U6595 (N_6595,N_5240,N_5281);
and U6596 (N_6596,N_5225,N_5491);
or U6597 (N_6597,N_5256,N_5392);
xnor U6598 (N_6598,N_5087,N_5052);
xor U6599 (N_6599,N_5618,N_5605);
nor U6600 (N_6600,N_5464,N_5805);
and U6601 (N_6601,N_5992,N_5998);
nor U6602 (N_6602,N_5158,N_5967);
or U6603 (N_6603,N_5185,N_5279);
nand U6604 (N_6604,N_5395,N_5368);
xnor U6605 (N_6605,N_5702,N_5877);
nor U6606 (N_6606,N_5348,N_5197);
and U6607 (N_6607,N_5204,N_5136);
and U6608 (N_6608,N_5162,N_5289);
or U6609 (N_6609,N_5837,N_5972);
or U6610 (N_6610,N_5373,N_5590);
nor U6611 (N_6611,N_5312,N_5716);
and U6612 (N_6612,N_5143,N_5565);
nor U6613 (N_6613,N_5166,N_5329);
nor U6614 (N_6614,N_5718,N_5074);
and U6615 (N_6615,N_5260,N_5940);
or U6616 (N_6616,N_5974,N_5298);
nor U6617 (N_6617,N_5128,N_5419);
nor U6618 (N_6618,N_5554,N_5216);
or U6619 (N_6619,N_5468,N_5641);
xnor U6620 (N_6620,N_5304,N_5749);
or U6621 (N_6621,N_5427,N_5579);
nand U6622 (N_6622,N_5043,N_5164);
and U6623 (N_6623,N_5763,N_5043);
and U6624 (N_6624,N_5949,N_5484);
nor U6625 (N_6625,N_5135,N_5051);
nor U6626 (N_6626,N_5929,N_5504);
nand U6627 (N_6627,N_5912,N_5375);
and U6628 (N_6628,N_5223,N_5612);
nand U6629 (N_6629,N_5104,N_5979);
xnor U6630 (N_6630,N_5111,N_5262);
nand U6631 (N_6631,N_5454,N_5364);
nand U6632 (N_6632,N_5695,N_5333);
and U6633 (N_6633,N_5182,N_5702);
or U6634 (N_6634,N_5608,N_5533);
or U6635 (N_6635,N_5961,N_5467);
or U6636 (N_6636,N_5055,N_5272);
nor U6637 (N_6637,N_5161,N_5163);
nor U6638 (N_6638,N_5499,N_5649);
nor U6639 (N_6639,N_5262,N_5374);
or U6640 (N_6640,N_5983,N_5159);
xor U6641 (N_6641,N_5215,N_5007);
or U6642 (N_6642,N_5234,N_5232);
and U6643 (N_6643,N_5623,N_5417);
or U6644 (N_6644,N_5252,N_5061);
xor U6645 (N_6645,N_5238,N_5955);
and U6646 (N_6646,N_5895,N_5938);
nand U6647 (N_6647,N_5917,N_5636);
nand U6648 (N_6648,N_5038,N_5864);
xor U6649 (N_6649,N_5080,N_5522);
nand U6650 (N_6650,N_5138,N_5533);
nor U6651 (N_6651,N_5177,N_5520);
xor U6652 (N_6652,N_5346,N_5052);
xor U6653 (N_6653,N_5636,N_5710);
nor U6654 (N_6654,N_5056,N_5900);
or U6655 (N_6655,N_5582,N_5436);
nand U6656 (N_6656,N_5189,N_5854);
or U6657 (N_6657,N_5070,N_5222);
or U6658 (N_6658,N_5041,N_5921);
or U6659 (N_6659,N_5572,N_5622);
or U6660 (N_6660,N_5451,N_5948);
xor U6661 (N_6661,N_5114,N_5766);
xor U6662 (N_6662,N_5050,N_5128);
nor U6663 (N_6663,N_5967,N_5677);
nand U6664 (N_6664,N_5205,N_5204);
and U6665 (N_6665,N_5769,N_5792);
nor U6666 (N_6666,N_5903,N_5771);
nand U6667 (N_6667,N_5064,N_5048);
or U6668 (N_6668,N_5413,N_5333);
nand U6669 (N_6669,N_5491,N_5498);
nand U6670 (N_6670,N_5819,N_5215);
xnor U6671 (N_6671,N_5861,N_5612);
or U6672 (N_6672,N_5845,N_5101);
nor U6673 (N_6673,N_5616,N_5600);
or U6674 (N_6674,N_5272,N_5941);
nand U6675 (N_6675,N_5845,N_5337);
or U6676 (N_6676,N_5888,N_5620);
or U6677 (N_6677,N_5109,N_5913);
or U6678 (N_6678,N_5978,N_5506);
nor U6679 (N_6679,N_5242,N_5562);
or U6680 (N_6680,N_5043,N_5548);
nor U6681 (N_6681,N_5396,N_5078);
or U6682 (N_6682,N_5419,N_5820);
and U6683 (N_6683,N_5422,N_5367);
nand U6684 (N_6684,N_5969,N_5054);
or U6685 (N_6685,N_5618,N_5896);
and U6686 (N_6686,N_5090,N_5616);
nand U6687 (N_6687,N_5506,N_5821);
nor U6688 (N_6688,N_5860,N_5759);
and U6689 (N_6689,N_5242,N_5955);
nor U6690 (N_6690,N_5149,N_5484);
and U6691 (N_6691,N_5547,N_5351);
xor U6692 (N_6692,N_5117,N_5470);
nand U6693 (N_6693,N_5672,N_5938);
xnor U6694 (N_6694,N_5912,N_5304);
nor U6695 (N_6695,N_5500,N_5543);
nor U6696 (N_6696,N_5951,N_5948);
and U6697 (N_6697,N_5495,N_5512);
and U6698 (N_6698,N_5586,N_5538);
or U6699 (N_6699,N_5535,N_5686);
nor U6700 (N_6700,N_5065,N_5590);
xor U6701 (N_6701,N_5418,N_5760);
or U6702 (N_6702,N_5348,N_5096);
nor U6703 (N_6703,N_5226,N_5175);
xnor U6704 (N_6704,N_5325,N_5788);
and U6705 (N_6705,N_5168,N_5596);
and U6706 (N_6706,N_5375,N_5740);
xnor U6707 (N_6707,N_5664,N_5611);
nor U6708 (N_6708,N_5355,N_5945);
nor U6709 (N_6709,N_5011,N_5009);
xnor U6710 (N_6710,N_5044,N_5882);
or U6711 (N_6711,N_5044,N_5342);
xnor U6712 (N_6712,N_5947,N_5575);
nor U6713 (N_6713,N_5780,N_5259);
and U6714 (N_6714,N_5546,N_5425);
xor U6715 (N_6715,N_5154,N_5480);
and U6716 (N_6716,N_5389,N_5573);
or U6717 (N_6717,N_5174,N_5705);
and U6718 (N_6718,N_5062,N_5782);
and U6719 (N_6719,N_5562,N_5367);
or U6720 (N_6720,N_5516,N_5186);
nand U6721 (N_6721,N_5502,N_5622);
nand U6722 (N_6722,N_5789,N_5105);
and U6723 (N_6723,N_5023,N_5997);
xor U6724 (N_6724,N_5335,N_5343);
xnor U6725 (N_6725,N_5032,N_5997);
or U6726 (N_6726,N_5099,N_5952);
xnor U6727 (N_6727,N_5530,N_5340);
or U6728 (N_6728,N_5332,N_5532);
xnor U6729 (N_6729,N_5675,N_5429);
or U6730 (N_6730,N_5639,N_5057);
nor U6731 (N_6731,N_5939,N_5773);
or U6732 (N_6732,N_5028,N_5186);
xnor U6733 (N_6733,N_5122,N_5290);
nor U6734 (N_6734,N_5490,N_5382);
and U6735 (N_6735,N_5206,N_5459);
nor U6736 (N_6736,N_5764,N_5908);
nor U6737 (N_6737,N_5312,N_5709);
nand U6738 (N_6738,N_5737,N_5945);
xnor U6739 (N_6739,N_5000,N_5178);
and U6740 (N_6740,N_5751,N_5390);
or U6741 (N_6741,N_5584,N_5754);
xor U6742 (N_6742,N_5233,N_5483);
and U6743 (N_6743,N_5633,N_5110);
xnor U6744 (N_6744,N_5734,N_5385);
or U6745 (N_6745,N_5565,N_5525);
nor U6746 (N_6746,N_5480,N_5332);
or U6747 (N_6747,N_5360,N_5711);
and U6748 (N_6748,N_5441,N_5446);
xnor U6749 (N_6749,N_5998,N_5097);
or U6750 (N_6750,N_5725,N_5393);
nor U6751 (N_6751,N_5277,N_5863);
xnor U6752 (N_6752,N_5513,N_5631);
nand U6753 (N_6753,N_5346,N_5457);
nand U6754 (N_6754,N_5275,N_5497);
nand U6755 (N_6755,N_5980,N_5035);
xor U6756 (N_6756,N_5793,N_5669);
xor U6757 (N_6757,N_5933,N_5478);
and U6758 (N_6758,N_5236,N_5366);
and U6759 (N_6759,N_5547,N_5456);
nand U6760 (N_6760,N_5786,N_5972);
nand U6761 (N_6761,N_5085,N_5224);
xor U6762 (N_6762,N_5316,N_5523);
nand U6763 (N_6763,N_5123,N_5813);
nand U6764 (N_6764,N_5603,N_5618);
or U6765 (N_6765,N_5661,N_5808);
and U6766 (N_6766,N_5637,N_5965);
or U6767 (N_6767,N_5026,N_5327);
or U6768 (N_6768,N_5111,N_5976);
nand U6769 (N_6769,N_5534,N_5508);
and U6770 (N_6770,N_5959,N_5162);
nand U6771 (N_6771,N_5781,N_5137);
nand U6772 (N_6772,N_5222,N_5639);
xor U6773 (N_6773,N_5511,N_5466);
or U6774 (N_6774,N_5332,N_5213);
or U6775 (N_6775,N_5283,N_5581);
or U6776 (N_6776,N_5564,N_5472);
or U6777 (N_6777,N_5162,N_5675);
nor U6778 (N_6778,N_5005,N_5556);
and U6779 (N_6779,N_5402,N_5793);
or U6780 (N_6780,N_5456,N_5802);
xor U6781 (N_6781,N_5986,N_5229);
or U6782 (N_6782,N_5015,N_5390);
nand U6783 (N_6783,N_5717,N_5820);
xnor U6784 (N_6784,N_5479,N_5604);
nand U6785 (N_6785,N_5088,N_5259);
nand U6786 (N_6786,N_5885,N_5253);
and U6787 (N_6787,N_5189,N_5691);
or U6788 (N_6788,N_5965,N_5897);
xnor U6789 (N_6789,N_5037,N_5742);
nand U6790 (N_6790,N_5952,N_5491);
nor U6791 (N_6791,N_5415,N_5172);
nand U6792 (N_6792,N_5961,N_5402);
or U6793 (N_6793,N_5060,N_5698);
and U6794 (N_6794,N_5553,N_5258);
nor U6795 (N_6795,N_5237,N_5288);
and U6796 (N_6796,N_5111,N_5982);
nand U6797 (N_6797,N_5173,N_5410);
or U6798 (N_6798,N_5070,N_5425);
xor U6799 (N_6799,N_5225,N_5464);
xnor U6800 (N_6800,N_5412,N_5738);
or U6801 (N_6801,N_5975,N_5417);
or U6802 (N_6802,N_5741,N_5932);
nor U6803 (N_6803,N_5192,N_5164);
or U6804 (N_6804,N_5737,N_5634);
nand U6805 (N_6805,N_5648,N_5366);
and U6806 (N_6806,N_5554,N_5787);
and U6807 (N_6807,N_5398,N_5710);
nand U6808 (N_6808,N_5513,N_5538);
xnor U6809 (N_6809,N_5577,N_5470);
and U6810 (N_6810,N_5384,N_5922);
xor U6811 (N_6811,N_5054,N_5115);
xor U6812 (N_6812,N_5606,N_5963);
xnor U6813 (N_6813,N_5737,N_5982);
and U6814 (N_6814,N_5844,N_5159);
xor U6815 (N_6815,N_5454,N_5390);
xor U6816 (N_6816,N_5507,N_5566);
or U6817 (N_6817,N_5433,N_5226);
and U6818 (N_6818,N_5806,N_5732);
or U6819 (N_6819,N_5940,N_5437);
xnor U6820 (N_6820,N_5491,N_5545);
or U6821 (N_6821,N_5789,N_5209);
or U6822 (N_6822,N_5876,N_5797);
and U6823 (N_6823,N_5961,N_5794);
xnor U6824 (N_6824,N_5407,N_5829);
xor U6825 (N_6825,N_5097,N_5318);
xor U6826 (N_6826,N_5565,N_5462);
or U6827 (N_6827,N_5473,N_5858);
nor U6828 (N_6828,N_5306,N_5696);
nor U6829 (N_6829,N_5130,N_5993);
nand U6830 (N_6830,N_5806,N_5312);
xnor U6831 (N_6831,N_5136,N_5288);
or U6832 (N_6832,N_5235,N_5483);
and U6833 (N_6833,N_5315,N_5603);
xnor U6834 (N_6834,N_5338,N_5059);
xnor U6835 (N_6835,N_5670,N_5256);
or U6836 (N_6836,N_5478,N_5677);
and U6837 (N_6837,N_5248,N_5877);
or U6838 (N_6838,N_5720,N_5849);
and U6839 (N_6839,N_5777,N_5604);
and U6840 (N_6840,N_5657,N_5102);
or U6841 (N_6841,N_5735,N_5255);
nor U6842 (N_6842,N_5958,N_5717);
nor U6843 (N_6843,N_5490,N_5509);
xnor U6844 (N_6844,N_5014,N_5582);
nand U6845 (N_6845,N_5278,N_5196);
nand U6846 (N_6846,N_5014,N_5552);
xor U6847 (N_6847,N_5386,N_5002);
nor U6848 (N_6848,N_5727,N_5222);
and U6849 (N_6849,N_5695,N_5231);
and U6850 (N_6850,N_5738,N_5515);
or U6851 (N_6851,N_5192,N_5486);
xor U6852 (N_6852,N_5856,N_5018);
xnor U6853 (N_6853,N_5994,N_5902);
or U6854 (N_6854,N_5950,N_5923);
or U6855 (N_6855,N_5683,N_5053);
nand U6856 (N_6856,N_5220,N_5862);
nand U6857 (N_6857,N_5797,N_5896);
nor U6858 (N_6858,N_5531,N_5491);
and U6859 (N_6859,N_5714,N_5848);
and U6860 (N_6860,N_5099,N_5643);
and U6861 (N_6861,N_5164,N_5572);
or U6862 (N_6862,N_5865,N_5192);
nor U6863 (N_6863,N_5862,N_5990);
nor U6864 (N_6864,N_5658,N_5908);
and U6865 (N_6865,N_5089,N_5963);
or U6866 (N_6866,N_5525,N_5900);
xnor U6867 (N_6867,N_5163,N_5291);
or U6868 (N_6868,N_5498,N_5164);
and U6869 (N_6869,N_5030,N_5467);
or U6870 (N_6870,N_5995,N_5383);
or U6871 (N_6871,N_5866,N_5020);
nand U6872 (N_6872,N_5132,N_5365);
or U6873 (N_6873,N_5412,N_5977);
or U6874 (N_6874,N_5616,N_5786);
or U6875 (N_6875,N_5470,N_5388);
or U6876 (N_6876,N_5587,N_5695);
and U6877 (N_6877,N_5677,N_5470);
nand U6878 (N_6878,N_5822,N_5409);
xnor U6879 (N_6879,N_5048,N_5791);
or U6880 (N_6880,N_5175,N_5277);
xor U6881 (N_6881,N_5967,N_5165);
or U6882 (N_6882,N_5996,N_5762);
xnor U6883 (N_6883,N_5900,N_5587);
xnor U6884 (N_6884,N_5563,N_5454);
or U6885 (N_6885,N_5720,N_5690);
nand U6886 (N_6886,N_5010,N_5875);
nand U6887 (N_6887,N_5339,N_5038);
nor U6888 (N_6888,N_5993,N_5576);
and U6889 (N_6889,N_5075,N_5439);
or U6890 (N_6890,N_5558,N_5764);
nor U6891 (N_6891,N_5677,N_5723);
xnor U6892 (N_6892,N_5292,N_5602);
or U6893 (N_6893,N_5962,N_5918);
or U6894 (N_6894,N_5426,N_5090);
xor U6895 (N_6895,N_5077,N_5144);
and U6896 (N_6896,N_5423,N_5674);
nor U6897 (N_6897,N_5473,N_5406);
xor U6898 (N_6898,N_5385,N_5559);
or U6899 (N_6899,N_5147,N_5343);
xnor U6900 (N_6900,N_5744,N_5764);
nor U6901 (N_6901,N_5002,N_5433);
nand U6902 (N_6902,N_5026,N_5286);
nand U6903 (N_6903,N_5911,N_5747);
nor U6904 (N_6904,N_5058,N_5659);
and U6905 (N_6905,N_5129,N_5636);
or U6906 (N_6906,N_5394,N_5537);
nor U6907 (N_6907,N_5024,N_5297);
xnor U6908 (N_6908,N_5136,N_5681);
nor U6909 (N_6909,N_5780,N_5877);
nand U6910 (N_6910,N_5919,N_5462);
and U6911 (N_6911,N_5689,N_5399);
nand U6912 (N_6912,N_5600,N_5404);
or U6913 (N_6913,N_5582,N_5251);
or U6914 (N_6914,N_5985,N_5861);
and U6915 (N_6915,N_5993,N_5590);
and U6916 (N_6916,N_5863,N_5040);
xor U6917 (N_6917,N_5848,N_5006);
and U6918 (N_6918,N_5969,N_5790);
xnor U6919 (N_6919,N_5347,N_5297);
nand U6920 (N_6920,N_5356,N_5991);
nor U6921 (N_6921,N_5009,N_5991);
or U6922 (N_6922,N_5742,N_5417);
xor U6923 (N_6923,N_5064,N_5307);
and U6924 (N_6924,N_5201,N_5190);
and U6925 (N_6925,N_5038,N_5769);
or U6926 (N_6926,N_5448,N_5948);
nand U6927 (N_6927,N_5301,N_5780);
or U6928 (N_6928,N_5397,N_5120);
nand U6929 (N_6929,N_5730,N_5642);
nand U6930 (N_6930,N_5047,N_5866);
and U6931 (N_6931,N_5117,N_5532);
and U6932 (N_6932,N_5487,N_5849);
or U6933 (N_6933,N_5957,N_5363);
xor U6934 (N_6934,N_5664,N_5577);
nor U6935 (N_6935,N_5546,N_5492);
or U6936 (N_6936,N_5733,N_5412);
xor U6937 (N_6937,N_5685,N_5960);
nor U6938 (N_6938,N_5092,N_5464);
or U6939 (N_6939,N_5027,N_5112);
nor U6940 (N_6940,N_5251,N_5737);
and U6941 (N_6941,N_5595,N_5063);
xor U6942 (N_6942,N_5976,N_5962);
xor U6943 (N_6943,N_5938,N_5422);
xor U6944 (N_6944,N_5834,N_5553);
and U6945 (N_6945,N_5155,N_5456);
xor U6946 (N_6946,N_5907,N_5819);
or U6947 (N_6947,N_5612,N_5842);
xnor U6948 (N_6948,N_5902,N_5254);
and U6949 (N_6949,N_5340,N_5174);
and U6950 (N_6950,N_5048,N_5482);
and U6951 (N_6951,N_5301,N_5979);
nand U6952 (N_6952,N_5656,N_5671);
and U6953 (N_6953,N_5547,N_5499);
or U6954 (N_6954,N_5640,N_5858);
or U6955 (N_6955,N_5509,N_5052);
xnor U6956 (N_6956,N_5202,N_5746);
xor U6957 (N_6957,N_5268,N_5094);
or U6958 (N_6958,N_5929,N_5555);
and U6959 (N_6959,N_5482,N_5059);
nor U6960 (N_6960,N_5654,N_5312);
or U6961 (N_6961,N_5900,N_5485);
or U6962 (N_6962,N_5515,N_5715);
xor U6963 (N_6963,N_5576,N_5727);
nand U6964 (N_6964,N_5483,N_5822);
or U6965 (N_6965,N_5876,N_5970);
xnor U6966 (N_6966,N_5671,N_5239);
xnor U6967 (N_6967,N_5809,N_5177);
xnor U6968 (N_6968,N_5080,N_5020);
xor U6969 (N_6969,N_5032,N_5291);
and U6970 (N_6970,N_5786,N_5524);
nand U6971 (N_6971,N_5667,N_5787);
or U6972 (N_6972,N_5433,N_5443);
and U6973 (N_6973,N_5033,N_5453);
xor U6974 (N_6974,N_5126,N_5951);
nand U6975 (N_6975,N_5533,N_5846);
and U6976 (N_6976,N_5249,N_5645);
and U6977 (N_6977,N_5956,N_5915);
nand U6978 (N_6978,N_5912,N_5172);
xnor U6979 (N_6979,N_5462,N_5263);
nor U6980 (N_6980,N_5078,N_5664);
or U6981 (N_6981,N_5995,N_5634);
or U6982 (N_6982,N_5088,N_5700);
or U6983 (N_6983,N_5063,N_5873);
xor U6984 (N_6984,N_5530,N_5733);
nor U6985 (N_6985,N_5294,N_5581);
or U6986 (N_6986,N_5234,N_5856);
nor U6987 (N_6987,N_5622,N_5529);
and U6988 (N_6988,N_5906,N_5833);
nand U6989 (N_6989,N_5600,N_5388);
nand U6990 (N_6990,N_5535,N_5122);
nand U6991 (N_6991,N_5073,N_5054);
nand U6992 (N_6992,N_5464,N_5789);
nor U6993 (N_6993,N_5394,N_5947);
xor U6994 (N_6994,N_5732,N_5068);
xor U6995 (N_6995,N_5041,N_5866);
nor U6996 (N_6996,N_5804,N_5816);
xor U6997 (N_6997,N_5642,N_5158);
nor U6998 (N_6998,N_5104,N_5913);
nor U6999 (N_6999,N_5467,N_5673);
and U7000 (N_7000,N_6642,N_6441);
nor U7001 (N_7001,N_6274,N_6883);
or U7002 (N_7002,N_6045,N_6471);
nor U7003 (N_7003,N_6127,N_6941);
xor U7004 (N_7004,N_6726,N_6478);
xor U7005 (N_7005,N_6961,N_6142);
nor U7006 (N_7006,N_6589,N_6493);
nor U7007 (N_7007,N_6149,N_6007);
and U7008 (N_7008,N_6617,N_6359);
nand U7009 (N_7009,N_6430,N_6926);
xnor U7010 (N_7010,N_6998,N_6939);
nor U7011 (N_7011,N_6599,N_6831);
or U7012 (N_7012,N_6345,N_6691);
nand U7013 (N_7013,N_6635,N_6675);
and U7014 (N_7014,N_6191,N_6767);
xor U7015 (N_7015,N_6841,N_6571);
nand U7016 (N_7016,N_6836,N_6062);
xnor U7017 (N_7017,N_6426,N_6550);
nor U7018 (N_7018,N_6111,N_6473);
and U7019 (N_7019,N_6396,N_6777);
or U7020 (N_7020,N_6099,N_6217);
nand U7021 (N_7021,N_6268,N_6079);
and U7022 (N_7022,N_6468,N_6663);
xnor U7023 (N_7023,N_6917,N_6555);
and U7024 (N_7024,N_6188,N_6046);
nor U7025 (N_7025,N_6623,N_6710);
and U7026 (N_7026,N_6826,N_6522);
xnor U7027 (N_7027,N_6202,N_6332);
or U7028 (N_7028,N_6439,N_6338);
and U7029 (N_7029,N_6908,N_6243);
xor U7030 (N_7030,N_6829,N_6198);
nand U7031 (N_7031,N_6795,N_6234);
nor U7032 (N_7032,N_6715,N_6145);
and U7033 (N_7033,N_6669,N_6254);
nor U7034 (N_7034,N_6762,N_6236);
nand U7035 (N_7035,N_6492,N_6641);
and U7036 (N_7036,N_6511,N_6671);
and U7037 (N_7037,N_6108,N_6905);
xnor U7038 (N_7038,N_6933,N_6415);
xor U7039 (N_7039,N_6469,N_6867);
or U7040 (N_7040,N_6739,N_6838);
nor U7041 (N_7041,N_6649,N_6117);
or U7042 (N_7042,N_6516,N_6043);
or U7043 (N_7043,N_6814,N_6624);
nand U7044 (N_7044,N_6030,N_6593);
or U7045 (N_7045,N_6159,N_6660);
nand U7046 (N_7046,N_6993,N_6713);
or U7047 (N_7047,N_6677,N_6432);
nand U7048 (N_7048,N_6152,N_6333);
nand U7049 (N_7049,N_6765,N_6886);
and U7050 (N_7050,N_6971,N_6869);
nand U7051 (N_7051,N_6833,N_6271);
nand U7052 (N_7052,N_6906,N_6056);
xor U7053 (N_7053,N_6741,N_6573);
or U7054 (N_7054,N_6800,N_6832);
xnor U7055 (N_7055,N_6881,N_6900);
and U7056 (N_7056,N_6028,N_6760);
nand U7057 (N_7057,N_6298,N_6358);
xnor U7058 (N_7058,N_6746,N_6651);
xor U7059 (N_7059,N_6125,N_6895);
nand U7060 (N_7060,N_6798,N_6576);
xor U7061 (N_7061,N_6557,N_6411);
xnor U7062 (N_7062,N_6784,N_6343);
or U7063 (N_7063,N_6205,N_6954);
or U7064 (N_7064,N_6627,N_6957);
or U7065 (N_7065,N_6891,N_6199);
or U7066 (N_7066,N_6357,N_6636);
nor U7067 (N_7067,N_6534,N_6040);
and U7068 (N_7068,N_6364,N_6153);
or U7069 (N_7069,N_6779,N_6059);
or U7070 (N_7070,N_6240,N_6248);
xor U7071 (N_7071,N_6082,N_6500);
nand U7072 (N_7072,N_6318,N_6595);
and U7073 (N_7073,N_6950,N_6283);
nand U7074 (N_7074,N_6690,N_6705);
and U7075 (N_7075,N_6857,N_6241);
nor U7076 (N_7076,N_6170,N_6858);
nand U7077 (N_7077,N_6012,N_6928);
or U7078 (N_7078,N_6370,N_6383);
or U7079 (N_7079,N_6786,N_6897);
and U7080 (N_7080,N_6503,N_6376);
nand U7081 (N_7081,N_6309,N_6321);
and U7082 (N_7082,N_6868,N_6233);
xor U7083 (N_7083,N_6618,N_6119);
or U7084 (N_7084,N_6700,N_6899);
and U7085 (N_7085,N_6302,N_6490);
nand U7086 (N_7086,N_6425,N_6808);
nor U7087 (N_7087,N_6583,N_6666);
or U7088 (N_7088,N_6247,N_6614);
and U7089 (N_7089,N_6259,N_6262);
nand U7090 (N_7090,N_6404,N_6440);
nand U7091 (N_7091,N_6398,N_6165);
nor U7092 (N_7092,N_6818,N_6051);
and U7093 (N_7093,N_6619,N_6532);
and U7094 (N_7094,N_6512,N_6066);
and U7095 (N_7095,N_6904,N_6923);
nor U7096 (N_7096,N_6171,N_6050);
xor U7097 (N_7097,N_6434,N_6197);
nor U7098 (N_7098,N_6265,N_6123);
or U7099 (N_7099,N_6437,N_6184);
or U7100 (N_7100,N_6393,N_6982);
nand U7101 (N_7101,N_6355,N_6470);
xnor U7102 (N_7102,N_6385,N_6633);
xor U7103 (N_7103,N_6342,N_6545);
and U7104 (N_7104,N_6179,N_6730);
or U7105 (N_7105,N_6443,N_6284);
and U7106 (N_7106,N_6257,N_6520);
xnor U7107 (N_7107,N_6922,N_6005);
and U7108 (N_7108,N_6166,N_6769);
or U7109 (N_7109,N_6102,N_6055);
nand U7110 (N_7110,N_6572,N_6825);
nor U7111 (N_7111,N_6788,N_6094);
xnor U7112 (N_7112,N_6584,N_6901);
nand U7113 (N_7113,N_6187,N_6547);
nand U7114 (N_7114,N_6266,N_6350);
or U7115 (N_7115,N_6994,N_6965);
nor U7116 (N_7116,N_6960,N_6681);
nand U7117 (N_7117,N_6065,N_6429);
nand U7118 (N_7118,N_6120,N_6275);
nor U7119 (N_7119,N_6602,N_6820);
nor U7120 (N_7120,N_6725,N_6804);
nor U7121 (N_7121,N_6568,N_6272);
and U7122 (N_7122,N_6768,N_6962);
or U7123 (N_7123,N_6027,N_6390);
xor U7124 (N_7124,N_6448,N_6122);
nand U7125 (N_7125,N_6776,N_6421);
and U7126 (N_7126,N_6981,N_6916);
nor U7127 (N_7127,N_6774,N_6112);
xor U7128 (N_7128,N_6626,N_6653);
or U7129 (N_7129,N_6023,N_6016);
or U7130 (N_7130,N_6796,N_6377);
or U7131 (N_7131,N_6173,N_6537);
nand U7132 (N_7132,N_6308,N_6061);
nor U7133 (N_7133,N_6544,N_6577);
or U7134 (N_7134,N_6615,N_6267);
nand U7135 (N_7135,N_6146,N_6920);
and U7136 (N_7136,N_6925,N_6458);
or U7137 (N_7137,N_6356,N_6080);
or U7138 (N_7138,N_6255,N_6387);
nor U7139 (N_7139,N_6608,N_6542);
nor U7140 (N_7140,N_6174,N_6032);
or U7141 (N_7141,N_6201,N_6932);
and U7142 (N_7142,N_6540,N_6766);
or U7143 (N_7143,N_6610,N_6935);
or U7144 (N_7144,N_6348,N_6835);
or U7145 (N_7145,N_6455,N_6505);
and U7146 (N_7146,N_6067,N_6481);
nor U7147 (N_7147,N_6620,N_6562);
xor U7148 (N_7148,N_6854,N_6687);
nand U7149 (N_7149,N_6491,N_6802);
and U7150 (N_7150,N_6222,N_6477);
xnor U7151 (N_7151,N_6015,N_6495);
nand U7152 (N_7152,N_6402,N_6246);
nand U7153 (N_7153,N_6893,N_6116);
xnor U7154 (N_7154,N_6316,N_6890);
nor U7155 (N_7155,N_6462,N_6674);
nor U7156 (N_7156,N_6979,N_6315);
or U7157 (N_7157,N_6987,N_6305);
nand U7158 (N_7158,N_6209,N_6888);
nor U7159 (N_7159,N_6752,N_6931);
nand U7160 (N_7160,N_6031,N_6238);
xnor U7161 (N_7161,N_6380,N_6706);
xor U7162 (N_7162,N_6510,N_6001);
or U7163 (N_7163,N_6162,N_6239);
nand U7164 (N_7164,N_6025,N_6938);
or U7165 (N_7165,N_6499,N_6929);
or U7166 (N_7166,N_6978,N_6852);
nor U7167 (N_7167,N_6183,N_6092);
xnor U7168 (N_7168,N_6704,N_6693);
xor U7169 (N_7169,N_6943,N_6422);
and U7170 (N_7170,N_6919,N_6724);
nor U7171 (N_7171,N_6256,N_6759);
nand U7172 (N_7172,N_6349,N_6328);
xnor U7173 (N_7173,N_6812,N_6264);
nand U7174 (N_7174,N_6639,N_6678);
or U7175 (N_7175,N_6698,N_6394);
and U7176 (N_7176,N_6322,N_6541);
and U7177 (N_7177,N_6090,N_6634);
xnor U7178 (N_7178,N_6719,N_6320);
or U7179 (N_7179,N_6172,N_6083);
or U7180 (N_7180,N_6021,N_6531);
xor U7181 (N_7181,N_6915,N_6995);
nand U7182 (N_7182,N_6294,N_6058);
and U7183 (N_7183,N_6530,N_6223);
xor U7184 (N_7184,N_6974,N_6096);
xor U7185 (N_7185,N_6068,N_6446);
and U7186 (N_7186,N_6772,N_6087);
and U7187 (N_7187,N_6278,N_6151);
or U7188 (N_7188,N_6983,N_6871);
and U7189 (N_7189,N_6399,N_6970);
nand U7190 (N_7190,N_6301,N_6417);
and U7191 (N_7191,N_6386,N_6181);
and U7192 (N_7192,N_6646,N_6819);
xor U7193 (N_7193,N_6594,N_6219);
and U7194 (N_7194,N_6064,N_6753);
or U7195 (N_7195,N_6934,N_6029);
and U7196 (N_7196,N_6466,N_6848);
or U7197 (N_7197,N_6269,N_6996);
or U7198 (N_7198,N_6295,N_6579);
or U7199 (N_7199,N_6228,N_6310);
and U7200 (N_7200,N_6427,N_6770);
xnor U7201 (N_7201,N_6709,N_6980);
and U7202 (N_7202,N_6258,N_6161);
or U7203 (N_7203,N_6940,N_6442);
xor U7204 (N_7204,N_6003,N_6840);
nand U7205 (N_7205,N_6862,N_6740);
and U7206 (N_7206,N_6711,N_6379);
xor U7207 (N_7207,N_6504,N_6086);
or U7208 (N_7208,N_6569,N_6823);
and U7209 (N_7209,N_6176,N_6733);
or U7210 (N_7210,N_6876,N_6720);
or U7211 (N_7211,N_6661,N_6887);
or U7212 (N_7212,N_6323,N_6780);
xor U7213 (N_7213,N_6955,N_6578);
nand U7214 (N_7214,N_6115,N_6643);
nand U7215 (N_7215,N_6699,N_6963);
nand U7216 (N_7216,N_6597,N_6607);
and U7217 (N_7217,N_6375,N_6200);
or U7218 (N_7218,N_6898,N_6910);
nand U7219 (N_7219,N_6793,N_6482);
or U7220 (N_7220,N_6433,N_6894);
and U7221 (N_7221,N_6628,N_6913);
xor U7222 (N_7222,N_6975,N_6076);
or U7223 (N_7223,N_6559,N_6882);
nand U7224 (N_7224,N_6344,N_6889);
nor U7225 (N_7225,N_6276,N_6009);
nor U7226 (N_7226,N_6892,N_6684);
nor U7227 (N_7227,N_6973,N_6590);
nor U7228 (N_7228,N_6985,N_6093);
and U7229 (N_7229,N_6141,N_6231);
nor U7230 (N_7230,N_6324,N_6750);
nor U7231 (N_7231,N_6423,N_6290);
or U7232 (N_7232,N_6736,N_6697);
or U7233 (N_7233,N_6655,N_6834);
or U7234 (N_7234,N_6822,N_6874);
nor U7235 (N_7235,N_6453,N_6790);
or U7236 (N_7236,N_6483,N_6091);
xnor U7237 (N_7237,N_6523,N_6077);
and U7238 (N_7238,N_6103,N_6054);
nor U7239 (N_7239,N_6476,N_6461);
or U7240 (N_7240,N_6797,N_6845);
and U7241 (N_7241,N_6403,N_6743);
nor U7242 (N_7242,N_6964,N_6409);
xor U7243 (N_7243,N_6060,N_6944);
nand U7244 (N_7244,N_6778,N_6870);
nor U7245 (N_7245,N_6033,N_6182);
nand U7246 (N_7246,N_6053,N_6738);
nand U7247 (N_7247,N_6185,N_6539);
nor U7248 (N_7248,N_6273,N_6824);
nor U7249 (N_7249,N_6037,N_6659);
nand U7250 (N_7250,N_6175,N_6177);
xnor U7251 (N_7251,N_6723,N_6878);
xnor U7252 (N_7252,N_6405,N_6853);
nand U7253 (N_7253,N_6407,N_6128);
and U7254 (N_7254,N_6391,N_6992);
nand U7255 (N_7255,N_6519,N_6563);
and U7256 (N_7256,N_6842,N_6137);
xor U7257 (N_7257,N_6914,N_6327);
nor U7258 (N_7258,N_6603,N_6412);
nor U7259 (N_7259,N_6098,N_6810);
nor U7260 (N_7260,N_6416,N_6424);
nor U7261 (N_7261,N_6131,N_6261);
and U7262 (N_7262,N_6606,N_6070);
nand U7263 (N_7263,N_6817,N_6097);
or U7264 (N_7264,N_6279,N_6947);
nor U7265 (N_7265,N_6764,N_6783);
or U7266 (N_7266,N_6121,N_6625);
and U7267 (N_7267,N_6480,N_6196);
or U7268 (N_7268,N_6075,N_6586);
xnor U7269 (N_7269,N_6664,N_6937);
and U7270 (N_7270,N_6160,N_6361);
and U7271 (N_7271,N_6095,N_6968);
nor U7272 (N_7272,N_6558,N_6863);
or U7273 (N_7273,N_6972,N_6803);
nand U7274 (N_7274,N_6263,N_6360);
or U7275 (N_7275,N_6549,N_6525);
xnor U7276 (N_7276,N_6210,N_6341);
and U7277 (N_7277,N_6419,N_6872);
nand U7278 (N_7278,N_6044,N_6002);
xnor U7279 (N_7279,N_6019,N_6648);
xor U7280 (N_7280,N_6336,N_6751);
or U7281 (N_7281,N_6976,N_6670);
or U7282 (N_7282,N_6877,N_6337);
xor U7283 (N_7283,N_6775,N_6211);
or U7284 (N_7284,N_6368,N_6585);
or U7285 (N_7285,N_6745,N_6289);
nor U7286 (N_7286,N_6124,N_6507);
nor U7287 (N_7287,N_6143,N_6132);
nor U7288 (N_7288,N_6156,N_6144);
and U7289 (N_7289,N_6758,N_6304);
nand U7290 (N_7290,N_6846,N_6085);
xor U7291 (N_7291,N_6335,N_6942);
xor U7292 (N_7292,N_6498,N_6331);
and U7293 (N_7293,N_6186,N_6017);
xnor U7294 (N_7294,N_6388,N_6133);
nor U7295 (N_7295,N_6526,N_6456);
and U7296 (N_7296,N_6508,N_6397);
nor U7297 (N_7297,N_6229,N_6673);
nand U7298 (N_7298,N_6130,N_6588);
and U7299 (N_7299,N_6896,N_6856);
nand U7300 (N_7300,N_6712,N_6582);
and U7301 (N_7301,N_6683,N_6249);
nor U7302 (N_7302,N_6297,N_6069);
or U7303 (N_7303,N_6212,N_6296);
and U7304 (N_7304,N_6773,N_6850);
xor U7305 (N_7305,N_6536,N_6638);
xnor U7306 (N_7306,N_6138,N_6300);
or U7307 (N_7307,N_6224,N_6420);
nand U7308 (N_7308,N_6966,N_6849);
or U7309 (N_7309,N_6533,N_6689);
or U7310 (N_7310,N_6564,N_6598);
nand U7311 (N_7311,N_6311,N_6613);
or U7312 (N_7312,N_6809,N_6591);
and U7313 (N_7313,N_6727,N_6821);
and U7314 (N_7314,N_6018,N_6286);
or U7315 (N_7315,N_6629,N_6535);
xnor U7316 (N_7316,N_6517,N_6109);
and U7317 (N_7317,N_6630,N_6215);
nand U7318 (N_7318,N_6190,N_6761);
xnor U7319 (N_7319,N_6662,N_6592);
xor U7320 (N_7320,N_6195,N_6837);
nand U7321 (N_7321,N_6672,N_6918);
or U7322 (N_7322,N_6650,N_6218);
xnor U7323 (N_7323,N_6039,N_6460);
nor U7324 (N_7324,N_6986,N_6688);
and U7325 (N_7325,N_6789,N_6969);
nand U7326 (N_7326,N_6959,N_6155);
and U7327 (N_7327,N_6347,N_6911);
nand U7328 (N_7328,N_6782,N_6365);
nor U7329 (N_7329,N_6363,N_6521);
or U7330 (N_7330,N_6792,N_6253);
or U7331 (N_7331,N_6227,N_6656);
xnor U7332 (N_7332,N_6281,N_6967);
nand U7333 (N_7333,N_6408,N_6884);
and U7334 (N_7334,N_6484,N_6596);
nor U7335 (N_7335,N_6637,N_6885);
nor U7336 (N_7336,N_6047,N_6502);
xor U7337 (N_7337,N_6612,N_6912);
or U7338 (N_7338,N_6527,N_6497);
or U7339 (N_7339,N_6251,N_6611);
xor U7340 (N_7340,N_6680,N_6406);
nor U7341 (N_7341,N_6285,N_6575);
nor U7342 (N_7342,N_6990,N_6313);
xor U7343 (N_7343,N_6204,N_6860);
nor U7344 (N_7344,N_6787,N_6381);
and U7345 (N_7345,N_6806,N_6873);
or U7346 (N_7346,N_6042,N_6828);
nor U7347 (N_7347,N_6757,N_6515);
nor U7348 (N_7348,N_6552,N_6107);
and U7349 (N_7349,N_6529,N_6464);
and U7350 (N_7350,N_6494,N_6011);
nor U7351 (N_7351,N_6509,N_6465);
nor U7352 (N_7352,N_6049,N_6078);
xor U7353 (N_7353,N_6604,N_6104);
nor U7354 (N_7354,N_6609,N_6560);
nand U7355 (N_7355,N_6682,N_6319);
or U7356 (N_7356,N_6815,N_6864);
or U7357 (N_7357,N_6556,N_6071);
nand U7358 (N_7358,N_6435,N_6794);
and U7359 (N_7359,N_6785,N_6513);
nand U7360 (N_7360,N_6717,N_6647);
and U7361 (N_7361,N_6811,N_6807);
xnor U7362 (N_7362,N_6644,N_6260);
or U7363 (N_7363,N_6252,N_6317);
nand U7364 (N_7364,N_6036,N_6048);
nor U7365 (N_7365,N_6192,N_6450);
nand U7366 (N_7366,N_6158,N_6668);
and U7367 (N_7367,N_6667,N_6488);
xor U7368 (N_7368,N_6946,N_6354);
xor U7369 (N_7369,N_6024,N_6139);
xnor U7370 (N_7370,N_6756,N_6528);
or U7371 (N_7371,N_6487,N_6581);
and U7372 (N_7372,N_6574,N_6169);
xnor U7373 (N_7373,N_6570,N_6728);
nor U7374 (N_7374,N_6395,N_6444);
nor U7375 (N_7375,N_6951,N_6392);
and U7376 (N_7376,N_6148,N_6734);
xnor U7377 (N_7377,N_6861,N_6449);
or U7378 (N_7378,N_6921,N_6230);
or U7379 (N_7379,N_6496,N_6189);
nand U7380 (N_7380,N_6312,N_6126);
xor U7381 (N_7381,N_6718,N_6057);
xor U7382 (N_7382,N_6372,N_6984);
nand U7383 (N_7383,N_6721,N_6518);
and U7384 (N_7384,N_6695,N_6288);
nor U7385 (N_7385,N_6755,N_6479);
nand U7386 (N_7386,N_6292,N_6366);
nor U7387 (N_7387,N_6110,N_6006);
or U7388 (N_7388,N_6180,N_6194);
nand U7389 (N_7389,N_6244,N_6506);
and U7390 (N_7390,N_6731,N_6008);
or U7391 (N_7391,N_6676,N_6084);
xnor U7392 (N_7392,N_6866,N_6135);
or U7393 (N_7393,N_6129,N_6371);
nand U7394 (N_7394,N_6543,N_6708);
xor U7395 (N_7395,N_6168,N_6351);
nand U7396 (N_7396,N_6105,N_6454);
or U7397 (N_7397,N_6287,N_6022);
or U7398 (N_7398,N_6474,N_6277);
xor U7399 (N_7399,N_6501,N_6207);
xor U7400 (N_7400,N_6418,N_6221);
and U7401 (N_7401,N_6791,N_6213);
xor U7402 (N_7402,N_6843,N_6459);
nor U7403 (N_7403,N_6113,N_6485);
nand U7404 (N_7404,N_6216,N_6136);
nand U7405 (N_7405,N_6551,N_6410);
or U7406 (N_7406,N_6631,N_6088);
xnor U7407 (N_7407,N_6714,N_6467);
or U7408 (N_7408,N_6118,N_6924);
nor U7409 (N_7409,N_6428,N_6438);
nand U7410 (N_7410,N_6193,N_6329);
nand U7411 (N_7411,N_6384,N_6373);
or U7412 (N_7412,N_6089,N_6340);
or U7413 (N_7413,N_6805,N_6352);
and U7414 (N_7414,N_6781,N_6548);
and U7415 (N_7415,N_6431,N_6801);
nand U7416 (N_7416,N_6334,N_6561);
xor U7417 (N_7417,N_6208,N_6902);
nor U7418 (N_7418,N_6686,N_6553);
xnor U7419 (N_7419,N_6367,N_6270);
and U7420 (N_7420,N_6665,N_6707);
or U7421 (N_7421,N_6679,N_6605);
nand U7422 (N_7422,N_6685,N_6744);
nor U7423 (N_7423,N_6991,N_6010);
nand U7424 (N_7424,N_6977,N_6657);
or U7425 (N_7425,N_6632,N_6203);
xnor U7426 (N_7426,N_6014,N_6038);
nand U7427 (N_7427,N_6134,N_6353);
and U7428 (N_7428,N_6303,N_6930);
xnor U7429 (N_7429,N_6035,N_6447);
or U7430 (N_7430,N_6859,N_6622);
and U7431 (N_7431,N_6074,N_6701);
xor U7432 (N_7432,N_6830,N_6538);
and U7433 (N_7433,N_6742,N_6280);
xor U7434 (N_7434,N_6703,N_6226);
nor U7435 (N_7435,N_6771,N_6401);
nor U7436 (N_7436,N_6475,N_6953);
or U7437 (N_7437,N_6600,N_6106);
or U7438 (N_7438,N_6729,N_6952);
or U7439 (N_7439,N_6851,N_6601);
and U7440 (N_7440,N_6847,N_6073);
nand U7441 (N_7441,N_6554,N_6999);
nor U7442 (N_7442,N_6763,N_6645);
xnor U7443 (N_7443,N_6716,N_6989);
and U7444 (N_7444,N_6063,N_6855);
nand U7445 (N_7445,N_6445,N_6880);
and U7446 (N_7446,N_6307,N_6214);
nand U7447 (N_7447,N_6546,N_6654);
or U7448 (N_7448,N_6293,N_6514);
xnor U7449 (N_7449,N_6378,N_6747);
nand U7450 (N_7450,N_6114,N_6652);
nand U7451 (N_7451,N_6000,N_6206);
nor U7452 (N_7452,N_6524,N_6242);
or U7453 (N_7453,N_6722,N_6816);
nor U7454 (N_7454,N_6346,N_6565);
xor U7455 (N_7455,N_6903,N_6580);
nor U7456 (N_7456,N_6640,N_6694);
or U7457 (N_7457,N_6400,N_6299);
xnor U7458 (N_7458,N_6147,N_6749);
nor U7459 (N_7459,N_6732,N_6457);
nand U7460 (N_7460,N_6369,N_6909);
and U7461 (N_7461,N_6314,N_6988);
and U7462 (N_7462,N_6326,N_6382);
nand U7463 (N_7463,N_6339,N_6330);
and U7464 (N_7464,N_6948,N_6232);
or U7465 (N_7465,N_6167,N_6052);
xnor U7466 (N_7466,N_6844,N_6567);
nor U7467 (N_7467,N_6927,N_6154);
nand U7468 (N_7468,N_6452,N_6735);
nor U7469 (N_7469,N_6362,N_6486);
nor U7470 (N_7470,N_6026,N_6306);
nand U7471 (N_7471,N_6827,N_6587);
or U7472 (N_7472,N_6013,N_6949);
xor U7473 (N_7473,N_6150,N_6839);
nand U7474 (N_7474,N_6250,N_6958);
nand U7475 (N_7475,N_6436,N_6696);
xnor U7476 (N_7476,N_6956,N_6225);
or U7477 (N_7477,N_6748,N_6034);
nand U7478 (N_7478,N_6936,N_6463);
or U7479 (N_7479,N_6245,N_6389);
nand U7480 (N_7480,N_6235,N_6472);
nand U7481 (N_7481,N_6692,N_6157);
and U7482 (N_7482,N_6237,N_6072);
nand U7483 (N_7483,N_6945,N_6879);
or U7484 (N_7484,N_6004,N_6621);
nand U7485 (N_7485,N_6754,N_6020);
nand U7486 (N_7486,N_6813,N_6101);
nor U7487 (N_7487,N_6140,N_6702);
or U7488 (N_7488,N_6566,N_6220);
xor U7489 (N_7489,N_6489,N_6282);
and U7490 (N_7490,N_6325,N_6413);
nand U7491 (N_7491,N_6737,N_6163);
or U7492 (N_7492,N_6414,N_6451);
nand U7493 (N_7493,N_6081,N_6164);
or U7494 (N_7494,N_6100,N_6178);
xnor U7495 (N_7495,N_6799,N_6997);
nor U7496 (N_7496,N_6616,N_6291);
xnor U7497 (N_7497,N_6907,N_6658);
or U7498 (N_7498,N_6865,N_6041);
or U7499 (N_7499,N_6875,N_6374);
nand U7500 (N_7500,N_6237,N_6844);
and U7501 (N_7501,N_6928,N_6626);
nor U7502 (N_7502,N_6061,N_6738);
or U7503 (N_7503,N_6625,N_6784);
or U7504 (N_7504,N_6319,N_6068);
nand U7505 (N_7505,N_6159,N_6962);
and U7506 (N_7506,N_6760,N_6630);
xnor U7507 (N_7507,N_6116,N_6963);
xor U7508 (N_7508,N_6841,N_6847);
nand U7509 (N_7509,N_6301,N_6476);
or U7510 (N_7510,N_6720,N_6673);
xor U7511 (N_7511,N_6164,N_6060);
nor U7512 (N_7512,N_6658,N_6592);
nor U7513 (N_7513,N_6856,N_6139);
nand U7514 (N_7514,N_6315,N_6745);
nand U7515 (N_7515,N_6576,N_6754);
and U7516 (N_7516,N_6584,N_6749);
xnor U7517 (N_7517,N_6225,N_6348);
and U7518 (N_7518,N_6255,N_6337);
nand U7519 (N_7519,N_6781,N_6537);
xnor U7520 (N_7520,N_6321,N_6503);
and U7521 (N_7521,N_6426,N_6075);
and U7522 (N_7522,N_6279,N_6744);
nand U7523 (N_7523,N_6403,N_6275);
or U7524 (N_7524,N_6536,N_6558);
nor U7525 (N_7525,N_6938,N_6516);
nor U7526 (N_7526,N_6102,N_6924);
nand U7527 (N_7527,N_6804,N_6310);
nand U7528 (N_7528,N_6839,N_6584);
and U7529 (N_7529,N_6616,N_6698);
and U7530 (N_7530,N_6917,N_6671);
nand U7531 (N_7531,N_6896,N_6169);
xnor U7532 (N_7532,N_6969,N_6069);
xnor U7533 (N_7533,N_6103,N_6077);
nand U7534 (N_7534,N_6598,N_6557);
xnor U7535 (N_7535,N_6037,N_6241);
and U7536 (N_7536,N_6119,N_6933);
xnor U7537 (N_7537,N_6905,N_6251);
or U7538 (N_7538,N_6234,N_6491);
nor U7539 (N_7539,N_6189,N_6492);
xor U7540 (N_7540,N_6381,N_6038);
nor U7541 (N_7541,N_6751,N_6366);
nand U7542 (N_7542,N_6151,N_6612);
and U7543 (N_7543,N_6761,N_6530);
xor U7544 (N_7544,N_6676,N_6591);
and U7545 (N_7545,N_6149,N_6638);
nor U7546 (N_7546,N_6723,N_6242);
and U7547 (N_7547,N_6496,N_6438);
nor U7548 (N_7548,N_6998,N_6749);
nor U7549 (N_7549,N_6861,N_6302);
and U7550 (N_7550,N_6746,N_6035);
and U7551 (N_7551,N_6014,N_6001);
xor U7552 (N_7552,N_6420,N_6340);
nand U7553 (N_7553,N_6959,N_6474);
or U7554 (N_7554,N_6675,N_6591);
nor U7555 (N_7555,N_6282,N_6433);
xnor U7556 (N_7556,N_6287,N_6789);
xor U7557 (N_7557,N_6904,N_6466);
nand U7558 (N_7558,N_6834,N_6341);
and U7559 (N_7559,N_6631,N_6429);
and U7560 (N_7560,N_6264,N_6707);
nand U7561 (N_7561,N_6600,N_6205);
and U7562 (N_7562,N_6247,N_6412);
nand U7563 (N_7563,N_6910,N_6546);
nor U7564 (N_7564,N_6636,N_6692);
xor U7565 (N_7565,N_6045,N_6007);
nand U7566 (N_7566,N_6304,N_6427);
xnor U7567 (N_7567,N_6463,N_6759);
nand U7568 (N_7568,N_6641,N_6640);
nand U7569 (N_7569,N_6568,N_6977);
nor U7570 (N_7570,N_6779,N_6617);
nor U7571 (N_7571,N_6131,N_6596);
nor U7572 (N_7572,N_6654,N_6506);
or U7573 (N_7573,N_6049,N_6660);
xnor U7574 (N_7574,N_6039,N_6029);
nand U7575 (N_7575,N_6641,N_6485);
nor U7576 (N_7576,N_6149,N_6496);
nor U7577 (N_7577,N_6240,N_6306);
or U7578 (N_7578,N_6983,N_6707);
nor U7579 (N_7579,N_6642,N_6366);
nand U7580 (N_7580,N_6715,N_6899);
and U7581 (N_7581,N_6044,N_6313);
or U7582 (N_7582,N_6274,N_6924);
or U7583 (N_7583,N_6761,N_6311);
nor U7584 (N_7584,N_6608,N_6836);
and U7585 (N_7585,N_6129,N_6584);
nor U7586 (N_7586,N_6440,N_6582);
and U7587 (N_7587,N_6273,N_6402);
xnor U7588 (N_7588,N_6616,N_6080);
and U7589 (N_7589,N_6297,N_6740);
xnor U7590 (N_7590,N_6022,N_6693);
nand U7591 (N_7591,N_6373,N_6266);
and U7592 (N_7592,N_6905,N_6885);
xnor U7593 (N_7593,N_6565,N_6468);
nand U7594 (N_7594,N_6391,N_6691);
nor U7595 (N_7595,N_6692,N_6644);
nor U7596 (N_7596,N_6518,N_6314);
nand U7597 (N_7597,N_6929,N_6354);
nor U7598 (N_7598,N_6144,N_6344);
or U7599 (N_7599,N_6500,N_6954);
xor U7600 (N_7600,N_6382,N_6064);
and U7601 (N_7601,N_6993,N_6844);
and U7602 (N_7602,N_6823,N_6303);
nor U7603 (N_7603,N_6079,N_6307);
xnor U7604 (N_7604,N_6605,N_6684);
or U7605 (N_7605,N_6653,N_6918);
or U7606 (N_7606,N_6569,N_6266);
nor U7607 (N_7607,N_6149,N_6606);
nand U7608 (N_7608,N_6479,N_6622);
nor U7609 (N_7609,N_6977,N_6444);
xnor U7610 (N_7610,N_6742,N_6253);
xor U7611 (N_7611,N_6809,N_6934);
or U7612 (N_7612,N_6256,N_6706);
nor U7613 (N_7613,N_6118,N_6437);
or U7614 (N_7614,N_6877,N_6297);
nand U7615 (N_7615,N_6504,N_6998);
and U7616 (N_7616,N_6602,N_6044);
nor U7617 (N_7617,N_6572,N_6785);
or U7618 (N_7618,N_6871,N_6058);
xor U7619 (N_7619,N_6557,N_6804);
nand U7620 (N_7620,N_6067,N_6498);
nor U7621 (N_7621,N_6954,N_6801);
and U7622 (N_7622,N_6731,N_6718);
and U7623 (N_7623,N_6506,N_6227);
xnor U7624 (N_7624,N_6576,N_6386);
xnor U7625 (N_7625,N_6708,N_6153);
xnor U7626 (N_7626,N_6199,N_6325);
or U7627 (N_7627,N_6472,N_6428);
nor U7628 (N_7628,N_6910,N_6886);
nand U7629 (N_7629,N_6239,N_6233);
nand U7630 (N_7630,N_6523,N_6508);
nand U7631 (N_7631,N_6878,N_6130);
and U7632 (N_7632,N_6890,N_6146);
nand U7633 (N_7633,N_6530,N_6233);
xnor U7634 (N_7634,N_6493,N_6526);
nand U7635 (N_7635,N_6196,N_6719);
or U7636 (N_7636,N_6695,N_6046);
nor U7637 (N_7637,N_6586,N_6077);
nand U7638 (N_7638,N_6166,N_6634);
and U7639 (N_7639,N_6631,N_6966);
nor U7640 (N_7640,N_6875,N_6937);
and U7641 (N_7641,N_6471,N_6354);
nand U7642 (N_7642,N_6694,N_6122);
and U7643 (N_7643,N_6851,N_6449);
and U7644 (N_7644,N_6491,N_6422);
xor U7645 (N_7645,N_6955,N_6038);
nor U7646 (N_7646,N_6228,N_6515);
and U7647 (N_7647,N_6541,N_6504);
or U7648 (N_7648,N_6348,N_6622);
and U7649 (N_7649,N_6325,N_6002);
nand U7650 (N_7650,N_6397,N_6698);
nand U7651 (N_7651,N_6044,N_6961);
and U7652 (N_7652,N_6711,N_6320);
xnor U7653 (N_7653,N_6604,N_6892);
and U7654 (N_7654,N_6564,N_6043);
xor U7655 (N_7655,N_6015,N_6196);
nand U7656 (N_7656,N_6158,N_6943);
nor U7657 (N_7657,N_6512,N_6199);
or U7658 (N_7658,N_6958,N_6653);
and U7659 (N_7659,N_6849,N_6074);
xor U7660 (N_7660,N_6091,N_6092);
nand U7661 (N_7661,N_6893,N_6800);
nand U7662 (N_7662,N_6245,N_6711);
nand U7663 (N_7663,N_6453,N_6561);
nor U7664 (N_7664,N_6406,N_6986);
nand U7665 (N_7665,N_6162,N_6356);
or U7666 (N_7666,N_6331,N_6471);
xor U7667 (N_7667,N_6911,N_6872);
xnor U7668 (N_7668,N_6406,N_6468);
or U7669 (N_7669,N_6094,N_6397);
xnor U7670 (N_7670,N_6782,N_6798);
xnor U7671 (N_7671,N_6903,N_6105);
or U7672 (N_7672,N_6378,N_6278);
xnor U7673 (N_7673,N_6502,N_6136);
nor U7674 (N_7674,N_6484,N_6266);
or U7675 (N_7675,N_6608,N_6907);
and U7676 (N_7676,N_6236,N_6544);
or U7677 (N_7677,N_6418,N_6409);
nand U7678 (N_7678,N_6036,N_6434);
xnor U7679 (N_7679,N_6078,N_6925);
or U7680 (N_7680,N_6045,N_6547);
and U7681 (N_7681,N_6477,N_6591);
nand U7682 (N_7682,N_6490,N_6335);
nand U7683 (N_7683,N_6992,N_6416);
and U7684 (N_7684,N_6099,N_6621);
xor U7685 (N_7685,N_6344,N_6332);
nand U7686 (N_7686,N_6797,N_6875);
nand U7687 (N_7687,N_6905,N_6825);
and U7688 (N_7688,N_6597,N_6520);
nand U7689 (N_7689,N_6092,N_6968);
or U7690 (N_7690,N_6670,N_6819);
and U7691 (N_7691,N_6200,N_6104);
nor U7692 (N_7692,N_6648,N_6394);
xnor U7693 (N_7693,N_6167,N_6099);
or U7694 (N_7694,N_6498,N_6553);
nor U7695 (N_7695,N_6719,N_6961);
nor U7696 (N_7696,N_6733,N_6119);
nor U7697 (N_7697,N_6779,N_6596);
nand U7698 (N_7698,N_6409,N_6773);
nor U7699 (N_7699,N_6851,N_6334);
nor U7700 (N_7700,N_6022,N_6832);
and U7701 (N_7701,N_6657,N_6402);
nand U7702 (N_7702,N_6170,N_6181);
nand U7703 (N_7703,N_6416,N_6387);
nor U7704 (N_7704,N_6146,N_6260);
or U7705 (N_7705,N_6238,N_6093);
or U7706 (N_7706,N_6946,N_6407);
nor U7707 (N_7707,N_6743,N_6102);
nand U7708 (N_7708,N_6368,N_6975);
nand U7709 (N_7709,N_6636,N_6412);
nor U7710 (N_7710,N_6617,N_6331);
or U7711 (N_7711,N_6394,N_6110);
or U7712 (N_7712,N_6808,N_6009);
nand U7713 (N_7713,N_6616,N_6794);
nand U7714 (N_7714,N_6017,N_6656);
or U7715 (N_7715,N_6183,N_6376);
and U7716 (N_7716,N_6704,N_6528);
xor U7717 (N_7717,N_6517,N_6221);
nand U7718 (N_7718,N_6625,N_6010);
nand U7719 (N_7719,N_6343,N_6049);
xnor U7720 (N_7720,N_6891,N_6978);
or U7721 (N_7721,N_6890,N_6493);
or U7722 (N_7722,N_6360,N_6796);
nor U7723 (N_7723,N_6475,N_6156);
or U7724 (N_7724,N_6044,N_6919);
or U7725 (N_7725,N_6387,N_6801);
xor U7726 (N_7726,N_6393,N_6926);
and U7727 (N_7727,N_6014,N_6699);
and U7728 (N_7728,N_6557,N_6840);
and U7729 (N_7729,N_6778,N_6146);
xnor U7730 (N_7730,N_6551,N_6884);
xnor U7731 (N_7731,N_6391,N_6767);
and U7732 (N_7732,N_6551,N_6924);
nand U7733 (N_7733,N_6776,N_6172);
xnor U7734 (N_7734,N_6998,N_6834);
xnor U7735 (N_7735,N_6766,N_6762);
nor U7736 (N_7736,N_6995,N_6114);
xor U7737 (N_7737,N_6175,N_6753);
nor U7738 (N_7738,N_6747,N_6083);
nand U7739 (N_7739,N_6230,N_6582);
nand U7740 (N_7740,N_6475,N_6137);
nor U7741 (N_7741,N_6884,N_6359);
nor U7742 (N_7742,N_6938,N_6837);
nand U7743 (N_7743,N_6090,N_6362);
and U7744 (N_7744,N_6313,N_6671);
xnor U7745 (N_7745,N_6041,N_6228);
nor U7746 (N_7746,N_6707,N_6253);
or U7747 (N_7747,N_6871,N_6589);
or U7748 (N_7748,N_6568,N_6082);
nor U7749 (N_7749,N_6610,N_6011);
and U7750 (N_7750,N_6816,N_6455);
or U7751 (N_7751,N_6329,N_6298);
and U7752 (N_7752,N_6342,N_6129);
or U7753 (N_7753,N_6863,N_6485);
or U7754 (N_7754,N_6371,N_6362);
nand U7755 (N_7755,N_6808,N_6817);
nor U7756 (N_7756,N_6991,N_6002);
xor U7757 (N_7757,N_6699,N_6305);
xor U7758 (N_7758,N_6056,N_6342);
or U7759 (N_7759,N_6148,N_6139);
xor U7760 (N_7760,N_6694,N_6089);
and U7761 (N_7761,N_6464,N_6305);
nand U7762 (N_7762,N_6071,N_6852);
nor U7763 (N_7763,N_6561,N_6348);
or U7764 (N_7764,N_6781,N_6927);
and U7765 (N_7765,N_6002,N_6093);
and U7766 (N_7766,N_6891,N_6743);
xor U7767 (N_7767,N_6629,N_6557);
xor U7768 (N_7768,N_6309,N_6711);
xor U7769 (N_7769,N_6333,N_6029);
and U7770 (N_7770,N_6454,N_6791);
and U7771 (N_7771,N_6495,N_6004);
and U7772 (N_7772,N_6047,N_6684);
nor U7773 (N_7773,N_6729,N_6311);
or U7774 (N_7774,N_6785,N_6601);
or U7775 (N_7775,N_6282,N_6678);
nand U7776 (N_7776,N_6498,N_6703);
nor U7777 (N_7777,N_6863,N_6237);
or U7778 (N_7778,N_6305,N_6545);
xnor U7779 (N_7779,N_6891,N_6075);
or U7780 (N_7780,N_6093,N_6730);
xnor U7781 (N_7781,N_6373,N_6735);
xnor U7782 (N_7782,N_6284,N_6113);
nand U7783 (N_7783,N_6622,N_6273);
and U7784 (N_7784,N_6354,N_6141);
nand U7785 (N_7785,N_6842,N_6278);
nor U7786 (N_7786,N_6732,N_6615);
xnor U7787 (N_7787,N_6056,N_6974);
or U7788 (N_7788,N_6852,N_6583);
and U7789 (N_7789,N_6850,N_6812);
xnor U7790 (N_7790,N_6372,N_6649);
nand U7791 (N_7791,N_6213,N_6218);
xnor U7792 (N_7792,N_6875,N_6413);
xor U7793 (N_7793,N_6059,N_6742);
xnor U7794 (N_7794,N_6259,N_6207);
or U7795 (N_7795,N_6194,N_6010);
or U7796 (N_7796,N_6192,N_6616);
nand U7797 (N_7797,N_6301,N_6840);
and U7798 (N_7798,N_6773,N_6329);
or U7799 (N_7799,N_6889,N_6605);
xor U7800 (N_7800,N_6585,N_6980);
and U7801 (N_7801,N_6539,N_6447);
nor U7802 (N_7802,N_6214,N_6921);
and U7803 (N_7803,N_6721,N_6661);
and U7804 (N_7804,N_6290,N_6928);
and U7805 (N_7805,N_6922,N_6110);
and U7806 (N_7806,N_6811,N_6212);
or U7807 (N_7807,N_6347,N_6444);
xor U7808 (N_7808,N_6784,N_6811);
and U7809 (N_7809,N_6194,N_6674);
or U7810 (N_7810,N_6916,N_6731);
or U7811 (N_7811,N_6780,N_6691);
nand U7812 (N_7812,N_6046,N_6406);
or U7813 (N_7813,N_6451,N_6405);
and U7814 (N_7814,N_6594,N_6514);
and U7815 (N_7815,N_6716,N_6289);
nand U7816 (N_7816,N_6674,N_6809);
nand U7817 (N_7817,N_6794,N_6966);
or U7818 (N_7818,N_6364,N_6147);
or U7819 (N_7819,N_6256,N_6026);
or U7820 (N_7820,N_6561,N_6530);
and U7821 (N_7821,N_6642,N_6639);
nand U7822 (N_7822,N_6567,N_6202);
nor U7823 (N_7823,N_6880,N_6325);
or U7824 (N_7824,N_6917,N_6235);
nor U7825 (N_7825,N_6264,N_6617);
xor U7826 (N_7826,N_6316,N_6299);
and U7827 (N_7827,N_6631,N_6937);
and U7828 (N_7828,N_6569,N_6994);
or U7829 (N_7829,N_6913,N_6248);
xnor U7830 (N_7830,N_6011,N_6450);
nor U7831 (N_7831,N_6275,N_6532);
or U7832 (N_7832,N_6341,N_6046);
nand U7833 (N_7833,N_6593,N_6719);
nor U7834 (N_7834,N_6370,N_6734);
nand U7835 (N_7835,N_6700,N_6767);
and U7836 (N_7836,N_6827,N_6930);
nor U7837 (N_7837,N_6971,N_6042);
nand U7838 (N_7838,N_6688,N_6995);
xnor U7839 (N_7839,N_6579,N_6989);
xor U7840 (N_7840,N_6761,N_6897);
nor U7841 (N_7841,N_6433,N_6288);
nor U7842 (N_7842,N_6333,N_6630);
and U7843 (N_7843,N_6909,N_6800);
nor U7844 (N_7844,N_6144,N_6123);
nor U7845 (N_7845,N_6190,N_6959);
nand U7846 (N_7846,N_6374,N_6996);
and U7847 (N_7847,N_6464,N_6418);
nor U7848 (N_7848,N_6695,N_6335);
nand U7849 (N_7849,N_6706,N_6660);
xor U7850 (N_7850,N_6009,N_6830);
xnor U7851 (N_7851,N_6380,N_6703);
nor U7852 (N_7852,N_6534,N_6596);
xor U7853 (N_7853,N_6163,N_6945);
or U7854 (N_7854,N_6068,N_6628);
nand U7855 (N_7855,N_6933,N_6878);
xnor U7856 (N_7856,N_6982,N_6478);
and U7857 (N_7857,N_6704,N_6550);
or U7858 (N_7858,N_6627,N_6792);
xnor U7859 (N_7859,N_6068,N_6872);
nand U7860 (N_7860,N_6127,N_6785);
xor U7861 (N_7861,N_6231,N_6092);
xnor U7862 (N_7862,N_6950,N_6949);
or U7863 (N_7863,N_6393,N_6090);
nor U7864 (N_7864,N_6507,N_6553);
xor U7865 (N_7865,N_6353,N_6175);
xnor U7866 (N_7866,N_6444,N_6427);
and U7867 (N_7867,N_6201,N_6910);
xnor U7868 (N_7868,N_6112,N_6278);
and U7869 (N_7869,N_6948,N_6711);
nor U7870 (N_7870,N_6201,N_6880);
nor U7871 (N_7871,N_6291,N_6374);
or U7872 (N_7872,N_6625,N_6551);
nand U7873 (N_7873,N_6723,N_6565);
xor U7874 (N_7874,N_6384,N_6150);
and U7875 (N_7875,N_6073,N_6792);
nor U7876 (N_7876,N_6058,N_6600);
or U7877 (N_7877,N_6289,N_6331);
nand U7878 (N_7878,N_6158,N_6693);
and U7879 (N_7879,N_6714,N_6085);
xor U7880 (N_7880,N_6139,N_6692);
or U7881 (N_7881,N_6746,N_6933);
nand U7882 (N_7882,N_6930,N_6161);
and U7883 (N_7883,N_6873,N_6545);
and U7884 (N_7884,N_6096,N_6543);
and U7885 (N_7885,N_6985,N_6029);
nand U7886 (N_7886,N_6399,N_6310);
nor U7887 (N_7887,N_6280,N_6420);
and U7888 (N_7888,N_6231,N_6509);
or U7889 (N_7889,N_6696,N_6263);
and U7890 (N_7890,N_6471,N_6786);
and U7891 (N_7891,N_6268,N_6090);
nand U7892 (N_7892,N_6548,N_6406);
and U7893 (N_7893,N_6535,N_6311);
xnor U7894 (N_7894,N_6772,N_6871);
nor U7895 (N_7895,N_6080,N_6622);
nor U7896 (N_7896,N_6876,N_6682);
nor U7897 (N_7897,N_6278,N_6663);
xor U7898 (N_7898,N_6110,N_6281);
xor U7899 (N_7899,N_6708,N_6892);
or U7900 (N_7900,N_6586,N_6560);
nand U7901 (N_7901,N_6365,N_6473);
xor U7902 (N_7902,N_6091,N_6446);
and U7903 (N_7903,N_6065,N_6211);
nor U7904 (N_7904,N_6832,N_6672);
or U7905 (N_7905,N_6491,N_6899);
nor U7906 (N_7906,N_6902,N_6402);
or U7907 (N_7907,N_6193,N_6550);
nand U7908 (N_7908,N_6560,N_6101);
or U7909 (N_7909,N_6729,N_6827);
nand U7910 (N_7910,N_6707,N_6741);
nor U7911 (N_7911,N_6447,N_6636);
xnor U7912 (N_7912,N_6429,N_6375);
nor U7913 (N_7913,N_6586,N_6171);
nor U7914 (N_7914,N_6308,N_6266);
and U7915 (N_7915,N_6906,N_6309);
xnor U7916 (N_7916,N_6337,N_6630);
and U7917 (N_7917,N_6794,N_6396);
nand U7918 (N_7918,N_6301,N_6600);
nand U7919 (N_7919,N_6716,N_6787);
and U7920 (N_7920,N_6519,N_6904);
nor U7921 (N_7921,N_6478,N_6717);
nand U7922 (N_7922,N_6569,N_6818);
and U7923 (N_7923,N_6148,N_6513);
and U7924 (N_7924,N_6908,N_6736);
nor U7925 (N_7925,N_6671,N_6942);
nor U7926 (N_7926,N_6827,N_6276);
or U7927 (N_7927,N_6335,N_6421);
or U7928 (N_7928,N_6066,N_6575);
xor U7929 (N_7929,N_6896,N_6053);
and U7930 (N_7930,N_6171,N_6610);
and U7931 (N_7931,N_6550,N_6339);
and U7932 (N_7932,N_6974,N_6989);
xnor U7933 (N_7933,N_6576,N_6516);
or U7934 (N_7934,N_6665,N_6532);
nand U7935 (N_7935,N_6449,N_6915);
nor U7936 (N_7936,N_6113,N_6009);
or U7937 (N_7937,N_6829,N_6317);
and U7938 (N_7938,N_6487,N_6809);
xnor U7939 (N_7939,N_6193,N_6726);
xor U7940 (N_7940,N_6404,N_6058);
xnor U7941 (N_7941,N_6589,N_6244);
or U7942 (N_7942,N_6248,N_6078);
or U7943 (N_7943,N_6954,N_6935);
xor U7944 (N_7944,N_6387,N_6236);
xor U7945 (N_7945,N_6313,N_6142);
and U7946 (N_7946,N_6469,N_6906);
nor U7947 (N_7947,N_6609,N_6521);
nor U7948 (N_7948,N_6214,N_6810);
xor U7949 (N_7949,N_6690,N_6527);
xor U7950 (N_7950,N_6997,N_6467);
nor U7951 (N_7951,N_6411,N_6373);
and U7952 (N_7952,N_6345,N_6496);
or U7953 (N_7953,N_6293,N_6240);
and U7954 (N_7954,N_6540,N_6654);
and U7955 (N_7955,N_6773,N_6383);
nand U7956 (N_7956,N_6376,N_6575);
and U7957 (N_7957,N_6328,N_6782);
xor U7958 (N_7958,N_6138,N_6261);
nand U7959 (N_7959,N_6322,N_6821);
xor U7960 (N_7960,N_6485,N_6355);
xnor U7961 (N_7961,N_6790,N_6820);
xor U7962 (N_7962,N_6027,N_6454);
and U7963 (N_7963,N_6908,N_6434);
xor U7964 (N_7964,N_6840,N_6145);
or U7965 (N_7965,N_6117,N_6266);
nand U7966 (N_7966,N_6378,N_6792);
nor U7967 (N_7967,N_6424,N_6569);
nor U7968 (N_7968,N_6645,N_6597);
and U7969 (N_7969,N_6160,N_6916);
xnor U7970 (N_7970,N_6111,N_6246);
xor U7971 (N_7971,N_6905,N_6399);
xnor U7972 (N_7972,N_6546,N_6653);
and U7973 (N_7973,N_6073,N_6798);
nand U7974 (N_7974,N_6860,N_6593);
or U7975 (N_7975,N_6284,N_6477);
xor U7976 (N_7976,N_6841,N_6007);
nand U7977 (N_7977,N_6906,N_6915);
xor U7978 (N_7978,N_6779,N_6820);
xor U7979 (N_7979,N_6901,N_6516);
nand U7980 (N_7980,N_6969,N_6456);
or U7981 (N_7981,N_6752,N_6025);
nand U7982 (N_7982,N_6879,N_6747);
xnor U7983 (N_7983,N_6052,N_6412);
or U7984 (N_7984,N_6274,N_6262);
xnor U7985 (N_7985,N_6407,N_6759);
nand U7986 (N_7986,N_6485,N_6668);
xor U7987 (N_7987,N_6321,N_6260);
or U7988 (N_7988,N_6734,N_6949);
nand U7989 (N_7989,N_6657,N_6419);
nand U7990 (N_7990,N_6717,N_6879);
and U7991 (N_7991,N_6239,N_6024);
nor U7992 (N_7992,N_6289,N_6696);
or U7993 (N_7993,N_6569,N_6440);
or U7994 (N_7994,N_6449,N_6426);
nor U7995 (N_7995,N_6758,N_6628);
or U7996 (N_7996,N_6785,N_6586);
and U7997 (N_7997,N_6470,N_6220);
and U7998 (N_7998,N_6206,N_6389);
nand U7999 (N_7999,N_6285,N_6685);
nor U8000 (N_8000,N_7750,N_7257);
nor U8001 (N_8001,N_7616,N_7506);
nand U8002 (N_8002,N_7555,N_7442);
xor U8003 (N_8003,N_7038,N_7647);
and U8004 (N_8004,N_7181,N_7448);
nand U8005 (N_8005,N_7211,N_7546);
and U8006 (N_8006,N_7351,N_7797);
xnor U8007 (N_8007,N_7146,N_7652);
nor U8008 (N_8008,N_7645,N_7269);
nor U8009 (N_8009,N_7423,N_7260);
or U8010 (N_8010,N_7853,N_7514);
nand U8011 (N_8011,N_7457,N_7337);
or U8012 (N_8012,N_7524,N_7928);
nand U8013 (N_8013,N_7094,N_7069);
xnor U8014 (N_8014,N_7238,N_7954);
nor U8015 (N_8015,N_7931,N_7678);
nor U8016 (N_8016,N_7341,N_7716);
nor U8017 (N_8017,N_7128,N_7218);
or U8018 (N_8018,N_7193,N_7733);
nor U8019 (N_8019,N_7771,N_7032);
or U8020 (N_8020,N_7608,N_7274);
and U8021 (N_8021,N_7400,N_7369);
xor U8022 (N_8022,N_7386,N_7730);
nor U8023 (N_8023,N_7018,N_7511);
nand U8024 (N_8024,N_7809,N_7941);
or U8025 (N_8025,N_7075,N_7398);
nor U8026 (N_8026,N_7603,N_7317);
xnor U8027 (N_8027,N_7751,N_7049);
and U8028 (N_8028,N_7946,N_7587);
xnor U8029 (N_8029,N_7714,N_7474);
or U8030 (N_8030,N_7254,N_7418);
or U8031 (N_8031,N_7168,N_7549);
nor U8032 (N_8032,N_7694,N_7986);
nor U8033 (N_8033,N_7695,N_7158);
and U8034 (N_8034,N_7329,N_7842);
xnor U8035 (N_8035,N_7190,N_7342);
nor U8036 (N_8036,N_7405,N_7642);
nor U8037 (N_8037,N_7911,N_7082);
nand U8038 (N_8038,N_7489,N_7131);
nand U8039 (N_8039,N_7718,N_7106);
or U8040 (N_8040,N_7175,N_7536);
and U8041 (N_8041,N_7999,N_7530);
or U8042 (N_8042,N_7803,N_7284);
and U8043 (N_8043,N_7787,N_7255);
nor U8044 (N_8044,N_7452,N_7960);
and U8045 (N_8045,N_7854,N_7490);
and U8046 (N_8046,N_7163,N_7118);
xor U8047 (N_8047,N_7836,N_7942);
nor U8048 (N_8048,N_7039,N_7611);
or U8049 (N_8049,N_7592,N_7785);
or U8050 (N_8050,N_7811,N_7015);
and U8051 (N_8051,N_7129,N_7174);
nand U8052 (N_8052,N_7844,N_7164);
xnor U8053 (N_8053,N_7302,N_7731);
nand U8054 (N_8054,N_7690,N_7055);
or U8055 (N_8055,N_7562,N_7689);
and U8056 (N_8056,N_7330,N_7240);
nand U8057 (N_8057,N_7320,N_7065);
or U8058 (N_8058,N_7793,N_7145);
or U8059 (N_8059,N_7265,N_7207);
or U8060 (N_8060,N_7304,N_7824);
or U8061 (N_8061,N_7570,N_7821);
and U8062 (N_8062,N_7961,N_7684);
nand U8063 (N_8063,N_7060,N_7826);
xor U8064 (N_8064,N_7007,N_7185);
and U8065 (N_8065,N_7888,N_7495);
and U8066 (N_8066,N_7743,N_7875);
nor U8067 (N_8067,N_7250,N_7231);
nor U8068 (N_8068,N_7076,N_7768);
nand U8069 (N_8069,N_7140,N_7825);
nand U8070 (N_8070,N_7117,N_7576);
and U8071 (N_8071,N_7995,N_7027);
nor U8072 (N_8072,N_7899,N_7370);
and U8073 (N_8073,N_7701,N_7124);
or U8074 (N_8074,N_7479,N_7962);
and U8075 (N_8075,N_7557,N_7155);
nand U8076 (N_8076,N_7385,N_7650);
xnor U8077 (N_8077,N_7191,N_7580);
and U8078 (N_8078,N_7368,N_7982);
nand U8079 (N_8079,N_7979,N_7219);
nand U8080 (N_8080,N_7827,N_7139);
xnor U8081 (N_8081,N_7950,N_7513);
nand U8082 (N_8082,N_7331,N_7992);
nor U8083 (N_8083,N_7275,N_7727);
xnor U8084 (N_8084,N_7379,N_7522);
nand U8085 (N_8085,N_7217,N_7291);
nor U8086 (N_8086,N_7981,N_7382);
xnor U8087 (N_8087,N_7905,N_7829);
nor U8088 (N_8088,N_7259,N_7841);
nor U8089 (N_8089,N_7098,N_7700);
xnor U8090 (N_8090,N_7212,N_7309);
or U8091 (N_8091,N_7907,N_7074);
xor U8092 (N_8092,N_7741,N_7553);
nand U8093 (N_8093,N_7802,N_7560);
and U8094 (N_8094,N_7444,N_7441);
xor U8095 (N_8095,N_7092,N_7728);
nand U8096 (N_8096,N_7850,N_7769);
nor U8097 (N_8097,N_7569,N_7437);
and U8098 (N_8098,N_7738,N_7571);
nor U8099 (N_8099,N_7066,N_7481);
nor U8100 (N_8100,N_7160,N_7749);
xnor U8101 (N_8101,N_7097,N_7040);
nor U8102 (N_8102,N_7804,N_7293);
or U8103 (N_8103,N_7088,N_7206);
nor U8104 (N_8104,N_7488,N_7313);
nand U8105 (N_8105,N_7149,N_7294);
and U8106 (N_8106,N_7162,N_7770);
nand U8107 (N_8107,N_7396,N_7390);
nand U8108 (N_8108,N_7817,N_7619);
and U8109 (N_8109,N_7394,N_7093);
nor U8110 (N_8110,N_7624,N_7438);
and U8111 (N_8111,N_7552,N_7846);
nor U8112 (N_8112,N_7063,N_7432);
xnor U8113 (N_8113,N_7648,N_7053);
xnor U8114 (N_8114,N_7409,N_7073);
xor U8115 (N_8115,N_7614,N_7711);
and U8116 (N_8116,N_7148,N_7556);
and U8117 (N_8117,N_7970,N_7510);
or U8118 (N_8118,N_7737,N_7115);
nor U8119 (N_8119,N_7504,N_7980);
nand U8120 (N_8120,N_7143,N_7508);
xnor U8121 (N_8121,N_7675,N_7515);
xnor U8122 (N_8122,N_7589,N_7189);
and U8123 (N_8123,N_7558,N_7984);
or U8124 (N_8124,N_7110,N_7713);
xnor U8125 (N_8125,N_7554,N_7201);
xor U8126 (N_8126,N_7141,N_7917);
nand U8127 (N_8127,N_7563,N_7296);
nand U8128 (N_8128,N_7280,N_7107);
and U8129 (N_8129,N_7402,N_7381);
or U8130 (N_8130,N_7828,N_7346);
nor U8131 (N_8131,N_7584,N_7748);
and U8132 (N_8132,N_7134,N_7273);
xnor U8133 (N_8133,N_7879,N_7739);
xnor U8134 (N_8134,N_7318,N_7985);
or U8135 (N_8135,N_7401,N_7864);
and U8136 (N_8136,N_7550,N_7976);
and U8137 (N_8137,N_7865,N_7615);
nand U8138 (N_8138,N_7677,N_7334);
or U8139 (N_8139,N_7876,N_7968);
nand U8140 (N_8140,N_7416,N_7077);
nor U8141 (N_8141,N_7732,N_7095);
xor U8142 (N_8142,N_7578,N_7159);
nor U8143 (N_8143,N_7637,N_7367);
xnor U8144 (N_8144,N_7268,N_7167);
or U8145 (N_8145,N_7012,N_7539);
nor U8146 (N_8146,N_7877,N_7216);
nand U8147 (N_8147,N_7453,N_7639);
xnor U8148 (N_8148,N_7500,N_7165);
and U8149 (N_8149,N_7655,N_7610);
nand U8150 (N_8150,N_7724,N_7236);
nand U8151 (N_8151,N_7150,N_7109);
nor U8152 (N_8152,N_7031,N_7043);
or U8153 (N_8153,N_7246,N_7096);
or U8154 (N_8154,N_7990,N_7964);
and U8155 (N_8155,N_7901,N_7264);
and U8156 (N_8156,N_7994,N_7204);
nor U8157 (N_8157,N_7213,N_7757);
or U8158 (N_8158,N_7256,N_7154);
nor U8159 (N_8159,N_7956,N_7064);
or U8160 (N_8160,N_7358,N_7832);
or U8161 (N_8161,N_7224,N_7443);
or U8162 (N_8162,N_7988,N_7362);
or U8163 (N_8163,N_7262,N_7178);
xnor U8164 (N_8164,N_7407,N_7940);
xnor U8165 (N_8165,N_7326,N_7860);
or U8166 (N_8166,N_7532,N_7779);
nand U8167 (N_8167,N_7023,N_7475);
nor U8168 (N_8168,N_7035,N_7322);
xnor U8169 (N_8169,N_7818,N_7881);
xor U8170 (N_8170,N_7679,N_7458);
nand U8171 (N_8171,N_7121,N_7799);
nand U8172 (N_8172,N_7024,N_7340);
nand U8173 (N_8173,N_7004,N_7062);
or U8174 (N_8174,N_7450,N_7108);
nor U8175 (N_8175,N_7674,N_7939);
nand U8176 (N_8176,N_7840,N_7235);
nand U8177 (N_8177,N_7632,N_7891);
or U8178 (N_8178,N_7210,N_7788);
nor U8179 (N_8179,N_7903,N_7391);
nor U8180 (N_8180,N_7355,N_7525);
and U8181 (N_8181,N_7133,N_7651);
nand U8182 (N_8182,N_7130,N_7449);
nand U8183 (N_8183,N_7923,N_7858);
or U8184 (N_8184,N_7173,N_7104);
nor U8185 (N_8185,N_7503,N_7314);
nand U8186 (N_8186,N_7087,N_7435);
nand U8187 (N_8187,N_7482,N_7215);
or U8188 (N_8188,N_7719,N_7880);
nand U8189 (N_8189,N_7413,N_7883);
nand U8190 (N_8190,N_7561,N_7627);
xor U8191 (N_8191,N_7581,N_7372);
nor U8192 (N_8192,N_7758,N_7237);
and U8193 (N_8193,N_7792,N_7323);
nor U8194 (N_8194,N_7930,N_7755);
or U8195 (N_8195,N_7760,N_7568);
and U8196 (N_8196,N_7430,N_7297);
and U8197 (N_8197,N_7278,N_7308);
xor U8198 (N_8198,N_7166,N_7312);
or U8199 (N_8199,N_7955,N_7464);
nor U8200 (N_8200,N_7815,N_7017);
and U8201 (N_8201,N_7798,N_7182);
or U8202 (N_8202,N_7873,N_7483);
nor U8203 (N_8203,N_7411,N_7629);
or U8204 (N_8204,N_7292,N_7279);
or U8205 (N_8205,N_7099,N_7664);
and U8206 (N_8206,N_7068,N_7991);
xnor U8207 (N_8207,N_7285,N_7969);
nand U8208 (N_8208,N_7567,N_7574);
and U8209 (N_8209,N_7239,N_7606);
nor U8210 (N_8210,N_7671,N_7915);
and U8211 (N_8211,N_7157,N_7541);
nand U8212 (N_8212,N_7693,N_7277);
nor U8213 (N_8213,N_7203,N_7445);
nand U8214 (N_8214,N_7467,N_7335);
xnor U8215 (N_8215,N_7670,N_7625);
xnor U8216 (N_8216,N_7517,N_7975);
or U8217 (N_8217,N_7963,N_7559);
xnor U8218 (N_8218,N_7820,N_7360);
nor U8219 (N_8219,N_7747,N_7564);
xnor U8220 (N_8220,N_7319,N_7226);
nand U8221 (N_8221,N_7593,N_7338);
nor U8222 (N_8222,N_7813,N_7753);
nor U8223 (N_8223,N_7949,N_7583);
xnor U8224 (N_8224,N_7666,N_7710);
xor U8225 (N_8225,N_7657,N_7433);
xor U8226 (N_8226,N_7344,N_7894);
nand U8227 (N_8227,N_7228,N_7403);
nand U8228 (N_8228,N_7626,N_7686);
or U8229 (N_8229,N_7659,N_7126);
nand U8230 (N_8230,N_7003,N_7512);
xor U8231 (N_8231,N_7878,N_7653);
and U8232 (N_8232,N_7925,N_7588);
and U8233 (N_8233,N_7208,N_7046);
nor U8234 (N_8234,N_7597,N_7912);
nor U8235 (N_8235,N_7451,N_7465);
xor U8236 (N_8236,N_7786,N_7889);
xnor U8237 (N_8237,N_7740,N_7113);
nor U8238 (N_8238,N_7663,N_7658);
nand U8239 (N_8239,N_7998,N_7183);
nand U8240 (N_8240,N_7026,N_7882);
and U8241 (N_8241,N_7350,N_7058);
and U8242 (N_8242,N_7456,N_7951);
and U8243 (N_8243,N_7699,N_7544);
and U8244 (N_8244,N_7623,N_7682);
xor U8245 (N_8245,N_7518,N_7742);
and U8246 (N_8246,N_7520,N_7725);
or U8247 (N_8247,N_7874,N_7127);
or U8248 (N_8248,N_7989,N_7596);
or U8249 (N_8249,N_7598,N_7373);
or U8250 (N_8250,N_7047,N_7287);
nor U8251 (N_8251,N_7766,N_7784);
nand U8252 (N_8252,N_7180,N_7849);
xor U8253 (N_8253,N_7387,N_7052);
and U8254 (N_8254,N_7202,N_7871);
nor U8255 (N_8255,N_7920,N_7276);
and U8256 (N_8256,N_7646,N_7656);
nor U8257 (N_8257,N_7487,N_7613);
nand U8258 (N_8258,N_7491,N_7927);
nor U8259 (N_8259,N_7848,N_7136);
or U8260 (N_8260,N_7147,N_7466);
nand U8261 (N_8261,N_7997,N_7958);
nand U8262 (N_8262,N_7186,N_7179);
and U8263 (N_8263,N_7683,N_7311);
nor U8264 (N_8264,N_7702,N_7575);
xnor U8265 (N_8265,N_7234,N_7298);
or U8266 (N_8266,N_7953,N_7199);
and U8267 (N_8267,N_7486,N_7295);
or U8268 (N_8268,N_7404,N_7347);
and U8269 (N_8269,N_7762,N_7187);
nor U8270 (N_8270,N_7359,N_7460);
or U8271 (N_8271,N_7484,N_7688);
or U8272 (N_8272,N_7054,N_7408);
or U8273 (N_8273,N_7778,N_7170);
and U8274 (N_8274,N_7957,N_7116);
or U8275 (N_8275,N_7735,N_7498);
nand U8276 (N_8276,N_7943,N_7783);
or U8277 (N_8277,N_7644,N_7703);
xnor U8278 (N_8278,N_7230,N_7083);
nor U8279 (N_8279,N_7222,N_7469);
or U8280 (N_8280,N_7566,N_7947);
xnor U8281 (N_8281,N_7497,N_7843);
nand U8282 (N_8282,N_7636,N_7764);
xor U8283 (N_8283,N_7041,N_7025);
nor U8284 (N_8284,N_7904,N_7196);
nor U8285 (N_8285,N_7021,N_7022);
nor U8286 (N_8286,N_7414,N_7717);
nand U8287 (N_8287,N_7343,N_7691);
nand U8288 (N_8288,N_7253,N_7286);
or U8289 (N_8289,N_7014,N_7934);
and U8290 (N_8290,N_7005,N_7908);
and U8291 (N_8291,N_7290,N_7833);
or U8292 (N_8292,N_7258,N_7084);
nand U8293 (N_8293,N_7805,N_7902);
or U8294 (N_8294,N_7247,N_7667);
and U8295 (N_8295,N_7744,N_7363);
and U8296 (N_8296,N_7153,N_7807);
nor U8297 (N_8297,N_7507,N_7527);
and U8298 (N_8298,N_7072,N_7922);
and U8299 (N_8299,N_7897,N_7161);
and U8300 (N_8300,N_7938,N_7845);
or U8301 (N_8301,N_7348,N_7135);
or U8302 (N_8302,N_7471,N_7333);
and U8303 (N_8303,N_7967,N_7537);
and U8304 (N_8304,N_7673,N_7123);
or U8305 (N_8305,N_7654,N_7241);
nand U8306 (N_8306,N_7209,N_7051);
xnor U8307 (N_8307,N_7971,N_7493);
nand U8308 (N_8308,N_7707,N_7214);
nor U8309 (N_8309,N_7582,N_7519);
or U8310 (N_8310,N_7529,N_7754);
and U8311 (N_8311,N_7371,N_7364);
xnor U8312 (N_8312,N_7502,N_7983);
xor U8313 (N_8313,N_7472,N_7188);
nand U8314 (N_8314,N_7775,N_7959);
and U8315 (N_8315,N_7781,N_7079);
and U8316 (N_8316,N_7426,N_7057);
nand U8317 (N_8317,N_7125,N_7013);
nor U8318 (N_8318,N_7044,N_7756);
nand U8319 (N_8319,N_7872,N_7061);
and U8320 (N_8320,N_7800,N_7447);
or U8321 (N_8321,N_7281,N_7223);
xor U8322 (N_8322,N_7195,N_7263);
or U8323 (N_8323,N_7708,N_7352);
nand U8324 (N_8324,N_7892,N_7114);
nor U8325 (N_8325,N_7509,N_7933);
and U8326 (N_8326,N_7085,N_7814);
xnor U8327 (N_8327,N_7631,N_7974);
nor U8328 (N_8328,N_7336,N_7847);
and U8329 (N_8329,N_7726,N_7151);
nand U8330 (N_8330,N_7070,N_7916);
xnor U8331 (N_8331,N_7935,N_7325);
xor U8332 (N_8332,N_7577,N_7937);
nand U8333 (N_8333,N_7729,N_7704);
nor U8334 (N_8334,N_7019,N_7119);
or U8335 (N_8335,N_7425,N_7384);
nor U8336 (N_8336,N_7028,N_7410);
or U8337 (N_8337,N_7723,N_7374);
nor U8338 (N_8338,N_7638,N_7676);
nor U8339 (N_8339,N_7122,N_7299);
and U8340 (N_8340,N_7176,N_7830);
nand U8341 (N_8341,N_7565,N_7378);
xnor U8342 (N_8342,N_7806,N_7965);
nand U8343 (N_8343,N_7339,N_7000);
and U8344 (N_8344,N_7777,N_7412);
nor U8345 (N_8345,N_7890,N_7857);
xnor U8346 (N_8346,N_7305,N_7137);
or U8347 (N_8347,N_7669,N_7324);
and U8348 (N_8348,N_7542,N_7528);
or U8349 (N_8349,N_7680,N_7586);
xnor U8350 (N_8350,N_7245,N_7681);
and U8351 (N_8351,N_7184,N_7869);
nand U8352 (N_8352,N_7697,N_7609);
and U8353 (N_8353,N_7138,N_7823);
and U8354 (N_8354,N_7790,N_7885);
nor U8355 (N_8355,N_7945,N_7480);
nor U8356 (N_8356,N_7037,N_7105);
or U8357 (N_8357,N_7835,N_7103);
xnor U8358 (N_8358,N_7421,N_7884);
and U8359 (N_8359,N_7436,N_7100);
nand U8360 (N_8360,N_7029,N_7251);
xor U8361 (N_8361,N_7628,N_7776);
nand U8362 (N_8362,N_7831,N_7789);
nand U8363 (N_8363,N_7643,N_7243);
and U8364 (N_8364,N_7056,N_7288);
nor U8365 (N_8365,N_7289,N_7476);
and U8366 (N_8366,N_7492,N_7392);
and U8367 (N_8367,N_7895,N_7399);
and U8368 (N_8368,N_7198,N_7604);
nor U8369 (N_8369,N_7081,N_7966);
or U8370 (N_8370,N_7548,N_7855);
or U8371 (N_8371,N_7194,N_7270);
and U8372 (N_8372,N_7551,N_7376);
nand U8373 (N_8373,N_7242,N_7887);
nor U8374 (N_8374,N_7948,N_7759);
and U8375 (N_8375,N_7709,N_7516);
nor U8376 (N_8376,N_7361,N_7746);
and U8377 (N_8377,N_7761,N_7910);
and U8378 (N_8378,N_7266,N_7635);
xor U8379 (N_8379,N_7712,N_7540);
nor U8380 (N_8380,N_7071,N_7812);
nand U8381 (N_8381,N_7220,N_7594);
nor U8382 (N_8382,N_7819,N_7306);
nor U8383 (N_8383,N_7354,N_7200);
xnor U8384 (N_8384,N_7283,N_7692);
or U8385 (N_8385,N_7868,N_7389);
or U8386 (N_8386,N_7687,N_7091);
and U8387 (N_8387,N_7132,N_7048);
xor U8388 (N_8388,N_7303,N_7356);
or U8389 (N_8389,N_7112,N_7822);
nor U8390 (N_8390,N_7630,N_7375);
nor U8391 (N_8391,N_7834,N_7328);
nor U8392 (N_8392,N_7042,N_7993);
nor U8393 (N_8393,N_7459,N_7377);
and U8394 (N_8394,N_7271,N_7810);
xnor U8395 (N_8395,N_7605,N_7649);
and U8396 (N_8396,N_7366,N_7030);
nand U8397 (N_8397,N_7696,N_7660);
or U8398 (N_8398,N_7485,N_7856);
nand U8399 (N_8399,N_7547,N_7745);
or U8400 (N_8400,N_7365,N_7601);
xnor U8401 (N_8401,N_7316,N_7417);
xor U8402 (N_8402,N_7415,N_7918);
nor U8403 (N_8403,N_7705,N_7461);
nand U8404 (N_8404,N_7397,N_7668);
xnor U8405 (N_8405,N_7380,N_7078);
nor U8406 (N_8406,N_7919,N_7244);
and U8407 (N_8407,N_7016,N_7431);
nor U8408 (N_8408,N_7229,N_7617);
xor U8409 (N_8409,N_7538,N_7393);
and U8410 (N_8410,N_7607,N_7543);
nor U8411 (N_8411,N_7462,N_7221);
nand U8412 (N_8412,N_7863,N_7932);
xnor U8413 (N_8413,N_7591,N_7838);
and U8414 (N_8414,N_7439,N_7177);
nand U8415 (N_8415,N_7996,N_7172);
or U8416 (N_8416,N_7102,N_7535);
nand U8417 (N_8417,N_7205,N_7252);
nand U8418 (N_8418,N_7101,N_7752);
nand U8419 (N_8419,N_7672,N_7620);
xor U8420 (N_8420,N_7767,N_7531);
nand U8421 (N_8421,N_7698,N_7736);
xor U8422 (N_8422,N_7795,N_7913);
xnor U8423 (N_8423,N_7248,N_7307);
xor U8424 (N_8424,N_7640,N_7440);
and U8425 (N_8425,N_7893,N_7772);
xnor U8426 (N_8426,N_7156,N_7020);
and U8427 (N_8427,N_7357,N_7470);
xor U8428 (N_8428,N_7816,N_7010);
or U8429 (N_8429,N_7595,N_7142);
or U8430 (N_8430,N_7232,N_7225);
nor U8431 (N_8431,N_7169,N_7978);
or U8432 (N_8432,N_7249,N_7120);
nand U8433 (N_8433,N_7050,N_7590);
or U8434 (N_8434,N_7089,N_7427);
or U8435 (N_8435,N_7977,N_7987);
or U8436 (N_8436,N_7936,N_7267);
xor U8437 (N_8437,N_7523,N_7633);
and U8438 (N_8438,N_7715,N_7765);
and U8439 (N_8439,N_7473,N_7090);
or U8440 (N_8440,N_7321,N_7002);
and U8441 (N_8441,N_7463,N_7327);
nand U8442 (N_8442,N_7197,N_7429);
nor U8443 (N_8443,N_7454,N_7921);
and U8444 (N_8444,N_7661,N_7599);
nand U8445 (N_8445,N_7272,N_7045);
nand U8446 (N_8446,N_7009,N_7349);
nand U8447 (N_8447,N_7900,N_7796);
xnor U8448 (N_8448,N_7862,N_7300);
nand U8449 (N_8449,N_7634,N_7434);
or U8450 (N_8450,N_7791,N_7420);
and U8451 (N_8451,N_7034,N_7067);
xnor U8452 (N_8452,N_7944,N_7315);
nand U8453 (N_8453,N_7001,N_7395);
xnor U8454 (N_8454,N_7706,N_7774);
xnor U8455 (N_8455,N_7388,N_7924);
and U8456 (N_8456,N_7233,N_7780);
or U8457 (N_8457,N_7861,N_7641);
nor U8458 (N_8458,N_7721,N_7496);
or U8459 (N_8459,N_7621,N_7618);
nand U8460 (N_8460,N_7144,N_7353);
nor U8461 (N_8461,N_7906,N_7870);
nand U8462 (N_8462,N_7383,N_7036);
nor U8463 (N_8463,N_7763,N_7533);
or U8464 (N_8464,N_7782,N_7494);
xor U8465 (N_8465,N_7428,N_7499);
xnor U8466 (N_8466,N_7866,N_7801);
or U8467 (N_8467,N_7406,N_7111);
or U8468 (N_8468,N_7973,N_7622);
xor U8469 (N_8469,N_7886,N_7579);
nor U8470 (N_8470,N_7837,N_7505);
and U8471 (N_8471,N_7851,N_7468);
or U8472 (N_8472,N_7612,N_7534);
nand U8473 (N_8473,N_7720,N_7080);
and U8474 (N_8474,N_7794,N_7867);
nor U8475 (N_8475,N_7477,N_7585);
or U8476 (N_8476,N_7929,N_7808);
nand U8477 (N_8477,N_7859,N_7310);
and U8478 (N_8478,N_7192,N_7773);
and U8479 (N_8479,N_7526,N_7059);
or U8480 (N_8480,N_7722,N_7227);
or U8481 (N_8481,N_7545,N_7914);
nor U8482 (N_8482,N_7839,N_7332);
and U8483 (N_8483,N_7455,N_7419);
nand U8484 (N_8484,N_7662,N_7152);
nor U8485 (N_8485,N_7952,N_7926);
or U8486 (N_8486,N_7008,N_7602);
or U8487 (N_8487,N_7261,N_7572);
nand U8488 (N_8488,N_7345,N_7898);
and U8489 (N_8489,N_7033,N_7896);
nand U8490 (N_8490,N_7909,N_7422);
or U8491 (N_8491,N_7685,N_7501);
nand U8492 (N_8492,N_7282,N_7301);
nand U8493 (N_8493,N_7478,N_7600);
nor U8494 (N_8494,N_7972,N_7446);
and U8495 (N_8495,N_7852,N_7734);
xor U8496 (N_8496,N_7011,N_7171);
xor U8497 (N_8497,N_7665,N_7424);
or U8498 (N_8498,N_7573,N_7006);
or U8499 (N_8499,N_7521,N_7086);
and U8500 (N_8500,N_7931,N_7288);
nor U8501 (N_8501,N_7536,N_7741);
and U8502 (N_8502,N_7806,N_7611);
xnor U8503 (N_8503,N_7729,N_7914);
nor U8504 (N_8504,N_7434,N_7403);
or U8505 (N_8505,N_7980,N_7272);
nand U8506 (N_8506,N_7584,N_7800);
xor U8507 (N_8507,N_7628,N_7075);
and U8508 (N_8508,N_7744,N_7100);
xnor U8509 (N_8509,N_7610,N_7418);
and U8510 (N_8510,N_7385,N_7902);
xnor U8511 (N_8511,N_7474,N_7285);
nand U8512 (N_8512,N_7646,N_7008);
and U8513 (N_8513,N_7683,N_7764);
nor U8514 (N_8514,N_7729,N_7214);
xor U8515 (N_8515,N_7865,N_7464);
nor U8516 (N_8516,N_7588,N_7709);
nor U8517 (N_8517,N_7422,N_7758);
nor U8518 (N_8518,N_7939,N_7435);
nor U8519 (N_8519,N_7191,N_7173);
xnor U8520 (N_8520,N_7814,N_7854);
nor U8521 (N_8521,N_7209,N_7156);
or U8522 (N_8522,N_7904,N_7526);
xor U8523 (N_8523,N_7203,N_7198);
xnor U8524 (N_8524,N_7859,N_7671);
nand U8525 (N_8525,N_7789,N_7314);
or U8526 (N_8526,N_7925,N_7618);
nand U8527 (N_8527,N_7654,N_7053);
xor U8528 (N_8528,N_7886,N_7939);
nand U8529 (N_8529,N_7704,N_7420);
or U8530 (N_8530,N_7554,N_7978);
and U8531 (N_8531,N_7707,N_7588);
xor U8532 (N_8532,N_7997,N_7517);
nand U8533 (N_8533,N_7843,N_7617);
nand U8534 (N_8534,N_7844,N_7155);
xnor U8535 (N_8535,N_7437,N_7174);
nand U8536 (N_8536,N_7077,N_7511);
or U8537 (N_8537,N_7594,N_7847);
nand U8538 (N_8538,N_7580,N_7796);
nor U8539 (N_8539,N_7717,N_7284);
nor U8540 (N_8540,N_7130,N_7064);
or U8541 (N_8541,N_7088,N_7356);
xor U8542 (N_8542,N_7795,N_7377);
xnor U8543 (N_8543,N_7303,N_7153);
nand U8544 (N_8544,N_7323,N_7098);
and U8545 (N_8545,N_7492,N_7240);
nand U8546 (N_8546,N_7756,N_7553);
nor U8547 (N_8547,N_7956,N_7947);
nor U8548 (N_8548,N_7598,N_7694);
and U8549 (N_8549,N_7360,N_7569);
and U8550 (N_8550,N_7453,N_7875);
xnor U8551 (N_8551,N_7992,N_7201);
nor U8552 (N_8552,N_7458,N_7330);
xnor U8553 (N_8553,N_7194,N_7201);
nor U8554 (N_8554,N_7202,N_7106);
nor U8555 (N_8555,N_7087,N_7976);
and U8556 (N_8556,N_7078,N_7898);
or U8557 (N_8557,N_7534,N_7925);
or U8558 (N_8558,N_7591,N_7874);
or U8559 (N_8559,N_7110,N_7116);
nand U8560 (N_8560,N_7929,N_7966);
xor U8561 (N_8561,N_7431,N_7130);
or U8562 (N_8562,N_7525,N_7308);
xor U8563 (N_8563,N_7696,N_7570);
and U8564 (N_8564,N_7618,N_7571);
and U8565 (N_8565,N_7856,N_7892);
xnor U8566 (N_8566,N_7094,N_7832);
xnor U8567 (N_8567,N_7769,N_7257);
xnor U8568 (N_8568,N_7611,N_7379);
and U8569 (N_8569,N_7569,N_7045);
nor U8570 (N_8570,N_7371,N_7800);
nor U8571 (N_8571,N_7801,N_7396);
xor U8572 (N_8572,N_7634,N_7717);
and U8573 (N_8573,N_7826,N_7086);
and U8574 (N_8574,N_7791,N_7778);
nor U8575 (N_8575,N_7428,N_7641);
and U8576 (N_8576,N_7915,N_7152);
and U8577 (N_8577,N_7268,N_7161);
xor U8578 (N_8578,N_7506,N_7672);
nor U8579 (N_8579,N_7950,N_7362);
xnor U8580 (N_8580,N_7963,N_7378);
or U8581 (N_8581,N_7515,N_7283);
or U8582 (N_8582,N_7845,N_7170);
or U8583 (N_8583,N_7997,N_7554);
and U8584 (N_8584,N_7887,N_7684);
nand U8585 (N_8585,N_7677,N_7658);
nor U8586 (N_8586,N_7615,N_7958);
or U8587 (N_8587,N_7801,N_7779);
xor U8588 (N_8588,N_7110,N_7120);
and U8589 (N_8589,N_7679,N_7991);
nand U8590 (N_8590,N_7349,N_7113);
and U8591 (N_8591,N_7991,N_7548);
or U8592 (N_8592,N_7128,N_7040);
nor U8593 (N_8593,N_7262,N_7575);
and U8594 (N_8594,N_7247,N_7413);
xor U8595 (N_8595,N_7578,N_7277);
or U8596 (N_8596,N_7173,N_7163);
nor U8597 (N_8597,N_7962,N_7113);
nand U8598 (N_8598,N_7641,N_7199);
nor U8599 (N_8599,N_7288,N_7249);
or U8600 (N_8600,N_7129,N_7224);
and U8601 (N_8601,N_7455,N_7104);
or U8602 (N_8602,N_7890,N_7242);
or U8603 (N_8603,N_7790,N_7767);
and U8604 (N_8604,N_7408,N_7211);
nor U8605 (N_8605,N_7866,N_7555);
nor U8606 (N_8606,N_7301,N_7690);
or U8607 (N_8607,N_7619,N_7652);
nand U8608 (N_8608,N_7782,N_7556);
or U8609 (N_8609,N_7594,N_7741);
nand U8610 (N_8610,N_7526,N_7154);
nor U8611 (N_8611,N_7876,N_7086);
xor U8612 (N_8612,N_7736,N_7016);
nor U8613 (N_8613,N_7598,N_7350);
nor U8614 (N_8614,N_7942,N_7520);
nor U8615 (N_8615,N_7047,N_7332);
and U8616 (N_8616,N_7980,N_7302);
or U8617 (N_8617,N_7275,N_7247);
nand U8618 (N_8618,N_7096,N_7918);
or U8619 (N_8619,N_7801,N_7736);
nor U8620 (N_8620,N_7638,N_7016);
nor U8621 (N_8621,N_7007,N_7520);
nor U8622 (N_8622,N_7704,N_7467);
and U8623 (N_8623,N_7579,N_7671);
and U8624 (N_8624,N_7311,N_7851);
and U8625 (N_8625,N_7527,N_7586);
nand U8626 (N_8626,N_7634,N_7889);
and U8627 (N_8627,N_7159,N_7464);
and U8628 (N_8628,N_7606,N_7175);
and U8629 (N_8629,N_7561,N_7005);
and U8630 (N_8630,N_7649,N_7337);
nand U8631 (N_8631,N_7427,N_7014);
or U8632 (N_8632,N_7632,N_7526);
or U8633 (N_8633,N_7631,N_7786);
nand U8634 (N_8634,N_7736,N_7722);
nand U8635 (N_8635,N_7235,N_7971);
xnor U8636 (N_8636,N_7398,N_7423);
xor U8637 (N_8637,N_7720,N_7645);
and U8638 (N_8638,N_7927,N_7047);
xor U8639 (N_8639,N_7176,N_7935);
and U8640 (N_8640,N_7106,N_7804);
xnor U8641 (N_8641,N_7229,N_7714);
and U8642 (N_8642,N_7219,N_7180);
or U8643 (N_8643,N_7375,N_7845);
nor U8644 (N_8644,N_7601,N_7280);
and U8645 (N_8645,N_7630,N_7855);
nor U8646 (N_8646,N_7492,N_7286);
nand U8647 (N_8647,N_7047,N_7401);
and U8648 (N_8648,N_7350,N_7803);
xor U8649 (N_8649,N_7372,N_7556);
nand U8650 (N_8650,N_7057,N_7544);
or U8651 (N_8651,N_7820,N_7392);
nor U8652 (N_8652,N_7455,N_7968);
and U8653 (N_8653,N_7664,N_7636);
or U8654 (N_8654,N_7056,N_7272);
nand U8655 (N_8655,N_7241,N_7343);
nand U8656 (N_8656,N_7395,N_7394);
or U8657 (N_8657,N_7307,N_7309);
nor U8658 (N_8658,N_7191,N_7873);
xnor U8659 (N_8659,N_7170,N_7880);
nand U8660 (N_8660,N_7008,N_7142);
nor U8661 (N_8661,N_7089,N_7790);
and U8662 (N_8662,N_7707,N_7888);
nand U8663 (N_8663,N_7394,N_7338);
and U8664 (N_8664,N_7733,N_7659);
xnor U8665 (N_8665,N_7286,N_7922);
nand U8666 (N_8666,N_7115,N_7888);
nor U8667 (N_8667,N_7724,N_7596);
nand U8668 (N_8668,N_7510,N_7841);
nor U8669 (N_8669,N_7436,N_7541);
xnor U8670 (N_8670,N_7888,N_7798);
nor U8671 (N_8671,N_7318,N_7802);
nor U8672 (N_8672,N_7022,N_7754);
xnor U8673 (N_8673,N_7871,N_7564);
nor U8674 (N_8674,N_7698,N_7706);
nand U8675 (N_8675,N_7181,N_7652);
nor U8676 (N_8676,N_7870,N_7536);
xnor U8677 (N_8677,N_7826,N_7797);
xor U8678 (N_8678,N_7895,N_7787);
xnor U8679 (N_8679,N_7375,N_7045);
or U8680 (N_8680,N_7910,N_7448);
xnor U8681 (N_8681,N_7877,N_7206);
and U8682 (N_8682,N_7323,N_7369);
nor U8683 (N_8683,N_7721,N_7831);
or U8684 (N_8684,N_7710,N_7615);
nor U8685 (N_8685,N_7385,N_7115);
nand U8686 (N_8686,N_7068,N_7382);
nand U8687 (N_8687,N_7113,N_7913);
or U8688 (N_8688,N_7097,N_7959);
xnor U8689 (N_8689,N_7023,N_7509);
xor U8690 (N_8690,N_7073,N_7572);
and U8691 (N_8691,N_7239,N_7427);
and U8692 (N_8692,N_7269,N_7452);
nor U8693 (N_8693,N_7312,N_7070);
and U8694 (N_8694,N_7061,N_7352);
xor U8695 (N_8695,N_7099,N_7480);
or U8696 (N_8696,N_7061,N_7482);
nand U8697 (N_8697,N_7267,N_7634);
and U8698 (N_8698,N_7436,N_7325);
xor U8699 (N_8699,N_7482,N_7375);
xnor U8700 (N_8700,N_7404,N_7483);
and U8701 (N_8701,N_7667,N_7217);
and U8702 (N_8702,N_7295,N_7281);
and U8703 (N_8703,N_7714,N_7870);
or U8704 (N_8704,N_7469,N_7997);
nor U8705 (N_8705,N_7252,N_7258);
or U8706 (N_8706,N_7839,N_7546);
nand U8707 (N_8707,N_7857,N_7910);
or U8708 (N_8708,N_7831,N_7311);
xnor U8709 (N_8709,N_7597,N_7751);
nand U8710 (N_8710,N_7223,N_7370);
xor U8711 (N_8711,N_7523,N_7916);
xor U8712 (N_8712,N_7118,N_7071);
nand U8713 (N_8713,N_7286,N_7882);
xor U8714 (N_8714,N_7127,N_7824);
xor U8715 (N_8715,N_7725,N_7005);
nor U8716 (N_8716,N_7959,N_7168);
or U8717 (N_8717,N_7620,N_7986);
or U8718 (N_8718,N_7282,N_7453);
nand U8719 (N_8719,N_7472,N_7307);
or U8720 (N_8720,N_7598,N_7243);
and U8721 (N_8721,N_7760,N_7774);
or U8722 (N_8722,N_7217,N_7972);
and U8723 (N_8723,N_7702,N_7618);
or U8724 (N_8724,N_7061,N_7931);
nand U8725 (N_8725,N_7858,N_7550);
or U8726 (N_8726,N_7210,N_7945);
and U8727 (N_8727,N_7744,N_7961);
xor U8728 (N_8728,N_7392,N_7018);
xor U8729 (N_8729,N_7666,N_7867);
nor U8730 (N_8730,N_7430,N_7061);
or U8731 (N_8731,N_7198,N_7329);
nor U8732 (N_8732,N_7795,N_7836);
and U8733 (N_8733,N_7641,N_7464);
or U8734 (N_8734,N_7631,N_7666);
and U8735 (N_8735,N_7463,N_7722);
nand U8736 (N_8736,N_7697,N_7061);
xnor U8737 (N_8737,N_7933,N_7597);
and U8738 (N_8738,N_7757,N_7581);
nor U8739 (N_8739,N_7379,N_7342);
xor U8740 (N_8740,N_7644,N_7497);
xor U8741 (N_8741,N_7106,N_7308);
nand U8742 (N_8742,N_7587,N_7252);
nand U8743 (N_8743,N_7641,N_7548);
and U8744 (N_8744,N_7761,N_7244);
and U8745 (N_8745,N_7961,N_7226);
nand U8746 (N_8746,N_7459,N_7134);
or U8747 (N_8747,N_7529,N_7380);
and U8748 (N_8748,N_7316,N_7798);
nand U8749 (N_8749,N_7536,N_7202);
or U8750 (N_8750,N_7850,N_7016);
xor U8751 (N_8751,N_7740,N_7998);
xor U8752 (N_8752,N_7351,N_7232);
nand U8753 (N_8753,N_7937,N_7179);
xor U8754 (N_8754,N_7330,N_7782);
nand U8755 (N_8755,N_7079,N_7839);
xor U8756 (N_8756,N_7969,N_7846);
xnor U8757 (N_8757,N_7938,N_7682);
nand U8758 (N_8758,N_7325,N_7789);
nor U8759 (N_8759,N_7290,N_7794);
nor U8760 (N_8760,N_7695,N_7565);
xor U8761 (N_8761,N_7362,N_7096);
xnor U8762 (N_8762,N_7454,N_7516);
and U8763 (N_8763,N_7914,N_7780);
nor U8764 (N_8764,N_7375,N_7036);
xnor U8765 (N_8765,N_7442,N_7258);
xnor U8766 (N_8766,N_7192,N_7250);
and U8767 (N_8767,N_7999,N_7513);
nand U8768 (N_8768,N_7204,N_7241);
xor U8769 (N_8769,N_7201,N_7805);
or U8770 (N_8770,N_7861,N_7105);
xor U8771 (N_8771,N_7141,N_7383);
nor U8772 (N_8772,N_7916,N_7202);
nand U8773 (N_8773,N_7401,N_7973);
and U8774 (N_8774,N_7983,N_7902);
nand U8775 (N_8775,N_7487,N_7969);
xnor U8776 (N_8776,N_7649,N_7664);
nor U8777 (N_8777,N_7112,N_7904);
or U8778 (N_8778,N_7049,N_7860);
nand U8779 (N_8779,N_7754,N_7251);
or U8780 (N_8780,N_7792,N_7765);
or U8781 (N_8781,N_7507,N_7861);
nor U8782 (N_8782,N_7858,N_7486);
nor U8783 (N_8783,N_7283,N_7871);
xor U8784 (N_8784,N_7852,N_7628);
nor U8785 (N_8785,N_7421,N_7174);
and U8786 (N_8786,N_7114,N_7499);
nand U8787 (N_8787,N_7914,N_7708);
xor U8788 (N_8788,N_7556,N_7635);
nor U8789 (N_8789,N_7230,N_7592);
nor U8790 (N_8790,N_7667,N_7888);
and U8791 (N_8791,N_7272,N_7050);
or U8792 (N_8792,N_7059,N_7067);
xor U8793 (N_8793,N_7093,N_7454);
and U8794 (N_8794,N_7779,N_7960);
or U8795 (N_8795,N_7119,N_7148);
nor U8796 (N_8796,N_7190,N_7324);
or U8797 (N_8797,N_7038,N_7567);
nor U8798 (N_8798,N_7637,N_7661);
xnor U8799 (N_8799,N_7000,N_7541);
nor U8800 (N_8800,N_7782,N_7612);
nand U8801 (N_8801,N_7842,N_7130);
xor U8802 (N_8802,N_7427,N_7027);
and U8803 (N_8803,N_7769,N_7572);
nor U8804 (N_8804,N_7188,N_7311);
xnor U8805 (N_8805,N_7676,N_7284);
xnor U8806 (N_8806,N_7710,N_7471);
xor U8807 (N_8807,N_7191,N_7034);
nor U8808 (N_8808,N_7480,N_7821);
xnor U8809 (N_8809,N_7351,N_7217);
nor U8810 (N_8810,N_7844,N_7659);
xnor U8811 (N_8811,N_7555,N_7128);
or U8812 (N_8812,N_7693,N_7978);
nor U8813 (N_8813,N_7925,N_7794);
or U8814 (N_8814,N_7259,N_7749);
and U8815 (N_8815,N_7036,N_7457);
or U8816 (N_8816,N_7876,N_7378);
and U8817 (N_8817,N_7456,N_7479);
nand U8818 (N_8818,N_7541,N_7485);
or U8819 (N_8819,N_7499,N_7509);
nand U8820 (N_8820,N_7726,N_7722);
nand U8821 (N_8821,N_7444,N_7072);
xnor U8822 (N_8822,N_7002,N_7144);
and U8823 (N_8823,N_7008,N_7217);
xor U8824 (N_8824,N_7190,N_7192);
nor U8825 (N_8825,N_7633,N_7110);
nand U8826 (N_8826,N_7794,N_7577);
and U8827 (N_8827,N_7585,N_7511);
or U8828 (N_8828,N_7357,N_7788);
xnor U8829 (N_8829,N_7055,N_7960);
and U8830 (N_8830,N_7021,N_7743);
xnor U8831 (N_8831,N_7794,N_7360);
or U8832 (N_8832,N_7472,N_7517);
nand U8833 (N_8833,N_7197,N_7325);
nand U8834 (N_8834,N_7593,N_7007);
or U8835 (N_8835,N_7107,N_7179);
or U8836 (N_8836,N_7937,N_7743);
and U8837 (N_8837,N_7560,N_7381);
nor U8838 (N_8838,N_7972,N_7664);
or U8839 (N_8839,N_7297,N_7816);
or U8840 (N_8840,N_7917,N_7065);
nor U8841 (N_8841,N_7054,N_7357);
and U8842 (N_8842,N_7131,N_7410);
xor U8843 (N_8843,N_7790,N_7707);
or U8844 (N_8844,N_7333,N_7143);
or U8845 (N_8845,N_7438,N_7439);
xnor U8846 (N_8846,N_7576,N_7433);
or U8847 (N_8847,N_7161,N_7771);
xnor U8848 (N_8848,N_7352,N_7383);
xor U8849 (N_8849,N_7369,N_7141);
nand U8850 (N_8850,N_7106,N_7179);
xor U8851 (N_8851,N_7826,N_7149);
and U8852 (N_8852,N_7974,N_7394);
xor U8853 (N_8853,N_7626,N_7909);
nor U8854 (N_8854,N_7803,N_7151);
nand U8855 (N_8855,N_7492,N_7701);
and U8856 (N_8856,N_7091,N_7767);
nand U8857 (N_8857,N_7393,N_7955);
or U8858 (N_8858,N_7628,N_7580);
nand U8859 (N_8859,N_7951,N_7984);
and U8860 (N_8860,N_7843,N_7454);
xor U8861 (N_8861,N_7431,N_7577);
or U8862 (N_8862,N_7589,N_7071);
xnor U8863 (N_8863,N_7169,N_7893);
nand U8864 (N_8864,N_7886,N_7209);
or U8865 (N_8865,N_7489,N_7613);
xor U8866 (N_8866,N_7865,N_7231);
xor U8867 (N_8867,N_7158,N_7816);
and U8868 (N_8868,N_7172,N_7854);
xor U8869 (N_8869,N_7232,N_7100);
nor U8870 (N_8870,N_7971,N_7663);
xnor U8871 (N_8871,N_7947,N_7120);
xnor U8872 (N_8872,N_7529,N_7942);
or U8873 (N_8873,N_7235,N_7930);
and U8874 (N_8874,N_7313,N_7783);
or U8875 (N_8875,N_7227,N_7301);
or U8876 (N_8876,N_7726,N_7252);
nor U8877 (N_8877,N_7925,N_7842);
xor U8878 (N_8878,N_7583,N_7584);
xor U8879 (N_8879,N_7124,N_7524);
nor U8880 (N_8880,N_7724,N_7042);
nor U8881 (N_8881,N_7204,N_7895);
and U8882 (N_8882,N_7903,N_7234);
and U8883 (N_8883,N_7160,N_7851);
xor U8884 (N_8884,N_7925,N_7560);
nand U8885 (N_8885,N_7890,N_7986);
and U8886 (N_8886,N_7447,N_7579);
nor U8887 (N_8887,N_7449,N_7943);
or U8888 (N_8888,N_7971,N_7368);
nand U8889 (N_8889,N_7782,N_7104);
or U8890 (N_8890,N_7036,N_7736);
xnor U8891 (N_8891,N_7237,N_7915);
or U8892 (N_8892,N_7436,N_7034);
nand U8893 (N_8893,N_7417,N_7139);
nand U8894 (N_8894,N_7858,N_7538);
or U8895 (N_8895,N_7049,N_7310);
and U8896 (N_8896,N_7343,N_7301);
xor U8897 (N_8897,N_7727,N_7247);
or U8898 (N_8898,N_7011,N_7692);
nand U8899 (N_8899,N_7577,N_7304);
xnor U8900 (N_8900,N_7030,N_7170);
nor U8901 (N_8901,N_7151,N_7268);
and U8902 (N_8902,N_7907,N_7166);
xor U8903 (N_8903,N_7600,N_7288);
and U8904 (N_8904,N_7352,N_7936);
and U8905 (N_8905,N_7901,N_7131);
nand U8906 (N_8906,N_7275,N_7619);
xnor U8907 (N_8907,N_7298,N_7056);
nor U8908 (N_8908,N_7337,N_7299);
xnor U8909 (N_8909,N_7425,N_7819);
xor U8910 (N_8910,N_7423,N_7642);
and U8911 (N_8911,N_7572,N_7256);
and U8912 (N_8912,N_7342,N_7763);
or U8913 (N_8913,N_7743,N_7981);
or U8914 (N_8914,N_7770,N_7573);
xnor U8915 (N_8915,N_7024,N_7288);
and U8916 (N_8916,N_7109,N_7192);
xor U8917 (N_8917,N_7927,N_7799);
and U8918 (N_8918,N_7748,N_7625);
xor U8919 (N_8919,N_7960,N_7908);
nor U8920 (N_8920,N_7870,N_7459);
or U8921 (N_8921,N_7894,N_7139);
xor U8922 (N_8922,N_7718,N_7912);
and U8923 (N_8923,N_7560,N_7204);
nand U8924 (N_8924,N_7018,N_7802);
or U8925 (N_8925,N_7713,N_7443);
nand U8926 (N_8926,N_7514,N_7085);
or U8927 (N_8927,N_7923,N_7634);
xor U8928 (N_8928,N_7533,N_7298);
xor U8929 (N_8929,N_7374,N_7437);
and U8930 (N_8930,N_7313,N_7434);
xor U8931 (N_8931,N_7531,N_7964);
nor U8932 (N_8932,N_7936,N_7457);
or U8933 (N_8933,N_7391,N_7812);
nand U8934 (N_8934,N_7021,N_7356);
nor U8935 (N_8935,N_7128,N_7497);
and U8936 (N_8936,N_7987,N_7179);
nand U8937 (N_8937,N_7163,N_7767);
nand U8938 (N_8938,N_7515,N_7633);
and U8939 (N_8939,N_7130,N_7402);
xor U8940 (N_8940,N_7948,N_7621);
nand U8941 (N_8941,N_7693,N_7490);
nand U8942 (N_8942,N_7539,N_7627);
or U8943 (N_8943,N_7354,N_7552);
or U8944 (N_8944,N_7504,N_7008);
or U8945 (N_8945,N_7298,N_7596);
or U8946 (N_8946,N_7315,N_7299);
xnor U8947 (N_8947,N_7631,N_7945);
or U8948 (N_8948,N_7563,N_7745);
and U8949 (N_8949,N_7483,N_7747);
and U8950 (N_8950,N_7600,N_7630);
nand U8951 (N_8951,N_7494,N_7931);
or U8952 (N_8952,N_7562,N_7997);
nor U8953 (N_8953,N_7227,N_7056);
nand U8954 (N_8954,N_7067,N_7857);
nor U8955 (N_8955,N_7211,N_7314);
and U8956 (N_8956,N_7863,N_7592);
nor U8957 (N_8957,N_7523,N_7898);
nand U8958 (N_8958,N_7790,N_7664);
nor U8959 (N_8959,N_7469,N_7996);
nor U8960 (N_8960,N_7029,N_7832);
or U8961 (N_8961,N_7930,N_7748);
nor U8962 (N_8962,N_7520,N_7627);
and U8963 (N_8963,N_7761,N_7926);
xor U8964 (N_8964,N_7456,N_7457);
nor U8965 (N_8965,N_7190,N_7745);
and U8966 (N_8966,N_7132,N_7103);
or U8967 (N_8967,N_7100,N_7807);
xor U8968 (N_8968,N_7625,N_7194);
xnor U8969 (N_8969,N_7985,N_7979);
and U8970 (N_8970,N_7368,N_7962);
nor U8971 (N_8971,N_7732,N_7262);
or U8972 (N_8972,N_7770,N_7675);
and U8973 (N_8973,N_7536,N_7221);
nand U8974 (N_8974,N_7788,N_7479);
xnor U8975 (N_8975,N_7540,N_7361);
nor U8976 (N_8976,N_7220,N_7659);
xor U8977 (N_8977,N_7094,N_7983);
nor U8978 (N_8978,N_7614,N_7915);
or U8979 (N_8979,N_7035,N_7331);
or U8980 (N_8980,N_7020,N_7993);
or U8981 (N_8981,N_7348,N_7308);
nor U8982 (N_8982,N_7509,N_7053);
or U8983 (N_8983,N_7704,N_7187);
xnor U8984 (N_8984,N_7906,N_7827);
nand U8985 (N_8985,N_7816,N_7065);
nand U8986 (N_8986,N_7687,N_7251);
nand U8987 (N_8987,N_7035,N_7608);
and U8988 (N_8988,N_7687,N_7800);
xor U8989 (N_8989,N_7821,N_7159);
nand U8990 (N_8990,N_7551,N_7650);
nand U8991 (N_8991,N_7639,N_7945);
and U8992 (N_8992,N_7972,N_7767);
or U8993 (N_8993,N_7885,N_7832);
and U8994 (N_8994,N_7613,N_7072);
or U8995 (N_8995,N_7665,N_7686);
or U8996 (N_8996,N_7549,N_7878);
nand U8997 (N_8997,N_7870,N_7141);
xnor U8998 (N_8998,N_7610,N_7986);
xor U8999 (N_8999,N_7022,N_7376);
nor U9000 (N_9000,N_8540,N_8324);
or U9001 (N_9001,N_8495,N_8979);
nand U9002 (N_9002,N_8021,N_8816);
nand U9003 (N_9003,N_8125,N_8367);
and U9004 (N_9004,N_8048,N_8394);
nand U9005 (N_9005,N_8253,N_8607);
nor U9006 (N_9006,N_8918,N_8202);
and U9007 (N_9007,N_8981,N_8598);
or U9008 (N_9008,N_8881,N_8501);
or U9009 (N_9009,N_8600,N_8705);
xor U9010 (N_9010,N_8387,N_8870);
nand U9011 (N_9011,N_8409,N_8817);
nand U9012 (N_9012,N_8217,N_8086);
nor U9013 (N_9013,N_8199,N_8397);
nor U9014 (N_9014,N_8398,N_8335);
and U9015 (N_9015,N_8123,N_8514);
or U9016 (N_9016,N_8887,N_8510);
xnor U9017 (N_9017,N_8458,N_8189);
nor U9018 (N_9018,N_8908,N_8952);
or U9019 (N_9019,N_8194,N_8126);
nand U9020 (N_9020,N_8522,N_8005);
xnor U9021 (N_9021,N_8143,N_8803);
nand U9022 (N_9022,N_8873,N_8897);
xor U9023 (N_9023,N_8186,N_8311);
nor U9024 (N_9024,N_8808,N_8699);
nor U9025 (N_9025,N_8532,N_8434);
and U9026 (N_9026,N_8275,N_8382);
and U9027 (N_9027,N_8717,N_8737);
nand U9028 (N_9028,N_8450,N_8622);
xnor U9029 (N_9029,N_8488,N_8401);
nor U9030 (N_9030,N_8337,N_8754);
nand U9031 (N_9031,N_8082,N_8869);
and U9032 (N_9032,N_8057,N_8166);
and U9033 (N_9033,N_8624,N_8861);
xnor U9034 (N_9034,N_8513,N_8019);
nand U9035 (N_9035,N_8593,N_8637);
and U9036 (N_9036,N_8411,N_8316);
xnor U9037 (N_9037,N_8105,N_8489);
xnor U9038 (N_9038,N_8215,N_8378);
or U9039 (N_9039,N_8960,N_8493);
nor U9040 (N_9040,N_8693,N_8244);
or U9041 (N_9041,N_8366,N_8516);
and U9042 (N_9042,N_8216,N_8565);
nand U9043 (N_9043,N_8414,N_8563);
or U9044 (N_9044,N_8708,N_8961);
xor U9045 (N_9045,N_8174,N_8201);
nor U9046 (N_9046,N_8261,N_8212);
nand U9047 (N_9047,N_8996,N_8172);
nor U9048 (N_9048,N_8112,N_8904);
nand U9049 (N_9049,N_8104,N_8884);
and U9050 (N_9050,N_8278,N_8103);
xor U9051 (N_9051,N_8913,N_8950);
and U9052 (N_9052,N_8994,N_8219);
nor U9053 (N_9053,N_8702,N_8851);
xnor U9054 (N_9054,N_8121,N_8774);
nand U9055 (N_9055,N_8460,N_8403);
nor U9056 (N_9056,N_8056,N_8505);
nor U9057 (N_9057,N_8590,N_8257);
and U9058 (N_9058,N_8896,N_8660);
nor U9059 (N_9059,N_8033,N_8597);
nor U9060 (N_9060,N_8667,N_8188);
nand U9061 (N_9061,N_8964,N_8471);
nand U9062 (N_9062,N_8207,N_8814);
nand U9063 (N_9063,N_8351,N_8615);
xnor U9064 (N_9064,N_8346,N_8308);
nand U9065 (N_9065,N_8511,N_8746);
xor U9066 (N_9066,N_8003,N_8327);
and U9067 (N_9067,N_8046,N_8646);
nor U9068 (N_9068,N_8425,N_8974);
nand U9069 (N_9069,N_8771,N_8862);
and U9070 (N_9070,N_8154,N_8901);
xor U9071 (N_9071,N_8921,N_8858);
and U9072 (N_9072,N_8476,N_8907);
nand U9073 (N_9073,N_8825,N_8747);
or U9074 (N_9074,N_8148,N_8496);
nand U9075 (N_9075,N_8878,N_8250);
nand U9076 (N_9076,N_8359,N_8684);
nand U9077 (N_9077,N_8054,N_8799);
nor U9078 (N_9078,N_8534,N_8474);
xnor U9079 (N_9079,N_8765,N_8785);
xor U9080 (N_9080,N_8138,N_8070);
and U9081 (N_9081,N_8585,N_8305);
xnor U9082 (N_9082,N_8139,N_8779);
nand U9083 (N_9083,N_8859,N_8567);
and U9084 (N_9084,N_8776,N_8420);
nand U9085 (N_9085,N_8323,N_8834);
or U9086 (N_9086,N_8784,N_8947);
nor U9087 (N_9087,N_8587,N_8821);
nor U9088 (N_9088,N_8438,N_8628);
nor U9089 (N_9089,N_8369,N_8014);
nor U9090 (N_9090,N_8772,N_8299);
or U9091 (N_9091,N_8355,N_8022);
nand U9092 (N_9092,N_8927,N_8617);
nand U9093 (N_9093,N_8012,N_8594);
xor U9094 (N_9094,N_8109,N_8936);
nand U9095 (N_9095,N_8446,N_8910);
nand U9096 (N_9096,N_8924,N_8318);
nand U9097 (N_9097,N_8042,N_8130);
nor U9098 (N_9098,N_8868,N_8214);
nor U9099 (N_9099,N_8578,N_8704);
nand U9100 (N_9100,N_8963,N_8399);
or U9101 (N_9101,N_8065,N_8179);
nand U9102 (N_9102,N_8447,N_8011);
nand U9103 (N_9103,N_8762,N_8051);
nor U9104 (N_9104,N_8620,N_8644);
nor U9105 (N_9105,N_8716,N_8156);
and U9106 (N_9106,N_8674,N_8454);
and U9107 (N_9107,N_8502,N_8701);
nor U9108 (N_9108,N_8309,N_8601);
or U9109 (N_9109,N_8481,N_8743);
or U9110 (N_9110,N_8364,N_8016);
or U9111 (N_9111,N_8824,N_8358);
xnor U9112 (N_9112,N_8835,N_8004);
and U9113 (N_9113,N_8856,N_8204);
xor U9114 (N_9114,N_8240,N_8722);
xnor U9115 (N_9115,N_8052,N_8020);
xor U9116 (N_9116,N_8114,N_8231);
or U9117 (N_9117,N_8827,N_8891);
nand U9118 (N_9118,N_8857,N_8755);
nor U9119 (N_9119,N_8494,N_8234);
nor U9120 (N_9120,N_8549,N_8060);
nand U9121 (N_9121,N_8256,N_8221);
or U9122 (N_9122,N_8725,N_8676);
xor U9123 (N_9123,N_8252,N_8338);
xor U9124 (N_9124,N_8006,N_8357);
xor U9125 (N_9125,N_8304,N_8491);
and U9126 (N_9126,N_8553,N_8110);
or U9127 (N_9127,N_8889,N_8745);
xor U9128 (N_9128,N_8595,N_8241);
nor U9129 (N_9129,N_8026,N_8182);
nor U9130 (N_9130,N_8649,N_8749);
xor U9131 (N_9131,N_8180,N_8662);
and U9132 (N_9132,N_8322,N_8625);
nand U9133 (N_9133,N_8426,N_8223);
nor U9134 (N_9134,N_8937,N_8018);
nand U9135 (N_9135,N_8621,N_8354);
nor U9136 (N_9136,N_8059,N_8064);
xnor U9137 (N_9137,N_8612,N_8572);
or U9138 (N_9138,N_8589,N_8376);
nor U9139 (N_9139,N_8102,N_8744);
xor U9140 (N_9140,N_8766,N_8657);
xor U9141 (N_9141,N_8757,N_8957);
and U9142 (N_9142,N_8912,N_8271);
or U9143 (N_9143,N_8506,N_8599);
nor U9144 (N_9144,N_8412,N_8332);
and U9145 (N_9145,N_8696,N_8120);
nand U9146 (N_9146,N_8473,N_8678);
or U9147 (N_9147,N_8789,N_8523);
and U9148 (N_9148,N_8984,N_8047);
nand U9149 (N_9149,N_8552,N_8395);
and U9150 (N_9150,N_8062,N_8209);
and U9151 (N_9151,N_8078,N_8437);
xor U9152 (N_9152,N_8160,N_8239);
nand U9153 (N_9153,N_8805,N_8988);
xnor U9154 (N_9154,N_8456,N_8431);
and U9155 (N_9155,N_8185,N_8571);
nor U9156 (N_9156,N_8373,N_8880);
nor U9157 (N_9157,N_8976,N_8142);
xor U9158 (N_9158,N_8486,N_8654);
and U9159 (N_9159,N_8575,N_8117);
or U9160 (N_9160,N_8811,N_8392);
xor U9161 (N_9161,N_8883,N_8507);
nor U9162 (N_9162,N_8002,N_8876);
nor U9163 (N_9163,N_8832,N_8273);
nor U9164 (N_9164,N_8475,N_8459);
or U9165 (N_9165,N_8410,N_8153);
nand U9166 (N_9166,N_8030,N_8238);
and U9167 (N_9167,N_8661,N_8728);
nor U9168 (N_9168,N_8529,N_8379);
nor U9169 (N_9169,N_8085,N_8158);
nor U9170 (N_9170,N_8652,N_8890);
or U9171 (N_9171,N_8849,N_8417);
nor U9172 (N_9172,N_8769,N_8246);
nand U9173 (N_9173,N_8451,N_8647);
nand U9174 (N_9174,N_8569,N_8951);
and U9175 (N_9175,N_8967,N_8993);
and U9176 (N_9176,N_8756,N_8067);
nand U9177 (N_9177,N_8365,N_8719);
nor U9178 (N_9178,N_8551,N_8902);
or U9179 (N_9179,N_8101,N_8445);
nand U9180 (N_9180,N_8455,N_8340);
nand U9181 (N_9181,N_8732,N_8429);
xor U9182 (N_9182,N_8911,N_8822);
or U9183 (N_9183,N_8049,N_8225);
and U9184 (N_9184,N_8886,N_8838);
nand U9185 (N_9185,N_8132,N_8758);
or U9186 (N_9186,N_8797,N_8282);
xor U9187 (N_9187,N_8509,N_8222);
and U9188 (N_9188,N_8916,N_8260);
or U9189 (N_9189,N_8462,N_8436);
nor U9190 (N_9190,N_8404,N_8605);
or U9191 (N_9191,N_8263,N_8955);
xnor U9192 (N_9192,N_8350,N_8543);
and U9193 (N_9193,N_8579,N_8203);
nor U9194 (N_9194,N_8470,N_8711);
nand U9195 (N_9195,N_8925,N_8008);
xnor U9196 (N_9196,N_8794,N_8267);
nand U9197 (N_9197,N_8694,N_8424);
or U9198 (N_9198,N_8363,N_8682);
or U9199 (N_9199,N_8592,N_8508);
and U9200 (N_9200,N_8812,N_8770);
nand U9201 (N_9201,N_8570,N_8609);
nor U9202 (N_9202,N_8945,N_8413);
nand U9203 (N_9203,N_8650,N_8229);
xor U9204 (N_9204,N_8653,N_8632);
xnor U9205 (N_9205,N_8196,N_8091);
nand U9206 (N_9206,N_8007,N_8530);
or U9207 (N_9207,N_8141,N_8251);
xor U9208 (N_9208,N_8561,N_8798);
nand U9209 (N_9209,N_8800,N_8089);
or U9210 (N_9210,N_8150,N_8991);
nand U9211 (N_9211,N_8129,N_8035);
or U9212 (N_9212,N_8917,N_8272);
or U9213 (N_9213,N_8029,N_8761);
nand U9214 (N_9214,N_8277,N_8736);
and U9215 (N_9215,N_8027,N_8407);
or U9216 (N_9216,N_8715,N_8683);
nand U9217 (N_9217,N_8131,N_8844);
and U9218 (N_9218,N_8293,N_8145);
or U9219 (N_9219,N_8689,N_8804);
xor U9220 (N_9220,N_8441,N_8058);
xnor U9221 (N_9221,N_8288,N_8793);
and U9222 (N_9222,N_8813,N_8767);
nand U9223 (N_9223,N_8232,N_8959);
or U9224 (N_9224,N_8381,N_8384);
xnor U9225 (N_9225,N_8941,N_8442);
nand U9226 (N_9226,N_8727,N_8464);
and U9227 (N_9227,N_8707,N_8712);
xnor U9228 (N_9228,N_8692,N_8671);
nor U9229 (N_9229,N_8205,N_8349);
nor U9230 (N_9230,N_8448,N_8393);
nor U9231 (N_9231,N_8792,N_8919);
or U9232 (N_9232,N_8619,N_8479);
and U9233 (N_9233,N_8371,N_8564);
xor U9234 (N_9234,N_8069,N_8391);
and U9235 (N_9235,N_8839,N_8882);
nor U9236 (N_9236,N_8230,N_8374);
nor U9237 (N_9237,N_8245,N_8562);
nand U9238 (N_9238,N_8247,N_8266);
nand U9239 (N_9239,N_8806,N_8533);
or U9240 (N_9240,N_8922,N_8985);
or U9241 (N_9241,N_8405,N_8721);
and U9242 (N_9242,N_8954,N_8328);
nand U9243 (N_9243,N_8764,N_8140);
or U9244 (N_9244,N_8249,N_8815);
xnor U9245 (N_9245,N_8433,N_8942);
or U9246 (N_9246,N_8929,N_8164);
xnor U9247 (N_9247,N_8935,N_8852);
and U9248 (N_9248,N_8790,N_8482);
and U9249 (N_9249,N_8220,N_8934);
nand U9250 (N_9250,N_8170,N_8894);
or U9251 (N_9251,N_8648,N_8990);
nor U9252 (N_9252,N_8738,N_8828);
xnor U9253 (N_9253,N_8187,N_8877);
nand U9254 (N_9254,N_8968,N_8375);
xnor U9255 (N_9255,N_8276,N_8163);
and U9256 (N_9256,N_8487,N_8149);
xnor U9257 (N_9257,N_8040,N_8422);
xor U9258 (N_9258,N_8467,N_8780);
nor U9259 (N_9259,N_8541,N_8698);
xor U9260 (N_9260,N_8372,N_8439);
xor U9261 (N_9261,N_8243,N_8184);
or U9262 (N_9262,N_8146,N_8173);
xor U9263 (N_9263,N_8402,N_8453);
and U9264 (N_9264,N_8210,N_8932);
and U9265 (N_9265,N_8097,N_8666);
nor U9266 (N_9266,N_8321,N_8385);
xor U9267 (N_9267,N_8080,N_8301);
xnor U9268 (N_9268,N_8759,N_8183);
nor U9269 (N_9269,N_8037,N_8686);
nand U9270 (N_9270,N_8748,N_8226);
xnor U9271 (N_9271,N_8206,N_8900);
and U9272 (N_9272,N_8400,N_8171);
nor U9273 (N_9273,N_8075,N_8665);
nor U9274 (N_9274,N_8452,N_8457);
nor U9275 (N_9275,N_8015,N_8608);
or U9276 (N_9276,N_8076,N_8281);
nand U9277 (N_9277,N_8289,N_8830);
and U9278 (N_9278,N_8041,N_8500);
and U9279 (N_9279,N_8840,N_8307);
nand U9280 (N_9280,N_8630,N_8591);
and U9281 (N_9281,N_8837,N_8681);
and U9282 (N_9282,N_8083,N_8664);
xor U9283 (N_9283,N_8915,N_8953);
or U9284 (N_9284,N_8368,N_8264);
or U9285 (N_9285,N_8108,N_8558);
or U9286 (N_9286,N_8545,N_8973);
xor U9287 (N_9287,N_8997,N_8001);
nand U9288 (N_9288,N_8312,N_8833);
xnor U9289 (N_9289,N_8053,N_8415);
nor U9290 (N_9290,N_8290,N_8478);
xnor U9291 (N_9291,N_8291,N_8144);
nand U9292 (N_9292,N_8819,N_8284);
nor U9293 (N_9293,N_8867,N_8344);
or U9294 (N_9294,N_8962,N_8408);
nor U9295 (N_9295,N_8864,N_8136);
xnor U9296 (N_9296,N_8497,N_8325);
nand U9297 (N_9297,N_8675,N_8836);
xor U9298 (N_9298,N_8866,N_8406);
nand U9299 (N_9299,N_8634,N_8228);
and U9300 (N_9300,N_8208,N_8390);
xnor U9301 (N_9301,N_8658,N_8465);
nor U9302 (N_9302,N_8641,N_8262);
nand U9303 (N_9303,N_8559,N_8099);
or U9304 (N_9304,N_8259,N_8469);
and U9305 (N_9305,N_8706,N_8602);
and U9306 (N_9306,N_8731,N_8610);
and U9307 (N_9307,N_8720,N_8389);
xnor U9308 (N_9308,N_8874,N_8557);
and U9309 (N_9309,N_8775,N_8419);
or U9310 (N_9310,N_8872,N_8377);
nor U9311 (N_9311,N_8227,N_8848);
nand U9312 (N_9312,N_8198,N_8865);
or U9313 (N_9313,N_8440,N_8636);
or U9314 (N_9314,N_8023,N_8948);
nor U9315 (N_9315,N_8842,N_8544);
xnor U9316 (N_9316,N_8733,N_8192);
or U9317 (N_9317,N_8695,N_8635);
xor U9318 (N_9318,N_8485,N_8643);
nor U9319 (N_9319,N_8697,N_8560);
nor U9320 (N_9320,N_8061,N_8127);
and U9321 (N_9321,N_8669,N_8236);
nand U9322 (N_9322,N_8383,N_8656);
nor U9323 (N_9323,N_8159,N_8483);
xor U9324 (N_9324,N_8193,N_8200);
xor U9325 (N_9325,N_8729,N_8971);
nor U9326 (N_9326,N_8539,N_8124);
xnor U9327 (N_9327,N_8845,N_8038);
nor U9328 (N_9328,N_8663,N_8361);
and U9329 (N_9329,N_8039,N_8317);
xor U9330 (N_9330,N_8155,N_8242);
nor U9331 (N_9331,N_8633,N_8518);
xor U9332 (N_9332,N_8531,N_8034);
or U9333 (N_9333,N_8360,N_8999);
nor U9334 (N_9334,N_8418,N_8168);
nor U9335 (N_9335,N_8255,N_8685);
nand U9336 (N_9336,N_8554,N_8626);
nand U9337 (N_9337,N_8074,N_8463);
nor U9338 (N_9338,N_8568,N_8449);
nor U9339 (N_9339,N_8167,N_8938);
xnor U9340 (N_9340,N_8386,N_8331);
xor U9341 (N_9341,N_8972,N_8970);
nor U9342 (N_9342,N_8098,N_8017);
xnor U9343 (N_9343,N_8169,N_8659);
xnor U9344 (N_9344,N_8892,N_8655);
and U9345 (N_9345,N_8987,N_8863);
nand U9346 (N_9346,N_8546,N_8542);
nor U9347 (N_9347,N_8783,N_8477);
xnor U9348 (N_9348,N_8709,N_8000);
nand U9349 (N_9349,N_8740,N_8499);
xor U9350 (N_9350,N_8843,N_8213);
xnor U9351 (N_9351,N_8137,N_8718);
xor U9352 (N_9352,N_8586,N_8115);
or U9353 (N_9353,N_8965,N_8796);
and U9354 (N_9354,N_8829,N_8092);
nand U9355 (N_9355,N_8781,N_8248);
and U9356 (N_9356,N_8690,N_8432);
nand U9357 (N_9357,N_8352,N_8670);
nand U9358 (N_9358,N_8430,N_8980);
and U9359 (N_9359,N_8691,N_8928);
or U9360 (N_9360,N_8875,N_8280);
xor U9361 (N_9361,N_8818,N_8931);
nand U9362 (N_9362,N_8730,N_8673);
xnor U9363 (N_9363,N_8116,N_8315);
xor U9364 (N_9364,N_8940,N_8298);
xor U9365 (N_9365,N_8472,N_8946);
or U9366 (N_9366,N_8966,N_8978);
xor U9367 (N_9367,N_8254,N_8521);
nor U9368 (N_9368,N_8939,N_8119);
nor U9369 (N_9369,N_8606,N_8975);
nor U9370 (N_9370,N_8898,N_8760);
nor U9371 (N_9371,N_8283,N_8627);
nand U9372 (N_9372,N_8713,N_8093);
nand U9373 (N_9373,N_8314,N_8933);
nor U9374 (N_9374,N_8631,N_8850);
or U9375 (N_9375,N_8871,N_8914);
nor U9376 (N_9376,N_8287,N_8370);
or U9377 (N_9377,N_8700,N_8895);
nand U9378 (N_9378,N_8768,N_8128);
nand U9379 (N_9379,N_8416,N_8032);
nor U9380 (N_9380,N_8677,N_8944);
nand U9381 (N_9381,N_8050,N_8345);
nor U9382 (N_9382,N_8045,N_8161);
or U9383 (N_9383,N_8580,N_8977);
and U9384 (N_9384,N_8009,N_8165);
nand U9385 (N_9385,N_8724,N_8286);
nor U9386 (N_9386,N_8444,N_8274);
nand U9387 (N_9387,N_8503,N_8854);
xnor U9388 (N_9388,N_8787,N_8157);
nand U9389 (N_9389,N_8396,N_8071);
or U9390 (N_9390,N_8319,N_8435);
and U9391 (N_9391,N_8135,N_8548);
or U9392 (N_9392,N_8742,N_8603);
and U9393 (N_9393,N_8888,N_8613);
xnor U9394 (N_9394,N_8639,N_8484);
xnor U9395 (N_9395,N_8909,N_8068);
xor U9396 (N_9396,N_8268,N_8986);
nand U9397 (N_9397,N_8629,N_8788);
nor U9398 (N_9398,N_8336,N_8920);
xnor U9399 (N_9399,N_8292,N_8750);
or U9400 (N_9400,N_8177,N_8958);
nor U9401 (N_9401,N_8714,N_8853);
nand U9402 (N_9402,N_8492,N_8306);
nand U9403 (N_9403,N_8356,N_8823);
or U9404 (N_9404,N_8992,N_8735);
and U9405 (N_9405,N_8342,N_8341);
xnor U9406 (N_9406,N_8846,N_8296);
nor U9407 (N_9407,N_8111,N_8777);
and U9408 (N_9408,N_8703,N_8588);
xor U9409 (N_9409,N_8512,N_8515);
and U9410 (N_9410,N_8031,N_8334);
nand U9411 (N_9411,N_8380,N_8461);
or U9412 (N_9412,N_8982,N_8949);
and U9413 (N_9413,N_8723,N_8573);
xor U9414 (N_9414,N_8751,N_8066);
nand U9415 (N_9415,N_8640,N_8998);
or U9416 (N_9416,N_8339,N_8726);
or U9417 (N_9417,N_8604,N_8094);
or U9418 (N_9418,N_8055,N_8106);
or U9419 (N_9419,N_8147,N_8537);
nor U9420 (N_9420,N_8584,N_8906);
nor U9421 (N_9421,N_8237,N_8320);
nor U9422 (N_9422,N_8044,N_8778);
xor U9423 (N_9423,N_8763,N_8191);
xor U9424 (N_9424,N_8810,N_8923);
nand U9425 (N_9425,N_8480,N_8423);
nor U9426 (N_9426,N_8879,N_8195);
nand U9427 (N_9427,N_8218,N_8388);
or U9428 (N_9428,N_8893,N_8081);
nand U9429 (N_9429,N_8087,N_8343);
nand U9430 (N_9430,N_8073,N_8134);
or U9431 (N_9431,N_8190,N_8826);
or U9432 (N_9432,N_8680,N_8905);
nor U9433 (N_9433,N_8013,N_8943);
or U9434 (N_9434,N_8989,N_8734);
xnor U9435 (N_9435,N_8084,N_8090);
xnor U9436 (N_9436,N_8490,N_8297);
or U9437 (N_9437,N_8072,N_8556);
nand U9438 (N_9438,N_8596,N_8739);
nor U9439 (N_9439,N_8197,N_8795);
or U9440 (N_9440,N_8550,N_8773);
nand U9441 (N_9441,N_8528,N_8362);
nand U9442 (N_9442,N_8847,N_8224);
xnor U9443 (N_9443,N_8801,N_8151);
nor U9444 (N_9444,N_8028,N_8903);
and U9445 (N_9445,N_8427,N_8024);
and U9446 (N_9446,N_8095,N_8524);
xor U9447 (N_9447,N_8983,N_8645);
xnor U9448 (N_9448,N_8113,N_8235);
xor U9449 (N_9449,N_8133,N_8995);
xnor U9450 (N_9450,N_8100,N_8302);
and U9451 (N_9451,N_8538,N_8841);
or U9452 (N_9452,N_8176,N_8079);
nand U9453 (N_9453,N_8178,N_8536);
nand U9454 (N_9454,N_8638,N_8270);
nor U9455 (N_9455,N_8162,N_8581);
or U9456 (N_9456,N_8611,N_8303);
xor U9457 (N_9457,N_8088,N_8258);
nand U9458 (N_9458,N_8300,N_8330);
or U9459 (N_9459,N_8118,N_8468);
and U9460 (N_9460,N_8096,N_8582);
xnor U9461 (N_9461,N_8527,N_8831);
and U9462 (N_9462,N_8519,N_8498);
and U9463 (N_9463,N_8443,N_8265);
xnor U9464 (N_9464,N_8687,N_8025);
or U9465 (N_9465,N_8526,N_8535);
nand U9466 (N_9466,N_8043,N_8623);
nor U9467 (N_9467,N_8574,N_8956);
nor U9468 (N_9468,N_8295,N_8421);
nand U9469 (N_9469,N_8329,N_8791);
and U9470 (N_9470,N_8466,N_8310);
nor U9471 (N_9471,N_8583,N_8525);
nand U9472 (N_9472,N_8651,N_8353);
nand U9473 (N_9473,N_8077,N_8555);
and U9474 (N_9474,N_8930,N_8152);
nand U9475 (N_9475,N_8860,N_8211);
nor U9476 (N_9476,N_8679,N_8269);
xnor U9477 (N_9477,N_8279,N_8855);
nand U9478 (N_9478,N_8741,N_8504);
or U9479 (N_9479,N_8969,N_8614);
or U9480 (N_9480,N_8752,N_8107);
nand U9481 (N_9481,N_8885,N_8122);
nand U9482 (N_9482,N_8175,N_8753);
or U9483 (N_9483,N_8782,N_8517);
xnor U9484 (N_9484,N_8688,N_8802);
and U9485 (N_9485,N_8063,N_8520);
nor U9486 (N_9486,N_8181,N_8348);
nand U9487 (N_9487,N_8326,N_8285);
nor U9488 (N_9488,N_8547,N_8616);
nand U9489 (N_9489,N_8668,N_8618);
and U9490 (N_9490,N_8820,N_8809);
nor U9491 (N_9491,N_8807,N_8313);
or U9492 (N_9492,N_8233,N_8333);
and U9493 (N_9493,N_8566,N_8010);
and U9494 (N_9494,N_8347,N_8428);
xor U9495 (N_9495,N_8899,N_8577);
xnor U9496 (N_9496,N_8642,N_8672);
and U9497 (N_9497,N_8036,N_8710);
xor U9498 (N_9498,N_8294,N_8786);
xnor U9499 (N_9499,N_8576,N_8926);
nor U9500 (N_9500,N_8033,N_8846);
nor U9501 (N_9501,N_8646,N_8267);
and U9502 (N_9502,N_8904,N_8752);
nand U9503 (N_9503,N_8348,N_8162);
nor U9504 (N_9504,N_8671,N_8306);
nor U9505 (N_9505,N_8597,N_8559);
nand U9506 (N_9506,N_8386,N_8056);
or U9507 (N_9507,N_8784,N_8624);
nand U9508 (N_9508,N_8018,N_8365);
nor U9509 (N_9509,N_8672,N_8470);
nor U9510 (N_9510,N_8979,N_8159);
nand U9511 (N_9511,N_8675,N_8834);
or U9512 (N_9512,N_8615,N_8743);
nand U9513 (N_9513,N_8318,N_8300);
nand U9514 (N_9514,N_8080,N_8592);
or U9515 (N_9515,N_8469,N_8938);
or U9516 (N_9516,N_8810,N_8617);
xnor U9517 (N_9517,N_8149,N_8719);
and U9518 (N_9518,N_8509,N_8571);
nor U9519 (N_9519,N_8853,N_8540);
nand U9520 (N_9520,N_8546,N_8486);
nor U9521 (N_9521,N_8706,N_8962);
or U9522 (N_9522,N_8832,N_8327);
or U9523 (N_9523,N_8225,N_8078);
xnor U9524 (N_9524,N_8257,N_8634);
xor U9525 (N_9525,N_8895,N_8361);
xor U9526 (N_9526,N_8767,N_8101);
nand U9527 (N_9527,N_8593,N_8566);
or U9528 (N_9528,N_8769,N_8807);
nor U9529 (N_9529,N_8072,N_8000);
and U9530 (N_9530,N_8300,N_8699);
xnor U9531 (N_9531,N_8042,N_8519);
nand U9532 (N_9532,N_8308,N_8259);
nand U9533 (N_9533,N_8626,N_8397);
nand U9534 (N_9534,N_8915,N_8383);
nor U9535 (N_9535,N_8221,N_8536);
or U9536 (N_9536,N_8952,N_8156);
xnor U9537 (N_9537,N_8129,N_8289);
nand U9538 (N_9538,N_8310,N_8298);
and U9539 (N_9539,N_8394,N_8536);
nand U9540 (N_9540,N_8924,N_8626);
xor U9541 (N_9541,N_8691,N_8907);
or U9542 (N_9542,N_8267,N_8920);
and U9543 (N_9543,N_8773,N_8026);
xnor U9544 (N_9544,N_8636,N_8128);
xor U9545 (N_9545,N_8703,N_8415);
xnor U9546 (N_9546,N_8882,N_8807);
or U9547 (N_9547,N_8105,N_8664);
or U9548 (N_9548,N_8639,N_8703);
or U9549 (N_9549,N_8452,N_8721);
xor U9550 (N_9550,N_8589,N_8524);
nand U9551 (N_9551,N_8470,N_8070);
or U9552 (N_9552,N_8666,N_8398);
or U9553 (N_9553,N_8466,N_8992);
nor U9554 (N_9554,N_8600,N_8535);
or U9555 (N_9555,N_8665,N_8936);
xor U9556 (N_9556,N_8218,N_8485);
nand U9557 (N_9557,N_8212,N_8775);
nand U9558 (N_9558,N_8691,N_8033);
nand U9559 (N_9559,N_8897,N_8214);
and U9560 (N_9560,N_8053,N_8236);
or U9561 (N_9561,N_8434,N_8489);
and U9562 (N_9562,N_8821,N_8172);
xnor U9563 (N_9563,N_8744,N_8119);
nand U9564 (N_9564,N_8533,N_8127);
nor U9565 (N_9565,N_8397,N_8268);
or U9566 (N_9566,N_8832,N_8350);
or U9567 (N_9567,N_8080,N_8320);
nor U9568 (N_9568,N_8679,N_8053);
or U9569 (N_9569,N_8719,N_8310);
nand U9570 (N_9570,N_8107,N_8086);
or U9571 (N_9571,N_8242,N_8274);
or U9572 (N_9572,N_8688,N_8085);
xor U9573 (N_9573,N_8735,N_8689);
or U9574 (N_9574,N_8059,N_8863);
nand U9575 (N_9575,N_8647,N_8320);
nor U9576 (N_9576,N_8286,N_8455);
nor U9577 (N_9577,N_8703,N_8387);
nand U9578 (N_9578,N_8806,N_8985);
nor U9579 (N_9579,N_8983,N_8614);
and U9580 (N_9580,N_8128,N_8272);
and U9581 (N_9581,N_8993,N_8274);
nor U9582 (N_9582,N_8835,N_8478);
or U9583 (N_9583,N_8166,N_8071);
xor U9584 (N_9584,N_8986,N_8627);
nor U9585 (N_9585,N_8459,N_8059);
or U9586 (N_9586,N_8380,N_8425);
or U9587 (N_9587,N_8984,N_8012);
nor U9588 (N_9588,N_8699,N_8440);
xnor U9589 (N_9589,N_8886,N_8098);
nand U9590 (N_9590,N_8779,N_8057);
nand U9591 (N_9591,N_8958,N_8465);
nand U9592 (N_9592,N_8430,N_8141);
nand U9593 (N_9593,N_8287,N_8865);
xnor U9594 (N_9594,N_8081,N_8592);
xnor U9595 (N_9595,N_8798,N_8471);
and U9596 (N_9596,N_8902,N_8806);
xnor U9597 (N_9597,N_8024,N_8822);
xor U9598 (N_9598,N_8505,N_8612);
or U9599 (N_9599,N_8665,N_8921);
nand U9600 (N_9600,N_8763,N_8080);
nand U9601 (N_9601,N_8642,N_8618);
nor U9602 (N_9602,N_8007,N_8996);
and U9603 (N_9603,N_8568,N_8553);
and U9604 (N_9604,N_8215,N_8711);
and U9605 (N_9605,N_8932,N_8966);
or U9606 (N_9606,N_8446,N_8578);
nand U9607 (N_9607,N_8333,N_8503);
nor U9608 (N_9608,N_8385,N_8887);
or U9609 (N_9609,N_8277,N_8104);
nor U9610 (N_9610,N_8299,N_8785);
xor U9611 (N_9611,N_8064,N_8143);
or U9612 (N_9612,N_8833,N_8506);
or U9613 (N_9613,N_8697,N_8452);
xnor U9614 (N_9614,N_8086,N_8659);
nand U9615 (N_9615,N_8444,N_8052);
or U9616 (N_9616,N_8463,N_8157);
nor U9617 (N_9617,N_8768,N_8974);
xnor U9618 (N_9618,N_8632,N_8598);
or U9619 (N_9619,N_8374,N_8993);
nor U9620 (N_9620,N_8712,N_8557);
or U9621 (N_9621,N_8125,N_8339);
or U9622 (N_9622,N_8203,N_8624);
xnor U9623 (N_9623,N_8718,N_8507);
and U9624 (N_9624,N_8113,N_8257);
and U9625 (N_9625,N_8983,N_8913);
nand U9626 (N_9626,N_8774,N_8725);
nand U9627 (N_9627,N_8838,N_8113);
nand U9628 (N_9628,N_8982,N_8436);
or U9629 (N_9629,N_8540,N_8150);
nand U9630 (N_9630,N_8070,N_8371);
nand U9631 (N_9631,N_8146,N_8124);
or U9632 (N_9632,N_8597,N_8497);
nor U9633 (N_9633,N_8988,N_8525);
and U9634 (N_9634,N_8234,N_8353);
xnor U9635 (N_9635,N_8790,N_8218);
nand U9636 (N_9636,N_8040,N_8041);
and U9637 (N_9637,N_8777,N_8772);
nor U9638 (N_9638,N_8464,N_8058);
nand U9639 (N_9639,N_8076,N_8975);
nor U9640 (N_9640,N_8732,N_8135);
xor U9641 (N_9641,N_8039,N_8290);
and U9642 (N_9642,N_8370,N_8798);
and U9643 (N_9643,N_8437,N_8473);
or U9644 (N_9644,N_8599,N_8401);
and U9645 (N_9645,N_8373,N_8334);
nand U9646 (N_9646,N_8560,N_8127);
or U9647 (N_9647,N_8702,N_8708);
or U9648 (N_9648,N_8030,N_8634);
nand U9649 (N_9649,N_8780,N_8169);
and U9650 (N_9650,N_8267,N_8498);
nand U9651 (N_9651,N_8706,N_8229);
and U9652 (N_9652,N_8841,N_8225);
nor U9653 (N_9653,N_8796,N_8227);
nand U9654 (N_9654,N_8379,N_8040);
and U9655 (N_9655,N_8385,N_8109);
or U9656 (N_9656,N_8529,N_8067);
xor U9657 (N_9657,N_8160,N_8202);
nor U9658 (N_9658,N_8062,N_8500);
xnor U9659 (N_9659,N_8556,N_8829);
nor U9660 (N_9660,N_8083,N_8486);
xor U9661 (N_9661,N_8580,N_8588);
and U9662 (N_9662,N_8840,N_8691);
and U9663 (N_9663,N_8615,N_8642);
nand U9664 (N_9664,N_8837,N_8669);
nand U9665 (N_9665,N_8750,N_8994);
or U9666 (N_9666,N_8565,N_8836);
xor U9667 (N_9667,N_8882,N_8729);
and U9668 (N_9668,N_8896,N_8543);
xor U9669 (N_9669,N_8886,N_8580);
nand U9670 (N_9670,N_8581,N_8193);
nor U9671 (N_9671,N_8294,N_8838);
xor U9672 (N_9672,N_8199,N_8475);
xnor U9673 (N_9673,N_8810,N_8569);
or U9674 (N_9674,N_8885,N_8834);
nand U9675 (N_9675,N_8875,N_8387);
nor U9676 (N_9676,N_8246,N_8289);
nand U9677 (N_9677,N_8278,N_8600);
and U9678 (N_9678,N_8686,N_8096);
nor U9679 (N_9679,N_8417,N_8261);
and U9680 (N_9680,N_8841,N_8603);
xnor U9681 (N_9681,N_8374,N_8846);
or U9682 (N_9682,N_8208,N_8566);
xnor U9683 (N_9683,N_8303,N_8429);
xor U9684 (N_9684,N_8695,N_8092);
or U9685 (N_9685,N_8240,N_8594);
or U9686 (N_9686,N_8018,N_8708);
nor U9687 (N_9687,N_8447,N_8793);
and U9688 (N_9688,N_8423,N_8765);
and U9689 (N_9689,N_8875,N_8596);
or U9690 (N_9690,N_8545,N_8210);
and U9691 (N_9691,N_8780,N_8516);
and U9692 (N_9692,N_8046,N_8042);
and U9693 (N_9693,N_8314,N_8217);
xnor U9694 (N_9694,N_8746,N_8432);
nand U9695 (N_9695,N_8079,N_8058);
and U9696 (N_9696,N_8963,N_8001);
nor U9697 (N_9697,N_8503,N_8225);
and U9698 (N_9698,N_8116,N_8284);
nor U9699 (N_9699,N_8639,N_8709);
xor U9700 (N_9700,N_8186,N_8395);
or U9701 (N_9701,N_8340,N_8596);
and U9702 (N_9702,N_8389,N_8406);
or U9703 (N_9703,N_8477,N_8040);
nor U9704 (N_9704,N_8524,N_8718);
nor U9705 (N_9705,N_8749,N_8048);
nand U9706 (N_9706,N_8021,N_8123);
nand U9707 (N_9707,N_8426,N_8417);
or U9708 (N_9708,N_8342,N_8767);
nand U9709 (N_9709,N_8939,N_8006);
and U9710 (N_9710,N_8677,N_8002);
nand U9711 (N_9711,N_8784,N_8605);
or U9712 (N_9712,N_8793,N_8951);
or U9713 (N_9713,N_8258,N_8568);
xnor U9714 (N_9714,N_8345,N_8673);
or U9715 (N_9715,N_8100,N_8850);
xnor U9716 (N_9716,N_8215,N_8726);
or U9717 (N_9717,N_8004,N_8770);
nor U9718 (N_9718,N_8061,N_8580);
nor U9719 (N_9719,N_8871,N_8722);
nand U9720 (N_9720,N_8240,N_8601);
nand U9721 (N_9721,N_8187,N_8258);
nor U9722 (N_9722,N_8623,N_8663);
xor U9723 (N_9723,N_8396,N_8299);
nor U9724 (N_9724,N_8656,N_8463);
nor U9725 (N_9725,N_8075,N_8466);
xor U9726 (N_9726,N_8367,N_8681);
nand U9727 (N_9727,N_8547,N_8112);
nor U9728 (N_9728,N_8766,N_8435);
nand U9729 (N_9729,N_8647,N_8276);
xor U9730 (N_9730,N_8760,N_8641);
or U9731 (N_9731,N_8787,N_8147);
xor U9732 (N_9732,N_8342,N_8291);
nor U9733 (N_9733,N_8128,N_8962);
nand U9734 (N_9734,N_8926,N_8150);
xnor U9735 (N_9735,N_8988,N_8771);
nand U9736 (N_9736,N_8460,N_8004);
and U9737 (N_9737,N_8560,N_8461);
nand U9738 (N_9738,N_8371,N_8910);
xnor U9739 (N_9739,N_8257,N_8097);
nand U9740 (N_9740,N_8456,N_8743);
nand U9741 (N_9741,N_8000,N_8253);
and U9742 (N_9742,N_8088,N_8506);
xnor U9743 (N_9743,N_8668,N_8585);
nor U9744 (N_9744,N_8988,N_8785);
or U9745 (N_9745,N_8656,N_8180);
xor U9746 (N_9746,N_8569,N_8775);
xnor U9747 (N_9747,N_8075,N_8235);
nor U9748 (N_9748,N_8123,N_8669);
xor U9749 (N_9749,N_8171,N_8549);
xor U9750 (N_9750,N_8308,N_8855);
or U9751 (N_9751,N_8457,N_8963);
xor U9752 (N_9752,N_8076,N_8550);
nor U9753 (N_9753,N_8195,N_8476);
nand U9754 (N_9754,N_8345,N_8957);
and U9755 (N_9755,N_8968,N_8555);
and U9756 (N_9756,N_8821,N_8949);
xor U9757 (N_9757,N_8250,N_8189);
and U9758 (N_9758,N_8551,N_8975);
xor U9759 (N_9759,N_8969,N_8250);
xor U9760 (N_9760,N_8451,N_8342);
nor U9761 (N_9761,N_8931,N_8780);
nand U9762 (N_9762,N_8091,N_8002);
or U9763 (N_9763,N_8511,N_8215);
or U9764 (N_9764,N_8706,N_8994);
xnor U9765 (N_9765,N_8202,N_8292);
nor U9766 (N_9766,N_8756,N_8539);
nand U9767 (N_9767,N_8615,N_8669);
nand U9768 (N_9768,N_8691,N_8927);
nor U9769 (N_9769,N_8912,N_8267);
or U9770 (N_9770,N_8229,N_8971);
or U9771 (N_9771,N_8240,N_8083);
nand U9772 (N_9772,N_8676,N_8528);
xnor U9773 (N_9773,N_8742,N_8131);
nor U9774 (N_9774,N_8454,N_8486);
and U9775 (N_9775,N_8636,N_8574);
and U9776 (N_9776,N_8947,N_8219);
nand U9777 (N_9777,N_8598,N_8313);
xor U9778 (N_9778,N_8536,N_8768);
and U9779 (N_9779,N_8818,N_8853);
nor U9780 (N_9780,N_8630,N_8007);
nand U9781 (N_9781,N_8273,N_8964);
and U9782 (N_9782,N_8023,N_8204);
or U9783 (N_9783,N_8168,N_8018);
nor U9784 (N_9784,N_8563,N_8552);
and U9785 (N_9785,N_8258,N_8260);
or U9786 (N_9786,N_8988,N_8390);
or U9787 (N_9787,N_8080,N_8474);
or U9788 (N_9788,N_8519,N_8778);
nand U9789 (N_9789,N_8628,N_8310);
xnor U9790 (N_9790,N_8765,N_8197);
nor U9791 (N_9791,N_8429,N_8332);
xnor U9792 (N_9792,N_8298,N_8273);
and U9793 (N_9793,N_8445,N_8045);
nor U9794 (N_9794,N_8619,N_8992);
or U9795 (N_9795,N_8246,N_8916);
xnor U9796 (N_9796,N_8575,N_8163);
xnor U9797 (N_9797,N_8732,N_8808);
nor U9798 (N_9798,N_8676,N_8421);
or U9799 (N_9799,N_8631,N_8300);
xor U9800 (N_9800,N_8533,N_8258);
nand U9801 (N_9801,N_8486,N_8837);
xnor U9802 (N_9802,N_8819,N_8961);
nor U9803 (N_9803,N_8344,N_8650);
xor U9804 (N_9804,N_8791,N_8345);
xor U9805 (N_9805,N_8664,N_8742);
nor U9806 (N_9806,N_8868,N_8172);
and U9807 (N_9807,N_8717,N_8977);
and U9808 (N_9808,N_8647,N_8928);
or U9809 (N_9809,N_8553,N_8679);
and U9810 (N_9810,N_8721,N_8099);
nand U9811 (N_9811,N_8643,N_8437);
or U9812 (N_9812,N_8900,N_8148);
nor U9813 (N_9813,N_8638,N_8689);
xor U9814 (N_9814,N_8184,N_8350);
xnor U9815 (N_9815,N_8625,N_8166);
nor U9816 (N_9816,N_8428,N_8869);
xnor U9817 (N_9817,N_8429,N_8040);
or U9818 (N_9818,N_8548,N_8651);
xnor U9819 (N_9819,N_8835,N_8051);
xor U9820 (N_9820,N_8266,N_8628);
and U9821 (N_9821,N_8497,N_8056);
or U9822 (N_9822,N_8281,N_8577);
xnor U9823 (N_9823,N_8155,N_8527);
xnor U9824 (N_9824,N_8293,N_8313);
nand U9825 (N_9825,N_8643,N_8790);
nor U9826 (N_9826,N_8423,N_8290);
xnor U9827 (N_9827,N_8871,N_8234);
nor U9828 (N_9828,N_8861,N_8881);
and U9829 (N_9829,N_8580,N_8157);
or U9830 (N_9830,N_8151,N_8385);
nor U9831 (N_9831,N_8819,N_8908);
or U9832 (N_9832,N_8487,N_8693);
xor U9833 (N_9833,N_8160,N_8110);
and U9834 (N_9834,N_8314,N_8625);
and U9835 (N_9835,N_8318,N_8125);
xor U9836 (N_9836,N_8262,N_8577);
xor U9837 (N_9837,N_8426,N_8909);
nor U9838 (N_9838,N_8812,N_8970);
xor U9839 (N_9839,N_8954,N_8633);
xnor U9840 (N_9840,N_8132,N_8280);
nand U9841 (N_9841,N_8357,N_8106);
or U9842 (N_9842,N_8819,N_8923);
nor U9843 (N_9843,N_8365,N_8753);
or U9844 (N_9844,N_8579,N_8013);
nand U9845 (N_9845,N_8733,N_8529);
xor U9846 (N_9846,N_8041,N_8423);
or U9847 (N_9847,N_8215,N_8304);
nor U9848 (N_9848,N_8066,N_8212);
nor U9849 (N_9849,N_8689,N_8289);
and U9850 (N_9850,N_8348,N_8101);
nor U9851 (N_9851,N_8604,N_8428);
and U9852 (N_9852,N_8501,N_8476);
and U9853 (N_9853,N_8360,N_8097);
nor U9854 (N_9854,N_8908,N_8460);
and U9855 (N_9855,N_8412,N_8450);
xnor U9856 (N_9856,N_8077,N_8934);
or U9857 (N_9857,N_8730,N_8694);
nand U9858 (N_9858,N_8299,N_8607);
and U9859 (N_9859,N_8120,N_8296);
xor U9860 (N_9860,N_8233,N_8816);
nor U9861 (N_9861,N_8441,N_8453);
nor U9862 (N_9862,N_8201,N_8381);
or U9863 (N_9863,N_8422,N_8744);
nor U9864 (N_9864,N_8222,N_8665);
nor U9865 (N_9865,N_8907,N_8264);
and U9866 (N_9866,N_8292,N_8935);
nor U9867 (N_9867,N_8111,N_8282);
or U9868 (N_9868,N_8867,N_8579);
or U9869 (N_9869,N_8725,N_8772);
nor U9870 (N_9870,N_8897,N_8032);
xor U9871 (N_9871,N_8403,N_8057);
nor U9872 (N_9872,N_8679,N_8239);
nor U9873 (N_9873,N_8891,N_8929);
nor U9874 (N_9874,N_8115,N_8970);
nand U9875 (N_9875,N_8913,N_8143);
xnor U9876 (N_9876,N_8356,N_8897);
xnor U9877 (N_9877,N_8567,N_8832);
nor U9878 (N_9878,N_8596,N_8762);
xor U9879 (N_9879,N_8578,N_8348);
nand U9880 (N_9880,N_8664,N_8855);
nor U9881 (N_9881,N_8012,N_8877);
and U9882 (N_9882,N_8013,N_8726);
nor U9883 (N_9883,N_8494,N_8328);
xnor U9884 (N_9884,N_8629,N_8966);
xor U9885 (N_9885,N_8841,N_8449);
nand U9886 (N_9886,N_8904,N_8341);
nand U9887 (N_9887,N_8360,N_8393);
and U9888 (N_9888,N_8312,N_8377);
nand U9889 (N_9889,N_8861,N_8747);
and U9890 (N_9890,N_8096,N_8385);
or U9891 (N_9891,N_8982,N_8655);
xor U9892 (N_9892,N_8873,N_8475);
nand U9893 (N_9893,N_8772,N_8824);
or U9894 (N_9894,N_8066,N_8819);
or U9895 (N_9895,N_8104,N_8711);
xor U9896 (N_9896,N_8037,N_8310);
nand U9897 (N_9897,N_8376,N_8239);
or U9898 (N_9898,N_8163,N_8768);
or U9899 (N_9899,N_8111,N_8070);
nand U9900 (N_9900,N_8604,N_8653);
xnor U9901 (N_9901,N_8507,N_8906);
nor U9902 (N_9902,N_8142,N_8612);
and U9903 (N_9903,N_8760,N_8749);
nor U9904 (N_9904,N_8335,N_8627);
or U9905 (N_9905,N_8353,N_8671);
or U9906 (N_9906,N_8862,N_8050);
xnor U9907 (N_9907,N_8354,N_8464);
xor U9908 (N_9908,N_8563,N_8786);
and U9909 (N_9909,N_8269,N_8155);
nand U9910 (N_9910,N_8655,N_8851);
or U9911 (N_9911,N_8975,N_8592);
or U9912 (N_9912,N_8769,N_8327);
xnor U9913 (N_9913,N_8595,N_8743);
nor U9914 (N_9914,N_8991,N_8332);
xnor U9915 (N_9915,N_8670,N_8347);
and U9916 (N_9916,N_8431,N_8872);
and U9917 (N_9917,N_8703,N_8908);
xor U9918 (N_9918,N_8389,N_8515);
nand U9919 (N_9919,N_8456,N_8274);
nand U9920 (N_9920,N_8688,N_8887);
or U9921 (N_9921,N_8657,N_8304);
or U9922 (N_9922,N_8671,N_8189);
or U9923 (N_9923,N_8301,N_8705);
nor U9924 (N_9924,N_8153,N_8490);
nand U9925 (N_9925,N_8501,N_8745);
and U9926 (N_9926,N_8013,N_8650);
xnor U9927 (N_9927,N_8430,N_8638);
or U9928 (N_9928,N_8561,N_8006);
nand U9929 (N_9929,N_8290,N_8168);
nand U9930 (N_9930,N_8305,N_8798);
or U9931 (N_9931,N_8712,N_8933);
nand U9932 (N_9932,N_8088,N_8585);
nor U9933 (N_9933,N_8282,N_8703);
and U9934 (N_9934,N_8191,N_8331);
or U9935 (N_9935,N_8237,N_8624);
nor U9936 (N_9936,N_8799,N_8443);
nor U9937 (N_9937,N_8029,N_8208);
nor U9938 (N_9938,N_8324,N_8780);
nand U9939 (N_9939,N_8081,N_8518);
or U9940 (N_9940,N_8073,N_8784);
or U9941 (N_9941,N_8915,N_8030);
or U9942 (N_9942,N_8713,N_8192);
or U9943 (N_9943,N_8339,N_8611);
nor U9944 (N_9944,N_8884,N_8716);
xnor U9945 (N_9945,N_8281,N_8979);
xor U9946 (N_9946,N_8406,N_8552);
or U9947 (N_9947,N_8070,N_8546);
nand U9948 (N_9948,N_8601,N_8620);
and U9949 (N_9949,N_8862,N_8489);
nand U9950 (N_9950,N_8144,N_8582);
nor U9951 (N_9951,N_8434,N_8463);
nand U9952 (N_9952,N_8033,N_8952);
and U9953 (N_9953,N_8050,N_8940);
and U9954 (N_9954,N_8398,N_8876);
nor U9955 (N_9955,N_8309,N_8565);
and U9956 (N_9956,N_8472,N_8351);
or U9957 (N_9957,N_8000,N_8299);
nand U9958 (N_9958,N_8842,N_8433);
nor U9959 (N_9959,N_8414,N_8572);
nor U9960 (N_9960,N_8296,N_8475);
or U9961 (N_9961,N_8210,N_8193);
and U9962 (N_9962,N_8251,N_8167);
and U9963 (N_9963,N_8815,N_8260);
nand U9964 (N_9964,N_8396,N_8695);
nor U9965 (N_9965,N_8614,N_8062);
xor U9966 (N_9966,N_8930,N_8026);
xnor U9967 (N_9967,N_8142,N_8439);
or U9968 (N_9968,N_8862,N_8791);
or U9969 (N_9969,N_8629,N_8142);
nand U9970 (N_9970,N_8609,N_8543);
or U9971 (N_9971,N_8996,N_8831);
nor U9972 (N_9972,N_8294,N_8765);
nor U9973 (N_9973,N_8502,N_8807);
xnor U9974 (N_9974,N_8113,N_8242);
nand U9975 (N_9975,N_8382,N_8452);
xor U9976 (N_9976,N_8263,N_8421);
and U9977 (N_9977,N_8892,N_8425);
nand U9978 (N_9978,N_8710,N_8705);
or U9979 (N_9979,N_8660,N_8750);
xnor U9980 (N_9980,N_8289,N_8742);
nand U9981 (N_9981,N_8227,N_8806);
or U9982 (N_9982,N_8118,N_8164);
and U9983 (N_9983,N_8814,N_8419);
and U9984 (N_9984,N_8035,N_8721);
or U9985 (N_9985,N_8438,N_8478);
nor U9986 (N_9986,N_8781,N_8795);
and U9987 (N_9987,N_8628,N_8475);
xor U9988 (N_9988,N_8689,N_8727);
nand U9989 (N_9989,N_8283,N_8997);
nor U9990 (N_9990,N_8456,N_8620);
xor U9991 (N_9991,N_8117,N_8876);
xnor U9992 (N_9992,N_8363,N_8699);
xnor U9993 (N_9993,N_8645,N_8873);
xor U9994 (N_9994,N_8624,N_8311);
or U9995 (N_9995,N_8498,N_8592);
nor U9996 (N_9996,N_8431,N_8594);
and U9997 (N_9997,N_8135,N_8775);
nor U9998 (N_9998,N_8188,N_8454);
or U9999 (N_9999,N_8779,N_8468);
xor U10000 (N_10000,N_9734,N_9560);
nand U10001 (N_10001,N_9995,N_9593);
and U10002 (N_10002,N_9456,N_9379);
and U10003 (N_10003,N_9415,N_9159);
nand U10004 (N_10004,N_9578,N_9248);
xor U10005 (N_10005,N_9189,N_9943);
or U10006 (N_10006,N_9769,N_9154);
and U10007 (N_10007,N_9236,N_9253);
or U10008 (N_10008,N_9360,N_9685);
nand U10009 (N_10009,N_9766,N_9941);
and U10010 (N_10010,N_9750,N_9588);
nand U10011 (N_10011,N_9779,N_9031);
and U10012 (N_10012,N_9243,N_9126);
nand U10013 (N_10013,N_9891,N_9717);
nand U10014 (N_10014,N_9896,N_9876);
nand U10015 (N_10015,N_9352,N_9382);
and U10016 (N_10016,N_9036,N_9858);
and U10017 (N_10017,N_9881,N_9129);
nand U10018 (N_10018,N_9116,N_9540);
nor U10019 (N_10019,N_9491,N_9216);
nand U10020 (N_10020,N_9393,N_9019);
and U10021 (N_10021,N_9577,N_9017);
xor U10022 (N_10022,N_9230,N_9339);
nand U10023 (N_10023,N_9543,N_9933);
and U10024 (N_10024,N_9186,N_9797);
xor U10025 (N_10025,N_9217,N_9956);
nor U10026 (N_10026,N_9403,N_9887);
xor U10027 (N_10027,N_9961,N_9803);
or U10028 (N_10028,N_9653,N_9760);
and U10029 (N_10029,N_9369,N_9520);
xnor U10030 (N_10030,N_9582,N_9408);
and U10031 (N_10031,N_9747,N_9917);
or U10032 (N_10032,N_9002,N_9982);
or U10033 (N_10033,N_9203,N_9938);
and U10034 (N_10034,N_9093,N_9185);
nand U10035 (N_10035,N_9856,N_9892);
or U10036 (N_10036,N_9077,N_9525);
or U10037 (N_10037,N_9380,N_9849);
nor U10038 (N_10038,N_9325,N_9712);
nand U10039 (N_10039,N_9549,N_9206);
and U10040 (N_10040,N_9710,N_9903);
or U10041 (N_10041,N_9402,N_9953);
nand U10042 (N_10042,N_9249,N_9628);
xnor U10043 (N_10043,N_9460,N_9333);
or U10044 (N_10044,N_9478,N_9099);
xnor U10045 (N_10045,N_9764,N_9058);
or U10046 (N_10046,N_9562,N_9187);
nor U10047 (N_10047,N_9356,N_9962);
xnor U10048 (N_10048,N_9072,N_9798);
nand U10049 (N_10049,N_9361,N_9479);
nor U10050 (N_10050,N_9032,N_9544);
nor U10051 (N_10051,N_9513,N_9056);
xnor U10052 (N_10052,N_9191,N_9699);
nor U10053 (N_10053,N_9272,N_9518);
nand U10054 (N_10054,N_9314,N_9390);
nand U10055 (N_10055,N_9472,N_9133);
and U10056 (N_10056,N_9844,N_9312);
nand U10057 (N_10057,N_9346,N_9698);
and U10058 (N_10058,N_9771,N_9895);
or U10059 (N_10059,N_9992,N_9709);
nand U10060 (N_10060,N_9886,N_9322);
or U10061 (N_10061,N_9649,N_9737);
nand U10062 (N_10062,N_9494,N_9413);
and U10063 (N_10063,N_9125,N_9984);
xor U10064 (N_10064,N_9008,N_9433);
or U10065 (N_10065,N_9111,N_9283);
or U10066 (N_10066,N_9527,N_9502);
nor U10067 (N_10067,N_9662,N_9626);
xor U10068 (N_10068,N_9024,N_9557);
or U10069 (N_10069,N_9137,N_9752);
nand U10070 (N_10070,N_9865,N_9607);
or U10071 (N_10071,N_9081,N_9120);
and U10072 (N_10072,N_9336,N_9681);
nand U10073 (N_10073,N_9400,N_9815);
xnor U10074 (N_10074,N_9439,N_9783);
nor U10075 (N_10075,N_9556,N_9347);
and U10076 (N_10076,N_9633,N_9666);
and U10077 (N_10077,N_9700,N_9595);
or U10078 (N_10078,N_9065,N_9515);
or U10079 (N_10079,N_9138,N_9384);
or U10080 (N_10080,N_9637,N_9220);
or U10081 (N_10081,N_9447,N_9660);
nor U10082 (N_10082,N_9970,N_9250);
nand U10083 (N_10083,N_9761,N_9714);
xnor U10084 (N_10084,N_9343,N_9028);
xnor U10085 (N_10085,N_9535,N_9173);
nor U10086 (N_10086,N_9772,N_9328);
or U10087 (N_10087,N_9365,N_9062);
xor U10088 (N_10088,N_9565,N_9959);
nand U10089 (N_10089,N_9857,N_9353);
or U10090 (N_10090,N_9840,N_9027);
or U10091 (N_10091,N_9420,N_9350);
or U10092 (N_10092,N_9949,N_9241);
and U10093 (N_10093,N_9988,N_9642);
and U10094 (N_10094,N_9348,N_9590);
xnor U10095 (N_10095,N_9997,N_9960);
or U10096 (N_10096,N_9923,N_9668);
or U10097 (N_10097,N_9921,N_9966);
nor U10098 (N_10098,N_9499,N_9102);
xor U10099 (N_10099,N_9483,N_9894);
xnor U10100 (N_10100,N_9276,N_9287);
nor U10101 (N_10101,N_9204,N_9680);
nor U10102 (N_10102,N_9300,N_9768);
nand U10103 (N_10103,N_9945,N_9324);
nand U10104 (N_10104,N_9304,N_9257);
nor U10105 (N_10105,N_9405,N_9208);
xor U10106 (N_10106,N_9273,N_9452);
nor U10107 (N_10107,N_9808,N_9545);
nand U10108 (N_10108,N_9449,N_9197);
and U10109 (N_10109,N_9282,N_9237);
or U10110 (N_10110,N_9068,N_9155);
xnor U10111 (N_10111,N_9824,N_9222);
nand U10112 (N_10112,N_9316,N_9880);
nor U10113 (N_10113,N_9848,N_9615);
nor U10114 (N_10114,N_9829,N_9758);
nand U10115 (N_10115,N_9147,N_9057);
nor U10116 (N_10116,N_9647,N_9519);
or U10117 (N_10117,N_9823,N_9799);
nand U10118 (N_10118,N_9014,N_9931);
or U10119 (N_10119,N_9684,N_9211);
and U10120 (N_10120,N_9210,N_9445);
nand U10121 (N_10121,N_9127,N_9431);
or U10122 (N_10122,N_9916,N_9158);
nor U10123 (N_10123,N_9184,N_9354);
nand U10124 (N_10124,N_9115,N_9335);
xnor U10125 (N_10125,N_9994,N_9381);
nand U10126 (N_10126,N_9996,N_9410);
nor U10127 (N_10127,N_9188,N_9991);
or U10128 (N_10128,N_9288,N_9142);
nand U10129 (N_10129,N_9897,N_9985);
xor U10130 (N_10130,N_9073,N_9207);
xor U10131 (N_10131,N_9118,N_9367);
nand U10132 (N_10132,N_9134,N_9429);
xnor U10133 (N_10133,N_9476,N_9161);
and U10134 (N_10134,N_9167,N_9832);
nor U10135 (N_10135,N_9745,N_9725);
nor U10136 (N_10136,N_9192,N_9157);
nand U10137 (N_10137,N_9374,N_9526);
nand U10138 (N_10138,N_9516,N_9029);
or U10139 (N_10139,N_9845,N_9821);
nor U10140 (N_10140,N_9226,N_9292);
xnor U10141 (N_10141,N_9162,N_9837);
nand U10142 (N_10142,N_9890,N_9968);
nor U10143 (N_10143,N_9366,N_9268);
xor U10144 (N_10144,N_9568,N_9487);
nor U10145 (N_10145,N_9025,N_9691);
or U10146 (N_10146,N_9980,N_9804);
or U10147 (N_10147,N_9201,N_9874);
xnor U10148 (N_10148,N_9198,N_9655);
nand U10149 (N_10149,N_9735,N_9561);
nor U10150 (N_10150,N_9807,N_9825);
nand U10151 (N_10151,N_9475,N_9852);
nor U10152 (N_10152,N_9117,N_9317);
nor U10153 (N_10153,N_9862,N_9101);
or U10154 (N_10154,N_9703,N_9645);
xor U10155 (N_10155,N_9442,N_9489);
or U10156 (N_10156,N_9052,N_9656);
nand U10157 (N_10157,N_9376,N_9464);
and U10158 (N_10158,N_9567,N_9508);
and U10159 (N_10159,N_9199,N_9688);
nand U10160 (N_10160,N_9939,N_9501);
nor U10161 (N_10161,N_9496,N_9524);
nand U10162 (N_10162,N_9898,N_9753);
and U10163 (N_10163,N_9785,N_9235);
nor U10164 (N_10164,N_9830,N_9040);
nor U10165 (N_10165,N_9541,N_9539);
or U10166 (N_10166,N_9678,N_9861);
nor U10167 (N_10167,N_9884,N_9121);
xnor U10168 (N_10168,N_9667,N_9835);
nand U10169 (N_10169,N_9926,N_9602);
xnor U10170 (N_10170,N_9109,N_9190);
and U10171 (N_10171,N_9462,N_9048);
or U10172 (N_10172,N_9802,N_9981);
xnor U10173 (N_10173,N_9695,N_9875);
nor U10174 (N_10174,N_9964,N_9811);
nor U10175 (N_10175,N_9289,N_9906);
xor U10176 (N_10176,N_9486,N_9899);
or U10177 (N_10177,N_9076,N_9603);
or U10178 (N_10178,N_9227,N_9573);
or U10179 (N_10179,N_9935,N_9426);
nand U10180 (N_10180,N_9416,N_9912);
and U10181 (N_10181,N_9853,N_9090);
nor U10182 (N_10182,N_9748,N_9720);
xor U10183 (N_10183,N_9687,N_9529);
or U10184 (N_10184,N_9428,N_9739);
and U10185 (N_10185,N_9087,N_9046);
nand U10186 (N_10186,N_9746,N_9682);
xor U10187 (N_10187,N_9389,N_9570);
nand U10188 (N_10188,N_9311,N_9869);
and U10189 (N_10189,N_9728,N_9003);
nor U10190 (N_10190,N_9796,N_9706);
nor U10191 (N_10191,N_9094,N_9993);
and U10192 (N_10192,N_9587,N_9601);
nor U10193 (N_10193,N_9910,N_9175);
and U10194 (N_10194,N_9592,N_9630);
nand U10195 (N_10195,N_9636,N_9122);
or U10196 (N_10196,N_9605,N_9377);
and U10197 (N_10197,N_9900,N_9221);
nor U10198 (N_10198,N_9332,N_9233);
nand U10199 (N_10199,N_9329,N_9533);
nand U10200 (N_10200,N_9051,N_9517);
nand U10201 (N_10201,N_9523,N_9394);
or U10202 (N_10202,N_9107,N_9885);
xor U10203 (N_10203,N_9432,N_9690);
xnor U10204 (N_10204,N_9412,N_9275);
xor U10205 (N_10205,N_9528,N_9757);
nor U10206 (N_10206,N_9911,N_9741);
xnor U10207 (N_10207,N_9218,N_9139);
xor U10208 (N_10208,N_9124,N_9296);
nor U10209 (N_10209,N_9291,N_9414);
nor U10210 (N_10210,N_9879,N_9174);
and U10211 (N_10211,N_9045,N_9385);
nand U10212 (N_10212,N_9473,N_9418);
nor U10213 (N_10213,N_9098,N_9397);
xor U10214 (N_10214,N_9512,N_9484);
and U10215 (N_10215,N_9537,N_9256);
or U10216 (N_10216,N_9244,N_9168);
nand U10217 (N_10217,N_9708,N_9437);
and U10218 (N_10218,N_9041,N_9671);
and U10219 (N_10219,N_9454,N_9215);
xor U10220 (N_10220,N_9140,N_9676);
or U10221 (N_10221,N_9063,N_9532);
and U10222 (N_10222,N_9877,N_9049);
xor U10223 (N_10223,N_9702,N_9580);
nor U10224 (N_10224,N_9707,N_9552);
nand U10225 (N_10225,N_9178,N_9306);
xor U10226 (N_10226,N_9463,N_9831);
xor U10227 (N_10227,N_9599,N_9337);
or U10228 (N_10228,N_9301,N_9809);
or U10229 (N_10229,N_9182,N_9978);
or U10230 (N_10230,N_9144,N_9621);
nor U10231 (N_10231,N_9088,N_9310);
and U10232 (N_10232,N_9242,N_9972);
and U10233 (N_10233,N_9606,N_9011);
and U10234 (N_10234,N_9100,N_9971);
and U10235 (N_10235,N_9751,N_9225);
nor U10236 (N_10236,N_9983,N_9097);
or U10237 (N_10237,N_9617,N_9375);
and U10238 (N_10238,N_9266,N_9181);
and U10239 (N_10239,N_9631,N_9451);
nor U10240 (N_10240,N_9183,N_9500);
and U10241 (N_10241,N_9547,N_9979);
xnor U10242 (N_10242,N_9318,N_9816);
and U10243 (N_10243,N_9836,N_9723);
and U10244 (N_10244,N_9789,N_9929);
and U10245 (N_10245,N_9818,N_9534);
nor U10246 (N_10246,N_9672,N_9870);
nand U10247 (N_10247,N_9294,N_9860);
or U10248 (N_10248,N_9326,N_9531);
and U10249 (N_10249,N_9998,N_9850);
nor U10250 (N_10250,N_9349,N_9736);
or U10251 (N_10251,N_9613,N_9510);
and U10252 (N_10252,N_9434,N_9039);
nor U10253 (N_10253,N_9705,N_9654);
and U10254 (N_10254,N_9932,N_9006);
or U10255 (N_10255,N_9240,N_9915);
xor U10256 (N_10256,N_9872,N_9990);
and U10257 (N_10257,N_9293,N_9214);
nor U10258 (N_10258,N_9364,N_9265);
and U10259 (N_10259,N_9370,N_9004);
xor U10260 (N_10260,N_9387,N_9503);
xor U10261 (N_10261,N_9080,N_9612);
or U10262 (N_10262,N_9228,N_9563);
nor U10263 (N_10263,N_9308,N_9866);
and U10264 (N_10264,N_9947,N_9195);
nand U10265 (N_10265,N_9999,N_9893);
and U10266 (N_10266,N_9194,N_9648);
xor U10267 (N_10267,N_9149,N_9696);
or U10268 (N_10268,N_9148,N_9022);
or U10269 (N_10269,N_9135,N_9609);
xor U10270 (N_10270,N_9812,N_9341);
nand U10271 (N_10271,N_9948,N_9677);
and U10272 (N_10272,N_9665,N_9247);
nand U10273 (N_10273,N_9784,N_9430);
nor U10274 (N_10274,N_9686,N_9363);
nor U10275 (N_10275,N_9571,N_9061);
or U10276 (N_10276,N_9123,N_9722);
nand U10277 (N_10277,N_9007,N_9095);
and U10278 (N_10278,N_9566,N_9596);
nor U10279 (N_10279,N_9298,N_9112);
xnor U10280 (N_10280,N_9373,N_9509);
nor U10281 (N_10281,N_9559,N_9659);
or U10282 (N_10282,N_9105,N_9200);
nand U10283 (N_10283,N_9744,N_9608);
xnor U10284 (N_10284,N_9594,N_9160);
nand U10285 (N_10285,N_9574,N_9641);
nand U10286 (N_10286,N_9152,N_9600);
and U10287 (N_10287,N_9251,N_9584);
nand U10288 (N_10288,N_9987,N_9012);
and U10289 (N_10289,N_9542,N_9827);
and U10290 (N_10290,N_9833,N_9918);
nor U10291 (N_10291,N_9224,N_9407);
xnor U10292 (N_10292,N_9842,N_9650);
nand U10293 (N_10293,N_9424,N_9975);
and U10294 (N_10294,N_9013,N_9822);
nand U10295 (N_10295,N_9330,N_9794);
nand U10296 (N_10296,N_9787,N_9342);
xnor U10297 (N_10297,N_9765,N_9793);
and U10298 (N_10298,N_9719,N_9309);
nor U10299 (N_10299,N_9651,N_9422);
and U10300 (N_10300,N_9358,N_9092);
or U10301 (N_10301,N_9740,N_9023);
or U10302 (N_10302,N_9619,N_9132);
nand U10303 (N_10303,N_9942,N_9806);
nand U10304 (N_10304,N_9924,N_9963);
nand U10305 (N_10305,N_9082,N_9558);
and U10306 (N_10306,N_9481,N_9927);
xnor U10307 (N_10307,N_9469,N_9466);
and U10308 (N_10308,N_9172,N_9009);
or U10309 (N_10309,N_9277,N_9461);
and U10310 (N_10310,N_9435,N_9792);
nand U10311 (N_10311,N_9675,N_9863);
nor U10312 (N_10312,N_9086,N_9320);
nor U10313 (N_10313,N_9713,N_9219);
nand U10314 (N_10314,N_9327,N_9589);
xnor U10315 (N_10315,N_9554,N_9069);
and U10316 (N_10316,N_9193,N_9604);
or U10317 (N_10317,N_9391,N_9493);
and U10318 (N_10318,N_9245,N_9733);
nor U10319 (N_10319,N_9085,N_9334);
nor U10320 (N_10320,N_9362,N_9773);
nor U10321 (N_10321,N_9694,N_9670);
or U10322 (N_10322,N_9169,N_9357);
nor U10323 (N_10323,N_9331,N_9954);
and U10324 (N_10324,N_9726,N_9967);
nor U10325 (N_10325,N_9059,N_9839);
xnor U10326 (N_10326,N_9620,N_9550);
nor U10327 (N_10327,N_9388,N_9922);
nand U10328 (N_10328,N_9313,N_9171);
nand U10329 (N_10329,N_9826,N_9634);
nand U10330 (N_10330,N_9583,N_9021);
nor U10331 (N_10331,N_9438,N_9854);
or U10332 (N_10332,N_9020,N_9141);
or U10333 (N_10333,N_9598,N_9864);
or U10334 (N_10334,N_9788,N_9297);
xor U10335 (N_10335,N_9444,N_9944);
nor U10336 (N_10336,N_9450,N_9396);
xor U10337 (N_10337,N_9791,N_9411);
and U10338 (N_10338,N_9506,N_9170);
or U10339 (N_10339,N_9718,N_9474);
or U10340 (N_10340,N_9538,N_9303);
or U10341 (N_10341,N_9946,N_9646);
xor U10342 (N_10342,N_9103,N_9627);
xor U10343 (N_10343,N_9759,N_9958);
and U10344 (N_10344,N_9813,N_9934);
nor U10345 (N_10345,N_9778,N_9905);
or U10346 (N_10346,N_9477,N_9459);
nand U10347 (N_10347,N_9805,N_9401);
xor U10348 (N_10348,N_9252,N_9883);
nand U10349 (N_10349,N_9673,N_9406);
and U10350 (N_10350,N_9371,N_9427);
or U10351 (N_10351,N_9205,N_9913);
nand U10352 (N_10352,N_9624,N_9457);
or U10353 (N_10353,N_9258,N_9470);
nor U10354 (N_10354,N_9034,N_9530);
nand U10355 (N_10355,N_9471,N_9255);
nand U10356 (N_10356,N_9576,N_9820);
or U10357 (N_10357,N_9498,N_9035);
nand U10358 (N_10358,N_9930,N_9037);
xor U10359 (N_10359,N_9777,N_9693);
and U10360 (N_10360,N_9492,N_9986);
xnor U10361 (N_10361,N_9841,N_9867);
nand U10362 (N_10362,N_9398,N_9421);
xnor U10363 (N_10363,N_9553,N_9066);
nor U10364 (N_10364,N_9404,N_9919);
nor U10365 (N_10365,N_9351,N_9392);
and U10366 (N_10366,N_9033,N_9482);
xor U10367 (N_10367,N_9724,N_9060);
and U10368 (N_10368,N_9378,N_9131);
nand U10369 (N_10369,N_9467,N_9321);
nand U10370 (N_10370,N_9128,N_9239);
nor U10371 (N_10371,N_9639,N_9212);
and U10372 (N_10372,N_9585,N_9026);
or U10373 (N_10373,N_9231,N_9974);
xnor U10374 (N_10374,N_9743,N_9071);
nand U10375 (N_10375,N_9089,N_9260);
nor U10376 (N_10376,N_9368,N_9622);
nor U10377 (N_10377,N_9704,N_9762);
nand U10378 (N_10378,N_9838,N_9106);
and U10379 (N_10379,N_9078,N_9755);
and U10380 (N_10380,N_9868,N_9043);
nor U10381 (N_10381,N_9232,N_9164);
nor U10382 (N_10382,N_9267,N_9495);
or U10383 (N_10383,N_9146,N_9180);
nand U10384 (N_10384,N_9281,N_9610);
and U10385 (N_10385,N_9950,N_9638);
and U10386 (N_10386,N_9716,N_9914);
nor U10387 (N_10387,N_9074,N_9871);
and U10388 (N_10388,N_9730,N_9928);
and U10389 (N_10389,N_9108,N_9448);
xor U10390 (N_10390,N_9399,N_9644);
xnor U10391 (N_10391,N_9458,N_9096);
and U10392 (N_10392,N_9419,N_9658);
and U10393 (N_10393,N_9774,N_9262);
or U10394 (N_10394,N_9738,N_9047);
nand U10395 (N_10395,N_9521,N_9480);
nand U10396 (N_10396,N_9555,N_9163);
nor U10397 (N_10397,N_9177,N_9591);
or U10398 (N_10398,N_9079,N_9279);
xor U10399 (N_10399,N_9721,N_9338);
xnor U10400 (N_10400,N_9067,N_9286);
nand U10401 (N_10401,N_9679,N_9781);
or U10402 (N_10402,N_9130,N_9957);
xor U10403 (N_10403,N_9345,N_9075);
and U10404 (N_10404,N_9423,N_9767);
or U10405 (N_10405,N_9828,N_9150);
or U10406 (N_10406,N_9763,N_9005);
xnor U10407 (N_10407,N_9223,N_9937);
nand U10408 (N_10408,N_9455,N_9661);
and U10409 (N_10409,N_9446,N_9453);
and U10410 (N_10410,N_9302,N_9018);
xor U10411 (N_10411,N_9973,N_9618);
or U10412 (N_10412,N_9151,N_9729);
nor U10413 (N_10413,N_9110,N_9909);
nand U10414 (N_10414,N_9153,N_9569);
nor U10415 (N_10415,N_9664,N_9878);
and U10416 (N_10416,N_9643,N_9113);
xor U10417 (N_10417,N_9846,N_9640);
xnor U10418 (N_10418,N_9114,N_9522);
or U10419 (N_10419,N_9632,N_9269);
xor U10420 (N_10420,N_9409,N_9278);
xnor U10421 (N_10421,N_9834,N_9775);
or U10422 (N_10422,N_9902,N_9507);
nand U10423 (N_10423,N_9091,N_9010);
and U10424 (N_10424,N_9340,N_9254);
xor U10425 (N_10425,N_9742,N_9104);
nor U10426 (N_10426,N_9372,N_9000);
and U10427 (N_10427,N_9165,N_9786);
nand U10428 (N_10428,N_9083,N_9050);
nand U10429 (N_10429,N_9485,N_9851);
nor U10430 (N_10430,N_9070,N_9546);
nand U10431 (N_10431,N_9689,N_9614);
and U10432 (N_10432,N_9586,N_9234);
and U10433 (N_10433,N_9038,N_9727);
xor U10434 (N_10434,N_9908,N_9951);
xnor U10435 (N_10435,N_9145,N_9383);
nor U10436 (N_10436,N_9166,N_9754);
nand U10437 (N_10437,N_9888,N_9443);
or U10438 (N_10438,N_9855,N_9270);
nand U10439 (N_10439,N_9976,N_9355);
and U10440 (N_10440,N_9652,N_9054);
nand U10441 (N_10441,N_9490,N_9196);
xnor U10442 (N_10442,N_9299,N_9136);
and U10443 (N_10443,N_9889,N_9989);
or U10444 (N_10444,N_9616,N_9505);
and U10445 (N_10445,N_9468,N_9064);
or U10446 (N_10446,N_9465,N_9882);
and U10447 (N_10447,N_9209,N_9001);
or U10448 (N_10448,N_9579,N_9732);
or U10449 (N_10449,N_9536,N_9016);
and U10450 (N_10450,N_9623,N_9044);
and U10451 (N_10451,N_9042,N_9575);
nor U10452 (N_10452,N_9843,N_9817);
nor U10453 (N_10453,N_9261,N_9859);
xor U10454 (N_10454,N_9323,N_9611);
and U10455 (N_10455,N_9635,N_9213);
or U10456 (N_10456,N_9504,N_9440);
nor U10457 (N_10457,N_9901,N_9629);
and U10458 (N_10458,N_9084,N_9436);
xnor U10459 (N_10459,N_9597,N_9683);
and U10460 (N_10460,N_9497,N_9156);
xor U10461 (N_10461,N_9246,N_9030);
nor U10462 (N_10462,N_9711,N_9814);
and U10463 (N_10463,N_9285,N_9307);
xnor U10464 (N_10464,N_9770,N_9119);
xnor U10465 (N_10465,N_9819,N_9179);
nand U10466 (N_10466,N_9749,N_9229);
or U10467 (N_10467,N_9977,N_9055);
or U10468 (N_10468,N_9053,N_9952);
and U10469 (N_10469,N_9202,N_9441);
nand U10470 (N_10470,N_9715,N_9940);
and U10471 (N_10471,N_9319,N_9315);
or U10472 (N_10472,N_9572,N_9259);
and U10473 (N_10473,N_9425,N_9548);
xor U10474 (N_10474,N_9359,N_9625);
and U10475 (N_10475,N_9143,N_9674);
nor U10476 (N_10476,N_9692,N_9669);
or U10477 (N_10477,N_9290,N_9936);
nor U10478 (N_10478,N_9801,N_9581);
nor U10479 (N_10479,N_9969,N_9271);
xnor U10480 (N_10480,N_9847,N_9756);
nor U10481 (N_10481,N_9295,N_9965);
and U10482 (N_10482,N_9514,N_9511);
or U10483 (N_10483,N_9488,N_9264);
and U10484 (N_10484,N_9663,N_9564);
xnor U10485 (N_10485,N_9344,N_9701);
or U10486 (N_10486,N_9657,N_9800);
nor U10487 (N_10487,N_9955,N_9417);
nand U10488 (N_10488,N_9731,N_9795);
nor U10489 (N_10489,N_9697,N_9780);
xor U10490 (N_10490,N_9284,N_9782);
and U10491 (N_10491,N_9263,N_9925);
nor U10492 (N_10492,N_9551,N_9904);
nor U10493 (N_10493,N_9280,N_9907);
and U10494 (N_10494,N_9776,N_9810);
nand U10495 (N_10495,N_9176,N_9386);
nor U10496 (N_10496,N_9873,N_9920);
nor U10497 (N_10497,N_9305,N_9238);
and U10498 (N_10498,N_9015,N_9274);
nor U10499 (N_10499,N_9395,N_9790);
or U10500 (N_10500,N_9555,N_9342);
or U10501 (N_10501,N_9585,N_9133);
nor U10502 (N_10502,N_9587,N_9418);
or U10503 (N_10503,N_9664,N_9311);
xnor U10504 (N_10504,N_9785,N_9039);
or U10505 (N_10505,N_9838,N_9206);
and U10506 (N_10506,N_9420,N_9508);
or U10507 (N_10507,N_9236,N_9935);
nor U10508 (N_10508,N_9045,N_9244);
nor U10509 (N_10509,N_9840,N_9518);
and U10510 (N_10510,N_9723,N_9510);
and U10511 (N_10511,N_9784,N_9168);
xor U10512 (N_10512,N_9084,N_9239);
or U10513 (N_10513,N_9843,N_9362);
xor U10514 (N_10514,N_9072,N_9142);
nor U10515 (N_10515,N_9297,N_9947);
nor U10516 (N_10516,N_9822,N_9759);
nor U10517 (N_10517,N_9851,N_9389);
xnor U10518 (N_10518,N_9573,N_9593);
nand U10519 (N_10519,N_9134,N_9296);
and U10520 (N_10520,N_9470,N_9464);
xnor U10521 (N_10521,N_9373,N_9846);
and U10522 (N_10522,N_9381,N_9909);
nand U10523 (N_10523,N_9555,N_9016);
nor U10524 (N_10524,N_9066,N_9278);
nor U10525 (N_10525,N_9566,N_9902);
and U10526 (N_10526,N_9430,N_9420);
nor U10527 (N_10527,N_9994,N_9563);
and U10528 (N_10528,N_9377,N_9208);
or U10529 (N_10529,N_9010,N_9139);
nor U10530 (N_10530,N_9679,N_9167);
nor U10531 (N_10531,N_9870,N_9476);
and U10532 (N_10532,N_9251,N_9413);
nor U10533 (N_10533,N_9084,N_9552);
and U10534 (N_10534,N_9107,N_9739);
nor U10535 (N_10535,N_9751,N_9883);
and U10536 (N_10536,N_9049,N_9606);
or U10537 (N_10537,N_9847,N_9514);
nor U10538 (N_10538,N_9002,N_9618);
nand U10539 (N_10539,N_9346,N_9292);
and U10540 (N_10540,N_9762,N_9483);
nor U10541 (N_10541,N_9976,N_9776);
and U10542 (N_10542,N_9824,N_9049);
nand U10543 (N_10543,N_9476,N_9210);
nor U10544 (N_10544,N_9100,N_9320);
nand U10545 (N_10545,N_9773,N_9391);
nand U10546 (N_10546,N_9404,N_9260);
nor U10547 (N_10547,N_9220,N_9175);
and U10548 (N_10548,N_9253,N_9401);
nand U10549 (N_10549,N_9117,N_9663);
and U10550 (N_10550,N_9153,N_9915);
nor U10551 (N_10551,N_9697,N_9434);
nor U10552 (N_10552,N_9385,N_9441);
and U10553 (N_10553,N_9583,N_9323);
nor U10554 (N_10554,N_9458,N_9437);
and U10555 (N_10555,N_9143,N_9943);
xnor U10556 (N_10556,N_9445,N_9694);
or U10557 (N_10557,N_9750,N_9992);
and U10558 (N_10558,N_9211,N_9450);
xnor U10559 (N_10559,N_9617,N_9337);
nor U10560 (N_10560,N_9507,N_9940);
and U10561 (N_10561,N_9400,N_9613);
and U10562 (N_10562,N_9937,N_9990);
nand U10563 (N_10563,N_9031,N_9450);
and U10564 (N_10564,N_9213,N_9500);
xnor U10565 (N_10565,N_9046,N_9605);
and U10566 (N_10566,N_9938,N_9603);
nand U10567 (N_10567,N_9640,N_9397);
nor U10568 (N_10568,N_9884,N_9788);
or U10569 (N_10569,N_9494,N_9294);
and U10570 (N_10570,N_9876,N_9170);
or U10571 (N_10571,N_9773,N_9752);
xnor U10572 (N_10572,N_9400,N_9188);
and U10573 (N_10573,N_9598,N_9033);
and U10574 (N_10574,N_9884,N_9295);
or U10575 (N_10575,N_9278,N_9852);
nand U10576 (N_10576,N_9265,N_9753);
or U10577 (N_10577,N_9734,N_9404);
xnor U10578 (N_10578,N_9940,N_9295);
xor U10579 (N_10579,N_9713,N_9928);
and U10580 (N_10580,N_9144,N_9862);
xor U10581 (N_10581,N_9621,N_9762);
xnor U10582 (N_10582,N_9517,N_9125);
nor U10583 (N_10583,N_9435,N_9199);
and U10584 (N_10584,N_9580,N_9216);
nand U10585 (N_10585,N_9066,N_9595);
nor U10586 (N_10586,N_9595,N_9022);
nand U10587 (N_10587,N_9552,N_9502);
and U10588 (N_10588,N_9766,N_9996);
nand U10589 (N_10589,N_9518,N_9705);
and U10590 (N_10590,N_9019,N_9458);
nand U10591 (N_10591,N_9198,N_9014);
nand U10592 (N_10592,N_9553,N_9786);
and U10593 (N_10593,N_9153,N_9969);
xor U10594 (N_10594,N_9171,N_9713);
xor U10595 (N_10595,N_9568,N_9118);
nand U10596 (N_10596,N_9123,N_9384);
and U10597 (N_10597,N_9089,N_9520);
and U10598 (N_10598,N_9684,N_9394);
nand U10599 (N_10599,N_9193,N_9882);
nor U10600 (N_10600,N_9750,N_9599);
nor U10601 (N_10601,N_9773,N_9035);
nor U10602 (N_10602,N_9160,N_9255);
or U10603 (N_10603,N_9158,N_9850);
or U10604 (N_10604,N_9422,N_9925);
xor U10605 (N_10605,N_9294,N_9248);
nor U10606 (N_10606,N_9190,N_9695);
or U10607 (N_10607,N_9109,N_9754);
nor U10608 (N_10608,N_9093,N_9978);
and U10609 (N_10609,N_9608,N_9153);
xnor U10610 (N_10610,N_9638,N_9233);
nor U10611 (N_10611,N_9577,N_9181);
and U10612 (N_10612,N_9708,N_9913);
nand U10613 (N_10613,N_9882,N_9425);
and U10614 (N_10614,N_9950,N_9401);
nor U10615 (N_10615,N_9437,N_9090);
nand U10616 (N_10616,N_9948,N_9872);
or U10617 (N_10617,N_9547,N_9005);
nor U10618 (N_10618,N_9239,N_9294);
and U10619 (N_10619,N_9457,N_9645);
or U10620 (N_10620,N_9676,N_9634);
and U10621 (N_10621,N_9985,N_9877);
xor U10622 (N_10622,N_9394,N_9771);
or U10623 (N_10623,N_9577,N_9327);
nor U10624 (N_10624,N_9915,N_9743);
or U10625 (N_10625,N_9992,N_9848);
xor U10626 (N_10626,N_9563,N_9041);
xor U10627 (N_10627,N_9199,N_9781);
nand U10628 (N_10628,N_9068,N_9058);
nor U10629 (N_10629,N_9726,N_9453);
or U10630 (N_10630,N_9210,N_9547);
xnor U10631 (N_10631,N_9865,N_9476);
nand U10632 (N_10632,N_9941,N_9140);
nand U10633 (N_10633,N_9326,N_9873);
or U10634 (N_10634,N_9969,N_9810);
xor U10635 (N_10635,N_9073,N_9859);
nor U10636 (N_10636,N_9767,N_9425);
nand U10637 (N_10637,N_9983,N_9063);
nand U10638 (N_10638,N_9908,N_9485);
nor U10639 (N_10639,N_9790,N_9957);
nor U10640 (N_10640,N_9977,N_9091);
xnor U10641 (N_10641,N_9617,N_9430);
nor U10642 (N_10642,N_9339,N_9494);
nor U10643 (N_10643,N_9858,N_9353);
nor U10644 (N_10644,N_9571,N_9668);
or U10645 (N_10645,N_9591,N_9198);
and U10646 (N_10646,N_9879,N_9964);
or U10647 (N_10647,N_9057,N_9318);
nor U10648 (N_10648,N_9122,N_9942);
and U10649 (N_10649,N_9009,N_9372);
and U10650 (N_10650,N_9631,N_9891);
and U10651 (N_10651,N_9086,N_9299);
or U10652 (N_10652,N_9430,N_9552);
and U10653 (N_10653,N_9561,N_9871);
nand U10654 (N_10654,N_9773,N_9342);
xor U10655 (N_10655,N_9216,N_9099);
nand U10656 (N_10656,N_9929,N_9875);
nand U10657 (N_10657,N_9885,N_9518);
and U10658 (N_10658,N_9019,N_9460);
and U10659 (N_10659,N_9303,N_9261);
or U10660 (N_10660,N_9206,N_9379);
nand U10661 (N_10661,N_9848,N_9466);
xor U10662 (N_10662,N_9772,N_9648);
xnor U10663 (N_10663,N_9037,N_9103);
and U10664 (N_10664,N_9222,N_9939);
xor U10665 (N_10665,N_9171,N_9410);
nand U10666 (N_10666,N_9809,N_9138);
xor U10667 (N_10667,N_9725,N_9671);
and U10668 (N_10668,N_9063,N_9855);
and U10669 (N_10669,N_9214,N_9838);
nand U10670 (N_10670,N_9561,N_9366);
nand U10671 (N_10671,N_9423,N_9498);
nand U10672 (N_10672,N_9711,N_9714);
nor U10673 (N_10673,N_9623,N_9882);
and U10674 (N_10674,N_9636,N_9996);
or U10675 (N_10675,N_9667,N_9649);
xnor U10676 (N_10676,N_9524,N_9825);
and U10677 (N_10677,N_9513,N_9254);
and U10678 (N_10678,N_9025,N_9252);
or U10679 (N_10679,N_9241,N_9754);
nor U10680 (N_10680,N_9903,N_9522);
or U10681 (N_10681,N_9737,N_9218);
xor U10682 (N_10682,N_9235,N_9060);
xnor U10683 (N_10683,N_9974,N_9544);
nand U10684 (N_10684,N_9937,N_9748);
and U10685 (N_10685,N_9824,N_9864);
or U10686 (N_10686,N_9241,N_9638);
nor U10687 (N_10687,N_9412,N_9102);
or U10688 (N_10688,N_9829,N_9915);
nand U10689 (N_10689,N_9261,N_9808);
nand U10690 (N_10690,N_9479,N_9436);
and U10691 (N_10691,N_9581,N_9041);
nand U10692 (N_10692,N_9399,N_9729);
nand U10693 (N_10693,N_9990,N_9214);
and U10694 (N_10694,N_9151,N_9532);
or U10695 (N_10695,N_9653,N_9056);
xor U10696 (N_10696,N_9314,N_9249);
nor U10697 (N_10697,N_9167,N_9421);
nand U10698 (N_10698,N_9163,N_9213);
nor U10699 (N_10699,N_9187,N_9918);
or U10700 (N_10700,N_9226,N_9003);
and U10701 (N_10701,N_9233,N_9948);
nand U10702 (N_10702,N_9813,N_9524);
nand U10703 (N_10703,N_9147,N_9679);
xnor U10704 (N_10704,N_9403,N_9189);
or U10705 (N_10705,N_9566,N_9962);
and U10706 (N_10706,N_9269,N_9361);
nand U10707 (N_10707,N_9983,N_9313);
nor U10708 (N_10708,N_9254,N_9229);
and U10709 (N_10709,N_9496,N_9205);
nand U10710 (N_10710,N_9083,N_9314);
nor U10711 (N_10711,N_9305,N_9760);
and U10712 (N_10712,N_9366,N_9580);
nand U10713 (N_10713,N_9305,N_9378);
nor U10714 (N_10714,N_9354,N_9293);
nand U10715 (N_10715,N_9699,N_9139);
xnor U10716 (N_10716,N_9728,N_9524);
xor U10717 (N_10717,N_9231,N_9299);
or U10718 (N_10718,N_9559,N_9303);
and U10719 (N_10719,N_9433,N_9072);
nand U10720 (N_10720,N_9256,N_9752);
and U10721 (N_10721,N_9893,N_9077);
and U10722 (N_10722,N_9684,N_9900);
or U10723 (N_10723,N_9824,N_9822);
and U10724 (N_10724,N_9734,N_9603);
nand U10725 (N_10725,N_9248,N_9010);
nand U10726 (N_10726,N_9965,N_9583);
or U10727 (N_10727,N_9983,N_9103);
nor U10728 (N_10728,N_9387,N_9203);
or U10729 (N_10729,N_9416,N_9315);
nor U10730 (N_10730,N_9575,N_9456);
xor U10731 (N_10731,N_9355,N_9292);
xor U10732 (N_10732,N_9921,N_9407);
nor U10733 (N_10733,N_9621,N_9527);
nand U10734 (N_10734,N_9190,N_9395);
nor U10735 (N_10735,N_9993,N_9291);
and U10736 (N_10736,N_9185,N_9372);
nor U10737 (N_10737,N_9862,N_9132);
or U10738 (N_10738,N_9413,N_9607);
and U10739 (N_10739,N_9827,N_9258);
xnor U10740 (N_10740,N_9598,N_9168);
and U10741 (N_10741,N_9392,N_9693);
nor U10742 (N_10742,N_9174,N_9283);
xnor U10743 (N_10743,N_9844,N_9469);
nor U10744 (N_10744,N_9216,N_9495);
nand U10745 (N_10745,N_9157,N_9282);
or U10746 (N_10746,N_9694,N_9259);
or U10747 (N_10747,N_9262,N_9240);
nand U10748 (N_10748,N_9951,N_9109);
nor U10749 (N_10749,N_9495,N_9532);
nand U10750 (N_10750,N_9017,N_9044);
or U10751 (N_10751,N_9256,N_9084);
xor U10752 (N_10752,N_9849,N_9225);
nand U10753 (N_10753,N_9229,N_9152);
nand U10754 (N_10754,N_9560,N_9972);
nand U10755 (N_10755,N_9475,N_9641);
xor U10756 (N_10756,N_9538,N_9190);
xor U10757 (N_10757,N_9508,N_9702);
nor U10758 (N_10758,N_9471,N_9248);
nand U10759 (N_10759,N_9317,N_9794);
nand U10760 (N_10760,N_9586,N_9293);
and U10761 (N_10761,N_9853,N_9364);
nand U10762 (N_10762,N_9927,N_9030);
or U10763 (N_10763,N_9178,N_9046);
nand U10764 (N_10764,N_9160,N_9956);
xor U10765 (N_10765,N_9618,N_9177);
nor U10766 (N_10766,N_9214,N_9728);
or U10767 (N_10767,N_9001,N_9454);
and U10768 (N_10768,N_9700,N_9763);
and U10769 (N_10769,N_9120,N_9039);
nor U10770 (N_10770,N_9539,N_9591);
nor U10771 (N_10771,N_9718,N_9125);
or U10772 (N_10772,N_9483,N_9298);
xor U10773 (N_10773,N_9445,N_9052);
nor U10774 (N_10774,N_9210,N_9687);
nand U10775 (N_10775,N_9909,N_9775);
or U10776 (N_10776,N_9435,N_9816);
nor U10777 (N_10777,N_9306,N_9313);
nor U10778 (N_10778,N_9970,N_9142);
xnor U10779 (N_10779,N_9097,N_9836);
xnor U10780 (N_10780,N_9088,N_9490);
or U10781 (N_10781,N_9108,N_9103);
nand U10782 (N_10782,N_9984,N_9217);
xor U10783 (N_10783,N_9723,N_9719);
or U10784 (N_10784,N_9855,N_9435);
nor U10785 (N_10785,N_9439,N_9081);
nand U10786 (N_10786,N_9611,N_9575);
and U10787 (N_10787,N_9283,N_9919);
nand U10788 (N_10788,N_9925,N_9198);
and U10789 (N_10789,N_9427,N_9968);
nor U10790 (N_10790,N_9782,N_9582);
nor U10791 (N_10791,N_9708,N_9401);
or U10792 (N_10792,N_9055,N_9497);
nand U10793 (N_10793,N_9382,N_9629);
xor U10794 (N_10794,N_9000,N_9288);
or U10795 (N_10795,N_9548,N_9840);
and U10796 (N_10796,N_9669,N_9741);
xor U10797 (N_10797,N_9715,N_9616);
nand U10798 (N_10798,N_9048,N_9350);
nor U10799 (N_10799,N_9950,N_9493);
nor U10800 (N_10800,N_9520,N_9508);
nor U10801 (N_10801,N_9427,N_9574);
nor U10802 (N_10802,N_9922,N_9176);
or U10803 (N_10803,N_9011,N_9849);
nor U10804 (N_10804,N_9873,N_9476);
nand U10805 (N_10805,N_9438,N_9756);
and U10806 (N_10806,N_9306,N_9372);
nand U10807 (N_10807,N_9555,N_9238);
nand U10808 (N_10808,N_9096,N_9357);
nand U10809 (N_10809,N_9263,N_9539);
and U10810 (N_10810,N_9790,N_9948);
nand U10811 (N_10811,N_9841,N_9746);
xor U10812 (N_10812,N_9136,N_9851);
nor U10813 (N_10813,N_9049,N_9602);
nand U10814 (N_10814,N_9192,N_9576);
and U10815 (N_10815,N_9706,N_9831);
and U10816 (N_10816,N_9958,N_9647);
nand U10817 (N_10817,N_9741,N_9935);
or U10818 (N_10818,N_9055,N_9807);
and U10819 (N_10819,N_9080,N_9544);
xor U10820 (N_10820,N_9314,N_9573);
xnor U10821 (N_10821,N_9751,N_9301);
xnor U10822 (N_10822,N_9494,N_9483);
nand U10823 (N_10823,N_9826,N_9123);
nand U10824 (N_10824,N_9434,N_9981);
and U10825 (N_10825,N_9522,N_9021);
and U10826 (N_10826,N_9001,N_9512);
nand U10827 (N_10827,N_9897,N_9663);
nor U10828 (N_10828,N_9302,N_9570);
nand U10829 (N_10829,N_9426,N_9190);
or U10830 (N_10830,N_9708,N_9714);
xor U10831 (N_10831,N_9758,N_9947);
nand U10832 (N_10832,N_9395,N_9697);
nand U10833 (N_10833,N_9016,N_9168);
xor U10834 (N_10834,N_9765,N_9555);
and U10835 (N_10835,N_9436,N_9992);
xnor U10836 (N_10836,N_9375,N_9259);
or U10837 (N_10837,N_9043,N_9403);
nand U10838 (N_10838,N_9549,N_9777);
nor U10839 (N_10839,N_9353,N_9871);
xor U10840 (N_10840,N_9730,N_9355);
or U10841 (N_10841,N_9049,N_9941);
or U10842 (N_10842,N_9529,N_9325);
nand U10843 (N_10843,N_9507,N_9492);
nand U10844 (N_10844,N_9894,N_9093);
nand U10845 (N_10845,N_9827,N_9517);
nor U10846 (N_10846,N_9915,N_9906);
xnor U10847 (N_10847,N_9832,N_9736);
nand U10848 (N_10848,N_9325,N_9455);
and U10849 (N_10849,N_9426,N_9565);
and U10850 (N_10850,N_9885,N_9049);
nor U10851 (N_10851,N_9155,N_9516);
or U10852 (N_10852,N_9179,N_9602);
or U10853 (N_10853,N_9248,N_9547);
and U10854 (N_10854,N_9482,N_9154);
nor U10855 (N_10855,N_9811,N_9320);
nand U10856 (N_10856,N_9749,N_9901);
or U10857 (N_10857,N_9707,N_9583);
and U10858 (N_10858,N_9892,N_9974);
nor U10859 (N_10859,N_9298,N_9791);
xor U10860 (N_10860,N_9743,N_9163);
xor U10861 (N_10861,N_9596,N_9626);
or U10862 (N_10862,N_9235,N_9124);
and U10863 (N_10863,N_9274,N_9367);
or U10864 (N_10864,N_9806,N_9727);
xnor U10865 (N_10865,N_9686,N_9401);
nor U10866 (N_10866,N_9607,N_9480);
and U10867 (N_10867,N_9463,N_9454);
nor U10868 (N_10868,N_9217,N_9973);
xor U10869 (N_10869,N_9719,N_9823);
xor U10870 (N_10870,N_9226,N_9535);
and U10871 (N_10871,N_9265,N_9153);
or U10872 (N_10872,N_9030,N_9530);
xnor U10873 (N_10873,N_9763,N_9072);
or U10874 (N_10874,N_9712,N_9839);
xor U10875 (N_10875,N_9567,N_9935);
nand U10876 (N_10876,N_9123,N_9785);
xnor U10877 (N_10877,N_9593,N_9478);
xnor U10878 (N_10878,N_9323,N_9118);
nand U10879 (N_10879,N_9096,N_9878);
xnor U10880 (N_10880,N_9907,N_9565);
or U10881 (N_10881,N_9526,N_9697);
or U10882 (N_10882,N_9792,N_9283);
and U10883 (N_10883,N_9830,N_9064);
xnor U10884 (N_10884,N_9442,N_9952);
or U10885 (N_10885,N_9908,N_9704);
and U10886 (N_10886,N_9616,N_9941);
and U10887 (N_10887,N_9828,N_9384);
nor U10888 (N_10888,N_9842,N_9565);
xnor U10889 (N_10889,N_9788,N_9135);
xor U10890 (N_10890,N_9541,N_9899);
nand U10891 (N_10891,N_9685,N_9384);
xor U10892 (N_10892,N_9187,N_9313);
nor U10893 (N_10893,N_9446,N_9673);
or U10894 (N_10894,N_9448,N_9489);
xnor U10895 (N_10895,N_9941,N_9458);
or U10896 (N_10896,N_9767,N_9524);
nand U10897 (N_10897,N_9443,N_9933);
nor U10898 (N_10898,N_9171,N_9614);
and U10899 (N_10899,N_9182,N_9990);
nand U10900 (N_10900,N_9764,N_9763);
or U10901 (N_10901,N_9868,N_9310);
nor U10902 (N_10902,N_9930,N_9210);
nand U10903 (N_10903,N_9098,N_9123);
and U10904 (N_10904,N_9615,N_9993);
and U10905 (N_10905,N_9893,N_9190);
nor U10906 (N_10906,N_9213,N_9558);
nor U10907 (N_10907,N_9421,N_9053);
or U10908 (N_10908,N_9908,N_9965);
nand U10909 (N_10909,N_9850,N_9429);
xnor U10910 (N_10910,N_9617,N_9507);
nor U10911 (N_10911,N_9669,N_9557);
xnor U10912 (N_10912,N_9538,N_9735);
xnor U10913 (N_10913,N_9396,N_9896);
nor U10914 (N_10914,N_9977,N_9265);
xor U10915 (N_10915,N_9739,N_9159);
nand U10916 (N_10916,N_9087,N_9762);
and U10917 (N_10917,N_9254,N_9754);
nand U10918 (N_10918,N_9608,N_9699);
xor U10919 (N_10919,N_9129,N_9350);
or U10920 (N_10920,N_9699,N_9798);
nor U10921 (N_10921,N_9281,N_9056);
nand U10922 (N_10922,N_9469,N_9049);
or U10923 (N_10923,N_9390,N_9599);
xor U10924 (N_10924,N_9368,N_9732);
and U10925 (N_10925,N_9203,N_9582);
and U10926 (N_10926,N_9123,N_9048);
or U10927 (N_10927,N_9050,N_9704);
xor U10928 (N_10928,N_9080,N_9633);
nor U10929 (N_10929,N_9791,N_9805);
nand U10930 (N_10930,N_9466,N_9307);
and U10931 (N_10931,N_9999,N_9205);
nor U10932 (N_10932,N_9188,N_9936);
nor U10933 (N_10933,N_9614,N_9889);
and U10934 (N_10934,N_9220,N_9989);
xor U10935 (N_10935,N_9961,N_9890);
nand U10936 (N_10936,N_9972,N_9213);
nand U10937 (N_10937,N_9768,N_9951);
nand U10938 (N_10938,N_9064,N_9298);
nand U10939 (N_10939,N_9459,N_9675);
nor U10940 (N_10940,N_9394,N_9932);
and U10941 (N_10941,N_9152,N_9737);
xnor U10942 (N_10942,N_9859,N_9537);
or U10943 (N_10943,N_9935,N_9190);
xnor U10944 (N_10944,N_9348,N_9803);
xnor U10945 (N_10945,N_9406,N_9970);
nor U10946 (N_10946,N_9591,N_9134);
or U10947 (N_10947,N_9133,N_9978);
or U10948 (N_10948,N_9751,N_9440);
xnor U10949 (N_10949,N_9565,N_9452);
nand U10950 (N_10950,N_9561,N_9149);
nor U10951 (N_10951,N_9716,N_9564);
and U10952 (N_10952,N_9591,N_9692);
or U10953 (N_10953,N_9778,N_9631);
or U10954 (N_10954,N_9228,N_9135);
nand U10955 (N_10955,N_9044,N_9060);
nor U10956 (N_10956,N_9462,N_9927);
nor U10957 (N_10957,N_9292,N_9829);
xor U10958 (N_10958,N_9200,N_9274);
nand U10959 (N_10959,N_9381,N_9392);
nor U10960 (N_10960,N_9057,N_9973);
or U10961 (N_10961,N_9832,N_9844);
and U10962 (N_10962,N_9819,N_9156);
xor U10963 (N_10963,N_9115,N_9579);
nor U10964 (N_10964,N_9783,N_9906);
nand U10965 (N_10965,N_9864,N_9389);
nor U10966 (N_10966,N_9472,N_9865);
nand U10967 (N_10967,N_9676,N_9542);
xnor U10968 (N_10968,N_9756,N_9058);
nor U10969 (N_10969,N_9695,N_9861);
xnor U10970 (N_10970,N_9755,N_9232);
or U10971 (N_10971,N_9810,N_9351);
or U10972 (N_10972,N_9064,N_9721);
or U10973 (N_10973,N_9552,N_9575);
xnor U10974 (N_10974,N_9495,N_9632);
or U10975 (N_10975,N_9987,N_9181);
nor U10976 (N_10976,N_9426,N_9287);
nand U10977 (N_10977,N_9457,N_9271);
xor U10978 (N_10978,N_9368,N_9434);
nor U10979 (N_10979,N_9553,N_9826);
xnor U10980 (N_10980,N_9433,N_9617);
or U10981 (N_10981,N_9733,N_9653);
or U10982 (N_10982,N_9199,N_9814);
nand U10983 (N_10983,N_9457,N_9940);
and U10984 (N_10984,N_9036,N_9758);
and U10985 (N_10985,N_9508,N_9544);
and U10986 (N_10986,N_9535,N_9496);
and U10987 (N_10987,N_9596,N_9729);
or U10988 (N_10988,N_9032,N_9843);
nand U10989 (N_10989,N_9348,N_9740);
nand U10990 (N_10990,N_9859,N_9048);
nand U10991 (N_10991,N_9934,N_9175);
nand U10992 (N_10992,N_9799,N_9770);
xnor U10993 (N_10993,N_9903,N_9995);
xnor U10994 (N_10994,N_9883,N_9479);
or U10995 (N_10995,N_9125,N_9105);
nand U10996 (N_10996,N_9425,N_9707);
xor U10997 (N_10997,N_9175,N_9552);
xor U10998 (N_10998,N_9153,N_9234);
or U10999 (N_10999,N_9386,N_9393);
nand U11000 (N_11000,N_10095,N_10027);
xor U11001 (N_11001,N_10149,N_10313);
or U11002 (N_11002,N_10425,N_10742);
nand U11003 (N_11003,N_10104,N_10227);
nor U11004 (N_11004,N_10760,N_10271);
nor U11005 (N_11005,N_10502,N_10590);
nand U11006 (N_11006,N_10993,N_10430);
nand U11007 (N_11007,N_10439,N_10209);
nor U11008 (N_11008,N_10044,N_10967);
or U11009 (N_11009,N_10112,N_10142);
xor U11010 (N_11010,N_10306,N_10648);
nor U11011 (N_11011,N_10485,N_10900);
nor U11012 (N_11012,N_10922,N_10554);
or U11013 (N_11013,N_10806,N_10193);
and U11014 (N_11014,N_10756,N_10436);
nor U11015 (N_11015,N_10917,N_10228);
and U11016 (N_11016,N_10492,N_10162);
xnor U11017 (N_11017,N_10921,N_10605);
nor U11018 (N_11018,N_10048,N_10717);
nand U11019 (N_11019,N_10270,N_10217);
xnor U11020 (N_11020,N_10232,N_10643);
or U11021 (N_11021,N_10873,N_10132);
or U11022 (N_11022,N_10121,N_10595);
or U11023 (N_11023,N_10958,N_10723);
or U11024 (N_11024,N_10317,N_10931);
nand U11025 (N_11025,N_10100,N_10429);
or U11026 (N_11026,N_10542,N_10081);
nand U11027 (N_11027,N_10692,N_10892);
xor U11028 (N_11028,N_10389,N_10582);
or U11029 (N_11029,N_10600,N_10196);
xnor U11030 (N_11030,N_10072,N_10418);
or U11031 (N_11031,N_10963,N_10062);
nand U11032 (N_11032,N_10634,N_10224);
xnor U11033 (N_11033,N_10949,N_10693);
nor U11034 (N_11034,N_10729,N_10243);
nand U11035 (N_11035,N_10663,N_10879);
and U11036 (N_11036,N_10122,N_10810);
nand U11037 (N_11037,N_10221,N_10655);
nor U11038 (N_11038,N_10844,N_10627);
and U11039 (N_11039,N_10177,N_10744);
xnor U11040 (N_11040,N_10906,N_10815);
or U11041 (N_11041,N_10323,N_10514);
nand U11042 (N_11042,N_10036,N_10866);
nor U11043 (N_11043,N_10803,N_10608);
xor U11044 (N_11044,N_10630,N_10666);
nor U11045 (N_11045,N_10686,N_10998);
xor U11046 (N_11046,N_10965,N_10423);
nand U11047 (N_11047,N_10982,N_10901);
and U11048 (N_11048,N_10312,N_10195);
and U11049 (N_11049,N_10083,N_10335);
or U11050 (N_11050,N_10570,N_10918);
or U11051 (N_11051,N_10898,N_10645);
and U11052 (N_11052,N_10356,N_10461);
nand U11053 (N_11053,N_10286,N_10792);
nor U11054 (N_11054,N_10427,N_10457);
nand U11055 (N_11055,N_10831,N_10626);
and U11056 (N_11056,N_10651,N_10490);
nor U11057 (N_11057,N_10962,N_10231);
nand U11058 (N_11058,N_10416,N_10604);
nor U11059 (N_11059,N_10825,N_10518);
xnor U11060 (N_11060,N_10254,N_10843);
and U11061 (N_11061,N_10333,N_10936);
and U11062 (N_11062,N_10449,N_10813);
and U11063 (N_11063,N_10611,N_10226);
xnor U11064 (N_11064,N_10888,N_10442);
or U11065 (N_11065,N_10020,N_10212);
and U11066 (N_11066,N_10553,N_10732);
nand U11067 (N_11067,N_10262,N_10008);
xnor U11068 (N_11068,N_10240,N_10956);
xnor U11069 (N_11069,N_10566,N_10580);
and U11070 (N_11070,N_10688,N_10373);
and U11071 (N_11071,N_10598,N_10509);
or U11072 (N_11072,N_10417,N_10755);
nor U11073 (N_11073,N_10158,N_10536);
nand U11074 (N_11074,N_10491,N_10804);
xor U11075 (N_11075,N_10948,N_10912);
xnor U11076 (N_11076,N_10871,N_10839);
xnor U11077 (N_11077,N_10125,N_10239);
or U11078 (N_11078,N_10853,N_10404);
or U11079 (N_11079,N_10781,N_10156);
xor U11080 (N_11080,N_10776,N_10043);
nand U11081 (N_11081,N_10073,N_10143);
nand U11082 (N_11082,N_10650,N_10618);
nor U11083 (N_11083,N_10159,N_10926);
or U11084 (N_11084,N_10510,N_10690);
nor U11085 (N_11085,N_10077,N_10585);
nor U11086 (N_11086,N_10710,N_10068);
or U11087 (N_11087,N_10625,N_10620);
and U11088 (N_11088,N_10471,N_10876);
nor U11089 (N_11089,N_10127,N_10896);
or U11090 (N_11090,N_10115,N_10444);
nand U11091 (N_11091,N_10574,N_10205);
nor U11092 (N_11092,N_10953,N_10552);
and U11093 (N_11093,N_10376,N_10114);
or U11094 (N_11094,N_10285,N_10550);
or U11095 (N_11095,N_10342,N_10406);
or U11096 (N_11096,N_10653,N_10292);
xor U11097 (N_11097,N_10378,N_10654);
and U11098 (N_11098,N_10332,N_10836);
nand U11099 (N_11099,N_10116,N_10517);
xor U11100 (N_11100,N_10622,N_10768);
nor U11101 (N_11101,N_10434,N_10652);
or U11102 (N_11102,N_10204,N_10763);
xnor U11103 (N_11103,N_10206,N_10208);
or U11104 (N_11104,N_10414,N_10327);
nor U11105 (N_11105,N_10002,N_10991);
nand U11106 (N_11106,N_10636,N_10034);
and U11107 (N_11107,N_10004,N_10396);
and U11108 (N_11108,N_10950,N_10326);
and U11109 (N_11109,N_10191,N_10802);
or U11110 (N_11110,N_10555,N_10472);
nand U11111 (N_11111,N_10097,N_10631);
or U11112 (N_11112,N_10338,N_10042);
nor U11113 (N_11113,N_10126,N_10280);
and U11114 (N_11114,N_10040,N_10828);
nor U11115 (N_11115,N_10798,N_10111);
xor U11116 (N_11116,N_10784,N_10137);
or U11117 (N_11117,N_10054,N_10747);
or U11118 (N_11118,N_10371,N_10259);
and U11119 (N_11119,N_10632,N_10103);
nor U11120 (N_11120,N_10479,N_10568);
and U11121 (N_11121,N_10001,N_10189);
and U11122 (N_11122,N_10129,N_10109);
or U11123 (N_11123,N_10211,N_10973);
or U11124 (N_11124,N_10702,N_10320);
xnor U11125 (N_11125,N_10261,N_10529);
nor U11126 (N_11126,N_10319,N_10697);
nand U11127 (N_11127,N_10420,N_10375);
xor U11128 (N_11128,N_10558,N_10025);
nor U11129 (N_11129,N_10885,N_10505);
and U11130 (N_11130,N_10685,N_10119);
xor U11131 (N_11131,N_10220,N_10593);
nor U11132 (N_11132,N_10513,N_10790);
xor U11133 (N_11133,N_10173,N_10775);
nor U11134 (N_11134,N_10454,N_10480);
xnor U11135 (N_11135,N_10250,N_10266);
nand U11136 (N_11136,N_10037,N_10599);
or U11137 (N_11137,N_10551,N_10021);
and U11138 (N_11138,N_10123,N_10175);
or U11139 (N_11139,N_10233,N_10242);
nand U11140 (N_11140,N_10387,N_10355);
and U11141 (N_11141,N_10649,N_10791);
xor U11142 (N_11142,N_10561,N_10924);
nand U11143 (N_11143,N_10886,N_10464);
or U11144 (N_11144,N_10833,N_10624);
or U11145 (N_11145,N_10909,N_10656);
and U11146 (N_11146,N_10283,N_10672);
nor U11147 (N_11147,N_10153,N_10665);
nor U11148 (N_11148,N_10481,N_10889);
and U11149 (N_11149,N_10238,N_10374);
xnor U11150 (N_11150,N_10782,N_10074);
xnor U11151 (N_11151,N_10493,N_10904);
nand U11152 (N_11152,N_10017,N_10222);
and U11153 (N_11153,N_10758,N_10812);
and U11154 (N_11154,N_10110,N_10639);
and U11155 (N_11155,N_10161,N_10659);
xor U11156 (N_11156,N_10694,N_10579);
nand U11157 (N_11157,N_10478,N_10779);
nor U11158 (N_11158,N_10171,N_10365);
and U11159 (N_11159,N_10923,N_10916);
and U11160 (N_11160,N_10386,N_10977);
nand U11161 (N_11161,N_10287,N_10989);
or U11162 (N_11162,N_10470,N_10051);
xnor U11163 (N_11163,N_10557,N_10133);
or U11164 (N_11164,N_10411,N_10390);
xor U11165 (N_11165,N_10487,N_10468);
nor U11166 (N_11166,N_10296,N_10052);
nand U11167 (N_11167,N_10276,N_10304);
nor U11168 (N_11168,N_10180,N_10147);
or U11169 (N_11169,N_10847,N_10006);
nand U11170 (N_11170,N_10391,N_10541);
nor U11171 (N_11171,N_10264,N_10683);
xnor U11172 (N_11172,N_10814,N_10325);
xor U11173 (N_11173,N_10858,N_10562);
xor U11174 (N_11174,N_10745,N_10281);
nor U11175 (N_11175,N_10489,N_10548);
nand U11176 (N_11176,N_10298,N_10169);
or U11177 (N_11177,N_10671,N_10070);
or U11178 (N_11178,N_10805,N_10015);
xnor U11179 (N_11179,N_10668,N_10609);
and U11180 (N_11180,N_10832,N_10155);
and U11181 (N_11181,N_10684,N_10988);
or U11182 (N_11182,N_10398,N_10720);
nand U11183 (N_11183,N_10533,N_10932);
and U11184 (N_11184,N_10762,N_10951);
and U11185 (N_11185,N_10503,N_10571);
nand U11186 (N_11186,N_10738,N_10640);
nor U11187 (N_11187,N_10165,N_10310);
xnor U11188 (N_11188,N_10474,N_10978);
xnor U11189 (N_11189,N_10249,N_10018);
or U11190 (N_11190,N_10394,N_10026);
nor U11191 (N_11191,N_10340,N_10714);
or U11192 (N_11192,N_10446,N_10199);
xnor U11193 (N_11193,N_10352,N_10531);
or U11194 (N_11194,N_10564,N_10862);
nor U11195 (N_11195,N_10282,N_10581);
nand U11196 (N_11196,N_10065,N_10603);
and U11197 (N_11197,N_10056,N_10475);
nand U11198 (N_11198,N_10589,N_10236);
nand U11199 (N_11199,N_10854,N_10410);
xor U11200 (N_11200,N_10086,N_10361);
and U11201 (N_11201,N_10800,N_10878);
or U11202 (N_11202,N_10687,N_10185);
nor U11203 (N_11203,N_10947,N_10251);
or U11204 (N_11204,N_10178,N_10576);
xnor U11205 (N_11205,N_10013,N_10565);
nand U11206 (N_11206,N_10882,N_10329);
and U11207 (N_11207,N_10827,N_10076);
and U11208 (N_11208,N_10868,N_10028);
nand U11209 (N_11209,N_10770,N_10187);
nor U11210 (N_11210,N_10587,N_10445);
or U11211 (N_11211,N_10560,N_10456);
nand U11212 (N_11212,N_10759,N_10362);
and U11213 (N_11213,N_10269,N_10029);
or U11214 (N_11214,N_10314,N_10786);
and U11215 (N_11215,N_10160,N_10891);
or U11216 (N_11216,N_10368,N_10899);
and U11217 (N_11217,N_10422,N_10294);
and U11218 (N_11218,N_10725,N_10606);
xnor U11219 (N_11219,N_10841,N_10197);
nor U11220 (N_11220,N_10032,N_10709);
xor U11221 (N_11221,N_10999,N_10811);
and U11222 (N_11222,N_10384,N_10537);
nand U11223 (N_11223,N_10107,N_10821);
xnor U11224 (N_11224,N_10145,N_10303);
nor U11225 (N_11225,N_10426,N_10360);
or U11226 (N_11226,N_10834,N_10483);
xor U11227 (N_11227,N_10366,N_10093);
nor U11228 (N_11228,N_10789,N_10733);
or U11229 (N_11229,N_10438,N_10328);
nand U11230 (N_11230,N_10010,N_10230);
and U11231 (N_11231,N_10279,N_10452);
nor U11232 (N_11232,N_10141,N_10954);
or U11233 (N_11233,N_10617,N_10099);
xnor U11234 (N_11234,N_10079,N_10055);
nor U11235 (N_11235,N_10315,N_10996);
or U11236 (N_11236,N_10872,N_10867);
xor U11237 (N_11237,N_10321,N_10014);
xor U11238 (N_11238,N_10987,N_10223);
nand U11239 (N_11239,N_10830,N_10247);
nor U11240 (N_11240,N_10397,N_10381);
xor U11241 (N_11241,N_10621,N_10556);
and U11242 (N_11242,N_10465,N_10731);
xnor U11243 (N_11243,N_10678,N_10563);
or U11244 (N_11244,N_10619,N_10664);
and U11245 (N_11245,N_10754,N_10737);
xor U11246 (N_11246,N_10382,N_10289);
xnor U11247 (N_11247,N_10975,N_10401);
nor U11248 (N_11248,N_10877,N_10824);
xor U11249 (N_11249,N_10504,N_10772);
nand U11250 (N_11250,N_10938,N_10752);
xor U11251 (N_11251,N_10940,N_10154);
or U11252 (N_11252,N_10615,N_10660);
xnor U11253 (N_11253,N_10372,N_10903);
xnor U11254 (N_11254,N_10749,N_10275);
nor U11255 (N_11255,N_10897,N_10740);
or U11256 (N_11256,N_10435,N_10713);
or U11257 (N_11257,N_10496,N_10351);
or U11258 (N_11258,N_10431,N_10202);
nand U11259 (N_11259,N_10937,N_10911);
nand U11260 (N_11260,N_10380,N_10573);
or U11261 (N_11261,N_10458,N_10229);
xnor U11262 (N_11262,N_10089,N_10213);
xnor U11263 (N_11263,N_10979,N_10819);
or U11264 (N_11264,N_10252,N_10681);
or U11265 (N_11265,N_10150,N_10060);
nor U11266 (N_11266,N_10644,N_10511);
nor U11267 (N_11267,N_10348,N_10787);
xnor U11268 (N_11268,N_10735,N_10596);
nand U11269 (N_11269,N_10263,N_10905);
nand U11270 (N_11270,N_10441,N_10030);
nand U11271 (N_11271,N_10117,N_10190);
nand U11272 (N_11272,N_10091,N_10234);
or U11273 (N_11273,N_10712,N_10174);
xnor U11274 (N_11274,N_10476,N_10377);
or U11275 (N_11275,N_10842,N_10895);
or U11276 (N_11276,N_10347,N_10751);
nor U11277 (N_11277,N_10494,N_10090);
nor U11278 (N_11278,N_10440,N_10267);
and U11279 (N_11279,N_10852,N_10567);
nand U11280 (N_11280,N_10920,N_10075);
nand U11281 (N_11281,N_10085,N_10255);
xor U11282 (N_11282,N_10750,N_10796);
or U11283 (N_11283,N_10935,N_10961);
and U11284 (N_11284,N_10592,N_10176);
nor U11285 (N_11285,N_10495,N_10715);
xor U11286 (N_11286,N_10370,N_10290);
nand U11287 (N_11287,N_10363,N_10146);
xnor U11288 (N_11288,N_10767,N_10499);
and U11289 (N_11289,N_10437,N_10736);
or U11290 (N_11290,N_10860,N_10945);
nand U11291 (N_11291,N_10983,N_10837);
nand U11292 (N_11292,N_10219,N_10817);
nor U11293 (N_11293,N_10293,N_10501);
nand U11294 (N_11294,N_10788,N_10486);
xnor U11295 (N_11295,N_10730,N_10395);
nor U11296 (N_11296,N_10064,N_10894);
or U11297 (N_11297,N_10746,N_10711);
xnor U11298 (N_11298,N_10534,N_10322);
or U11299 (N_11299,N_10801,N_10766);
nand U11300 (N_11300,N_10863,N_10272);
nor U11301 (N_11301,N_10602,N_10614);
and U11302 (N_11302,N_10577,N_10295);
xor U11303 (N_11303,N_10874,N_10148);
xnor U11304 (N_11304,N_10344,N_10482);
or U11305 (N_11305,N_10955,N_10726);
nor U11306 (N_11306,N_10392,N_10284);
nand U11307 (N_11307,N_10704,N_10641);
and U11308 (N_11308,N_10019,N_10628);
or U11309 (N_11309,N_10818,N_10244);
or U11310 (N_11310,N_10336,N_10339);
or U11311 (N_11311,N_10635,N_10288);
xnor U11312 (N_11312,N_10402,N_10637);
or U11313 (N_11313,N_10033,N_10638);
xnor U11314 (N_11314,N_10192,N_10623);
and U11315 (N_11315,N_10972,N_10260);
or U11316 (N_11316,N_10172,N_10268);
or U11317 (N_11317,N_10383,N_10274);
nand U11318 (N_11318,N_10584,N_10743);
or U11319 (N_11319,N_10976,N_10588);
xor U11320 (N_11320,N_10661,N_10960);
xnor U11321 (N_11321,N_10741,N_10113);
and U11322 (N_11322,N_10941,N_10428);
nor U11323 (N_11323,N_10981,N_10957);
nor U11324 (N_11324,N_10547,N_10400);
xor U11325 (N_11325,N_10011,N_10990);
and U11326 (N_11326,N_10861,N_10607);
or U11327 (N_11327,N_10035,N_10188);
nor U11328 (N_11328,N_10408,N_10012);
nand U11329 (N_11329,N_10771,N_10067);
and U11330 (N_11330,N_10078,N_10939);
nand U11331 (N_11331,N_10722,N_10902);
xnor U11332 (N_11332,N_10179,N_10676);
nor U11333 (N_11333,N_10186,N_10848);
nand U11334 (N_11334,N_10181,N_10210);
and U11335 (N_11335,N_10265,N_10970);
and U11336 (N_11336,N_10535,N_10345);
or U11337 (N_11337,N_10305,N_10783);
and U11338 (N_11338,N_10785,N_10773);
xor U11339 (N_11339,N_10850,N_10718);
or U11340 (N_11340,N_10307,N_10009);
nor U11341 (N_11341,N_10412,N_10933);
and U11342 (N_11342,N_10913,N_10049);
xor U11343 (N_11343,N_10703,N_10108);
or U11344 (N_11344,N_10246,N_10597);
nand U11345 (N_11345,N_10058,N_10807);
and U11346 (N_11346,N_10102,N_10721);
xnor U11347 (N_11347,N_10545,N_10118);
nor U11348 (N_11348,N_10708,N_10583);
xor U11349 (N_11349,N_10105,N_10524);
nor U11350 (N_11350,N_10024,N_10256);
xnor U11351 (N_11351,N_10748,N_10066);
nand U11352 (N_11352,N_10248,N_10670);
nand U11353 (N_11353,N_10856,N_10995);
xnor U11354 (N_11354,N_10498,N_10946);
nand U11355 (N_11355,N_10353,N_10082);
or U11356 (N_11356,N_10539,N_10890);
xnor U11357 (N_11357,N_10469,N_10059);
xor U11358 (N_11358,N_10135,N_10308);
or U11359 (N_11359,N_10591,N_10727);
xor U11360 (N_11360,N_10851,N_10405);
nand U11361 (N_11361,N_10151,N_10413);
nand U11362 (N_11362,N_10170,N_10098);
nand U11363 (N_11363,N_10448,N_10559);
xnor U11364 (N_11364,N_10450,N_10069);
and U11365 (N_11365,N_10930,N_10350);
nand U11366 (N_11366,N_10466,N_10144);
and U11367 (N_11367,N_10183,N_10969);
nor U11368 (N_11368,N_10297,N_10061);
nor U11369 (N_11369,N_10612,N_10633);
or U11370 (N_11370,N_10207,N_10106);
or U11371 (N_11371,N_10527,N_10447);
xnor U11372 (N_11372,N_10257,N_10519);
and U11373 (N_11373,N_10358,N_10092);
xor U11374 (N_11374,N_10764,N_10543);
and U11375 (N_11375,N_10433,N_10544);
xnor U11376 (N_11376,N_10152,N_10041);
nor U11377 (N_11377,N_10120,N_10875);
nor U11378 (N_11378,N_10330,N_10334);
xnor U11379 (N_11379,N_10964,N_10942);
nand U11380 (N_11380,N_10761,N_10379);
or U11381 (N_11381,N_10453,N_10910);
or U11382 (N_11382,N_10388,N_10237);
nand U11383 (N_11383,N_10245,N_10515);
or U11384 (N_11384,N_10797,N_10331);
nor U11385 (N_11385,N_10003,N_10369);
and U11386 (N_11386,N_10403,N_10616);
nor U11387 (N_11387,N_10728,N_10488);
nor U11388 (N_11388,N_10657,N_10443);
and U11389 (N_11389,N_10128,N_10415);
and U11390 (N_11390,N_10984,N_10484);
xnor U11391 (N_11391,N_10838,N_10341);
and U11392 (N_11392,N_10809,N_10927);
nand U11393 (N_11393,N_10716,N_10864);
or U11394 (N_11394,N_10887,N_10005);
nand U11395 (N_11395,N_10167,N_10698);
xnor U11396 (N_11396,N_10816,N_10201);
or U11397 (N_11397,N_10318,N_10087);
xor U11398 (N_11398,N_10053,N_10166);
and U11399 (N_11399,N_10467,N_10050);
and U11400 (N_11400,N_10521,N_10667);
or U11401 (N_11401,N_10575,N_10399);
nand U11402 (N_11402,N_10980,N_10808);
and U11403 (N_11403,N_10080,N_10451);
or U11404 (N_11404,N_10278,N_10022);
nor U11405 (N_11405,N_10164,N_10594);
nand U11406 (N_11406,N_10038,N_10522);
xnor U11407 (N_11407,N_10138,N_10689);
nand U11408 (N_11408,N_10675,N_10455);
nor U11409 (N_11409,N_10163,N_10407);
and U11410 (N_11410,N_10849,N_10959);
xnor U11411 (N_11411,N_10463,N_10540);
xnor U11412 (N_11412,N_10695,N_10500);
nor U11413 (N_11413,N_10610,N_10706);
or U11414 (N_11414,N_10908,N_10302);
xnor U11415 (N_11415,N_10734,N_10884);
nor U11416 (N_11416,N_10324,N_10944);
nor U11417 (N_11417,N_10613,N_10432);
nor U11418 (N_11418,N_10506,N_10753);
nand U11419 (N_11419,N_10674,N_10023);
nand U11420 (N_11420,N_10131,N_10642);
or U11421 (N_11421,N_10699,N_10300);
nor U11422 (N_11422,N_10000,N_10357);
xnor U11423 (N_11423,N_10094,N_10780);
or U11424 (N_11424,N_10497,N_10757);
and U11425 (N_11425,N_10845,N_10291);
and U11426 (N_11426,N_10794,N_10601);
xor U11427 (N_11427,N_10934,N_10719);
nor U11428 (N_11428,N_10393,N_10870);
xnor U11429 (N_11429,N_10662,N_10994);
or U11430 (N_11430,N_10691,N_10578);
xor U11431 (N_11431,N_10840,N_10700);
and U11432 (N_11432,N_10907,N_10214);
nor U11433 (N_11433,N_10777,N_10855);
and U11434 (N_11434,N_10273,N_10724);
xor U11435 (N_11435,N_10016,N_10349);
nor U11436 (N_11436,N_10778,N_10857);
nor U11437 (N_11437,N_10367,N_10508);
and U11438 (N_11438,N_10952,N_10462);
xor U11439 (N_11439,N_10992,N_10299);
or U11440 (N_11440,N_10235,N_10943);
and U11441 (N_11441,N_10046,N_10538);
or U11442 (N_11442,N_10549,N_10215);
or U11443 (N_11443,N_10512,N_10419);
or U11444 (N_11444,N_10459,N_10184);
xnor U11445 (N_11445,N_10629,N_10799);
or U11446 (N_11446,N_10507,N_10409);
and U11447 (N_11447,N_10203,N_10820);
nand U11448 (N_11448,N_10218,N_10859);
xnor U11449 (N_11449,N_10765,N_10823);
xnor U11450 (N_11450,N_10919,N_10354);
or U11451 (N_11451,N_10739,N_10669);
nand U11452 (N_11452,N_10084,N_10477);
nor U11453 (N_11453,N_10346,N_10793);
xnor U11454 (N_11454,N_10881,N_10139);
nor U11455 (N_11455,N_10822,N_10680);
and U11456 (N_11456,N_10101,N_10646);
or U11457 (N_11457,N_10039,N_10124);
or U11458 (N_11458,N_10516,N_10974);
nor U11459 (N_11459,N_10971,N_10045);
or U11460 (N_11460,N_10134,N_10586);
or U11461 (N_11461,N_10880,N_10200);
and U11462 (N_11462,N_10835,N_10473);
nand U11463 (N_11463,N_10096,N_10658);
xor U11464 (N_11464,N_10309,N_10679);
nand U11465 (N_11465,N_10893,N_10865);
xor U11466 (N_11466,N_10301,N_10168);
nor U11467 (N_11467,N_10057,N_10677);
and U11468 (N_11468,N_10031,N_10985);
xor U11469 (N_11469,N_10925,N_10569);
xnor U11470 (N_11470,N_10385,N_10928);
nand U11471 (N_11471,N_10424,N_10337);
nand U11472 (N_11472,N_10572,N_10071);
nor U11473 (N_11473,N_10007,N_10157);
nor U11474 (N_11474,N_10364,N_10546);
xnor U11475 (N_11475,N_10696,N_10774);
xnor U11476 (N_11476,N_10915,N_10526);
xnor U11477 (N_11477,N_10316,N_10829);
nor U11478 (N_11478,N_10258,N_10846);
and U11479 (N_11479,N_10088,N_10277);
and U11480 (N_11480,N_10795,N_10705);
or U11481 (N_11481,N_10530,N_10707);
and U11482 (N_11482,N_10769,N_10520);
or U11483 (N_11483,N_10673,N_10682);
or U11484 (N_11484,N_10198,N_10986);
or U11485 (N_11485,N_10968,N_10311);
nor U11486 (N_11486,N_10966,N_10929);
or U11487 (N_11487,N_10525,N_10216);
nor U11488 (N_11488,N_10343,N_10523);
xor U11489 (N_11489,N_10869,N_10528);
xor U11490 (N_11490,N_10883,N_10253);
and U11491 (N_11491,N_10047,N_10359);
xor U11492 (N_11492,N_10914,N_10241);
nand U11493 (N_11493,N_10130,N_10701);
nand U11494 (N_11494,N_10063,N_10136);
or U11495 (N_11495,N_10826,N_10460);
or U11496 (N_11496,N_10194,N_10997);
nor U11497 (N_11497,N_10421,N_10532);
xor U11498 (N_11498,N_10647,N_10140);
and U11499 (N_11499,N_10225,N_10182);
or U11500 (N_11500,N_10963,N_10269);
nor U11501 (N_11501,N_10193,N_10058);
xor U11502 (N_11502,N_10087,N_10239);
xor U11503 (N_11503,N_10044,N_10922);
xor U11504 (N_11504,N_10008,N_10074);
nor U11505 (N_11505,N_10095,N_10646);
xnor U11506 (N_11506,N_10921,N_10452);
xor U11507 (N_11507,N_10354,N_10435);
xnor U11508 (N_11508,N_10048,N_10255);
xor U11509 (N_11509,N_10234,N_10073);
and U11510 (N_11510,N_10287,N_10791);
and U11511 (N_11511,N_10772,N_10982);
nand U11512 (N_11512,N_10994,N_10324);
and U11513 (N_11513,N_10297,N_10608);
or U11514 (N_11514,N_10887,N_10612);
and U11515 (N_11515,N_10324,N_10625);
and U11516 (N_11516,N_10593,N_10290);
or U11517 (N_11517,N_10394,N_10278);
and U11518 (N_11518,N_10657,N_10468);
or U11519 (N_11519,N_10825,N_10248);
and U11520 (N_11520,N_10378,N_10258);
xor U11521 (N_11521,N_10309,N_10887);
nor U11522 (N_11522,N_10594,N_10970);
nand U11523 (N_11523,N_10043,N_10641);
and U11524 (N_11524,N_10206,N_10411);
or U11525 (N_11525,N_10220,N_10072);
nand U11526 (N_11526,N_10793,N_10418);
xnor U11527 (N_11527,N_10387,N_10266);
xnor U11528 (N_11528,N_10074,N_10322);
or U11529 (N_11529,N_10836,N_10934);
and U11530 (N_11530,N_10601,N_10818);
and U11531 (N_11531,N_10856,N_10313);
and U11532 (N_11532,N_10049,N_10842);
nor U11533 (N_11533,N_10489,N_10770);
or U11534 (N_11534,N_10277,N_10772);
xor U11535 (N_11535,N_10952,N_10097);
nand U11536 (N_11536,N_10926,N_10936);
and U11537 (N_11537,N_10222,N_10683);
and U11538 (N_11538,N_10617,N_10549);
nor U11539 (N_11539,N_10337,N_10989);
nand U11540 (N_11540,N_10526,N_10724);
xor U11541 (N_11541,N_10072,N_10067);
nor U11542 (N_11542,N_10472,N_10529);
xor U11543 (N_11543,N_10691,N_10007);
and U11544 (N_11544,N_10862,N_10104);
and U11545 (N_11545,N_10953,N_10738);
nor U11546 (N_11546,N_10200,N_10631);
or U11547 (N_11547,N_10844,N_10479);
or U11548 (N_11548,N_10699,N_10599);
or U11549 (N_11549,N_10447,N_10645);
nand U11550 (N_11550,N_10704,N_10814);
nor U11551 (N_11551,N_10000,N_10668);
and U11552 (N_11552,N_10578,N_10385);
and U11553 (N_11553,N_10512,N_10043);
nand U11554 (N_11554,N_10841,N_10546);
or U11555 (N_11555,N_10838,N_10902);
and U11556 (N_11556,N_10240,N_10843);
or U11557 (N_11557,N_10556,N_10341);
nand U11558 (N_11558,N_10449,N_10232);
nand U11559 (N_11559,N_10048,N_10074);
xnor U11560 (N_11560,N_10316,N_10211);
and U11561 (N_11561,N_10711,N_10695);
nand U11562 (N_11562,N_10948,N_10590);
xnor U11563 (N_11563,N_10051,N_10469);
and U11564 (N_11564,N_10458,N_10362);
or U11565 (N_11565,N_10604,N_10331);
nor U11566 (N_11566,N_10254,N_10266);
or U11567 (N_11567,N_10865,N_10609);
xor U11568 (N_11568,N_10591,N_10870);
or U11569 (N_11569,N_10707,N_10071);
and U11570 (N_11570,N_10803,N_10986);
xor U11571 (N_11571,N_10783,N_10759);
and U11572 (N_11572,N_10707,N_10856);
or U11573 (N_11573,N_10936,N_10387);
and U11574 (N_11574,N_10981,N_10403);
nand U11575 (N_11575,N_10226,N_10416);
and U11576 (N_11576,N_10567,N_10856);
and U11577 (N_11577,N_10337,N_10812);
and U11578 (N_11578,N_10279,N_10491);
nand U11579 (N_11579,N_10172,N_10185);
nor U11580 (N_11580,N_10408,N_10010);
and U11581 (N_11581,N_10896,N_10813);
nor U11582 (N_11582,N_10981,N_10724);
and U11583 (N_11583,N_10893,N_10569);
and U11584 (N_11584,N_10552,N_10821);
nand U11585 (N_11585,N_10258,N_10362);
and U11586 (N_11586,N_10241,N_10593);
xnor U11587 (N_11587,N_10498,N_10214);
nor U11588 (N_11588,N_10582,N_10560);
or U11589 (N_11589,N_10640,N_10469);
or U11590 (N_11590,N_10275,N_10911);
or U11591 (N_11591,N_10414,N_10737);
and U11592 (N_11592,N_10583,N_10007);
nand U11593 (N_11593,N_10600,N_10745);
nor U11594 (N_11594,N_10500,N_10549);
nand U11595 (N_11595,N_10423,N_10205);
and U11596 (N_11596,N_10079,N_10573);
nand U11597 (N_11597,N_10861,N_10481);
nand U11598 (N_11598,N_10652,N_10366);
nand U11599 (N_11599,N_10511,N_10290);
xor U11600 (N_11600,N_10683,N_10953);
nand U11601 (N_11601,N_10684,N_10566);
and U11602 (N_11602,N_10591,N_10372);
nand U11603 (N_11603,N_10765,N_10829);
xor U11604 (N_11604,N_10548,N_10797);
and U11605 (N_11605,N_10253,N_10811);
xor U11606 (N_11606,N_10925,N_10071);
and U11607 (N_11607,N_10520,N_10464);
or U11608 (N_11608,N_10491,N_10081);
or U11609 (N_11609,N_10000,N_10312);
nand U11610 (N_11610,N_10749,N_10311);
or U11611 (N_11611,N_10050,N_10763);
xnor U11612 (N_11612,N_10715,N_10520);
and U11613 (N_11613,N_10645,N_10349);
or U11614 (N_11614,N_10273,N_10636);
nor U11615 (N_11615,N_10850,N_10149);
nand U11616 (N_11616,N_10146,N_10654);
or U11617 (N_11617,N_10925,N_10305);
xor U11618 (N_11618,N_10125,N_10747);
nand U11619 (N_11619,N_10355,N_10881);
xor U11620 (N_11620,N_10363,N_10465);
nor U11621 (N_11621,N_10382,N_10242);
nand U11622 (N_11622,N_10864,N_10785);
or U11623 (N_11623,N_10693,N_10960);
or U11624 (N_11624,N_10338,N_10381);
and U11625 (N_11625,N_10593,N_10109);
or U11626 (N_11626,N_10002,N_10992);
nor U11627 (N_11627,N_10082,N_10209);
and U11628 (N_11628,N_10369,N_10732);
nor U11629 (N_11629,N_10473,N_10735);
or U11630 (N_11630,N_10855,N_10652);
nor U11631 (N_11631,N_10789,N_10251);
xor U11632 (N_11632,N_10376,N_10718);
nand U11633 (N_11633,N_10519,N_10544);
and U11634 (N_11634,N_10989,N_10295);
or U11635 (N_11635,N_10539,N_10248);
nand U11636 (N_11636,N_10857,N_10995);
or U11637 (N_11637,N_10708,N_10640);
nor U11638 (N_11638,N_10906,N_10943);
nor U11639 (N_11639,N_10707,N_10130);
and U11640 (N_11640,N_10255,N_10532);
nor U11641 (N_11641,N_10904,N_10133);
nand U11642 (N_11642,N_10347,N_10638);
and U11643 (N_11643,N_10616,N_10291);
xnor U11644 (N_11644,N_10220,N_10955);
and U11645 (N_11645,N_10015,N_10307);
nor U11646 (N_11646,N_10296,N_10789);
xnor U11647 (N_11647,N_10847,N_10883);
xnor U11648 (N_11648,N_10086,N_10295);
and U11649 (N_11649,N_10326,N_10835);
nand U11650 (N_11650,N_10242,N_10082);
xnor U11651 (N_11651,N_10165,N_10683);
or U11652 (N_11652,N_10892,N_10574);
nor U11653 (N_11653,N_10691,N_10113);
nor U11654 (N_11654,N_10146,N_10818);
nor U11655 (N_11655,N_10883,N_10141);
nand U11656 (N_11656,N_10818,N_10853);
or U11657 (N_11657,N_10466,N_10853);
or U11658 (N_11658,N_10100,N_10973);
or U11659 (N_11659,N_10375,N_10306);
or U11660 (N_11660,N_10302,N_10030);
xor U11661 (N_11661,N_10592,N_10849);
nor U11662 (N_11662,N_10448,N_10895);
and U11663 (N_11663,N_10455,N_10178);
and U11664 (N_11664,N_10810,N_10481);
and U11665 (N_11665,N_10047,N_10277);
nand U11666 (N_11666,N_10030,N_10040);
nand U11667 (N_11667,N_10554,N_10865);
xnor U11668 (N_11668,N_10316,N_10062);
nor U11669 (N_11669,N_10424,N_10922);
or U11670 (N_11670,N_10847,N_10619);
or U11671 (N_11671,N_10695,N_10879);
nor U11672 (N_11672,N_10558,N_10504);
nor U11673 (N_11673,N_10545,N_10168);
and U11674 (N_11674,N_10120,N_10699);
or U11675 (N_11675,N_10085,N_10266);
or U11676 (N_11676,N_10783,N_10573);
nand U11677 (N_11677,N_10283,N_10831);
xnor U11678 (N_11678,N_10504,N_10551);
nand U11679 (N_11679,N_10523,N_10165);
and U11680 (N_11680,N_10962,N_10934);
or U11681 (N_11681,N_10599,N_10697);
nand U11682 (N_11682,N_10608,N_10968);
nand U11683 (N_11683,N_10364,N_10970);
and U11684 (N_11684,N_10278,N_10776);
nand U11685 (N_11685,N_10099,N_10656);
and U11686 (N_11686,N_10293,N_10103);
or U11687 (N_11687,N_10777,N_10736);
nand U11688 (N_11688,N_10679,N_10864);
nand U11689 (N_11689,N_10421,N_10023);
nand U11690 (N_11690,N_10059,N_10333);
and U11691 (N_11691,N_10374,N_10963);
nor U11692 (N_11692,N_10503,N_10589);
xor U11693 (N_11693,N_10667,N_10464);
xor U11694 (N_11694,N_10080,N_10550);
or U11695 (N_11695,N_10539,N_10183);
or U11696 (N_11696,N_10435,N_10756);
and U11697 (N_11697,N_10931,N_10402);
nand U11698 (N_11698,N_10639,N_10936);
xor U11699 (N_11699,N_10401,N_10942);
nor U11700 (N_11700,N_10534,N_10684);
nand U11701 (N_11701,N_10139,N_10634);
or U11702 (N_11702,N_10125,N_10716);
xnor U11703 (N_11703,N_10863,N_10797);
nor U11704 (N_11704,N_10205,N_10567);
xnor U11705 (N_11705,N_10951,N_10774);
nor U11706 (N_11706,N_10385,N_10848);
xnor U11707 (N_11707,N_10235,N_10230);
or U11708 (N_11708,N_10358,N_10127);
xor U11709 (N_11709,N_10713,N_10182);
or U11710 (N_11710,N_10687,N_10434);
nand U11711 (N_11711,N_10204,N_10554);
nand U11712 (N_11712,N_10620,N_10315);
xnor U11713 (N_11713,N_10735,N_10528);
xor U11714 (N_11714,N_10015,N_10615);
xor U11715 (N_11715,N_10109,N_10348);
nand U11716 (N_11716,N_10255,N_10177);
or U11717 (N_11717,N_10932,N_10747);
and U11718 (N_11718,N_10022,N_10158);
and U11719 (N_11719,N_10816,N_10107);
nand U11720 (N_11720,N_10393,N_10324);
and U11721 (N_11721,N_10417,N_10109);
nand U11722 (N_11722,N_10659,N_10640);
nand U11723 (N_11723,N_10733,N_10925);
and U11724 (N_11724,N_10729,N_10305);
nand U11725 (N_11725,N_10793,N_10184);
or U11726 (N_11726,N_10387,N_10174);
and U11727 (N_11727,N_10113,N_10800);
nand U11728 (N_11728,N_10046,N_10741);
nand U11729 (N_11729,N_10902,N_10776);
xor U11730 (N_11730,N_10049,N_10480);
or U11731 (N_11731,N_10089,N_10818);
nand U11732 (N_11732,N_10591,N_10988);
xnor U11733 (N_11733,N_10735,N_10322);
and U11734 (N_11734,N_10714,N_10582);
nand U11735 (N_11735,N_10813,N_10945);
nor U11736 (N_11736,N_10431,N_10257);
or U11737 (N_11737,N_10163,N_10057);
and U11738 (N_11738,N_10708,N_10560);
and U11739 (N_11739,N_10859,N_10865);
and U11740 (N_11740,N_10409,N_10954);
xor U11741 (N_11741,N_10963,N_10144);
xnor U11742 (N_11742,N_10731,N_10140);
xor U11743 (N_11743,N_10940,N_10386);
nand U11744 (N_11744,N_10774,N_10173);
or U11745 (N_11745,N_10519,N_10091);
or U11746 (N_11746,N_10640,N_10897);
nand U11747 (N_11747,N_10423,N_10866);
nor U11748 (N_11748,N_10287,N_10877);
or U11749 (N_11749,N_10291,N_10147);
and U11750 (N_11750,N_10423,N_10883);
nor U11751 (N_11751,N_10652,N_10064);
or U11752 (N_11752,N_10557,N_10066);
xor U11753 (N_11753,N_10798,N_10009);
and U11754 (N_11754,N_10746,N_10090);
and U11755 (N_11755,N_10497,N_10598);
or U11756 (N_11756,N_10706,N_10372);
nand U11757 (N_11757,N_10543,N_10097);
xor U11758 (N_11758,N_10012,N_10837);
xor U11759 (N_11759,N_10702,N_10524);
and U11760 (N_11760,N_10244,N_10658);
xnor U11761 (N_11761,N_10599,N_10047);
and U11762 (N_11762,N_10155,N_10289);
nor U11763 (N_11763,N_10114,N_10529);
nand U11764 (N_11764,N_10436,N_10760);
xnor U11765 (N_11765,N_10956,N_10733);
or U11766 (N_11766,N_10330,N_10737);
nand U11767 (N_11767,N_10437,N_10408);
and U11768 (N_11768,N_10969,N_10461);
or U11769 (N_11769,N_10007,N_10751);
nand U11770 (N_11770,N_10754,N_10514);
nor U11771 (N_11771,N_10793,N_10799);
xor U11772 (N_11772,N_10841,N_10422);
and U11773 (N_11773,N_10154,N_10493);
or U11774 (N_11774,N_10239,N_10317);
nor U11775 (N_11775,N_10767,N_10746);
or U11776 (N_11776,N_10738,N_10022);
xnor U11777 (N_11777,N_10919,N_10620);
xnor U11778 (N_11778,N_10662,N_10926);
nand U11779 (N_11779,N_10380,N_10040);
or U11780 (N_11780,N_10140,N_10928);
nor U11781 (N_11781,N_10111,N_10223);
or U11782 (N_11782,N_10906,N_10890);
xnor U11783 (N_11783,N_10604,N_10967);
nand U11784 (N_11784,N_10037,N_10591);
or U11785 (N_11785,N_10644,N_10474);
or U11786 (N_11786,N_10984,N_10610);
or U11787 (N_11787,N_10514,N_10624);
and U11788 (N_11788,N_10521,N_10134);
nand U11789 (N_11789,N_10426,N_10788);
nand U11790 (N_11790,N_10488,N_10224);
or U11791 (N_11791,N_10906,N_10206);
nor U11792 (N_11792,N_10039,N_10163);
nor U11793 (N_11793,N_10295,N_10453);
or U11794 (N_11794,N_10099,N_10486);
nand U11795 (N_11795,N_10582,N_10743);
nor U11796 (N_11796,N_10723,N_10342);
nand U11797 (N_11797,N_10287,N_10095);
xnor U11798 (N_11798,N_10680,N_10633);
nor U11799 (N_11799,N_10252,N_10762);
and U11800 (N_11800,N_10548,N_10521);
xnor U11801 (N_11801,N_10545,N_10638);
and U11802 (N_11802,N_10029,N_10823);
nand U11803 (N_11803,N_10216,N_10226);
or U11804 (N_11804,N_10334,N_10409);
nand U11805 (N_11805,N_10859,N_10470);
and U11806 (N_11806,N_10912,N_10506);
nand U11807 (N_11807,N_10542,N_10915);
nor U11808 (N_11808,N_10647,N_10739);
and U11809 (N_11809,N_10629,N_10644);
xnor U11810 (N_11810,N_10561,N_10761);
nand U11811 (N_11811,N_10991,N_10934);
and U11812 (N_11812,N_10007,N_10628);
xor U11813 (N_11813,N_10936,N_10357);
xnor U11814 (N_11814,N_10707,N_10010);
xor U11815 (N_11815,N_10635,N_10764);
or U11816 (N_11816,N_10813,N_10500);
xnor U11817 (N_11817,N_10392,N_10539);
xor U11818 (N_11818,N_10951,N_10375);
and U11819 (N_11819,N_10019,N_10737);
xor U11820 (N_11820,N_10753,N_10062);
nand U11821 (N_11821,N_10112,N_10409);
nor U11822 (N_11822,N_10273,N_10924);
and U11823 (N_11823,N_10027,N_10298);
and U11824 (N_11824,N_10980,N_10109);
xor U11825 (N_11825,N_10543,N_10713);
nor U11826 (N_11826,N_10618,N_10123);
nand U11827 (N_11827,N_10930,N_10809);
xnor U11828 (N_11828,N_10109,N_10397);
or U11829 (N_11829,N_10554,N_10777);
xor U11830 (N_11830,N_10618,N_10289);
or U11831 (N_11831,N_10172,N_10769);
and U11832 (N_11832,N_10288,N_10904);
and U11833 (N_11833,N_10868,N_10063);
nor U11834 (N_11834,N_10917,N_10312);
and U11835 (N_11835,N_10036,N_10120);
xor U11836 (N_11836,N_10647,N_10127);
nor U11837 (N_11837,N_10420,N_10386);
or U11838 (N_11838,N_10641,N_10764);
nor U11839 (N_11839,N_10967,N_10606);
xnor U11840 (N_11840,N_10828,N_10558);
xor U11841 (N_11841,N_10817,N_10928);
and U11842 (N_11842,N_10228,N_10337);
xnor U11843 (N_11843,N_10841,N_10272);
nand U11844 (N_11844,N_10351,N_10871);
xor U11845 (N_11845,N_10377,N_10820);
nand U11846 (N_11846,N_10171,N_10393);
nand U11847 (N_11847,N_10037,N_10760);
and U11848 (N_11848,N_10553,N_10396);
xnor U11849 (N_11849,N_10692,N_10094);
xnor U11850 (N_11850,N_10883,N_10344);
and U11851 (N_11851,N_10230,N_10270);
nor U11852 (N_11852,N_10590,N_10230);
or U11853 (N_11853,N_10593,N_10160);
nor U11854 (N_11854,N_10031,N_10744);
nor U11855 (N_11855,N_10372,N_10683);
nand U11856 (N_11856,N_10804,N_10287);
nand U11857 (N_11857,N_10069,N_10140);
and U11858 (N_11858,N_10170,N_10002);
and U11859 (N_11859,N_10455,N_10690);
nand U11860 (N_11860,N_10628,N_10753);
nand U11861 (N_11861,N_10292,N_10274);
xor U11862 (N_11862,N_10650,N_10948);
or U11863 (N_11863,N_10768,N_10972);
nor U11864 (N_11864,N_10558,N_10220);
or U11865 (N_11865,N_10834,N_10602);
and U11866 (N_11866,N_10453,N_10385);
xor U11867 (N_11867,N_10403,N_10024);
or U11868 (N_11868,N_10872,N_10723);
xor U11869 (N_11869,N_10415,N_10478);
xnor U11870 (N_11870,N_10521,N_10596);
or U11871 (N_11871,N_10953,N_10190);
nor U11872 (N_11872,N_10998,N_10493);
nand U11873 (N_11873,N_10503,N_10816);
nor U11874 (N_11874,N_10588,N_10383);
xor U11875 (N_11875,N_10981,N_10907);
and U11876 (N_11876,N_10474,N_10376);
nor U11877 (N_11877,N_10459,N_10007);
nor U11878 (N_11878,N_10753,N_10235);
nand U11879 (N_11879,N_10646,N_10803);
and U11880 (N_11880,N_10974,N_10730);
and U11881 (N_11881,N_10025,N_10783);
or U11882 (N_11882,N_10894,N_10116);
xor U11883 (N_11883,N_10015,N_10258);
nand U11884 (N_11884,N_10011,N_10629);
nand U11885 (N_11885,N_10731,N_10455);
nor U11886 (N_11886,N_10553,N_10404);
nor U11887 (N_11887,N_10991,N_10940);
nor U11888 (N_11888,N_10747,N_10230);
nor U11889 (N_11889,N_10072,N_10603);
or U11890 (N_11890,N_10370,N_10690);
or U11891 (N_11891,N_10108,N_10902);
xor U11892 (N_11892,N_10690,N_10567);
xnor U11893 (N_11893,N_10613,N_10361);
nor U11894 (N_11894,N_10354,N_10013);
or U11895 (N_11895,N_10772,N_10335);
and U11896 (N_11896,N_10085,N_10689);
xnor U11897 (N_11897,N_10377,N_10037);
and U11898 (N_11898,N_10126,N_10732);
and U11899 (N_11899,N_10174,N_10541);
nor U11900 (N_11900,N_10477,N_10258);
nand U11901 (N_11901,N_10148,N_10318);
xor U11902 (N_11902,N_10419,N_10455);
or U11903 (N_11903,N_10503,N_10555);
or U11904 (N_11904,N_10378,N_10084);
nand U11905 (N_11905,N_10602,N_10781);
xnor U11906 (N_11906,N_10326,N_10380);
and U11907 (N_11907,N_10311,N_10089);
xor U11908 (N_11908,N_10919,N_10655);
or U11909 (N_11909,N_10640,N_10072);
nand U11910 (N_11910,N_10109,N_10440);
nand U11911 (N_11911,N_10394,N_10943);
nor U11912 (N_11912,N_10021,N_10588);
or U11913 (N_11913,N_10090,N_10172);
and U11914 (N_11914,N_10733,N_10682);
nor U11915 (N_11915,N_10394,N_10674);
and U11916 (N_11916,N_10923,N_10745);
nand U11917 (N_11917,N_10711,N_10053);
nor U11918 (N_11918,N_10712,N_10861);
and U11919 (N_11919,N_10357,N_10836);
or U11920 (N_11920,N_10816,N_10184);
nor U11921 (N_11921,N_10122,N_10854);
and U11922 (N_11922,N_10778,N_10556);
nor U11923 (N_11923,N_10042,N_10501);
or U11924 (N_11924,N_10987,N_10303);
nand U11925 (N_11925,N_10368,N_10535);
nor U11926 (N_11926,N_10601,N_10821);
xor U11927 (N_11927,N_10727,N_10758);
nor U11928 (N_11928,N_10863,N_10598);
nand U11929 (N_11929,N_10692,N_10981);
nand U11930 (N_11930,N_10537,N_10237);
nand U11931 (N_11931,N_10838,N_10878);
xnor U11932 (N_11932,N_10278,N_10740);
or U11933 (N_11933,N_10700,N_10509);
xnor U11934 (N_11934,N_10290,N_10009);
or U11935 (N_11935,N_10671,N_10352);
and U11936 (N_11936,N_10036,N_10214);
xnor U11937 (N_11937,N_10710,N_10816);
nor U11938 (N_11938,N_10866,N_10889);
nand U11939 (N_11939,N_10441,N_10447);
and U11940 (N_11940,N_10717,N_10505);
or U11941 (N_11941,N_10494,N_10467);
nand U11942 (N_11942,N_10812,N_10632);
nor U11943 (N_11943,N_10650,N_10486);
xor U11944 (N_11944,N_10264,N_10296);
and U11945 (N_11945,N_10222,N_10750);
nand U11946 (N_11946,N_10935,N_10821);
or U11947 (N_11947,N_10430,N_10473);
nor U11948 (N_11948,N_10101,N_10119);
nor U11949 (N_11949,N_10185,N_10765);
and U11950 (N_11950,N_10392,N_10167);
xor U11951 (N_11951,N_10512,N_10842);
or U11952 (N_11952,N_10260,N_10785);
nor U11953 (N_11953,N_10632,N_10415);
or U11954 (N_11954,N_10026,N_10208);
nor U11955 (N_11955,N_10903,N_10214);
xnor U11956 (N_11956,N_10708,N_10616);
xnor U11957 (N_11957,N_10669,N_10730);
and U11958 (N_11958,N_10697,N_10570);
xor U11959 (N_11959,N_10138,N_10844);
or U11960 (N_11960,N_10473,N_10050);
or U11961 (N_11961,N_10507,N_10254);
or U11962 (N_11962,N_10355,N_10023);
nand U11963 (N_11963,N_10983,N_10558);
nor U11964 (N_11964,N_10706,N_10602);
or U11965 (N_11965,N_10412,N_10279);
and U11966 (N_11966,N_10356,N_10378);
nand U11967 (N_11967,N_10079,N_10784);
or U11968 (N_11968,N_10037,N_10582);
nand U11969 (N_11969,N_10189,N_10163);
xnor U11970 (N_11970,N_10351,N_10433);
and U11971 (N_11971,N_10823,N_10897);
or U11972 (N_11972,N_10363,N_10060);
or U11973 (N_11973,N_10620,N_10083);
nand U11974 (N_11974,N_10887,N_10392);
nor U11975 (N_11975,N_10697,N_10834);
nor U11976 (N_11976,N_10583,N_10569);
nor U11977 (N_11977,N_10620,N_10038);
xnor U11978 (N_11978,N_10641,N_10378);
nor U11979 (N_11979,N_10827,N_10024);
xnor U11980 (N_11980,N_10661,N_10610);
xor U11981 (N_11981,N_10081,N_10236);
nor U11982 (N_11982,N_10183,N_10308);
xor U11983 (N_11983,N_10075,N_10520);
xor U11984 (N_11984,N_10527,N_10044);
and U11985 (N_11985,N_10077,N_10944);
nand U11986 (N_11986,N_10376,N_10192);
xnor U11987 (N_11987,N_10703,N_10779);
or U11988 (N_11988,N_10482,N_10942);
and U11989 (N_11989,N_10359,N_10078);
nand U11990 (N_11990,N_10371,N_10570);
xnor U11991 (N_11991,N_10545,N_10930);
nor U11992 (N_11992,N_10613,N_10210);
nand U11993 (N_11993,N_10615,N_10674);
nor U11994 (N_11994,N_10584,N_10321);
or U11995 (N_11995,N_10782,N_10826);
nand U11996 (N_11996,N_10314,N_10112);
or U11997 (N_11997,N_10163,N_10326);
and U11998 (N_11998,N_10372,N_10478);
nor U11999 (N_11999,N_10499,N_10045);
or U12000 (N_12000,N_11773,N_11990);
nor U12001 (N_12001,N_11984,N_11770);
nor U12002 (N_12002,N_11896,N_11333);
nor U12003 (N_12003,N_11190,N_11015);
and U12004 (N_12004,N_11911,N_11674);
xnor U12005 (N_12005,N_11640,N_11747);
nand U12006 (N_12006,N_11650,N_11681);
or U12007 (N_12007,N_11698,N_11223);
nand U12008 (N_12008,N_11332,N_11638);
nand U12009 (N_12009,N_11013,N_11185);
nor U12010 (N_12010,N_11504,N_11292);
or U12011 (N_12011,N_11104,N_11056);
nand U12012 (N_12012,N_11878,N_11270);
or U12013 (N_12013,N_11012,N_11246);
nand U12014 (N_12014,N_11094,N_11230);
or U12015 (N_12015,N_11314,N_11168);
and U12016 (N_12016,N_11272,N_11508);
and U12017 (N_12017,N_11520,N_11478);
xnor U12018 (N_12018,N_11622,N_11918);
or U12019 (N_12019,N_11330,N_11566);
nor U12020 (N_12020,N_11473,N_11624);
nor U12021 (N_12021,N_11629,N_11052);
xor U12022 (N_12022,N_11999,N_11714);
or U12023 (N_12023,N_11832,N_11704);
or U12024 (N_12024,N_11291,N_11317);
and U12025 (N_12025,N_11891,N_11528);
or U12026 (N_12026,N_11467,N_11746);
xor U12027 (N_12027,N_11644,N_11919);
or U12028 (N_12028,N_11838,N_11120);
or U12029 (N_12029,N_11290,N_11108);
nor U12030 (N_12030,N_11582,N_11413);
nand U12031 (N_12031,N_11836,N_11772);
and U12032 (N_12032,N_11194,N_11533);
or U12033 (N_12033,N_11002,N_11577);
xor U12034 (N_12034,N_11822,N_11149);
nand U12035 (N_12035,N_11811,N_11204);
and U12036 (N_12036,N_11509,N_11008);
or U12037 (N_12037,N_11670,N_11360);
nor U12038 (N_12038,N_11496,N_11084);
xor U12039 (N_12039,N_11229,N_11461);
nand U12040 (N_12040,N_11396,N_11534);
nor U12041 (N_12041,N_11046,N_11620);
nor U12042 (N_12042,N_11962,N_11655);
xor U12043 (N_12043,N_11584,N_11725);
xor U12044 (N_12044,N_11817,N_11585);
and U12045 (N_12045,N_11265,N_11445);
xnor U12046 (N_12046,N_11551,N_11414);
and U12047 (N_12047,N_11139,N_11831);
nand U12048 (N_12048,N_11182,N_11814);
nor U12049 (N_12049,N_11144,N_11019);
nor U12050 (N_12050,N_11448,N_11180);
nand U12051 (N_12051,N_11479,N_11404);
xor U12052 (N_12052,N_11952,N_11712);
and U12053 (N_12053,N_11973,N_11258);
and U12054 (N_12054,N_11557,N_11549);
nand U12055 (N_12055,N_11524,N_11102);
nor U12056 (N_12056,N_11976,N_11320);
nand U12057 (N_12057,N_11124,N_11932);
or U12058 (N_12058,N_11064,N_11938);
or U12059 (N_12059,N_11819,N_11188);
nor U12060 (N_12060,N_11410,N_11059);
and U12061 (N_12061,N_11697,N_11484);
and U12062 (N_12062,N_11486,N_11334);
nor U12063 (N_12063,N_11529,N_11009);
nor U12064 (N_12064,N_11312,N_11894);
and U12065 (N_12065,N_11022,N_11153);
nand U12066 (N_12066,N_11284,N_11730);
xnor U12067 (N_12067,N_11550,N_11512);
nand U12068 (N_12068,N_11535,N_11239);
xnor U12069 (N_12069,N_11540,N_11489);
nand U12070 (N_12070,N_11800,N_11175);
nor U12071 (N_12071,N_11611,N_11235);
or U12072 (N_12072,N_11379,N_11957);
xnor U12073 (N_12073,N_11845,N_11151);
nand U12074 (N_12074,N_11623,N_11868);
and U12075 (N_12075,N_11498,N_11543);
nand U12076 (N_12076,N_11386,N_11858);
nor U12077 (N_12077,N_11892,N_11327);
nor U12078 (N_12078,N_11606,N_11202);
or U12079 (N_12079,N_11726,N_11179);
or U12080 (N_12080,N_11067,N_11460);
and U12081 (N_12081,N_11925,N_11572);
nor U12082 (N_12082,N_11830,N_11118);
nor U12083 (N_12083,N_11693,N_11308);
and U12084 (N_12084,N_11542,N_11200);
nand U12085 (N_12085,N_11567,N_11574);
nand U12086 (N_12086,N_11942,N_11571);
and U12087 (N_12087,N_11752,N_11370);
nand U12088 (N_12088,N_11329,N_11824);
nand U12089 (N_12089,N_11127,N_11956);
nand U12090 (N_12090,N_11851,N_11782);
nor U12091 (N_12091,N_11017,N_11420);
or U12092 (N_12092,N_11287,N_11384);
or U12093 (N_12093,N_11864,N_11672);
nand U12094 (N_12094,N_11183,N_11625);
nand U12095 (N_12095,N_11676,N_11391);
xnor U12096 (N_12096,N_11684,N_11328);
nand U12097 (N_12097,N_11702,N_11429);
or U12098 (N_12098,N_11117,N_11724);
xor U12099 (N_12099,N_11169,N_11545);
xor U12100 (N_12100,N_11361,N_11283);
or U12101 (N_12101,N_11197,N_11663);
or U12102 (N_12102,N_11598,N_11835);
nand U12103 (N_12103,N_11152,N_11771);
nand U12104 (N_12104,N_11458,N_11218);
nand U12105 (N_12105,N_11281,N_11307);
or U12106 (N_12106,N_11341,N_11854);
nor U12107 (N_12107,N_11846,N_11616);
nor U12108 (N_12108,N_11259,N_11887);
xnor U12109 (N_12109,N_11761,N_11743);
nor U12110 (N_12110,N_11751,N_11121);
xnor U12111 (N_12111,N_11285,N_11485);
and U12112 (N_12112,N_11129,N_11807);
xnor U12113 (N_12113,N_11353,N_11048);
nand U12114 (N_12114,N_11289,N_11377);
xor U12115 (N_12115,N_11254,N_11493);
nor U12116 (N_12116,N_11089,N_11740);
nor U12117 (N_12117,N_11546,N_11221);
and U12118 (N_12118,N_11621,N_11599);
nor U12119 (N_12119,N_11395,N_11555);
or U12120 (N_12120,N_11727,N_11749);
nand U12121 (N_12121,N_11898,N_11348);
and U12122 (N_12122,N_11558,N_11977);
nand U12123 (N_12123,N_11596,N_11499);
and U12124 (N_12124,N_11459,N_11145);
xnor U12125 (N_12125,N_11619,N_11216);
nand U12126 (N_12126,N_11220,N_11424);
xnor U12127 (N_12127,N_11701,N_11658);
nand U12128 (N_12128,N_11427,N_11742);
nand U12129 (N_12129,N_11939,N_11541);
or U12130 (N_12130,N_11306,N_11736);
xnor U12131 (N_12131,N_11989,N_11931);
xnor U12132 (N_12132,N_11393,N_11037);
nand U12133 (N_12133,N_11958,N_11767);
or U12134 (N_12134,N_11828,N_11913);
nand U12135 (N_12135,N_11159,N_11853);
xor U12136 (N_12136,N_11447,N_11648);
and U12137 (N_12137,N_11516,N_11100);
nand U12138 (N_12138,N_11641,N_11031);
xnor U12139 (N_12139,N_11798,N_11081);
xor U12140 (N_12140,N_11791,N_11109);
xnor U12141 (N_12141,N_11649,N_11967);
nand U12142 (N_12142,N_11829,N_11131);
and U12143 (N_12143,N_11148,N_11126);
or U12144 (N_12144,N_11722,N_11612);
nand U12145 (N_12145,N_11464,N_11385);
nand U12146 (N_12146,N_11095,N_11038);
xor U12147 (N_12147,N_11039,N_11293);
nand U12148 (N_12148,N_11021,N_11902);
nor U12149 (N_12149,N_11273,N_11440);
nand U12150 (N_12150,N_11774,N_11001);
xnor U12151 (N_12151,N_11214,N_11586);
or U12152 (N_12152,N_11613,N_11369);
or U12153 (N_12153,N_11786,N_11449);
xor U12154 (N_12154,N_11940,N_11071);
or U12155 (N_12155,N_11716,N_11494);
nor U12156 (N_12156,N_11300,N_11346);
nor U12157 (N_12157,N_11174,N_11355);
or U12158 (N_12158,N_11115,N_11881);
xnor U12159 (N_12159,N_11441,N_11004);
nand U12160 (N_12160,N_11438,N_11732);
xor U12161 (N_12161,N_11871,N_11257);
xnor U12162 (N_12162,N_11161,N_11975);
nand U12163 (N_12163,N_11968,N_11321);
nand U12164 (N_12164,N_11390,N_11705);
or U12165 (N_12165,N_11575,N_11238);
nand U12166 (N_12166,N_11818,N_11433);
nor U12167 (N_12167,N_11368,N_11793);
nor U12168 (N_12168,N_11924,N_11895);
and U12169 (N_12169,N_11883,N_11518);
nor U12170 (N_12170,N_11792,N_11759);
nand U12171 (N_12171,N_11122,N_11322);
or U12172 (N_12172,N_11389,N_11787);
xnor U12173 (N_12173,N_11600,N_11994);
xnor U12174 (N_12174,N_11343,N_11316);
nand U12175 (N_12175,N_11646,N_11462);
xor U12176 (N_12176,N_11267,N_11633);
xor U12177 (N_12177,N_11850,N_11176);
xor U12178 (N_12178,N_11339,N_11847);
xor U12179 (N_12179,N_11852,N_11337);
or U12180 (N_12180,N_11177,N_11796);
nand U12181 (N_12181,N_11626,N_11991);
nand U12182 (N_12182,N_11526,N_11603);
xor U12183 (N_12183,N_11816,N_11682);
nor U12184 (N_12184,N_11690,N_11136);
nor U12185 (N_12185,N_11114,N_11418);
nand U12186 (N_12186,N_11735,N_11490);
xnor U12187 (N_12187,N_11073,N_11812);
and U12188 (N_12188,N_11592,N_11423);
and U12189 (N_12189,N_11451,N_11146);
nor U12190 (N_12190,N_11750,N_11488);
nand U12191 (N_12191,N_11699,N_11416);
nor U12192 (N_12192,N_11856,N_11125);
and U12193 (N_12193,N_11930,N_11375);
and U12194 (N_12194,N_11301,N_11405);
or U12195 (N_12195,N_11589,N_11869);
xor U12196 (N_12196,N_11247,N_11966);
nand U12197 (N_12197,N_11899,N_11442);
nand U12198 (N_12198,N_11315,N_11910);
nor U12199 (N_12199,N_11789,N_11628);
and U12200 (N_12200,N_11820,N_11474);
and U12201 (N_12201,N_11237,N_11452);
nand U12202 (N_12202,N_11262,N_11591);
or U12203 (N_12203,N_11454,N_11143);
nor U12204 (N_12204,N_11318,N_11335);
nor U12205 (N_12205,N_11981,N_11784);
and U12206 (N_12206,N_11406,N_11371);
or U12207 (N_12207,N_11799,N_11745);
or U12208 (N_12208,N_11402,N_11134);
or U12209 (N_12209,N_11839,N_11047);
or U12210 (N_12210,N_11744,N_11949);
nor U12211 (N_12211,N_11664,N_11242);
nor U12212 (N_12212,N_11196,N_11758);
or U12213 (N_12213,N_11036,N_11072);
or U12214 (N_12214,N_11155,N_11500);
nand U12215 (N_12215,N_11615,N_11062);
xnor U12216 (N_12216,N_11519,N_11656);
and U12217 (N_12217,N_11965,N_11921);
xnor U12218 (N_12218,N_11453,N_11003);
nand U12219 (N_12219,N_11662,N_11525);
or U12220 (N_12220,N_11797,N_11739);
nor U12221 (N_12221,N_11045,N_11954);
xnor U12222 (N_12222,N_11282,N_11186);
nor U12223 (N_12223,N_11815,N_11480);
nor U12224 (N_12224,N_11502,N_11434);
nor U12225 (N_12225,N_11936,N_11078);
nor U12226 (N_12226,N_11671,N_11189);
nor U12227 (N_12227,N_11298,N_11431);
or U12228 (N_12228,N_11680,N_11184);
or U12229 (N_12229,N_11154,N_11167);
xor U12230 (N_12230,N_11521,N_11844);
nor U12231 (N_12231,N_11760,N_11268);
or U12232 (N_12232,N_11610,N_11495);
nor U12233 (N_12233,N_11843,N_11205);
xor U12234 (N_12234,N_11419,N_11753);
or U12235 (N_12235,N_11354,N_11795);
nand U12236 (N_12236,N_11092,N_11906);
nand U12237 (N_12237,N_11252,N_11934);
or U12238 (N_12238,N_11988,N_11688);
nor U12239 (N_12239,N_11594,N_11119);
and U12240 (N_12240,N_11979,N_11703);
nor U12241 (N_12241,N_11953,N_11618);
and U12242 (N_12242,N_11138,N_11425);
nor U12243 (N_12243,N_11547,N_11455);
or U12244 (N_12244,N_11099,N_11400);
or U12245 (N_12245,N_11779,N_11997);
nor U12246 (N_12246,N_11914,N_11863);
nor U12247 (N_12247,N_11077,N_11028);
and U12248 (N_12248,N_11006,N_11764);
or U12249 (N_12249,N_11082,N_11707);
and U12250 (N_12250,N_11227,N_11388);
xor U12251 (N_12251,N_11741,N_11193);
xnor U12252 (N_12252,N_11859,N_11042);
xor U12253 (N_12253,N_11723,N_11808);
xnor U12254 (N_12254,N_11016,N_11980);
nand U12255 (N_12255,N_11647,N_11497);
or U12256 (N_12256,N_11201,N_11040);
and U12257 (N_12257,N_11691,N_11860);
xnor U12258 (N_12258,N_11356,N_11948);
xor U12259 (N_12259,N_11232,N_11280);
xor U12260 (N_12260,N_11351,N_11130);
nor U12261 (N_12261,N_11399,N_11675);
nor U12262 (N_12262,N_11432,N_11228);
nand U12263 (N_12263,N_11950,N_11033);
nor U12264 (N_12264,N_11576,N_11565);
xor U12265 (N_12265,N_11358,N_11706);
or U12266 (N_12266,N_11086,N_11855);
nand U12267 (N_12267,N_11443,N_11068);
nand U12268 (N_12268,N_11849,N_11349);
xor U12269 (N_12269,N_11187,N_11861);
xnor U12270 (N_12270,N_11527,N_11178);
xor U12271 (N_12271,N_11310,N_11032);
xnor U12272 (N_12272,N_11556,N_11970);
or U12273 (N_12273,N_11909,N_11236);
and U12274 (N_12274,N_11049,N_11063);
xor U12275 (N_12275,N_11171,N_11827);
or U12276 (N_12276,N_11901,N_11392);
nand U12277 (N_12277,N_11244,N_11279);
nand U12278 (N_12278,N_11935,N_11700);
or U12279 (N_12279,N_11605,N_11561);
xnor U12280 (N_12280,N_11874,N_11826);
xor U12281 (N_12281,N_11995,N_11061);
or U12282 (N_12282,N_11435,N_11054);
and U12283 (N_12283,N_11780,N_11945);
xnor U12284 (N_12284,N_11436,N_11053);
nand U12285 (N_12285,N_11133,N_11276);
nand U12286 (N_12286,N_11407,N_11079);
and U12287 (N_12287,N_11769,N_11987);
nor U12288 (N_12288,N_11444,N_11872);
or U12289 (N_12289,N_11960,N_11587);
xnor U12290 (N_12290,N_11837,N_11217);
and U12291 (N_12291,N_11677,N_11207);
or U12292 (N_12292,N_11614,N_11098);
nand U12293 (N_12293,N_11409,N_11324);
or U12294 (N_12294,N_11581,N_11304);
nor U12295 (N_12295,N_11477,N_11755);
nand U12296 (N_12296,N_11050,N_11415);
or U12297 (N_12297,N_11173,N_11364);
xnor U12298 (N_12298,N_11692,N_11717);
and U12299 (N_12299,N_11069,N_11421);
nor U12300 (N_12300,N_11366,N_11135);
xor U12301 (N_12301,N_11381,N_11476);
xnor U12302 (N_12302,N_11199,N_11920);
or U12303 (N_12303,N_11070,N_11890);
or U12304 (N_12304,N_11972,N_11785);
xor U12305 (N_12305,N_11877,N_11790);
or U12306 (N_12306,N_11969,N_11757);
and U12307 (N_12307,N_11294,N_11020);
nand U12308 (N_12308,N_11998,N_11470);
or U12309 (N_12309,N_11029,N_11922);
nand U12310 (N_12310,N_11687,N_11231);
or U12311 (N_12311,N_11737,N_11466);
and U12312 (N_12312,N_11588,N_11927);
nor U12313 (N_12313,N_11274,N_11044);
nand U12314 (N_12314,N_11645,N_11570);
nor U12315 (N_12315,N_11014,N_11142);
and U12316 (N_12316,N_11107,N_11568);
xnor U12317 (N_12317,N_11532,N_11733);
and U12318 (N_12318,N_11642,N_11195);
nor U12319 (N_12319,N_11209,N_11673);
xor U12320 (N_12320,N_11842,N_11720);
or U12321 (N_12321,N_11666,N_11403);
nor U12322 (N_12322,N_11492,N_11000);
nand U12323 (N_12323,N_11051,N_11721);
xor U12324 (N_12324,N_11889,N_11810);
nand U12325 (N_12325,N_11713,N_11065);
and U12326 (N_12326,N_11275,N_11249);
nand U12327 (N_12327,N_11766,N_11465);
and U12328 (N_12328,N_11531,N_11437);
nand U12329 (N_12329,N_11536,N_11057);
and U12330 (N_12330,N_11422,N_11163);
or U12331 (N_12331,N_11296,N_11578);
and U12332 (N_12332,N_11768,N_11709);
and U12333 (N_12333,N_11295,N_11522);
or U12334 (N_12334,N_11251,N_11657);
and U12335 (N_12335,N_11794,N_11560);
nand U12336 (N_12336,N_11141,N_11277);
nand U12337 (N_12337,N_11539,N_11491);
or U12338 (N_12338,N_11222,N_11537);
and U12339 (N_12339,N_11963,N_11659);
or U12340 (N_12340,N_11066,N_11240);
xor U12341 (N_12341,N_11781,N_11926);
nand U12342 (N_12342,N_11487,N_11311);
nand U12343 (N_12343,N_11030,N_11456);
xor U12344 (N_12344,N_11034,N_11103);
nand U12345 (N_12345,N_11916,N_11026);
or U12346 (N_12346,N_11695,N_11158);
xnor U12347 (N_12347,N_11783,N_11515);
and U12348 (N_12348,N_11562,N_11563);
nor U12349 (N_12349,N_11668,N_11170);
or U12350 (N_12350,N_11915,N_11215);
or U12351 (N_12351,N_11778,N_11689);
or U12352 (N_12352,N_11111,N_11601);
nand U12353 (N_12353,N_11996,N_11959);
and U12354 (N_12354,N_11338,N_11097);
xor U12355 (N_12355,N_11928,N_11867);
nor U12356 (N_12356,N_11503,N_11912);
and U12357 (N_12357,N_11093,N_11475);
or U12358 (N_12358,N_11893,N_11669);
nor U12359 (N_12359,N_11595,N_11683);
nand U12360 (N_12360,N_11469,N_11635);
xor U12361 (N_12361,N_11482,N_11181);
or U12362 (N_12362,N_11643,N_11250);
or U12363 (N_12363,N_11233,N_11686);
or U12364 (N_12364,N_11352,N_11471);
nor U12365 (N_12365,N_11823,N_11806);
nor U12366 (N_12366,N_11297,N_11765);
and U12367 (N_12367,N_11105,N_11261);
nor U12368 (N_12368,N_11840,N_11088);
nand U12369 (N_12369,N_11880,N_11593);
xor U12370 (N_12370,N_11080,N_11210);
nor U12371 (N_12371,N_11363,N_11374);
and U12372 (N_12372,N_11708,N_11719);
nand U12373 (N_12373,N_11754,N_11472);
nor U12374 (N_12374,N_11224,N_11803);
and U12375 (N_12375,N_11336,N_11580);
xor U12376 (N_12376,N_11331,N_11937);
nand U12377 (N_12377,N_11166,N_11573);
xnor U12378 (N_12378,N_11617,N_11654);
nor U12379 (N_12379,N_11678,N_11198);
and U12380 (N_12380,N_11357,N_11825);
nand U12381 (N_12381,N_11943,N_11777);
xor U12382 (N_12382,N_11933,N_11160);
or U12383 (N_12383,N_11096,N_11417);
and U12384 (N_12384,N_11192,N_11213);
or U12385 (N_12385,N_11203,N_11961);
and U12386 (N_12386,N_11821,N_11340);
nand U12387 (N_12387,N_11430,N_11075);
and U12388 (N_12388,N_11652,N_11661);
nand U12389 (N_12389,N_11986,N_11162);
or U12390 (N_12390,N_11060,N_11660);
or U12391 (N_12391,N_11885,N_11775);
nor U12392 (N_12392,N_11408,N_11763);
or U12393 (N_12393,N_11005,N_11110);
or U12394 (N_12394,N_11091,N_11834);
xnor U12395 (N_12395,N_11597,N_11382);
xor U12396 (N_12396,N_11225,N_11523);
xor U12397 (N_12397,N_11964,N_11245);
nor U12398 (N_12398,N_11234,N_11731);
and U12399 (N_12399,N_11362,N_11376);
nor U12400 (N_12400,N_11211,N_11041);
xnor U12401 (N_12401,N_11554,N_11866);
nand U12402 (N_12402,N_11865,N_11380);
or U12403 (N_12403,N_11501,N_11255);
xnor U12404 (N_12404,N_11372,N_11450);
nand U12405 (N_12405,N_11299,N_11929);
nand U12406 (N_12406,N_11505,N_11944);
or U12407 (N_12407,N_11288,N_11564);
and U12408 (N_12408,N_11457,N_11264);
xnor U12409 (N_12409,N_11090,N_11637);
xor U12410 (N_12410,N_11112,N_11888);
nor U12411 (N_12411,N_11665,N_11553);
nor U12412 (N_12412,N_11286,N_11241);
and U12413 (N_12413,N_11908,N_11513);
and U12414 (N_12414,N_11776,N_11848);
nor U12415 (N_12415,N_11696,N_11667);
or U12416 (N_12416,N_11359,N_11035);
xnor U12417 (N_12417,N_11323,N_11510);
nand U12418 (N_12418,N_11715,N_11982);
or U12419 (N_12419,N_11172,N_11801);
and U12420 (N_12420,N_11278,N_11305);
or U12421 (N_12421,N_11303,N_11983);
nor U12422 (N_12422,N_11862,N_11788);
xor U12423 (N_12423,N_11992,N_11344);
and U12424 (N_12424,N_11347,N_11651);
nand U12425 (N_12425,N_11609,N_11870);
or U12426 (N_12426,N_11007,N_11085);
nand U12427 (N_12427,N_11813,N_11428);
and U12428 (N_12428,N_11212,N_11248);
nor U12429 (N_12429,N_11905,N_11917);
nand U12430 (N_12430,N_11378,N_11260);
and U12431 (N_12431,N_11468,N_11514);
nand U12432 (N_12432,N_11506,N_11023);
or U12433 (N_12433,N_11411,N_11165);
or U12434 (N_12434,N_11367,N_11653);
and U12435 (N_12435,N_11718,N_11140);
or U12436 (N_12436,N_11446,N_11156);
or U12437 (N_12437,N_11398,N_11627);
and U12438 (N_12438,N_11271,N_11639);
and U12439 (N_12439,N_11027,N_11302);
nand U12440 (N_12440,N_11876,N_11269);
and U12441 (N_12441,N_11941,N_11907);
xnor U12442 (N_12442,N_11325,N_11463);
nor U12443 (N_12443,N_11552,N_11951);
xnor U12444 (N_12444,N_11756,N_11632);
or U12445 (N_12445,N_11087,N_11946);
or U12446 (N_12446,N_11569,N_11882);
nor U12447 (N_12447,N_11128,N_11630);
and U12448 (N_12448,N_11538,N_11309);
nand U12449 (N_12449,N_11685,N_11365);
nand U12450 (N_12450,N_11833,N_11857);
and U12451 (N_12451,N_11694,N_11728);
xnor U12452 (N_12452,N_11342,N_11147);
and U12453 (N_12453,N_11256,N_11383);
or U12454 (N_12454,N_11394,N_11439);
and U12455 (N_12455,N_11043,N_11879);
nor U12456 (N_12456,N_11884,N_11971);
nand U12457 (N_12457,N_11074,N_11710);
nor U12458 (N_12458,N_11544,N_11010);
nor U12459 (N_12459,N_11226,N_11583);
nand U12460 (N_12460,N_11955,N_11904);
nand U12461 (N_12461,N_11679,N_11738);
or U12462 (N_12462,N_11018,N_11058);
nand U12463 (N_12463,N_11157,N_11507);
or U12464 (N_12464,N_11101,N_11530);
nand U12465 (N_12465,N_11219,N_11634);
or U12466 (N_12466,N_11083,N_11313);
or U12467 (N_12467,N_11345,N_11604);
or U12468 (N_12468,N_11024,N_11636);
nand U12469 (N_12469,N_11511,N_11900);
nor U12470 (N_12470,N_11809,N_11397);
or U12471 (N_12471,N_11025,N_11748);
or U12472 (N_12472,N_11802,N_11150);
xnor U12473 (N_12473,N_11164,N_11113);
or U12474 (N_12474,N_11243,N_11903);
nor U12475 (N_12475,N_11387,N_11373);
or U12476 (N_12476,N_11805,N_11734);
or U12477 (N_12477,N_11076,N_11974);
xnor U12478 (N_12478,N_11055,N_11116);
xnor U12479 (N_12479,N_11993,N_11875);
nor U12480 (N_12480,N_11401,N_11985);
nor U12481 (N_12481,N_11481,N_11319);
xor U12482 (N_12482,N_11631,N_11266);
nand U12483 (N_12483,N_11579,N_11608);
and U12484 (N_12484,N_11137,N_11548);
nor U12485 (N_12485,N_11412,N_11559);
nor U12486 (N_12486,N_11132,N_11426);
or U12487 (N_12487,N_11326,N_11263);
nor U12488 (N_12488,N_11729,N_11897);
nor U12489 (N_12489,N_11804,N_11762);
nor U12490 (N_12490,N_11253,N_11208);
or U12491 (N_12491,N_11191,N_11590);
nand U12492 (N_12492,N_11350,N_11123);
nor U12493 (N_12493,N_11206,N_11978);
nand U12494 (N_12494,N_11607,N_11711);
xnor U12495 (N_12495,N_11947,N_11106);
and U12496 (N_12496,N_11517,N_11923);
nor U12497 (N_12497,N_11011,N_11873);
or U12498 (N_12498,N_11841,N_11483);
nor U12499 (N_12499,N_11886,N_11602);
or U12500 (N_12500,N_11507,N_11258);
and U12501 (N_12501,N_11075,N_11944);
nor U12502 (N_12502,N_11912,N_11218);
nand U12503 (N_12503,N_11479,N_11326);
nand U12504 (N_12504,N_11706,N_11833);
or U12505 (N_12505,N_11371,N_11010);
nand U12506 (N_12506,N_11268,N_11846);
or U12507 (N_12507,N_11126,N_11382);
and U12508 (N_12508,N_11595,N_11024);
nor U12509 (N_12509,N_11587,N_11403);
or U12510 (N_12510,N_11357,N_11638);
or U12511 (N_12511,N_11407,N_11918);
xnor U12512 (N_12512,N_11259,N_11669);
or U12513 (N_12513,N_11264,N_11118);
xor U12514 (N_12514,N_11952,N_11651);
or U12515 (N_12515,N_11292,N_11570);
nand U12516 (N_12516,N_11023,N_11041);
xnor U12517 (N_12517,N_11594,N_11827);
and U12518 (N_12518,N_11316,N_11635);
or U12519 (N_12519,N_11607,N_11776);
nor U12520 (N_12520,N_11828,N_11404);
nand U12521 (N_12521,N_11245,N_11573);
nor U12522 (N_12522,N_11590,N_11425);
xor U12523 (N_12523,N_11328,N_11774);
or U12524 (N_12524,N_11273,N_11407);
xnor U12525 (N_12525,N_11579,N_11444);
and U12526 (N_12526,N_11632,N_11457);
xnor U12527 (N_12527,N_11385,N_11214);
nand U12528 (N_12528,N_11968,N_11852);
nand U12529 (N_12529,N_11315,N_11533);
nor U12530 (N_12530,N_11920,N_11792);
or U12531 (N_12531,N_11569,N_11354);
xnor U12532 (N_12532,N_11809,N_11944);
and U12533 (N_12533,N_11697,N_11718);
nor U12534 (N_12534,N_11480,N_11507);
nor U12535 (N_12535,N_11256,N_11564);
and U12536 (N_12536,N_11558,N_11727);
or U12537 (N_12537,N_11354,N_11424);
and U12538 (N_12538,N_11589,N_11949);
and U12539 (N_12539,N_11514,N_11959);
nand U12540 (N_12540,N_11668,N_11237);
nand U12541 (N_12541,N_11590,N_11608);
and U12542 (N_12542,N_11343,N_11358);
and U12543 (N_12543,N_11117,N_11262);
and U12544 (N_12544,N_11574,N_11064);
and U12545 (N_12545,N_11226,N_11822);
nor U12546 (N_12546,N_11383,N_11863);
or U12547 (N_12547,N_11740,N_11955);
xor U12548 (N_12548,N_11706,N_11699);
xor U12549 (N_12549,N_11311,N_11209);
xnor U12550 (N_12550,N_11071,N_11186);
nor U12551 (N_12551,N_11761,N_11633);
nor U12552 (N_12552,N_11865,N_11620);
or U12553 (N_12553,N_11341,N_11807);
nand U12554 (N_12554,N_11853,N_11179);
and U12555 (N_12555,N_11475,N_11567);
and U12556 (N_12556,N_11616,N_11999);
xnor U12557 (N_12557,N_11727,N_11833);
or U12558 (N_12558,N_11123,N_11713);
or U12559 (N_12559,N_11304,N_11741);
nand U12560 (N_12560,N_11761,N_11874);
and U12561 (N_12561,N_11175,N_11761);
and U12562 (N_12562,N_11493,N_11356);
nand U12563 (N_12563,N_11514,N_11479);
nor U12564 (N_12564,N_11003,N_11156);
nand U12565 (N_12565,N_11607,N_11576);
and U12566 (N_12566,N_11558,N_11282);
nand U12567 (N_12567,N_11759,N_11928);
nand U12568 (N_12568,N_11836,N_11809);
nor U12569 (N_12569,N_11826,N_11239);
xor U12570 (N_12570,N_11031,N_11423);
nor U12571 (N_12571,N_11608,N_11943);
or U12572 (N_12572,N_11174,N_11668);
or U12573 (N_12573,N_11113,N_11818);
and U12574 (N_12574,N_11148,N_11509);
nand U12575 (N_12575,N_11480,N_11961);
nand U12576 (N_12576,N_11558,N_11822);
nor U12577 (N_12577,N_11279,N_11483);
nand U12578 (N_12578,N_11688,N_11885);
nand U12579 (N_12579,N_11249,N_11154);
or U12580 (N_12580,N_11257,N_11235);
nor U12581 (N_12581,N_11092,N_11495);
or U12582 (N_12582,N_11505,N_11140);
nor U12583 (N_12583,N_11111,N_11555);
nor U12584 (N_12584,N_11521,N_11887);
xor U12585 (N_12585,N_11483,N_11967);
nor U12586 (N_12586,N_11698,N_11213);
or U12587 (N_12587,N_11743,N_11605);
nor U12588 (N_12588,N_11264,N_11816);
and U12589 (N_12589,N_11825,N_11921);
xor U12590 (N_12590,N_11284,N_11578);
nand U12591 (N_12591,N_11582,N_11360);
nor U12592 (N_12592,N_11194,N_11054);
nor U12593 (N_12593,N_11942,N_11505);
nand U12594 (N_12594,N_11452,N_11794);
and U12595 (N_12595,N_11602,N_11134);
nor U12596 (N_12596,N_11994,N_11437);
or U12597 (N_12597,N_11544,N_11594);
or U12598 (N_12598,N_11766,N_11893);
xor U12599 (N_12599,N_11056,N_11726);
and U12600 (N_12600,N_11844,N_11075);
nand U12601 (N_12601,N_11609,N_11460);
nand U12602 (N_12602,N_11463,N_11217);
or U12603 (N_12603,N_11377,N_11251);
or U12604 (N_12604,N_11237,N_11157);
nor U12605 (N_12605,N_11778,N_11823);
or U12606 (N_12606,N_11037,N_11643);
and U12607 (N_12607,N_11357,N_11118);
nor U12608 (N_12608,N_11682,N_11921);
and U12609 (N_12609,N_11383,N_11852);
nor U12610 (N_12610,N_11583,N_11273);
or U12611 (N_12611,N_11549,N_11783);
or U12612 (N_12612,N_11518,N_11891);
or U12613 (N_12613,N_11483,N_11426);
nand U12614 (N_12614,N_11389,N_11576);
nand U12615 (N_12615,N_11159,N_11066);
nand U12616 (N_12616,N_11265,N_11121);
or U12617 (N_12617,N_11302,N_11109);
xor U12618 (N_12618,N_11665,N_11901);
or U12619 (N_12619,N_11027,N_11445);
or U12620 (N_12620,N_11665,N_11598);
nand U12621 (N_12621,N_11805,N_11870);
nand U12622 (N_12622,N_11721,N_11213);
nand U12623 (N_12623,N_11562,N_11446);
nand U12624 (N_12624,N_11485,N_11289);
xor U12625 (N_12625,N_11655,N_11782);
nor U12626 (N_12626,N_11885,N_11098);
nand U12627 (N_12627,N_11353,N_11532);
nand U12628 (N_12628,N_11587,N_11493);
xor U12629 (N_12629,N_11733,N_11556);
xnor U12630 (N_12630,N_11762,N_11035);
nand U12631 (N_12631,N_11681,N_11080);
nand U12632 (N_12632,N_11505,N_11541);
nor U12633 (N_12633,N_11249,N_11117);
nand U12634 (N_12634,N_11934,N_11349);
nand U12635 (N_12635,N_11426,N_11373);
nor U12636 (N_12636,N_11733,N_11933);
nand U12637 (N_12637,N_11598,N_11808);
and U12638 (N_12638,N_11512,N_11193);
nand U12639 (N_12639,N_11808,N_11734);
or U12640 (N_12640,N_11240,N_11441);
or U12641 (N_12641,N_11913,N_11765);
nor U12642 (N_12642,N_11872,N_11236);
and U12643 (N_12643,N_11195,N_11746);
nand U12644 (N_12644,N_11425,N_11000);
nor U12645 (N_12645,N_11144,N_11637);
xnor U12646 (N_12646,N_11214,N_11007);
xnor U12647 (N_12647,N_11309,N_11063);
xor U12648 (N_12648,N_11483,N_11320);
nand U12649 (N_12649,N_11669,N_11399);
xnor U12650 (N_12650,N_11783,N_11651);
xor U12651 (N_12651,N_11859,N_11696);
nand U12652 (N_12652,N_11489,N_11722);
or U12653 (N_12653,N_11813,N_11278);
nand U12654 (N_12654,N_11440,N_11231);
nand U12655 (N_12655,N_11726,N_11048);
nand U12656 (N_12656,N_11535,N_11420);
xor U12657 (N_12657,N_11294,N_11609);
and U12658 (N_12658,N_11753,N_11062);
nor U12659 (N_12659,N_11596,N_11610);
and U12660 (N_12660,N_11102,N_11851);
nor U12661 (N_12661,N_11761,N_11576);
nand U12662 (N_12662,N_11715,N_11849);
nor U12663 (N_12663,N_11793,N_11563);
nand U12664 (N_12664,N_11251,N_11931);
xnor U12665 (N_12665,N_11629,N_11475);
and U12666 (N_12666,N_11576,N_11408);
or U12667 (N_12667,N_11494,N_11926);
nand U12668 (N_12668,N_11717,N_11679);
xor U12669 (N_12669,N_11670,N_11559);
and U12670 (N_12670,N_11501,N_11976);
or U12671 (N_12671,N_11693,N_11265);
xor U12672 (N_12672,N_11326,N_11704);
or U12673 (N_12673,N_11226,N_11209);
or U12674 (N_12674,N_11292,N_11056);
nor U12675 (N_12675,N_11545,N_11073);
and U12676 (N_12676,N_11314,N_11287);
and U12677 (N_12677,N_11508,N_11606);
xnor U12678 (N_12678,N_11467,N_11597);
and U12679 (N_12679,N_11428,N_11425);
and U12680 (N_12680,N_11005,N_11021);
xor U12681 (N_12681,N_11650,N_11260);
or U12682 (N_12682,N_11689,N_11853);
nor U12683 (N_12683,N_11176,N_11863);
or U12684 (N_12684,N_11507,N_11485);
and U12685 (N_12685,N_11001,N_11820);
nor U12686 (N_12686,N_11749,N_11402);
xor U12687 (N_12687,N_11616,N_11873);
nor U12688 (N_12688,N_11401,N_11254);
and U12689 (N_12689,N_11812,N_11504);
or U12690 (N_12690,N_11477,N_11314);
nor U12691 (N_12691,N_11558,N_11083);
nor U12692 (N_12692,N_11499,N_11330);
nand U12693 (N_12693,N_11234,N_11706);
or U12694 (N_12694,N_11129,N_11314);
nor U12695 (N_12695,N_11903,N_11239);
or U12696 (N_12696,N_11500,N_11150);
and U12697 (N_12697,N_11995,N_11430);
and U12698 (N_12698,N_11795,N_11399);
nor U12699 (N_12699,N_11498,N_11926);
xor U12700 (N_12700,N_11810,N_11229);
or U12701 (N_12701,N_11621,N_11733);
or U12702 (N_12702,N_11202,N_11601);
or U12703 (N_12703,N_11363,N_11908);
nand U12704 (N_12704,N_11250,N_11850);
nor U12705 (N_12705,N_11297,N_11441);
nor U12706 (N_12706,N_11372,N_11644);
or U12707 (N_12707,N_11183,N_11576);
xnor U12708 (N_12708,N_11178,N_11364);
xnor U12709 (N_12709,N_11640,N_11623);
xor U12710 (N_12710,N_11693,N_11304);
nor U12711 (N_12711,N_11251,N_11924);
nand U12712 (N_12712,N_11631,N_11743);
nor U12713 (N_12713,N_11166,N_11913);
nand U12714 (N_12714,N_11503,N_11928);
nor U12715 (N_12715,N_11630,N_11566);
xnor U12716 (N_12716,N_11359,N_11711);
and U12717 (N_12717,N_11430,N_11150);
and U12718 (N_12718,N_11343,N_11016);
nor U12719 (N_12719,N_11863,N_11264);
or U12720 (N_12720,N_11553,N_11594);
nand U12721 (N_12721,N_11532,N_11831);
or U12722 (N_12722,N_11035,N_11614);
nand U12723 (N_12723,N_11560,N_11207);
nor U12724 (N_12724,N_11934,N_11056);
and U12725 (N_12725,N_11619,N_11304);
nand U12726 (N_12726,N_11465,N_11348);
nor U12727 (N_12727,N_11409,N_11704);
xnor U12728 (N_12728,N_11561,N_11846);
nand U12729 (N_12729,N_11529,N_11349);
or U12730 (N_12730,N_11839,N_11927);
or U12731 (N_12731,N_11004,N_11728);
nand U12732 (N_12732,N_11226,N_11554);
and U12733 (N_12733,N_11267,N_11766);
or U12734 (N_12734,N_11832,N_11195);
or U12735 (N_12735,N_11487,N_11360);
nand U12736 (N_12736,N_11457,N_11798);
or U12737 (N_12737,N_11497,N_11465);
or U12738 (N_12738,N_11936,N_11178);
and U12739 (N_12739,N_11892,N_11951);
xnor U12740 (N_12740,N_11900,N_11153);
nor U12741 (N_12741,N_11327,N_11326);
nor U12742 (N_12742,N_11398,N_11953);
or U12743 (N_12743,N_11607,N_11430);
nand U12744 (N_12744,N_11360,N_11375);
xnor U12745 (N_12745,N_11018,N_11766);
nor U12746 (N_12746,N_11884,N_11297);
nor U12747 (N_12747,N_11136,N_11252);
xnor U12748 (N_12748,N_11596,N_11898);
or U12749 (N_12749,N_11378,N_11779);
nand U12750 (N_12750,N_11773,N_11493);
and U12751 (N_12751,N_11570,N_11196);
or U12752 (N_12752,N_11227,N_11295);
or U12753 (N_12753,N_11882,N_11583);
or U12754 (N_12754,N_11446,N_11093);
and U12755 (N_12755,N_11681,N_11188);
xnor U12756 (N_12756,N_11956,N_11161);
or U12757 (N_12757,N_11999,N_11770);
nor U12758 (N_12758,N_11965,N_11123);
nor U12759 (N_12759,N_11821,N_11994);
or U12760 (N_12760,N_11969,N_11577);
and U12761 (N_12761,N_11449,N_11219);
or U12762 (N_12762,N_11267,N_11947);
and U12763 (N_12763,N_11686,N_11977);
nor U12764 (N_12764,N_11948,N_11307);
and U12765 (N_12765,N_11570,N_11615);
or U12766 (N_12766,N_11422,N_11166);
nor U12767 (N_12767,N_11900,N_11094);
and U12768 (N_12768,N_11563,N_11324);
xor U12769 (N_12769,N_11685,N_11513);
nor U12770 (N_12770,N_11990,N_11478);
nand U12771 (N_12771,N_11078,N_11663);
nor U12772 (N_12772,N_11636,N_11040);
and U12773 (N_12773,N_11038,N_11305);
nor U12774 (N_12774,N_11018,N_11981);
and U12775 (N_12775,N_11104,N_11609);
and U12776 (N_12776,N_11517,N_11362);
nand U12777 (N_12777,N_11812,N_11325);
xnor U12778 (N_12778,N_11050,N_11212);
or U12779 (N_12779,N_11386,N_11581);
and U12780 (N_12780,N_11788,N_11245);
or U12781 (N_12781,N_11985,N_11662);
or U12782 (N_12782,N_11785,N_11451);
nand U12783 (N_12783,N_11038,N_11742);
nor U12784 (N_12784,N_11753,N_11746);
xor U12785 (N_12785,N_11284,N_11835);
nand U12786 (N_12786,N_11898,N_11208);
nand U12787 (N_12787,N_11499,N_11707);
nand U12788 (N_12788,N_11200,N_11823);
nor U12789 (N_12789,N_11353,N_11826);
nand U12790 (N_12790,N_11189,N_11766);
or U12791 (N_12791,N_11751,N_11187);
or U12792 (N_12792,N_11506,N_11020);
nor U12793 (N_12793,N_11362,N_11855);
nor U12794 (N_12794,N_11076,N_11586);
xnor U12795 (N_12795,N_11092,N_11103);
xor U12796 (N_12796,N_11085,N_11050);
xor U12797 (N_12797,N_11580,N_11508);
and U12798 (N_12798,N_11767,N_11070);
nor U12799 (N_12799,N_11049,N_11914);
nor U12800 (N_12800,N_11159,N_11999);
or U12801 (N_12801,N_11156,N_11843);
xor U12802 (N_12802,N_11659,N_11464);
or U12803 (N_12803,N_11263,N_11775);
and U12804 (N_12804,N_11375,N_11132);
xnor U12805 (N_12805,N_11161,N_11355);
and U12806 (N_12806,N_11938,N_11112);
or U12807 (N_12807,N_11032,N_11148);
nor U12808 (N_12808,N_11013,N_11798);
nand U12809 (N_12809,N_11925,N_11548);
and U12810 (N_12810,N_11262,N_11569);
and U12811 (N_12811,N_11485,N_11212);
and U12812 (N_12812,N_11582,N_11814);
xor U12813 (N_12813,N_11462,N_11890);
and U12814 (N_12814,N_11772,N_11150);
xor U12815 (N_12815,N_11454,N_11552);
and U12816 (N_12816,N_11779,N_11455);
xnor U12817 (N_12817,N_11599,N_11515);
and U12818 (N_12818,N_11115,N_11064);
nand U12819 (N_12819,N_11994,N_11484);
nor U12820 (N_12820,N_11247,N_11634);
nand U12821 (N_12821,N_11921,N_11833);
nand U12822 (N_12822,N_11368,N_11778);
and U12823 (N_12823,N_11174,N_11908);
nand U12824 (N_12824,N_11919,N_11904);
nand U12825 (N_12825,N_11487,N_11877);
nand U12826 (N_12826,N_11429,N_11053);
and U12827 (N_12827,N_11826,N_11727);
xor U12828 (N_12828,N_11574,N_11258);
nand U12829 (N_12829,N_11517,N_11441);
xnor U12830 (N_12830,N_11769,N_11006);
xnor U12831 (N_12831,N_11104,N_11809);
nand U12832 (N_12832,N_11604,N_11265);
nor U12833 (N_12833,N_11828,N_11779);
or U12834 (N_12834,N_11305,N_11783);
xor U12835 (N_12835,N_11101,N_11470);
nor U12836 (N_12836,N_11800,N_11119);
xor U12837 (N_12837,N_11492,N_11924);
xor U12838 (N_12838,N_11812,N_11796);
nand U12839 (N_12839,N_11203,N_11637);
nor U12840 (N_12840,N_11405,N_11469);
nand U12841 (N_12841,N_11173,N_11355);
xor U12842 (N_12842,N_11365,N_11464);
and U12843 (N_12843,N_11422,N_11329);
or U12844 (N_12844,N_11709,N_11113);
and U12845 (N_12845,N_11807,N_11552);
and U12846 (N_12846,N_11920,N_11177);
nor U12847 (N_12847,N_11476,N_11570);
nor U12848 (N_12848,N_11248,N_11550);
xor U12849 (N_12849,N_11976,N_11496);
nor U12850 (N_12850,N_11178,N_11855);
nor U12851 (N_12851,N_11669,N_11677);
and U12852 (N_12852,N_11845,N_11920);
nor U12853 (N_12853,N_11511,N_11248);
and U12854 (N_12854,N_11424,N_11671);
nor U12855 (N_12855,N_11085,N_11396);
or U12856 (N_12856,N_11520,N_11784);
and U12857 (N_12857,N_11466,N_11434);
and U12858 (N_12858,N_11298,N_11650);
xor U12859 (N_12859,N_11990,N_11504);
and U12860 (N_12860,N_11146,N_11457);
xnor U12861 (N_12861,N_11872,N_11508);
or U12862 (N_12862,N_11334,N_11890);
nand U12863 (N_12863,N_11248,N_11569);
nor U12864 (N_12864,N_11666,N_11277);
xor U12865 (N_12865,N_11637,N_11599);
or U12866 (N_12866,N_11047,N_11304);
xnor U12867 (N_12867,N_11859,N_11723);
nand U12868 (N_12868,N_11245,N_11448);
and U12869 (N_12869,N_11612,N_11027);
or U12870 (N_12870,N_11072,N_11618);
nor U12871 (N_12871,N_11908,N_11800);
nor U12872 (N_12872,N_11622,N_11017);
nand U12873 (N_12873,N_11206,N_11600);
nor U12874 (N_12874,N_11642,N_11257);
nor U12875 (N_12875,N_11118,N_11956);
or U12876 (N_12876,N_11270,N_11016);
nor U12877 (N_12877,N_11590,N_11058);
and U12878 (N_12878,N_11398,N_11317);
or U12879 (N_12879,N_11520,N_11227);
nor U12880 (N_12880,N_11089,N_11692);
or U12881 (N_12881,N_11955,N_11725);
and U12882 (N_12882,N_11489,N_11195);
nor U12883 (N_12883,N_11700,N_11155);
nand U12884 (N_12884,N_11702,N_11660);
and U12885 (N_12885,N_11061,N_11088);
or U12886 (N_12886,N_11894,N_11402);
xor U12887 (N_12887,N_11193,N_11698);
nor U12888 (N_12888,N_11575,N_11582);
and U12889 (N_12889,N_11670,N_11979);
or U12890 (N_12890,N_11653,N_11072);
nor U12891 (N_12891,N_11985,N_11728);
nor U12892 (N_12892,N_11284,N_11616);
and U12893 (N_12893,N_11478,N_11840);
xor U12894 (N_12894,N_11450,N_11249);
xor U12895 (N_12895,N_11097,N_11383);
nor U12896 (N_12896,N_11514,N_11310);
xor U12897 (N_12897,N_11037,N_11091);
or U12898 (N_12898,N_11431,N_11739);
and U12899 (N_12899,N_11147,N_11519);
xor U12900 (N_12900,N_11647,N_11191);
xor U12901 (N_12901,N_11252,N_11393);
nor U12902 (N_12902,N_11447,N_11446);
xor U12903 (N_12903,N_11285,N_11454);
nor U12904 (N_12904,N_11678,N_11447);
and U12905 (N_12905,N_11163,N_11961);
nor U12906 (N_12906,N_11839,N_11980);
nand U12907 (N_12907,N_11527,N_11369);
or U12908 (N_12908,N_11092,N_11271);
or U12909 (N_12909,N_11088,N_11505);
xor U12910 (N_12910,N_11085,N_11145);
nor U12911 (N_12911,N_11716,N_11637);
nand U12912 (N_12912,N_11738,N_11964);
or U12913 (N_12913,N_11788,N_11946);
or U12914 (N_12914,N_11726,N_11088);
nor U12915 (N_12915,N_11417,N_11044);
and U12916 (N_12916,N_11266,N_11323);
nor U12917 (N_12917,N_11593,N_11564);
nor U12918 (N_12918,N_11833,N_11814);
and U12919 (N_12919,N_11048,N_11454);
xnor U12920 (N_12920,N_11303,N_11746);
nand U12921 (N_12921,N_11127,N_11370);
or U12922 (N_12922,N_11397,N_11028);
nand U12923 (N_12923,N_11004,N_11336);
xnor U12924 (N_12924,N_11472,N_11046);
nor U12925 (N_12925,N_11156,N_11475);
nand U12926 (N_12926,N_11684,N_11777);
nor U12927 (N_12927,N_11581,N_11096);
or U12928 (N_12928,N_11781,N_11861);
nor U12929 (N_12929,N_11727,N_11753);
or U12930 (N_12930,N_11500,N_11667);
nor U12931 (N_12931,N_11109,N_11157);
nor U12932 (N_12932,N_11645,N_11322);
xnor U12933 (N_12933,N_11106,N_11677);
nor U12934 (N_12934,N_11398,N_11144);
nand U12935 (N_12935,N_11423,N_11189);
nand U12936 (N_12936,N_11806,N_11590);
or U12937 (N_12937,N_11645,N_11419);
and U12938 (N_12938,N_11413,N_11096);
xor U12939 (N_12939,N_11566,N_11744);
or U12940 (N_12940,N_11703,N_11287);
nor U12941 (N_12941,N_11912,N_11229);
nor U12942 (N_12942,N_11975,N_11054);
nand U12943 (N_12943,N_11597,N_11551);
nand U12944 (N_12944,N_11081,N_11552);
nor U12945 (N_12945,N_11437,N_11988);
or U12946 (N_12946,N_11078,N_11330);
nor U12947 (N_12947,N_11422,N_11998);
nand U12948 (N_12948,N_11897,N_11936);
xnor U12949 (N_12949,N_11522,N_11676);
nand U12950 (N_12950,N_11731,N_11708);
nand U12951 (N_12951,N_11887,N_11833);
and U12952 (N_12952,N_11942,N_11966);
nand U12953 (N_12953,N_11290,N_11891);
nand U12954 (N_12954,N_11496,N_11486);
or U12955 (N_12955,N_11378,N_11477);
nor U12956 (N_12956,N_11368,N_11440);
xor U12957 (N_12957,N_11130,N_11596);
nand U12958 (N_12958,N_11858,N_11430);
nand U12959 (N_12959,N_11589,N_11526);
and U12960 (N_12960,N_11327,N_11133);
and U12961 (N_12961,N_11683,N_11760);
nor U12962 (N_12962,N_11179,N_11603);
and U12963 (N_12963,N_11631,N_11491);
or U12964 (N_12964,N_11216,N_11707);
and U12965 (N_12965,N_11501,N_11610);
or U12966 (N_12966,N_11976,N_11533);
or U12967 (N_12967,N_11375,N_11770);
or U12968 (N_12968,N_11396,N_11566);
and U12969 (N_12969,N_11804,N_11644);
and U12970 (N_12970,N_11663,N_11253);
and U12971 (N_12971,N_11582,N_11497);
nand U12972 (N_12972,N_11088,N_11226);
or U12973 (N_12973,N_11861,N_11303);
nor U12974 (N_12974,N_11920,N_11143);
xor U12975 (N_12975,N_11437,N_11672);
nand U12976 (N_12976,N_11005,N_11272);
or U12977 (N_12977,N_11013,N_11758);
or U12978 (N_12978,N_11997,N_11935);
nand U12979 (N_12979,N_11855,N_11013);
or U12980 (N_12980,N_11981,N_11548);
and U12981 (N_12981,N_11797,N_11205);
and U12982 (N_12982,N_11356,N_11431);
xnor U12983 (N_12983,N_11242,N_11455);
nor U12984 (N_12984,N_11416,N_11163);
and U12985 (N_12985,N_11707,N_11698);
nor U12986 (N_12986,N_11480,N_11986);
or U12987 (N_12987,N_11940,N_11752);
nand U12988 (N_12988,N_11721,N_11090);
nand U12989 (N_12989,N_11197,N_11603);
and U12990 (N_12990,N_11804,N_11923);
and U12991 (N_12991,N_11229,N_11751);
xor U12992 (N_12992,N_11400,N_11278);
and U12993 (N_12993,N_11592,N_11288);
xor U12994 (N_12994,N_11091,N_11669);
nand U12995 (N_12995,N_11751,N_11805);
or U12996 (N_12996,N_11077,N_11832);
or U12997 (N_12997,N_11896,N_11362);
and U12998 (N_12998,N_11248,N_11031);
nand U12999 (N_12999,N_11185,N_11401);
or U13000 (N_13000,N_12689,N_12196);
or U13001 (N_13001,N_12106,N_12650);
xnor U13002 (N_13002,N_12765,N_12772);
nor U13003 (N_13003,N_12861,N_12289);
or U13004 (N_13004,N_12680,N_12438);
nand U13005 (N_13005,N_12967,N_12397);
nand U13006 (N_13006,N_12691,N_12775);
or U13007 (N_13007,N_12928,N_12527);
nand U13008 (N_13008,N_12159,N_12790);
xnor U13009 (N_13009,N_12748,N_12989);
nand U13010 (N_13010,N_12164,N_12589);
nor U13011 (N_13011,N_12509,N_12107);
nor U13012 (N_13012,N_12126,N_12912);
nand U13013 (N_13013,N_12666,N_12962);
or U13014 (N_13014,N_12905,N_12312);
xor U13015 (N_13015,N_12080,N_12430);
nor U13016 (N_13016,N_12632,N_12668);
nand U13017 (N_13017,N_12693,N_12324);
and U13018 (N_13018,N_12971,N_12092);
nand U13019 (N_13019,N_12182,N_12955);
and U13020 (N_13020,N_12858,N_12373);
nand U13021 (N_13021,N_12402,N_12352);
xnor U13022 (N_13022,N_12079,N_12291);
or U13023 (N_13023,N_12115,N_12619);
or U13024 (N_13024,N_12348,N_12728);
nor U13025 (N_13025,N_12094,N_12747);
or U13026 (N_13026,N_12843,N_12207);
xor U13027 (N_13027,N_12276,N_12097);
nand U13028 (N_13028,N_12902,N_12481);
nand U13029 (N_13029,N_12633,N_12778);
nand U13030 (N_13030,N_12796,N_12114);
nand U13031 (N_13031,N_12354,N_12317);
and U13032 (N_13032,N_12646,N_12046);
xor U13033 (N_13033,N_12030,N_12878);
and U13034 (N_13034,N_12978,N_12952);
and U13035 (N_13035,N_12282,N_12837);
nor U13036 (N_13036,N_12547,N_12724);
xor U13037 (N_13037,N_12785,N_12740);
nand U13038 (N_13038,N_12839,N_12720);
xnor U13039 (N_13039,N_12382,N_12970);
nor U13040 (N_13040,N_12745,N_12241);
nand U13041 (N_13041,N_12514,N_12395);
xnor U13042 (N_13042,N_12715,N_12223);
or U13043 (N_13043,N_12679,N_12766);
or U13044 (N_13044,N_12059,N_12564);
or U13045 (N_13045,N_12303,N_12009);
and U13046 (N_13046,N_12227,N_12625);
and U13047 (N_13047,N_12371,N_12937);
or U13048 (N_13048,N_12256,N_12587);
xnor U13049 (N_13049,N_12469,N_12802);
nand U13050 (N_13050,N_12898,N_12375);
or U13051 (N_13051,N_12511,N_12882);
nand U13052 (N_13052,N_12670,N_12119);
nor U13053 (N_13053,N_12322,N_12661);
nand U13054 (N_13054,N_12866,N_12501);
nor U13055 (N_13055,N_12873,N_12914);
and U13056 (N_13056,N_12355,N_12151);
nor U13057 (N_13057,N_12200,N_12684);
nor U13058 (N_13058,N_12815,N_12268);
nor U13059 (N_13059,N_12518,N_12368);
and U13060 (N_13060,N_12083,N_12822);
nand U13061 (N_13061,N_12489,N_12176);
and U13062 (N_13062,N_12433,N_12797);
nor U13063 (N_13063,N_12440,N_12338);
and U13064 (N_13064,N_12102,N_12480);
xor U13065 (N_13065,N_12854,N_12627);
nand U13066 (N_13066,N_12285,N_12571);
nor U13067 (N_13067,N_12408,N_12038);
xnor U13068 (N_13068,N_12321,N_12769);
or U13069 (N_13069,N_12135,N_12683);
nor U13070 (N_13070,N_12148,N_12770);
xnor U13071 (N_13071,N_12892,N_12346);
nor U13072 (N_13072,N_12064,N_12620);
xnor U13073 (N_13073,N_12697,N_12942);
and U13074 (N_13074,N_12434,N_12936);
and U13075 (N_13075,N_12795,N_12213);
nand U13076 (N_13076,N_12677,N_12019);
nor U13077 (N_13077,N_12474,N_12713);
nand U13078 (N_13078,N_12893,N_12144);
and U13079 (N_13079,N_12238,N_12570);
or U13080 (N_13080,N_12170,N_12737);
xor U13081 (N_13081,N_12246,N_12362);
nor U13082 (N_13082,N_12986,N_12486);
nor U13083 (N_13083,N_12572,N_12202);
or U13084 (N_13084,N_12002,N_12876);
xnor U13085 (N_13085,N_12593,N_12130);
nand U13086 (N_13086,N_12027,N_12350);
nand U13087 (N_13087,N_12215,N_12051);
and U13088 (N_13088,N_12807,N_12789);
or U13089 (N_13089,N_12628,N_12143);
or U13090 (N_13090,N_12274,N_12603);
nand U13091 (N_13091,N_12476,N_12911);
or U13092 (N_13092,N_12386,N_12872);
or U13093 (N_13093,N_12310,N_12655);
or U13094 (N_13094,N_12738,N_12688);
nand U13095 (N_13095,N_12602,N_12886);
and U13096 (N_13096,N_12071,N_12442);
or U13097 (N_13097,N_12311,N_12743);
nand U13098 (N_13098,N_12584,N_12423);
nand U13099 (N_13099,N_12218,N_12733);
nand U13100 (N_13100,N_12913,N_12762);
nor U13101 (N_13101,N_12831,N_12718);
xnor U13102 (N_13102,N_12384,N_12431);
xor U13103 (N_13103,N_12337,N_12214);
nor U13104 (N_13104,N_12596,N_12190);
nand U13105 (N_13105,N_12921,N_12543);
nand U13106 (N_13106,N_12884,N_12128);
nor U13107 (N_13107,N_12754,N_12640);
nor U13108 (N_13108,N_12172,N_12869);
or U13109 (N_13109,N_12178,N_12923);
nor U13110 (N_13110,N_12709,N_12675);
xor U13111 (N_13111,N_12468,N_12700);
and U13112 (N_13112,N_12297,N_12294);
xor U13113 (N_13113,N_12193,N_12774);
nand U13114 (N_13114,N_12209,N_12407);
nand U13115 (N_13115,N_12611,N_12577);
xnor U13116 (N_13116,N_12216,N_12544);
xor U13117 (N_13117,N_12055,N_12562);
and U13118 (N_13118,N_12483,N_12413);
or U13119 (N_13119,N_12281,N_12336);
nand U13120 (N_13120,N_12567,N_12755);
nand U13121 (N_13121,N_12284,N_12290);
and U13122 (N_13122,N_12982,N_12706);
xor U13123 (N_13123,N_12864,N_12805);
xor U13124 (N_13124,N_12053,N_12592);
nand U13125 (N_13125,N_12934,N_12113);
or U13126 (N_13126,N_12824,N_12141);
and U13127 (N_13127,N_12887,N_12503);
or U13128 (N_13128,N_12367,N_12445);
nand U13129 (N_13129,N_12192,N_12441);
nor U13130 (N_13130,N_12663,N_12535);
nor U13131 (N_13131,N_12808,N_12605);
or U13132 (N_13132,N_12764,N_12767);
and U13133 (N_13133,N_12149,N_12761);
or U13134 (N_13134,N_12492,N_12272);
nor U13135 (N_13135,N_12449,N_12418);
xor U13136 (N_13136,N_12964,N_12615);
nand U13137 (N_13137,N_12819,N_12933);
nand U13138 (N_13138,N_12183,N_12590);
nor U13139 (N_13139,N_12333,N_12366);
or U13140 (N_13140,N_12278,N_12206);
nand U13141 (N_13141,N_12653,N_12614);
nand U13142 (N_13142,N_12062,N_12205);
or U13143 (N_13143,N_12283,N_12542);
nor U13144 (N_13144,N_12990,N_12957);
nor U13145 (N_13145,N_12944,N_12198);
xor U13146 (N_13146,N_12123,N_12217);
or U13147 (N_13147,N_12604,N_12082);
and U13148 (N_13148,N_12341,N_12788);
nor U13149 (N_13149,N_12125,N_12648);
nand U13150 (N_13150,N_12034,N_12457);
nand U13151 (N_13151,N_12105,N_12001);
or U13152 (N_13152,N_12070,N_12409);
nand U13153 (N_13153,N_12383,N_12996);
nor U13154 (N_13154,N_12950,N_12003);
or U13155 (N_13155,N_12818,N_12085);
nor U13156 (N_13156,N_12557,N_12103);
or U13157 (N_13157,N_12353,N_12129);
nor U13158 (N_13158,N_12906,N_12484);
xnor U13159 (N_13159,N_12553,N_12840);
or U13160 (N_13160,N_12307,N_12545);
nor U13161 (N_13161,N_12581,N_12953);
or U13162 (N_13162,N_12502,N_12154);
nor U13163 (N_13163,N_12041,N_12271);
xor U13164 (N_13164,N_12412,N_12191);
and U13165 (N_13165,N_12047,N_12237);
nor U13166 (N_13166,N_12983,N_12320);
xor U13167 (N_13167,N_12393,N_12617);
nand U13168 (N_13168,N_12210,N_12540);
and U13169 (N_13169,N_12050,N_12758);
or U13170 (N_13170,N_12834,N_12612);
xor U13171 (N_13171,N_12479,N_12220);
nand U13172 (N_13172,N_12351,N_12376);
or U13173 (N_13173,N_12226,N_12088);
and U13174 (N_13174,N_12736,N_12844);
or U13175 (N_13175,N_12969,N_12782);
or U13176 (N_13176,N_12756,N_12139);
or U13177 (N_13177,N_12156,N_12018);
and U13178 (N_13178,N_12915,N_12414);
nor U13179 (N_13179,N_12500,N_12069);
xor U13180 (N_13180,N_12781,N_12599);
nand U13181 (N_13181,N_12702,N_12812);
or U13182 (N_13182,N_12232,N_12949);
xor U13183 (N_13183,N_12157,N_12314);
or U13184 (N_13184,N_12254,N_12568);
nor U13185 (N_13185,N_12258,N_12426);
nor U13186 (N_13186,N_12332,N_12823);
xor U13187 (N_13187,N_12270,N_12832);
nor U13188 (N_13188,N_12305,N_12561);
xnor U13189 (N_13189,N_12750,N_12842);
nor U13190 (N_13190,N_12794,N_12120);
nand U13191 (N_13191,N_12012,N_12968);
nand U13192 (N_13192,N_12095,N_12931);
or U13193 (N_13193,N_12856,N_12877);
xor U13194 (N_13194,N_12828,N_12536);
xor U13195 (N_13195,N_12826,N_12731);
nand U13196 (N_13196,N_12777,N_12188);
nand U13197 (N_13197,N_12173,N_12954);
xor U13198 (N_13198,N_12017,N_12171);
nand U13199 (N_13199,N_12401,N_12405);
nand U13200 (N_13200,N_12394,N_12998);
nand U13201 (N_13201,N_12028,N_12516);
nand U13202 (N_13202,N_12779,N_12265);
or U13203 (N_13203,N_12185,N_12037);
nor U13204 (N_13204,N_12043,N_12885);
or U13205 (N_13205,N_12669,N_12259);
or U13206 (N_13206,N_12380,N_12287);
and U13207 (N_13207,N_12415,N_12879);
xor U13208 (N_13208,N_12626,N_12428);
nor U13209 (N_13209,N_12391,N_12867);
or U13210 (N_13210,N_12150,N_12871);
nand U13211 (N_13211,N_12077,N_12065);
nor U13212 (N_13212,N_12644,N_12586);
or U13213 (N_13213,N_12707,N_12630);
or U13214 (N_13214,N_12240,N_12916);
or U13215 (N_13215,N_12965,N_12497);
nor U13216 (N_13216,N_12865,N_12918);
nor U13217 (N_13217,N_12498,N_12058);
nor U13218 (N_13218,N_12298,N_12494);
nand U13219 (N_13219,N_12846,N_12506);
and U13220 (N_13220,N_12784,N_12345);
and U13221 (N_13221,N_12569,N_12624);
nor U13222 (N_13222,N_12253,N_12111);
nand U13223 (N_13223,N_12868,N_12277);
xor U13224 (N_13224,N_12881,N_12904);
xnor U13225 (N_13225,N_12061,N_12326);
xnor U13226 (N_13226,N_12295,N_12184);
and U13227 (N_13227,N_12145,N_12076);
nand U13228 (N_13228,N_12976,N_12450);
nand U13229 (N_13229,N_12255,N_12424);
and U13230 (N_13230,N_12711,N_12752);
nor U13231 (N_13231,N_12563,N_12180);
nor U13232 (N_13232,N_12153,N_12899);
or U13233 (N_13233,N_12610,N_12979);
nor U13234 (N_13234,N_12487,N_12600);
nor U13235 (N_13235,N_12629,N_12493);
nand U13236 (N_13236,N_12559,N_12725);
xor U13237 (N_13237,N_12531,N_12851);
xor U13238 (N_13238,N_12212,N_12883);
xnor U13239 (N_13239,N_12020,N_12045);
xor U13240 (N_13240,N_12089,N_12991);
or U13241 (N_13241,N_12806,N_12980);
xor U13242 (N_13242,N_12472,N_12809);
and U13243 (N_13243,N_12040,N_12390);
nand U13244 (N_13244,N_12467,N_12739);
and U13245 (N_13245,N_12512,N_12730);
and U13246 (N_13246,N_12452,N_12665);
or U13247 (N_13247,N_12727,N_12168);
nand U13248 (N_13248,N_12793,N_12301);
or U13249 (N_13249,N_12072,N_12427);
xnor U13250 (N_13250,N_12288,N_12901);
nor U13251 (N_13251,N_12521,N_12622);
nor U13252 (N_13252,N_12895,N_12201);
or U13253 (N_13253,N_12654,N_12676);
or U13254 (N_13254,N_12437,N_12233);
and U13255 (N_13255,N_12133,N_12786);
or U13256 (N_13256,N_12685,N_12993);
xor U13257 (N_13257,N_12313,N_12532);
nor U13258 (N_13258,N_12455,N_12147);
nor U13259 (N_13259,N_12499,N_12121);
and U13260 (N_13260,N_12652,N_12664);
and U13261 (N_13261,N_12162,N_12091);
xnor U13262 (N_13262,N_12432,N_12349);
xor U13263 (N_13263,N_12546,N_12267);
nor U13264 (N_13264,N_12098,N_12800);
xnor U13265 (N_13265,N_12101,N_12835);
or U13266 (N_13266,N_12946,N_12035);
nand U13267 (N_13267,N_12396,N_12451);
and U13268 (N_13268,N_12379,N_12330);
nand U13269 (N_13269,N_12328,N_12538);
nand U13270 (N_13270,N_12810,N_12732);
xnor U13271 (N_13271,N_12565,N_12029);
nor U13272 (N_13272,N_12453,N_12146);
or U13273 (N_13273,N_12616,N_12613);
xor U13274 (N_13274,N_12224,N_12066);
xor U13275 (N_13275,N_12174,N_12308);
nand U13276 (N_13276,N_12473,N_12932);
xnor U13277 (N_13277,N_12465,N_12903);
nand U13278 (N_13278,N_12024,N_12109);
or U13279 (N_13279,N_12334,N_12852);
xnor U13280 (N_13280,N_12554,N_12853);
and U13281 (N_13281,N_12021,N_12874);
nand U13282 (N_13282,N_12358,N_12672);
or U13283 (N_13283,N_12257,N_12327);
xor U13284 (N_13284,N_12813,N_12791);
or U13285 (N_13285,N_12300,N_12023);
nor U13286 (N_13286,N_12890,N_12959);
xnor U13287 (N_13287,N_12988,N_12639);
nor U13288 (N_13288,N_12179,N_12995);
xnor U13289 (N_13289,N_12555,N_12010);
or U13290 (N_13290,N_12588,N_12578);
or U13291 (N_13291,N_12695,N_12768);
or U13292 (N_13292,N_12122,N_12016);
or U13293 (N_13293,N_12804,N_12448);
xnor U13294 (N_13294,N_12471,N_12690);
and U13295 (N_13295,N_12504,N_12722);
nor U13296 (N_13296,N_12054,N_12712);
and U13297 (N_13297,N_12817,N_12529);
nor U13298 (N_13298,N_12015,N_12667);
and U13299 (N_13299,N_12389,N_12920);
or U13300 (N_13300,N_12533,N_12436);
or U13301 (N_13301,N_12658,N_12703);
nand U13302 (N_13302,N_12994,N_12651);
and U13303 (N_13303,N_12787,N_12435);
and U13304 (N_13304,N_12574,N_12007);
or U13305 (N_13305,N_12771,N_12721);
nor U13306 (N_13306,N_12325,N_12236);
nor U13307 (N_13307,N_12378,N_12673);
nand U13308 (N_13308,N_12042,N_12696);
xnor U13309 (N_13309,N_12419,N_12573);
or U13310 (N_13310,N_12595,N_12166);
xnor U13311 (N_13311,N_12365,N_12929);
nor U13312 (N_13312,N_12385,N_12943);
or U13313 (N_13313,N_12249,N_12845);
or U13314 (N_13314,N_12520,N_12678);
and U13315 (N_13315,N_12919,N_12264);
nand U13316 (N_13316,N_12359,N_12636);
nand U13317 (N_13317,N_12247,N_12369);
xnor U13318 (N_13318,N_12411,N_12894);
xor U13319 (N_13319,N_12275,N_12907);
nand U13320 (N_13320,N_12960,N_12470);
nor U13321 (N_13321,N_12075,N_12136);
and U13322 (N_13322,N_12243,N_12086);
xor U13323 (N_13323,N_12643,N_12485);
and U13324 (N_13324,N_12203,N_12177);
and U13325 (N_13325,N_12909,N_12165);
or U13326 (N_13326,N_12692,N_12124);
nor U13327 (N_13327,N_12211,N_12974);
xnor U13328 (N_13328,N_12608,N_12235);
or U13329 (N_13329,N_12776,N_12958);
nor U13330 (N_13330,N_12081,N_12830);
xor U13331 (N_13331,N_12742,N_12416);
nand U13332 (N_13332,N_12033,N_12558);
or U13333 (N_13333,N_12269,N_12780);
nor U13334 (N_13334,N_12112,N_12187);
nor U13335 (N_13335,N_12403,N_12726);
xnor U13336 (N_13336,N_12528,N_12744);
xor U13337 (N_13337,N_12118,N_12841);
and U13338 (N_13338,N_12025,N_12985);
and U13339 (N_13339,N_12134,N_12838);
nand U13340 (N_13340,N_12517,N_12417);
or U13341 (N_13341,N_12930,N_12621);
or U13342 (N_13342,N_12260,N_12585);
xnor U13343 (N_13343,N_12387,N_12420);
xor U13344 (N_13344,N_12821,N_12142);
and U13345 (N_13345,N_12251,N_12701);
or U13346 (N_13346,N_12548,N_12011);
or U13347 (N_13347,N_12292,N_12347);
xnor U13348 (N_13348,N_12315,N_12847);
or U13349 (N_13349,N_12078,N_12488);
nor U13350 (N_13350,N_12456,N_12963);
xnor U13351 (N_13351,N_12231,N_12250);
and U13352 (N_13352,N_12704,N_12048);
nand U13353 (N_13353,N_12917,N_12645);
and U13354 (N_13354,N_12461,N_12541);
nand U13355 (N_13355,N_12763,N_12671);
xor U13356 (N_13356,N_12863,N_12977);
xor U13357 (N_13357,N_12966,N_12792);
nor U13358 (N_13358,N_12972,N_12399);
nand U13359 (N_13359,N_12642,N_12381);
and U13360 (N_13360,N_12199,N_12374);
and U13361 (N_13361,N_12222,N_12910);
and U13362 (N_13362,N_12344,N_12013);
nor U13363 (N_13363,N_12576,N_12656);
nand U13364 (N_13364,N_12286,N_12049);
xnor U13365 (N_13365,N_12039,N_12490);
nor U13366 (N_13366,N_12195,N_12219);
or U13367 (N_13367,N_12137,N_12044);
and U13368 (N_13368,N_12496,N_12753);
nand U13369 (N_13369,N_12956,N_12108);
nand U13370 (N_13370,N_12947,N_12400);
nor U13371 (N_13371,N_12244,N_12388);
xor U13372 (N_13372,N_12908,N_12896);
xor U13373 (N_13373,N_12729,N_12623);
nor U13374 (N_13374,N_12659,N_12221);
xnor U13375 (N_13375,N_12507,N_12860);
and U13376 (N_13376,N_12634,N_12783);
nand U13377 (N_13377,N_12060,N_12579);
or U13378 (N_13378,N_12997,N_12372);
xnor U13379 (N_13379,N_12052,N_12463);
and U13380 (N_13380,N_12951,N_12719);
nor U13381 (N_13381,N_12454,N_12682);
xor U13382 (N_13382,N_12252,N_12318);
nand U13383 (N_13383,N_12132,N_12361);
nor U13384 (N_13384,N_12100,N_12022);
xor U13385 (N_13385,N_12938,N_12566);
xor U13386 (N_13386,N_12900,N_12889);
xnor U13387 (N_13387,N_12342,N_12186);
and U13388 (N_13388,N_12716,N_12591);
and U13389 (N_13389,N_12825,N_12421);
and U13390 (N_13390,N_12710,N_12984);
nand U13391 (N_13391,N_12006,N_12466);
xnor U13392 (N_13392,N_12439,N_12228);
and U13393 (N_13393,N_12104,N_12127);
nor U13394 (N_13394,N_12096,N_12773);
and U13395 (N_13395,N_12340,N_12987);
and U13396 (N_13396,N_12891,N_12357);
nor U13397 (N_13397,N_12302,N_12057);
xor U13398 (N_13398,N_12973,N_12681);
and U13399 (N_13399,N_12849,N_12087);
nand U13400 (N_13400,N_12945,N_12000);
and U13401 (N_13401,N_12309,N_12870);
xnor U13402 (N_13402,N_12491,N_12935);
nor U13403 (N_13403,N_12940,N_12140);
nand U13404 (N_13404,N_12152,N_12525);
nor U13405 (N_13405,N_12687,N_12036);
and U13406 (N_13406,N_12981,N_12827);
nand U13407 (N_13407,N_12117,N_12280);
and U13408 (N_13408,N_12723,N_12647);
xnor U13409 (N_13409,N_12460,N_12759);
or U13410 (N_13410,N_12194,N_12008);
or U13411 (N_13411,N_12167,N_12074);
nor U13412 (N_13412,N_12638,N_12410);
nor U13413 (N_13413,N_12458,N_12601);
and U13414 (N_13414,N_12635,N_12475);
nor U13415 (N_13415,N_12530,N_12422);
nor U13416 (N_13416,N_12641,N_12926);
and U13417 (N_13417,N_12245,N_12478);
xor U13418 (N_13418,N_12161,N_12404);
nor U13419 (N_13419,N_12927,N_12698);
or U13420 (N_13420,N_12263,N_12319);
nor U13421 (N_13421,N_12948,N_12110);
nand U13422 (N_13422,N_12848,N_12556);
and U13423 (N_13423,N_12299,N_12004);
and U13424 (N_13424,N_12099,N_12513);
and U13425 (N_13425,N_12462,N_12163);
xnor U13426 (N_13426,N_12444,N_12924);
nand U13427 (N_13427,N_12293,N_12551);
and U13428 (N_13428,N_12522,N_12406);
or U13429 (N_13429,N_12583,N_12734);
nor U13430 (N_13430,N_12741,N_12242);
nor U13431 (N_13431,N_12014,N_12446);
or U13432 (N_13432,N_12005,N_12888);
and U13433 (N_13433,N_12582,N_12803);
and U13434 (N_13434,N_12814,N_12477);
nand U13435 (N_13435,N_12032,N_12735);
nand U13436 (N_13436,N_12816,N_12580);
or U13437 (N_13437,N_12631,N_12594);
or U13438 (N_13438,N_12699,N_12534);
nand U13439 (N_13439,N_12859,N_12537);
xnor U13440 (N_13440,N_12833,N_12811);
or U13441 (N_13441,N_12248,N_12169);
or U13442 (N_13442,N_12155,N_12686);
nor U13443 (N_13443,N_12597,N_12464);
xnor U13444 (N_13444,N_12515,N_12550);
nand U13445 (N_13445,N_12660,N_12181);
nor U13446 (N_13446,N_12850,N_12575);
nand U13447 (N_13447,N_12875,N_12356);
or U13448 (N_13448,N_12552,N_12459);
or U13449 (N_13449,N_12961,N_12799);
nor U13450 (N_13450,N_12539,N_12234);
xnor U13451 (N_13451,N_12829,N_12992);
or U13452 (N_13452,N_12225,N_12158);
or U13453 (N_13453,N_12801,N_12067);
nor U13454 (N_13454,N_12197,N_12939);
and U13455 (N_13455,N_12377,N_12323);
or U13456 (N_13456,N_12273,N_12482);
or U13457 (N_13457,N_12363,N_12922);
nand U13458 (N_13458,N_12261,N_12714);
nand U13459 (N_13459,N_12266,N_12549);
or U13460 (N_13460,N_12068,N_12607);
nand U13461 (N_13461,N_12116,N_12370);
nor U13462 (N_13462,N_12598,N_12090);
nand U13463 (N_13463,N_12708,N_12523);
xnor U13464 (N_13464,N_12606,N_12508);
and U13465 (N_13465,N_12757,N_12398);
nand U13466 (N_13466,N_12609,N_12857);
nand U13467 (N_13467,N_12204,N_12510);
nand U13468 (N_13468,N_12335,N_12073);
xor U13469 (N_13469,N_12084,N_12443);
nand U13470 (N_13470,N_12798,N_12208);
nor U13471 (N_13471,N_12694,N_12705);
nor U13472 (N_13472,N_12749,N_12392);
nor U13473 (N_13473,N_12160,N_12239);
and U13474 (N_13474,N_12031,N_12138);
xnor U13475 (N_13475,N_12560,N_12279);
nor U13476 (N_13476,N_12820,N_12093);
or U13477 (N_13477,N_12760,N_12316);
xor U13478 (N_13478,N_12425,N_12526);
nor U13479 (N_13479,N_12505,N_12339);
nand U13480 (N_13480,N_12855,N_12999);
nand U13481 (N_13481,N_12674,N_12941);
and U13482 (N_13482,N_12447,N_12331);
xor U13483 (N_13483,N_12056,N_12495);
xor U13484 (N_13484,N_12262,N_12230);
nor U13485 (N_13485,N_12897,N_12662);
nor U13486 (N_13486,N_12519,N_12925);
nor U13487 (N_13487,N_12296,N_12429);
nor U13488 (N_13488,N_12751,N_12229);
xor U13489 (N_13489,N_12880,N_12329);
and U13490 (N_13490,N_12063,N_12836);
xnor U13491 (N_13491,N_12862,N_12746);
and U13492 (N_13492,N_12649,N_12306);
and U13493 (N_13493,N_12026,N_12524);
and U13494 (N_13494,N_12364,N_12618);
nor U13495 (N_13495,N_12304,N_12637);
nand U13496 (N_13496,N_12131,N_12975);
xor U13497 (N_13497,N_12717,N_12189);
xor U13498 (N_13498,N_12175,N_12657);
nor U13499 (N_13499,N_12360,N_12343);
xnor U13500 (N_13500,N_12426,N_12966);
xor U13501 (N_13501,N_12973,N_12824);
nor U13502 (N_13502,N_12638,N_12077);
xor U13503 (N_13503,N_12469,N_12449);
nor U13504 (N_13504,N_12055,N_12537);
or U13505 (N_13505,N_12614,N_12801);
nor U13506 (N_13506,N_12059,N_12720);
or U13507 (N_13507,N_12589,N_12597);
or U13508 (N_13508,N_12297,N_12524);
nand U13509 (N_13509,N_12070,N_12412);
xnor U13510 (N_13510,N_12645,N_12283);
or U13511 (N_13511,N_12088,N_12353);
nand U13512 (N_13512,N_12100,N_12775);
xor U13513 (N_13513,N_12304,N_12106);
or U13514 (N_13514,N_12589,N_12484);
nand U13515 (N_13515,N_12576,N_12628);
nor U13516 (N_13516,N_12452,N_12798);
and U13517 (N_13517,N_12866,N_12541);
nor U13518 (N_13518,N_12866,N_12821);
xor U13519 (N_13519,N_12611,N_12409);
xnor U13520 (N_13520,N_12247,N_12165);
nor U13521 (N_13521,N_12882,N_12242);
or U13522 (N_13522,N_12560,N_12383);
nor U13523 (N_13523,N_12766,N_12271);
or U13524 (N_13524,N_12351,N_12852);
or U13525 (N_13525,N_12515,N_12199);
and U13526 (N_13526,N_12983,N_12931);
nor U13527 (N_13527,N_12478,N_12694);
nor U13528 (N_13528,N_12707,N_12846);
and U13529 (N_13529,N_12389,N_12240);
xor U13530 (N_13530,N_12837,N_12495);
xnor U13531 (N_13531,N_12721,N_12901);
or U13532 (N_13532,N_12630,N_12550);
and U13533 (N_13533,N_12337,N_12564);
nand U13534 (N_13534,N_12499,N_12363);
nand U13535 (N_13535,N_12028,N_12576);
or U13536 (N_13536,N_12690,N_12093);
or U13537 (N_13537,N_12656,N_12657);
or U13538 (N_13538,N_12484,N_12028);
nand U13539 (N_13539,N_12526,N_12320);
and U13540 (N_13540,N_12351,N_12375);
and U13541 (N_13541,N_12313,N_12901);
nor U13542 (N_13542,N_12693,N_12987);
nor U13543 (N_13543,N_12065,N_12932);
nand U13544 (N_13544,N_12117,N_12671);
xnor U13545 (N_13545,N_12576,N_12877);
or U13546 (N_13546,N_12811,N_12683);
and U13547 (N_13547,N_12804,N_12480);
or U13548 (N_13548,N_12219,N_12691);
nand U13549 (N_13549,N_12591,N_12691);
nand U13550 (N_13550,N_12986,N_12889);
nand U13551 (N_13551,N_12459,N_12070);
and U13552 (N_13552,N_12705,N_12901);
and U13553 (N_13553,N_12585,N_12780);
xor U13554 (N_13554,N_12475,N_12153);
or U13555 (N_13555,N_12869,N_12178);
or U13556 (N_13556,N_12848,N_12942);
and U13557 (N_13557,N_12729,N_12456);
xor U13558 (N_13558,N_12577,N_12137);
and U13559 (N_13559,N_12305,N_12225);
and U13560 (N_13560,N_12015,N_12206);
nor U13561 (N_13561,N_12179,N_12141);
or U13562 (N_13562,N_12554,N_12692);
and U13563 (N_13563,N_12099,N_12366);
or U13564 (N_13564,N_12948,N_12576);
nor U13565 (N_13565,N_12367,N_12726);
nand U13566 (N_13566,N_12695,N_12039);
nor U13567 (N_13567,N_12309,N_12700);
nor U13568 (N_13568,N_12150,N_12794);
and U13569 (N_13569,N_12481,N_12644);
and U13570 (N_13570,N_12488,N_12100);
nand U13571 (N_13571,N_12121,N_12407);
nor U13572 (N_13572,N_12896,N_12814);
xnor U13573 (N_13573,N_12899,N_12137);
xor U13574 (N_13574,N_12165,N_12005);
or U13575 (N_13575,N_12902,N_12030);
nor U13576 (N_13576,N_12425,N_12424);
nor U13577 (N_13577,N_12919,N_12696);
nor U13578 (N_13578,N_12559,N_12308);
nor U13579 (N_13579,N_12023,N_12471);
nor U13580 (N_13580,N_12403,N_12426);
nand U13581 (N_13581,N_12695,N_12672);
xor U13582 (N_13582,N_12745,N_12369);
nand U13583 (N_13583,N_12916,N_12885);
and U13584 (N_13584,N_12867,N_12467);
or U13585 (N_13585,N_12258,N_12211);
and U13586 (N_13586,N_12410,N_12686);
and U13587 (N_13587,N_12119,N_12960);
nor U13588 (N_13588,N_12513,N_12185);
and U13589 (N_13589,N_12834,N_12455);
or U13590 (N_13590,N_12202,N_12794);
nand U13591 (N_13591,N_12407,N_12752);
nor U13592 (N_13592,N_12353,N_12152);
nand U13593 (N_13593,N_12124,N_12863);
xnor U13594 (N_13594,N_12622,N_12708);
and U13595 (N_13595,N_12625,N_12358);
or U13596 (N_13596,N_12378,N_12246);
nor U13597 (N_13597,N_12877,N_12733);
and U13598 (N_13598,N_12154,N_12712);
nand U13599 (N_13599,N_12945,N_12641);
and U13600 (N_13600,N_12670,N_12935);
nor U13601 (N_13601,N_12841,N_12946);
nor U13602 (N_13602,N_12992,N_12661);
xnor U13603 (N_13603,N_12532,N_12933);
and U13604 (N_13604,N_12303,N_12687);
nand U13605 (N_13605,N_12779,N_12952);
and U13606 (N_13606,N_12156,N_12103);
nand U13607 (N_13607,N_12768,N_12794);
or U13608 (N_13608,N_12309,N_12685);
xor U13609 (N_13609,N_12438,N_12821);
or U13610 (N_13610,N_12063,N_12481);
nand U13611 (N_13611,N_12693,N_12610);
xor U13612 (N_13612,N_12777,N_12027);
nand U13613 (N_13613,N_12433,N_12794);
xor U13614 (N_13614,N_12357,N_12877);
xnor U13615 (N_13615,N_12256,N_12628);
nand U13616 (N_13616,N_12631,N_12695);
and U13617 (N_13617,N_12437,N_12963);
and U13618 (N_13618,N_12695,N_12512);
xnor U13619 (N_13619,N_12544,N_12792);
nand U13620 (N_13620,N_12664,N_12340);
nand U13621 (N_13621,N_12479,N_12219);
and U13622 (N_13622,N_12914,N_12519);
and U13623 (N_13623,N_12234,N_12059);
xnor U13624 (N_13624,N_12648,N_12919);
and U13625 (N_13625,N_12819,N_12021);
and U13626 (N_13626,N_12740,N_12012);
or U13627 (N_13627,N_12627,N_12236);
nand U13628 (N_13628,N_12567,N_12788);
nand U13629 (N_13629,N_12526,N_12355);
and U13630 (N_13630,N_12961,N_12095);
nor U13631 (N_13631,N_12588,N_12118);
xnor U13632 (N_13632,N_12738,N_12891);
or U13633 (N_13633,N_12134,N_12692);
or U13634 (N_13634,N_12498,N_12714);
and U13635 (N_13635,N_12280,N_12692);
nand U13636 (N_13636,N_12017,N_12495);
xor U13637 (N_13637,N_12603,N_12043);
or U13638 (N_13638,N_12301,N_12531);
nor U13639 (N_13639,N_12438,N_12271);
nand U13640 (N_13640,N_12367,N_12285);
nand U13641 (N_13641,N_12910,N_12067);
or U13642 (N_13642,N_12523,N_12870);
and U13643 (N_13643,N_12636,N_12134);
and U13644 (N_13644,N_12910,N_12879);
and U13645 (N_13645,N_12750,N_12784);
nand U13646 (N_13646,N_12573,N_12248);
and U13647 (N_13647,N_12813,N_12532);
nor U13648 (N_13648,N_12648,N_12949);
xnor U13649 (N_13649,N_12308,N_12939);
nand U13650 (N_13650,N_12889,N_12161);
nor U13651 (N_13651,N_12681,N_12895);
nand U13652 (N_13652,N_12975,N_12053);
nand U13653 (N_13653,N_12857,N_12840);
nor U13654 (N_13654,N_12521,N_12350);
nand U13655 (N_13655,N_12026,N_12942);
xor U13656 (N_13656,N_12303,N_12824);
nand U13657 (N_13657,N_12895,N_12421);
xor U13658 (N_13658,N_12715,N_12188);
and U13659 (N_13659,N_12350,N_12615);
or U13660 (N_13660,N_12103,N_12480);
or U13661 (N_13661,N_12936,N_12973);
xnor U13662 (N_13662,N_12173,N_12361);
nand U13663 (N_13663,N_12865,N_12526);
nor U13664 (N_13664,N_12647,N_12061);
nand U13665 (N_13665,N_12325,N_12151);
and U13666 (N_13666,N_12712,N_12010);
nand U13667 (N_13667,N_12051,N_12751);
xnor U13668 (N_13668,N_12212,N_12388);
nor U13669 (N_13669,N_12195,N_12016);
xnor U13670 (N_13670,N_12836,N_12412);
nor U13671 (N_13671,N_12680,N_12603);
or U13672 (N_13672,N_12935,N_12795);
nand U13673 (N_13673,N_12557,N_12422);
xor U13674 (N_13674,N_12312,N_12293);
nand U13675 (N_13675,N_12461,N_12315);
and U13676 (N_13676,N_12716,N_12310);
or U13677 (N_13677,N_12847,N_12102);
nand U13678 (N_13678,N_12638,N_12219);
xor U13679 (N_13679,N_12005,N_12751);
xor U13680 (N_13680,N_12384,N_12227);
nor U13681 (N_13681,N_12408,N_12946);
or U13682 (N_13682,N_12748,N_12594);
or U13683 (N_13683,N_12449,N_12742);
and U13684 (N_13684,N_12004,N_12789);
and U13685 (N_13685,N_12157,N_12102);
xor U13686 (N_13686,N_12745,N_12663);
nand U13687 (N_13687,N_12914,N_12652);
xor U13688 (N_13688,N_12159,N_12949);
or U13689 (N_13689,N_12630,N_12678);
nor U13690 (N_13690,N_12827,N_12636);
nor U13691 (N_13691,N_12367,N_12072);
nor U13692 (N_13692,N_12566,N_12029);
xnor U13693 (N_13693,N_12688,N_12457);
xor U13694 (N_13694,N_12232,N_12156);
or U13695 (N_13695,N_12284,N_12610);
nand U13696 (N_13696,N_12254,N_12708);
nand U13697 (N_13697,N_12030,N_12558);
xor U13698 (N_13698,N_12694,N_12168);
nor U13699 (N_13699,N_12446,N_12687);
nor U13700 (N_13700,N_12316,N_12941);
or U13701 (N_13701,N_12847,N_12021);
nor U13702 (N_13702,N_12382,N_12505);
nor U13703 (N_13703,N_12322,N_12788);
and U13704 (N_13704,N_12392,N_12106);
or U13705 (N_13705,N_12515,N_12281);
and U13706 (N_13706,N_12742,N_12711);
nand U13707 (N_13707,N_12942,N_12380);
nor U13708 (N_13708,N_12759,N_12510);
nand U13709 (N_13709,N_12294,N_12394);
xor U13710 (N_13710,N_12276,N_12080);
xor U13711 (N_13711,N_12657,N_12391);
nand U13712 (N_13712,N_12327,N_12640);
and U13713 (N_13713,N_12146,N_12312);
and U13714 (N_13714,N_12454,N_12482);
nand U13715 (N_13715,N_12355,N_12041);
nor U13716 (N_13716,N_12452,N_12138);
nand U13717 (N_13717,N_12276,N_12419);
xor U13718 (N_13718,N_12029,N_12552);
nand U13719 (N_13719,N_12887,N_12499);
xnor U13720 (N_13720,N_12782,N_12668);
nor U13721 (N_13721,N_12409,N_12873);
nor U13722 (N_13722,N_12818,N_12380);
nand U13723 (N_13723,N_12425,N_12242);
or U13724 (N_13724,N_12651,N_12407);
nor U13725 (N_13725,N_12749,N_12025);
nand U13726 (N_13726,N_12284,N_12355);
and U13727 (N_13727,N_12293,N_12108);
nand U13728 (N_13728,N_12807,N_12644);
nand U13729 (N_13729,N_12031,N_12425);
nor U13730 (N_13730,N_12849,N_12922);
nor U13731 (N_13731,N_12546,N_12609);
or U13732 (N_13732,N_12412,N_12455);
and U13733 (N_13733,N_12370,N_12258);
and U13734 (N_13734,N_12160,N_12766);
xor U13735 (N_13735,N_12250,N_12267);
nor U13736 (N_13736,N_12328,N_12031);
or U13737 (N_13737,N_12619,N_12185);
nand U13738 (N_13738,N_12306,N_12020);
or U13739 (N_13739,N_12994,N_12452);
xor U13740 (N_13740,N_12215,N_12435);
nor U13741 (N_13741,N_12623,N_12881);
nor U13742 (N_13742,N_12000,N_12148);
nor U13743 (N_13743,N_12425,N_12684);
and U13744 (N_13744,N_12288,N_12388);
or U13745 (N_13745,N_12622,N_12618);
and U13746 (N_13746,N_12389,N_12520);
nor U13747 (N_13747,N_12805,N_12990);
xor U13748 (N_13748,N_12420,N_12814);
and U13749 (N_13749,N_12814,N_12495);
xnor U13750 (N_13750,N_12761,N_12930);
xor U13751 (N_13751,N_12034,N_12760);
xor U13752 (N_13752,N_12988,N_12664);
nand U13753 (N_13753,N_12376,N_12923);
and U13754 (N_13754,N_12751,N_12025);
or U13755 (N_13755,N_12949,N_12619);
nand U13756 (N_13756,N_12184,N_12571);
or U13757 (N_13757,N_12707,N_12299);
xor U13758 (N_13758,N_12789,N_12329);
nor U13759 (N_13759,N_12788,N_12036);
xnor U13760 (N_13760,N_12901,N_12589);
or U13761 (N_13761,N_12833,N_12333);
nand U13762 (N_13762,N_12917,N_12842);
nor U13763 (N_13763,N_12277,N_12579);
and U13764 (N_13764,N_12624,N_12658);
and U13765 (N_13765,N_12646,N_12173);
xor U13766 (N_13766,N_12716,N_12287);
or U13767 (N_13767,N_12493,N_12736);
xor U13768 (N_13768,N_12999,N_12359);
nand U13769 (N_13769,N_12237,N_12751);
and U13770 (N_13770,N_12234,N_12665);
xnor U13771 (N_13771,N_12404,N_12667);
or U13772 (N_13772,N_12415,N_12611);
nor U13773 (N_13773,N_12599,N_12579);
nand U13774 (N_13774,N_12549,N_12777);
or U13775 (N_13775,N_12731,N_12491);
nor U13776 (N_13776,N_12223,N_12819);
and U13777 (N_13777,N_12971,N_12732);
xor U13778 (N_13778,N_12384,N_12724);
and U13779 (N_13779,N_12072,N_12395);
nand U13780 (N_13780,N_12961,N_12360);
nor U13781 (N_13781,N_12695,N_12950);
and U13782 (N_13782,N_12711,N_12246);
and U13783 (N_13783,N_12344,N_12117);
nand U13784 (N_13784,N_12265,N_12806);
nor U13785 (N_13785,N_12574,N_12317);
nand U13786 (N_13786,N_12166,N_12471);
nor U13787 (N_13787,N_12199,N_12714);
or U13788 (N_13788,N_12265,N_12697);
or U13789 (N_13789,N_12694,N_12047);
xor U13790 (N_13790,N_12601,N_12662);
and U13791 (N_13791,N_12972,N_12690);
nor U13792 (N_13792,N_12437,N_12717);
xor U13793 (N_13793,N_12295,N_12387);
nand U13794 (N_13794,N_12790,N_12324);
and U13795 (N_13795,N_12064,N_12391);
and U13796 (N_13796,N_12351,N_12418);
nand U13797 (N_13797,N_12787,N_12932);
xnor U13798 (N_13798,N_12944,N_12502);
and U13799 (N_13799,N_12960,N_12633);
xnor U13800 (N_13800,N_12306,N_12777);
and U13801 (N_13801,N_12707,N_12497);
and U13802 (N_13802,N_12235,N_12193);
xnor U13803 (N_13803,N_12449,N_12815);
nand U13804 (N_13804,N_12330,N_12890);
xnor U13805 (N_13805,N_12812,N_12157);
or U13806 (N_13806,N_12795,N_12745);
xor U13807 (N_13807,N_12573,N_12209);
xnor U13808 (N_13808,N_12049,N_12302);
nor U13809 (N_13809,N_12750,N_12967);
nand U13810 (N_13810,N_12411,N_12451);
or U13811 (N_13811,N_12989,N_12792);
xnor U13812 (N_13812,N_12307,N_12891);
xnor U13813 (N_13813,N_12586,N_12293);
nor U13814 (N_13814,N_12263,N_12030);
nor U13815 (N_13815,N_12411,N_12753);
xor U13816 (N_13816,N_12518,N_12608);
nand U13817 (N_13817,N_12015,N_12830);
nand U13818 (N_13818,N_12637,N_12799);
nor U13819 (N_13819,N_12692,N_12168);
and U13820 (N_13820,N_12944,N_12513);
nor U13821 (N_13821,N_12877,N_12204);
or U13822 (N_13822,N_12032,N_12469);
or U13823 (N_13823,N_12198,N_12252);
nor U13824 (N_13824,N_12352,N_12661);
or U13825 (N_13825,N_12184,N_12449);
nand U13826 (N_13826,N_12559,N_12066);
nand U13827 (N_13827,N_12413,N_12916);
nand U13828 (N_13828,N_12001,N_12211);
xnor U13829 (N_13829,N_12295,N_12055);
xnor U13830 (N_13830,N_12917,N_12211);
xnor U13831 (N_13831,N_12998,N_12087);
nor U13832 (N_13832,N_12666,N_12700);
or U13833 (N_13833,N_12574,N_12180);
nor U13834 (N_13834,N_12506,N_12386);
xnor U13835 (N_13835,N_12450,N_12302);
xnor U13836 (N_13836,N_12267,N_12324);
xnor U13837 (N_13837,N_12193,N_12528);
nor U13838 (N_13838,N_12375,N_12100);
xor U13839 (N_13839,N_12406,N_12797);
and U13840 (N_13840,N_12754,N_12802);
nand U13841 (N_13841,N_12548,N_12460);
nand U13842 (N_13842,N_12508,N_12058);
and U13843 (N_13843,N_12675,N_12301);
nand U13844 (N_13844,N_12765,N_12494);
nor U13845 (N_13845,N_12448,N_12884);
or U13846 (N_13846,N_12014,N_12106);
and U13847 (N_13847,N_12859,N_12596);
nor U13848 (N_13848,N_12449,N_12077);
nand U13849 (N_13849,N_12394,N_12951);
nor U13850 (N_13850,N_12611,N_12301);
xor U13851 (N_13851,N_12774,N_12653);
xnor U13852 (N_13852,N_12754,N_12461);
or U13853 (N_13853,N_12736,N_12438);
xnor U13854 (N_13854,N_12516,N_12182);
nor U13855 (N_13855,N_12330,N_12917);
and U13856 (N_13856,N_12300,N_12908);
or U13857 (N_13857,N_12573,N_12609);
xor U13858 (N_13858,N_12481,N_12558);
nand U13859 (N_13859,N_12511,N_12297);
nor U13860 (N_13860,N_12059,N_12433);
or U13861 (N_13861,N_12002,N_12435);
nor U13862 (N_13862,N_12407,N_12399);
or U13863 (N_13863,N_12436,N_12563);
xnor U13864 (N_13864,N_12572,N_12418);
nand U13865 (N_13865,N_12410,N_12326);
xnor U13866 (N_13866,N_12655,N_12937);
nand U13867 (N_13867,N_12085,N_12801);
and U13868 (N_13868,N_12902,N_12225);
and U13869 (N_13869,N_12479,N_12865);
and U13870 (N_13870,N_12487,N_12061);
or U13871 (N_13871,N_12393,N_12795);
or U13872 (N_13872,N_12512,N_12907);
nor U13873 (N_13873,N_12355,N_12097);
or U13874 (N_13874,N_12872,N_12940);
or U13875 (N_13875,N_12956,N_12433);
nand U13876 (N_13876,N_12304,N_12429);
and U13877 (N_13877,N_12698,N_12526);
xnor U13878 (N_13878,N_12562,N_12400);
or U13879 (N_13879,N_12587,N_12315);
or U13880 (N_13880,N_12171,N_12658);
xor U13881 (N_13881,N_12625,N_12935);
nand U13882 (N_13882,N_12744,N_12043);
nand U13883 (N_13883,N_12131,N_12902);
xor U13884 (N_13884,N_12944,N_12412);
nor U13885 (N_13885,N_12891,N_12343);
nand U13886 (N_13886,N_12360,N_12204);
nand U13887 (N_13887,N_12370,N_12512);
and U13888 (N_13888,N_12595,N_12885);
nand U13889 (N_13889,N_12453,N_12400);
nand U13890 (N_13890,N_12241,N_12475);
or U13891 (N_13891,N_12340,N_12674);
or U13892 (N_13892,N_12888,N_12507);
nor U13893 (N_13893,N_12003,N_12160);
and U13894 (N_13894,N_12803,N_12040);
and U13895 (N_13895,N_12474,N_12944);
nor U13896 (N_13896,N_12779,N_12792);
and U13897 (N_13897,N_12282,N_12172);
or U13898 (N_13898,N_12170,N_12246);
and U13899 (N_13899,N_12308,N_12488);
nor U13900 (N_13900,N_12661,N_12003);
nor U13901 (N_13901,N_12067,N_12323);
xnor U13902 (N_13902,N_12000,N_12724);
or U13903 (N_13903,N_12135,N_12231);
and U13904 (N_13904,N_12023,N_12020);
xnor U13905 (N_13905,N_12537,N_12831);
xnor U13906 (N_13906,N_12850,N_12157);
xnor U13907 (N_13907,N_12396,N_12176);
nor U13908 (N_13908,N_12039,N_12549);
nand U13909 (N_13909,N_12411,N_12362);
nor U13910 (N_13910,N_12457,N_12413);
and U13911 (N_13911,N_12442,N_12662);
nor U13912 (N_13912,N_12191,N_12860);
nor U13913 (N_13913,N_12961,N_12294);
xnor U13914 (N_13914,N_12412,N_12918);
nor U13915 (N_13915,N_12320,N_12068);
nand U13916 (N_13916,N_12947,N_12036);
or U13917 (N_13917,N_12342,N_12281);
nor U13918 (N_13918,N_12919,N_12506);
nor U13919 (N_13919,N_12867,N_12633);
xor U13920 (N_13920,N_12708,N_12533);
nor U13921 (N_13921,N_12567,N_12038);
nor U13922 (N_13922,N_12875,N_12862);
nor U13923 (N_13923,N_12261,N_12033);
xnor U13924 (N_13924,N_12892,N_12308);
xor U13925 (N_13925,N_12591,N_12217);
xnor U13926 (N_13926,N_12233,N_12501);
and U13927 (N_13927,N_12679,N_12536);
nor U13928 (N_13928,N_12237,N_12479);
nand U13929 (N_13929,N_12385,N_12104);
xnor U13930 (N_13930,N_12700,N_12074);
and U13931 (N_13931,N_12089,N_12629);
or U13932 (N_13932,N_12284,N_12860);
nor U13933 (N_13933,N_12349,N_12425);
and U13934 (N_13934,N_12840,N_12528);
nor U13935 (N_13935,N_12188,N_12169);
nand U13936 (N_13936,N_12017,N_12932);
xnor U13937 (N_13937,N_12504,N_12752);
and U13938 (N_13938,N_12540,N_12343);
and U13939 (N_13939,N_12543,N_12375);
and U13940 (N_13940,N_12184,N_12908);
and U13941 (N_13941,N_12424,N_12566);
or U13942 (N_13942,N_12931,N_12968);
or U13943 (N_13943,N_12992,N_12967);
and U13944 (N_13944,N_12401,N_12801);
or U13945 (N_13945,N_12708,N_12139);
and U13946 (N_13946,N_12968,N_12919);
nor U13947 (N_13947,N_12501,N_12437);
xnor U13948 (N_13948,N_12943,N_12302);
nor U13949 (N_13949,N_12046,N_12080);
nor U13950 (N_13950,N_12390,N_12474);
or U13951 (N_13951,N_12829,N_12312);
or U13952 (N_13952,N_12407,N_12112);
and U13953 (N_13953,N_12060,N_12727);
nor U13954 (N_13954,N_12311,N_12853);
xor U13955 (N_13955,N_12508,N_12706);
xor U13956 (N_13956,N_12953,N_12833);
xnor U13957 (N_13957,N_12812,N_12671);
nor U13958 (N_13958,N_12470,N_12529);
and U13959 (N_13959,N_12571,N_12591);
or U13960 (N_13960,N_12743,N_12292);
xor U13961 (N_13961,N_12909,N_12254);
xnor U13962 (N_13962,N_12993,N_12892);
nand U13963 (N_13963,N_12588,N_12226);
nor U13964 (N_13964,N_12825,N_12656);
xor U13965 (N_13965,N_12127,N_12826);
or U13966 (N_13966,N_12012,N_12463);
nand U13967 (N_13967,N_12580,N_12808);
xor U13968 (N_13968,N_12140,N_12864);
nand U13969 (N_13969,N_12644,N_12699);
nand U13970 (N_13970,N_12082,N_12827);
nor U13971 (N_13971,N_12032,N_12843);
nand U13972 (N_13972,N_12951,N_12215);
and U13973 (N_13973,N_12327,N_12661);
nor U13974 (N_13974,N_12811,N_12817);
xor U13975 (N_13975,N_12473,N_12171);
xor U13976 (N_13976,N_12415,N_12158);
or U13977 (N_13977,N_12800,N_12040);
nand U13978 (N_13978,N_12870,N_12329);
and U13979 (N_13979,N_12099,N_12634);
or U13980 (N_13980,N_12297,N_12587);
nor U13981 (N_13981,N_12223,N_12982);
nor U13982 (N_13982,N_12484,N_12888);
xor U13983 (N_13983,N_12342,N_12782);
nand U13984 (N_13984,N_12042,N_12628);
xor U13985 (N_13985,N_12274,N_12459);
nand U13986 (N_13986,N_12773,N_12339);
nor U13987 (N_13987,N_12312,N_12975);
or U13988 (N_13988,N_12433,N_12819);
xor U13989 (N_13989,N_12887,N_12872);
xnor U13990 (N_13990,N_12007,N_12875);
nor U13991 (N_13991,N_12149,N_12141);
nand U13992 (N_13992,N_12168,N_12528);
nor U13993 (N_13993,N_12106,N_12750);
and U13994 (N_13994,N_12987,N_12439);
or U13995 (N_13995,N_12997,N_12239);
nand U13996 (N_13996,N_12002,N_12522);
nor U13997 (N_13997,N_12603,N_12507);
or U13998 (N_13998,N_12548,N_12000);
or U13999 (N_13999,N_12751,N_12148);
or U14000 (N_14000,N_13242,N_13636);
nand U14001 (N_14001,N_13177,N_13779);
or U14002 (N_14002,N_13412,N_13154);
xnor U14003 (N_14003,N_13045,N_13228);
or U14004 (N_14004,N_13968,N_13085);
and U14005 (N_14005,N_13034,N_13068);
and U14006 (N_14006,N_13709,N_13086);
nor U14007 (N_14007,N_13274,N_13103);
or U14008 (N_14008,N_13468,N_13434);
or U14009 (N_14009,N_13815,N_13942);
nor U14010 (N_14010,N_13165,N_13006);
nor U14011 (N_14011,N_13643,N_13637);
or U14012 (N_14012,N_13837,N_13343);
xor U14013 (N_14013,N_13507,N_13748);
xor U14014 (N_14014,N_13858,N_13883);
or U14015 (N_14015,N_13078,N_13382);
xor U14016 (N_14016,N_13769,N_13459);
nand U14017 (N_14017,N_13024,N_13393);
xnor U14018 (N_14018,N_13601,N_13819);
nand U14019 (N_14019,N_13607,N_13183);
xnor U14020 (N_14020,N_13612,N_13606);
and U14021 (N_14021,N_13625,N_13480);
nand U14022 (N_14022,N_13881,N_13135);
xnor U14023 (N_14023,N_13557,N_13053);
nor U14024 (N_14024,N_13860,N_13947);
xnor U14025 (N_14025,N_13443,N_13181);
nand U14026 (N_14026,N_13953,N_13452);
nand U14027 (N_14027,N_13584,N_13221);
nand U14028 (N_14028,N_13275,N_13256);
or U14029 (N_14029,N_13658,N_13395);
xor U14030 (N_14030,N_13277,N_13499);
or U14031 (N_14031,N_13156,N_13640);
or U14032 (N_14032,N_13429,N_13717);
nand U14033 (N_14033,N_13394,N_13582);
nor U14034 (N_14034,N_13123,N_13916);
nand U14035 (N_14035,N_13014,N_13448);
nand U14036 (N_14036,N_13843,N_13767);
xnor U14037 (N_14037,N_13320,N_13080);
xnor U14038 (N_14038,N_13004,N_13096);
or U14039 (N_14039,N_13492,N_13380);
nand U14040 (N_14040,N_13617,N_13095);
or U14041 (N_14041,N_13990,N_13891);
and U14042 (N_14042,N_13983,N_13593);
or U14043 (N_14043,N_13441,N_13941);
nand U14044 (N_14044,N_13125,N_13365);
or U14045 (N_14045,N_13351,N_13759);
nand U14046 (N_14046,N_13138,N_13475);
xor U14047 (N_14047,N_13190,N_13250);
and U14048 (N_14048,N_13620,N_13110);
or U14049 (N_14049,N_13496,N_13802);
nand U14050 (N_14050,N_13806,N_13783);
nand U14051 (N_14051,N_13554,N_13733);
nand U14052 (N_14052,N_13535,N_13464);
or U14053 (N_14053,N_13513,N_13195);
xnor U14054 (N_14054,N_13244,N_13831);
nand U14055 (N_14055,N_13375,N_13400);
and U14056 (N_14056,N_13545,N_13627);
or U14057 (N_14057,N_13927,N_13101);
nand U14058 (N_14058,N_13547,N_13706);
and U14059 (N_14059,N_13703,N_13404);
and U14060 (N_14060,N_13425,N_13321);
nand U14061 (N_14061,N_13337,N_13340);
and U14062 (N_14062,N_13648,N_13057);
or U14063 (N_14063,N_13628,N_13764);
nand U14064 (N_14064,N_13901,N_13885);
nor U14065 (N_14065,N_13349,N_13234);
nand U14066 (N_14066,N_13933,N_13996);
and U14067 (N_14067,N_13911,N_13809);
xnor U14068 (N_14068,N_13174,N_13671);
or U14069 (N_14069,N_13820,N_13923);
nor U14070 (N_14070,N_13795,N_13659);
and U14071 (N_14071,N_13836,N_13962);
nor U14072 (N_14072,N_13846,N_13555);
and U14073 (N_14073,N_13909,N_13986);
xnor U14074 (N_14074,N_13192,N_13127);
xor U14075 (N_14075,N_13863,N_13598);
nand U14076 (N_14076,N_13470,N_13852);
xnor U14077 (N_14077,N_13534,N_13419);
and U14078 (N_14078,N_13610,N_13134);
nand U14079 (N_14079,N_13537,N_13835);
and U14080 (N_14080,N_13528,N_13205);
nor U14081 (N_14081,N_13295,N_13089);
nand U14082 (N_14082,N_13090,N_13976);
or U14083 (N_14083,N_13482,N_13444);
and U14084 (N_14084,N_13511,N_13245);
or U14085 (N_14085,N_13150,N_13463);
and U14086 (N_14086,N_13532,N_13278);
nor U14087 (N_14087,N_13546,N_13600);
nand U14088 (N_14088,N_13445,N_13211);
nor U14089 (N_14089,N_13818,N_13169);
and U14090 (N_14090,N_13680,N_13841);
xnor U14091 (N_14091,N_13999,N_13258);
xnor U14092 (N_14092,N_13991,N_13855);
or U14093 (N_14093,N_13253,N_13611);
nand U14094 (N_14094,N_13568,N_13196);
nor U14095 (N_14095,N_13974,N_13776);
and U14096 (N_14096,N_13410,N_13925);
nor U14097 (N_14097,N_13741,N_13294);
nor U14098 (N_14098,N_13527,N_13227);
xor U14099 (N_14099,N_13398,N_13873);
xnor U14100 (N_14100,N_13710,N_13536);
nand U14101 (N_14101,N_13426,N_13887);
xor U14102 (N_14102,N_13220,N_13893);
or U14103 (N_14103,N_13289,N_13868);
nand U14104 (N_14104,N_13170,N_13987);
nor U14105 (N_14105,N_13029,N_13414);
or U14106 (N_14106,N_13692,N_13193);
or U14107 (N_14107,N_13478,N_13094);
or U14108 (N_14108,N_13235,N_13411);
nor U14109 (N_14109,N_13564,N_13455);
or U14110 (N_14110,N_13450,N_13689);
xor U14111 (N_14111,N_13222,N_13905);
and U14112 (N_14112,N_13218,N_13039);
xnor U14113 (N_14113,N_13940,N_13629);
nor U14114 (N_14114,N_13240,N_13804);
nor U14115 (N_14115,N_13614,N_13880);
xor U14116 (N_14116,N_13063,N_13727);
or U14117 (N_14117,N_13267,N_13148);
and U14118 (N_14118,N_13072,N_13178);
or U14119 (N_14119,N_13531,N_13409);
nor U14120 (N_14120,N_13296,N_13416);
xnor U14121 (N_14121,N_13206,N_13142);
xor U14122 (N_14122,N_13615,N_13907);
and U14123 (N_14123,N_13202,N_13171);
nor U14124 (N_14124,N_13297,N_13396);
nor U14125 (N_14125,N_13525,N_13644);
or U14126 (N_14126,N_13969,N_13918);
nand U14127 (N_14127,N_13229,N_13702);
nor U14128 (N_14128,N_13265,N_13377);
xor U14129 (N_14129,N_13930,N_13383);
and U14130 (N_14130,N_13001,N_13675);
and U14131 (N_14131,N_13575,N_13862);
nand U14132 (N_14132,N_13427,N_13924);
xor U14133 (N_14133,N_13867,N_13803);
nor U14134 (N_14134,N_13008,N_13097);
and U14135 (N_14135,N_13782,N_13403);
xnor U14136 (N_14136,N_13116,N_13257);
xor U14137 (N_14137,N_13826,N_13965);
xnor U14138 (N_14138,N_13255,N_13466);
nor U14139 (N_14139,N_13037,N_13808);
xor U14140 (N_14140,N_13543,N_13254);
nand U14141 (N_14141,N_13269,N_13904);
and U14142 (N_14142,N_13318,N_13332);
xor U14143 (N_14143,N_13370,N_13460);
nor U14144 (N_14144,N_13609,N_13500);
nor U14145 (N_14145,N_13203,N_13249);
nand U14146 (N_14146,N_13736,N_13864);
or U14147 (N_14147,N_13757,N_13437);
and U14148 (N_14148,N_13363,N_13345);
nand U14149 (N_14149,N_13408,N_13739);
nor U14150 (N_14150,N_13216,N_13955);
and U14151 (N_14151,N_13019,N_13565);
and U14152 (N_14152,N_13642,N_13457);
or U14153 (N_14153,N_13728,N_13280);
xnor U14154 (N_14154,N_13538,N_13824);
xor U14155 (N_14155,N_13071,N_13886);
nand U14156 (N_14156,N_13497,N_13752);
xnor U14157 (N_14157,N_13786,N_13963);
or U14158 (N_14158,N_13422,N_13632);
xor U14159 (N_14159,N_13921,N_13721);
nor U14160 (N_14160,N_13672,N_13998);
nand U14161 (N_14161,N_13260,N_13099);
nor U14162 (N_14162,N_13477,N_13239);
and U14163 (N_14163,N_13505,N_13413);
xnor U14164 (N_14164,N_13719,N_13122);
and U14165 (N_14165,N_13934,N_13981);
nor U14166 (N_14166,N_13281,N_13420);
xnor U14167 (N_14167,N_13041,N_13327);
or U14168 (N_14168,N_13772,N_13453);
xnor U14169 (N_14169,N_13185,N_13027);
or U14170 (N_14170,N_13487,N_13483);
and U14171 (N_14171,N_13421,N_13028);
or U14172 (N_14172,N_13677,N_13111);
or U14173 (N_14173,N_13773,N_13679);
and U14174 (N_14174,N_13491,N_13875);
xnor U14175 (N_14175,N_13724,N_13010);
and U14176 (N_14176,N_13032,N_13775);
or U14177 (N_14177,N_13553,N_13261);
and U14178 (N_14178,N_13417,N_13428);
and U14179 (N_14179,N_13081,N_13336);
xnor U14180 (N_14180,N_13950,N_13931);
nor U14181 (N_14181,N_13451,N_13179);
xnor U14182 (N_14182,N_13124,N_13397);
nor U14183 (N_14183,N_13816,N_13023);
or U14184 (N_14184,N_13026,N_13005);
or U14185 (N_14185,N_13742,N_13108);
nor U14186 (N_14186,N_13935,N_13760);
and U14187 (N_14187,N_13523,N_13722);
and U14188 (N_14188,N_13517,N_13884);
nor U14189 (N_14189,N_13133,N_13360);
nor U14190 (N_14190,N_13530,N_13371);
or U14191 (N_14191,N_13364,N_13781);
nand U14192 (N_14192,N_13621,N_13346);
and U14193 (N_14193,N_13376,N_13339);
xnor U14194 (N_14194,N_13272,N_13882);
and U14195 (N_14195,N_13390,N_13871);
and U14196 (N_14196,N_13472,N_13687);
nor U14197 (N_14197,N_13755,N_13697);
or U14198 (N_14198,N_13812,N_13303);
or U14199 (N_14199,N_13385,N_13874);
or U14200 (N_14200,N_13995,N_13715);
and U14201 (N_14201,N_13971,N_13763);
nand U14202 (N_14202,N_13287,N_13391);
xnor U14203 (N_14203,N_13853,N_13599);
nand U14204 (N_14204,N_13797,N_13114);
and U14205 (N_14205,N_13624,N_13811);
xnor U14206 (N_14206,N_13288,N_13681);
xor U14207 (N_14207,N_13569,N_13248);
nand U14208 (N_14208,N_13007,N_13054);
or U14209 (N_14209,N_13838,N_13619);
nand U14210 (N_14210,N_13857,N_13978);
nor U14211 (N_14211,N_13237,N_13246);
xor U14212 (N_14212,N_13159,N_13481);
xor U14213 (N_14213,N_13737,N_13056);
xnor U14214 (N_14214,N_13092,N_13262);
or U14215 (N_14215,N_13328,N_13333);
xor U14216 (N_14216,N_13866,N_13731);
nand U14217 (N_14217,N_13319,N_13276);
and U14218 (N_14218,N_13641,N_13406);
nor U14219 (N_14219,N_13347,N_13194);
nor U14220 (N_14220,N_13259,N_13059);
nor U14221 (N_14221,N_13791,N_13524);
nand U14222 (N_14222,N_13018,N_13247);
or U14223 (N_14223,N_13566,N_13407);
nor U14224 (N_14224,N_13372,N_13577);
nor U14225 (N_14225,N_13512,N_13898);
xnor U14226 (N_14226,N_13152,N_13330);
nor U14227 (N_14227,N_13967,N_13009);
or U14228 (N_14228,N_13839,N_13042);
xor U14229 (N_14229,N_13794,N_13494);
nand U14230 (N_14230,N_13653,N_13338);
and U14231 (N_14231,N_13979,N_13226);
and U14232 (N_14232,N_13712,N_13115);
nor U14233 (N_14233,N_13851,N_13186);
or U14234 (N_14234,N_13065,N_13827);
xnor U14235 (N_14235,N_13066,N_13798);
nand U14236 (N_14236,N_13305,N_13630);
nand U14237 (N_14237,N_13163,N_13574);
or U14238 (N_14238,N_13424,N_13521);
and U14239 (N_14239,N_13489,N_13430);
nor U14240 (N_14240,N_13075,N_13673);
xnor U14241 (N_14241,N_13369,N_13572);
nor U14242 (N_14242,N_13243,N_13067);
nand U14243 (N_14243,N_13106,N_13334);
and U14244 (N_14244,N_13490,N_13929);
and U14245 (N_14245,N_13622,N_13501);
xnor U14246 (N_14246,N_13777,N_13964);
and U14247 (N_14247,N_13432,N_13188);
nand U14248 (N_14248,N_13015,N_13074);
xor U14249 (N_14249,N_13449,N_13633);
nor U14250 (N_14250,N_13310,N_13355);
or U14251 (N_14251,N_13268,N_13645);
nor U14252 (N_14252,N_13718,N_13936);
nand U14253 (N_14253,N_13581,N_13635);
and U14254 (N_14254,N_13879,N_13693);
xor U14255 (N_14255,N_13686,N_13102);
nand U14256 (N_14256,N_13638,N_13785);
nand U14257 (N_14257,N_13842,N_13302);
xor U14258 (N_14258,N_13354,N_13676);
nor U14259 (N_14259,N_13168,N_13506);
nand U14260 (N_14260,N_13442,N_13002);
or U14261 (N_14261,N_13823,N_13113);
or U14262 (N_14262,N_13859,N_13164);
nand U14263 (N_14263,N_13865,N_13016);
and U14264 (N_14264,N_13588,N_13603);
nand U14265 (N_14265,N_13145,N_13022);
xnor U14266 (N_14266,N_13939,N_13402);
nand U14267 (N_14267,N_13896,N_13469);
or U14268 (N_14268,N_13548,N_13960);
and U14269 (N_14269,N_13201,N_13596);
xor U14270 (N_14270,N_13342,N_13052);
nor U14271 (N_14271,N_13198,N_13064);
and U14272 (N_14272,N_13465,N_13570);
or U14273 (N_14273,N_13307,N_13112);
or U14274 (N_14274,N_13932,N_13695);
xnor U14275 (N_14275,N_13314,N_13821);
and U14276 (N_14276,N_13701,N_13273);
nor U14277 (N_14277,N_13230,N_13539);
and U14278 (N_14278,N_13694,N_13146);
and U14279 (N_14279,N_13583,N_13540);
nor U14280 (N_14280,N_13848,N_13560);
xnor U14281 (N_14281,N_13730,N_13176);
nand U14282 (N_14282,N_13980,N_13691);
and U14283 (N_14283,N_13415,N_13439);
and U14284 (N_14284,N_13224,N_13605);
or U14285 (N_14285,N_13660,N_13304);
nand U14286 (N_14286,N_13219,N_13038);
nor U14287 (N_14287,N_13914,N_13667);
xor U14288 (N_14288,N_13761,N_13126);
nor U14289 (N_14289,N_13132,N_13571);
nor U14290 (N_14290,N_13140,N_13750);
and U14291 (N_14291,N_13479,N_13503);
nor U14292 (N_14292,N_13647,N_13559);
xor U14293 (N_14293,N_13191,N_13668);
nand U14294 (N_14294,N_13073,N_13051);
and U14295 (N_14295,N_13822,N_13985);
nor U14296 (N_14296,N_13509,N_13817);
xor U14297 (N_14297,N_13952,N_13335);
nand U14298 (N_14298,N_13814,N_13738);
xnor U14299 (N_14299,N_13043,N_13292);
or U14300 (N_14300,N_13590,N_13184);
nor U14301 (N_14301,N_13845,N_13118);
xor U14302 (N_14302,N_13341,N_13768);
or U14303 (N_14303,N_13199,N_13972);
and U14304 (N_14304,N_13661,N_13943);
nand U14305 (N_14305,N_13060,N_13498);
xnor U14306 (N_14306,N_13913,N_13740);
xor U14307 (N_14307,N_13549,N_13604);
or U14308 (N_14308,N_13747,N_13754);
nor U14309 (N_14309,N_13495,N_13849);
nor U14310 (N_14310,N_13107,N_13084);
nand U14311 (N_14311,N_13353,N_13079);
nor U14312 (N_14312,N_13088,N_13121);
or U14313 (N_14313,N_13238,N_13161);
and U14314 (N_14314,N_13561,N_13308);
xor U14315 (N_14315,N_13970,N_13563);
or U14316 (N_14316,N_13670,N_13129);
or U14317 (N_14317,N_13994,N_13374);
and U14318 (N_14318,N_13362,N_13473);
nor U14319 (N_14319,N_13889,N_13172);
nor U14320 (N_14320,N_13350,N_13988);
and U14321 (N_14321,N_13324,N_13279);
xnor U14322 (N_14322,N_13306,N_13580);
nor U14323 (N_14323,N_13180,N_13562);
nand U14324 (N_14324,N_13799,N_13046);
and U14325 (N_14325,N_13358,N_13387);
or U14326 (N_14326,N_13945,N_13519);
or U14327 (N_14327,N_13418,N_13212);
xnor U14328 (N_14328,N_13602,N_13241);
nor U14329 (N_14329,N_13392,N_13937);
nand U14330 (N_14330,N_13825,N_13231);
or U14331 (N_14331,N_13698,N_13800);
or U14332 (N_14332,N_13151,N_13894);
nor U14333 (N_14333,N_13213,N_13440);
nand U14334 (N_14334,N_13993,N_13682);
nand U14335 (N_14335,N_13771,N_13688);
nor U14336 (N_14336,N_13232,N_13951);
xor U14337 (N_14337,N_13264,N_13368);
and U14338 (N_14338,N_13888,N_13616);
and U14339 (N_14339,N_13109,N_13446);
or U14340 (N_14340,N_13902,N_13013);
or U14341 (N_14341,N_13098,N_13542);
and U14342 (N_14342,N_13585,N_13379);
and U14343 (N_14343,N_13147,N_13699);
nand U14344 (N_14344,N_13801,N_13117);
nor U14345 (N_14345,N_13522,N_13309);
nand U14346 (N_14346,N_13725,N_13646);
and U14347 (N_14347,N_13832,N_13726);
xor U14348 (N_14348,N_13591,N_13083);
xnor U14349 (N_14349,N_13317,N_13788);
xnor U14350 (N_14350,N_13664,N_13510);
xor U14351 (N_14351,N_13665,N_13723);
xor U14352 (N_14352,N_13579,N_13946);
and U14353 (N_14353,N_13313,N_13137);
xnor U14354 (N_14354,N_13926,N_13251);
nor U14355 (N_14355,N_13631,N_13751);
or U14356 (N_14356,N_13100,N_13529);
and U14357 (N_14357,N_13977,N_13223);
xor U14358 (N_14358,N_13910,N_13020);
nor U14359 (N_14359,N_13716,N_13683);
and U14360 (N_14360,N_13705,N_13903);
nand U14361 (N_14361,N_13650,N_13533);
xor U14362 (N_14362,N_13870,N_13618);
nand U14363 (N_14363,N_13356,N_13966);
nor U14364 (N_14364,N_13070,N_13160);
xnor U14365 (N_14365,N_13055,N_13869);
xor U14366 (N_14366,N_13373,N_13131);
nor U14367 (N_14367,N_13649,N_13899);
and U14368 (N_14368,N_13476,N_13919);
xnor U14369 (N_14369,N_13187,N_13743);
and U14370 (N_14370,N_13040,N_13587);
or U14371 (N_14371,N_13141,N_13669);
and U14372 (N_14372,N_13366,N_13435);
nand U14373 (N_14373,N_13576,N_13592);
or U14374 (N_14374,N_13556,N_13711);
nand U14375 (N_14375,N_13105,N_13854);
and U14376 (N_14376,N_13290,N_13447);
and U14377 (N_14377,N_13149,N_13613);
or U14378 (N_14378,N_13878,N_13384);
xnor U14379 (N_14379,N_13762,N_13516);
nand U14380 (N_14380,N_13595,N_13745);
or U14381 (N_14381,N_13770,N_13182);
or U14382 (N_14382,N_13900,N_13423);
nand U14383 (N_14383,N_13158,N_13805);
and U14384 (N_14384,N_13299,N_13961);
nand U14385 (N_14385,N_13957,N_13329);
and U14386 (N_14386,N_13634,N_13544);
xnor U14387 (N_14387,N_13714,N_13550);
nand U14388 (N_14388,N_13657,N_13285);
and U14389 (N_14389,N_13597,N_13515);
xor U14390 (N_14390,N_13352,N_13359);
xor U14391 (N_14391,N_13486,N_13061);
xnor U14392 (N_14392,N_13077,N_13796);
nor U14393 (N_14393,N_13120,N_13992);
xor U14394 (N_14394,N_13959,N_13076);
nand U14395 (N_14395,N_13144,N_13514);
nor U14396 (N_14396,N_13401,N_13922);
nor U14397 (N_14397,N_13944,N_13143);
nor U14398 (N_14398,N_13069,N_13300);
xor U14399 (N_14399,N_13488,N_13948);
nand U14400 (N_14400,N_13003,N_13856);
or U14401 (N_14401,N_13485,N_13734);
xnor U14402 (N_14402,N_13789,N_13793);
nor U14403 (N_14403,N_13508,N_13233);
nand U14404 (N_14404,N_13685,N_13104);
nand U14405 (N_14405,N_13093,N_13062);
or U14406 (N_14406,N_13316,N_13284);
nor U14407 (N_14407,N_13312,N_13036);
or U14408 (N_14408,N_13048,N_13674);
or U14409 (N_14409,N_13892,N_13784);
nand U14410 (N_14410,N_13830,N_13058);
and U14411 (N_14411,N_13541,N_13850);
xor U14412 (N_14412,N_13700,N_13438);
and U14413 (N_14413,N_13890,N_13928);
and U14414 (N_14414,N_13917,N_13984);
nand U14415 (N_14415,N_13087,N_13436);
or U14416 (N_14416,N_13139,N_13707);
or U14417 (N_14417,N_13197,N_13774);
and U14418 (N_14418,N_13807,N_13467);
and U14419 (N_14419,N_13044,N_13348);
or U14420 (N_14420,N_13756,N_13047);
and U14421 (N_14421,N_13997,N_13204);
nand U14422 (N_14422,N_13626,N_13502);
and U14423 (N_14423,N_13749,N_13678);
and U14424 (N_14424,N_13526,N_13704);
or U14425 (N_14425,N_13958,N_13908);
nor U14426 (N_14426,N_13652,N_13035);
or U14427 (N_14427,N_13214,N_13000);
nand U14428 (N_14428,N_13291,N_13357);
nand U14429 (N_14429,N_13847,N_13623);
nand U14430 (N_14430,N_13298,N_13225);
nor U14431 (N_14431,N_13753,N_13270);
or U14432 (N_14432,N_13315,N_13252);
nor U14433 (N_14433,N_13662,N_13033);
xnor U14434 (N_14434,N_13323,N_13130);
xor U14435 (N_14435,N_13829,N_13973);
and U14436 (N_14436,N_13790,N_13031);
nand U14437 (N_14437,N_13167,N_13573);
nand U14438 (N_14438,N_13949,N_13840);
and U14439 (N_14439,N_13558,N_13200);
nor U14440 (N_14440,N_13518,N_13266);
or U14441 (N_14441,N_13344,N_13938);
or U14442 (N_14442,N_13906,N_13861);
and U14443 (N_14443,N_13325,N_13666);
or U14444 (N_14444,N_13552,N_13732);
and U14445 (N_14445,N_13283,N_13975);
nand U14446 (N_14446,N_13895,N_13690);
nor U14447 (N_14447,N_13025,N_13876);
nand U14448 (N_14448,N_13388,N_13454);
nor U14449 (N_14449,N_13157,N_13217);
or U14450 (N_14450,N_13386,N_13173);
xnor U14451 (N_14451,N_13431,N_13215);
and U14452 (N_14452,N_13461,N_13735);
nand U14453 (N_14453,N_13684,N_13920);
nor U14454 (N_14454,N_13810,N_13663);
and U14455 (N_14455,N_13162,N_13136);
or U14456 (N_14456,N_13520,N_13282);
nor U14457 (N_14457,N_13456,N_13766);
nand U14458 (N_14458,N_13017,N_13049);
and U14459 (N_14459,N_13236,N_13208);
or U14460 (N_14460,N_13897,N_13271);
nor U14461 (N_14461,N_13746,N_13639);
xor U14462 (N_14462,N_13030,N_13912);
and U14463 (N_14463,N_13872,N_13433);
xor U14464 (N_14464,N_13493,N_13050);
nand U14465 (N_14465,N_13462,N_13378);
or U14466 (N_14466,N_13119,N_13331);
or U14467 (N_14467,N_13458,N_13210);
nand U14468 (N_14468,N_13578,N_13322);
and U14469 (N_14469,N_13361,N_13091);
xor U14470 (N_14470,N_13155,N_13209);
xor U14471 (N_14471,N_13082,N_13877);
or U14472 (N_14472,N_13651,N_13915);
or U14473 (N_14473,N_13813,N_13567);
xor U14474 (N_14474,N_13021,N_13982);
xor U14475 (N_14475,N_13311,N_13399);
nor U14476 (N_14476,N_13778,N_13828);
and U14477 (N_14477,N_13654,N_13608);
and U14478 (N_14478,N_13787,N_13474);
xnor U14479 (N_14479,N_13765,N_13833);
nand U14480 (N_14480,N_13286,N_13484);
nor U14481 (N_14481,N_13128,N_13708);
and U14482 (N_14482,N_13189,N_13586);
xor U14483 (N_14483,N_13989,N_13471);
nand U14484 (N_14484,N_13263,N_13956);
and U14485 (N_14485,N_13153,N_13720);
xor U14486 (N_14486,N_13834,N_13326);
or U14487 (N_14487,N_13844,N_13954);
nand U14488 (N_14488,N_13713,N_13293);
or U14489 (N_14489,N_13166,N_13792);
nor U14490 (N_14490,N_13729,N_13207);
xor U14491 (N_14491,N_13367,N_13594);
and U14492 (N_14492,N_13744,N_13504);
and U14493 (N_14493,N_13758,N_13780);
or U14494 (N_14494,N_13389,N_13011);
nor U14495 (N_14495,N_13381,N_13301);
and U14496 (N_14496,N_13589,N_13656);
and U14497 (N_14497,N_13175,N_13405);
and U14498 (N_14498,N_13551,N_13012);
or U14499 (N_14499,N_13696,N_13655);
nor U14500 (N_14500,N_13194,N_13713);
nand U14501 (N_14501,N_13312,N_13149);
nor U14502 (N_14502,N_13472,N_13393);
and U14503 (N_14503,N_13752,N_13836);
or U14504 (N_14504,N_13620,N_13494);
xor U14505 (N_14505,N_13527,N_13535);
or U14506 (N_14506,N_13241,N_13899);
xnor U14507 (N_14507,N_13137,N_13098);
nand U14508 (N_14508,N_13688,N_13267);
nor U14509 (N_14509,N_13619,N_13460);
and U14510 (N_14510,N_13561,N_13261);
and U14511 (N_14511,N_13920,N_13685);
xnor U14512 (N_14512,N_13838,N_13759);
and U14513 (N_14513,N_13897,N_13778);
nand U14514 (N_14514,N_13629,N_13342);
nand U14515 (N_14515,N_13487,N_13322);
and U14516 (N_14516,N_13579,N_13607);
or U14517 (N_14517,N_13116,N_13956);
and U14518 (N_14518,N_13307,N_13702);
or U14519 (N_14519,N_13401,N_13054);
xor U14520 (N_14520,N_13989,N_13082);
and U14521 (N_14521,N_13062,N_13747);
nand U14522 (N_14522,N_13047,N_13917);
nor U14523 (N_14523,N_13215,N_13691);
xnor U14524 (N_14524,N_13104,N_13048);
or U14525 (N_14525,N_13019,N_13536);
nand U14526 (N_14526,N_13399,N_13576);
nor U14527 (N_14527,N_13516,N_13447);
nor U14528 (N_14528,N_13981,N_13374);
or U14529 (N_14529,N_13651,N_13201);
nor U14530 (N_14530,N_13080,N_13477);
nand U14531 (N_14531,N_13976,N_13262);
nand U14532 (N_14532,N_13580,N_13444);
and U14533 (N_14533,N_13483,N_13531);
and U14534 (N_14534,N_13441,N_13740);
nand U14535 (N_14535,N_13216,N_13934);
or U14536 (N_14536,N_13717,N_13995);
or U14537 (N_14537,N_13128,N_13636);
and U14538 (N_14538,N_13242,N_13231);
nor U14539 (N_14539,N_13619,N_13075);
nor U14540 (N_14540,N_13155,N_13201);
xor U14541 (N_14541,N_13624,N_13755);
and U14542 (N_14542,N_13481,N_13166);
and U14543 (N_14543,N_13140,N_13449);
nor U14544 (N_14544,N_13276,N_13806);
nand U14545 (N_14545,N_13666,N_13802);
or U14546 (N_14546,N_13646,N_13412);
xnor U14547 (N_14547,N_13703,N_13642);
and U14548 (N_14548,N_13387,N_13564);
xnor U14549 (N_14549,N_13716,N_13868);
and U14550 (N_14550,N_13811,N_13004);
nor U14551 (N_14551,N_13014,N_13848);
xnor U14552 (N_14552,N_13155,N_13609);
nor U14553 (N_14553,N_13072,N_13526);
or U14554 (N_14554,N_13190,N_13815);
nand U14555 (N_14555,N_13743,N_13410);
and U14556 (N_14556,N_13466,N_13594);
nand U14557 (N_14557,N_13121,N_13072);
nor U14558 (N_14558,N_13755,N_13193);
or U14559 (N_14559,N_13352,N_13598);
or U14560 (N_14560,N_13596,N_13565);
xor U14561 (N_14561,N_13953,N_13711);
or U14562 (N_14562,N_13847,N_13932);
or U14563 (N_14563,N_13048,N_13384);
nor U14564 (N_14564,N_13038,N_13084);
and U14565 (N_14565,N_13751,N_13470);
or U14566 (N_14566,N_13435,N_13500);
nand U14567 (N_14567,N_13709,N_13353);
or U14568 (N_14568,N_13669,N_13076);
nor U14569 (N_14569,N_13227,N_13397);
and U14570 (N_14570,N_13743,N_13163);
or U14571 (N_14571,N_13381,N_13743);
nand U14572 (N_14572,N_13357,N_13349);
nand U14573 (N_14573,N_13440,N_13384);
nor U14574 (N_14574,N_13102,N_13365);
or U14575 (N_14575,N_13986,N_13044);
and U14576 (N_14576,N_13021,N_13423);
xnor U14577 (N_14577,N_13676,N_13254);
nor U14578 (N_14578,N_13539,N_13838);
xor U14579 (N_14579,N_13738,N_13655);
nor U14580 (N_14580,N_13925,N_13417);
or U14581 (N_14581,N_13604,N_13873);
nor U14582 (N_14582,N_13052,N_13063);
nor U14583 (N_14583,N_13301,N_13001);
xor U14584 (N_14584,N_13709,N_13923);
or U14585 (N_14585,N_13216,N_13990);
xnor U14586 (N_14586,N_13346,N_13217);
or U14587 (N_14587,N_13472,N_13779);
nor U14588 (N_14588,N_13612,N_13018);
and U14589 (N_14589,N_13773,N_13811);
nand U14590 (N_14590,N_13834,N_13220);
xnor U14591 (N_14591,N_13881,N_13461);
or U14592 (N_14592,N_13279,N_13869);
nor U14593 (N_14593,N_13350,N_13910);
xnor U14594 (N_14594,N_13300,N_13380);
xor U14595 (N_14595,N_13007,N_13243);
and U14596 (N_14596,N_13112,N_13159);
and U14597 (N_14597,N_13996,N_13768);
xor U14598 (N_14598,N_13538,N_13279);
nor U14599 (N_14599,N_13305,N_13841);
and U14600 (N_14600,N_13817,N_13197);
nor U14601 (N_14601,N_13268,N_13703);
nand U14602 (N_14602,N_13905,N_13750);
and U14603 (N_14603,N_13847,N_13737);
nand U14604 (N_14604,N_13373,N_13494);
xnor U14605 (N_14605,N_13246,N_13111);
or U14606 (N_14606,N_13907,N_13412);
or U14607 (N_14607,N_13228,N_13402);
xor U14608 (N_14608,N_13279,N_13212);
nor U14609 (N_14609,N_13112,N_13319);
nand U14610 (N_14610,N_13802,N_13160);
nand U14611 (N_14611,N_13392,N_13167);
nor U14612 (N_14612,N_13845,N_13347);
nand U14613 (N_14613,N_13427,N_13866);
nor U14614 (N_14614,N_13709,N_13200);
nand U14615 (N_14615,N_13325,N_13939);
nor U14616 (N_14616,N_13114,N_13336);
and U14617 (N_14617,N_13202,N_13058);
nor U14618 (N_14618,N_13367,N_13024);
or U14619 (N_14619,N_13551,N_13260);
nand U14620 (N_14620,N_13350,N_13308);
and U14621 (N_14621,N_13621,N_13565);
nand U14622 (N_14622,N_13816,N_13154);
nor U14623 (N_14623,N_13043,N_13081);
or U14624 (N_14624,N_13119,N_13028);
or U14625 (N_14625,N_13270,N_13202);
nor U14626 (N_14626,N_13076,N_13284);
xnor U14627 (N_14627,N_13952,N_13575);
and U14628 (N_14628,N_13122,N_13017);
xnor U14629 (N_14629,N_13406,N_13731);
and U14630 (N_14630,N_13350,N_13778);
and U14631 (N_14631,N_13314,N_13768);
nor U14632 (N_14632,N_13230,N_13061);
xnor U14633 (N_14633,N_13850,N_13588);
xnor U14634 (N_14634,N_13247,N_13804);
xor U14635 (N_14635,N_13338,N_13507);
nand U14636 (N_14636,N_13918,N_13651);
or U14637 (N_14637,N_13434,N_13917);
nor U14638 (N_14638,N_13404,N_13141);
nor U14639 (N_14639,N_13839,N_13186);
xnor U14640 (N_14640,N_13479,N_13259);
or U14641 (N_14641,N_13430,N_13572);
or U14642 (N_14642,N_13395,N_13206);
nor U14643 (N_14643,N_13258,N_13613);
nor U14644 (N_14644,N_13346,N_13731);
xnor U14645 (N_14645,N_13578,N_13686);
and U14646 (N_14646,N_13239,N_13119);
xnor U14647 (N_14647,N_13669,N_13004);
nor U14648 (N_14648,N_13951,N_13583);
nor U14649 (N_14649,N_13385,N_13132);
or U14650 (N_14650,N_13073,N_13980);
or U14651 (N_14651,N_13515,N_13332);
or U14652 (N_14652,N_13545,N_13359);
xor U14653 (N_14653,N_13199,N_13346);
or U14654 (N_14654,N_13113,N_13322);
or U14655 (N_14655,N_13237,N_13212);
or U14656 (N_14656,N_13658,N_13322);
or U14657 (N_14657,N_13002,N_13644);
or U14658 (N_14658,N_13399,N_13874);
and U14659 (N_14659,N_13380,N_13818);
or U14660 (N_14660,N_13037,N_13768);
xnor U14661 (N_14661,N_13856,N_13459);
or U14662 (N_14662,N_13301,N_13722);
xnor U14663 (N_14663,N_13728,N_13477);
nand U14664 (N_14664,N_13446,N_13867);
nor U14665 (N_14665,N_13295,N_13104);
nand U14666 (N_14666,N_13363,N_13301);
or U14667 (N_14667,N_13668,N_13407);
and U14668 (N_14668,N_13685,N_13554);
nor U14669 (N_14669,N_13567,N_13735);
nand U14670 (N_14670,N_13762,N_13989);
xnor U14671 (N_14671,N_13805,N_13354);
nand U14672 (N_14672,N_13598,N_13888);
nand U14673 (N_14673,N_13411,N_13902);
and U14674 (N_14674,N_13820,N_13359);
and U14675 (N_14675,N_13357,N_13530);
nor U14676 (N_14676,N_13266,N_13675);
nor U14677 (N_14677,N_13638,N_13148);
nand U14678 (N_14678,N_13692,N_13633);
nor U14679 (N_14679,N_13269,N_13612);
or U14680 (N_14680,N_13436,N_13609);
xnor U14681 (N_14681,N_13773,N_13817);
and U14682 (N_14682,N_13860,N_13530);
and U14683 (N_14683,N_13091,N_13386);
nor U14684 (N_14684,N_13920,N_13866);
or U14685 (N_14685,N_13425,N_13914);
xor U14686 (N_14686,N_13563,N_13314);
nor U14687 (N_14687,N_13004,N_13939);
and U14688 (N_14688,N_13611,N_13426);
nand U14689 (N_14689,N_13491,N_13549);
xnor U14690 (N_14690,N_13321,N_13998);
or U14691 (N_14691,N_13778,N_13978);
nand U14692 (N_14692,N_13454,N_13673);
nor U14693 (N_14693,N_13908,N_13993);
nand U14694 (N_14694,N_13628,N_13391);
or U14695 (N_14695,N_13788,N_13203);
or U14696 (N_14696,N_13955,N_13989);
nand U14697 (N_14697,N_13971,N_13080);
xnor U14698 (N_14698,N_13582,N_13874);
nand U14699 (N_14699,N_13229,N_13576);
and U14700 (N_14700,N_13657,N_13099);
or U14701 (N_14701,N_13868,N_13741);
nor U14702 (N_14702,N_13242,N_13380);
or U14703 (N_14703,N_13753,N_13006);
nand U14704 (N_14704,N_13152,N_13338);
or U14705 (N_14705,N_13425,N_13677);
and U14706 (N_14706,N_13766,N_13779);
nor U14707 (N_14707,N_13639,N_13915);
nand U14708 (N_14708,N_13218,N_13845);
xnor U14709 (N_14709,N_13063,N_13894);
nand U14710 (N_14710,N_13314,N_13499);
nor U14711 (N_14711,N_13243,N_13270);
and U14712 (N_14712,N_13228,N_13374);
or U14713 (N_14713,N_13097,N_13000);
nand U14714 (N_14714,N_13860,N_13170);
nand U14715 (N_14715,N_13643,N_13676);
or U14716 (N_14716,N_13193,N_13469);
xor U14717 (N_14717,N_13300,N_13800);
nor U14718 (N_14718,N_13588,N_13484);
xnor U14719 (N_14719,N_13363,N_13774);
and U14720 (N_14720,N_13869,N_13206);
or U14721 (N_14721,N_13356,N_13763);
and U14722 (N_14722,N_13647,N_13951);
nand U14723 (N_14723,N_13702,N_13725);
or U14724 (N_14724,N_13975,N_13437);
or U14725 (N_14725,N_13730,N_13750);
xor U14726 (N_14726,N_13162,N_13237);
and U14727 (N_14727,N_13558,N_13133);
xor U14728 (N_14728,N_13691,N_13091);
xnor U14729 (N_14729,N_13433,N_13940);
nand U14730 (N_14730,N_13857,N_13976);
xor U14731 (N_14731,N_13944,N_13359);
xnor U14732 (N_14732,N_13508,N_13246);
nand U14733 (N_14733,N_13074,N_13417);
and U14734 (N_14734,N_13033,N_13160);
nand U14735 (N_14735,N_13976,N_13029);
xnor U14736 (N_14736,N_13548,N_13123);
nand U14737 (N_14737,N_13621,N_13253);
nor U14738 (N_14738,N_13598,N_13961);
or U14739 (N_14739,N_13359,N_13538);
and U14740 (N_14740,N_13865,N_13653);
and U14741 (N_14741,N_13645,N_13109);
or U14742 (N_14742,N_13222,N_13814);
nand U14743 (N_14743,N_13208,N_13478);
or U14744 (N_14744,N_13540,N_13104);
or U14745 (N_14745,N_13564,N_13958);
nor U14746 (N_14746,N_13130,N_13616);
nor U14747 (N_14747,N_13277,N_13594);
or U14748 (N_14748,N_13174,N_13811);
nand U14749 (N_14749,N_13735,N_13297);
nand U14750 (N_14750,N_13916,N_13576);
nand U14751 (N_14751,N_13456,N_13989);
nor U14752 (N_14752,N_13983,N_13616);
nand U14753 (N_14753,N_13019,N_13637);
or U14754 (N_14754,N_13657,N_13166);
nand U14755 (N_14755,N_13885,N_13344);
nand U14756 (N_14756,N_13067,N_13529);
and U14757 (N_14757,N_13263,N_13450);
or U14758 (N_14758,N_13866,N_13965);
xnor U14759 (N_14759,N_13712,N_13330);
nor U14760 (N_14760,N_13984,N_13157);
xnor U14761 (N_14761,N_13527,N_13875);
xnor U14762 (N_14762,N_13689,N_13785);
xor U14763 (N_14763,N_13383,N_13911);
and U14764 (N_14764,N_13269,N_13842);
nand U14765 (N_14765,N_13296,N_13644);
xnor U14766 (N_14766,N_13606,N_13870);
and U14767 (N_14767,N_13591,N_13116);
nor U14768 (N_14768,N_13931,N_13862);
or U14769 (N_14769,N_13533,N_13426);
or U14770 (N_14770,N_13343,N_13889);
nand U14771 (N_14771,N_13203,N_13041);
xnor U14772 (N_14772,N_13021,N_13118);
nand U14773 (N_14773,N_13519,N_13674);
nand U14774 (N_14774,N_13889,N_13183);
nand U14775 (N_14775,N_13751,N_13065);
or U14776 (N_14776,N_13632,N_13369);
or U14777 (N_14777,N_13694,N_13809);
xnor U14778 (N_14778,N_13967,N_13510);
nand U14779 (N_14779,N_13370,N_13277);
or U14780 (N_14780,N_13014,N_13538);
or U14781 (N_14781,N_13491,N_13252);
or U14782 (N_14782,N_13997,N_13052);
xor U14783 (N_14783,N_13733,N_13922);
nor U14784 (N_14784,N_13960,N_13196);
or U14785 (N_14785,N_13489,N_13807);
nor U14786 (N_14786,N_13298,N_13649);
nand U14787 (N_14787,N_13186,N_13938);
or U14788 (N_14788,N_13609,N_13538);
nor U14789 (N_14789,N_13407,N_13155);
nand U14790 (N_14790,N_13917,N_13040);
xnor U14791 (N_14791,N_13840,N_13200);
nand U14792 (N_14792,N_13045,N_13503);
or U14793 (N_14793,N_13385,N_13673);
xnor U14794 (N_14794,N_13285,N_13216);
and U14795 (N_14795,N_13598,N_13331);
nor U14796 (N_14796,N_13261,N_13837);
or U14797 (N_14797,N_13143,N_13945);
and U14798 (N_14798,N_13656,N_13793);
nor U14799 (N_14799,N_13728,N_13116);
and U14800 (N_14800,N_13674,N_13709);
nand U14801 (N_14801,N_13916,N_13513);
and U14802 (N_14802,N_13388,N_13881);
or U14803 (N_14803,N_13041,N_13466);
nand U14804 (N_14804,N_13290,N_13136);
nor U14805 (N_14805,N_13562,N_13902);
nor U14806 (N_14806,N_13480,N_13403);
nor U14807 (N_14807,N_13780,N_13922);
nor U14808 (N_14808,N_13470,N_13083);
nor U14809 (N_14809,N_13329,N_13680);
or U14810 (N_14810,N_13903,N_13668);
nor U14811 (N_14811,N_13712,N_13033);
and U14812 (N_14812,N_13476,N_13938);
nor U14813 (N_14813,N_13791,N_13086);
and U14814 (N_14814,N_13231,N_13899);
xor U14815 (N_14815,N_13306,N_13378);
and U14816 (N_14816,N_13939,N_13890);
and U14817 (N_14817,N_13367,N_13343);
xnor U14818 (N_14818,N_13844,N_13395);
or U14819 (N_14819,N_13450,N_13848);
nand U14820 (N_14820,N_13449,N_13855);
xnor U14821 (N_14821,N_13539,N_13878);
and U14822 (N_14822,N_13273,N_13543);
xnor U14823 (N_14823,N_13997,N_13880);
nand U14824 (N_14824,N_13899,N_13923);
xnor U14825 (N_14825,N_13061,N_13490);
or U14826 (N_14826,N_13759,N_13497);
nor U14827 (N_14827,N_13740,N_13180);
xnor U14828 (N_14828,N_13937,N_13856);
nand U14829 (N_14829,N_13466,N_13717);
or U14830 (N_14830,N_13868,N_13569);
or U14831 (N_14831,N_13941,N_13306);
nand U14832 (N_14832,N_13257,N_13653);
and U14833 (N_14833,N_13977,N_13001);
or U14834 (N_14834,N_13659,N_13167);
nand U14835 (N_14835,N_13673,N_13461);
or U14836 (N_14836,N_13280,N_13219);
xnor U14837 (N_14837,N_13526,N_13651);
nand U14838 (N_14838,N_13876,N_13576);
xor U14839 (N_14839,N_13087,N_13665);
xor U14840 (N_14840,N_13492,N_13689);
and U14841 (N_14841,N_13548,N_13962);
or U14842 (N_14842,N_13629,N_13361);
xnor U14843 (N_14843,N_13522,N_13880);
and U14844 (N_14844,N_13608,N_13764);
nor U14845 (N_14845,N_13506,N_13745);
or U14846 (N_14846,N_13492,N_13004);
xor U14847 (N_14847,N_13832,N_13589);
nor U14848 (N_14848,N_13444,N_13230);
nand U14849 (N_14849,N_13665,N_13737);
xnor U14850 (N_14850,N_13220,N_13651);
xor U14851 (N_14851,N_13775,N_13755);
nor U14852 (N_14852,N_13942,N_13204);
nand U14853 (N_14853,N_13588,N_13515);
nand U14854 (N_14854,N_13974,N_13142);
or U14855 (N_14855,N_13309,N_13304);
nor U14856 (N_14856,N_13689,N_13342);
xnor U14857 (N_14857,N_13866,N_13053);
nand U14858 (N_14858,N_13596,N_13618);
or U14859 (N_14859,N_13451,N_13431);
or U14860 (N_14860,N_13842,N_13277);
or U14861 (N_14861,N_13754,N_13003);
and U14862 (N_14862,N_13935,N_13575);
nor U14863 (N_14863,N_13983,N_13806);
xnor U14864 (N_14864,N_13282,N_13934);
nand U14865 (N_14865,N_13504,N_13164);
xnor U14866 (N_14866,N_13190,N_13129);
and U14867 (N_14867,N_13566,N_13696);
nor U14868 (N_14868,N_13237,N_13591);
nand U14869 (N_14869,N_13245,N_13703);
xnor U14870 (N_14870,N_13222,N_13495);
nand U14871 (N_14871,N_13673,N_13749);
nand U14872 (N_14872,N_13573,N_13069);
nor U14873 (N_14873,N_13910,N_13716);
or U14874 (N_14874,N_13364,N_13225);
and U14875 (N_14875,N_13890,N_13954);
nand U14876 (N_14876,N_13909,N_13902);
nand U14877 (N_14877,N_13054,N_13017);
nor U14878 (N_14878,N_13097,N_13375);
xnor U14879 (N_14879,N_13854,N_13596);
or U14880 (N_14880,N_13759,N_13915);
or U14881 (N_14881,N_13798,N_13479);
or U14882 (N_14882,N_13048,N_13444);
xnor U14883 (N_14883,N_13941,N_13664);
nor U14884 (N_14884,N_13362,N_13687);
nor U14885 (N_14885,N_13918,N_13892);
or U14886 (N_14886,N_13321,N_13606);
nand U14887 (N_14887,N_13362,N_13026);
or U14888 (N_14888,N_13266,N_13064);
or U14889 (N_14889,N_13238,N_13748);
nand U14890 (N_14890,N_13361,N_13610);
or U14891 (N_14891,N_13791,N_13786);
nor U14892 (N_14892,N_13056,N_13544);
xnor U14893 (N_14893,N_13440,N_13949);
xnor U14894 (N_14894,N_13466,N_13293);
or U14895 (N_14895,N_13299,N_13889);
xnor U14896 (N_14896,N_13216,N_13123);
and U14897 (N_14897,N_13140,N_13830);
nor U14898 (N_14898,N_13375,N_13848);
nand U14899 (N_14899,N_13553,N_13395);
nand U14900 (N_14900,N_13615,N_13446);
xnor U14901 (N_14901,N_13505,N_13387);
or U14902 (N_14902,N_13881,N_13700);
xor U14903 (N_14903,N_13546,N_13369);
or U14904 (N_14904,N_13283,N_13127);
or U14905 (N_14905,N_13568,N_13504);
nor U14906 (N_14906,N_13547,N_13459);
nor U14907 (N_14907,N_13221,N_13607);
and U14908 (N_14908,N_13415,N_13101);
nand U14909 (N_14909,N_13923,N_13806);
or U14910 (N_14910,N_13994,N_13666);
and U14911 (N_14911,N_13849,N_13216);
nand U14912 (N_14912,N_13283,N_13096);
or U14913 (N_14913,N_13882,N_13104);
nand U14914 (N_14914,N_13821,N_13489);
or U14915 (N_14915,N_13504,N_13324);
xnor U14916 (N_14916,N_13887,N_13702);
nor U14917 (N_14917,N_13552,N_13546);
nand U14918 (N_14918,N_13240,N_13942);
or U14919 (N_14919,N_13209,N_13416);
nand U14920 (N_14920,N_13635,N_13424);
or U14921 (N_14921,N_13168,N_13383);
xor U14922 (N_14922,N_13849,N_13859);
nor U14923 (N_14923,N_13264,N_13454);
and U14924 (N_14924,N_13516,N_13833);
or U14925 (N_14925,N_13386,N_13739);
xor U14926 (N_14926,N_13673,N_13370);
and U14927 (N_14927,N_13828,N_13217);
and U14928 (N_14928,N_13672,N_13992);
nor U14929 (N_14929,N_13033,N_13996);
nor U14930 (N_14930,N_13283,N_13959);
or U14931 (N_14931,N_13225,N_13763);
or U14932 (N_14932,N_13063,N_13102);
or U14933 (N_14933,N_13747,N_13047);
xnor U14934 (N_14934,N_13302,N_13375);
or U14935 (N_14935,N_13664,N_13957);
xnor U14936 (N_14936,N_13082,N_13021);
nor U14937 (N_14937,N_13090,N_13354);
xor U14938 (N_14938,N_13635,N_13795);
nand U14939 (N_14939,N_13205,N_13859);
and U14940 (N_14940,N_13140,N_13698);
nor U14941 (N_14941,N_13732,N_13037);
nor U14942 (N_14942,N_13379,N_13400);
or U14943 (N_14943,N_13124,N_13507);
nor U14944 (N_14944,N_13764,N_13080);
and U14945 (N_14945,N_13045,N_13710);
nand U14946 (N_14946,N_13706,N_13736);
or U14947 (N_14947,N_13609,N_13825);
xnor U14948 (N_14948,N_13233,N_13643);
nand U14949 (N_14949,N_13163,N_13156);
nand U14950 (N_14950,N_13059,N_13341);
and U14951 (N_14951,N_13091,N_13238);
and U14952 (N_14952,N_13213,N_13696);
or U14953 (N_14953,N_13259,N_13932);
and U14954 (N_14954,N_13971,N_13326);
xnor U14955 (N_14955,N_13137,N_13750);
and U14956 (N_14956,N_13431,N_13551);
nor U14957 (N_14957,N_13670,N_13532);
and U14958 (N_14958,N_13304,N_13787);
or U14959 (N_14959,N_13027,N_13710);
and U14960 (N_14960,N_13938,N_13940);
or U14961 (N_14961,N_13271,N_13357);
xor U14962 (N_14962,N_13774,N_13368);
xnor U14963 (N_14963,N_13302,N_13579);
or U14964 (N_14964,N_13782,N_13516);
nand U14965 (N_14965,N_13071,N_13841);
and U14966 (N_14966,N_13752,N_13693);
nor U14967 (N_14967,N_13334,N_13855);
nor U14968 (N_14968,N_13760,N_13004);
xor U14969 (N_14969,N_13574,N_13113);
nor U14970 (N_14970,N_13059,N_13008);
and U14971 (N_14971,N_13732,N_13454);
and U14972 (N_14972,N_13557,N_13732);
nor U14973 (N_14973,N_13942,N_13563);
xor U14974 (N_14974,N_13625,N_13446);
or U14975 (N_14975,N_13616,N_13037);
and U14976 (N_14976,N_13083,N_13067);
and U14977 (N_14977,N_13164,N_13043);
or U14978 (N_14978,N_13665,N_13116);
nor U14979 (N_14979,N_13429,N_13243);
and U14980 (N_14980,N_13533,N_13594);
or U14981 (N_14981,N_13064,N_13310);
and U14982 (N_14982,N_13161,N_13977);
nor U14983 (N_14983,N_13573,N_13497);
nor U14984 (N_14984,N_13407,N_13471);
and U14985 (N_14985,N_13391,N_13042);
nand U14986 (N_14986,N_13892,N_13018);
xnor U14987 (N_14987,N_13410,N_13358);
nand U14988 (N_14988,N_13032,N_13901);
nor U14989 (N_14989,N_13714,N_13308);
nor U14990 (N_14990,N_13867,N_13499);
nor U14991 (N_14991,N_13031,N_13225);
xor U14992 (N_14992,N_13715,N_13859);
and U14993 (N_14993,N_13524,N_13171);
nand U14994 (N_14994,N_13939,N_13791);
nor U14995 (N_14995,N_13131,N_13531);
or U14996 (N_14996,N_13800,N_13402);
xnor U14997 (N_14997,N_13812,N_13019);
or U14998 (N_14998,N_13751,N_13927);
and U14999 (N_14999,N_13954,N_13898);
nor U15000 (N_15000,N_14293,N_14516);
nor U15001 (N_15001,N_14152,N_14762);
and U15002 (N_15002,N_14462,N_14554);
nor U15003 (N_15003,N_14242,N_14454);
and U15004 (N_15004,N_14286,N_14647);
and U15005 (N_15005,N_14822,N_14206);
or U15006 (N_15006,N_14795,N_14075);
nor U15007 (N_15007,N_14529,N_14494);
nand U15008 (N_15008,N_14411,N_14291);
xor U15009 (N_15009,N_14926,N_14547);
and U15010 (N_15010,N_14840,N_14079);
nor U15011 (N_15011,N_14819,N_14791);
nand U15012 (N_15012,N_14948,N_14330);
nor U15013 (N_15013,N_14639,N_14222);
or U15014 (N_15014,N_14219,N_14004);
nand U15015 (N_15015,N_14017,N_14631);
and U15016 (N_15016,N_14747,N_14183);
nand U15017 (N_15017,N_14685,N_14969);
or U15018 (N_15018,N_14146,N_14843);
and U15019 (N_15019,N_14193,N_14739);
nand U15020 (N_15020,N_14419,N_14629);
xor U15021 (N_15021,N_14560,N_14883);
nand U15022 (N_15022,N_14596,N_14216);
nand U15023 (N_15023,N_14913,N_14750);
nand U15024 (N_15024,N_14717,N_14113);
and U15025 (N_15025,N_14887,N_14586);
or U15026 (N_15026,N_14395,N_14888);
or U15027 (N_15027,N_14059,N_14711);
xnor U15028 (N_15028,N_14583,N_14775);
nand U15029 (N_15029,N_14846,N_14692);
and U15030 (N_15030,N_14285,N_14910);
and U15031 (N_15031,N_14294,N_14947);
and U15032 (N_15032,N_14087,N_14379);
and U15033 (N_15033,N_14437,N_14319);
nor U15034 (N_15034,N_14140,N_14618);
nand U15035 (N_15035,N_14033,N_14155);
and U15036 (N_15036,N_14986,N_14442);
xor U15037 (N_15037,N_14545,N_14557);
nor U15038 (N_15038,N_14011,N_14720);
or U15039 (N_15039,N_14591,N_14849);
xnor U15040 (N_15040,N_14376,N_14231);
and U15041 (N_15041,N_14387,N_14686);
xor U15042 (N_15042,N_14851,N_14946);
nand U15043 (N_15043,N_14299,N_14177);
nor U15044 (N_15044,N_14374,N_14654);
or U15045 (N_15045,N_14148,N_14467);
or U15046 (N_15046,N_14570,N_14649);
and U15047 (N_15047,N_14452,N_14905);
xor U15048 (N_15048,N_14798,N_14069);
nand U15049 (N_15049,N_14042,N_14809);
nand U15050 (N_15050,N_14154,N_14701);
and U15051 (N_15051,N_14725,N_14919);
nor U15052 (N_15052,N_14641,N_14471);
or U15053 (N_15053,N_14517,N_14036);
nor U15054 (N_15054,N_14492,N_14681);
or U15055 (N_15055,N_14901,N_14027);
or U15056 (N_15056,N_14116,N_14716);
nor U15057 (N_15057,N_14198,N_14574);
and U15058 (N_15058,N_14035,N_14498);
nor U15059 (N_15059,N_14766,N_14745);
nor U15060 (N_15060,N_14223,N_14371);
nor U15061 (N_15061,N_14857,N_14131);
xor U15062 (N_15062,N_14007,N_14125);
or U15063 (N_15063,N_14663,N_14207);
nor U15064 (N_15064,N_14126,N_14705);
and U15065 (N_15065,N_14553,N_14549);
or U15066 (N_15066,N_14904,N_14331);
nand U15067 (N_15067,N_14671,N_14267);
and U15068 (N_15068,N_14665,N_14963);
xor U15069 (N_15069,N_14160,N_14188);
xor U15070 (N_15070,N_14891,N_14759);
nor U15071 (N_15071,N_14501,N_14070);
nor U15072 (N_15072,N_14251,N_14730);
and U15073 (N_15073,N_14388,N_14072);
nand U15074 (N_15074,N_14412,N_14834);
and U15075 (N_15075,N_14302,N_14831);
nor U15076 (N_15076,N_14788,N_14200);
and U15077 (N_15077,N_14226,N_14953);
nor U15078 (N_15078,N_14082,N_14472);
and U15079 (N_15079,N_14392,N_14264);
xor U15080 (N_15080,N_14550,N_14425);
xnor U15081 (N_15081,N_14078,N_14559);
or U15082 (N_15082,N_14732,N_14579);
or U15083 (N_15083,N_14839,N_14039);
or U15084 (N_15084,N_14777,N_14165);
nor U15085 (N_15085,N_14841,N_14714);
xor U15086 (N_15086,N_14283,N_14312);
nand U15087 (N_15087,N_14358,N_14627);
xor U15088 (N_15088,N_14185,N_14749);
or U15089 (N_15089,N_14748,N_14523);
nand U15090 (N_15090,N_14785,N_14053);
nor U15091 (N_15091,N_14490,N_14751);
nand U15092 (N_15092,N_14172,N_14088);
nor U15093 (N_15093,N_14334,N_14943);
and U15094 (N_15094,N_14847,N_14562);
xor U15095 (N_15095,N_14384,N_14908);
xnor U15096 (N_15096,N_14459,N_14248);
nor U15097 (N_15097,N_14932,N_14451);
nor U15098 (N_15098,N_14608,N_14658);
or U15099 (N_15099,N_14994,N_14449);
and U15100 (N_15100,N_14230,N_14531);
nand U15101 (N_15101,N_14651,N_14962);
nand U15102 (N_15102,N_14724,N_14060);
or U15103 (N_15103,N_14927,N_14588);
or U15104 (N_15104,N_14166,N_14244);
nand U15105 (N_15105,N_14202,N_14611);
nand U15106 (N_15106,N_14619,N_14266);
and U15107 (N_15107,N_14170,N_14130);
xor U15108 (N_15108,N_14333,N_14793);
or U15109 (N_15109,N_14678,N_14563);
nor U15110 (N_15110,N_14282,N_14105);
nand U15111 (N_15111,N_14068,N_14213);
nand U15112 (N_15112,N_14998,N_14773);
and U15113 (N_15113,N_14741,N_14316);
nor U15114 (N_15114,N_14979,N_14199);
and U15115 (N_15115,N_14045,N_14761);
or U15116 (N_15116,N_14044,N_14561);
nand U15117 (N_15117,N_14061,N_14102);
and U15118 (N_15118,N_14900,N_14378);
or U15119 (N_15119,N_14505,N_14295);
xor U15120 (N_15120,N_14178,N_14504);
or U15121 (N_15121,N_14642,N_14881);
nor U15122 (N_15122,N_14852,N_14546);
nor U15123 (N_15123,N_14210,N_14957);
and U15124 (N_15124,N_14694,N_14578);
xnor U15125 (N_15125,N_14783,N_14342);
nand U15126 (N_15126,N_14931,N_14071);
and U15127 (N_15127,N_14814,N_14643);
nor U15128 (N_15128,N_14424,N_14744);
nand U15129 (N_15129,N_14280,N_14365);
and U15130 (N_15130,N_14799,N_14848);
or U15131 (N_15131,N_14622,N_14488);
nand U15132 (N_15132,N_14593,N_14487);
and U15133 (N_15133,N_14753,N_14014);
xor U15134 (N_15134,N_14037,N_14010);
nor U15135 (N_15135,N_14434,N_14854);
nor U15136 (N_15136,N_14975,N_14604);
nor U15137 (N_15137,N_14229,N_14301);
nor U15138 (N_15138,N_14176,N_14917);
nor U15139 (N_15139,N_14179,N_14268);
nor U15140 (N_15140,N_14461,N_14064);
nor U15141 (N_15141,N_14278,N_14988);
nand U15142 (N_15142,N_14617,N_14247);
xor U15143 (N_15143,N_14405,N_14937);
or U15144 (N_15144,N_14009,N_14048);
or U15145 (N_15145,N_14811,N_14101);
nand U15146 (N_15146,N_14606,N_14237);
or U15147 (N_15147,N_14086,N_14275);
nor U15148 (N_15148,N_14427,N_14001);
or U15149 (N_15149,N_14352,N_14112);
nor U15150 (N_15150,N_14477,N_14043);
nor U15151 (N_15151,N_14544,N_14907);
and U15152 (N_15152,N_14916,N_14510);
nor U15153 (N_15153,N_14702,N_14002);
nand U15154 (N_15154,N_14174,N_14952);
or U15155 (N_15155,N_14095,N_14245);
xnor U15156 (N_15156,N_14710,N_14008);
or U15157 (N_15157,N_14463,N_14816);
nand U15158 (N_15158,N_14934,N_14699);
and U15159 (N_15159,N_14191,N_14965);
nand U15160 (N_15160,N_14215,N_14922);
nand U15161 (N_15161,N_14738,N_14339);
nor U15162 (N_15162,N_14406,N_14889);
and U15163 (N_15163,N_14933,N_14401);
and U15164 (N_15164,N_14864,N_14423);
nor U15165 (N_15165,N_14465,N_14915);
xnor U15166 (N_15166,N_14296,N_14813);
or U15167 (N_15167,N_14448,N_14089);
xnor U15168 (N_15168,N_14515,N_14566);
xnor U15169 (N_15169,N_14225,N_14599);
nand U15170 (N_15170,N_14478,N_14391);
and U15171 (N_15171,N_14169,N_14197);
xnor U15172 (N_15172,N_14511,N_14802);
xor U15173 (N_15173,N_14496,N_14259);
and U15174 (N_15174,N_14743,N_14398);
nor U15175 (N_15175,N_14346,N_14019);
and U15176 (N_15176,N_14149,N_14127);
xnor U15177 (N_15177,N_14196,N_14500);
xor U15178 (N_15178,N_14984,N_14866);
nand U15179 (N_15179,N_14956,N_14661);
or U15180 (N_15180,N_14964,N_14855);
nand U15181 (N_15181,N_14117,N_14790);
xor U15182 (N_15182,N_14313,N_14603);
and U15183 (N_15183,N_14484,N_14537);
xnor U15184 (N_15184,N_14114,N_14343);
xnor U15185 (N_15185,N_14800,N_14836);
xnor U15186 (N_15186,N_14145,N_14897);
or U15187 (N_15187,N_14370,N_14135);
or U15188 (N_15188,N_14568,N_14949);
and U15189 (N_15189,N_14491,N_14094);
nor U15190 (N_15190,N_14779,N_14447);
and U15191 (N_15191,N_14960,N_14616);
nand U15192 (N_15192,N_14122,N_14914);
and U15193 (N_15193,N_14390,N_14065);
or U15194 (N_15194,N_14119,N_14729);
xor U15195 (N_15195,N_14679,N_14203);
and U15196 (N_15196,N_14826,N_14414);
xnor U15197 (N_15197,N_14756,N_14921);
nor U15198 (N_15198,N_14438,N_14375);
and U15199 (N_15199,N_14935,N_14718);
and U15200 (N_15200,N_14522,N_14805);
and U15201 (N_15201,N_14763,N_14228);
nor U15202 (N_15202,N_14520,N_14476);
and U15203 (N_15203,N_14277,N_14723);
xnor U15204 (N_15204,N_14046,N_14107);
and U15205 (N_15205,N_14415,N_14542);
nor U15206 (N_15206,N_14524,N_14493);
nand U15207 (N_15207,N_14156,N_14354);
xor U15208 (N_15208,N_14909,N_14697);
xor U15209 (N_15209,N_14689,N_14509);
and U15210 (N_15210,N_14249,N_14551);
xor U15211 (N_15211,N_14121,N_14640);
nor U15212 (N_15212,N_14458,N_14066);
and U15213 (N_15213,N_14784,N_14351);
xnor U15214 (N_15214,N_14539,N_14162);
or U15215 (N_15215,N_14924,N_14828);
nor U15216 (N_15216,N_14413,N_14092);
xnor U15217 (N_15217,N_14818,N_14115);
or U15218 (N_15218,N_14556,N_14304);
nor U15219 (N_15219,N_14499,N_14440);
xnor U15220 (N_15220,N_14298,N_14151);
nor U15221 (N_15221,N_14409,N_14276);
and U15222 (N_15222,N_14896,N_14049);
nor U15223 (N_15223,N_14138,N_14625);
nor U15224 (N_15224,N_14817,N_14845);
nand U15225 (N_15225,N_14677,N_14977);
and U15226 (N_15226,N_14990,N_14605);
nor U15227 (N_15227,N_14360,N_14860);
xnor U15228 (N_15228,N_14533,N_14704);
nand U15229 (N_15229,N_14912,N_14644);
or U15230 (N_15230,N_14770,N_14450);
xor U15231 (N_15231,N_14621,N_14534);
xor U15232 (N_15232,N_14980,N_14576);
nor U15233 (N_15233,N_14161,N_14722);
and U15234 (N_15234,N_14205,N_14595);
nand U15235 (N_15235,N_14584,N_14133);
xnor U15236 (N_15236,N_14587,N_14754);
or U15237 (N_15237,N_14815,N_14755);
or U15238 (N_15238,N_14309,N_14292);
nand U15239 (N_15239,N_14103,N_14399);
or U15240 (N_15240,N_14243,N_14760);
and U15241 (N_15241,N_14324,N_14380);
xnor U15242 (N_15242,N_14961,N_14232);
and U15243 (N_15243,N_14804,N_14526);
xnor U15244 (N_15244,N_14950,N_14527);
nand U15245 (N_15245,N_14981,N_14862);
and U15246 (N_15246,N_14633,N_14382);
and U15247 (N_15247,N_14297,N_14322);
xnor U15248 (N_15248,N_14323,N_14073);
nor U15249 (N_15249,N_14973,N_14485);
nor U15250 (N_15250,N_14077,N_14925);
xor U15251 (N_15251,N_14429,N_14320);
and U15252 (N_15252,N_14090,N_14967);
nor U15253 (N_15253,N_14212,N_14218);
or U15254 (N_15254,N_14991,N_14564);
xnor U15255 (N_15255,N_14664,N_14827);
or U15256 (N_15256,N_14894,N_14270);
and U15257 (N_15257,N_14794,N_14483);
or U15258 (N_15258,N_14100,N_14480);
nor U15259 (N_15259,N_14000,N_14305);
nand U15260 (N_15260,N_14335,N_14361);
nand U15261 (N_15261,N_14288,N_14274);
or U15262 (N_15262,N_14428,N_14796);
nor U15263 (N_15263,N_14396,N_14648);
nor U15264 (N_15264,N_14159,N_14792);
and U15265 (N_15265,N_14475,N_14938);
and U15266 (N_15266,N_14650,N_14863);
or U15267 (N_15267,N_14700,N_14022);
or U15268 (N_15268,N_14110,N_14431);
or U15269 (N_15269,N_14150,N_14164);
or U15270 (N_15270,N_14441,N_14466);
nand U15271 (N_15271,N_14672,N_14257);
or U15272 (N_15272,N_14613,N_14808);
or U15273 (N_15273,N_14347,N_14646);
and U15274 (N_15274,N_14377,N_14186);
nor U15275 (N_15275,N_14328,N_14246);
nor U15276 (N_15276,N_14781,N_14120);
nor U15277 (N_15277,N_14404,N_14735);
nand U15278 (N_15278,N_14632,N_14688);
nand U15279 (N_15279,N_14989,N_14337);
or U15280 (N_15280,N_14364,N_14942);
xor U15281 (N_15281,N_14940,N_14873);
or U15282 (N_15282,N_14582,N_14870);
xor U15283 (N_15283,N_14250,N_14820);
nand U15284 (N_15284,N_14996,N_14951);
nand U15285 (N_15285,N_14778,N_14659);
xnor U15286 (N_15286,N_14992,N_14410);
or U15287 (N_15287,N_14163,N_14684);
and U15288 (N_15288,N_14945,N_14597);
and U15289 (N_15289,N_14740,N_14728);
and U15290 (N_15290,N_14056,N_14106);
nor U15291 (N_15291,N_14696,N_14012);
nor U15292 (N_15292,N_14669,N_14468);
nand U15293 (N_15293,N_14372,N_14108);
and U15294 (N_15294,N_14709,N_14030);
nand U15295 (N_15295,N_14580,N_14332);
nand U15296 (N_15296,N_14006,N_14906);
nor U15297 (N_15297,N_14139,N_14607);
and U15298 (N_15298,N_14939,N_14682);
nor U15299 (N_15299,N_14217,N_14124);
or U15300 (N_15300,N_14220,N_14464);
xor U15301 (N_15301,N_14143,N_14407);
nand U15302 (N_15302,N_14832,N_14084);
xor U15303 (N_15303,N_14667,N_14572);
or U15304 (N_15304,N_14201,N_14063);
nand U15305 (N_15305,N_14005,N_14569);
nand U15306 (N_15306,N_14214,N_14144);
or U15307 (N_15307,N_14512,N_14235);
nor U15308 (N_15308,N_14444,N_14928);
xor U15309 (N_15309,N_14470,N_14902);
nand U15310 (N_15310,N_14047,N_14879);
nand U15311 (N_15311,N_14742,N_14706);
nand U15312 (N_15312,N_14898,N_14041);
nor U15313 (N_15313,N_14211,N_14055);
or U15314 (N_15314,N_14944,N_14054);
or U15315 (N_15315,N_14460,N_14136);
nor U15316 (N_15316,N_14999,N_14703);
xnor U15317 (N_15317,N_14978,N_14971);
xnor U15318 (N_15318,N_14393,N_14726);
nand U15319 (N_15319,N_14349,N_14708);
xnor U15320 (N_15320,N_14880,N_14737);
nand U15321 (N_15321,N_14344,N_14624);
or U15322 (N_15322,N_14481,N_14474);
nand U15323 (N_15323,N_14363,N_14421);
or U15324 (N_15324,N_14394,N_14872);
nor U15325 (N_15325,N_14532,N_14966);
or U15326 (N_15326,N_14445,N_14920);
or U15327 (N_15327,N_14776,N_14194);
or U15328 (N_15328,N_14565,N_14208);
nor U15329 (N_15329,N_14356,N_14204);
and U15330 (N_15330,N_14609,N_14080);
and U15331 (N_15331,N_14638,N_14034);
and U15332 (N_15332,N_14098,N_14308);
and U15333 (N_15333,N_14752,N_14540);
or U15334 (N_15334,N_14495,N_14029);
nor U15335 (N_15335,N_14837,N_14683);
or U15336 (N_15336,N_14013,N_14600);
nor U15337 (N_15337,N_14408,N_14081);
nor U15338 (N_15338,N_14987,N_14221);
nor U15339 (N_15339,N_14167,N_14719);
or U15340 (N_15340,N_14571,N_14626);
or U15341 (N_15341,N_14918,N_14757);
or U15342 (N_15342,N_14536,N_14543);
nand U15343 (N_15343,N_14353,N_14040);
or U15344 (N_15344,N_14224,N_14861);
nand U15345 (N_15345,N_14653,N_14015);
or U15346 (N_15346,N_14974,N_14782);
xnor U15347 (N_15347,N_14713,N_14687);
nor U15348 (N_15348,N_14209,N_14253);
nand U15349 (N_15349,N_14340,N_14830);
nor U15350 (N_15350,N_14585,N_14118);
and U15351 (N_15351,N_14676,N_14482);
nor U15352 (N_15352,N_14525,N_14637);
nor U15353 (N_15353,N_14182,N_14284);
or U15354 (N_15354,N_14123,N_14195);
xor U15355 (N_15355,N_14051,N_14656);
or U15356 (N_15356,N_14435,N_14137);
nor U15357 (N_15357,N_14290,N_14801);
nor U15358 (N_15358,N_14469,N_14109);
xnor U15359 (N_15359,N_14911,N_14016);
and U15360 (N_15360,N_14263,N_14385);
nand U15361 (N_15361,N_14670,N_14780);
and U15362 (N_15362,N_14997,N_14258);
xnor U15363 (N_15363,N_14976,N_14882);
nor U15364 (N_15364,N_14521,N_14577);
xnor U15365 (N_15365,N_14479,N_14317);
and U15366 (N_15366,N_14812,N_14180);
nor U15367 (N_15367,N_14329,N_14628);
and U15368 (N_15368,N_14623,N_14844);
or U15369 (N_15369,N_14003,N_14503);
and U15370 (N_15370,N_14765,N_14955);
xnor U15371 (N_15371,N_14386,N_14307);
and U15372 (N_15372,N_14303,N_14367);
or U15373 (N_15373,N_14548,N_14573);
nor U15374 (N_15374,N_14240,N_14610);
xor U15375 (N_15375,N_14734,N_14239);
or U15376 (N_15376,N_14985,N_14675);
nor U15377 (N_15377,N_14026,N_14567);
and U15378 (N_15378,N_14050,N_14514);
or U15379 (N_15379,N_14803,N_14318);
or U15380 (N_15380,N_14829,N_14530);
and U15381 (N_15381,N_14129,N_14528);
or U15382 (N_15382,N_14052,N_14764);
xor U15383 (N_15383,N_14327,N_14128);
and U15384 (N_15384,N_14097,N_14995);
nand U15385 (N_15385,N_14903,N_14457);
and U15386 (N_15386,N_14300,N_14456);
and U15387 (N_15387,N_14721,N_14733);
and U15388 (N_15388,N_14368,N_14581);
nand U15389 (N_15389,N_14345,N_14189);
nor U15390 (N_15390,N_14262,N_14173);
and U15391 (N_15391,N_14134,N_14400);
or U15392 (N_15392,N_14810,N_14338);
xor U15393 (N_15393,N_14871,N_14383);
nor U15394 (N_15394,N_14104,N_14083);
and U15395 (N_15395,N_14707,N_14321);
and U15396 (N_15396,N_14359,N_14031);
nor U15397 (N_15397,N_14892,N_14858);
or U15398 (N_15398,N_14555,N_14418);
or U15399 (N_15399,N_14954,N_14727);
nand U15400 (N_15400,N_14369,N_14612);
and U15401 (N_15401,N_14575,N_14184);
xor U15402 (N_15402,N_14715,N_14168);
and U15403 (N_15403,N_14630,N_14673);
xor U15404 (N_15404,N_14772,N_14662);
xnor U15405 (N_15405,N_14899,N_14306);
nand U15406 (N_15406,N_14153,N_14513);
and U15407 (N_15407,N_14142,N_14789);
nor U15408 (N_15408,N_14859,N_14256);
nand U15409 (N_15409,N_14381,N_14970);
nand U15410 (N_15410,N_14806,N_14497);
nand U15411 (N_15411,N_14227,N_14698);
or U15412 (N_15412,N_14020,N_14397);
xor U15413 (N_15413,N_14238,N_14175);
nor U15414 (N_15414,N_14786,N_14355);
nand U15415 (N_15415,N_14091,N_14265);
nand U15416 (N_15416,N_14348,N_14652);
xor U15417 (N_15417,N_14821,N_14455);
nor U15418 (N_15418,N_14538,N_14787);
xnor U15419 (N_15419,N_14062,N_14635);
nor U15420 (N_15420,N_14807,N_14972);
nor U15421 (N_15421,N_14453,N_14272);
and U15422 (N_15422,N_14058,N_14645);
or U15423 (N_15423,N_14096,N_14132);
and U15424 (N_15424,N_14326,N_14982);
nor U15425 (N_15425,N_14634,N_14325);
or U15426 (N_15426,N_14430,N_14590);
and U15427 (N_15427,N_14422,N_14993);
nor U15428 (N_15428,N_14067,N_14691);
and U15429 (N_15429,N_14518,N_14885);
nor U15430 (N_15430,N_14731,N_14594);
nand U15431 (N_15431,N_14833,N_14024);
nand U15432 (N_15432,N_14158,N_14157);
or U15433 (N_15433,N_14884,N_14099);
and U15434 (N_15434,N_14025,N_14038);
or U15435 (N_15435,N_14983,N_14366);
nand U15436 (N_15436,N_14655,N_14416);
nor U15437 (N_15437,N_14959,N_14190);
xnor U15438 (N_15438,N_14602,N_14271);
and U15439 (N_15439,N_14028,N_14236);
nor U15440 (N_15440,N_14535,N_14598);
nor U15441 (N_15441,N_14233,N_14433);
nand U15442 (N_15442,N_14774,N_14085);
nor U15443 (N_15443,N_14680,N_14824);
or U15444 (N_15444,N_14620,N_14552);
nand U15445 (N_15445,N_14666,N_14660);
and U15446 (N_15446,N_14032,N_14234);
nor U15447 (N_15447,N_14187,N_14838);
and U15448 (N_15448,N_14171,N_14695);
or U15449 (N_15449,N_14893,N_14402);
or U15450 (N_15450,N_14023,N_14289);
and U15451 (N_15451,N_14519,N_14758);
and U15452 (N_15452,N_14436,N_14111);
xor U15453 (N_15453,N_14541,N_14823);
xnor U15454 (N_15454,N_14769,N_14426);
and U15455 (N_15455,N_14506,N_14875);
and U15456 (N_15456,N_14507,N_14315);
nand U15457 (N_15457,N_14417,N_14601);
nor U15458 (N_15458,N_14941,N_14432);
or U15459 (N_15459,N_14141,N_14850);
and U15460 (N_15460,N_14657,N_14252);
or U15461 (N_15461,N_14825,N_14181);
nor U15462 (N_15462,N_14868,N_14895);
or U15463 (N_15463,N_14968,N_14403);
nand U15464 (N_15464,N_14261,N_14260);
and U15465 (N_15465,N_14362,N_14508);
nand U15466 (N_15466,N_14877,N_14615);
nor U15467 (N_15467,N_14269,N_14254);
and U15468 (N_15468,N_14093,N_14736);
or U15469 (N_15469,N_14929,N_14958);
or U15470 (N_15470,N_14771,N_14865);
or U15471 (N_15471,N_14446,N_14768);
nor U15472 (N_15472,N_14473,N_14668);
nor U15473 (N_15473,N_14018,N_14878);
nand U15474 (N_15474,N_14021,N_14592);
nor U15475 (N_15475,N_14502,N_14890);
and U15476 (N_15476,N_14074,N_14057);
xnor U15477 (N_15477,N_14923,N_14336);
nand U15478 (N_15478,N_14357,N_14853);
or U15479 (N_15479,N_14930,N_14876);
and U15480 (N_15480,N_14341,N_14746);
nand U15481 (N_15481,N_14373,N_14255);
nand U15482 (N_15482,N_14486,N_14439);
xnor U15483 (N_15483,N_14936,N_14674);
and U15484 (N_15484,N_14389,N_14241);
nand U15485 (N_15485,N_14712,N_14589);
nor U15486 (N_15486,N_14281,N_14310);
nand U15487 (N_15487,N_14867,N_14874);
nand U15488 (N_15488,N_14311,N_14076);
nand U15489 (N_15489,N_14835,N_14636);
and U15490 (N_15490,N_14690,N_14279);
or U15491 (N_15491,N_14614,N_14273);
xor U15492 (N_15492,N_14558,N_14869);
and U15493 (N_15493,N_14489,N_14350);
nand U15494 (N_15494,N_14767,N_14856);
nand U15495 (N_15495,N_14886,N_14287);
nor U15496 (N_15496,N_14147,N_14420);
nor U15497 (N_15497,N_14797,N_14693);
nand U15498 (N_15498,N_14443,N_14314);
nand U15499 (N_15499,N_14842,N_14192);
and U15500 (N_15500,N_14322,N_14439);
xor U15501 (N_15501,N_14942,N_14823);
nand U15502 (N_15502,N_14397,N_14737);
and U15503 (N_15503,N_14278,N_14172);
xor U15504 (N_15504,N_14129,N_14878);
nand U15505 (N_15505,N_14017,N_14572);
nand U15506 (N_15506,N_14805,N_14229);
xnor U15507 (N_15507,N_14143,N_14264);
or U15508 (N_15508,N_14125,N_14617);
nand U15509 (N_15509,N_14198,N_14832);
nor U15510 (N_15510,N_14315,N_14870);
nor U15511 (N_15511,N_14753,N_14500);
xnor U15512 (N_15512,N_14561,N_14249);
nand U15513 (N_15513,N_14259,N_14805);
nand U15514 (N_15514,N_14599,N_14907);
nand U15515 (N_15515,N_14658,N_14897);
xnor U15516 (N_15516,N_14598,N_14995);
or U15517 (N_15517,N_14468,N_14690);
xor U15518 (N_15518,N_14273,N_14666);
or U15519 (N_15519,N_14032,N_14518);
and U15520 (N_15520,N_14367,N_14907);
nand U15521 (N_15521,N_14133,N_14235);
nand U15522 (N_15522,N_14553,N_14838);
xor U15523 (N_15523,N_14668,N_14765);
or U15524 (N_15524,N_14192,N_14400);
and U15525 (N_15525,N_14194,N_14155);
or U15526 (N_15526,N_14843,N_14856);
or U15527 (N_15527,N_14380,N_14165);
nor U15528 (N_15528,N_14841,N_14528);
or U15529 (N_15529,N_14099,N_14893);
and U15530 (N_15530,N_14591,N_14915);
nand U15531 (N_15531,N_14673,N_14136);
and U15532 (N_15532,N_14726,N_14579);
nor U15533 (N_15533,N_14815,N_14201);
or U15534 (N_15534,N_14659,N_14629);
nand U15535 (N_15535,N_14277,N_14695);
and U15536 (N_15536,N_14184,N_14841);
and U15537 (N_15537,N_14345,N_14236);
or U15538 (N_15538,N_14557,N_14964);
or U15539 (N_15539,N_14011,N_14862);
or U15540 (N_15540,N_14063,N_14738);
nor U15541 (N_15541,N_14684,N_14483);
nand U15542 (N_15542,N_14730,N_14238);
xnor U15543 (N_15543,N_14571,N_14685);
and U15544 (N_15544,N_14456,N_14563);
nor U15545 (N_15545,N_14404,N_14057);
nor U15546 (N_15546,N_14111,N_14810);
and U15547 (N_15547,N_14718,N_14953);
and U15548 (N_15548,N_14839,N_14913);
and U15549 (N_15549,N_14583,N_14952);
nand U15550 (N_15550,N_14470,N_14399);
nand U15551 (N_15551,N_14767,N_14550);
xor U15552 (N_15552,N_14969,N_14923);
and U15553 (N_15553,N_14544,N_14817);
nor U15554 (N_15554,N_14049,N_14736);
nor U15555 (N_15555,N_14015,N_14611);
or U15556 (N_15556,N_14102,N_14059);
or U15557 (N_15557,N_14926,N_14750);
or U15558 (N_15558,N_14652,N_14270);
nor U15559 (N_15559,N_14026,N_14404);
nor U15560 (N_15560,N_14841,N_14974);
nand U15561 (N_15561,N_14176,N_14784);
and U15562 (N_15562,N_14800,N_14040);
or U15563 (N_15563,N_14886,N_14254);
xor U15564 (N_15564,N_14469,N_14283);
and U15565 (N_15565,N_14766,N_14778);
or U15566 (N_15566,N_14970,N_14867);
xor U15567 (N_15567,N_14720,N_14924);
or U15568 (N_15568,N_14637,N_14330);
nand U15569 (N_15569,N_14893,N_14781);
and U15570 (N_15570,N_14632,N_14842);
and U15571 (N_15571,N_14747,N_14743);
nor U15572 (N_15572,N_14956,N_14121);
and U15573 (N_15573,N_14971,N_14445);
xnor U15574 (N_15574,N_14837,N_14595);
nor U15575 (N_15575,N_14091,N_14555);
nor U15576 (N_15576,N_14209,N_14191);
xnor U15577 (N_15577,N_14414,N_14756);
xnor U15578 (N_15578,N_14897,N_14015);
nor U15579 (N_15579,N_14647,N_14370);
or U15580 (N_15580,N_14286,N_14237);
nand U15581 (N_15581,N_14704,N_14316);
nand U15582 (N_15582,N_14065,N_14003);
or U15583 (N_15583,N_14677,N_14967);
xor U15584 (N_15584,N_14458,N_14625);
nand U15585 (N_15585,N_14194,N_14620);
or U15586 (N_15586,N_14685,N_14180);
or U15587 (N_15587,N_14316,N_14329);
xnor U15588 (N_15588,N_14318,N_14888);
or U15589 (N_15589,N_14177,N_14484);
or U15590 (N_15590,N_14922,N_14456);
nand U15591 (N_15591,N_14783,N_14354);
and U15592 (N_15592,N_14716,N_14146);
and U15593 (N_15593,N_14901,N_14561);
nor U15594 (N_15594,N_14723,N_14072);
or U15595 (N_15595,N_14763,N_14755);
xnor U15596 (N_15596,N_14558,N_14086);
xnor U15597 (N_15597,N_14585,N_14062);
nor U15598 (N_15598,N_14147,N_14027);
or U15599 (N_15599,N_14354,N_14253);
and U15600 (N_15600,N_14225,N_14573);
nand U15601 (N_15601,N_14844,N_14001);
nor U15602 (N_15602,N_14603,N_14258);
or U15603 (N_15603,N_14950,N_14149);
and U15604 (N_15604,N_14951,N_14035);
and U15605 (N_15605,N_14543,N_14496);
nor U15606 (N_15606,N_14446,N_14744);
nor U15607 (N_15607,N_14209,N_14669);
nor U15608 (N_15608,N_14693,N_14820);
or U15609 (N_15609,N_14781,N_14440);
or U15610 (N_15610,N_14596,N_14030);
and U15611 (N_15611,N_14885,N_14145);
nor U15612 (N_15612,N_14855,N_14021);
nand U15613 (N_15613,N_14554,N_14147);
or U15614 (N_15614,N_14924,N_14735);
xor U15615 (N_15615,N_14202,N_14503);
xnor U15616 (N_15616,N_14589,N_14745);
or U15617 (N_15617,N_14836,N_14316);
xor U15618 (N_15618,N_14630,N_14788);
nand U15619 (N_15619,N_14932,N_14133);
nor U15620 (N_15620,N_14001,N_14993);
or U15621 (N_15621,N_14331,N_14717);
nor U15622 (N_15622,N_14454,N_14336);
xnor U15623 (N_15623,N_14528,N_14412);
nand U15624 (N_15624,N_14447,N_14053);
nor U15625 (N_15625,N_14742,N_14416);
nand U15626 (N_15626,N_14225,N_14795);
and U15627 (N_15627,N_14218,N_14364);
nor U15628 (N_15628,N_14380,N_14289);
nor U15629 (N_15629,N_14714,N_14152);
xnor U15630 (N_15630,N_14308,N_14485);
or U15631 (N_15631,N_14394,N_14256);
or U15632 (N_15632,N_14986,N_14559);
and U15633 (N_15633,N_14221,N_14737);
nor U15634 (N_15634,N_14085,N_14591);
nor U15635 (N_15635,N_14149,N_14990);
or U15636 (N_15636,N_14464,N_14440);
nand U15637 (N_15637,N_14047,N_14384);
nor U15638 (N_15638,N_14175,N_14061);
and U15639 (N_15639,N_14686,N_14797);
nand U15640 (N_15640,N_14966,N_14742);
nor U15641 (N_15641,N_14035,N_14594);
and U15642 (N_15642,N_14735,N_14722);
nand U15643 (N_15643,N_14136,N_14061);
nor U15644 (N_15644,N_14856,N_14044);
nand U15645 (N_15645,N_14428,N_14200);
nand U15646 (N_15646,N_14650,N_14570);
xnor U15647 (N_15647,N_14442,N_14418);
or U15648 (N_15648,N_14757,N_14189);
or U15649 (N_15649,N_14862,N_14888);
xor U15650 (N_15650,N_14402,N_14787);
nand U15651 (N_15651,N_14639,N_14127);
nor U15652 (N_15652,N_14305,N_14350);
nand U15653 (N_15653,N_14845,N_14554);
nand U15654 (N_15654,N_14314,N_14947);
nor U15655 (N_15655,N_14597,N_14794);
xnor U15656 (N_15656,N_14004,N_14477);
or U15657 (N_15657,N_14408,N_14127);
nor U15658 (N_15658,N_14037,N_14062);
or U15659 (N_15659,N_14702,N_14805);
nor U15660 (N_15660,N_14651,N_14104);
xnor U15661 (N_15661,N_14295,N_14634);
or U15662 (N_15662,N_14644,N_14143);
xnor U15663 (N_15663,N_14965,N_14496);
and U15664 (N_15664,N_14342,N_14541);
nor U15665 (N_15665,N_14040,N_14066);
nand U15666 (N_15666,N_14789,N_14262);
nor U15667 (N_15667,N_14309,N_14748);
xnor U15668 (N_15668,N_14772,N_14904);
or U15669 (N_15669,N_14165,N_14635);
nor U15670 (N_15670,N_14997,N_14054);
xor U15671 (N_15671,N_14466,N_14130);
nor U15672 (N_15672,N_14939,N_14020);
xor U15673 (N_15673,N_14816,N_14324);
nand U15674 (N_15674,N_14558,N_14938);
nand U15675 (N_15675,N_14973,N_14143);
or U15676 (N_15676,N_14118,N_14645);
or U15677 (N_15677,N_14101,N_14657);
nand U15678 (N_15678,N_14385,N_14314);
nand U15679 (N_15679,N_14688,N_14105);
nor U15680 (N_15680,N_14384,N_14929);
nand U15681 (N_15681,N_14846,N_14694);
xor U15682 (N_15682,N_14998,N_14630);
nor U15683 (N_15683,N_14295,N_14154);
or U15684 (N_15684,N_14512,N_14425);
nor U15685 (N_15685,N_14245,N_14359);
or U15686 (N_15686,N_14212,N_14640);
and U15687 (N_15687,N_14615,N_14596);
nand U15688 (N_15688,N_14083,N_14858);
nor U15689 (N_15689,N_14050,N_14309);
nor U15690 (N_15690,N_14557,N_14341);
and U15691 (N_15691,N_14284,N_14426);
nor U15692 (N_15692,N_14464,N_14413);
nor U15693 (N_15693,N_14855,N_14352);
and U15694 (N_15694,N_14478,N_14729);
xor U15695 (N_15695,N_14660,N_14817);
nor U15696 (N_15696,N_14097,N_14548);
or U15697 (N_15697,N_14420,N_14621);
nor U15698 (N_15698,N_14127,N_14440);
and U15699 (N_15699,N_14691,N_14549);
nand U15700 (N_15700,N_14048,N_14222);
nand U15701 (N_15701,N_14670,N_14881);
and U15702 (N_15702,N_14186,N_14312);
xor U15703 (N_15703,N_14266,N_14215);
nand U15704 (N_15704,N_14860,N_14175);
or U15705 (N_15705,N_14803,N_14769);
nand U15706 (N_15706,N_14591,N_14152);
or U15707 (N_15707,N_14068,N_14509);
and U15708 (N_15708,N_14909,N_14793);
or U15709 (N_15709,N_14255,N_14574);
nor U15710 (N_15710,N_14947,N_14548);
nor U15711 (N_15711,N_14227,N_14348);
and U15712 (N_15712,N_14248,N_14403);
nand U15713 (N_15713,N_14609,N_14316);
nand U15714 (N_15714,N_14895,N_14389);
xnor U15715 (N_15715,N_14519,N_14304);
nand U15716 (N_15716,N_14945,N_14796);
nand U15717 (N_15717,N_14029,N_14210);
and U15718 (N_15718,N_14311,N_14911);
nand U15719 (N_15719,N_14201,N_14590);
or U15720 (N_15720,N_14785,N_14911);
xor U15721 (N_15721,N_14478,N_14572);
nand U15722 (N_15722,N_14021,N_14202);
xor U15723 (N_15723,N_14326,N_14773);
and U15724 (N_15724,N_14036,N_14775);
or U15725 (N_15725,N_14689,N_14712);
or U15726 (N_15726,N_14236,N_14669);
nand U15727 (N_15727,N_14970,N_14694);
xnor U15728 (N_15728,N_14798,N_14829);
nor U15729 (N_15729,N_14534,N_14963);
nand U15730 (N_15730,N_14881,N_14043);
nand U15731 (N_15731,N_14783,N_14663);
and U15732 (N_15732,N_14202,N_14986);
nand U15733 (N_15733,N_14778,N_14769);
and U15734 (N_15734,N_14354,N_14982);
xnor U15735 (N_15735,N_14379,N_14118);
or U15736 (N_15736,N_14271,N_14604);
and U15737 (N_15737,N_14008,N_14707);
xor U15738 (N_15738,N_14941,N_14833);
xor U15739 (N_15739,N_14281,N_14769);
nand U15740 (N_15740,N_14672,N_14172);
and U15741 (N_15741,N_14652,N_14534);
nor U15742 (N_15742,N_14623,N_14697);
nand U15743 (N_15743,N_14142,N_14739);
and U15744 (N_15744,N_14444,N_14180);
and U15745 (N_15745,N_14150,N_14839);
xor U15746 (N_15746,N_14148,N_14348);
nor U15747 (N_15747,N_14714,N_14230);
and U15748 (N_15748,N_14567,N_14560);
xor U15749 (N_15749,N_14466,N_14066);
xnor U15750 (N_15750,N_14981,N_14189);
xor U15751 (N_15751,N_14516,N_14636);
nand U15752 (N_15752,N_14066,N_14803);
or U15753 (N_15753,N_14927,N_14475);
nand U15754 (N_15754,N_14175,N_14124);
nor U15755 (N_15755,N_14971,N_14481);
xnor U15756 (N_15756,N_14048,N_14393);
xor U15757 (N_15757,N_14147,N_14328);
nor U15758 (N_15758,N_14312,N_14797);
nor U15759 (N_15759,N_14697,N_14702);
and U15760 (N_15760,N_14577,N_14362);
nand U15761 (N_15761,N_14672,N_14777);
and U15762 (N_15762,N_14414,N_14786);
or U15763 (N_15763,N_14465,N_14857);
and U15764 (N_15764,N_14635,N_14307);
nand U15765 (N_15765,N_14973,N_14566);
nor U15766 (N_15766,N_14258,N_14213);
or U15767 (N_15767,N_14838,N_14524);
nor U15768 (N_15768,N_14757,N_14086);
or U15769 (N_15769,N_14730,N_14708);
xnor U15770 (N_15770,N_14918,N_14256);
nand U15771 (N_15771,N_14704,N_14706);
nor U15772 (N_15772,N_14524,N_14503);
nand U15773 (N_15773,N_14844,N_14317);
and U15774 (N_15774,N_14170,N_14570);
nand U15775 (N_15775,N_14031,N_14219);
nand U15776 (N_15776,N_14783,N_14341);
and U15777 (N_15777,N_14365,N_14355);
or U15778 (N_15778,N_14743,N_14035);
and U15779 (N_15779,N_14537,N_14879);
nor U15780 (N_15780,N_14401,N_14711);
or U15781 (N_15781,N_14868,N_14496);
nor U15782 (N_15782,N_14909,N_14925);
or U15783 (N_15783,N_14663,N_14287);
xor U15784 (N_15784,N_14631,N_14974);
and U15785 (N_15785,N_14611,N_14590);
or U15786 (N_15786,N_14800,N_14811);
nand U15787 (N_15787,N_14863,N_14830);
nand U15788 (N_15788,N_14485,N_14180);
nor U15789 (N_15789,N_14932,N_14843);
and U15790 (N_15790,N_14339,N_14327);
xnor U15791 (N_15791,N_14845,N_14023);
nand U15792 (N_15792,N_14880,N_14262);
xor U15793 (N_15793,N_14644,N_14938);
xnor U15794 (N_15794,N_14421,N_14700);
nand U15795 (N_15795,N_14892,N_14308);
or U15796 (N_15796,N_14900,N_14140);
or U15797 (N_15797,N_14684,N_14258);
xnor U15798 (N_15798,N_14118,N_14711);
xnor U15799 (N_15799,N_14723,N_14270);
nor U15800 (N_15800,N_14699,N_14819);
or U15801 (N_15801,N_14829,N_14750);
nor U15802 (N_15802,N_14091,N_14847);
xor U15803 (N_15803,N_14454,N_14023);
and U15804 (N_15804,N_14753,N_14872);
nand U15805 (N_15805,N_14334,N_14491);
xnor U15806 (N_15806,N_14760,N_14821);
and U15807 (N_15807,N_14766,N_14698);
or U15808 (N_15808,N_14046,N_14263);
xor U15809 (N_15809,N_14305,N_14217);
nor U15810 (N_15810,N_14427,N_14548);
nor U15811 (N_15811,N_14636,N_14968);
and U15812 (N_15812,N_14104,N_14010);
nand U15813 (N_15813,N_14964,N_14795);
nor U15814 (N_15814,N_14900,N_14879);
or U15815 (N_15815,N_14089,N_14733);
xnor U15816 (N_15816,N_14265,N_14242);
and U15817 (N_15817,N_14048,N_14200);
and U15818 (N_15818,N_14895,N_14168);
and U15819 (N_15819,N_14821,N_14509);
nand U15820 (N_15820,N_14780,N_14454);
or U15821 (N_15821,N_14387,N_14031);
nand U15822 (N_15822,N_14195,N_14655);
xnor U15823 (N_15823,N_14027,N_14254);
or U15824 (N_15824,N_14862,N_14830);
and U15825 (N_15825,N_14929,N_14497);
and U15826 (N_15826,N_14622,N_14217);
nor U15827 (N_15827,N_14862,N_14387);
nand U15828 (N_15828,N_14473,N_14377);
xnor U15829 (N_15829,N_14823,N_14453);
xor U15830 (N_15830,N_14306,N_14818);
nand U15831 (N_15831,N_14537,N_14320);
and U15832 (N_15832,N_14510,N_14935);
nand U15833 (N_15833,N_14344,N_14964);
or U15834 (N_15834,N_14550,N_14520);
or U15835 (N_15835,N_14317,N_14153);
nor U15836 (N_15836,N_14356,N_14197);
and U15837 (N_15837,N_14852,N_14093);
or U15838 (N_15838,N_14995,N_14773);
nor U15839 (N_15839,N_14304,N_14309);
nor U15840 (N_15840,N_14073,N_14726);
nand U15841 (N_15841,N_14738,N_14010);
or U15842 (N_15842,N_14748,N_14873);
nor U15843 (N_15843,N_14897,N_14344);
nand U15844 (N_15844,N_14402,N_14823);
xnor U15845 (N_15845,N_14745,N_14900);
xor U15846 (N_15846,N_14528,N_14788);
xor U15847 (N_15847,N_14158,N_14651);
nand U15848 (N_15848,N_14861,N_14890);
nand U15849 (N_15849,N_14607,N_14853);
xor U15850 (N_15850,N_14359,N_14505);
or U15851 (N_15851,N_14807,N_14284);
nor U15852 (N_15852,N_14952,N_14809);
or U15853 (N_15853,N_14484,N_14668);
nand U15854 (N_15854,N_14187,N_14691);
nand U15855 (N_15855,N_14866,N_14427);
or U15856 (N_15856,N_14278,N_14914);
nand U15857 (N_15857,N_14462,N_14475);
or U15858 (N_15858,N_14457,N_14727);
xnor U15859 (N_15859,N_14657,N_14887);
xnor U15860 (N_15860,N_14021,N_14392);
and U15861 (N_15861,N_14802,N_14837);
or U15862 (N_15862,N_14108,N_14850);
and U15863 (N_15863,N_14704,N_14150);
nand U15864 (N_15864,N_14153,N_14672);
nor U15865 (N_15865,N_14656,N_14995);
and U15866 (N_15866,N_14145,N_14873);
nand U15867 (N_15867,N_14777,N_14220);
nand U15868 (N_15868,N_14671,N_14043);
and U15869 (N_15869,N_14194,N_14102);
or U15870 (N_15870,N_14655,N_14764);
and U15871 (N_15871,N_14124,N_14593);
and U15872 (N_15872,N_14157,N_14517);
and U15873 (N_15873,N_14799,N_14913);
nand U15874 (N_15874,N_14302,N_14206);
xor U15875 (N_15875,N_14133,N_14674);
or U15876 (N_15876,N_14697,N_14839);
or U15877 (N_15877,N_14531,N_14809);
nor U15878 (N_15878,N_14527,N_14925);
or U15879 (N_15879,N_14151,N_14742);
or U15880 (N_15880,N_14544,N_14190);
or U15881 (N_15881,N_14738,N_14516);
or U15882 (N_15882,N_14489,N_14550);
xnor U15883 (N_15883,N_14748,N_14243);
nand U15884 (N_15884,N_14576,N_14249);
nand U15885 (N_15885,N_14821,N_14545);
xor U15886 (N_15886,N_14059,N_14713);
xor U15887 (N_15887,N_14423,N_14598);
xnor U15888 (N_15888,N_14000,N_14440);
xor U15889 (N_15889,N_14808,N_14169);
and U15890 (N_15890,N_14943,N_14208);
nor U15891 (N_15891,N_14768,N_14412);
and U15892 (N_15892,N_14414,N_14842);
nand U15893 (N_15893,N_14215,N_14280);
nand U15894 (N_15894,N_14383,N_14770);
nand U15895 (N_15895,N_14888,N_14123);
xor U15896 (N_15896,N_14273,N_14810);
or U15897 (N_15897,N_14843,N_14771);
or U15898 (N_15898,N_14368,N_14466);
or U15899 (N_15899,N_14621,N_14606);
nor U15900 (N_15900,N_14785,N_14315);
and U15901 (N_15901,N_14038,N_14218);
or U15902 (N_15902,N_14057,N_14183);
or U15903 (N_15903,N_14783,N_14152);
nor U15904 (N_15904,N_14480,N_14439);
or U15905 (N_15905,N_14607,N_14321);
and U15906 (N_15906,N_14565,N_14724);
nand U15907 (N_15907,N_14369,N_14746);
and U15908 (N_15908,N_14369,N_14676);
xor U15909 (N_15909,N_14857,N_14310);
xnor U15910 (N_15910,N_14633,N_14244);
nor U15911 (N_15911,N_14338,N_14537);
xor U15912 (N_15912,N_14885,N_14887);
xnor U15913 (N_15913,N_14964,N_14384);
nand U15914 (N_15914,N_14961,N_14638);
nand U15915 (N_15915,N_14441,N_14740);
xnor U15916 (N_15916,N_14319,N_14789);
or U15917 (N_15917,N_14011,N_14042);
xnor U15918 (N_15918,N_14028,N_14918);
nor U15919 (N_15919,N_14903,N_14087);
or U15920 (N_15920,N_14502,N_14261);
nand U15921 (N_15921,N_14559,N_14359);
nand U15922 (N_15922,N_14035,N_14324);
nor U15923 (N_15923,N_14571,N_14932);
xnor U15924 (N_15924,N_14247,N_14465);
nor U15925 (N_15925,N_14900,N_14225);
or U15926 (N_15926,N_14196,N_14876);
xor U15927 (N_15927,N_14901,N_14171);
xor U15928 (N_15928,N_14615,N_14821);
or U15929 (N_15929,N_14870,N_14824);
and U15930 (N_15930,N_14860,N_14932);
nor U15931 (N_15931,N_14139,N_14978);
nand U15932 (N_15932,N_14506,N_14680);
nand U15933 (N_15933,N_14958,N_14547);
xor U15934 (N_15934,N_14353,N_14973);
xnor U15935 (N_15935,N_14129,N_14599);
nand U15936 (N_15936,N_14086,N_14972);
or U15937 (N_15937,N_14157,N_14749);
or U15938 (N_15938,N_14900,N_14597);
nand U15939 (N_15939,N_14425,N_14890);
or U15940 (N_15940,N_14466,N_14077);
and U15941 (N_15941,N_14444,N_14469);
nand U15942 (N_15942,N_14755,N_14522);
xnor U15943 (N_15943,N_14235,N_14040);
nand U15944 (N_15944,N_14802,N_14977);
and U15945 (N_15945,N_14720,N_14562);
xnor U15946 (N_15946,N_14371,N_14590);
nand U15947 (N_15947,N_14692,N_14091);
or U15948 (N_15948,N_14522,N_14594);
nand U15949 (N_15949,N_14737,N_14592);
nand U15950 (N_15950,N_14964,N_14893);
or U15951 (N_15951,N_14274,N_14072);
xor U15952 (N_15952,N_14666,N_14062);
nor U15953 (N_15953,N_14839,N_14550);
nor U15954 (N_15954,N_14509,N_14196);
nor U15955 (N_15955,N_14618,N_14869);
and U15956 (N_15956,N_14476,N_14077);
or U15957 (N_15957,N_14630,N_14974);
nor U15958 (N_15958,N_14281,N_14504);
nor U15959 (N_15959,N_14147,N_14092);
xor U15960 (N_15960,N_14226,N_14087);
and U15961 (N_15961,N_14804,N_14191);
nand U15962 (N_15962,N_14598,N_14618);
xor U15963 (N_15963,N_14428,N_14411);
xnor U15964 (N_15964,N_14009,N_14066);
nor U15965 (N_15965,N_14730,N_14232);
nor U15966 (N_15966,N_14935,N_14019);
and U15967 (N_15967,N_14695,N_14222);
or U15968 (N_15968,N_14396,N_14475);
nor U15969 (N_15969,N_14894,N_14209);
and U15970 (N_15970,N_14982,N_14821);
xor U15971 (N_15971,N_14011,N_14930);
nand U15972 (N_15972,N_14634,N_14469);
nor U15973 (N_15973,N_14294,N_14072);
and U15974 (N_15974,N_14687,N_14203);
xor U15975 (N_15975,N_14971,N_14811);
and U15976 (N_15976,N_14203,N_14135);
xor U15977 (N_15977,N_14678,N_14755);
nor U15978 (N_15978,N_14254,N_14569);
and U15979 (N_15979,N_14343,N_14449);
or U15980 (N_15980,N_14429,N_14447);
nand U15981 (N_15981,N_14576,N_14839);
xnor U15982 (N_15982,N_14254,N_14144);
xnor U15983 (N_15983,N_14218,N_14184);
and U15984 (N_15984,N_14691,N_14034);
nor U15985 (N_15985,N_14833,N_14909);
xnor U15986 (N_15986,N_14744,N_14311);
and U15987 (N_15987,N_14436,N_14761);
nand U15988 (N_15988,N_14556,N_14398);
xnor U15989 (N_15989,N_14485,N_14122);
xor U15990 (N_15990,N_14700,N_14339);
nor U15991 (N_15991,N_14733,N_14489);
or U15992 (N_15992,N_14284,N_14691);
xnor U15993 (N_15993,N_14857,N_14405);
xor U15994 (N_15994,N_14514,N_14584);
nor U15995 (N_15995,N_14802,N_14559);
or U15996 (N_15996,N_14791,N_14921);
xnor U15997 (N_15997,N_14503,N_14109);
or U15998 (N_15998,N_14241,N_14983);
nand U15999 (N_15999,N_14083,N_14037);
nand U16000 (N_16000,N_15967,N_15013);
nand U16001 (N_16001,N_15690,N_15851);
and U16002 (N_16002,N_15774,N_15265);
and U16003 (N_16003,N_15442,N_15175);
xor U16004 (N_16004,N_15487,N_15418);
xnor U16005 (N_16005,N_15666,N_15952);
or U16006 (N_16006,N_15773,N_15923);
or U16007 (N_16007,N_15441,N_15722);
or U16008 (N_16008,N_15168,N_15628);
or U16009 (N_16009,N_15671,N_15513);
xor U16010 (N_16010,N_15351,N_15599);
xor U16011 (N_16011,N_15356,N_15314);
nor U16012 (N_16012,N_15656,N_15026);
xor U16013 (N_16013,N_15450,N_15883);
xor U16014 (N_16014,N_15543,N_15360);
or U16015 (N_16015,N_15262,N_15652);
or U16016 (N_16016,N_15367,N_15174);
or U16017 (N_16017,N_15447,N_15151);
and U16018 (N_16018,N_15597,N_15677);
nand U16019 (N_16019,N_15914,N_15377);
nor U16020 (N_16020,N_15925,N_15119);
or U16021 (N_16021,N_15612,N_15226);
xnor U16022 (N_16022,N_15193,N_15985);
or U16023 (N_16023,N_15010,N_15844);
nor U16024 (N_16024,N_15769,N_15427);
nand U16025 (N_16025,N_15782,N_15317);
and U16026 (N_16026,N_15555,N_15104);
xor U16027 (N_16027,N_15517,N_15941);
nor U16028 (N_16028,N_15056,N_15346);
nor U16029 (N_16029,N_15303,N_15281);
nand U16030 (N_16030,N_15827,N_15630);
nand U16031 (N_16031,N_15965,N_15014);
or U16032 (N_16032,N_15839,N_15876);
or U16033 (N_16033,N_15072,N_15412);
nand U16034 (N_16034,N_15768,N_15285);
and U16035 (N_16035,N_15017,N_15287);
xnor U16036 (N_16036,N_15407,N_15223);
xnor U16037 (N_16037,N_15255,N_15926);
nor U16038 (N_16038,N_15638,N_15854);
xor U16039 (N_16039,N_15050,N_15637);
nand U16040 (N_16040,N_15405,N_15519);
nand U16041 (N_16041,N_15887,N_15160);
xor U16042 (N_16042,N_15998,N_15270);
and U16043 (N_16043,N_15000,N_15957);
or U16044 (N_16044,N_15750,N_15188);
xnor U16045 (N_16045,N_15289,N_15847);
or U16046 (N_16046,N_15251,N_15958);
or U16047 (N_16047,N_15640,N_15058);
and U16048 (N_16048,N_15078,N_15059);
nor U16049 (N_16049,N_15974,N_15478);
or U16050 (N_16050,N_15197,N_15538);
nor U16051 (N_16051,N_15855,N_15100);
xor U16052 (N_16052,N_15537,N_15117);
and U16053 (N_16053,N_15269,N_15772);
nor U16054 (N_16054,N_15031,N_15254);
or U16055 (N_16055,N_15872,N_15863);
nand U16056 (N_16056,N_15426,N_15397);
nand U16057 (N_16057,N_15070,N_15027);
and U16058 (N_16058,N_15016,N_15483);
nand U16059 (N_16059,N_15961,N_15704);
nand U16060 (N_16060,N_15749,N_15936);
nor U16061 (N_16061,N_15260,N_15022);
nand U16062 (N_16062,N_15983,N_15569);
xnor U16063 (N_16063,N_15259,N_15329);
xnor U16064 (N_16064,N_15065,N_15869);
nand U16065 (N_16065,N_15499,N_15603);
and U16066 (N_16066,N_15445,N_15614);
nand U16067 (N_16067,N_15176,N_15993);
nand U16068 (N_16068,N_15158,N_15296);
or U16069 (N_16069,N_15906,N_15275);
or U16070 (N_16070,N_15258,N_15336);
nand U16071 (N_16071,N_15102,N_15280);
or U16072 (N_16072,N_15711,N_15837);
nor U16073 (N_16073,N_15292,N_15663);
nand U16074 (N_16074,N_15325,N_15374);
and U16075 (N_16075,N_15978,N_15520);
nor U16076 (N_16076,N_15139,N_15422);
or U16077 (N_16077,N_15803,N_15015);
or U16078 (N_16078,N_15306,N_15387);
nor U16079 (N_16079,N_15910,N_15747);
xor U16080 (N_16080,N_15693,N_15144);
nand U16081 (N_16081,N_15167,N_15786);
xnor U16082 (N_16082,N_15911,N_15766);
nor U16083 (N_16083,N_15846,N_15753);
xor U16084 (N_16084,N_15495,N_15856);
nand U16085 (N_16085,N_15283,N_15890);
and U16086 (N_16086,N_15934,N_15824);
nand U16087 (N_16087,N_15154,N_15865);
and U16088 (N_16088,N_15584,N_15632);
or U16089 (N_16089,N_15834,N_15195);
xnor U16090 (N_16090,N_15436,N_15635);
nor U16091 (N_16091,N_15939,N_15141);
nand U16092 (N_16092,N_15493,N_15045);
and U16093 (N_16093,N_15882,N_15467);
xnor U16094 (N_16094,N_15604,N_15205);
nor U16095 (N_16095,N_15033,N_15326);
and U16096 (N_16096,N_15942,N_15365);
and U16097 (N_16097,N_15217,N_15363);
or U16098 (N_16098,N_15931,N_15562);
nand U16099 (N_16099,N_15778,N_15173);
nor U16100 (N_16100,N_15123,N_15159);
and U16101 (N_16101,N_15540,N_15097);
xnor U16102 (N_16102,N_15049,N_15557);
nand U16103 (N_16103,N_15381,N_15721);
or U16104 (N_16104,N_15162,N_15645);
xor U16105 (N_16105,N_15791,N_15417);
nor U16106 (N_16106,N_15001,N_15596);
nor U16107 (N_16107,N_15145,N_15256);
nor U16108 (N_16108,N_15960,N_15044);
nor U16109 (N_16109,N_15190,N_15691);
nand U16110 (N_16110,N_15651,N_15886);
nor U16111 (N_16111,N_15479,N_15446);
xnor U16112 (N_16112,N_15085,N_15216);
and U16113 (N_16113,N_15528,N_15916);
or U16114 (N_16114,N_15807,N_15725);
or U16115 (N_16115,N_15615,N_15304);
or U16116 (N_16116,N_15634,N_15122);
nor U16117 (N_16117,N_15790,N_15309);
xor U16118 (N_16118,N_15730,N_15763);
and U16119 (N_16119,N_15047,N_15879);
or U16120 (N_16120,N_15054,N_15909);
xnor U16121 (N_16121,N_15115,N_15415);
nor U16122 (N_16122,N_15323,N_15740);
and U16123 (N_16123,N_15491,N_15420);
or U16124 (N_16124,N_15443,N_15613);
or U16125 (N_16125,N_15759,N_15267);
or U16126 (N_16126,N_15500,N_15735);
nand U16127 (N_16127,N_15347,N_15199);
and U16128 (N_16128,N_15813,N_15692);
xor U16129 (N_16129,N_15945,N_15271);
nand U16130 (N_16130,N_15187,N_15130);
nor U16131 (N_16131,N_15482,N_15764);
or U16132 (N_16132,N_15231,N_15522);
and U16133 (N_16133,N_15744,N_15464);
or U16134 (N_16134,N_15378,N_15966);
or U16135 (N_16135,N_15331,N_15274);
xnor U16136 (N_16136,N_15043,N_15496);
and U16137 (N_16137,N_15552,N_15793);
nand U16138 (N_16138,N_15308,N_15515);
or U16139 (N_16139,N_15071,N_15714);
xnor U16140 (N_16140,N_15792,N_15700);
and U16141 (N_16141,N_15781,N_15380);
xnor U16142 (N_16142,N_15787,N_15582);
xor U16143 (N_16143,N_15457,N_15452);
nor U16144 (N_16144,N_15897,N_15155);
and U16145 (N_16145,N_15818,N_15214);
xor U16146 (N_16146,N_15249,N_15776);
and U16147 (N_16147,N_15485,N_15732);
or U16148 (N_16148,N_15239,N_15736);
nand U16149 (N_16149,N_15424,N_15767);
nor U16150 (N_16150,N_15703,N_15196);
and U16151 (N_16151,N_15745,N_15946);
nand U16152 (N_16152,N_15598,N_15111);
nor U16153 (N_16153,N_15578,N_15619);
xnor U16154 (N_16154,N_15040,N_15076);
or U16155 (N_16155,N_15870,N_15060);
xnor U16156 (N_16156,N_15468,N_15607);
and U16157 (N_16157,N_15088,N_15244);
or U16158 (N_16158,N_15211,N_15889);
and U16159 (N_16159,N_15647,N_15293);
xor U16160 (N_16160,N_15246,N_15866);
xor U16161 (N_16161,N_15741,N_15696);
nor U16162 (N_16162,N_15840,N_15042);
or U16163 (N_16163,N_15364,N_15720);
xor U16164 (N_16164,N_15724,N_15206);
or U16165 (N_16165,N_15694,N_15913);
nand U16166 (N_16166,N_15590,N_15177);
and U16167 (N_16167,N_15698,N_15812);
nand U16168 (N_16168,N_15290,N_15083);
xor U16169 (N_16169,N_15497,N_15203);
nand U16170 (N_16170,N_15524,N_15697);
nand U16171 (N_16171,N_15006,N_15874);
xor U16172 (N_16172,N_15460,N_15215);
and U16173 (N_16173,N_15944,N_15621);
or U16174 (N_16174,N_15438,N_15760);
nand U16175 (N_16175,N_15875,N_15069);
or U16176 (N_16176,N_15376,N_15841);
or U16177 (N_16177,N_15298,N_15379);
nand U16178 (N_16178,N_15297,N_15172);
and U16179 (N_16179,N_15370,N_15534);
or U16180 (N_16180,N_15679,N_15324);
or U16181 (N_16181,N_15318,N_15751);
or U16182 (N_16182,N_15814,N_15333);
and U16183 (N_16183,N_15128,N_15976);
nor U16184 (N_16184,N_15316,N_15623);
or U16185 (N_16185,N_15547,N_15218);
or U16186 (N_16186,N_15392,N_15507);
nor U16187 (N_16187,N_15625,N_15660);
nor U16188 (N_16188,N_15579,N_15230);
nand U16189 (N_16189,N_15653,N_15617);
or U16190 (N_16190,N_15575,N_15066);
nor U16191 (N_16191,N_15963,N_15149);
nor U16192 (N_16192,N_15284,N_15899);
nand U16193 (N_16193,N_15109,N_15903);
xnor U16194 (N_16194,N_15166,N_15523);
or U16195 (N_16195,N_15550,N_15848);
xor U16196 (N_16196,N_15224,N_15502);
nor U16197 (N_16197,N_15798,N_15503);
and U16198 (N_16198,N_15797,N_15276);
and U16199 (N_16199,N_15343,N_15454);
or U16200 (N_16200,N_15997,N_15933);
or U16201 (N_16201,N_15439,N_15396);
xor U16202 (N_16202,N_15859,N_15532);
or U16203 (N_16203,N_15194,N_15905);
and U16204 (N_16204,N_15742,N_15340);
nor U16205 (N_16205,N_15877,N_15101);
xor U16206 (N_16206,N_15892,N_15286);
and U16207 (N_16207,N_15968,N_15157);
nand U16208 (N_16208,N_15972,N_15826);
nor U16209 (N_16209,N_15989,N_15871);
and U16210 (N_16210,N_15080,N_15456);
or U16211 (N_16211,N_15535,N_15444);
xor U16212 (N_16212,N_15964,N_15815);
nand U16213 (N_16213,N_15073,N_15935);
nand U16214 (N_16214,N_15036,N_15624);
nor U16215 (N_16215,N_15956,N_15801);
or U16216 (N_16216,N_15408,N_15842);
or U16217 (N_16217,N_15820,N_15981);
and U16218 (N_16218,N_15435,N_15559);
or U16219 (N_16219,N_15352,N_15150);
xor U16220 (N_16220,N_15606,N_15185);
and U16221 (N_16221,N_15400,N_15394);
nor U16222 (N_16222,N_15554,N_15147);
or U16223 (N_16223,N_15930,N_15061);
nor U16224 (N_16224,N_15810,N_15563);
xor U16225 (N_16225,N_15649,N_15170);
and U16226 (N_16226,N_15282,N_15809);
xnor U16227 (N_16227,N_15335,N_15712);
or U16228 (N_16228,N_15646,N_15838);
xor U16229 (N_16229,N_15025,N_15264);
nor U16230 (N_16230,N_15719,N_15095);
nand U16231 (N_16231,N_15542,N_15093);
xor U16232 (N_16232,N_15629,N_15002);
xor U16233 (N_16233,N_15079,N_15587);
nor U16234 (N_16234,N_15204,N_15954);
nor U16235 (N_16235,N_15404,N_15311);
and U16236 (N_16236,N_15734,N_15518);
and U16237 (N_16237,N_15738,N_15473);
xnor U16238 (N_16238,N_15893,N_15052);
or U16239 (N_16239,N_15112,N_15953);
or U16240 (N_16240,N_15191,N_15339);
xnor U16241 (N_16241,N_15928,N_15419);
xnor U16242 (N_16242,N_15683,N_15650);
xnor U16243 (N_16243,N_15067,N_15644);
and U16244 (N_16244,N_15568,N_15526);
or U16245 (N_16245,N_15337,N_15548);
and U16246 (N_16246,N_15146,N_15894);
or U16247 (N_16247,N_15948,N_15811);
or U16248 (N_16248,N_15631,N_15434);
nor U16249 (N_16249,N_15999,N_15682);
or U16250 (N_16250,N_15802,N_15881);
and U16251 (N_16251,N_15561,N_15019);
or U16252 (N_16252,N_15602,N_15429);
nor U16253 (N_16253,N_15577,N_15822);
xor U16254 (N_16254,N_15583,N_15062);
nand U16255 (N_16255,N_15618,N_15009);
nand U16256 (N_16256,N_15743,N_15567);
or U16257 (N_16257,N_15779,N_15761);
or U16258 (N_16258,N_15041,N_15121);
and U16259 (N_16259,N_15390,N_15943);
or U16260 (N_16260,N_15987,N_15137);
xor U16261 (N_16261,N_15636,N_15984);
and U16262 (N_16262,N_15996,N_15279);
nand U16263 (N_16263,N_15472,N_15375);
xor U16264 (N_16264,N_15234,N_15752);
xor U16265 (N_16265,N_15103,N_15701);
or U16266 (N_16266,N_15929,N_15090);
or U16267 (N_16267,N_15951,N_15676);
and U16268 (N_16268,N_15900,N_15564);
xor U16269 (N_16269,N_15754,N_15242);
and U16270 (N_16270,N_15278,N_15973);
nand U16271 (N_16271,N_15924,N_15488);
or U16272 (N_16272,N_15228,N_15475);
or U16273 (N_16273,N_15715,N_15341);
or U16274 (N_16274,N_15180,N_15344);
and U16275 (N_16275,N_15975,N_15867);
and U16276 (N_16276,N_15077,N_15332);
nor U16277 (N_16277,N_15825,N_15084);
nand U16278 (N_16278,N_15371,N_15247);
xnor U16279 (N_16279,N_15669,N_15868);
and U16280 (N_16280,N_15940,N_15560);
nor U16281 (N_16281,N_15573,N_15489);
nor U16282 (N_16282,N_15208,N_15648);
nor U16283 (N_16283,N_15558,N_15695);
or U16284 (N_16284,N_15536,N_15980);
and U16285 (N_16285,N_15108,N_15131);
nor U16286 (N_16286,N_15133,N_15035);
and U16287 (N_16287,N_15678,N_15539);
or U16288 (N_16288,N_15310,N_15135);
and U16289 (N_16289,N_15186,N_15800);
nand U16290 (N_16290,N_15046,N_15169);
nor U16291 (N_16291,N_15585,N_15182);
xor U16292 (N_16292,N_15055,N_15687);
nor U16293 (N_16293,N_15449,N_15248);
and U16294 (N_16294,N_15594,N_15366);
or U16295 (N_16295,N_15739,N_15771);
nor U16296 (N_16296,N_15138,N_15902);
xnor U16297 (N_16297,N_15233,N_15403);
and U16298 (N_16298,N_15416,N_15348);
xnor U16299 (N_16299,N_15428,N_15268);
or U16300 (N_16300,N_15498,N_15570);
and U16301 (N_16301,N_15592,N_15299);
nor U16302 (N_16302,N_15580,N_15470);
nor U16303 (N_16303,N_15857,N_15858);
nand U16304 (N_16304,N_15920,N_15300);
nor U16305 (N_16305,N_15219,N_15992);
nand U16306 (N_16306,N_15081,N_15737);
nand U16307 (N_16307,N_15406,N_15105);
nor U16308 (N_16308,N_15319,N_15880);
or U16309 (N_16309,N_15028,N_15708);
nor U16310 (N_16310,N_15626,N_15023);
nor U16311 (N_16311,N_15639,N_15490);
nor U16312 (N_16312,N_15358,N_15113);
and U16313 (N_16313,N_15124,N_15136);
and U16314 (N_16314,N_15345,N_15451);
xnor U16315 (N_16315,N_15970,N_15153);
or U16316 (N_16316,N_15453,N_15465);
nand U16317 (N_16317,N_15706,N_15142);
nor U16318 (N_16318,N_15589,N_15477);
xor U16319 (N_16319,N_15729,N_15556);
and U16320 (N_16320,N_15288,N_15605);
or U16321 (N_16321,N_15127,N_15029);
xor U16322 (N_16322,N_15235,N_15362);
nor U16323 (N_16323,N_15353,N_15393);
nand U16324 (N_16324,N_15201,N_15852);
nor U16325 (N_16325,N_15238,N_15448);
and U16326 (N_16326,N_15918,N_15225);
nor U16327 (N_16327,N_15202,N_15120);
nor U16328 (N_16328,N_15709,N_15440);
or U16329 (N_16329,N_15674,N_15272);
and U16330 (N_16330,N_15107,N_15295);
nand U16331 (N_16331,N_15633,N_15163);
nor U16332 (N_16332,N_15675,N_15184);
nand U16333 (N_16333,N_15904,N_15659);
or U16334 (N_16334,N_15595,N_15969);
nor U16335 (N_16335,N_15516,N_15302);
nor U16336 (N_16336,N_15183,N_15962);
xor U16337 (N_16337,N_15921,N_15699);
or U16338 (N_16338,N_15252,N_15971);
xor U16339 (N_16339,N_15198,N_15038);
xnor U16340 (N_16340,N_15593,N_15544);
xnor U16341 (N_16341,N_15305,N_15063);
nor U16342 (N_16342,N_15129,N_15571);
nor U16343 (N_16343,N_15783,N_15402);
or U16344 (N_16344,N_15389,N_15094);
or U16345 (N_16345,N_15126,N_15474);
xnor U16346 (N_16346,N_15853,N_15338);
nor U16347 (N_16347,N_15784,N_15034);
and U16348 (N_16348,N_15399,N_15553);
and U16349 (N_16349,N_15257,N_15549);
xor U16350 (N_16350,N_15830,N_15728);
xnor U16351 (N_16351,N_15873,N_15777);
and U16352 (N_16352,N_15134,N_15189);
xor U16353 (N_16353,N_15831,N_15668);
or U16354 (N_16354,N_15501,N_15243);
and U16355 (N_16355,N_15411,N_15600);
and U16356 (N_16356,N_15291,N_15106);
nor U16357 (N_16357,N_15301,N_15221);
or U16358 (N_16358,N_15148,N_15462);
nand U16359 (N_16359,N_15611,N_15461);
and U16360 (N_16360,N_15932,N_15885);
nand U16361 (N_16361,N_15373,N_15591);
or U16362 (N_16362,N_15414,N_15832);
and U16363 (N_16363,N_15616,N_15959);
nor U16364 (N_16364,N_15342,N_15907);
xor U16365 (N_16365,N_15116,N_15012);
or U16366 (N_16366,N_15051,N_15118);
or U16367 (N_16367,N_15756,N_15222);
nor U16368 (N_16368,N_15506,N_15328);
xor U16369 (N_16369,N_15401,N_15096);
nand U16370 (N_16370,N_15512,N_15988);
and U16371 (N_16371,N_15705,N_15261);
and U16372 (N_16372,N_15514,N_15642);
and U16373 (N_16373,N_15808,N_15032);
and U16374 (N_16374,N_15089,N_15327);
xnor U16375 (N_16375,N_15765,N_15008);
nand U16376 (N_16376,N_15836,N_15667);
nor U16377 (N_16377,N_15572,N_15775);
and U16378 (N_16378,N_15850,N_15171);
or U16379 (N_16379,N_15672,N_15086);
nand U16380 (N_16380,N_15207,N_15576);
or U16381 (N_16381,N_15463,N_15357);
nor U16382 (N_16382,N_15082,N_15240);
nor U16383 (N_16383,N_15455,N_15398);
nor U16384 (N_16384,N_15731,N_15670);
nor U16385 (N_16385,N_15210,N_15156);
nor U16386 (N_16386,N_15982,N_15368);
or U16387 (N_16387,N_15817,N_15209);
and U16388 (N_16388,N_15064,N_15164);
nor U16389 (N_16389,N_15213,N_15794);
nand U16390 (N_16390,N_15680,N_15685);
nand U16391 (N_16391,N_15466,N_15785);
and U16392 (N_16392,N_15391,N_15481);
nor U16393 (N_16393,N_15937,N_15132);
nor U16394 (N_16394,N_15266,N_15828);
and U16395 (N_16395,N_15901,N_15661);
nor U16396 (N_16396,N_15527,N_15702);
nor U16397 (N_16397,N_15245,N_15140);
nor U16398 (N_16398,N_15927,N_15229);
xnor U16399 (N_16399,N_15610,N_15891);
and U16400 (N_16400,N_15057,N_15733);
nand U16401 (N_16401,N_15321,N_15277);
or U16402 (N_16402,N_15382,N_15713);
nor U16403 (N_16403,N_15574,N_15908);
nor U16404 (N_16404,N_15717,N_15011);
nand U16405 (N_16405,N_15565,N_15566);
xnor U16406 (N_16406,N_15413,N_15098);
nor U16407 (N_16407,N_15313,N_15114);
and U16408 (N_16408,N_15895,N_15486);
xnor U16409 (N_16409,N_15330,N_15020);
and U16410 (N_16410,N_15684,N_15007);
and U16411 (N_16411,N_15409,N_15806);
and U16412 (N_16412,N_15110,N_15758);
or U16413 (N_16413,N_15322,N_15746);
nor U16414 (N_16414,N_15995,N_15263);
xor U16415 (N_16415,N_15480,N_15864);
and U16416 (N_16416,N_15757,N_15546);
nand U16417 (N_16417,N_15643,N_15586);
and U16418 (N_16418,N_15384,N_15048);
and U16419 (N_16419,N_15152,N_15833);
and U16420 (N_16420,N_15505,N_15074);
xor U16421 (N_16421,N_15253,N_15386);
xnor U16422 (N_16422,N_15125,N_15878);
nor U16423 (N_16423,N_15789,N_15664);
xnor U16424 (N_16424,N_15718,N_15979);
xor U16425 (N_16425,N_15821,N_15410);
xor U16426 (N_16426,N_15030,N_15021);
and U16427 (N_16427,N_15884,N_15250);
and U16428 (N_16428,N_15484,N_15947);
and U16429 (N_16429,N_15654,N_15977);
and U16430 (N_16430,N_15469,N_15385);
nor U16431 (N_16431,N_15723,N_15551);
nor U16432 (N_16432,N_15915,N_15681);
and U16433 (N_16433,N_15545,N_15200);
or U16434 (N_16434,N_15421,N_15541);
nor U16435 (N_16435,N_15430,N_15823);
or U16436 (N_16436,N_15509,N_15657);
and U16437 (N_16437,N_15179,N_15770);
and U16438 (N_16438,N_15504,N_15938);
or U16439 (N_16439,N_15241,N_15608);
nor U16440 (N_16440,N_15780,N_15432);
nor U16441 (N_16441,N_15688,N_15437);
or U16442 (N_16442,N_15431,N_15816);
xnor U16443 (N_16443,N_15227,N_15835);
and U16444 (N_16444,N_15796,N_15220);
nand U16445 (N_16445,N_15994,N_15788);
nor U16446 (N_16446,N_15917,N_15896);
and U16447 (N_16447,N_15039,N_15799);
nand U16448 (N_16448,N_15762,N_15805);
xor U16449 (N_16449,N_15369,N_15307);
and U16450 (N_16450,N_15092,N_15004);
xor U16451 (N_16451,N_15531,N_15087);
xnor U16452 (N_16452,N_15755,N_15726);
nand U16453 (N_16453,N_15143,N_15354);
nor U16454 (N_16454,N_15919,N_15601);
or U16455 (N_16455,N_15003,N_15627);
and U16456 (N_16456,N_15845,N_15425);
or U16457 (N_16457,N_15165,N_15458);
xor U16458 (N_16458,N_15689,N_15622);
xnor U16459 (N_16459,N_15508,N_15581);
nor U16460 (N_16460,N_15053,N_15620);
nor U16461 (N_16461,N_15068,N_15609);
xnor U16462 (N_16462,N_15862,N_15018);
and U16463 (N_16463,N_15349,N_15273);
xnor U16464 (N_16464,N_15510,N_15471);
xor U16465 (N_16465,N_15658,N_15986);
xor U16466 (N_16466,N_15423,N_15099);
or U16467 (N_16467,N_15181,N_15990);
nand U16468 (N_16468,N_15334,N_15991);
or U16469 (N_16469,N_15849,N_15819);
xor U16470 (N_16470,N_15716,N_15388);
nand U16471 (N_16471,N_15949,N_15005);
nand U16472 (N_16472,N_15533,N_15727);
nand U16473 (N_16473,N_15161,N_15037);
or U16474 (N_16474,N_15212,N_15662);
and U16475 (N_16475,N_15860,N_15655);
or U16476 (N_16476,N_15829,N_15075);
nand U16477 (N_16477,N_15494,N_15476);
or U16478 (N_16478,N_15912,N_15372);
nor U16479 (N_16479,N_15511,N_15312);
and U16480 (N_16480,N_15861,N_15315);
xnor U16481 (N_16481,N_15492,N_15359);
xor U16482 (N_16482,N_15192,N_15521);
or U16483 (N_16483,N_15673,N_15888);
and U16484 (N_16484,N_15530,N_15922);
nand U16485 (N_16485,N_15950,N_15383);
or U16486 (N_16486,N_15232,N_15804);
nor U16487 (N_16487,N_15178,N_15641);
xor U16488 (N_16488,N_15320,N_15459);
xor U16489 (N_16489,N_15707,N_15748);
nor U16490 (N_16490,N_15710,N_15843);
or U16491 (N_16491,N_15361,N_15294);
nand U16492 (N_16492,N_15529,N_15395);
nand U16493 (N_16493,N_15236,N_15091);
or U16494 (N_16494,N_15350,N_15588);
or U16495 (N_16495,N_15795,N_15686);
xnor U16496 (N_16496,N_15525,N_15898);
nand U16497 (N_16497,N_15433,N_15024);
and U16498 (N_16498,N_15355,N_15955);
nor U16499 (N_16499,N_15665,N_15237);
and U16500 (N_16500,N_15812,N_15919);
nand U16501 (N_16501,N_15224,N_15607);
or U16502 (N_16502,N_15311,N_15024);
and U16503 (N_16503,N_15318,N_15387);
or U16504 (N_16504,N_15773,N_15043);
or U16505 (N_16505,N_15622,N_15906);
or U16506 (N_16506,N_15650,N_15715);
nand U16507 (N_16507,N_15572,N_15263);
and U16508 (N_16508,N_15739,N_15091);
and U16509 (N_16509,N_15508,N_15930);
nand U16510 (N_16510,N_15687,N_15111);
or U16511 (N_16511,N_15756,N_15577);
and U16512 (N_16512,N_15389,N_15744);
or U16513 (N_16513,N_15411,N_15633);
or U16514 (N_16514,N_15359,N_15257);
xor U16515 (N_16515,N_15196,N_15276);
or U16516 (N_16516,N_15740,N_15395);
and U16517 (N_16517,N_15293,N_15166);
nand U16518 (N_16518,N_15639,N_15917);
nor U16519 (N_16519,N_15032,N_15097);
nand U16520 (N_16520,N_15033,N_15453);
xnor U16521 (N_16521,N_15638,N_15531);
nand U16522 (N_16522,N_15193,N_15245);
or U16523 (N_16523,N_15420,N_15366);
or U16524 (N_16524,N_15753,N_15468);
and U16525 (N_16525,N_15045,N_15900);
nor U16526 (N_16526,N_15874,N_15555);
nor U16527 (N_16527,N_15370,N_15132);
xnor U16528 (N_16528,N_15740,N_15322);
and U16529 (N_16529,N_15249,N_15823);
nor U16530 (N_16530,N_15653,N_15644);
or U16531 (N_16531,N_15222,N_15590);
nand U16532 (N_16532,N_15451,N_15195);
nor U16533 (N_16533,N_15933,N_15638);
and U16534 (N_16534,N_15055,N_15017);
nor U16535 (N_16535,N_15692,N_15410);
xor U16536 (N_16536,N_15988,N_15024);
or U16537 (N_16537,N_15058,N_15457);
xnor U16538 (N_16538,N_15422,N_15216);
and U16539 (N_16539,N_15904,N_15900);
or U16540 (N_16540,N_15487,N_15072);
and U16541 (N_16541,N_15580,N_15126);
xor U16542 (N_16542,N_15199,N_15093);
xnor U16543 (N_16543,N_15576,N_15594);
nand U16544 (N_16544,N_15531,N_15626);
nand U16545 (N_16545,N_15156,N_15819);
xnor U16546 (N_16546,N_15791,N_15853);
or U16547 (N_16547,N_15896,N_15354);
and U16548 (N_16548,N_15519,N_15397);
nand U16549 (N_16549,N_15897,N_15909);
nor U16550 (N_16550,N_15848,N_15935);
or U16551 (N_16551,N_15227,N_15135);
nand U16552 (N_16552,N_15613,N_15940);
nor U16553 (N_16553,N_15621,N_15401);
and U16554 (N_16554,N_15376,N_15976);
and U16555 (N_16555,N_15940,N_15789);
nand U16556 (N_16556,N_15561,N_15918);
and U16557 (N_16557,N_15772,N_15752);
and U16558 (N_16558,N_15935,N_15740);
nand U16559 (N_16559,N_15351,N_15801);
or U16560 (N_16560,N_15948,N_15464);
or U16561 (N_16561,N_15527,N_15517);
or U16562 (N_16562,N_15133,N_15589);
or U16563 (N_16563,N_15630,N_15190);
and U16564 (N_16564,N_15421,N_15011);
or U16565 (N_16565,N_15196,N_15150);
nand U16566 (N_16566,N_15825,N_15000);
nor U16567 (N_16567,N_15890,N_15502);
and U16568 (N_16568,N_15066,N_15921);
xnor U16569 (N_16569,N_15006,N_15464);
xor U16570 (N_16570,N_15377,N_15888);
or U16571 (N_16571,N_15159,N_15797);
nand U16572 (N_16572,N_15523,N_15664);
nor U16573 (N_16573,N_15114,N_15120);
xor U16574 (N_16574,N_15007,N_15107);
and U16575 (N_16575,N_15238,N_15272);
xnor U16576 (N_16576,N_15187,N_15804);
nor U16577 (N_16577,N_15686,N_15811);
xnor U16578 (N_16578,N_15715,N_15792);
and U16579 (N_16579,N_15626,N_15503);
xor U16580 (N_16580,N_15890,N_15562);
xor U16581 (N_16581,N_15102,N_15847);
nand U16582 (N_16582,N_15223,N_15615);
and U16583 (N_16583,N_15365,N_15792);
or U16584 (N_16584,N_15415,N_15631);
and U16585 (N_16585,N_15343,N_15684);
xnor U16586 (N_16586,N_15623,N_15256);
and U16587 (N_16587,N_15856,N_15766);
xnor U16588 (N_16588,N_15388,N_15504);
nor U16589 (N_16589,N_15629,N_15020);
nor U16590 (N_16590,N_15688,N_15916);
nor U16591 (N_16591,N_15947,N_15843);
nor U16592 (N_16592,N_15835,N_15717);
or U16593 (N_16593,N_15438,N_15614);
or U16594 (N_16594,N_15133,N_15150);
nor U16595 (N_16595,N_15375,N_15131);
nand U16596 (N_16596,N_15929,N_15941);
nand U16597 (N_16597,N_15510,N_15759);
and U16598 (N_16598,N_15276,N_15768);
or U16599 (N_16599,N_15934,N_15801);
nor U16600 (N_16600,N_15461,N_15783);
or U16601 (N_16601,N_15024,N_15244);
nand U16602 (N_16602,N_15838,N_15995);
nor U16603 (N_16603,N_15836,N_15886);
and U16604 (N_16604,N_15266,N_15078);
and U16605 (N_16605,N_15261,N_15281);
nand U16606 (N_16606,N_15867,N_15608);
xor U16607 (N_16607,N_15093,N_15791);
or U16608 (N_16608,N_15842,N_15410);
nand U16609 (N_16609,N_15110,N_15290);
nor U16610 (N_16610,N_15206,N_15782);
nor U16611 (N_16611,N_15239,N_15324);
nand U16612 (N_16612,N_15489,N_15051);
and U16613 (N_16613,N_15669,N_15497);
xnor U16614 (N_16614,N_15797,N_15351);
and U16615 (N_16615,N_15399,N_15641);
xor U16616 (N_16616,N_15539,N_15989);
nand U16617 (N_16617,N_15799,N_15022);
or U16618 (N_16618,N_15305,N_15610);
and U16619 (N_16619,N_15462,N_15972);
nor U16620 (N_16620,N_15299,N_15713);
and U16621 (N_16621,N_15524,N_15113);
and U16622 (N_16622,N_15019,N_15267);
or U16623 (N_16623,N_15676,N_15923);
xnor U16624 (N_16624,N_15974,N_15728);
nor U16625 (N_16625,N_15530,N_15639);
and U16626 (N_16626,N_15396,N_15127);
and U16627 (N_16627,N_15523,N_15544);
nor U16628 (N_16628,N_15078,N_15572);
xnor U16629 (N_16629,N_15449,N_15953);
nor U16630 (N_16630,N_15627,N_15623);
nor U16631 (N_16631,N_15457,N_15412);
or U16632 (N_16632,N_15593,N_15920);
or U16633 (N_16633,N_15700,N_15489);
or U16634 (N_16634,N_15016,N_15899);
and U16635 (N_16635,N_15812,N_15012);
or U16636 (N_16636,N_15559,N_15917);
nor U16637 (N_16637,N_15309,N_15734);
or U16638 (N_16638,N_15180,N_15972);
nor U16639 (N_16639,N_15099,N_15828);
nand U16640 (N_16640,N_15090,N_15884);
and U16641 (N_16641,N_15254,N_15726);
or U16642 (N_16642,N_15210,N_15628);
nand U16643 (N_16643,N_15825,N_15324);
nand U16644 (N_16644,N_15564,N_15692);
nand U16645 (N_16645,N_15005,N_15581);
and U16646 (N_16646,N_15812,N_15103);
and U16647 (N_16647,N_15204,N_15620);
xnor U16648 (N_16648,N_15816,N_15130);
nand U16649 (N_16649,N_15194,N_15718);
or U16650 (N_16650,N_15887,N_15990);
and U16651 (N_16651,N_15880,N_15412);
and U16652 (N_16652,N_15697,N_15959);
nor U16653 (N_16653,N_15881,N_15889);
xor U16654 (N_16654,N_15374,N_15140);
nor U16655 (N_16655,N_15076,N_15612);
nand U16656 (N_16656,N_15961,N_15122);
and U16657 (N_16657,N_15675,N_15964);
and U16658 (N_16658,N_15359,N_15136);
nor U16659 (N_16659,N_15661,N_15071);
nor U16660 (N_16660,N_15152,N_15476);
xor U16661 (N_16661,N_15006,N_15027);
xnor U16662 (N_16662,N_15237,N_15964);
nor U16663 (N_16663,N_15875,N_15910);
nor U16664 (N_16664,N_15547,N_15014);
and U16665 (N_16665,N_15994,N_15948);
and U16666 (N_16666,N_15964,N_15928);
nor U16667 (N_16667,N_15651,N_15856);
nor U16668 (N_16668,N_15450,N_15343);
xor U16669 (N_16669,N_15342,N_15468);
xor U16670 (N_16670,N_15119,N_15027);
nor U16671 (N_16671,N_15608,N_15516);
or U16672 (N_16672,N_15649,N_15112);
nand U16673 (N_16673,N_15061,N_15456);
or U16674 (N_16674,N_15236,N_15500);
and U16675 (N_16675,N_15971,N_15508);
nand U16676 (N_16676,N_15709,N_15055);
nor U16677 (N_16677,N_15041,N_15885);
and U16678 (N_16678,N_15711,N_15419);
xnor U16679 (N_16679,N_15776,N_15710);
and U16680 (N_16680,N_15064,N_15973);
nor U16681 (N_16681,N_15578,N_15876);
xor U16682 (N_16682,N_15757,N_15205);
or U16683 (N_16683,N_15130,N_15335);
and U16684 (N_16684,N_15116,N_15693);
xnor U16685 (N_16685,N_15541,N_15171);
or U16686 (N_16686,N_15642,N_15293);
xnor U16687 (N_16687,N_15218,N_15323);
nor U16688 (N_16688,N_15181,N_15056);
xnor U16689 (N_16689,N_15319,N_15383);
nor U16690 (N_16690,N_15946,N_15910);
or U16691 (N_16691,N_15110,N_15871);
xor U16692 (N_16692,N_15179,N_15842);
nand U16693 (N_16693,N_15273,N_15192);
xor U16694 (N_16694,N_15577,N_15316);
nor U16695 (N_16695,N_15369,N_15262);
nor U16696 (N_16696,N_15758,N_15495);
and U16697 (N_16697,N_15752,N_15520);
and U16698 (N_16698,N_15841,N_15829);
xnor U16699 (N_16699,N_15722,N_15696);
nand U16700 (N_16700,N_15768,N_15855);
nor U16701 (N_16701,N_15156,N_15454);
xnor U16702 (N_16702,N_15728,N_15155);
xnor U16703 (N_16703,N_15743,N_15713);
or U16704 (N_16704,N_15450,N_15515);
nand U16705 (N_16705,N_15013,N_15560);
nand U16706 (N_16706,N_15017,N_15390);
xor U16707 (N_16707,N_15069,N_15994);
or U16708 (N_16708,N_15438,N_15158);
or U16709 (N_16709,N_15805,N_15514);
nor U16710 (N_16710,N_15559,N_15412);
or U16711 (N_16711,N_15516,N_15140);
nor U16712 (N_16712,N_15523,N_15692);
xor U16713 (N_16713,N_15964,N_15810);
and U16714 (N_16714,N_15354,N_15344);
nand U16715 (N_16715,N_15757,N_15116);
and U16716 (N_16716,N_15788,N_15368);
nor U16717 (N_16717,N_15455,N_15471);
nor U16718 (N_16718,N_15598,N_15985);
or U16719 (N_16719,N_15538,N_15027);
nand U16720 (N_16720,N_15998,N_15093);
or U16721 (N_16721,N_15492,N_15439);
and U16722 (N_16722,N_15009,N_15706);
and U16723 (N_16723,N_15686,N_15466);
and U16724 (N_16724,N_15711,N_15560);
or U16725 (N_16725,N_15261,N_15616);
nand U16726 (N_16726,N_15900,N_15300);
or U16727 (N_16727,N_15141,N_15434);
nor U16728 (N_16728,N_15514,N_15809);
nand U16729 (N_16729,N_15679,N_15843);
and U16730 (N_16730,N_15210,N_15904);
or U16731 (N_16731,N_15158,N_15168);
and U16732 (N_16732,N_15095,N_15601);
nand U16733 (N_16733,N_15129,N_15276);
nand U16734 (N_16734,N_15487,N_15308);
nand U16735 (N_16735,N_15490,N_15210);
xnor U16736 (N_16736,N_15502,N_15595);
nand U16737 (N_16737,N_15100,N_15340);
or U16738 (N_16738,N_15043,N_15448);
xor U16739 (N_16739,N_15166,N_15739);
nor U16740 (N_16740,N_15647,N_15913);
or U16741 (N_16741,N_15646,N_15886);
or U16742 (N_16742,N_15862,N_15464);
xnor U16743 (N_16743,N_15313,N_15817);
or U16744 (N_16744,N_15020,N_15259);
nand U16745 (N_16745,N_15727,N_15919);
nand U16746 (N_16746,N_15947,N_15377);
and U16747 (N_16747,N_15070,N_15330);
nor U16748 (N_16748,N_15211,N_15446);
and U16749 (N_16749,N_15908,N_15306);
xnor U16750 (N_16750,N_15984,N_15119);
or U16751 (N_16751,N_15982,N_15589);
nor U16752 (N_16752,N_15557,N_15025);
nand U16753 (N_16753,N_15529,N_15277);
or U16754 (N_16754,N_15054,N_15993);
xor U16755 (N_16755,N_15404,N_15160);
and U16756 (N_16756,N_15116,N_15458);
and U16757 (N_16757,N_15967,N_15027);
or U16758 (N_16758,N_15228,N_15924);
nand U16759 (N_16759,N_15038,N_15350);
and U16760 (N_16760,N_15831,N_15888);
or U16761 (N_16761,N_15834,N_15931);
nand U16762 (N_16762,N_15418,N_15519);
or U16763 (N_16763,N_15867,N_15713);
xor U16764 (N_16764,N_15353,N_15747);
nor U16765 (N_16765,N_15803,N_15183);
and U16766 (N_16766,N_15726,N_15411);
or U16767 (N_16767,N_15907,N_15769);
or U16768 (N_16768,N_15195,N_15674);
and U16769 (N_16769,N_15734,N_15340);
nand U16770 (N_16770,N_15870,N_15332);
nand U16771 (N_16771,N_15786,N_15323);
and U16772 (N_16772,N_15829,N_15763);
and U16773 (N_16773,N_15215,N_15012);
and U16774 (N_16774,N_15537,N_15446);
and U16775 (N_16775,N_15568,N_15660);
xor U16776 (N_16776,N_15121,N_15270);
nand U16777 (N_16777,N_15397,N_15145);
xor U16778 (N_16778,N_15595,N_15457);
xnor U16779 (N_16779,N_15984,N_15075);
nor U16780 (N_16780,N_15768,N_15354);
xnor U16781 (N_16781,N_15331,N_15676);
or U16782 (N_16782,N_15723,N_15612);
nor U16783 (N_16783,N_15071,N_15659);
xnor U16784 (N_16784,N_15048,N_15339);
xor U16785 (N_16785,N_15157,N_15006);
or U16786 (N_16786,N_15580,N_15683);
nor U16787 (N_16787,N_15418,N_15701);
or U16788 (N_16788,N_15006,N_15641);
or U16789 (N_16789,N_15678,N_15550);
nand U16790 (N_16790,N_15605,N_15608);
and U16791 (N_16791,N_15369,N_15211);
and U16792 (N_16792,N_15948,N_15664);
nor U16793 (N_16793,N_15788,N_15341);
and U16794 (N_16794,N_15835,N_15846);
or U16795 (N_16795,N_15145,N_15403);
nor U16796 (N_16796,N_15100,N_15207);
or U16797 (N_16797,N_15672,N_15304);
xor U16798 (N_16798,N_15016,N_15714);
xnor U16799 (N_16799,N_15222,N_15992);
nand U16800 (N_16800,N_15074,N_15344);
nand U16801 (N_16801,N_15689,N_15282);
and U16802 (N_16802,N_15351,N_15633);
nand U16803 (N_16803,N_15146,N_15871);
and U16804 (N_16804,N_15336,N_15695);
xnor U16805 (N_16805,N_15400,N_15230);
nand U16806 (N_16806,N_15814,N_15182);
or U16807 (N_16807,N_15082,N_15982);
or U16808 (N_16808,N_15801,N_15247);
and U16809 (N_16809,N_15675,N_15024);
and U16810 (N_16810,N_15744,N_15759);
or U16811 (N_16811,N_15916,N_15229);
and U16812 (N_16812,N_15325,N_15337);
nor U16813 (N_16813,N_15092,N_15857);
nand U16814 (N_16814,N_15356,N_15207);
and U16815 (N_16815,N_15763,N_15169);
nand U16816 (N_16816,N_15144,N_15031);
nand U16817 (N_16817,N_15236,N_15400);
or U16818 (N_16818,N_15658,N_15208);
xnor U16819 (N_16819,N_15466,N_15482);
or U16820 (N_16820,N_15600,N_15037);
or U16821 (N_16821,N_15823,N_15828);
or U16822 (N_16822,N_15447,N_15532);
xor U16823 (N_16823,N_15750,N_15455);
nor U16824 (N_16824,N_15059,N_15275);
and U16825 (N_16825,N_15613,N_15758);
or U16826 (N_16826,N_15199,N_15020);
nand U16827 (N_16827,N_15125,N_15104);
nand U16828 (N_16828,N_15862,N_15994);
nand U16829 (N_16829,N_15309,N_15034);
or U16830 (N_16830,N_15822,N_15965);
or U16831 (N_16831,N_15779,N_15994);
or U16832 (N_16832,N_15705,N_15293);
nor U16833 (N_16833,N_15015,N_15699);
xnor U16834 (N_16834,N_15009,N_15862);
or U16835 (N_16835,N_15333,N_15405);
nor U16836 (N_16836,N_15489,N_15329);
nor U16837 (N_16837,N_15053,N_15401);
nor U16838 (N_16838,N_15847,N_15985);
nor U16839 (N_16839,N_15651,N_15867);
nor U16840 (N_16840,N_15470,N_15407);
xnor U16841 (N_16841,N_15261,N_15128);
or U16842 (N_16842,N_15241,N_15722);
and U16843 (N_16843,N_15322,N_15263);
nor U16844 (N_16844,N_15755,N_15025);
nor U16845 (N_16845,N_15742,N_15776);
nand U16846 (N_16846,N_15239,N_15196);
xnor U16847 (N_16847,N_15455,N_15922);
or U16848 (N_16848,N_15018,N_15196);
nor U16849 (N_16849,N_15689,N_15382);
xnor U16850 (N_16850,N_15307,N_15859);
nor U16851 (N_16851,N_15859,N_15292);
and U16852 (N_16852,N_15825,N_15123);
nand U16853 (N_16853,N_15329,N_15971);
nor U16854 (N_16854,N_15586,N_15454);
or U16855 (N_16855,N_15910,N_15262);
and U16856 (N_16856,N_15729,N_15348);
nor U16857 (N_16857,N_15448,N_15339);
xnor U16858 (N_16858,N_15865,N_15195);
xor U16859 (N_16859,N_15030,N_15977);
or U16860 (N_16860,N_15524,N_15003);
nand U16861 (N_16861,N_15310,N_15659);
and U16862 (N_16862,N_15975,N_15967);
or U16863 (N_16863,N_15668,N_15047);
and U16864 (N_16864,N_15833,N_15298);
nand U16865 (N_16865,N_15891,N_15661);
and U16866 (N_16866,N_15917,N_15441);
xnor U16867 (N_16867,N_15669,N_15256);
nor U16868 (N_16868,N_15814,N_15768);
nor U16869 (N_16869,N_15481,N_15778);
xor U16870 (N_16870,N_15648,N_15331);
xor U16871 (N_16871,N_15254,N_15928);
nor U16872 (N_16872,N_15168,N_15115);
nand U16873 (N_16873,N_15134,N_15716);
or U16874 (N_16874,N_15752,N_15781);
and U16875 (N_16875,N_15177,N_15132);
and U16876 (N_16876,N_15699,N_15037);
nor U16877 (N_16877,N_15567,N_15858);
and U16878 (N_16878,N_15071,N_15379);
xnor U16879 (N_16879,N_15473,N_15257);
xor U16880 (N_16880,N_15302,N_15726);
and U16881 (N_16881,N_15956,N_15176);
and U16882 (N_16882,N_15898,N_15951);
and U16883 (N_16883,N_15227,N_15820);
and U16884 (N_16884,N_15544,N_15363);
and U16885 (N_16885,N_15192,N_15409);
nand U16886 (N_16886,N_15654,N_15004);
nor U16887 (N_16887,N_15067,N_15368);
or U16888 (N_16888,N_15703,N_15993);
nand U16889 (N_16889,N_15873,N_15494);
xor U16890 (N_16890,N_15479,N_15046);
xnor U16891 (N_16891,N_15507,N_15357);
nor U16892 (N_16892,N_15745,N_15266);
and U16893 (N_16893,N_15107,N_15588);
xor U16894 (N_16894,N_15608,N_15287);
nor U16895 (N_16895,N_15995,N_15004);
nand U16896 (N_16896,N_15147,N_15421);
nor U16897 (N_16897,N_15094,N_15285);
xor U16898 (N_16898,N_15286,N_15684);
xnor U16899 (N_16899,N_15109,N_15069);
xor U16900 (N_16900,N_15425,N_15327);
or U16901 (N_16901,N_15984,N_15935);
nor U16902 (N_16902,N_15635,N_15050);
nor U16903 (N_16903,N_15727,N_15217);
and U16904 (N_16904,N_15894,N_15825);
nor U16905 (N_16905,N_15497,N_15198);
nor U16906 (N_16906,N_15146,N_15730);
nand U16907 (N_16907,N_15201,N_15954);
nor U16908 (N_16908,N_15736,N_15217);
and U16909 (N_16909,N_15353,N_15013);
nand U16910 (N_16910,N_15571,N_15333);
or U16911 (N_16911,N_15398,N_15785);
nand U16912 (N_16912,N_15332,N_15392);
or U16913 (N_16913,N_15961,N_15417);
nand U16914 (N_16914,N_15077,N_15677);
nand U16915 (N_16915,N_15226,N_15759);
and U16916 (N_16916,N_15965,N_15745);
nor U16917 (N_16917,N_15172,N_15366);
and U16918 (N_16918,N_15183,N_15900);
xor U16919 (N_16919,N_15780,N_15728);
nand U16920 (N_16920,N_15599,N_15650);
or U16921 (N_16921,N_15481,N_15478);
nand U16922 (N_16922,N_15939,N_15601);
nand U16923 (N_16923,N_15088,N_15498);
or U16924 (N_16924,N_15647,N_15327);
or U16925 (N_16925,N_15932,N_15046);
or U16926 (N_16926,N_15076,N_15605);
or U16927 (N_16927,N_15428,N_15394);
xor U16928 (N_16928,N_15460,N_15113);
xor U16929 (N_16929,N_15138,N_15446);
and U16930 (N_16930,N_15102,N_15282);
and U16931 (N_16931,N_15998,N_15709);
xor U16932 (N_16932,N_15172,N_15934);
nor U16933 (N_16933,N_15034,N_15248);
nand U16934 (N_16934,N_15419,N_15169);
xor U16935 (N_16935,N_15071,N_15002);
nand U16936 (N_16936,N_15247,N_15918);
nand U16937 (N_16937,N_15221,N_15369);
nor U16938 (N_16938,N_15451,N_15117);
or U16939 (N_16939,N_15314,N_15323);
or U16940 (N_16940,N_15786,N_15799);
or U16941 (N_16941,N_15422,N_15251);
and U16942 (N_16942,N_15404,N_15363);
and U16943 (N_16943,N_15842,N_15473);
nor U16944 (N_16944,N_15187,N_15592);
and U16945 (N_16945,N_15936,N_15934);
or U16946 (N_16946,N_15527,N_15666);
nand U16947 (N_16947,N_15550,N_15399);
xnor U16948 (N_16948,N_15624,N_15445);
nor U16949 (N_16949,N_15250,N_15517);
or U16950 (N_16950,N_15637,N_15952);
nor U16951 (N_16951,N_15457,N_15493);
or U16952 (N_16952,N_15664,N_15861);
nand U16953 (N_16953,N_15807,N_15188);
xnor U16954 (N_16954,N_15491,N_15913);
or U16955 (N_16955,N_15194,N_15573);
nor U16956 (N_16956,N_15430,N_15953);
nor U16957 (N_16957,N_15415,N_15228);
or U16958 (N_16958,N_15641,N_15868);
or U16959 (N_16959,N_15777,N_15542);
or U16960 (N_16960,N_15162,N_15175);
and U16961 (N_16961,N_15561,N_15944);
nand U16962 (N_16962,N_15441,N_15116);
nor U16963 (N_16963,N_15232,N_15523);
and U16964 (N_16964,N_15005,N_15394);
and U16965 (N_16965,N_15238,N_15565);
nand U16966 (N_16966,N_15738,N_15277);
nor U16967 (N_16967,N_15104,N_15829);
or U16968 (N_16968,N_15655,N_15054);
and U16969 (N_16969,N_15030,N_15483);
xnor U16970 (N_16970,N_15369,N_15437);
nand U16971 (N_16971,N_15580,N_15448);
and U16972 (N_16972,N_15317,N_15289);
xnor U16973 (N_16973,N_15412,N_15829);
nand U16974 (N_16974,N_15661,N_15978);
and U16975 (N_16975,N_15036,N_15543);
nand U16976 (N_16976,N_15611,N_15799);
and U16977 (N_16977,N_15700,N_15602);
or U16978 (N_16978,N_15727,N_15718);
xor U16979 (N_16979,N_15212,N_15238);
nand U16980 (N_16980,N_15601,N_15937);
xor U16981 (N_16981,N_15438,N_15661);
and U16982 (N_16982,N_15999,N_15415);
nor U16983 (N_16983,N_15655,N_15881);
nor U16984 (N_16984,N_15515,N_15740);
or U16985 (N_16985,N_15998,N_15229);
xnor U16986 (N_16986,N_15205,N_15728);
xnor U16987 (N_16987,N_15261,N_15140);
nand U16988 (N_16988,N_15572,N_15561);
and U16989 (N_16989,N_15437,N_15441);
or U16990 (N_16990,N_15320,N_15380);
or U16991 (N_16991,N_15930,N_15964);
or U16992 (N_16992,N_15701,N_15128);
nand U16993 (N_16993,N_15004,N_15996);
or U16994 (N_16994,N_15577,N_15759);
and U16995 (N_16995,N_15616,N_15826);
and U16996 (N_16996,N_15670,N_15619);
or U16997 (N_16997,N_15950,N_15429);
and U16998 (N_16998,N_15769,N_15399);
xor U16999 (N_16999,N_15406,N_15501);
or U17000 (N_17000,N_16589,N_16969);
nand U17001 (N_17001,N_16242,N_16186);
nand U17002 (N_17002,N_16654,N_16060);
nor U17003 (N_17003,N_16885,N_16605);
and U17004 (N_17004,N_16041,N_16549);
nand U17005 (N_17005,N_16316,N_16446);
nor U17006 (N_17006,N_16964,N_16579);
nor U17007 (N_17007,N_16025,N_16855);
xor U17008 (N_17008,N_16232,N_16521);
nor U17009 (N_17009,N_16235,N_16016);
nor U17010 (N_17010,N_16121,N_16205);
xnor U17011 (N_17011,N_16619,N_16491);
nor U17012 (N_17012,N_16547,N_16126);
nor U17013 (N_17013,N_16601,N_16054);
xnor U17014 (N_17014,N_16865,N_16637);
and U17015 (N_17015,N_16529,N_16762);
nor U17016 (N_17016,N_16785,N_16646);
nand U17017 (N_17017,N_16071,N_16466);
nand U17018 (N_17018,N_16718,N_16449);
nand U17019 (N_17019,N_16586,N_16896);
nand U17020 (N_17020,N_16040,N_16608);
nor U17021 (N_17021,N_16631,N_16151);
xnor U17022 (N_17022,N_16685,N_16663);
nand U17023 (N_17023,N_16781,N_16502);
and U17024 (N_17024,N_16352,N_16972);
and U17025 (N_17025,N_16734,N_16345);
or U17026 (N_17026,N_16015,N_16265);
nor U17027 (N_17027,N_16091,N_16388);
nor U17028 (N_17028,N_16979,N_16409);
and U17029 (N_17029,N_16835,N_16639);
nand U17030 (N_17030,N_16609,N_16776);
nand U17031 (N_17031,N_16123,N_16084);
nor U17032 (N_17032,N_16289,N_16528);
xnor U17033 (N_17033,N_16450,N_16750);
and U17034 (N_17034,N_16523,N_16946);
nand U17035 (N_17035,N_16476,N_16161);
or U17036 (N_17036,N_16806,N_16413);
nor U17037 (N_17037,N_16485,N_16876);
and U17038 (N_17038,N_16249,N_16721);
nand U17039 (N_17039,N_16746,N_16583);
or U17040 (N_17040,N_16005,N_16200);
and U17041 (N_17041,N_16077,N_16907);
or U17042 (N_17042,N_16826,N_16953);
and U17043 (N_17043,N_16974,N_16560);
nand U17044 (N_17044,N_16612,N_16288);
or U17045 (N_17045,N_16083,N_16800);
and U17046 (N_17046,N_16769,N_16195);
or U17047 (N_17047,N_16952,N_16494);
and U17048 (N_17048,N_16606,N_16474);
nand U17049 (N_17049,N_16838,N_16839);
and U17050 (N_17050,N_16758,N_16965);
nand U17051 (N_17051,N_16088,N_16442);
nand U17052 (N_17052,N_16737,N_16498);
and U17053 (N_17053,N_16843,N_16164);
and U17054 (N_17054,N_16698,N_16134);
nor U17055 (N_17055,N_16807,N_16924);
or U17056 (N_17056,N_16338,N_16411);
nor U17057 (N_17057,N_16469,N_16346);
xnor U17058 (N_17058,N_16929,N_16994);
nand U17059 (N_17059,N_16453,N_16683);
nand U17060 (N_17060,N_16157,N_16389);
or U17061 (N_17061,N_16853,N_16185);
nand U17062 (N_17062,N_16640,N_16576);
and U17063 (N_17063,N_16690,N_16173);
xor U17064 (N_17064,N_16234,N_16099);
xnor U17065 (N_17065,N_16496,N_16436);
or U17066 (N_17066,N_16741,N_16543);
nand U17067 (N_17067,N_16271,N_16222);
nor U17068 (N_17068,N_16244,N_16171);
xor U17069 (N_17069,N_16784,N_16977);
nand U17070 (N_17070,N_16699,N_16920);
and U17071 (N_17071,N_16262,N_16796);
xnor U17072 (N_17072,N_16128,N_16405);
xnor U17073 (N_17073,N_16206,N_16532);
and U17074 (N_17074,N_16986,N_16331);
xor U17075 (N_17075,N_16666,N_16537);
or U17076 (N_17076,N_16361,N_16834);
xor U17077 (N_17077,N_16275,N_16792);
and U17078 (N_17078,N_16818,N_16634);
xor U17079 (N_17079,N_16643,N_16849);
xnor U17080 (N_17080,N_16754,N_16153);
and U17081 (N_17081,N_16795,N_16407);
or U17082 (N_17082,N_16517,N_16461);
xor U17083 (N_17083,N_16225,N_16548);
nand U17084 (N_17084,N_16152,N_16678);
or U17085 (N_17085,N_16661,N_16270);
or U17086 (N_17086,N_16836,N_16076);
and U17087 (N_17087,N_16221,N_16044);
xor U17088 (N_17088,N_16653,N_16909);
nand U17089 (N_17089,N_16810,N_16300);
nor U17090 (N_17090,N_16921,N_16651);
or U17091 (N_17091,N_16928,N_16714);
nand U17092 (N_17092,N_16456,N_16421);
and U17093 (N_17093,N_16108,N_16039);
or U17094 (N_17094,N_16854,N_16074);
and U17095 (N_17095,N_16172,N_16914);
xor U17096 (N_17096,N_16752,N_16359);
or U17097 (N_17097,N_16119,N_16933);
or U17098 (N_17098,N_16842,N_16281);
nand U17099 (N_17099,N_16512,N_16910);
and U17100 (N_17100,N_16291,N_16027);
and U17101 (N_17101,N_16382,N_16014);
and U17102 (N_17102,N_16379,N_16958);
or U17103 (N_17103,N_16429,N_16003);
and U17104 (N_17104,N_16012,N_16600);
or U17105 (N_17105,N_16645,N_16423);
and U17106 (N_17106,N_16627,N_16832);
nor U17107 (N_17107,N_16786,N_16577);
nor U17108 (N_17108,N_16742,N_16575);
xor U17109 (N_17109,N_16166,N_16845);
nor U17110 (N_17110,N_16387,N_16918);
nor U17111 (N_17111,N_16192,N_16967);
or U17112 (N_17112,N_16572,N_16727);
or U17113 (N_17113,N_16370,N_16709);
and U17114 (N_17114,N_16046,N_16309);
nand U17115 (N_17115,N_16671,N_16595);
nand U17116 (N_17116,N_16773,N_16793);
or U17117 (N_17117,N_16049,N_16481);
or U17118 (N_17118,N_16757,N_16497);
nor U17119 (N_17119,N_16383,N_16038);
nand U17120 (N_17120,N_16555,N_16542);
xnor U17121 (N_17121,N_16954,N_16694);
nand U17122 (N_17122,N_16692,N_16484);
or U17123 (N_17123,N_16454,N_16550);
nor U17124 (N_17124,N_16304,N_16884);
and U17125 (N_17125,N_16208,N_16238);
nand U17126 (N_17126,N_16169,N_16299);
nand U17127 (N_17127,N_16630,N_16131);
and U17128 (N_17128,N_16592,N_16940);
nand U17129 (N_17129,N_16417,N_16591);
xor U17130 (N_17130,N_16744,N_16691);
and U17131 (N_17131,N_16511,N_16895);
nand U17132 (N_17132,N_16625,N_16522);
xnor U17133 (N_17133,N_16008,N_16889);
or U17134 (N_17134,N_16822,N_16927);
nor U17135 (N_17135,N_16588,N_16216);
nor U17136 (N_17136,N_16023,N_16368);
nor U17137 (N_17137,N_16182,N_16158);
nand U17138 (N_17138,N_16080,N_16859);
xor U17139 (N_17139,N_16990,N_16391);
and U17140 (N_17140,N_16593,N_16086);
xnor U17141 (N_17141,N_16024,N_16725);
and U17142 (N_17142,N_16462,N_16254);
nand U17143 (N_17143,N_16693,N_16156);
or U17144 (N_17144,N_16022,N_16831);
nand U17145 (N_17145,N_16611,N_16312);
and U17146 (N_17146,N_16973,N_16770);
or U17147 (N_17147,N_16505,N_16194);
xor U17148 (N_17148,N_16350,N_16333);
nand U17149 (N_17149,N_16902,N_16351);
nand U17150 (N_17150,N_16059,N_16578);
or U17151 (N_17151,N_16478,N_16688);
nand U17152 (N_17152,N_16410,N_16852);
and U17153 (N_17153,N_16065,N_16679);
nor U17154 (N_17154,N_16129,N_16068);
or U17155 (N_17155,N_16228,N_16327);
xor U17156 (N_17156,N_16418,N_16603);
nand U17157 (N_17157,N_16004,N_16467);
xor U17158 (N_17158,N_16058,N_16841);
nor U17159 (N_17159,N_16212,N_16490);
and U17160 (N_17160,N_16636,N_16525);
and U17161 (N_17161,N_16524,N_16633);
nand U17162 (N_17162,N_16272,N_16148);
xor U17163 (N_17163,N_16697,N_16809);
xnor U17164 (N_17164,N_16115,N_16870);
nor U17165 (N_17165,N_16050,N_16802);
and U17166 (N_17166,N_16302,N_16989);
and U17167 (N_17167,N_16236,N_16133);
xnor U17168 (N_17168,N_16789,N_16251);
nand U17169 (N_17169,N_16749,N_16399);
and U17170 (N_17170,N_16125,N_16064);
and U17171 (N_17171,N_16961,N_16263);
xor U17172 (N_17172,N_16298,N_16787);
and U17173 (N_17173,N_16138,N_16401);
nor U17174 (N_17174,N_16923,N_16402);
nor U17175 (N_17175,N_16808,N_16110);
or U17176 (N_17176,N_16567,N_16486);
nand U17177 (N_17177,N_16011,N_16116);
xor U17178 (N_17178,N_16950,N_16915);
nor U17179 (N_17179,N_16867,N_16030);
xnor U17180 (N_17180,N_16293,N_16712);
or U17181 (N_17181,N_16563,N_16771);
xor U17182 (N_17182,N_16767,N_16294);
xnor U17183 (N_17183,N_16310,N_16955);
xor U17184 (N_17184,N_16167,N_16851);
xor U17185 (N_17185,N_16035,N_16956);
and U17186 (N_17186,N_16297,N_16067);
nor U17187 (N_17187,N_16912,N_16336);
nand U17188 (N_17188,N_16045,N_16573);
nor U17189 (N_17189,N_16878,N_16539);
or U17190 (N_17190,N_16439,N_16947);
xor U17191 (N_17191,N_16477,N_16730);
xnor U17192 (N_17192,N_16620,N_16507);
or U17193 (N_17193,N_16937,N_16193);
and U17194 (N_17194,N_16782,N_16540);
xor U17195 (N_17195,N_16873,N_16819);
nor U17196 (N_17196,N_16629,N_16055);
nand U17197 (N_17197,N_16570,N_16860);
nand U17198 (N_17198,N_16089,N_16279);
nor U17199 (N_17199,N_16901,N_16538);
nand U17200 (N_17200,N_16944,N_16602);
xnor U17201 (N_17201,N_16975,N_16949);
or U17202 (N_17202,N_16061,N_16286);
nor U17203 (N_17203,N_16211,N_16527);
xnor U17204 (N_17204,N_16069,N_16335);
nor U17205 (N_17205,N_16330,N_16136);
nand U17206 (N_17206,N_16638,N_16604);
or U17207 (N_17207,N_16483,N_16874);
nand U17208 (N_17208,N_16564,N_16662);
xnor U17209 (N_17209,N_16400,N_16150);
xnor U17210 (N_17210,N_16991,N_16305);
nor U17211 (N_17211,N_16916,N_16320);
and U17212 (N_17212,N_16034,N_16160);
or U17213 (N_17213,N_16266,N_16245);
and U17214 (N_17214,N_16715,N_16226);
and U17215 (N_17215,N_16743,N_16070);
nor U17216 (N_17216,N_16253,N_16259);
or U17217 (N_17217,N_16021,N_16696);
xnor U17218 (N_17218,N_16881,N_16057);
nand U17219 (N_17219,N_16328,N_16414);
nor U17220 (N_17220,N_16344,N_16203);
nand U17221 (N_17221,N_16376,N_16348);
nand U17222 (N_17222,N_16162,N_16624);
nor U17223 (N_17223,N_16282,N_16551);
nand U17224 (N_17224,N_16287,N_16778);
nor U17225 (N_17225,N_16056,N_16441);
xnor U17226 (N_17226,N_16180,N_16073);
and U17227 (N_17227,N_16188,N_16246);
or U17228 (N_17228,N_16433,N_16105);
nand U17229 (N_17229,N_16541,N_16412);
nand U17230 (N_17230,N_16581,N_16798);
nor U17231 (N_17231,N_16938,N_16117);
or U17232 (N_17232,N_16440,N_16392);
nor U17233 (N_17233,N_16426,N_16465);
nor U17234 (N_17234,N_16553,N_16913);
nand U17235 (N_17235,N_16610,N_16644);
or U17236 (N_17236,N_16170,N_16814);
nor U17237 (N_17237,N_16358,N_16085);
and U17238 (N_17238,N_16777,N_16102);
nor U17239 (N_17239,N_16658,N_16780);
nand U17240 (N_17240,N_16367,N_16660);
and U17241 (N_17241,N_16241,N_16783);
nor U17242 (N_17242,N_16768,N_16506);
nor U17243 (N_17243,N_16319,N_16791);
and U17244 (N_17244,N_16962,N_16616);
or U17245 (N_17245,N_16879,N_16455);
nor U17246 (N_17246,N_16670,N_16536);
nand U17247 (N_17247,N_16648,N_16464);
nand U17248 (N_17248,N_16930,N_16374);
xnor U17249 (N_17249,N_16719,N_16149);
xnor U17250 (N_17250,N_16472,N_16306);
xnor U17251 (N_17251,N_16817,N_16329);
nor U17252 (N_17252,N_16183,N_16710);
nor U17253 (N_17253,N_16393,N_16829);
xor U17254 (N_17254,N_16911,N_16499);
or U17255 (N_17255,N_16628,N_16992);
and U17256 (N_17256,N_16142,N_16104);
nor U17257 (N_17257,N_16354,N_16375);
nand U17258 (N_17258,N_16443,N_16501);
xnor U17259 (N_17259,N_16514,N_16273);
nor U17260 (N_17260,N_16945,N_16764);
nand U17261 (N_17261,N_16903,N_16313);
or U17262 (N_17262,N_16322,N_16480);
nor U17263 (N_17263,N_16130,N_16482);
nor U17264 (N_17264,N_16759,N_16763);
and U17265 (N_17265,N_16231,N_16363);
and U17266 (N_17266,N_16425,N_16794);
nand U17267 (N_17267,N_16120,N_16820);
nor U17268 (N_17268,N_16642,N_16078);
nor U17269 (N_17269,N_16470,N_16284);
nand U17270 (N_17270,N_16580,N_16090);
and U17271 (N_17271,N_16716,N_16428);
and U17272 (N_17272,N_16846,N_16983);
nor U17273 (N_17273,N_16966,N_16202);
and U17274 (N_17274,N_16775,N_16772);
or U17275 (N_17275,N_16504,N_16175);
or U17276 (N_17276,N_16479,N_16621);
nor U17277 (N_17277,N_16599,N_16657);
nor U17278 (N_17278,N_16204,N_16755);
xnor U17279 (N_17279,N_16647,N_16066);
xnor U17280 (N_17280,N_16665,N_16970);
xor U17281 (N_17281,N_16803,N_16676);
nand U17282 (N_17282,N_16364,N_16365);
nand U17283 (N_17283,N_16614,N_16939);
and U17284 (N_17284,N_16571,N_16668);
nand U17285 (N_17285,N_16308,N_16597);
nand U17286 (N_17286,N_16314,N_16176);
nand U17287 (N_17287,N_16520,N_16774);
nor U17288 (N_17288,N_16748,N_16096);
and U17289 (N_17289,N_16159,N_16324);
and U17290 (N_17290,N_16883,N_16706);
or U17291 (N_17291,N_16261,N_16968);
xor U17292 (N_17292,N_16866,N_16075);
xor U17293 (N_17293,N_16799,N_16987);
and U17294 (N_17294,N_16179,N_16165);
and U17295 (N_17295,N_16565,N_16509);
nand U17296 (N_17296,N_16437,N_16135);
nand U17297 (N_17297,N_16850,N_16618);
or U17298 (N_17298,N_16390,N_16558);
nand U17299 (N_17299,N_16394,N_16622);
nand U17300 (N_17300,N_16199,N_16451);
or U17301 (N_17301,N_16029,N_16875);
and U17302 (N_17302,N_16303,N_16406);
xnor U17303 (N_17303,N_16420,N_16111);
and U17304 (N_17304,N_16980,N_16274);
and U17305 (N_17305,N_16147,N_16230);
xor U17306 (N_17306,N_16681,N_16095);
or U17307 (N_17307,N_16317,N_16650);
or U17308 (N_17308,N_16594,N_16861);
or U17309 (N_17309,N_16857,N_16252);
nor U17310 (N_17310,N_16209,N_16936);
nand U17311 (N_17311,N_16386,N_16248);
xnor U17312 (N_17312,N_16037,N_16708);
nor U17313 (N_17313,N_16122,N_16877);
nor U17314 (N_17314,N_16998,N_16283);
or U17315 (N_17315,N_16277,N_16377);
nor U17316 (N_17316,N_16139,N_16174);
nor U17317 (N_17317,N_16043,N_16500);
or U17318 (N_17318,N_16941,N_16276);
or U17319 (N_17319,N_16546,N_16766);
nand U17320 (N_17320,N_16598,N_16756);
xnor U17321 (N_17321,N_16250,N_16184);
or U17322 (N_17322,N_16124,N_16247);
or U17323 (N_17323,N_16711,N_16686);
and U17324 (N_17324,N_16097,N_16471);
and U17325 (N_17325,N_16493,N_16419);
nand U17326 (N_17326,N_16655,N_16143);
or U17327 (N_17327,N_16168,N_16178);
or U17328 (N_17328,N_16761,N_16827);
nand U17329 (N_17329,N_16702,N_16632);
xnor U17330 (N_17330,N_16652,N_16227);
xor U17331 (N_17331,N_16740,N_16726);
nor U17332 (N_17332,N_16347,N_16371);
and U17333 (N_17333,N_16258,N_16201);
nor U17334 (N_17334,N_16243,N_16269);
xnor U17335 (N_17335,N_16978,N_16036);
or U17336 (N_17336,N_16880,N_16848);
or U17337 (N_17337,N_16459,N_16460);
xnor U17338 (N_17338,N_16444,N_16674);
xnor U17339 (N_17339,N_16408,N_16893);
nor U17340 (N_17340,N_16010,N_16519);
xor U17341 (N_17341,N_16863,N_16982);
xor U17342 (N_17342,N_16745,N_16334);
xor U17343 (N_17343,N_16815,N_16042);
and U17344 (N_17344,N_16340,N_16963);
or U17345 (N_17345,N_16475,N_16325);
or U17346 (N_17346,N_16452,N_16140);
xor U17347 (N_17347,N_16109,N_16535);
xor U17348 (N_17348,N_16448,N_16431);
and U17349 (N_17349,N_16118,N_16112);
nand U17350 (N_17350,N_16432,N_16001);
or U17351 (N_17351,N_16062,N_16488);
xor U17352 (N_17352,N_16584,N_16779);
xor U17353 (N_17353,N_16510,N_16033);
xnor U17354 (N_17354,N_16339,N_16240);
or U17355 (N_17355,N_16858,N_16137);
and U17356 (N_17356,N_16864,N_16682);
and U17357 (N_17357,N_16596,N_16380);
and U17358 (N_17358,N_16707,N_16659);
nand U17359 (N_17359,N_16031,N_16704);
or U17360 (N_17360,N_16951,N_16438);
nor U17361 (N_17361,N_16515,N_16720);
or U17362 (N_17362,N_16813,N_16531);
nand U17363 (N_17363,N_16268,N_16106);
nand U17364 (N_17364,N_16887,N_16356);
and U17365 (N_17365,N_16487,N_16569);
or U17366 (N_17366,N_16934,N_16518);
nand U17367 (N_17367,N_16053,N_16385);
and U17368 (N_17368,N_16002,N_16072);
xnor U17369 (N_17369,N_16641,N_16552);
nor U17370 (N_17370,N_16675,N_16526);
and U17371 (N_17371,N_16114,N_16213);
and U17372 (N_17372,N_16415,N_16932);
nand U17373 (N_17373,N_16590,N_16751);
nor U17374 (N_17374,N_16434,N_16957);
or U17375 (N_17375,N_16587,N_16530);
or U17376 (N_17376,N_16020,N_16190);
xnor U17377 (N_17377,N_16669,N_16447);
and U17378 (N_17378,N_16013,N_16871);
and U17379 (N_17379,N_16942,N_16713);
and U17380 (N_17380,N_16559,N_16424);
xnor U17381 (N_17381,N_16700,N_16296);
or U17382 (N_17382,N_16006,N_16366);
nor U17383 (N_17383,N_16705,N_16326);
and U17384 (N_17384,N_16856,N_16664);
or U17385 (N_17385,N_16574,N_16649);
or U17386 (N_17386,N_16191,N_16468);
nor U17387 (N_17387,N_16000,N_16894);
nand U17388 (N_17388,N_16673,N_16557);
nor U17389 (N_17389,N_16948,N_16680);
nor U17390 (N_17390,N_16508,N_16747);
nor U17391 (N_17391,N_16656,N_16256);
or U17392 (N_17392,N_16219,N_16985);
and U17393 (N_17393,N_16398,N_16626);
xor U17394 (N_17394,N_16318,N_16943);
and U17395 (N_17395,N_16739,N_16812);
and U17396 (N_17396,N_16804,N_16396);
nand U17397 (N_17397,N_16753,N_16556);
nand U17398 (N_17398,N_16307,N_16048);
and U17399 (N_17399,N_16931,N_16906);
nor U17400 (N_17400,N_16301,N_16360);
or U17401 (N_17401,N_16292,N_16215);
nand U17402 (N_17402,N_16353,N_16081);
or U17403 (N_17403,N_16919,N_16971);
nand U17404 (N_17404,N_16295,N_16667);
nand U17405 (N_17405,N_16239,N_16738);
nand U17406 (N_17406,N_16100,N_16760);
or U17407 (N_17407,N_16145,N_16092);
nor U17408 (N_17408,N_16458,N_16341);
nand U17409 (N_17409,N_16187,N_16823);
xnor U17410 (N_17410,N_16736,N_16492);
and U17411 (N_17411,N_16224,N_16534);
xor U17412 (N_17412,N_16237,N_16687);
or U17413 (N_17413,N_16290,N_16892);
and U17414 (N_17414,N_16445,N_16397);
xor U17415 (N_17415,N_16891,N_16255);
or U17416 (N_17416,N_16323,N_16554);
and U17417 (N_17417,N_16731,N_16765);
or U17418 (N_17418,N_16132,N_16427);
xor U17419 (N_17419,N_16585,N_16872);
nand U17420 (N_17420,N_16217,N_16198);
xnor U17421 (N_17421,N_16733,N_16908);
nor U17422 (N_17422,N_16533,N_16214);
nand U17423 (N_17423,N_16435,N_16082);
nand U17424 (N_17424,N_16372,N_16144);
nand U17425 (N_17425,N_16051,N_16904);
or U17426 (N_17426,N_16163,N_16028);
xnor U17427 (N_17427,N_16724,N_16993);
nor U17428 (N_17428,N_16196,N_16018);
nand U17429 (N_17429,N_16229,N_16103);
and U17430 (N_17430,N_16900,N_16722);
and U17431 (N_17431,N_16717,N_16922);
nand U17432 (N_17432,N_16960,N_16689);
and U17433 (N_17433,N_16801,N_16473);
or U17434 (N_17434,N_16278,N_16898);
nand U17435 (N_17435,N_16890,N_16189);
nor U17436 (N_17436,N_16107,N_16833);
and U17437 (N_17437,N_16899,N_16218);
and U17438 (N_17438,N_16695,N_16729);
or U17439 (N_17439,N_16797,N_16337);
and U17440 (N_17440,N_16343,N_16561);
or U17441 (N_17441,N_16177,N_16342);
and U17442 (N_17442,N_16355,N_16635);
nand U17443 (N_17443,N_16154,N_16079);
nor U17444 (N_17444,N_16997,N_16888);
and U17445 (N_17445,N_16844,N_16267);
xor U17446 (N_17446,N_16357,N_16463);
nand U17447 (N_17447,N_16223,N_16925);
and U17448 (N_17448,N_16677,N_16732);
nor U17449 (N_17449,N_16422,N_16996);
or U17450 (N_17450,N_16723,N_16009);
nand U17451 (N_17451,N_16617,N_16824);
or U17452 (N_17452,N_16544,N_16830);
nor U17453 (N_17453,N_16790,N_16311);
or U17454 (N_17454,N_16613,N_16052);
nand U17455 (N_17455,N_16260,N_16897);
and U17456 (N_17456,N_16141,N_16381);
nor U17457 (N_17457,N_16207,N_16988);
or U17458 (N_17458,N_16840,N_16384);
nand U17459 (N_17459,N_16430,N_16816);
nand U17460 (N_17460,N_16155,N_16210);
or U17461 (N_17461,N_16811,N_16032);
or U17462 (N_17462,N_16615,N_16181);
nor U17463 (N_17463,N_16562,N_16489);
nor U17464 (N_17464,N_16416,N_16017);
or U17465 (N_17465,N_16369,N_16735);
xnor U17466 (N_17466,N_16959,N_16995);
nor U17467 (N_17467,N_16127,N_16378);
and U17468 (N_17468,N_16926,N_16703);
nor U17469 (N_17469,N_16862,N_16981);
nand U17470 (N_17470,N_16087,N_16197);
or U17471 (N_17471,N_16976,N_16093);
and U17472 (N_17472,N_16280,N_16984);
xor U17473 (N_17473,N_16373,N_16321);
xnor U17474 (N_17474,N_16837,N_16728);
nor U17475 (N_17475,N_16233,N_16566);
and U17476 (N_17476,N_16098,N_16516);
nand U17477 (N_17477,N_16146,N_16905);
and U17478 (N_17478,N_16805,N_16869);
or U17479 (N_17479,N_16825,N_16362);
nor U17480 (N_17480,N_16007,N_16882);
or U17481 (N_17481,N_16220,N_16457);
or U17482 (N_17482,N_16019,N_16063);
xor U17483 (N_17483,N_16886,N_16264);
nand U17484 (N_17484,N_16935,N_16285);
nor U17485 (N_17485,N_16821,N_16999);
xnor U17486 (N_17486,N_16257,N_16315);
xor U17487 (N_17487,N_16607,N_16917);
xnor U17488 (N_17488,N_16701,N_16568);
or U17489 (N_17489,N_16684,N_16788);
nand U17490 (N_17490,N_16582,N_16101);
nor U17491 (N_17491,N_16513,N_16495);
and U17492 (N_17492,N_16545,N_16403);
nand U17493 (N_17493,N_16503,N_16395);
nand U17494 (N_17494,N_16868,N_16094);
nand U17495 (N_17495,N_16623,N_16349);
or U17496 (N_17496,N_16847,N_16026);
and U17497 (N_17497,N_16113,N_16047);
xor U17498 (N_17498,N_16828,N_16332);
nor U17499 (N_17499,N_16672,N_16404);
xor U17500 (N_17500,N_16782,N_16885);
or U17501 (N_17501,N_16641,N_16095);
xnor U17502 (N_17502,N_16195,N_16260);
nand U17503 (N_17503,N_16539,N_16375);
nand U17504 (N_17504,N_16180,N_16395);
xnor U17505 (N_17505,N_16215,N_16305);
and U17506 (N_17506,N_16825,N_16974);
xor U17507 (N_17507,N_16323,N_16584);
or U17508 (N_17508,N_16049,N_16874);
or U17509 (N_17509,N_16815,N_16258);
or U17510 (N_17510,N_16858,N_16892);
xor U17511 (N_17511,N_16674,N_16161);
nor U17512 (N_17512,N_16462,N_16943);
nand U17513 (N_17513,N_16219,N_16706);
or U17514 (N_17514,N_16997,N_16592);
and U17515 (N_17515,N_16402,N_16020);
nor U17516 (N_17516,N_16582,N_16201);
xnor U17517 (N_17517,N_16315,N_16410);
xor U17518 (N_17518,N_16477,N_16833);
nand U17519 (N_17519,N_16172,N_16526);
nor U17520 (N_17520,N_16958,N_16679);
nor U17521 (N_17521,N_16356,N_16776);
nand U17522 (N_17522,N_16021,N_16958);
nor U17523 (N_17523,N_16164,N_16057);
nor U17524 (N_17524,N_16891,N_16277);
nand U17525 (N_17525,N_16298,N_16029);
nand U17526 (N_17526,N_16769,N_16711);
nor U17527 (N_17527,N_16296,N_16382);
nor U17528 (N_17528,N_16205,N_16120);
and U17529 (N_17529,N_16242,N_16158);
nor U17530 (N_17530,N_16021,N_16846);
or U17531 (N_17531,N_16943,N_16665);
nand U17532 (N_17532,N_16547,N_16999);
xnor U17533 (N_17533,N_16226,N_16085);
and U17534 (N_17534,N_16702,N_16838);
nor U17535 (N_17535,N_16913,N_16579);
xnor U17536 (N_17536,N_16932,N_16987);
nor U17537 (N_17537,N_16847,N_16894);
or U17538 (N_17538,N_16040,N_16821);
nand U17539 (N_17539,N_16525,N_16947);
and U17540 (N_17540,N_16957,N_16071);
and U17541 (N_17541,N_16578,N_16789);
and U17542 (N_17542,N_16886,N_16302);
nand U17543 (N_17543,N_16051,N_16271);
and U17544 (N_17544,N_16711,N_16731);
or U17545 (N_17545,N_16961,N_16215);
or U17546 (N_17546,N_16857,N_16440);
xnor U17547 (N_17547,N_16922,N_16238);
or U17548 (N_17548,N_16325,N_16145);
or U17549 (N_17549,N_16645,N_16599);
nand U17550 (N_17550,N_16220,N_16545);
and U17551 (N_17551,N_16538,N_16165);
and U17552 (N_17552,N_16064,N_16798);
or U17553 (N_17553,N_16501,N_16060);
xnor U17554 (N_17554,N_16927,N_16655);
or U17555 (N_17555,N_16226,N_16172);
or U17556 (N_17556,N_16512,N_16029);
nor U17557 (N_17557,N_16378,N_16646);
xor U17558 (N_17558,N_16657,N_16239);
nand U17559 (N_17559,N_16929,N_16910);
and U17560 (N_17560,N_16771,N_16185);
nand U17561 (N_17561,N_16766,N_16949);
nand U17562 (N_17562,N_16626,N_16630);
xnor U17563 (N_17563,N_16124,N_16665);
nor U17564 (N_17564,N_16885,N_16358);
and U17565 (N_17565,N_16509,N_16975);
or U17566 (N_17566,N_16885,N_16329);
nand U17567 (N_17567,N_16504,N_16859);
or U17568 (N_17568,N_16105,N_16417);
nor U17569 (N_17569,N_16357,N_16848);
and U17570 (N_17570,N_16497,N_16814);
xor U17571 (N_17571,N_16355,N_16126);
nor U17572 (N_17572,N_16084,N_16476);
nor U17573 (N_17573,N_16196,N_16666);
and U17574 (N_17574,N_16972,N_16856);
or U17575 (N_17575,N_16836,N_16063);
xor U17576 (N_17576,N_16338,N_16013);
nand U17577 (N_17577,N_16870,N_16269);
xor U17578 (N_17578,N_16389,N_16216);
or U17579 (N_17579,N_16960,N_16519);
and U17580 (N_17580,N_16590,N_16482);
nand U17581 (N_17581,N_16340,N_16700);
nand U17582 (N_17582,N_16119,N_16736);
nor U17583 (N_17583,N_16986,N_16125);
or U17584 (N_17584,N_16890,N_16413);
nor U17585 (N_17585,N_16731,N_16161);
and U17586 (N_17586,N_16388,N_16461);
nor U17587 (N_17587,N_16213,N_16680);
xnor U17588 (N_17588,N_16511,N_16638);
or U17589 (N_17589,N_16033,N_16488);
xor U17590 (N_17590,N_16152,N_16705);
nor U17591 (N_17591,N_16093,N_16667);
and U17592 (N_17592,N_16002,N_16459);
nor U17593 (N_17593,N_16199,N_16782);
or U17594 (N_17594,N_16436,N_16939);
nand U17595 (N_17595,N_16362,N_16785);
and U17596 (N_17596,N_16462,N_16587);
nand U17597 (N_17597,N_16224,N_16808);
or U17598 (N_17598,N_16306,N_16490);
xor U17599 (N_17599,N_16688,N_16563);
xor U17600 (N_17600,N_16067,N_16148);
and U17601 (N_17601,N_16206,N_16213);
nor U17602 (N_17602,N_16392,N_16011);
or U17603 (N_17603,N_16605,N_16058);
or U17604 (N_17604,N_16704,N_16673);
nor U17605 (N_17605,N_16759,N_16366);
nor U17606 (N_17606,N_16121,N_16119);
nor U17607 (N_17607,N_16860,N_16839);
and U17608 (N_17608,N_16843,N_16439);
and U17609 (N_17609,N_16038,N_16408);
and U17610 (N_17610,N_16857,N_16357);
or U17611 (N_17611,N_16534,N_16659);
xor U17612 (N_17612,N_16618,N_16929);
xnor U17613 (N_17613,N_16301,N_16113);
or U17614 (N_17614,N_16585,N_16856);
nor U17615 (N_17615,N_16687,N_16126);
or U17616 (N_17616,N_16865,N_16988);
and U17617 (N_17617,N_16119,N_16603);
xor U17618 (N_17618,N_16178,N_16608);
or U17619 (N_17619,N_16963,N_16348);
and U17620 (N_17620,N_16474,N_16916);
or U17621 (N_17621,N_16414,N_16330);
nand U17622 (N_17622,N_16893,N_16443);
or U17623 (N_17623,N_16672,N_16395);
nor U17624 (N_17624,N_16142,N_16721);
nor U17625 (N_17625,N_16569,N_16080);
or U17626 (N_17626,N_16886,N_16625);
or U17627 (N_17627,N_16535,N_16149);
xor U17628 (N_17628,N_16829,N_16506);
or U17629 (N_17629,N_16816,N_16200);
nor U17630 (N_17630,N_16098,N_16795);
xnor U17631 (N_17631,N_16862,N_16227);
nand U17632 (N_17632,N_16983,N_16505);
xnor U17633 (N_17633,N_16963,N_16515);
xnor U17634 (N_17634,N_16486,N_16272);
nand U17635 (N_17635,N_16689,N_16305);
xnor U17636 (N_17636,N_16921,N_16831);
nor U17637 (N_17637,N_16159,N_16416);
or U17638 (N_17638,N_16440,N_16569);
nor U17639 (N_17639,N_16883,N_16641);
xor U17640 (N_17640,N_16008,N_16726);
xor U17641 (N_17641,N_16144,N_16268);
nor U17642 (N_17642,N_16362,N_16245);
xnor U17643 (N_17643,N_16966,N_16970);
nor U17644 (N_17644,N_16743,N_16424);
nor U17645 (N_17645,N_16360,N_16638);
xnor U17646 (N_17646,N_16338,N_16315);
nor U17647 (N_17647,N_16629,N_16081);
nor U17648 (N_17648,N_16336,N_16154);
or U17649 (N_17649,N_16482,N_16416);
nand U17650 (N_17650,N_16546,N_16221);
xor U17651 (N_17651,N_16198,N_16285);
nor U17652 (N_17652,N_16785,N_16128);
nor U17653 (N_17653,N_16349,N_16266);
nand U17654 (N_17654,N_16047,N_16712);
or U17655 (N_17655,N_16601,N_16134);
or U17656 (N_17656,N_16768,N_16104);
nor U17657 (N_17657,N_16805,N_16360);
and U17658 (N_17658,N_16254,N_16525);
xor U17659 (N_17659,N_16715,N_16560);
xnor U17660 (N_17660,N_16808,N_16924);
nor U17661 (N_17661,N_16730,N_16448);
or U17662 (N_17662,N_16577,N_16234);
and U17663 (N_17663,N_16277,N_16414);
xor U17664 (N_17664,N_16166,N_16884);
nor U17665 (N_17665,N_16131,N_16921);
nand U17666 (N_17666,N_16667,N_16599);
xor U17667 (N_17667,N_16176,N_16351);
xor U17668 (N_17668,N_16646,N_16831);
xor U17669 (N_17669,N_16767,N_16247);
nand U17670 (N_17670,N_16377,N_16515);
nand U17671 (N_17671,N_16179,N_16981);
xnor U17672 (N_17672,N_16524,N_16187);
nand U17673 (N_17673,N_16975,N_16682);
xor U17674 (N_17674,N_16805,N_16573);
xnor U17675 (N_17675,N_16591,N_16024);
nand U17676 (N_17676,N_16427,N_16743);
xor U17677 (N_17677,N_16434,N_16073);
nand U17678 (N_17678,N_16407,N_16815);
nor U17679 (N_17679,N_16449,N_16860);
or U17680 (N_17680,N_16168,N_16526);
nor U17681 (N_17681,N_16887,N_16669);
or U17682 (N_17682,N_16770,N_16719);
and U17683 (N_17683,N_16742,N_16702);
and U17684 (N_17684,N_16605,N_16283);
or U17685 (N_17685,N_16822,N_16771);
nand U17686 (N_17686,N_16233,N_16996);
xor U17687 (N_17687,N_16538,N_16829);
nand U17688 (N_17688,N_16445,N_16755);
xnor U17689 (N_17689,N_16129,N_16628);
nand U17690 (N_17690,N_16465,N_16222);
or U17691 (N_17691,N_16409,N_16253);
nor U17692 (N_17692,N_16985,N_16485);
nand U17693 (N_17693,N_16622,N_16036);
nor U17694 (N_17694,N_16378,N_16158);
and U17695 (N_17695,N_16532,N_16919);
nor U17696 (N_17696,N_16544,N_16223);
nand U17697 (N_17697,N_16495,N_16975);
xnor U17698 (N_17698,N_16792,N_16038);
or U17699 (N_17699,N_16373,N_16179);
nor U17700 (N_17700,N_16526,N_16021);
or U17701 (N_17701,N_16626,N_16950);
xor U17702 (N_17702,N_16591,N_16825);
nor U17703 (N_17703,N_16445,N_16513);
or U17704 (N_17704,N_16321,N_16368);
and U17705 (N_17705,N_16410,N_16821);
or U17706 (N_17706,N_16355,N_16191);
or U17707 (N_17707,N_16942,N_16841);
nand U17708 (N_17708,N_16711,N_16701);
and U17709 (N_17709,N_16380,N_16312);
and U17710 (N_17710,N_16760,N_16133);
xor U17711 (N_17711,N_16354,N_16237);
or U17712 (N_17712,N_16887,N_16281);
nor U17713 (N_17713,N_16409,N_16960);
or U17714 (N_17714,N_16577,N_16874);
xor U17715 (N_17715,N_16231,N_16671);
nor U17716 (N_17716,N_16591,N_16669);
xnor U17717 (N_17717,N_16555,N_16561);
nor U17718 (N_17718,N_16417,N_16004);
or U17719 (N_17719,N_16782,N_16399);
and U17720 (N_17720,N_16974,N_16827);
nor U17721 (N_17721,N_16962,N_16467);
and U17722 (N_17722,N_16287,N_16265);
nand U17723 (N_17723,N_16259,N_16231);
nor U17724 (N_17724,N_16973,N_16139);
nor U17725 (N_17725,N_16764,N_16659);
and U17726 (N_17726,N_16015,N_16310);
and U17727 (N_17727,N_16579,N_16883);
and U17728 (N_17728,N_16464,N_16609);
and U17729 (N_17729,N_16823,N_16748);
nand U17730 (N_17730,N_16327,N_16734);
nor U17731 (N_17731,N_16637,N_16718);
and U17732 (N_17732,N_16505,N_16298);
xnor U17733 (N_17733,N_16613,N_16838);
nor U17734 (N_17734,N_16540,N_16460);
xnor U17735 (N_17735,N_16814,N_16178);
xnor U17736 (N_17736,N_16931,N_16122);
nor U17737 (N_17737,N_16197,N_16462);
and U17738 (N_17738,N_16515,N_16746);
nand U17739 (N_17739,N_16498,N_16729);
and U17740 (N_17740,N_16307,N_16797);
xnor U17741 (N_17741,N_16709,N_16381);
nor U17742 (N_17742,N_16136,N_16650);
and U17743 (N_17743,N_16578,N_16316);
nor U17744 (N_17744,N_16500,N_16714);
or U17745 (N_17745,N_16002,N_16448);
nand U17746 (N_17746,N_16950,N_16545);
or U17747 (N_17747,N_16433,N_16119);
nor U17748 (N_17748,N_16935,N_16692);
nand U17749 (N_17749,N_16779,N_16602);
nor U17750 (N_17750,N_16282,N_16566);
or U17751 (N_17751,N_16684,N_16435);
nand U17752 (N_17752,N_16032,N_16027);
and U17753 (N_17753,N_16981,N_16135);
nor U17754 (N_17754,N_16528,N_16175);
or U17755 (N_17755,N_16193,N_16054);
nand U17756 (N_17756,N_16468,N_16111);
nor U17757 (N_17757,N_16964,N_16253);
or U17758 (N_17758,N_16922,N_16972);
nor U17759 (N_17759,N_16588,N_16948);
or U17760 (N_17760,N_16664,N_16210);
xor U17761 (N_17761,N_16329,N_16594);
nor U17762 (N_17762,N_16139,N_16035);
nand U17763 (N_17763,N_16046,N_16205);
nor U17764 (N_17764,N_16629,N_16203);
and U17765 (N_17765,N_16849,N_16845);
and U17766 (N_17766,N_16479,N_16486);
xnor U17767 (N_17767,N_16972,N_16802);
nor U17768 (N_17768,N_16668,N_16961);
and U17769 (N_17769,N_16811,N_16899);
nor U17770 (N_17770,N_16462,N_16128);
xnor U17771 (N_17771,N_16355,N_16360);
nand U17772 (N_17772,N_16002,N_16954);
nor U17773 (N_17773,N_16023,N_16489);
nor U17774 (N_17774,N_16976,N_16526);
and U17775 (N_17775,N_16017,N_16914);
nand U17776 (N_17776,N_16789,N_16753);
nand U17777 (N_17777,N_16430,N_16448);
nor U17778 (N_17778,N_16294,N_16648);
xnor U17779 (N_17779,N_16516,N_16484);
nand U17780 (N_17780,N_16021,N_16460);
xor U17781 (N_17781,N_16649,N_16423);
and U17782 (N_17782,N_16724,N_16355);
nand U17783 (N_17783,N_16463,N_16483);
nand U17784 (N_17784,N_16675,N_16755);
nor U17785 (N_17785,N_16101,N_16676);
nand U17786 (N_17786,N_16361,N_16723);
nor U17787 (N_17787,N_16153,N_16602);
nor U17788 (N_17788,N_16287,N_16349);
xor U17789 (N_17789,N_16548,N_16181);
and U17790 (N_17790,N_16404,N_16852);
xor U17791 (N_17791,N_16244,N_16238);
nand U17792 (N_17792,N_16484,N_16088);
nand U17793 (N_17793,N_16499,N_16684);
or U17794 (N_17794,N_16918,N_16773);
or U17795 (N_17795,N_16559,N_16040);
xnor U17796 (N_17796,N_16491,N_16666);
or U17797 (N_17797,N_16512,N_16702);
xnor U17798 (N_17798,N_16884,N_16901);
nand U17799 (N_17799,N_16648,N_16999);
nor U17800 (N_17800,N_16682,N_16541);
nor U17801 (N_17801,N_16404,N_16572);
nor U17802 (N_17802,N_16886,N_16253);
xor U17803 (N_17803,N_16639,N_16916);
nand U17804 (N_17804,N_16796,N_16922);
nand U17805 (N_17805,N_16667,N_16209);
xor U17806 (N_17806,N_16031,N_16411);
or U17807 (N_17807,N_16795,N_16605);
xnor U17808 (N_17808,N_16020,N_16621);
or U17809 (N_17809,N_16726,N_16613);
or U17810 (N_17810,N_16383,N_16406);
and U17811 (N_17811,N_16540,N_16711);
nand U17812 (N_17812,N_16253,N_16369);
xnor U17813 (N_17813,N_16541,N_16345);
nor U17814 (N_17814,N_16269,N_16217);
nand U17815 (N_17815,N_16378,N_16246);
xor U17816 (N_17816,N_16334,N_16369);
nand U17817 (N_17817,N_16866,N_16813);
or U17818 (N_17818,N_16460,N_16374);
or U17819 (N_17819,N_16300,N_16334);
xnor U17820 (N_17820,N_16713,N_16952);
nand U17821 (N_17821,N_16446,N_16623);
xnor U17822 (N_17822,N_16504,N_16379);
and U17823 (N_17823,N_16756,N_16704);
nand U17824 (N_17824,N_16175,N_16171);
xor U17825 (N_17825,N_16486,N_16823);
or U17826 (N_17826,N_16130,N_16888);
xor U17827 (N_17827,N_16205,N_16157);
nand U17828 (N_17828,N_16400,N_16362);
nand U17829 (N_17829,N_16923,N_16126);
nor U17830 (N_17830,N_16011,N_16699);
xnor U17831 (N_17831,N_16532,N_16072);
xor U17832 (N_17832,N_16740,N_16644);
nor U17833 (N_17833,N_16712,N_16224);
nor U17834 (N_17834,N_16717,N_16386);
or U17835 (N_17835,N_16000,N_16839);
xnor U17836 (N_17836,N_16382,N_16642);
nor U17837 (N_17837,N_16804,N_16269);
or U17838 (N_17838,N_16321,N_16527);
xnor U17839 (N_17839,N_16844,N_16718);
nor U17840 (N_17840,N_16905,N_16642);
and U17841 (N_17841,N_16144,N_16774);
nand U17842 (N_17842,N_16552,N_16109);
or U17843 (N_17843,N_16659,N_16924);
nor U17844 (N_17844,N_16776,N_16739);
and U17845 (N_17845,N_16143,N_16154);
nor U17846 (N_17846,N_16915,N_16735);
nand U17847 (N_17847,N_16744,N_16002);
nand U17848 (N_17848,N_16896,N_16385);
and U17849 (N_17849,N_16260,N_16368);
nand U17850 (N_17850,N_16700,N_16207);
nor U17851 (N_17851,N_16969,N_16362);
nand U17852 (N_17852,N_16611,N_16236);
or U17853 (N_17853,N_16024,N_16368);
nand U17854 (N_17854,N_16050,N_16742);
and U17855 (N_17855,N_16897,N_16389);
or U17856 (N_17856,N_16074,N_16096);
nand U17857 (N_17857,N_16489,N_16557);
xor U17858 (N_17858,N_16915,N_16884);
nand U17859 (N_17859,N_16364,N_16369);
and U17860 (N_17860,N_16959,N_16153);
nand U17861 (N_17861,N_16263,N_16634);
nor U17862 (N_17862,N_16250,N_16628);
or U17863 (N_17863,N_16336,N_16387);
nor U17864 (N_17864,N_16652,N_16391);
and U17865 (N_17865,N_16088,N_16745);
nor U17866 (N_17866,N_16992,N_16159);
and U17867 (N_17867,N_16913,N_16809);
and U17868 (N_17868,N_16944,N_16301);
xor U17869 (N_17869,N_16109,N_16973);
and U17870 (N_17870,N_16788,N_16277);
nor U17871 (N_17871,N_16889,N_16687);
xor U17872 (N_17872,N_16418,N_16651);
or U17873 (N_17873,N_16110,N_16243);
xnor U17874 (N_17874,N_16489,N_16947);
nor U17875 (N_17875,N_16642,N_16495);
xnor U17876 (N_17876,N_16471,N_16988);
nor U17877 (N_17877,N_16529,N_16576);
nor U17878 (N_17878,N_16983,N_16944);
and U17879 (N_17879,N_16433,N_16746);
nor U17880 (N_17880,N_16987,N_16341);
and U17881 (N_17881,N_16339,N_16180);
xor U17882 (N_17882,N_16889,N_16577);
nand U17883 (N_17883,N_16582,N_16561);
nor U17884 (N_17884,N_16264,N_16082);
or U17885 (N_17885,N_16278,N_16091);
nor U17886 (N_17886,N_16793,N_16039);
nand U17887 (N_17887,N_16184,N_16997);
nand U17888 (N_17888,N_16142,N_16476);
and U17889 (N_17889,N_16878,N_16716);
nor U17890 (N_17890,N_16391,N_16137);
and U17891 (N_17891,N_16802,N_16900);
xor U17892 (N_17892,N_16946,N_16953);
nand U17893 (N_17893,N_16411,N_16295);
and U17894 (N_17894,N_16874,N_16778);
xor U17895 (N_17895,N_16447,N_16346);
xor U17896 (N_17896,N_16680,N_16546);
and U17897 (N_17897,N_16185,N_16184);
and U17898 (N_17898,N_16965,N_16191);
xnor U17899 (N_17899,N_16325,N_16447);
nand U17900 (N_17900,N_16200,N_16221);
xnor U17901 (N_17901,N_16643,N_16673);
nand U17902 (N_17902,N_16269,N_16367);
and U17903 (N_17903,N_16923,N_16657);
nand U17904 (N_17904,N_16067,N_16525);
and U17905 (N_17905,N_16185,N_16088);
nor U17906 (N_17906,N_16939,N_16121);
xor U17907 (N_17907,N_16390,N_16909);
nand U17908 (N_17908,N_16735,N_16453);
and U17909 (N_17909,N_16665,N_16991);
nand U17910 (N_17910,N_16723,N_16887);
and U17911 (N_17911,N_16607,N_16636);
or U17912 (N_17912,N_16477,N_16176);
xor U17913 (N_17913,N_16573,N_16652);
xnor U17914 (N_17914,N_16407,N_16022);
xor U17915 (N_17915,N_16199,N_16502);
nand U17916 (N_17916,N_16522,N_16536);
and U17917 (N_17917,N_16780,N_16321);
xnor U17918 (N_17918,N_16487,N_16026);
and U17919 (N_17919,N_16866,N_16268);
xnor U17920 (N_17920,N_16349,N_16591);
and U17921 (N_17921,N_16799,N_16998);
nor U17922 (N_17922,N_16914,N_16646);
and U17923 (N_17923,N_16460,N_16605);
nand U17924 (N_17924,N_16070,N_16172);
nor U17925 (N_17925,N_16618,N_16664);
nand U17926 (N_17926,N_16456,N_16803);
or U17927 (N_17927,N_16023,N_16733);
nand U17928 (N_17928,N_16265,N_16419);
and U17929 (N_17929,N_16179,N_16785);
xnor U17930 (N_17930,N_16903,N_16222);
nor U17931 (N_17931,N_16333,N_16520);
or U17932 (N_17932,N_16622,N_16009);
or U17933 (N_17933,N_16867,N_16716);
nand U17934 (N_17934,N_16463,N_16763);
nor U17935 (N_17935,N_16346,N_16571);
nand U17936 (N_17936,N_16538,N_16204);
nand U17937 (N_17937,N_16587,N_16134);
and U17938 (N_17938,N_16942,N_16136);
nand U17939 (N_17939,N_16504,N_16368);
nand U17940 (N_17940,N_16162,N_16628);
nor U17941 (N_17941,N_16782,N_16966);
nor U17942 (N_17942,N_16947,N_16431);
and U17943 (N_17943,N_16704,N_16176);
nand U17944 (N_17944,N_16792,N_16500);
nand U17945 (N_17945,N_16224,N_16968);
xor U17946 (N_17946,N_16893,N_16199);
xor U17947 (N_17947,N_16975,N_16559);
nand U17948 (N_17948,N_16421,N_16029);
and U17949 (N_17949,N_16483,N_16290);
nor U17950 (N_17950,N_16073,N_16471);
nand U17951 (N_17951,N_16471,N_16729);
or U17952 (N_17952,N_16159,N_16137);
nor U17953 (N_17953,N_16538,N_16758);
nand U17954 (N_17954,N_16763,N_16668);
or U17955 (N_17955,N_16958,N_16243);
nand U17956 (N_17956,N_16240,N_16221);
nor U17957 (N_17957,N_16508,N_16776);
or U17958 (N_17958,N_16087,N_16953);
xnor U17959 (N_17959,N_16745,N_16636);
and U17960 (N_17960,N_16320,N_16522);
nor U17961 (N_17961,N_16252,N_16296);
xor U17962 (N_17962,N_16929,N_16132);
nor U17963 (N_17963,N_16446,N_16694);
xnor U17964 (N_17964,N_16625,N_16275);
or U17965 (N_17965,N_16811,N_16974);
nor U17966 (N_17966,N_16532,N_16767);
or U17967 (N_17967,N_16478,N_16448);
xor U17968 (N_17968,N_16052,N_16800);
or U17969 (N_17969,N_16356,N_16922);
and U17970 (N_17970,N_16915,N_16330);
nand U17971 (N_17971,N_16192,N_16164);
nand U17972 (N_17972,N_16488,N_16195);
or U17973 (N_17973,N_16158,N_16415);
nor U17974 (N_17974,N_16441,N_16966);
or U17975 (N_17975,N_16188,N_16591);
or U17976 (N_17976,N_16020,N_16891);
xnor U17977 (N_17977,N_16703,N_16943);
and U17978 (N_17978,N_16371,N_16220);
and U17979 (N_17979,N_16457,N_16060);
xor U17980 (N_17980,N_16980,N_16717);
or U17981 (N_17981,N_16928,N_16781);
xnor U17982 (N_17982,N_16386,N_16468);
and U17983 (N_17983,N_16507,N_16094);
nor U17984 (N_17984,N_16748,N_16077);
nor U17985 (N_17985,N_16890,N_16440);
and U17986 (N_17986,N_16378,N_16706);
nor U17987 (N_17987,N_16161,N_16020);
xor U17988 (N_17988,N_16932,N_16864);
xnor U17989 (N_17989,N_16122,N_16621);
xnor U17990 (N_17990,N_16620,N_16474);
or U17991 (N_17991,N_16759,N_16564);
or U17992 (N_17992,N_16625,N_16325);
nand U17993 (N_17993,N_16676,N_16111);
nor U17994 (N_17994,N_16727,N_16461);
or U17995 (N_17995,N_16780,N_16319);
nand U17996 (N_17996,N_16880,N_16491);
and U17997 (N_17997,N_16931,N_16433);
and U17998 (N_17998,N_16366,N_16662);
nand U17999 (N_17999,N_16598,N_16707);
xnor U18000 (N_18000,N_17673,N_17798);
and U18001 (N_18001,N_17781,N_17276);
nand U18002 (N_18002,N_17408,N_17419);
xor U18003 (N_18003,N_17200,N_17790);
and U18004 (N_18004,N_17969,N_17321);
nor U18005 (N_18005,N_17965,N_17873);
or U18006 (N_18006,N_17511,N_17393);
or U18007 (N_18007,N_17545,N_17930);
or U18008 (N_18008,N_17012,N_17436);
and U18009 (N_18009,N_17211,N_17556);
and U18010 (N_18010,N_17663,N_17234);
xor U18011 (N_18011,N_17426,N_17106);
or U18012 (N_18012,N_17523,N_17118);
nand U18013 (N_18013,N_17925,N_17631);
and U18014 (N_18014,N_17461,N_17845);
nor U18015 (N_18015,N_17140,N_17373);
and U18016 (N_18016,N_17616,N_17374);
nor U18017 (N_18017,N_17444,N_17213);
or U18018 (N_18018,N_17108,N_17534);
and U18019 (N_18019,N_17102,N_17991);
or U18020 (N_18020,N_17644,N_17089);
or U18021 (N_18021,N_17271,N_17660);
xnor U18022 (N_18022,N_17195,N_17286);
and U18023 (N_18023,N_17546,N_17875);
xnor U18024 (N_18024,N_17410,N_17893);
nor U18025 (N_18025,N_17957,N_17838);
nor U18026 (N_18026,N_17929,N_17208);
nand U18027 (N_18027,N_17993,N_17273);
or U18028 (N_18028,N_17020,N_17625);
xor U18029 (N_18029,N_17748,N_17265);
xnor U18030 (N_18030,N_17065,N_17127);
nand U18031 (N_18031,N_17695,N_17970);
nand U18032 (N_18032,N_17670,N_17716);
or U18033 (N_18033,N_17192,N_17193);
nand U18034 (N_18034,N_17752,N_17097);
and U18035 (N_18035,N_17242,N_17484);
and U18036 (N_18036,N_17185,N_17285);
nand U18037 (N_18037,N_17817,N_17754);
xor U18038 (N_18038,N_17569,N_17761);
nor U18039 (N_18039,N_17397,N_17221);
and U18040 (N_18040,N_17990,N_17119);
nor U18041 (N_18041,N_17908,N_17633);
xnor U18042 (N_18042,N_17805,N_17721);
and U18043 (N_18043,N_17451,N_17027);
and U18044 (N_18044,N_17601,N_17464);
and U18045 (N_18045,N_17979,N_17826);
xnor U18046 (N_18046,N_17103,N_17650);
xor U18047 (N_18047,N_17771,N_17478);
or U18048 (N_18048,N_17730,N_17096);
xor U18049 (N_18049,N_17704,N_17122);
xor U18050 (N_18050,N_17638,N_17043);
nand U18051 (N_18051,N_17528,N_17225);
xnor U18052 (N_18052,N_17220,N_17914);
and U18053 (N_18053,N_17270,N_17405);
and U18054 (N_18054,N_17927,N_17236);
xnor U18055 (N_18055,N_17376,N_17610);
or U18056 (N_18056,N_17843,N_17597);
nor U18057 (N_18057,N_17542,N_17206);
nand U18058 (N_18058,N_17115,N_17155);
or U18059 (N_18059,N_17057,N_17514);
and U18060 (N_18060,N_17722,N_17627);
nor U18061 (N_18061,N_17300,N_17475);
nand U18062 (N_18062,N_17310,N_17561);
nand U18063 (N_18063,N_17031,N_17825);
nor U18064 (N_18064,N_17256,N_17649);
nor U18065 (N_18065,N_17330,N_17414);
nand U18066 (N_18066,N_17656,N_17022);
nand U18067 (N_18067,N_17949,N_17657);
and U18068 (N_18068,N_17753,N_17009);
nand U18069 (N_18069,N_17053,N_17059);
and U18070 (N_18070,N_17175,N_17974);
xor U18071 (N_18071,N_17674,N_17164);
nor U18072 (N_18072,N_17928,N_17394);
or U18073 (N_18073,N_17341,N_17589);
xnor U18074 (N_18074,N_17223,N_17662);
xor U18075 (N_18075,N_17811,N_17703);
nand U18076 (N_18076,N_17731,N_17897);
or U18077 (N_18077,N_17110,N_17924);
and U18078 (N_18078,N_17622,N_17415);
xnor U18079 (N_18079,N_17564,N_17048);
and U18080 (N_18080,N_17168,N_17254);
xor U18081 (N_18081,N_17086,N_17491);
xor U18082 (N_18082,N_17485,N_17654);
nand U18083 (N_18083,N_17822,N_17462);
or U18084 (N_18084,N_17923,N_17258);
nor U18085 (N_18085,N_17447,N_17284);
nand U18086 (N_18086,N_17715,N_17204);
nand U18087 (N_18087,N_17816,N_17680);
or U18088 (N_18088,N_17350,N_17385);
and U18089 (N_18089,N_17777,N_17372);
nand U18090 (N_18090,N_17227,N_17324);
nor U18091 (N_18091,N_17091,N_17809);
nor U18092 (N_18092,N_17830,N_17418);
or U18093 (N_18093,N_17249,N_17019);
xnor U18094 (N_18094,N_17024,N_17483);
or U18095 (N_18095,N_17591,N_17869);
or U18096 (N_18096,N_17917,N_17603);
and U18097 (N_18097,N_17905,N_17322);
or U18098 (N_18098,N_17919,N_17573);
nor U18099 (N_18099,N_17301,N_17740);
nor U18100 (N_18100,N_17230,N_17335);
nand U18101 (N_18101,N_17782,N_17412);
xor U18102 (N_18102,N_17870,N_17750);
nor U18103 (N_18103,N_17100,N_17723);
xor U18104 (N_18104,N_17634,N_17554);
nand U18105 (N_18105,N_17763,N_17144);
xnor U18106 (N_18106,N_17506,N_17803);
xor U18107 (N_18107,N_17824,N_17686);
nor U18108 (N_18108,N_17567,N_17056);
or U18109 (N_18109,N_17593,N_17378);
xnor U18110 (N_18110,N_17398,N_17614);
or U18111 (N_18111,N_17643,N_17196);
xor U18112 (N_18112,N_17800,N_17689);
nand U18113 (N_18113,N_17712,N_17487);
or U18114 (N_18114,N_17467,N_17862);
and U18115 (N_18115,N_17481,N_17976);
xnor U18116 (N_18116,N_17525,N_17210);
xor U18117 (N_18117,N_17156,N_17309);
or U18118 (N_18118,N_17187,N_17125);
or U18119 (N_18119,N_17146,N_17113);
and U18120 (N_18120,N_17933,N_17456);
xor U18121 (N_18121,N_17519,N_17996);
nor U18122 (N_18122,N_17431,N_17819);
nand U18123 (N_18123,N_17305,N_17596);
nor U18124 (N_18124,N_17190,N_17453);
nand U18125 (N_18125,N_17320,N_17780);
or U18126 (N_18126,N_17263,N_17339);
nand U18127 (N_18127,N_17247,N_17241);
nor U18128 (N_18128,N_17380,N_17920);
xor U18129 (N_18129,N_17222,N_17030);
nor U18130 (N_18130,N_17584,N_17934);
xor U18131 (N_18131,N_17363,N_17445);
or U18132 (N_18132,N_17665,N_17326);
and U18133 (N_18133,N_17912,N_17726);
and U18134 (N_18134,N_17283,N_17961);
or U18135 (N_18135,N_17480,N_17804);
nand U18136 (N_18136,N_17913,N_17183);
and U18137 (N_18137,N_17989,N_17938);
or U18138 (N_18138,N_17666,N_17795);
and U18139 (N_18139,N_17992,N_17422);
nor U18140 (N_18140,N_17401,N_17492);
or U18141 (N_18141,N_17812,N_17717);
nor U18142 (N_18142,N_17571,N_17006);
xnor U18143 (N_18143,N_17972,N_17229);
and U18144 (N_18144,N_17852,N_17831);
nor U18145 (N_18145,N_17818,N_17297);
xor U18146 (N_18146,N_17355,N_17406);
xor U18147 (N_18147,N_17169,N_17797);
and U18148 (N_18148,N_17915,N_17783);
nand U18149 (N_18149,N_17560,N_17964);
nor U18150 (N_18150,N_17667,N_17068);
or U18151 (N_18151,N_17299,N_17944);
nor U18152 (N_18152,N_17742,N_17916);
xor U18153 (N_18153,N_17504,N_17720);
nand U18154 (N_18154,N_17566,N_17025);
xnor U18155 (N_18155,N_17617,N_17038);
and U18156 (N_18156,N_17232,N_17404);
nand U18157 (N_18157,N_17537,N_17147);
and U18158 (N_18158,N_17814,N_17592);
or U18159 (N_18159,N_17312,N_17553);
xor U18160 (N_18160,N_17931,N_17269);
xor U18161 (N_18161,N_17971,N_17706);
nand U18162 (N_18162,N_17774,N_17630);
and U18163 (N_18163,N_17779,N_17865);
nor U18164 (N_18164,N_17527,N_17016);
nor U18165 (N_18165,N_17651,N_17290);
nand U18166 (N_18166,N_17718,N_17294);
or U18167 (N_18167,N_17074,N_17264);
and U18168 (N_18168,N_17037,N_17648);
nor U18169 (N_18169,N_17538,N_17863);
and U18170 (N_18170,N_17946,N_17073);
nor U18171 (N_18171,N_17922,N_17551);
or U18172 (N_18172,N_17864,N_17732);
or U18173 (N_18173,N_17885,N_17116);
nor U18174 (N_18174,N_17375,N_17555);
and U18175 (N_18175,N_17751,N_17757);
nor U18176 (N_18176,N_17792,N_17203);
and U18177 (N_18177,N_17239,N_17951);
nand U18178 (N_18178,N_17623,N_17295);
nor U18179 (N_18179,N_17001,N_17423);
xnor U18180 (N_18180,N_17000,N_17835);
nor U18181 (N_18181,N_17072,N_17582);
or U18182 (N_18182,N_17468,N_17588);
xor U18183 (N_18183,N_17328,N_17936);
nand U18184 (N_18184,N_17980,N_17306);
nor U18185 (N_18185,N_17080,N_17543);
nor U18186 (N_18186,N_17823,N_17942);
and U18187 (N_18187,N_17035,N_17101);
xnor U18188 (N_18188,N_17207,N_17758);
or U18189 (N_18189,N_17984,N_17671);
xor U18190 (N_18190,N_17342,N_17581);
nand U18191 (N_18191,N_17463,N_17063);
nand U18192 (N_18192,N_17815,N_17713);
nor U18193 (N_18193,N_17540,N_17367);
xnor U18194 (N_18194,N_17956,N_17129);
and U18195 (N_18195,N_17386,N_17349);
nand U18196 (N_18196,N_17975,N_17132);
nand U18197 (N_18197,N_17973,N_17500);
or U18198 (N_18198,N_17503,N_17138);
xor U18199 (N_18199,N_17558,N_17871);
nand U18200 (N_18200,N_17259,N_17499);
xnor U18201 (N_18201,N_17252,N_17677);
nand U18202 (N_18202,N_17217,N_17067);
nor U18203 (N_18203,N_17784,N_17085);
nor U18204 (N_18204,N_17711,N_17120);
xnor U18205 (N_18205,N_17766,N_17641);
and U18206 (N_18206,N_17880,N_17600);
or U18207 (N_18207,N_17308,N_17455);
or U18208 (N_18208,N_17215,N_17495);
or U18209 (N_18209,N_17743,N_17281);
nand U18210 (N_18210,N_17435,N_17575);
xor U18211 (N_18211,N_17346,N_17162);
nand U18212 (N_18212,N_17157,N_17148);
xnor U18213 (N_18213,N_17248,N_17796);
nor U18214 (N_18214,N_17847,N_17585);
or U18215 (N_18215,N_17517,N_17608);
nor U18216 (N_18216,N_17997,N_17658);
or U18217 (N_18217,N_17637,N_17998);
xnor U18218 (N_18218,N_17848,N_17382);
xnor U18219 (N_18219,N_17186,N_17521);
nor U18220 (N_18220,N_17457,N_17939);
and U18221 (N_18221,N_17563,N_17010);
nor U18222 (N_18222,N_17676,N_17533);
or U18223 (N_18223,N_17520,N_17329);
nand U18224 (N_18224,N_17738,N_17856);
nand U18225 (N_18225,N_17609,N_17303);
and U18226 (N_18226,N_17531,N_17668);
or U18227 (N_18227,N_17327,N_17632);
nor U18228 (N_18228,N_17262,N_17598);
nor U18229 (N_18229,N_17090,N_17879);
nand U18230 (N_18230,N_17813,N_17081);
nand U18231 (N_18231,N_17449,N_17095);
and U18232 (N_18232,N_17945,N_17692);
or U18233 (N_18233,N_17522,N_17903);
nand U18234 (N_18234,N_17402,N_17443);
or U18235 (N_18235,N_17421,N_17047);
nand U18236 (N_18236,N_17014,N_17510);
and U18237 (N_18237,N_17338,N_17396);
or U18238 (N_18238,N_17189,N_17688);
and U18239 (N_18239,N_17141,N_17770);
nor U18240 (N_18240,N_17243,N_17895);
or U18241 (N_18241,N_17877,N_17371);
nor U18242 (N_18242,N_17586,N_17578);
and U18243 (N_18243,N_17887,N_17105);
nor U18244 (N_18244,N_17734,N_17690);
nor U18245 (N_18245,N_17199,N_17323);
xor U18246 (N_18246,N_17184,N_17383);
and U18247 (N_18247,N_17094,N_17767);
and U18248 (N_18248,N_17906,N_17724);
nor U18249 (N_18249,N_17032,N_17015);
nand U18250 (N_18250,N_17160,N_17550);
xor U18251 (N_18251,N_17182,N_17403);
nor U18252 (N_18252,N_17966,N_17696);
xnor U18253 (N_18253,N_17219,N_17867);
and U18254 (N_18254,N_17725,N_17701);
or U18255 (N_18255,N_17967,N_17868);
xor U18256 (N_18256,N_17749,N_17687);
or U18257 (N_18257,N_17621,N_17708);
nor U18258 (N_18258,N_17489,N_17034);
nor U18259 (N_18259,N_17051,N_17853);
nor U18260 (N_18260,N_17197,N_17982);
xor U18261 (N_18261,N_17054,N_17473);
or U18262 (N_18262,N_17802,N_17890);
nor U18263 (N_18263,N_17594,N_17829);
or U18264 (N_18264,N_17442,N_17710);
or U18265 (N_18265,N_17941,N_17859);
or U18266 (N_18266,N_17245,N_17559);
or U18267 (N_18267,N_17769,N_17036);
or U18268 (N_18268,N_17407,N_17154);
or U18269 (N_18269,N_17151,N_17858);
or U18270 (N_18270,N_17775,N_17505);
nand U18271 (N_18271,N_17250,N_17512);
and U18272 (N_18272,N_17828,N_17181);
and U18273 (N_18273,N_17707,N_17471);
or U18274 (N_18274,N_17785,N_17910);
or U18275 (N_18275,N_17071,N_17679);
nor U18276 (N_18276,N_17883,N_17011);
and U18277 (N_18277,N_17345,N_17469);
nand U18278 (N_18278,N_17678,N_17635);
xor U18279 (N_18279,N_17466,N_17257);
and U18280 (N_18280,N_17159,N_17188);
nand U18281 (N_18281,N_17778,N_17548);
and U18282 (N_18282,N_17166,N_17440);
or U18283 (N_18283,N_17152,N_17891);
nor U18284 (N_18284,N_17296,N_17178);
or U18285 (N_18285,N_17377,N_17420);
or U18286 (N_18286,N_17111,N_17476);
xor U18287 (N_18287,N_17963,N_17524);
nor U18288 (N_18288,N_17334,N_17107);
nand U18289 (N_18289,N_17918,N_17343);
xnor U18290 (N_18290,N_17465,N_17062);
nand U18291 (N_18291,N_17479,N_17502);
or U18292 (N_18292,N_17794,N_17293);
xor U18293 (N_18293,N_17907,N_17358);
nor U18294 (N_18294,N_17493,N_17759);
and U18295 (N_18295,N_17458,N_17488);
or U18296 (N_18296,N_17985,N_17599);
or U18297 (N_18297,N_17066,N_17955);
xor U18298 (N_18298,N_17983,N_17429);
or U18299 (N_18299,N_17552,N_17860);
nor U18300 (N_18300,N_17911,N_17477);
xnor U18301 (N_18301,N_17005,N_17018);
nor U18302 (N_18302,N_17866,N_17801);
xor U18303 (N_18303,N_17709,N_17639);
or U18304 (N_18304,N_17365,N_17126);
nor U18305 (N_18305,N_17216,N_17810);
nor U18306 (N_18306,N_17437,N_17170);
xnor U18307 (N_18307,N_17513,N_17180);
nand U18308 (N_18308,N_17958,N_17368);
nor U18309 (N_18309,N_17727,N_17021);
and U18310 (N_18310,N_17765,N_17557);
nor U18311 (N_18311,N_17900,N_17580);
nand U18312 (N_18312,N_17494,N_17149);
xnor U18313 (N_18313,N_17699,N_17092);
nor U18314 (N_18314,N_17882,N_17729);
xnor U18315 (N_18315,N_17736,N_17700);
xnor U18316 (N_18316,N_17351,N_17139);
or U18317 (N_18317,N_17395,N_17653);
xnor U18318 (N_18318,N_17077,N_17793);
or U18319 (N_18319,N_17082,N_17509);
nand U18320 (N_18320,N_17854,N_17399);
xor U18321 (N_18321,N_17433,N_17233);
and U18322 (N_18322,N_17606,N_17855);
nand U18323 (N_18323,N_17605,N_17516);
or U18324 (N_18324,N_17202,N_17124);
xor U18325 (N_18325,N_17347,N_17611);
xor U18326 (N_18326,N_17515,N_17088);
and U18327 (N_18327,N_17134,N_17109);
and U18328 (N_18328,N_17878,N_17806);
and U18329 (N_18329,N_17172,N_17041);
nor U18330 (N_18330,N_17507,N_17099);
and U18331 (N_18331,N_17776,N_17191);
nand U18332 (N_18332,N_17060,N_17595);
xor U18333 (N_18333,N_17369,N_17874);
xor U18334 (N_18334,N_17104,N_17846);
nand U18335 (N_18335,N_17194,N_17968);
xor U18336 (N_18336,N_17434,N_17645);
nor U18337 (N_18337,N_17612,N_17739);
or U18338 (N_18338,N_17379,N_17799);
xnor U18339 (N_18339,N_17390,N_17719);
nand U18340 (N_18340,N_17307,N_17093);
nor U18341 (N_18341,N_17255,N_17950);
and U18342 (N_18342,N_17583,N_17842);
or U18343 (N_18343,N_17251,N_17055);
xor U18344 (N_18344,N_17460,N_17218);
and U18345 (N_18345,N_17472,N_17360);
or U18346 (N_18346,N_17452,N_17052);
xnor U18347 (N_18347,N_17932,N_17384);
nor U18348 (N_18348,N_17827,N_17058);
or U18349 (N_18349,N_17762,N_17954);
xnor U18350 (N_18350,N_17881,N_17655);
and U18351 (N_18351,N_17112,N_17789);
or U18352 (N_18352,N_17568,N_17661);
or U18353 (N_18353,N_17788,N_17808);
xor U18354 (N_18354,N_17026,N_17470);
and U18355 (N_18355,N_17145,N_17176);
nand U18356 (N_18356,N_17143,N_17896);
or U18357 (N_18357,N_17807,N_17084);
xor U18358 (N_18358,N_17518,N_17987);
xnor U18359 (N_18359,N_17280,N_17231);
or U18360 (N_18360,N_17260,N_17023);
nand U18361 (N_18361,N_17131,N_17205);
nand U18362 (N_18362,N_17901,N_17697);
xnor U18363 (N_18363,N_17246,N_17424);
and U18364 (N_18364,N_17253,N_17045);
xnor U18365 (N_18365,N_17640,N_17174);
nor U18366 (N_18366,N_17508,N_17909);
or U18367 (N_18367,N_17960,N_17574);
xnor U18368 (N_18368,N_17007,N_17237);
xor U18369 (N_18369,N_17576,N_17943);
and U18370 (N_18370,N_17244,N_17008);
nand U18371 (N_18371,N_17275,N_17741);
and U18372 (N_18372,N_17391,N_17228);
nand U18373 (N_18373,N_17267,N_17033);
nor U18374 (N_18374,N_17642,N_17647);
nand U18375 (N_18375,N_17841,N_17133);
nand U18376 (N_18376,N_17142,N_17003);
or U18377 (N_18377,N_17889,N_17570);
xnor U18378 (N_18378,N_17675,N_17318);
or U18379 (N_18379,N_17441,N_17850);
or U18380 (N_18380,N_17044,N_17411);
and U18381 (N_18381,N_17702,N_17694);
or U18382 (N_18382,N_17198,N_17839);
nand U18383 (N_18383,N_17791,N_17620);
xnor U18384 (N_18384,N_17948,N_17413);
or U18385 (N_18385,N_17450,N_17833);
nand U18386 (N_18386,N_17136,N_17544);
nor U18387 (N_18387,N_17167,N_17314);
nand U18388 (N_18388,N_17772,N_17562);
and U18389 (N_18389,N_17636,N_17628);
or U18390 (N_18390,N_17837,N_17547);
or U18391 (N_18391,N_17691,N_17549);
nor U18392 (N_18392,N_17165,N_17438);
nand U18393 (N_18393,N_17004,N_17746);
xnor U18394 (N_18394,N_17040,N_17539);
xor U18395 (N_18395,N_17291,N_17114);
nor U18396 (N_18396,N_17618,N_17304);
xnor U18397 (N_18397,N_17070,N_17177);
nand U18398 (N_18398,N_17130,N_17298);
nand U18399 (N_18399,N_17171,N_17212);
nand U18400 (N_18400,N_17902,N_17947);
and U18401 (N_18401,N_17530,N_17526);
nor U18402 (N_18402,N_17333,N_17619);
and U18403 (N_18403,N_17400,N_17747);
xor U18404 (N_18404,N_17098,N_17268);
nor U18405 (N_18405,N_17075,N_17836);
and U18406 (N_18406,N_17952,N_17209);
nor U18407 (N_18407,N_17629,N_17899);
xnor U18408 (N_18408,N_17361,N_17898);
and U18409 (N_18409,N_17362,N_17459);
and U18410 (N_18410,N_17289,N_17076);
nand U18411 (N_18411,N_17353,N_17786);
nand U18412 (N_18412,N_17049,N_17240);
nand U18413 (N_18413,N_17921,N_17356);
or U18414 (N_18414,N_17937,N_17446);
and U18415 (N_18415,N_17387,N_17064);
or U18416 (N_18416,N_17755,N_17977);
xnor U18417 (N_18417,N_17432,N_17744);
nor U18418 (N_18418,N_17352,N_17613);
nand U18419 (N_18419,N_17735,N_17013);
or U18420 (N_18420,N_17501,N_17123);
or U18421 (N_18421,N_17354,N_17892);
or U18422 (N_18422,N_17364,N_17317);
nand U18423 (N_18423,N_17261,N_17872);
or U18424 (N_18424,N_17565,N_17454);
and U18425 (N_18425,N_17602,N_17953);
or U18426 (N_18426,N_17684,N_17672);
nand U18427 (N_18427,N_17894,N_17849);
xnor U18428 (N_18428,N_17926,N_17201);
or U18429 (N_18429,N_17287,N_17532);
xor U18430 (N_18430,N_17698,N_17029);
nand U18431 (N_18431,N_17173,N_17427);
nand U18432 (N_18432,N_17226,N_17981);
and U18433 (N_18433,N_17482,N_17274);
or U18434 (N_18434,N_17490,N_17417);
and U18435 (N_18435,N_17046,N_17768);
nand U18436 (N_18436,N_17137,N_17760);
and U18437 (N_18437,N_17238,N_17128);
nand U18438 (N_18438,N_17439,N_17028);
xnor U18439 (N_18439,N_17577,N_17388);
and U18440 (N_18440,N_17773,N_17756);
nand U18441 (N_18441,N_17529,N_17316);
and U18442 (N_18442,N_17821,N_17888);
and U18443 (N_18443,N_17940,N_17886);
and U18444 (N_18444,N_17615,N_17117);
nor U18445 (N_18445,N_17135,N_17579);
nor U18446 (N_18446,N_17986,N_17764);
and U18447 (N_18447,N_17039,N_17733);
nor U18448 (N_18448,N_17935,N_17535);
nand U18449 (N_18449,N_17425,N_17179);
nand U18450 (N_18450,N_17087,N_17042);
xnor U18451 (N_18451,N_17496,N_17161);
or U18452 (N_18452,N_17681,N_17282);
and U18453 (N_18453,N_17999,N_17745);
and U18454 (N_18454,N_17652,N_17313);
xor U18455 (N_18455,N_17714,N_17325);
xor U18456 (N_18456,N_17292,N_17683);
or U18457 (N_18457,N_17978,N_17150);
or U18458 (N_18458,N_17359,N_17876);
and U18459 (N_18459,N_17497,N_17448);
nor U18460 (N_18460,N_17607,N_17272);
nor U18461 (N_18461,N_17884,N_17604);
nor U18462 (N_18462,N_17536,N_17348);
and U18463 (N_18463,N_17541,N_17994);
or U18464 (N_18464,N_17079,N_17389);
xnor U18465 (N_18465,N_17962,N_17659);
or U18466 (N_18466,N_17121,N_17311);
xor U18467 (N_18467,N_17904,N_17685);
nand U18468 (N_18468,N_17959,N_17988);
and U18469 (N_18469,N_17820,N_17381);
or U18470 (N_18470,N_17235,N_17834);
or U18471 (N_18471,N_17340,N_17163);
nor U18472 (N_18472,N_17844,N_17153);
and U18473 (N_18473,N_17158,N_17995);
xor U18474 (N_18474,N_17279,N_17486);
nand U18475 (N_18475,N_17069,N_17288);
nand U18476 (N_18476,N_17693,N_17857);
nor U18477 (N_18477,N_17277,N_17428);
and U18478 (N_18478,N_17370,N_17266);
or U18479 (N_18479,N_17728,N_17705);
nor U18480 (N_18480,N_17315,N_17017);
nor U18481 (N_18481,N_17409,N_17416);
nor U18482 (N_18482,N_17669,N_17861);
or U18483 (N_18483,N_17646,N_17337);
nor U18484 (N_18484,N_17840,N_17050);
nand U18485 (N_18485,N_17278,N_17302);
or U18486 (N_18486,N_17214,N_17332);
or U18487 (N_18487,N_17832,N_17344);
or U18488 (N_18488,N_17664,N_17083);
xnor U18489 (N_18489,N_17851,N_17626);
xnor U18490 (N_18490,N_17474,N_17357);
or U18491 (N_18491,N_17061,N_17737);
and U18492 (N_18492,N_17587,N_17430);
and U18493 (N_18493,N_17787,N_17319);
xor U18494 (N_18494,N_17336,N_17078);
xnor U18495 (N_18495,N_17331,N_17624);
or U18496 (N_18496,N_17682,N_17392);
and U18497 (N_18497,N_17224,N_17590);
or U18498 (N_18498,N_17366,N_17498);
nand U18499 (N_18499,N_17572,N_17002);
or U18500 (N_18500,N_17778,N_17271);
or U18501 (N_18501,N_17205,N_17415);
xor U18502 (N_18502,N_17551,N_17667);
and U18503 (N_18503,N_17554,N_17564);
nand U18504 (N_18504,N_17307,N_17527);
and U18505 (N_18505,N_17078,N_17173);
and U18506 (N_18506,N_17626,N_17322);
or U18507 (N_18507,N_17852,N_17742);
nand U18508 (N_18508,N_17730,N_17894);
or U18509 (N_18509,N_17730,N_17278);
and U18510 (N_18510,N_17825,N_17012);
xnor U18511 (N_18511,N_17250,N_17378);
nand U18512 (N_18512,N_17826,N_17248);
and U18513 (N_18513,N_17556,N_17578);
xnor U18514 (N_18514,N_17442,N_17183);
and U18515 (N_18515,N_17205,N_17292);
or U18516 (N_18516,N_17209,N_17240);
nand U18517 (N_18517,N_17560,N_17698);
or U18518 (N_18518,N_17867,N_17971);
nor U18519 (N_18519,N_17713,N_17112);
or U18520 (N_18520,N_17484,N_17550);
nor U18521 (N_18521,N_17653,N_17858);
and U18522 (N_18522,N_17417,N_17149);
and U18523 (N_18523,N_17303,N_17374);
nand U18524 (N_18524,N_17317,N_17835);
or U18525 (N_18525,N_17940,N_17434);
nor U18526 (N_18526,N_17156,N_17417);
xor U18527 (N_18527,N_17722,N_17065);
nor U18528 (N_18528,N_17527,N_17207);
xnor U18529 (N_18529,N_17944,N_17591);
nor U18530 (N_18530,N_17609,N_17114);
and U18531 (N_18531,N_17898,N_17467);
or U18532 (N_18532,N_17178,N_17885);
xnor U18533 (N_18533,N_17074,N_17940);
and U18534 (N_18534,N_17538,N_17264);
xnor U18535 (N_18535,N_17787,N_17230);
nor U18536 (N_18536,N_17607,N_17110);
nor U18537 (N_18537,N_17845,N_17987);
xor U18538 (N_18538,N_17112,N_17392);
nor U18539 (N_18539,N_17495,N_17731);
nor U18540 (N_18540,N_17007,N_17828);
or U18541 (N_18541,N_17509,N_17590);
or U18542 (N_18542,N_17839,N_17849);
nor U18543 (N_18543,N_17201,N_17455);
nand U18544 (N_18544,N_17031,N_17942);
and U18545 (N_18545,N_17200,N_17276);
nor U18546 (N_18546,N_17420,N_17729);
and U18547 (N_18547,N_17965,N_17800);
xnor U18548 (N_18548,N_17732,N_17764);
xor U18549 (N_18549,N_17208,N_17013);
and U18550 (N_18550,N_17973,N_17235);
nand U18551 (N_18551,N_17877,N_17210);
xnor U18552 (N_18552,N_17207,N_17422);
nor U18553 (N_18553,N_17722,N_17655);
nor U18554 (N_18554,N_17301,N_17126);
or U18555 (N_18555,N_17034,N_17380);
xnor U18556 (N_18556,N_17113,N_17440);
nand U18557 (N_18557,N_17306,N_17969);
or U18558 (N_18558,N_17842,N_17874);
and U18559 (N_18559,N_17069,N_17877);
nor U18560 (N_18560,N_17665,N_17598);
nand U18561 (N_18561,N_17966,N_17843);
nand U18562 (N_18562,N_17915,N_17558);
nand U18563 (N_18563,N_17993,N_17978);
nor U18564 (N_18564,N_17582,N_17701);
xnor U18565 (N_18565,N_17438,N_17139);
or U18566 (N_18566,N_17763,N_17279);
nor U18567 (N_18567,N_17856,N_17942);
and U18568 (N_18568,N_17495,N_17757);
or U18569 (N_18569,N_17919,N_17732);
nand U18570 (N_18570,N_17076,N_17077);
nor U18571 (N_18571,N_17763,N_17467);
or U18572 (N_18572,N_17178,N_17509);
nand U18573 (N_18573,N_17563,N_17190);
nand U18574 (N_18574,N_17654,N_17106);
xor U18575 (N_18575,N_17096,N_17544);
and U18576 (N_18576,N_17607,N_17361);
xor U18577 (N_18577,N_17893,N_17127);
xor U18578 (N_18578,N_17779,N_17453);
nand U18579 (N_18579,N_17329,N_17540);
and U18580 (N_18580,N_17807,N_17755);
or U18581 (N_18581,N_17715,N_17555);
xor U18582 (N_18582,N_17803,N_17781);
nand U18583 (N_18583,N_17297,N_17478);
or U18584 (N_18584,N_17905,N_17153);
and U18585 (N_18585,N_17421,N_17352);
or U18586 (N_18586,N_17424,N_17722);
nand U18587 (N_18587,N_17372,N_17354);
nand U18588 (N_18588,N_17060,N_17307);
xnor U18589 (N_18589,N_17382,N_17022);
or U18590 (N_18590,N_17109,N_17775);
nand U18591 (N_18591,N_17841,N_17897);
and U18592 (N_18592,N_17977,N_17019);
nand U18593 (N_18593,N_17923,N_17763);
nand U18594 (N_18594,N_17798,N_17386);
xnor U18595 (N_18595,N_17768,N_17688);
and U18596 (N_18596,N_17875,N_17732);
nor U18597 (N_18597,N_17095,N_17616);
nor U18598 (N_18598,N_17538,N_17914);
nor U18599 (N_18599,N_17951,N_17885);
xor U18600 (N_18600,N_17458,N_17823);
and U18601 (N_18601,N_17411,N_17945);
nor U18602 (N_18602,N_17100,N_17214);
and U18603 (N_18603,N_17335,N_17691);
xor U18604 (N_18604,N_17576,N_17618);
nor U18605 (N_18605,N_17467,N_17735);
or U18606 (N_18606,N_17449,N_17804);
and U18607 (N_18607,N_17344,N_17494);
and U18608 (N_18608,N_17545,N_17355);
nor U18609 (N_18609,N_17177,N_17424);
or U18610 (N_18610,N_17738,N_17673);
and U18611 (N_18611,N_17443,N_17105);
and U18612 (N_18612,N_17872,N_17678);
or U18613 (N_18613,N_17863,N_17346);
nor U18614 (N_18614,N_17566,N_17125);
xnor U18615 (N_18615,N_17443,N_17972);
xnor U18616 (N_18616,N_17652,N_17861);
nand U18617 (N_18617,N_17792,N_17455);
and U18618 (N_18618,N_17257,N_17563);
xnor U18619 (N_18619,N_17622,N_17851);
nand U18620 (N_18620,N_17274,N_17334);
and U18621 (N_18621,N_17228,N_17742);
or U18622 (N_18622,N_17494,N_17591);
and U18623 (N_18623,N_17542,N_17085);
and U18624 (N_18624,N_17984,N_17486);
xnor U18625 (N_18625,N_17602,N_17370);
and U18626 (N_18626,N_17814,N_17834);
nor U18627 (N_18627,N_17040,N_17018);
nand U18628 (N_18628,N_17875,N_17231);
and U18629 (N_18629,N_17391,N_17502);
nor U18630 (N_18630,N_17210,N_17351);
or U18631 (N_18631,N_17230,N_17217);
or U18632 (N_18632,N_17309,N_17557);
nor U18633 (N_18633,N_17375,N_17103);
and U18634 (N_18634,N_17100,N_17032);
nand U18635 (N_18635,N_17228,N_17190);
xor U18636 (N_18636,N_17418,N_17216);
nor U18637 (N_18637,N_17475,N_17095);
or U18638 (N_18638,N_17478,N_17264);
nor U18639 (N_18639,N_17793,N_17134);
xnor U18640 (N_18640,N_17951,N_17314);
nand U18641 (N_18641,N_17555,N_17343);
xor U18642 (N_18642,N_17478,N_17743);
xor U18643 (N_18643,N_17025,N_17431);
and U18644 (N_18644,N_17203,N_17727);
nand U18645 (N_18645,N_17595,N_17313);
or U18646 (N_18646,N_17137,N_17507);
or U18647 (N_18647,N_17432,N_17388);
and U18648 (N_18648,N_17206,N_17268);
or U18649 (N_18649,N_17291,N_17056);
xor U18650 (N_18650,N_17177,N_17198);
or U18651 (N_18651,N_17928,N_17193);
xnor U18652 (N_18652,N_17247,N_17544);
or U18653 (N_18653,N_17631,N_17016);
and U18654 (N_18654,N_17936,N_17882);
or U18655 (N_18655,N_17359,N_17375);
xnor U18656 (N_18656,N_17428,N_17340);
nor U18657 (N_18657,N_17256,N_17073);
nor U18658 (N_18658,N_17668,N_17009);
nor U18659 (N_18659,N_17638,N_17763);
xor U18660 (N_18660,N_17097,N_17384);
xnor U18661 (N_18661,N_17801,N_17046);
nor U18662 (N_18662,N_17283,N_17622);
xnor U18663 (N_18663,N_17743,N_17260);
nor U18664 (N_18664,N_17696,N_17618);
xnor U18665 (N_18665,N_17571,N_17524);
nand U18666 (N_18666,N_17838,N_17006);
or U18667 (N_18667,N_17290,N_17519);
nor U18668 (N_18668,N_17963,N_17186);
or U18669 (N_18669,N_17821,N_17536);
or U18670 (N_18670,N_17378,N_17179);
xnor U18671 (N_18671,N_17940,N_17859);
and U18672 (N_18672,N_17710,N_17366);
and U18673 (N_18673,N_17614,N_17473);
xor U18674 (N_18674,N_17248,N_17009);
nand U18675 (N_18675,N_17657,N_17641);
nor U18676 (N_18676,N_17629,N_17780);
or U18677 (N_18677,N_17929,N_17382);
or U18678 (N_18678,N_17934,N_17831);
nor U18679 (N_18679,N_17571,N_17395);
or U18680 (N_18680,N_17632,N_17760);
nand U18681 (N_18681,N_17641,N_17114);
nand U18682 (N_18682,N_17264,N_17258);
and U18683 (N_18683,N_17080,N_17135);
xnor U18684 (N_18684,N_17263,N_17949);
and U18685 (N_18685,N_17993,N_17078);
nor U18686 (N_18686,N_17712,N_17729);
or U18687 (N_18687,N_17470,N_17694);
nor U18688 (N_18688,N_17995,N_17537);
xor U18689 (N_18689,N_17990,N_17600);
nand U18690 (N_18690,N_17032,N_17041);
nand U18691 (N_18691,N_17184,N_17640);
and U18692 (N_18692,N_17114,N_17044);
xnor U18693 (N_18693,N_17306,N_17931);
and U18694 (N_18694,N_17053,N_17120);
xnor U18695 (N_18695,N_17776,N_17497);
or U18696 (N_18696,N_17588,N_17745);
or U18697 (N_18697,N_17783,N_17361);
xnor U18698 (N_18698,N_17154,N_17101);
xnor U18699 (N_18699,N_17994,N_17486);
nor U18700 (N_18700,N_17383,N_17860);
or U18701 (N_18701,N_17225,N_17432);
nand U18702 (N_18702,N_17957,N_17632);
and U18703 (N_18703,N_17722,N_17355);
or U18704 (N_18704,N_17996,N_17583);
xor U18705 (N_18705,N_17626,N_17603);
nand U18706 (N_18706,N_17111,N_17638);
nand U18707 (N_18707,N_17327,N_17420);
or U18708 (N_18708,N_17060,N_17682);
nor U18709 (N_18709,N_17969,N_17778);
nor U18710 (N_18710,N_17145,N_17909);
or U18711 (N_18711,N_17396,N_17985);
nand U18712 (N_18712,N_17997,N_17617);
xor U18713 (N_18713,N_17597,N_17395);
xnor U18714 (N_18714,N_17608,N_17938);
nand U18715 (N_18715,N_17376,N_17334);
and U18716 (N_18716,N_17445,N_17503);
or U18717 (N_18717,N_17469,N_17898);
nand U18718 (N_18718,N_17832,N_17661);
xnor U18719 (N_18719,N_17371,N_17443);
nand U18720 (N_18720,N_17609,N_17331);
and U18721 (N_18721,N_17228,N_17863);
or U18722 (N_18722,N_17608,N_17086);
nor U18723 (N_18723,N_17973,N_17563);
nor U18724 (N_18724,N_17700,N_17359);
or U18725 (N_18725,N_17363,N_17494);
nor U18726 (N_18726,N_17485,N_17575);
nand U18727 (N_18727,N_17024,N_17188);
and U18728 (N_18728,N_17265,N_17484);
or U18729 (N_18729,N_17985,N_17246);
nor U18730 (N_18730,N_17911,N_17276);
nor U18731 (N_18731,N_17808,N_17534);
and U18732 (N_18732,N_17856,N_17345);
nand U18733 (N_18733,N_17236,N_17520);
nor U18734 (N_18734,N_17764,N_17577);
xnor U18735 (N_18735,N_17999,N_17842);
nor U18736 (N_18736,N_17713,N_17438);
nand U18737 (N_18737,N_17529,N_17109);
xor U18738 (N_18738,N_17716,N_17891);
and U18739 (N_18739,N_17835,N_17657);
nand U18740 (N_18740,N_17249,N_17652);
and U18741 (N_18741,N_17412,N_17934);
nand U18742 (N_18742,N_17122,N_17464);
xor U18743 (N_18743,N_17731,N_17146);
or U18744 (N_18744,N_17266,N_17738);
nor U18745 (N_18745,N_17071,N_17349);
nor U18746 (N_18746,N_17883,N_17983);
nor U18747 (N_18747,N_17793,N_17391);
and U18748 (N_18748,N_17719,N_17018);
xnor U18749 (N_18749,N_17310,N_17816);
nand U18750 (N_18750,N_17860,N_17872);
xor U18751 (N_18751,N_17026,N_17232);
nand U18752 (N_18752,N_17151,N_17943);
xnor U18753 (N_18753,N_17485,N_17526);
or U18754 (N_18754,N_17471,N_17489);
or U18755 (N_18755,N_17656,N_17401);
and U18756 (N_18756,N_17310,N_17642);
and U18757 (N_18757,N_17462,N_17639);
or U18758 (N_18758,N_17238,N_17124);
nand U18759 (N_18759,N_17350,N_17145);
and U18760 (N_18760,N_17329,N_17222);
or U18761 (N_18761,N_17583,N_17541);
nor U18762 (N_18762,N_17696,N_17085);
or U18763 (N_18763,N_17165,N_17846);
nor U18764 (N_18764,N_17264,N_17923);
nor U18765 (N_18765,N_17589,N_17285);
and U18766 (N_18766,N_17593,N_17117);
and U18767 (N_18767,N_17123,N_17692);
and U18768 (N_18768,N_17096,N_17713);
and U18769 (N_18769,N_17741,N_17855);
nor U18770 (N_18770,N_17241,N_17106);
xnor U18771 (N_18771,N_17134,N_17062);
and U18772 (N_18772,N_17718,N_17364);
nand U18773 (N_18773,N_17617,N_17055);
or U18774 (N_18774,N_17340,N_17077);
nor U18775 (N_18775,N_17681,N_17122);
xor U18776 (N_18776,N_17299,N_17355);
xnor U18777 (N_18777,N_17402,N_17138);
or U18778 (N_18778,N_17886,N_17495);
and U18779 (N_18779,N_17772,N_17868);
xor U18780 (N_18780,N_17665,N_17267);
or U18781 (N_18781,N_17303,N_17660);
xor U18782 (N_18782,N_17132,N_17855);
or U18783 (N_18783,N_17453,N_17192);
nand U18784 (N_18784,N_17972,N_17057);
nor U18785 (N_18785,N_17442,N_17556);
xnor U18786 (N_18786,N_17833,N_17092);
and U18787 (N_18787,N_17715,N_17020);
nor U18788 (N_18788,N_17099,N_17385);
or U18789 (N_18789,N_17835,N_17490);
and U18790 (N_18790,N_17102,N_17400);
or U18791 (N_18791,N_17738,N_17764);
xor U18792 (N_18792,N_17064,N_17076);
and U18793 (N_18793,N_17245,N_17903);
and U18794 (N_18794,N_17137,N_17874);
xor U18795 (N_18795,N_17523,N_17079);
and U18796 (N_18796,N_17692,N_17655);
and U18797 (N_18797,N_17223,N_17637);
nand U18798 (N_18798,N_17906,N_17099);
and U18799 (N_18799,N_17116,N_17467);
nand U18800 (N_18800,N_17395,N_17802);
and U18801 (N_18801,N_17167,N_17641);
xor U18802 (N_18802,N_17773,N_17478);
or U18803 (N_18803,N_17686,N_17204);
and U18804 (N_18804,N_17382,N_17524);
nor U18805 (N_18805,N_17730,N_17936);
or U18806 (N_18806,N_17315,N_17088);
nor U18807 (N_18807,N_17996,N_17948);
xnor U18808 (N_18808,N_17533,N_17069);
nand U18809 (N_18809,N_17481,N_17228);
and U18810 (N_18810,N_17512,N_17449);
or U18811 (N_18811,N_17034,N_17961);
xor U18812 (N_18812,N_17634,N_17489);
nor U18813 (N_18813,N_17666,N_17558);
nor U18814 (N_18814,N_17762,N_17163);
nand U18815 (N_18815,N_17127,N_17705);
or U18816 (N_18816,N_17670,N_17335);
xnor U18817 (N_18817,N_17601,N_17166);
xor U18818 (N_18818,N_17916,N_17855);
nand U18819 (N_18819,N_17047,N_17755);
and U18820 (N_18820,N_17795,N_17647);
or U18821 (N_18821,N_17199,N_17722);
nor U18822 (N_18822,N_17296,N_17911);
xnor U18823 (N_18823,N_17626,N_17726);
nand U18824 (N_18824,N_17744,N_17381);
xnor U18825 (N_18825,N_17640,N_17901);
nor U18826 (N_18826,N_17428,N_17892);
nand U18827 (N_18827,N_17511,N_17988);
xor U18828 (N_18828,N_17459,N_17951);
nor U18829 (N_18829,N_17938,N_17606);
nand U18830 (N_18830,N_17217,N_17829);
nor U18831 (N_18831,N_17294,N_17435);
and U18832 (N_18832,N_17714,N_17650);
nor U18833 (N_18833,N_17085,N_17504);
and U18834 (N_18834,N_17420,N_17581);
xnor U18835 (N_18835,N_17045,N_17661);
and U18836 (N_18836,N_17541,N_17348);
nand U18837 (N_18837,N_17423,N_17620);
and U18838 (N_18838,N_17170,N_17735);
xnor U18839 (N_18839,N_17119,N_17399);
nor U18840 (N_18840,N_17129,N_17985);
or U18841 (N_18841,N_17451,N_17053);
nor U18842 (N_18842,N_17965,N_17797);
or U18843 (N_18843,N_17660,N_17129);
or U18844 (N_18844,N_17194,N_17244);
or U18845 (N_18845,N_17137,N_17277);
xor U18846 (N_18846,N_17088,N_17893);
xnor U18847 (N_18847,N_17181,N_17527);
nor U18848 (N_18848,N_17897,N_17450);
nand U18849 (N_18849,N_17417,N_17533);
nor U18850 (N_18850,N_17718,N_17639);
nor U18851 (N_18851,N_17569,N_17510);
and U18852 (N_18852,N_17485,N_17696);
nor U18853 (N_18853,N_17652,N_17865);
or U18854 (N_18854,N_17975,N_17128);
xnor U18855 (N_18855,N_17829,N_17399);
or U18856 (N_18856,N_17064,N_17854);
nand U18857 (N_18857,N_17415,N_17457);
nand U18858 (N_18858,N_17165,N_17603);
or U18859 (N_18859,N_17618,N_17155);
and U18860 (N_18860,N_17629,N_17805);
xor U18861 (N_18861,N_17375,N_17755);
xnor U18862 (N_18862,N_17248,N_17181);
nand U18863 (N_18863,N_17346,N_17950);
nand U18864 (N_18864,N_17567,N_17113);
and U18865 (N_18865,N_17882,N_17359);
xnor U18866 (N_18866,N_17719,N_17910);
or U18867 (N_18867,N_17471,N_17630);
nand U18868 (N_18868,N_17311,N_17269);
nand U18869 (N_18869,N_17875,N_17726);
nand U18870 (N_18870,N_17171,N_17989);
and U18871 (N_18871,N_17157,N_17302);
or U18872 (N_18872,N_17017,N_17654);
nand U18873 (N_18873,N_17543,N_17770);
nor U18874 (N_18874,N_17054,N_17553);
nor U18875 (N_18875,N_17920,N_17990);
xnor U18876 (N_18876,N_17408,N_17547);
and U18877 (N_18877,N_17941,N_17973);
nor U18878 (N_18878,N_17951,N_17844);
nor U18879 (N_18879,N_17889,N_17362);
or U18880 (N_18880,N_17679,N_17971);
or U18881 (N_18881,N_17117,N_17790);
xnor U18882 (N_18882,N_17864,N_17296);
nor U18883 (N_18883,N_17583,N_17736);
nand U18884 (N_18884,N_17228,N_17772);
and U18885 (N_18885,N_17109,N_17812);
xor U18886 (N_18886,N_17100,N_17848);
xnor U18887 (N_18887,N_17414,N_17128);
and U18888 (N_18888,N_17743,N_17143);
xnor U18889 (N_18889,N_17700,N_17502);
xor U18890 (N_18890,N_17613,N_17674);
xnor U18891 (N_18891,N_17437,N_17500);
xnor U18892 (N_18892,N_17386,N_17611);
nor U18893 (N_18893,N_17103,N_17826);
nor U18894 (N_18894,N_17526,N_17502);
and U18895 (N_18895,N_17283,N_17691);
nand U18896 (N_18896,N_17704,N_17936);
nand U18897 (N_18897,N_17895,N_17279);
or U18898 (N_18898,N_17854,N_17034);
nor U18899 (N_18899,N_17085,N_17525);
nand U18900 (N_18900,N_17288,N_17815);
nand U18901 (N_18901,N_17546,N_17475);
nand U18902 (N_18902,N_17737,N_17188);
nand U18903 (N_18903,N_17915,N_17354);
xor U18904 (N_18904,N_17792,N_17305);
and U18905 (N_18905,N_17068,N_17037);
nor U18906 (N_18906,N_17111,N_17757);
nand U18907 (N_18907,N_17901,N_17074);
nor U18908 (N_18908,N_17259,N_17162);
or U18909 (N_18909,N_17906,N_17108);
nor U18910 (N_18910,N_17374,N_17171);
nor U18911 (N_18911,N_17908,N_17021);
and U18912 (N_18912,N_17046,N_17533);
nor U18913 (N_18913,N_17699,N_17044);
xnor U18914 (N_18914,N_17213,N_17989);
xor U18915 (N_18915,N_17248,N_17956);
xor U18916 (N_18916,N_17385,N_17782);
or U18917 (N_18917,N_17721,N_17284);
and U18918 (N_18918,N_17875,N_17871);
or U18919 (N_18919,N_17961,N_17191);
nor U18920 (N_18920,N_17437,N_17111);
and U18921 (N_18921,N_17409,N_17086);
or U18922 (N_18922,N_17178,N_17935);
and U18923 (N_18923,N_17660,N_17197);
nand U18924 (N_18924,N_17572,N_17510);
and U18925 (N_18925,N_17535,N_17941);
or U18926 (N_18926,N_17221,N_17970);
and U18927 (N_18927,N_17164,N_17717);
and U18928 (N_18928,N_17154,N_17060);
nor U18929 (N_18929,N_17188,N_17816);
nand U18930 (N_18930,N_17835,N_17755);
or U18931 (N_18931,N_17888,N_17016);
nor U18932 (N_18932,N_17779,N_17695);
and U18933 (N_18933,N_17129,N_17568);
or U18934 (N_18934,N_17296,N_17954);
nand U18935 (N_18935,N_17057,N_17134);
or U18936 (N_18936,N_17346,N_17922);
nor U18937 (N_18937,N_17497,N_17793);
nor U18938 (N_18938,N_17073,N_17527);
and U18939 (N_18939,N_17248,N_17454);
nor U18940 (N_18940,N_17231,N_17955);
and U18941 (N_18941,N_17101,N_17931);
or U18942 (N_18942,N_17127,N_17082);
and U18943 (N_18943,N_17989,N_17320);
xnor U18944 (N_18944,N_17481,N_17880);
xor U18945 (N_18945,N_17096,N_17315);
xor U18946 (N_18946,N_17472,N_17365);
nor U18947 (N_18947,N_17234,N_17158);
or U18948 (N_18948,N_17339,N_17050);
and U18949 (N_18949,N_17101,N_17724);
or U18950 (N_18950,N_17506,N_17835);
nand U18951 (N_18951,N_17606,N_17597);
xnor U18952 (N_18952,N_17970,N_17172);
xnor U18953 (N_18953,N_17090,N_17097);
nand U18954 (N_18954,N_17118,N_17473);
and U18955 (N_18955,N_17547,N_17509);
nor U18956 (N_18956,N_17614,N_17515);
nor U18957 (N_18957,N_17595,N_17606);
and U18958 (N_18958,N_17873,N_17500);
nand U18959 (N_18959,N_17508,N_17365);
nand U18960 (N_18960,N_17028,N_17308);
nand U18961 (N_18961,N_17384,N_17778);
nor U18962 (N_18962,N_17768,N_17875);
nand U18963 (N_18963,N_17292,N_17261);
and U18964 (N_18964,N_17601,N_17215);
or U18965 (N_18965,N_17004,N_17211);
xnor U18966 (N_18966,N_17125,N_17893);
and U18967 (N_18967,N_17071,N_17473);
xor U18968 (N_18968,N_17017,N_17262);
xnor U18969 (N_18969,N_17119,N_17934);
nand U18970 (N_18970,N_17870,N_17719);
nand U18971 (N_18971,N_17625,N_17811);
nor U18972 (N_18972,N_17169,N_17282);
or U18973 (N_18973,N_17114,N_17368);
nand U18974 (N_18974,N_17504,N_17311);
nor U18975 (N_18975,N_17917,N_17625);
nor U18976 (N_18976,N_17164,N_17363);
and U18977 (N_18977,N_17548,N_17626);
xnor U18978 (N_18978,N_17306,N_17311);
xor U18979 (N_18979,N_17405,N_17853);
nand U18980 (N_18980,N_17909,N_17395);
nor U18981 (N_18981,N_17805,N_17764);
nor U18982 (N_18982,N_17352,N_17687);
or U18983 (N_18983,N_17994,N_17264);
or U18984 (N_18984,N_17615,N_17787);
xnor U18985 (N_18985,N_17770,N_17862);
or U18986 (N_18986,N_17969,N_17473);
nand U18987 (N_18987,N_17206,N_17132);
and U18988 (N_18988,N_17628,N_17168);
or U18989 (N_18989,N_17332,N_17152);
xor U18990 (N_18990,N_17483,N_17918);
nor U18991 (N_18991,N_17241,N_17939);
xnor U18992 (N_18992,N_17127,N_17421);
nor U18993 (N_18993,N_17983,N_17803);
xnor U18994 (N_18994,N_17826,N_17304);
and U18995 (N_18995,N_17062,N_17470);
nand U18996 (N_18996,N_17776,N_17506);
or U18997 (N_18997,N_17816,N_17368);
nand U18998 (N_18998,N_17040,N_17605);
xnor U18999 (N_18999,N_17851,N_17133);
or U19000 (N_19000,N_18737,N_18025);
or U19001 (N_19001,N_18444,N_18030);
xnor U19002 (N_19002,N_18867,N_18521);
and U19003 (N_19003,N_18513,N_18223);
xnor U19004 (N_19004,N_18325,N_18280);
or U19005 (N_19005,N_18087,N_18984);
and U19006 (N_19006,N_18627,N_18118);
nor U19007 (N_19007,N_18157,N_18717);
xor U19008 (N_19008,N_18968,N_18750);
xor U19009 (N_19009,N_18208,N_18562);
and U19010 (N_19010,N_18662,N_18539);
nor U19011 (N_19011,N_18096,N_18593);
xor U19012 (N_19012,N_18209,N_18905);
or U19013 (N_19013,N_18457,N_18274);
and U19014 (N_19014,N_18155,N_18507);
nand U19015 (N_19015,N_18891,N_18917);
or U19016 (N_19016,N_18665,N_18842);
nor U19017 (N_19017,N_18983,N_18449);
or U19018 (N_19018,N_18699,N_18804);
nor U19019 (N_19019,N_18417,N_18973);
xor U19020 (N_19020,N_18017,N_18319);
or U19021 (N_19021,N_18954,N_18597);
xor U19022 (N_19022,N_18198,N_18471);
or U19023 (N_19023,N_18838,N_18048);
and U19024 (N_19024,N_18998,N_18163);
xnor U19025 (N_19025,N_18143,N_18920);
nor U19026 (N_19026,N_18035,N_18814);
nand U19027 (N_19027,N_18394,N_18367);
nand U19028 (N_19028,N_18359,N_18451);
nor U19029 (N_19029,N_18812,N_18124);
nor U19030 (N_19030,N_18523,N_18081);
and U19031 (N_19031,N_18279,N_18939);
nor U19032 (N_19032,N_18502,N_18055);
and U19033 (N_19033,N_18633,N_18706);
and U19034 (N_19034,N_18805,N_18037);
or U19035 (N_19035,N_18335,N_18254);
or U19036 (N_19036,N_18963,N_18635);
nand U19037 (N_19037,N_18168,N_18514);
nand U19038 (N_19038,N_18231,N_18606);
and U19039 (N_19039,N_18967,N_18650);
nand U19040 (N_19040,N_18546,N_18388);
nor U19041 (N_19041,N_18216,N_18074);
or U19042 (N_19042,N_18346,N_18385);
nor U19043 (N_19043,N_18815,N_18008);
and U19044 (N_19044,N_18895,N_18248);
xor U19045 (N_19045,N_18915,N_18570);
or U19046 (N_19046,N_18345,N_18578);
or U19047 (N_19047,N_18496,N_18205);
nand U19048 (N_19048,N_18360,N_18357);
nor U19049 (N_19049,N_18136,N_18363);
nand U19050 (N_19050,N_18387,N_18640);
nor U19051 (N_19051,N_18361,N_18820);
or U19052 (N_19052,N_18364,N_18906);
and U19053 (N_19053,N_18787,N_18158);
xor U19054 (N_19054,N_18889,N_18467);
or U19055 (N_19055,N_18308,N_18896);
nor U19056 (N_19056,N_18041,N_18641);
nor U19057 (N_19057,N_18951,N_18356);
nand U19058 (N_19058,N_18694,N_18749);
nor U19059 (N_19059,N_18621,N_18425);
xnor U19060 (N_19060,N_18292,N_18722);
and U19061 (N_19061,N_18605,N_18468);
or U19062 (N_19062,N_18721,N_18112);
or U19063 (N_19063,N_18407,N_18275);
nor U19064 (N_19064,N_18484,N_18372);
xnor U19065 (N_19065,N_18330,N_18454);
or U19066 (N_19066,N_18421,N_18224);
nor U19067 (N_19067,N_18202,N_18904);
nor U19068 (N_19068,N_18663,N_18064);
nor U19069 (N_19069,N_18545,N_18569);
or U19070 (N_19070,N_18376,N_18877);
or U19071 (N_19071,N_18918,N_18061);
nand U19072 (N_19072,N_18977,N_18647);
and U19073 (N_19073,N_18201,N_18206);
nand U19074 (N_19074,N_18255,N_18504);
nand U19075 (N_19075,N_18540,N_18594);
nor U19076 (N_19076,N_18549,N_18427);
xnor U19077 (N_19077,N_18798,N_18384);
nand U19078 (N_19078,N_18612,N_18241);
nor U19079 (N_19079,N_18347,N_18971);
or U19080 (N_19080,N_18887,N_18765);
nor U19081 (N_19081,N_18868,N_18464);
or U19082 (N_19082,N_18063,N_18192);
nor U19083 (N_19083,N_18290,N_18487);
and U19084 (N_19084,N_18581,N_18693);
and U19085 (N_19085,N_18799,N_18172);
xor U19086 (N_19086,N_18709,N_18398);
xnor U19087 (N_19087,N_18769,N_18832);
and U19088 (N_19088,N_18354,N_18092);
and U19089 (N_19089,N_18324,N_18207);
nand U19090 (N_19090,N_18826,N_18393);
xnor U19091 (N_19091,N_18448,N_18924);
xnor U19092 (N_19092,N_18953,N_18754);
nand U19093 (N_19093,N_18072,N_18733);
or U19094 (N_19094,N_18710,N_18433);
or U19095 (N_19095,N_18472,N_18459);
xnor U19096 (N_19096,N_18463,N_18078);
nor U19097 (N_19097,N_18674,N_18878);
nand U19098 (N_19098,N_18861,N_18145);
xor U19099 (N_19099,N_18188,N_18609);
xor U19100 (N_19100,N_18047,N_18858);
and U19101 (N_19101,N_18311,N_18135);
xor U19102 (N_19102,N_18727,N_18130);
or U19103 (N_19103,N_18149,N_18378);
or U19104 (N_19104,N_18256,N_18550);
or U19105 (N_19105,N_18723,N_18556);
xor U19106 (N_19106,N_18701,N_18196);
nor U19107 (N_19107,N_18980,N_18034);
nand U19108 (N_19108,N_18681,N_18309);
nand U19109 (N_19109,N_18894,N_18755);
or U19110 (N_19110,N_18529,N_18450);
and U19111 (N_19111,N_18422,N_18997);
nand U19112 (N_19112,N_18054,N_18420);
xnor U19113 (N_19113,N_18245,N_18966);
or U19114 (N_19114,N_18310,N_18560);
xor U19115 (N_19115,N_18910,N_18689);
or U19116 (N_19116,N_18132,N_18083);
or U19117 (N_19117,N_18718,N_18528);
nor U19118 (N_19118,N_18007,N_18775);
nand U19119 (N_19119,N_18673,N_18100);
nand U19120 (N_19120,N_18455,N_18713);
or U19121 (N_19121,N_18483,N_18584);
xor U19122 (N_19122,N_18297,N_18212);
nor U19123 (N_19123,N_18724,N_18270);
nor U19124 (N_19124,N_18850,N_18120);
nand U19125 (N_19125,N_18098,N_18604);
xor U19126 (N_19126,N_18505,N_18993);
nand U19127 (N_19127,N_18141,N_18613);
or U19128 (N_19128,N_18999,N_18883);
and U19129 (N_19129,N_18642,N_18180);
nor U19130 (N_19130,N_18049,N_18783);
xor U19131 (N_19131,N_18258,N_18461);
nand U19132 (N_19132,N_18511,N_18497);
xor U19133 (N_19133,N_18946,N_18801);
or U19134 (N_19134,N_18222,N_18732);
nand U19135 (N_19135,N_18106,N_18000);
and U19136 (N_19136,N_18848,N_18147);
and U19137 (N_19137,N_18866,N_18720);
nor U19138 (N_19138,N_18111,N_18683);
or U19139 (N_19139,N_18538,N_18987);
or U19140 (N_19140,N_18544,N_18304);
and U19141 (N_19141,N_18473,N_18389);
nand U19142 (N_19142,N_18036,N_18655);
nor U19143 (N_19143,N_18568,N_18856);
and U19144 (N_19144,N_18059,N_18476);
or U19145 (N_19145,N_18142,N_18789);
nor U19146 (N_19146,N_18014,N_18757);
nor U19147 (N_19147,N_18115,N_18088);
and U19148 (N_19148,N_18090,N_18257);
or U19149 (N_19149,N_18844,N_18328);
or U19150 (N_19150,N_18179,N_18992);
xnor U19151 (N_19151,N_18341,N_18520);
xnor U19152 (N_19152,N_18611,N_18171);
nand U19153 (N_19153,N_18602,N_18159);
or U19154 (N_19154,N_18784,N_18708);
nand U19155 (N_19155,N_18742,N_18499);
nand U19156 (N_19156,N_18622,N_18873);
xor U19157 (N_19157,N_18637,N_18936);
nand U19158 (N_19158,N_18161,N_18730);
xnor U19159 (N_19159,N_18091,N_18340);
xor U19160 (N_19160,N_18151,N_18751);
or U19161 (N_19161,N_18071,N_18728);
or U19162 (N_19162,N_18726,N_18006);
xnor U19163 (N_19163,N_18320,N_18571);
or U19164 (N_19164,N_18766,N_18339);
xor U19165 (N_19165,N_18630,N_18351);
xnor U19166 (N_19166,N_18288,N_18739);
nand U19167 (N_19167,N_18933,N_18767);
nor U19168 (N_19168,N_18313,N_18373);
and U19169 (N_19169,N_18186,N_18278);
nor U19170 (N_19170,N_18758,N_18862);
and U19171 (N_19171,N_18436,N_18958);
or U19172 (N_19172,N_18266,N_18317);
nand U19173 (N_19173,N_18780,N_18084);
or U19174 (N_19174,N_18534,N_18849);
nand U19175 (N_19175,N_18428,N_18975);
nand U19176 (N_19176,N_18104,N_18553);
nor U19177 (N_19177,N_18949,N_18580);
or U19178 (N_19178,N_18032,N_18247);
nand U19179 (N_19179,N_18276,N_18827);
and U19180 (N_19180,N_18770,N_18094);
nand U19181 (N_19181,N_18563,N_18719);
nand U19182 (N_19182,N_18919,N_18458);
and U19183 (N_19183,N_18964,N_18771);
and U19184 (N_19184,N_18267,N_18167);
and U19185 (N_19185,N_18183,N_18348);
nand U19186 (N_19186,N_18574,N_18854);
nor U19187 (N_19187,N_18934,N_18555);
nand U19188 (N_19188,N_18625,N_18995);
xor U19189 (N_19189,N_18986,N_18551);
and U19190 (N_19190,N_18139,N_18156);
or U19191 (N_19191,N_18038,N_18460);
xor U19192 (N_19192,N_18108,N_18860);
or U19193 (N_19193,N_18703,N_18774);
and U19194 (N_19194,N_18970,N_18636);
nor U19195 (N_19195,N_18644,N_18857);
nand U19196 (N_19196,N_18927,N_18039);
nor U19197 (N_19197,N_18137,N_18794);
xor U19198 (N_19198,N_18478,N_18731);
nand U19199 (N_19199,N_18073,N_18768);
nor U19200 (N_19200,N_18576,N_18316);
xor U19201 (N_19201,N_18044,N_18495);
xnor U19202 (N_19202,N_18148,N_18109);
and U19203 (N_19203,N_18876,N_18107);
xnor U19204 (N_19204,N_18489,N_18237);
nor U19205 (N_19205,N_18716,N_18649);
xor U19206 (N_19206,N_18023,N_18806);
or U19207 (N_19207,N_18045,N_18535);
or U19208 (N_19208,N_18065,N_18852);
or U19209 (N_19209,N_18518,N_18312);
xnor U19210 (N_19210,N_18485,N_18482);
nand U19211 (N_19211,N_18438,N_18705);
nand U19212 (N_19212,N_18976,N_18952);
or U19213 (N_19213,N_18575,N_18589);
xor U19214 (N_19214,N_18164,N_18371);
nor U19215 (N_19215,N_18283,N_18872);
and U19216 (N_19216,N_18401,N_18542);
nor U19217 (N_19217,N_18413,N_18796);
xnor U19218 (N_19218,N_18567,N_18989);
or U19219 (N_19219,N_18479,N_18797);
xnor U19220 (N_19220,N_18711,N_18572);
or U19221 (N_19221,N_18672,N_18800);
and U19222 (N_19222,N_18114,N_18639);
nor U19223 (N_19223,N_18591,N_18005);
xor U19224 (N_19224,N_18537,N_18380);
xnor U19225 (N_19225,N_18122,N_18391);
or U19226 (N_19226,N_18121,N_18592);
nand U19227 (N_19227,N_18969,N_18629);
nor U19228 (N_19228,N_18125,N_18903);
xor U19229 (N_19229,N_18807,N_18229);
nand U19230 (N_19230,N_18408,N_18029);
or U19231 (N_19231,N_18818,N_18300);
xor U19232 (N_19232,N_18493,N_18058);
nand U19233 (N_19233,N_18410,N_18645);
xnor U19234 (N_19234,N_18260,N_18790);
nor U19235 (N_19235,N_18874,N_18654);
or U19236 (N_19236,N_18264,N_18431);
and U19237 (N_19237,N_18618,N_18880);
nor U19238 (N_19238,N_18524,N_18439);
nand U19239 (N_19239,N_18187,N_18522);
and U19240 (N_19240,N_18286,N_18337);
or U19241 (N_19241,N_18203,N_18375);
nor U19242 (N_19242,N_18195,N_18501);
and U19243 (N_19243,N_18741,N_18344);
nand U19244 (N_19244,N_18558,N_18836);
xnor U19245 (N_19245,N_18955,N_18598);
nor U19246 (N_19246,N_18272,N_18412);
xor U19247 (N_19247,N_18819,N_18166);
and U19248 (N_19248,N_18123,N_18441);
or U19249 (N_19249,N_18102,N_18462);
xor U19250 (N_19250,N_18268,N_18326);
xnor U19251 (N_19251,N_18947,N_18001);
xor U19252 (N_19252,N_18698,N_18066);
nand U19253 (N_19253,N_18785,N_18046);
and U19254 (N_19254,N_18273,N_18128);
xnor U19255 (N_19255,N_18217,N_18251);
or U19256 (N_19256,N_18885,N_18442);
or U19257 (N_19257,N_18777,N_18808);
nor U19258 (N_19258,N_18822,N_18028);
nor U19259 (N_19259,N_18839,N_18051);
nand U19260 (N_19260,N_18079,N_18515);
nor U19261 (N_19261,N_18342,N_18194);
or U19262 (N_19262,N_18343,N_18435);
and U19263 (N_19263,N_18480,N_18956);
xnor U19264 (N_19264,N_18525,N_18855);
and U19265 (N_19265,N_18369,N_18676);
and U19266 (N_19266,N_18786,N_18791);
nand U19267 (N_19267,N_18670,N_18227);
or U19268 (N_19268,N_18093,N_18652);
nand U19269 (N_19269,N_18409,N_18923);
nand U19270 (N_19270,N_18871,N_18230);
or U19271 (N_19271,N_18293,N_18817);
xor U19272 (N_19272,N_18738,N_18491);
or U19273 (N_19273,N_18846,N_18825);
nor U19274 (N_19274,N_18829,N_18859);
nor U19275 (N_19275,N_18982,N_18447);
xor U19276 (N_19276,N_18557,N_18657);
or U19277 (N_19277,N_18469,N_18697);
and U19278 (N_19278,N_18162,N_18599);
xnor U19279 (N_19279,N_18010,N_18383);
and U19280 (N_19280,N_18884,N_18146);
xor U19281 (N_19281,N_18931,N_18870);
and U19282 (N_19282,N_18759,N_18620);
xor U19283 (N_19283,N_18185,N_18374);
or U19284 (N_19284,N_18013,N_18475);
nand U19285 (N_19285,N_18888,N_18176);
nand U19286 (N_19286,N_18299,N_18623);
nand U19287 (N_19287,N_18691,N_18498);
nand U19288 (N_19288,N_18875,N_18150);
nor U19289 (N_19289,N_18590,N_18062);
or U19290 (N_19290,N_18648,N_18748);
or U19291 (N_19291,N_18643,N_18453);
or U19292 (N_19292,N_18508,N_18138);
and U19293 (N_19293,N_18664,N_18811);
nand U19294 (N_19294,N_18991,N_18659);
nor U19295 (N_19295,N_18377,N_18190);
or U19296 (N_19296,N_18532,N_18835);
and U19297 (N_19297,N_18076,N_18752);
nand U19298 (N_19298,N_18821,N_18456);
xor U19299 (N_19299,N_18236,N_18680);
xnor U19300 (N_19300,N_18004,N_18285);
nor U19301 (N_19301,N_18828,N_18792);
and U19302 (N_19302,N_18651,N_18234);
xor U19303 (N_19303,N_18119,N_18715);
and U19304 (N_19304,N_18189,N_18333);
or U19305 (N_19305,N_18519,N_18295);
or U19306 (N_19306,N_18490,N_18116);
or U19307 (N_19307,N_18712,N_18960);
nor U19308 (N_19308,N_18153,N_18607);
or U19309 (N_19309,N_18579,N_18834);
or U19310 (N_19310,N_18466,N_18940);
or U19311 (N_19311,N_18200,N_18740);
or U19312 (N_19312,N_18253,N_18847);
or U19313 (N_19313,N_18327,N_18284);
or U19314 (N_19314,N_18583,N_18249);
or U19315 (N_19315,N_18303,N_18154);
nor U19316 (N_19316,N_18152,N_18486);
or U19317 (N_19317,N_18756,N_18117);
xor U19318 (N_19318,N_18926,N_18943);
nor U19319 (N_19319,N_18864,N_18988);
xor U19320 (N_19320,N_18778,N_18215);
xor U19321 (N_19321,N_18204,N_18688);
or U19322 (N_19322,N_18776,N_18133);
xnor U19323 (N_19323,N_18390,N_18305);
nor U19324 (N_19324,N_18684,N_18585);
nand U19325 (N_19325,N_18178,N_18003);
or U19326 (N_19326,N_18900,N_18331);
or U19327 (N_19327,N_18810,N_18281);
xor U19328 (N_19328,N_18907,N_18033);
nor U19329 (N_19329,N_18559,N_18452);
nor U19330 (N_19330,N_18669,N_18404);
xnor U19331 (N_19331,N_18773,N_18411);
nand U19332 (N_19332,N_18322,N_18024);
or U19333 (N_19333,N_18314,N_18400);
and U19334 (N_19334,N_18948,N_18911);
and U19335 (N_19335,N_18845,N_18077);
nand U19336 (N_19336,N_18879,N_18682);
nor U19337 (N_19337,N_18714,N_18517);
nor U19338 (N_19338,N_18886,N_18169);
nand U19339 (N_19339,N_18841,N_18961);
nor U19340 (N_19340,N_18582,N_18243);
or U19341 (N_19341,N_18653,N_18349);
nand U19342 (N_19342,N_18638,N_18586);
and U19343 (N_19343,N_18015,N_18823);
nor U19344 (N_19344,N_18282,N_18220);
nor U19345 (N_19345,N_18831,N_18541);
xnor U19346 (N_19346,N_18429,N_18628);
and U19347 (N_19347,N_18445,N_18210);
nand U19348 (N_19348,N_18397,N_18938);
nor U19349 (N_19349,N_18080,N_18901);
xor U19350 (N_19350,N_18941,N_18307);
xnor U19351 (N_19351,N_18430,N_18177);
nand U19352 (N_19352,N_18067,N_18909);
or U19353 (N_19353,N_18095,N_18082);
or U19354 (N_19354,N_18668,N_18837);
and U19355 (N_19355,N_18226,N_18959);
nor U19356 (N_19356,N_18577,N_18019);
or U19357 (N_19357,N_18702,N_18213);
and U19358 (N_19358,N_18779,N_18990);
or U19359 (N_19359,N_18443,N_18793);
nor U19360 (N_19360,N_18370,N_18908);
and U19361 (N_19361,N_18914,N_18211);
nor U19362 (N_19362,N_18350,N_18677);
xnor U19363 (N_19363,N_18050,N_18962);
or U19364 (N_19364,N_18671,N_18692);
xor U19365 (N_19365,N_18945,N_18890);
nand U19366 (N_19366,N_18631,N_18500);
nor U19367 (N_19367,N_18734,N_18040);
and U19368 (N_19368,N_18561,N_18965);
or U19369 (N_19369,N_18252,N_18761);
nand U19370 (N_19370,N_18503,N_18695);
nor U19371 (N_19371,N_18294,N_18181);
nor U19372 (N_19372,N_18246,N_18352);
xor U19373 (N_19373,N_18173,N_18746);
and U19374 (N_19374,N_18813,N_18830);
and U19375 (N_19375,N_18191,N_18685);
xnor U19376 (N_19376,N_18113,N_18552);
or U19377 (N_19377,N_18530,N_18418);
xor U19378 (N_19378,N_18446,N_18928);
nor U19379 (N_19379,N_18916,N_18735);
nor U19380 (N_19380,N_18396,N_18743);
and U19381 (N_19381,N_18573,N_18020);
and U19382 (N_19382,N_18686,N_18492);
nand U19383 (N_19383,N_18395,N_18564);
nand U19384 (N_19384,N_18996,N_18465);
nor U19385 (N_19385,N_18301,N_18921);
or U19386 (N_19386,N_18022,N_18233);
or U19387 (N_19387,N_18382,N_18239);
nand U19388 (N_19388,N_18182,N_18678);
xor U19389 (N_19389,N_18042,N_18772);
nand U19390 (N_19390,N_18160,N_18736);
and U19391 (N_19391,N_18565,N_18416);
xnor U19392 (N_19392,N_18296,N_18527);
nand U19393 (N_19393,N_18851,N_18932);
nand U19394 (N_19394,N_18103,N_18238);
nor U19395 (N_19395,N_18199,N_18610);
and U19396 (N_19396,N_18099,N_18614);
xnor U19397 (N_19397,N_18944,N_18291);
and U19398 (N_19398,N_18893,N_18235);
xor U19399 (N_19399,N_18057,N_18334);
xnor U19400 (N_19400,N_18543,N_18781);
and U19401 (N_19401,N_18240,N_18744);
and U19402 (N_19402,N_18603,N_18596);
nand U19403 (N_19403,N_18250,N_18379);
xor U19404 (N_19404,N_18753,N_18287);
nor U19405 (N_19405,N_18690,N_18009);
xnor U19406 (N_19406,N_18930,N_18175);
nand U19407 (N_19407,N_18228,N_18402);
nor U19408 (N_19408,N_18075,N_18437);
xnor U19409 (N_19409,N_18336,N_18060);
nand U19410 (N_19410,N_18666,N_18824);
nand U19411 (N_19411,N_18170,N_18184);
nor U19412 (N_19412,N_18424,N_18863);
xor U19413 (N_19413,N_18600,N_18085);
or U19414 (N_19414,N_18318,N_18419);
xor U19415 (N_19415,N_18833,N_18386);
nand U19416 (N_19416,N_18031,N_18488);
nor U19417 (N_19417,N_18432,N_18261);
nand U19418 (N_19418,N_18126,N_18018);
and U19419 (N_19419,N_18533,N_18302);
or U19420 (N_19420,N_18011,N_18667);
and U19421 (N_19421,N_18548,N_18747);
and U19422 (N_19422,N_18913,N_18840);
or U19423 (N_19423,N_18426,N_18110);
nand U19424 (N_19424,N_18381,N_18366);
and U19425 (N_19425,N_18788,N_18809);
nand U19426 (N_19426,N_18510,N_18957);
nand U19427 (N_19427,N_18089,N_18972);
or U19428 (N_19428,N_18803,N_18922);
nand U19429 (N_19429,N_18415,N_18547);
or U19430 (N_19430,N_18144,N_18134);
nand U19431 (N_19431,N_18843,N_18218);
xnor U19432 (N_19432,N_18232,N_18892);
nand U19433 (N_19433,N_18332,N_18225);
and U19434 (N_19434,N_18405,N_18289);
and U19435 (N_19435,N_18277,N_18974);
nand U19436 (N_19436,N_18271,N_18338);
nand U19437 (N_19437,N_18942,N_18595);
nand U19438 (N_19438,N_18242,N_18763);
nand U19439 (N_19439,N_18929,N_18566);
nand U19440 (N_19440,N_18687,N_18616);
or U19441 (N_19441,N_18069,N_18365);
nand U19442 (N_19442,N_18588,N_18129);
or U19443 (N_19443,N_18329,N_18392);
xor U19444 (N_19444,N_18626,N_18795);
and U19445 (N_19445,N_18259,N_18764);
xor U19446 (N_19446,N_18601,N_18745);
nand U19447 (N_19447,N_18937,N_18704);
nand U19448 (N_19448,N_18012,N_18898);
and U19449 (N_19449,N_18679,N_18086);
or U19450 (N_19450,N_18105,N_18950);
nor U19451 (N_19451,N_18002,N_18646);
nor U19452 (N_19452,N_18882,N_18509);
and U19453 (N_19453,N_18912,N_18516);
and U19454 (N_19454,N_18244,N_18262);
and U19455 (N_19455,N_18725,N_18782);
or U19456 (N_19456,N_18131,N_18634);
nand U19457 (N_19457,N_18174,N_18615);
or U19458 (N_19458,N_18403,N_18315);
nand U19459 (N_19459,N_18994,N_18608);
nor U19460 (N_19460,N_18869,N_18802);
nor U19461 (N_19461,N_18263,N_18700);
nor U19462 (N_19462,N_18554,N_18127);
nand U19463 (N_19463,N_18656,N_18056);
nor U19464 (N_19464,N_18865,N_18052);
or U19465 (N_19465,N_18140,N_18531);
nand U19466 (N_19466,N_18221,N_18043);
nor U19467 (N_19467,N_18368,N_18399);
nand U19468 (N_19468,N_18978,N_18306);
nand U19469 (N_19469,N_18026,N_18658);
or U19470 (N_19470,N_18925,N_18440);
or U19471 (N_19471,N_18477,N_18298);
nor U19472 (N_19472,N_18406,N_18536);
or U19473 (N_19473,N_18021,N_18587);
xnor U19474 (N_19474,N_18816,N_18512);
or U19475 (N_19475,N_18617,N_18101);
nor U19476 (N_19476,N_18899,N_18269);
nor U19477 (N_19477,N_18853,N_18624);
or U19478 (N_19478,N_18632,N_18353);
xnor U19479 (N_19479,N_18214,N_18661);
xor U19480 (N_19480,N_18619,N_18760);
and U19481 (N_19481,N_18165,N_18414);
or U19482 (N_19482,N_18707,N_18902);
nand U19483 (N_19483,N_18762,N_18729);
nor U19484 (N_19484,N_18494,N_18265);
or U19485 (N_19485,N_18474,N_18675);
nand U19486 (N_19486,N_18506,N_18985);
nor U19487 (N_19487,N_18470,N_18219);
and U19488 (N_19488,N_18423,N_18068);
nor U19489 (N_19489,N_18323,N_18660);
or U19490 (N_19490,N_18016,N_18097);
and U19491 (N_19491,N_18481,N_18979);
nor U19492 (N_19492,N_18897,N_18935);
nor U19493 (N_19493,N_18981,N_18053);
nor U19494 (N_19494,N_18362,N_18027);
and U19495 (N_19495,N_18358,N_18193);
nand U19496 (N_19496,N_18070,N_18355);
nand U19497 (N_19497,N_18321,N_18526);
nor U19498 (N_19498,N_18881,N_18197);
or U19499 (N_19499,N_18696,N_18434);
or U19500 (N_19500,N_18941,N_18743);
nand U19501 (N_19501,N_18537,N_18546);
or U19502 (N_19502,N_18899,N_18578);
nor U19503 (N_19503,N_18058,N_18368);
xnor U19504 (N_19504,N_18053,N_18828);
nor U19505 (N_19505,N_18953,N_18543);
nand U19506 (N_19506,N_18361,N_18765);
or U19507 (N_19507,N_18211,N_18366);
or U19508 (N_19508,N_18731,N_18397);
nand U19509 (N_19509,N_18328,N_18877);
and U19510 (N_19510,N_18849,N_18523);
nor U19511 (N_19511,N_18336,N_18992);
xor U19512 (N_19512,N_18071,N_18058);
nand U19513 (N_19513,N_18466,N_18865);
nand U19514 (N_19514,N_18934,N_18591);
xor U19515 (N_19515,N_18013,N_18693);
nor U19516 (N_19516,N_18020,N_18300);
and U19517 (N_19517,N_18945,N_18703);
and U19518 (N_19518,N_18631,N_18199);
or U19519 (N_19519,N_18027,N_18167);
nor U19520 (N_19520,N_18482,N_18650);
or U19521 (N_19521,N_18316,N_18813);
or U19522 (N_19522,N_18790,N_18177);
xor U19523 (N_19523,N_18336,N_18897);
and U19524 (N_19524,N_18069,N_18673);
and U19525 (N_19525,N_18594,N_18970);
xnor U19526 (N_19526,N_18485,N_18521);
nor U19527 (N_19527,N_18462,N_18292);
nor U19528 (N_19528,N_18385,N_18892);
or U19529 (N_19529,N_18028,N_18269);
nand U19530 (N_19530,N_18960,N_18403);
and U19531 (N_19531,N_18606,N_18647);
and U19532 (N_19532,N_18170,N_18314);
and U19533 (N_19533,N_18384,N_18470);
nand U19534 (N_19534,N_18045,N_18073);
nand U19535 (N_19535,N_18815,N_18689);
or U19536 (N_19536,N_18016,N_18715);
xor U19537 (N_19537,N_18986,N_18123);
and U19538 (N_19538,N_18150,N_18917);
xor U19539 (N_19539,N_18363,N_18642);
or U19540 (N_19540,N_18078,N_18409);
xnor U19541 (N_19541,N_18840,N_18087);
nor U19542 (N_19542,N_18807,N_18248);
xor U19543 (N_19543,N_18634,N_18537);
or U19544 (N_19544,N_18688,N_18399);
xor U19545 (N_19545,N_18385,N_18612);
nand U19546 (N_19546,N_18876,N_18012);
nor U19547 (N_19547,N_18051,N_18318);
xnor U19548 (N_19548,N_18450,N_18470);
and U19549 (N_19549,N_18586,N_18023);
nor U19550 (N_19550,N_18402,N_18129);
nor U19551 (N_19551,N_18094,N_18456);
nor U19552 (N_19552,N_18093,N_18083);
or U19553 (N_19553,N_18537,N_18427);
or U19554 (N_19554,N_18291,N_18279);
and U19555 (N_19555,N_18706,N_18520);
nor U19556 (N_19556,N_18907,N_18460);
xnor U19557 (N_19557,N_18097,N_18317);
nand U19558 (N_19558,N_18309,N_18699);
nor U19559 (N_19559,N_18557,N_18472);
or U19560 (N_19560,N_18674,N_18877);
or U19561 (N_19561,N_18230,N_18804);
nand U19562 (N_19562,N_18099,N_18383);
nand U19563 (N_19563,N_18683,N_18617);
nor U19564 (N_19564,N_18227,N_18195);
nand U19565 (N_19565,N_18531,N_18779);
nor U19566 (N_19566,N_18884,N_18419);
xor U19567 (N_19567,N_18490,N_18924);
xor U19568 (N_19568,N_18383,N_18686);
or U19569 (N_19569,N_18091,N_18110);
or U19570 (N_19570,N_18593,N_18427);
nand U19571 (N_19571,N_18920,N_18084);
nor U19572 (N_19572,N_18851,N_18551);
or U19573 (N_19573,N_18840,N_18269);
nor U19574 (N_19574,N_18937,N_18744);
and U19575 (N_19575,N_18305,N_18734);
or U19576 (N_19576,N_18485,N_18240);
or U19577 (N_19577,N_18813,N_18711);
nand U19578 (N_19578,N_18406,N_18444);
or U19579 (N_19579,N_18835,N_18833);
and U19580 (N_19580,N_18800,N_18913);
xor U19581 (N_19581,N_18871,N_18692);
nand U19582 (N_19582,N_18277,N_18787);
xnor U19583 (N_19583,N_18657,N_18844);
nand U19584 (N_19584,N_18091,N_18781);
nand U19585 (N_19585,N_18803,N_18658);
or U19586 (N_19586,N_18891,N_18483);
nand U19587 (N_19587,N_18439,N_18579);
nor U19588 (N_19588,N_18984,N_18737);
xnor U19589 (N_19589,N_18172,N_18307);
nand U19590 (N_19590,N_18318,N_18513);
or U19591 (N_19591,N_18216,N_18938);
nor U19592 (N_19592,N_18301,N_18961);
xor U19593 (N_19593,N_18028,N_18738);
nand U19594 (N_19594,N_18379,N_18774);
or U19595 (N_19595,N_18600,N_18547);
nor U19596 (N_19596,N_18905,N_18087);
and U19597 (N_19597,N_18878,N_18499);
nor U19598 (N_19598,N_18619,N_18602);
nor U19599 (N_19599,N_18805,N_18262);
xor U19600 (N_19600,N_18955,N_18968);
nand U19601 (N_19601,N_18932,N_18587);
or U19602 (N_19602,N_18093,N_18923);
xor U19603 (N_19603,N_18833,N_18117);
or U19604 (N_19604,N_18556,N_18466);
and U19605 (N_19605,N_18264,N_18242);
nor U19606 (N_19606,N_18881,N_18048);
or U19607 (N_19607,N_18932,N_18143);
and U19608 (N_19608,N_18101,N_18305);
nand U19609 (N_19609,N_18149,N_18831);
xor U19610 (N_19610,N_18615,N_18663);
nor U19611 (N_19611,N_18221,N_18942);
and U19612 (N_19612,N_18860,N_18710);
or U19613 (N_19613,N_18701,N_18418);
and U19614 (N_19614,N_18129,N_18309);
and U19615 (N_19615,N_18241,N_18704);
xor U19616 (N_19616,N_18652,N_18205);
and U19617 (N_19617,N_18906,N_18527);
nor U19618 (N_19618,N_18412,N_18525);
nor U19619 (N_19619,N_18245,N_18970);
or U19620 (N_19620,N_18734,N_18176);
nor U19621 (N_19621,N_18463,N_18960);
nand U19622 (N_19622,N_18388,N_18626);
xor U19623 (N_19623,N_18615,N_18632);
xor U19624 (N_19624,N_18966,N_18314);
xor U19625 (N_19625,N_18121,N_18796);
nor U19626 (N_19626,N_18260,N_18271);
or U19627 (N_19627,N_18338,N_18521);
xnor U19628 (N_19628,N_18483,N_18998);
nor U19629 (N_19629,N_18162,N_18047);
xor U19630 (N_19630,N_18569,N_18696);
or U19631 (N_19631,N_18212,N_18764);
nand U19632 (N_19632,N_18680,N_18111);
nand U19633 (N_19633,N_18113,N_18758);
or U19634 (N_19634,N_18524,N_18593);
nand U19635 (N_19635,N_18321,N_18874);
nand U19636 (N_19636,N_18455,N_18584);
xor U19637 (N_19637,N_18184,N_18808);
or U19638 (N_19638,N_18562,N_18444);
or U19639 (N_19639,N_18772,N_18964);
xnor U19640 (N_19640,N_18800,N_18421);
nor U19641 (N_19641,N_18567,N_18467);
nand U19642 (N_19642,N_18172,N_18860);
and U19643 (N_19643,N_18142,N_18494);
nor U19644 (N_19644,N_18861,N_18162);
and U19645 (N_19645,N_18003,N_18406);
or U19646 (N_19646,N_18274,N_18872);
nor U19647 (N_19647,N_18191,N_18828);
or U19648 (N_19648,N_18445,N_18318);
xor U19649 (N_19649,N_18041,N_18421);
and U19650 (N_19650,N_18611,N_18357);
and U19651 (N_19651,N_18194,N_18663);
nor U19652 (N_19652,N_18881,N_18490);
and U19653 (N_19653,N_18414,N_18489);
or U19654 (N_19654,N_18515,N_18293);
nor U19655 (N_19655,N_18429,N_18309);
or U19656 (N_19656,N_18605,N_18962);
and U19657 (N_19657,N_18606,N_18826);
and U19658 (N_19658,N_18420,N_18992);
or U19659 (N_19659,N_18578,N_18218);
nor U19660 (N_19660,N_18631,N_18028);
or U19661 (N_19661,N_18852,N_18560);
or U19662 (N_19662,N_18412,N_18926);
or U19663 (N_19663,N_18704,N_18543);
and U19664 (N_19664,N_18702,N_18942);
or U19665 (N_19665,N_18633,N_18467);
and U19666 (N_19666,N_18811,N_18401);
nand U19667 (N_19667,N_18380,N_18845);
nand U19668 (N_19668,N_18782,N_18705);
or U19669 (N_19669,N_18894,N_18890);
or U19670 (N_19670,N_18834,N_18388);
nor U19671 (N_19671,N_18658,N_18655);
xnor U19672 (N_19672,N_18287,N_18112);
and U19673 (N_19673,N_18612,N_18131);
nor U19674 (N_19674,N_18872,N_18592);
and U19675 (N_19675,N_18387,N_18862);
and U19676 (N_19676,N_18317,N_18635);
nor U19677 (N_19677,N_18875,N_18179);
and U19678 (N_19678,N_18333,N_18454);
nand U19679 (N_19679,N_18618,N_18557);
or U19680 (N_19680,N_18345,N_18713);
xnor U19681 (N_19681,N_18439,N_18657);
nor U19682 (N_19682,N_18994,N_18781);
and U19683 (N_19683,N_18445,N_18525);
or U19684 (N_19684,N_18944,N_18624);
xnor U19685 (N_19685,N_18008,N_18805);
xnor U19686 (N_19686,N_18240,N_18644);
nand U19687 (N_19687,N_18496,N_18914);
or U19688 (N_19688,N_18714,N_18381);
or U19689 (N_19689,N_18350,N_18965);
and U19690 (N_19690,N_18556,N_18860);
nor U19691 (N_19691,N_18109,N_18482);
or U19692 (N_19692,N_18492,N_18398);
nor U19693 (N_19693,N_18534,N_18039);
and U19694 (N_19694,N_18850,N_18681);
nand U19695 (N_19695,N_18982,N_18440);
xnor U19696 (N_19696,N_18815,N_18867);
and U19697 (N_19697,N_18654,N_18647);
or U19698 (N_19698,N_18656,N_18064);
nor U19699 (N_19699,N_18038,N_18829);
xor U19700 (N_19700,N_18978,N_18239);
xor U19701 (N_19701,N_18746,N_18972);
or U19702 (N_19702,N_18338,N_18335);
and U19703 (N_19703,N_18447,N_18672);
xor U19704 (N_19704,N_18436,N_18981);
and U19705 (N_19705,N_18837,N_18805);
or U19706 (N_19706,N_18458,N_18375);
and U19707 (N_19707,N_18167,N_18063);
or U19708 (N_19708,N_18574,N_18122);
nand U19709 (N_19709,N_18546,N_18676);
or U19710 (N_19710,N_18009,N_18542);
nand U19711 (N_19711,N_18341,N_18919);
xnor U19712 (N_19712,N_18216,N_18743);
nand U19713 (N_19713,N_18575,N_18086);
nand U19714 (N_19714,N_18968,N_18204);
nand U19715 (N_19715,N_18681,N_18297);
or U19716 (N_19716,N_18083,N_18737);
nand U19717 (N_19717,N_18954,N_18773);
or U19718 (N_19718,N_18986,N_18411);
nand U19719 (N_19719,N_18927,N_18090);
nor U19720 (N_19720,N_18847,N_18907);
xnor U19721 (N_19721,N_18476,N_18882);
or U19722 (N_19722,N_18008,N_18063);
nor U19723 (N_19723,N_18090,N_18453);
and U19724 (N_19724,N_18341,N_18349);
or U19725 (N_19725,N_18259,N_18918);
nor U19726 (N_19726,N_18203,N_18322);
nor U19727 (N_19727,N_18579,N_18054);
nand U19728 (N_19728,N_18792,N_18362);
and U19729 (N_19729,N_18245,N_18584);
or U19730 (N_19730,N_18868,N_18951);
xor U19731 (N_19731,N_18091,N_18015);
xnor U19732 (N_19732,N_18840,N_18433);
nor U19733 (N_19733,N_18237,N_18260);
or U19734 (N_19734,N_18819,N_18637);
or U19735 (N_19735,N_18140,N_18925);
or U19736 (N_19736,N_18857,N_18782);
xor U19737 (N_19737,N_18895,N_18785);
or U19738 (N_19738,N_18321,N_18729);
nor U19739 (N_19739,N_18695,N_18888);
or U19740 (N_19740,N_18062,N_18033);
or U19741 (N_19741,N_18950,N_18328);
and U19742 (N_19742,N_18161,N_18147);
or U19743 (N_19743,N_18270,N_18355);
xor U19744 (N_19744,N_18431,N_18094);
nor U19745 (N_19745,N_18689,N_18181);
nor U19746 (N_19746,N_18757,N_18800);
xor U19747 (N_19747,N_18744,N_18016);
or U19748 (N_19748,N_18342,N_18277);
nor U19749 (N_19749,N_18324,N_18960);
nand U19750 (N_19750,N_18060,N_18670);
nand U19751 (N_19751,N_18933,N_18502);
nor U19752 (N_19752,N_18489,N_18722);
or U19753 (N_19753,N_18068,N_18535);
nor U19754 (N_19754,N_18300,N_18756);
nor U19755 (N_19755,N_18410,N_18937);
xnor U19756 (N_19756,N_18893,N_18428);
or U19757 (N_19757,N_18551,N_18733);
and U19758 (N_19758,N_18224,N_18445);
and U19759 (N_19759,N_18751,N_18969);
and U19760 (N_19760,N_18232,N_18203);
nor U19761 (N_19761,N_18115,N_18335);
or U19762 (N_19762,N_18985,N_18651);
or U19763 (N_19763,N_18999,N_18236);
xor U19764 (N_19764,N_18475,N_18280);
or U19765 (N_19765,N_18333,N_18956);
xnor U19766 (N_19766,N_18779,N_18253);
nor U19767 (N_19767,N_18399,N_18842);
xor U19768 (N_19768,N_18150,N_18823);
nand U19769 (N_19769,N_18782,N_18695);
and U19770 (N_19770,N_18325,N_18530);
or U19771 (N_19771,N_18964,N_18308);
and U19772 (N_19772,N_18316,N_18044);
or U19773 (N_19773,N_18968,N_18655);
xor U19774 (N_19774,N_18162,N_18231);
nand U19775 (N_19775,N_18903,N_18618);
or U19776 (N_19776,N_18575,N_18056);
or U19777 (N_19777,N_18192,N_18598);
xnor U19778 (N_19778,N_18159,N_18305);
or U19779 (N_19779,N_18542,N_18620);
and U19780 (N_19780,N_18088,N_18600);
xnor U19781 (N_19781,N_18921,N_18379);
or U19782 (N_19782,N_18150,N_18953);
and U19783 (N_19783,N_18560,N_18424);
nand U19784 (N_19784,N_18677,N_18837);
nand U19785 (N_19785,N_18529,N_18470);
nor U19786 (N_19786,N_18155,N_18475);
and U19787 (N_19787,N_18083,N_18114);
or U19788 (N_19788,N_18106,N_18176);
xor U19789 (N_19789,N_18576,N_18488);
or U19790 (N_19790,N_18595,N_18973);
and U19791 (N_19791,N_18183,N_18493);
xor U19792 (N_19792,N_18480,N_18003);
or U19793 (N_19793,N_18672,N_18584);
nor U19794 (N_19794,N_18156,N_18892);
nor U19795 (N_19795,N_18771,N_18657);
nand U19796 (N_19796,N_18426,N_18822);
nor U19797 (N_19797,N_18785,N_18341);
nand U19798 (N_19798,N_18745,N_18721);
nor U19799 (N_19799,N_18228,N_18743);
or U19800 (N_19800,N_18054,N_18680);
and U19801 (N_19801,N_18162,N_18731);
nor U19802 (N_19802,N_18442,N_18021);
nor U19803 (N_19803,N_18796,N_18993);
xnor U19804 (N_19804,N_18191,N_18444);
nand U19805 (N_19805,N_18064,N_18667);
or U19806 (N_19806,N_18933,N_18975);
nand U19807 (N_19807,N_18362,N_18057);
nor U19808 (N_19808,N_18487,N_18221);
or U19809 (N_19809,N_18406,N_18708);
xnor U19810 (N_19810,N_18937,N_18763);
nand U19811 (N_19811,N_18624,N_18046);
and U19812 (N_19812,N_18781,N_18284);
nor U19813 (N_19813,N_18939,N_18133);
nand U19814 (N_19814,N_18965,N_18921);
or U19815 (N_19815,N_18673,N_18417);
nor U19816 (N_19816,N_18055,N_18014);
or U19817 (N_19817,N_18176,N_18104);
or U19818 (N_19818,N_18726,N_18005);
and U19819 (N_19819,N_18523,N_18726);
or U19820 (N_19820,N_18327,N_18152);
xor U19821 (N_19821,N_18958,N_18925);
xor U19822 (N_19822,N_18210,N_18510);
and U19823 (N_19823,N_18467,N_18424);
xnor U19824 (N_19824,N_18098,N_18223);
or U19825 (N_19825,N_18766,N_18356);
nand U19826 (N_19826,N_18524,N_18698);
or U19827 (N_19827,N_18704,N_18128);
and U19828 (N_19828,N_18215,N_18672);
nor U19829 (N_19829,N_18374,N_18695);
nor U19830 (N_19830,N_18595,N_18699);
nand U19831 (N_19831,N_18050,N_18733);
nand U19832 (N_19832,N_18226,N_18921);
xor U19833 (N_19833,N_18151,N_18082);
xnor U19834 (N_19834,N_18239,N_18856);
and U19835 (N_19835,N_18604,N_18352);
and U19836 (N_19836,N_18221,N_18708);
xnor U19837 (N_19837,N_18083,N_18321);
or U19838 (N_19838,N_18605,N_18247);
xnor U19839 (N_19839,N_18719,N_18999);
and U19840 (N_19840,N_18425,N_18189);
nand U19841 (N_19841,N_18570,N_18782);
or U19842 (N_19842,N_18653,N_18368);
nor U19843 (N_19843,N_18835,N_18480);
xor U19844 (N_19844,N_18754,N_18488);
xnor U19845 (N_19845,N_18257,N_18198);
or U19846 (N_19846,N_18347,N_18339);
nor U19847 (N_19847,N_18865,N_18309);
or U19848 (N_19848,N_18440,N_18152);
and U19849 (N_19849,N_18532,N_18463);
nand U19850 (N_19850,N_18222,N_18937);
and U19851 (N_19851,N_18813,N_18658);
and U19852 (N_19852,N_18584,N_18211);
and U19853 (N_19853,N_18328,N_18961);
or U19854 (N_19854,N_18415,N_18916);
and U19855 (N_19855,N_18278,N_18627);
nand U19856 (N_19856,N_18009,N_18160);
and U19857 (N_19857,N_18135,N_18837);
and U19858 (N_19858,N_18870,N_18347);
nand U19859 (N_19859,N_18840,N_18696);
xor U19860 (N_19860,N_18843,N_18442);
and U19861 (N_19861,N_18635,N_18792);
or U19862 (N_19862,N_18642,N_18653);
nor U19863 (N_19863,N_18851,N_18206);
and U19864 (N_19864,N_18185,N_18548);
nor U19865 (N_19865,N_18356,N_18281);
nand U19866 (N_19866,N_18424,N_18408);
xnor U19867 (N_19867,N_18095,N_18513);
nand U19868 (N_19868,N_18819,N_18477);
and U19869 (N_19869,N_18071,N_18147);
or U19870 (N_19870,N_18154,N_18846);
nand U19871 (N_19871,N_18101,N_18041);
or U19872 (N_19872,N_18266,N_18048);
nor U19873 (N_19873,N_18064,N_18278);
or U19874 (N_19874,N_18953,N_18473);
and U19875 (N_19875,N_18238,N_18874);
and U19876 (N_19876,N_18425,N_18585);
xor U19877 (N_19877,N_18329,N_18250);
nor U19878 (N_19878,N_18809,N_18044);
and U19879 (N_19879,N_18219,N_18447);
and U19880 (N_19880,N_18466,N_18707);
xnor U19881 (N_19881,N_18038,N_18068);
or U19882 (N_19882,N_18325,N_18463);
nand U19883 (N_19883,N_18304,N_18257);
nor U19884 (N_19884,N_18869,N_18560);
xor U19885 (N_19885,N_18344,N_18660);
and U19886 (N_19886,N_18269,N_18477);
and U19887 (N_19887,N_18880,N_18651);
and U19888 (N_19888,N_18899,N_18781);
and U19889 (N_19889,N_18983,N_18336);
and U19890 (N_19890,N_18044,N_18066);
and U19891 (N_19891,N_18728,N_18997);
nor U19892 (N_19892,N_18381,N_18131);
xnor U19893 (N_19893,N_18733,N_18314);
or U19894 (N_19894,N_18825,N_18551);
xor U19895 (N_19895,N_18598,N_18293);
and U19896 (N_19896,N_18721,N_18403);
or U19897 (N_19897,N_18158,N_18109);
and U19898 (N_19898,N_18094,N_18287);
nand U19899 (N_19899,N_18837,N_18301);
xor U19900 (N_19900,N_18722,N_18095);
xnor U19901 (N_19901,N_18253,N_18579);
or U19902 (N_19902,N_18145,N_18922);
nor U19903 (N_19903,N_18604,N_18174);
and U19904 (N_19904,N_18097,N_18444);
nor U19905 (N_19905,N_18782,N_18552);
xnor U19906 (N_19906,N_18460,N_18165);
nand U19907 (N_19907,N_18965,N_18378);
nor U19908 (N_19908,N_18470,N_18511);
and U19909 (N_19909,N_18612,N_18482);
xor U19910 (N_19910,N_18791,N_18748);
xnor U19911 (N_19911,N_18285,N_18721);
xor U19912 (N_19912,N_18857,N_18813);
and U19913 (N_19913,N_18038,N_18380);
or U19914 (N_19914,N_18169,N_18645);
xnor U19915 (N_19915,N_18871,N_18385);
nor U19916 (N_19916,N_18266,N_18275);
nor U19917 (N_19917,N_18868,N_18080);
and U19918 (N_19918,N_18423,N_18297);
or U19919 (N_19919,N_18580,N_18080);
nor U19920 (N_19920,N_18903,N_18049);
and U19921 (N_19921,N_18276,N_18220);
or U19922 (N_19922,N_18276,N_18645);
or U19923 (N_19923,N_18961,N_18546);
nor U19924 (N_19924,N_18793,N_18792);
nor U19925 (N_19925,N_18175,N_18733);
nand U19926 (N_19926,N_18639,N_18190);
and U19927 (N_19927,N_18275,N_18165);
nand U19928 (N_19928,N_18965,N_18182);
or U19929 (N_19929,N_18423,N_18146);
or U19930 (N_19930,N_18952,N_18305);
or U19931 (N_19931,N_18836,N_18675);
nand U19932 (N_19932,N_18401,N_18006);
nand U19933 (N_19933,N_18273,N_18332);
xnor U19934 (N_19934,N_18890,N_18260);
nand U19935 (N_19935,N_18874,N_18598);
xor U19936 (N_19936,N_18113,N_18789);
and U19937 (N_19937,N_18315,N_18027);
or U19938 (N_19938,N_18037,N_18441);
xor U19939 (N_19939,N_18715,N_18997);
and U19940 (N_19940,N_18260,N_18352);
or U19941 (N_19941,N_18540,N_18552);
nor U19942 (N_19942,N_18099,N_18008);
or U19943 (N_19943,N_18562,N_18839);
and U19944 (N_19944,N_18535,N_18156);
nand U19945 (N_19945,N_18075,N_18847);
xor U19946 (N_19946,N_18990,N_18036);
xor U19947 (N_19947,N_18296,N_18108);
nor U19948 (N_19948,N_18429,N_18523);
xnor U19949 (N_19949,N_18445,N_18032);
nand U19950 (N_19950,N_18505,N_18091);
xnor U19951 (N_19951,N_18209,N_18632);
and U19952 (N_19952,N_18409,N_18901);
nand U19953 (N_19953,N_18092,N_18944);
or U19954 (N_19954,N_18275,N_18399);
or U19955 (N_19955,N_18680,N_18451);
nand U19956 (N_19956,N_18638,N_18064);
nand U19957 (N_19957,N_18854,N_18628);
xnor U19958 (N_19958,N_18564,N_18033);
xnor U19959 (N_19959,N_18182,N_18313);
or U19960 (N_19960,N_18342,N_18765);
nand U19961 (N_19961,N_18443,N_18939);
nand U19962 (N_19962,N_18384,N_18271);
xnor U19963 (N_19963,N_18248,N_18086);
nand U19964 (N_19964,N_18507,N_18931);
and U19965 (N_19965,N_18349,N_18203);
nand U19966 (N_19966,N_18049,N_18395);
nor U19967 (N_19967,N_18965,N_18294);
nand U19968 (N_19968,N_18489,N_18590);
xnor U19969 (N_19969,N_18128,N_18691);
or U19970 (N_19970,N_18028,N_18602);
or U19971 (N_19971,N_18097,N_18009);
or U19972 (N_19972,N_18572,N_18175);
and U19973 (N_19973,N_18057,N_18816);
nand U19974 (N_19974,N_18237,N_18838);
or U19975 (N_19975,N_18009,N_18573);
nor U19976 (N_19976,N_18579,N_18501);
or U19977 (N_19977,N_18350,N_18216);
nor U19978 (N_19978,N_18668,N_18096);
xnor U19979 (N_19979,N_18626,N_18122);
nand U19980 (N_19980,N_18886,N_18862);
nand U19981 (N_19981,N_18161,N_18533);
xor U19982 (N_19982,N_18973,N_18554);
nor U19983 (N_19983,N_18730,N_18786);
nor U19984 (N_19984,N_18990,N_18102);
nor U19985 (N_19985,N_18389,N_18639);
and U19986 (N_19986,N_18352,N_18111);
nor U19987 (N_19987,N_18449,N_18860);
nor U19988 (N_19988,N_18986,N_18881);
nor U19989 (N_19989,N_18358,N_18190);
and U19990 (N_19990,N_18811,N_18425);
nor U19991 (N_19991,N_18988,N_18195);
nor U19992 (N_19992,N_18891,N_18539);
nor U19993 (N_19993,N_18407,N_18635);
nor U19994 (N_19994,N_18003,N_18118);
xor U19995 (N_19995,N_18621,N_18927);
nand U19996 (N_19996,N_18088,N_18547);
nand U19997 (N_19997,N_18485,N_18555);
and U19998 (N_19998,N_18936,N_18210);
nor U19999 (N_19999,N_18390,N_18997);
nor UO_0 (O_0,N_19843,N_19695);
and UO_1 (O_1,N_19103,N_19663);
xnor UO_2 (O_2,N_19683,N_19460);
xor UO_3 (O_3,N_19694,N_19349);
or UO_4 (O_4,N_19345,N_19706);
and UO_5 (O_5,N_19799,N_19909);
xnor UO_6 (O_6,N_19350,N_19403);
nand UO_7 (O_7,N_19541,N_19654);
nand UO_8 (O_8,N_19488,N_19729);
nor UO_9 (O_9,N_19508,N_19887);
or UO_10 (O_10,N_19859,N_19959);
and UO_11 (O_11,N_19133,N_19608);
and UO_12 (O_12,N_19090,N_19233);
nand UO_13 (O_13,N_19207,N_19225);
nand UO_14 (O_14,N_19626,N_19670);
and UO_15 (O_15,N_19879,N_19195);
nor UO_16 (O_16,N_19443,N_19392);
nand UO_17 (O_17,N_19389,N_19317);
or UO_18 (O_18,N_19358,N_19245);
nor UO_19 (O_19,N_19610,N_19682);
nor UO_20 (O_20,N_19364,N_19194);
or UO_21 (O_21,N_19014,N_19136);
and UO_22 (O_22,N_19641,N_19698);
nand UO_23 (O_23,N_19647,N_19660);
and UO_24 (O_24,N_19519,N_19646);
nand UO_25 (O_25,N_19015,N_19927);
nor UO_26 (O_26,N_19107,N_19946);
nor UO_27 (O_27,N_19562,N_19383);
nor UO_28 (O_28,N_19664,N_19065);
or UO_29 (O_29,N_19415,N_19411);
or UO_30 (O_30,N_19800,N_19168);
and UO_31 (O_31,N_19188,N_19692);
or UO_32 (O_32,N_19991,N_19412);
xor UO_33 (O_33,N_19330,N_19889);
and UO_34 (O_34,N_19475,N_19275);
or UO_35 (O_35,N_19602,N_19193);
nand UO_36 (O_36,N_19878,N_19972);
or UO_37 (O_37,N_19144,N_19752);
or UO_38 (O_38,N_19061,N_19622);
xor UO_39 (O_39,N_19224,N_19722);
or UO_40 (O_40,N_19551,N_19078);
or UO_41 (O_41,N_19053,N_19650);
and UO_42 (O_42,N_19669,N_19542);
and UO_43 (O_43,N_19156,N_19786);
nand UO_44 (O_44,N_19395,N_19416);
xor UO_45 (O_45,N_19742,N_19766);
or UO_46 (O_46,N_19322,N_19979);
nand UO_47 (O_47,N_19597,N_19110);
nand UO_48 (O_48,N_19578,N_19426);
nor UO_49 (O_49,N_19679,N_19268);
nor UO_50 (O_50,N_19405,N_19009);
or UO_51 (O_51,N_19720,N_19446);
xnor UO_52 (O_52,N_19221,N_19727);
nand UO_53 (O_53,N_19943,N_19662);
and UO_54 (O_54,N_19713,N_19584);
and UO_55 (O_55,N_19005,N_19814);
and UO_56 (O_56,N_19673,N_19655);
nor UO_57 (O_57,N_19604,N_19039);
nor UO_58 (O_58,N_19875,N_19234);
nand UO_59 (O_59,N_19605,N_19784);
nor UO_60 (O_60,N_19049,N_19585);
xor UO_61 (O_61,N_19920,N_19261);
or UO_62 (O_62,N_19581,N_19970);
nor UO_63 (O_63,N_19815,N_19924);
or UO_64 (O_64,N_19371,N_19677);
or UO_65 (O_65,N_19848,N_19525);
and UO_66 (O_66,N_19811,N_19229);
and UO_67 (O_67,N_19063,N_19068);
nor UO_68 (O_68,N_19201,N_19770);
or UO_69 (O_69,N_19771,N_19747);
or UO_70 (O_70,N_19950,N_19079);
nor UO_71 (O_71,N_19885,N_19262);
or UO_72 (O_72,N_19644,N_19387);
or UO_73 (O_73,N_19477,N_19997);
or UO_74 (O_74,N_19408,N_19466);
nand UO_75 (O_75,N_19746,N_19205);
or UO_76 (O_76,N_19938,N_19328);
and UO_77 (O_77,N_19034,N_19978);
or UO_78 (O_78,N_19686,N_19495);
and UO_79 (O_79,N_19560,N_19288);
or UO_80 (O_80,N_19779,N_19983);
nand UO_81 (O_81,N_19504,N_19627);
and UO_82 (O_82,N_19494,N_19896);
or UO_83 (O_83,N_19223,N_19247);
nand UO_84 (O_84,N_19098,N_19863);
and UO_85 (O_85,N_19829,N_19777);
nand UO_86 (O_86,N_19988,N_19294);
or UO_87 (O_87,N_19776,N_19457);
or UO_88 (O_88,N_19217,N_19666);
or UO_89 (O_89,N_19609,N_19081);
xor UO_90 (O_90,N_19115,N_19017);
and UO_91 (O_91,N_19105,N_19936);
xor UO_92 (O_92,N_19676,N_19952);
or UO_93 (O_93,N_19359,N_19678);
nand UO_94 (O_94,N_19296,N_19331);
or UO_95 (O_95,N_19892,N_19547);
or UO_96 (O_96,N_19523,N_19527);
xor UO_97 (O_97,N_19955,N_19071);
or UO_98 (O_98,N_19054,N_19282);
or UO_99 (O_99,N_19222,N_19621);
and UO_100 (O_100,N_19689,N_19113);
nand UO_101 (O_101,N_19376,N_19157);
nand UO_102 (O_102,N_19471,N_19176);
nand UO_103 (O_103,N_19351,N_19973);
xnor UO_104 (O_104,N_19898,N_19012);
nand UO_105 (O_105,N_19555,N_19391);
or UO_106 (O_106,N_19906,N_19763);
nor UO_107 (O_107,N_19515,N_19968);
and UO_108 (O_108,N_19084,N_19092);
or UO_109 (O_109,N_19482,N_19355);
and UO_110 (O_110,N_19088,N_19599);
xor UO_111 (O_111,N_19546,N_19553);
nor UO_112 (O_112,N_19214,N_19062);
xnor UO_113 (O_113,N_19064,N_19513);
xnor UO_114 (O_114,N_19143,N_19171);
and UO_115 (O_115,N_19883,N_19087);
nand UO_116 (O_116,N_19280,N_19452);
nor UO_117 (O_117,N_19458,N_19091);
and UO_118 (O_118,N_19192,N_19616);
and UO_119 (O_119,N_19321,N_19831);
or UO_120 (O_120,N_19998,N_19787);
nand UO_121 (O_121,N_19719,N_19919);
and UO_122 (O_122,N_19227,N_19797);
or UO_123 (O_123,N_19659,N_19051);
nand UO_124 (O_124,N_19667,N_19318);
or UO_125 (O_125,N_19394,N_19618);
or UO_126 (O_126,N_19963,N_19638);
nand UO_127 (O_127,N_19739,N_19237);
nor UO_128 (O_128,N_19570,N_19145);
or UO_129 (O_129,N_19612,N_19985);
nor UO_130 (O_130,N_19632,N_19196);
nor UO_131 (O_131,N_19880,N_19102);
and UO_132 (O_132,N_19400,N_19285);
xnor UO_133 (O_133,N_19147,N_19945);
nor UO_134 (O_134,N_19949,N_19661);
nor UO_135 (O_135,N_19552,N_19606);
nor UO_136 (O_136,N_19703,N_19451);
nand UO_137 (O_137,N_19002,N_19545);
and UO_138 (O_138,N_19381,N_19429);
and UO_139 (O_139,N_19165,N_19121);
nor UO_140 (O_140,N_19700,N_19559);
xnor UO_141 (O_141,N_19388,N_19530);
nand UO_142 (O_142,N_19208,N_19941);
and UO_143 (O_143,N_19158,N_19045);
nand UO_144 (O_144,N_19790,N_19709);
or UO_145 (O_145,N_19414,N_19750);
xor UO_146 (O_146,N_19272,N_19357);
nor UO_147 (O_147,N_19726,N_19639);
nor UO_148 (O_148,N_19109,N_19302);
and UO_149 (O_149,N_19010,N_19620);
xor UO_150 (O_150,N_19309,N_19827);
or UO_151 (O_151,N_19514,N_19636);
nor UO_152 (O_152,N_19303,N_19575);
and UO_153 (O_153,N_19313,N_19292);
xor UO_154 (O_154,N_19615,N_19888);
or UO_155 (O_155,N_19314,N_19837);
xor UO_156 (O_156,N_19436,N_19390);
nand UO_157 (O_157,N_19496,N_19561);
nor UO_158 (O_158,N_19821,N_19995);
xor UO_159 (O_159,N_19152,N_19286);
nand UO_160 (O_160,N_19339,N_19982);
and UO_161 (O_161,N_19824,N_19455);
nand UO_162 (O_162,N_19755,N_19297);
xnor UO_163 (O_163,N_19765,N_19178);
nor UO_164 (O_164,N_19693,N_19326);
and UO_165 (O_165,N_19440,N_19213);
and UO_166 (O_166,N_19465,N_19601);
and UO_167 (O_167,N_19377,N_19532);
or UO_168 (O_168,N_19928,N_19674);
or UO_169 (O_169,N_19238,N_19876);
nand UO_170 (O_170,N_19430,N_19834);
and UO_171 (O_171,N_19645,N_19424);
nand UO_172 (O_172,N_19707,N_19406);
xor UO_173 (O_173,N_19050,N_19806);
nor UO_174 (O_174,N_19839,N_19960);
or UO_175 (O_175,N_19220,N_19981);
and UO_176 (O_176,N_19454,N_19264);
xnor UO_177 (O_177,N_19069,N_19382);
xor UO_178 (O_178,N_19472,N_19628);
and UO_179 (O_179,N_19944,N_19492);
or UO_180 (O_180,N_19954,N_19582);
and UO_181 (O_181,N_19757,N_19200);
nand UO_182 (O_182,N_19187,N_19085);
nor UO_183 (O_183,N_19951,N_19183);
xor UO_184 (O_184,N_19315,N_19521);
nor UO_185 (O_185,N_19216,N_19431);
nor UO_186 (O_186,N_19059,N_19023);
or UO_187 (O_187,N_19930,N_19688);
and UO_188 (O_188,N_19191,N_19218);
nand UO_189 (O_189,N_19256,N_19625);
and UO_190 (O_190,N_19868,N_19587);
nor UO_191 (O_191,N_19802,N_19231);
and UO_192 (O_192,N_19818,N_19278);
xnor UO_193 (O_193,N_19796,N_19668);
xnor UO_194 (O_194,N_19869,N_19574);
or UO_195 (O_195,N_19226,N_19271);
nor UO_196 (O_196,N_19718,N_19461);
or UO_197 (O_197,N_19897,N_19600);
and UO_198 (O_198,N_19365,N_19798);
or UO_199 (O_199,N_19232,N_19576);
nand UO_200 (O_200,N_19864,N_19623);
and UO_201 (O_201,N_19816,N_19586);
nor UO_202 (O_202,N_19792,N_19011);
and UO_203 (O_203,N_19701,N_19146);
nand UO_204 (O_204,N_19439,N_19934);
xor UO_205 (O_205,N_19550,N_19476);
and UO_206 (O_206,N_19468,N_19409);
nand UO_207 (O_207,N_19912,N_19500);
and UO_208 (O_208,N_19535,N_19259);
xor UO_209 (O_209,N_19836,N_19298);
xor UO_210 (O_210,N_19649,N_19828);
nand UO_211 (O_211,N_19375,N_19048);
nor UO_212 (O_212,N_19691,N_19336);
or UO_213 (O_213,N_19164,N_19489);
or UO_214 (O_214,N_19994,N_19379);
nand UO_215 (O_215,N_19714,N_19179);
xor UO_216 (O_216,N_19058,N_19166);
and UO_217 (O_217,N_19738,N_19511);
and UO_218 (O_218,N_19258,N_19057);
nand UO_219 (O_219,N_19856,N_19823);
nand UO_220 (O_220,N_19710,N_19174);
nor UO_221 (O_221,N_19041,N_19253);
and UO_222 (O_222,N_19789,N_19175);
nand UO_223 (O_223,N_19520,N_19281);
xnor UO_224 (O_224,N_19373,N_19420);
xor UO_225 (O_225,N_19470,N_19252);
nand UO_226 (O_226,N_19717,N_19242);
xor UO_227 (O_227,N_19124,N_19347);
xnor UO_228 (O_228,N_19185,N_19913);
or UO_229 (O_229,N_19072,N_19751);
or UO_230 (O_230,N_19548,N_19544);
and UO_231 (O_231,N_19076,N_19246);
xnor UO_232 (O_232,N_19360,N_19055);
or UO_233 (O_233,N_19159,N_19918);
nand UO_234 (O_234,N_19337,N_19611);
nor UO_235 (O_235,N_19060,N_19731);
xnor UO_236 (O_236,N_19507,N_19239);
nor UO_237 (O_237,N_19533,N_19154);
or UO_238 (O_238,N_19635,N_19557);
or UO_239 (O_239,N_19130,N_19308);
and UO_240 (O_240,N_19228,N_19740);
or UO_241 (O_241,N_19704,N_19111);
or UO_242 (O_242,N_19984,N_19402);
or UO_243 (O_243,N_19480,N_19531);
or UO_244 (O_244,N_19840,N_19184);
and UO_245 (O_245,N_19456,N_19697);
xnor UO_246 (O_246,N_19453,N_19736);
or UO_247 (O_247,N_19029,N_19580);
or UO_248 (O_248,N_19172,N_19096);
xor UO_249 (O_249,N_19737,N_19540);
or UO_250 (O_250,N_19665,N_19131);
xor UO_251 (O_251,N_19760,N_19290);
nand UO_252 (O_252,N_19125,N_19181);
and UO_253 (O_253,N_19190,N_19528);
and UO_254 (O_254,N_19398,N_19120);
nand UO_255 (O_255,N_19705,N_19781);
nor UO_256 (O_256,N_19101,N_19594);
xnor UO_257 (O_257,N_19671,N_19043);
or UO_258 (O_258,N_19119,N_19539);
and UO_259 (O_259,N_19524,N_19442);
and UO_260 (O_260,N_19907,N_19648);
or UO_261 (O_261,N_19123,N_19969);
xnor UO_262 (O_262,N_19491,N_19447);
nor UO_263 (O_263,N_19329,N_19173);
or UO_264 (O_264,N_19073,N_19592);
nor UO_265 (O_265,N_19020,N_19316);
nor UO_266 (O_266,N_19013,N_19980);
nand UO_267 (O_267,N_19257,N_19761);
nor UO_268 (O_268,N_19947,N_19418);
nand UO_269 (O_269,N_19031,N_19803);
xnor UO_270 (O_270,N_19932,N_19813);
nor UO_271 (O_271,N_19445,N_19785);
nand UO_272 (O_272,N_19254,N_19826);
xnor UO_273 (O_273,N_19093,N_19744);
xnor UO_274 (O_274,N_19975,N_19342);
nor UO_275 (O_275,N_19128,N_19871);
xor UO_276 (O_276,N_19699,N_19853);
xnor UO_277 (O_277,N_19967,N_19835);
nand UO_278 (O_278,N_19203,N_19640);
nand UO_279 (O_279,N_19767,N_19681);
xor UO_280 (O_280,N_19267,N_19807);
nand UO_281 (O_281,N_19723,N_19596);
xnor UO_282 (O_282,N_19306,N_19624);
or UO_283 (O_283,N_19629,N_19884);
nand UO_284 (O_284,N_19464,N_19338);
nor UO_285 (O_285,N_19566,N_19872);
and UO_286 (O_286,N_19502,N_19046);
or UO_287 (O_287,N_19805,N_19086);
and UO_288 (O_288,N_19865,N_19895);
or UO_289 (O_289,N_19177,N_19385);
nand UO_290 (O_290,N_19774,N_19304);
and UO_291 (O_291,N_19240,N_19926);
and UO_292 (O_292,N_19450,N_19958);
nor UO_293 (O_293,N_19543,N_19916);
and UO_294 (O_294,N_19483,N_19095);
xor UO_295 (O_295,N_19211,N_19169);
nor UO_296 (O_296,N_19449,N_19287);
xor UO_297 (O_297,N_19501,N_19577);
nand UO_298 (O_298,N_19197,N_19487);
nand UO_299 (O_299,N_19685,N_19891);
xor UO_300 (O_300,N_19127,N_19044);
xor UO_301 (O_301,N_19432,N_19808);
and UO_302 (O_302,N_19966,N_19964);
nand UO_303 (O_303,N_19595,N_19914);
and UO_304 (O_304,N_19748,N_19343);
or UO_305 (O_305,N_19728,N_19003);
and UO_306 (O_306,N_19890,N_19858);
or UO_307 (O_307,N_19822,N_19617);
nor UO_308 (O_308,N_19568,N_19957);
nand UO_309 (O_309,N_19484,N_19516);
xnor UO_310 (O_310,N_19911,N_19499);
and UO_311 (O_311,N_19052,N_19032);
nand UO_312 (O_312,N_19354,N_19793);
nand UO_313 (O_313,N_19372,N_19633);
nand UO_314 (O_314,N_19311,N_19108);
or UO_315 (O_315,N_19490,N_19780);
and UO_316 (O_316,N_19850,N_19153);
nor UO_317 (O_317,N_19410,N_19841);
or UO_318 (O_318,N_19189,N_19022);
and UO_319 (O_319,N_19962,N_19462);
xor UO_320 (O_320,N_19348,N_19138);
nand UO_321 (O_321,N_19241,N_19986);
and UO_322 (O_322,N_19277,N_19830);
nand UO_323 (O_323,N_19270,N_19905);
xnor UO_324 (O_324,N_19293,N_19724);
xor UO_325 (O_325,N_19862,N_19929);
nor UO_326 (O_326,N_19142,N_19180);
and UO_327 (O_327,N_19680,N_19399);
xnor UO_328 (O_328,N_19769,N_19498);
xnor UO_329 (O_329,N_19260,N_19908);
xnor UO_330 (O_330,N_19025,N_19778);
nor UO_331 (O_331,N_19413,N_19099);
and UO_332 (O_332,N_19512,N_19937);
xor UO_333 (O_333,N_19572,N_19534);
and UO_334 (O_334,N_19922,N_19027);
nor UO_335 (O_335,N_19199,N_19732);
nand UO_336 (O_336,N_19097,N_19940);
nor UO_337 (O_337,N_19374,N_19782);
nor UO_338 (O_338,N_19148,N_19444);
nand UO_339 (O_339,N_19459,N_19506);
xor UO_340 (O_340,N_19000,N_19056);
nor UO_341 (O_341,N_19833,N_19401);
xnor UO_342 (O_342,N_19538,N_19642);
nor UO_343 (O_343,N_19448,N_19764);
nand UO_344 (O_344,N_19881,N_19104);
nand UO_345 (O_345,N_19526,N_19735);
xor UO_346 (O_346,N_19565,N_19289);
or UO_347 (O_347,N_19140,N_19588);
or UO_348 (O_348,N_19334,N_19652);
xor UO_349 (O_349,N_19441,N_19083);
and UO_350 (O_350,N_19637,N_19509);
nand UO_351 (O_351,N_19265,N_19522);
or UO_352 (O_352,N_19036,N_19900);
xor UO_353 (O_353,N_19033,N_19993);
xor UO_354 (O_354,N_19933,N_19310);
nor UO_355 (O_355,N_19404,N_19161);
and UO_356 (O_356,N_19743,N_19421);
or UO_357 (O_357,N_19077,N_19362);
and UO_358 (O_358,N_19861,N_19849);
and UO_359 (O_359,N_19753,N_19999);
nor UO_360 (O_360,N_19497,N_19899);
xor UO_361 (O_361,N_19614,N_19730);
nand UO_362 (O_362,N_19116,N_19368);
nand UO_363 (O_363,N_19361,N_19363);
or UO_364 (O_364,N_19935,N_19564);
nand UO_365 (O_365,N_19149,N_19437);
and UO_366 (O_366,N_19772,N_19035);
or UO_367 (O_367,N_19974,N_19094);
nor UO_368 (O_368,N_19817,N_19419);
nand UO_369 (O_369,N_19137,N_19019);
or UO_370 (O_370,N_19474,N_19276);
nand UO_371 (O_371,N_19026,N_19870);
and UO_372 (O_372,N_19505,N_19469);
and UO_373 (O_373,N_19163,N_19463);
nand UO_374 (O_374,N_19715,N_19536);
nor UO_375 (O_375,N_19135,N_19129);
nor UO_376 (O_376,N_19942,N_19971);
and UO_377 (O_377,N_19407,N_19956);
nor UO_378 (O_378,N_19204,N_19341);
nand UO_379 (O_379,N_19344,N_19921);
nor UO_380 (O_380,N_19367,N_19915);
or UO_381 (O_381,N_19589,N_19819);
and UO_382 (O_382,N_19518,N_19867);
nand UO_383 (O_383,N_19923,N_19684);
and UO_384 (O_384,N_19768,N_19040);
and UO_385 (O_385,N_19795,N_19579);
xnor UO_386 (O_386,N_19965,N_19283);
nand UO_387 (O_387,N_19007,N_19325);
nand UO_388 (O_388,N_19433,N_19571);
and UO_389 (O_389,N_19619,N_19734);
and UO_390 (O_390,N_19263,N_19209);
or UO_391 (O_391,N_19037,N_19300);
or UO_392 (O_392,N_19369,N_19340);
nor UO_393 (O_393,N_19866,N_19028);
or UO_394 (O_394,N_19366,N_19380);
and UO_395 (O_395,N_19593,N_19702);
or UO_396 (O_396,N_19549,N_19773);
or UO_397 (O_397,N_19687,N_19503);
nor UO_398 (O_398,N_19386,N_19352);
nand UO_399 (O_399,N_19801,N_19473);
and UO_400 (O_400,N_19001,N_19486);
nand UO_401 (O_401,N_19976,N_19070);
and UO_402 (O_402,N_19939,N_19151);
and UO_403 (O_403,N_19598,N_19809);
and UO_404 (O_404,N_19852,N_19112);
xnor UO_405 (O_405,N_19567,N_19591);
or UO_406 (O_406,N_19634,N_19716);
xnor UO_407 (O_407,N_19590,N_19990);
xnor UO_408 (O_408,N_19931,N_19255);
nand UO_409 (O_409,N_19467,N_19393);
nand UO_410 (O_410,N_19708,N_19008);
nand UO_411 (O_411,N_19160,N_19082);
xnor UO_412 (O_412,N_19122,N_19902);
nor UO_413 (O_413,N_19243,N_19904);
nor UO_414 (O_414,N_19977,N_19384);
xnor UO_415 (O_415,N_19794,N_19274);
and UO_416 (O_416,N_19741,N_19134);
and UO_417 (O_417,N_19016,N_19613);
and UO_418 (O_418,N_19106,N_19886);
or UO_419 (O_419,N_19810,N_19038);
nand UO_420 (O_420,N_19024,N_19435);
or UO_421 (O_421,N_19428,N_19485);
or UO_422 (O_422,N_19873,N_19832);
and UO_423 (O_423,N_19067,N_19117);
nor UO_424 (O_424,N_19855,N_19820);
nand UO_425 (O_425,N_19756,N_19877);
xnor UO_426 (O_426,N_19250,N_19917);
or UO_427 (O_427,N_19558,N_19307);
or UO_428 (O_428,N_19126,N_19854);
and UO_429 (O_429,N_19529,N_19248);
nor UO_430 (O_430,N_19847,N_19215);
nor UO_431 (O_431,N_19569,N_19517);
xnor UO_432 (O_432,N_19132,N_19754);
nor UO_433 (O_433,N_19733,N_19273);
nand UO_434 (O_434,N_19346,N_19857);
nor UO_435 (O_435,N_19783,N_19021);
or UO_436 (O_436,N_19324,N_19312);
or UO_437 (O_437,N_19295,N_19696);
xnor UO_438 (O_438,N_19825,N_19323);
xor UO_439 (O_439,N_19657,N_19675);
nand UO_440 (O_440,N_19269,N_19844);
and UO_441 (O_441,N_19987,N_19335);
and UO_442 (O_442,N_19478,N_19066);
nor UO_443 (O_443,N_19320,N_19249);
and UO_444 (O_444,N_19925,N_19235);
xor UO_445 (O_445,N_19251,N_19206);
nor UO_446 (O_446,N_19202,N_19370);
nor UO_447 (O_447,N_19948,N_19953);
or UO_448 (O_448,N_19651,N_19788);
nand UO_449 (O_449,N_19212,N_19846);
or UO_450 (O_450,N_19150,N_19284);
xor UO_451 (O_451,N_19658,N_19573);
xor UO_452 (O_452,N_19333,N_19299);
xor UO_453 (O_453,N_19631,N_19089);
xor UO_454 (O_454,N_19775,N_19356);
nand UO_455 (O_455,N_19901,N_19961);
nand UO_456 (O_456,N_19537,N_19989);
or UO_457 (O_457,N_19378,N_19479);
xnor UO_458 (O_458,N_19155,N_19004);
xnor UO_459 (O_459,N_19417,N_19236);
or UO_460 (O_460,N_19427,N_19860);
and UO_461 (O_461,N_19042,N_19100);
nand UO_462 (O_462,N_19080,N_19162);
nand UO_463 (O_463,N_19759,N_19118);
nor UO_464 (O_464,N_19291,N_19219);
or UO_465 (O_465,N_19423,N_19758);
nand UO_466 (O_466,N_19672,N_19047);
nor UO_467 (O_467,N_19279,N_19845);
xor UO_468 (O_468,N_19583,N_19141);
nand UO_469 (O_469,N_19198,N_19230);
xnor UO_470 (O_470,N_19425,N_19745);
and UO_471 (O_471,N_19327,N_19422);
and UO_472 (O_472,N_19186,N_19434);
or UO_473 (O_473,N_19170,N_19353);
or UO_474 (O_474,N_19030,N_19812);
nor UO_475 (O_475,N_19656,N_19438);
nand UO_476 (O_476,N_19653,N_19725);
nand UO_477 (O_477,N_19210,N_19114);
xnor UO_478 (O_478,N_19244,N_19996);
nor UO_479 (O_479,N_19712,N_19903);
xnor UO_480 (O_480,N_19711,N_19762);
or UO_481 (O_481,N_19167,N_19075);
or UO_482 (O_482,N_19396,N_19894);
and UO_483 (O_483,N_19319,N_19838);
and UO_484 (O_484,N_19305,N_19397);
or UO_485 (O_485,N_19266,N_19554);
and UO_486 (O_486,N_19301,N_19493);
and UO_487 (O_487,N_19690,N_19851);
or UO_488 (O_488,N_19791,N_19630);
and UO_489 (O_489,N_19603,N_19556);
or UO_490 (O_490,N_19893,N_19721);
or UO_491 (O_491,N_19018,N_19749);
and UO_492 (O_492,N_19563,N_19510);
or UO_493 (O_493,N_19804,N_19910);
and UO_494 (O_494,N_19992,N_19139);
nor UO_495 (O_495,N_19643,N_19332);
nor UO_496 (O_496,N_19074,N_19481);
nand UO_497 (O_497,N_19182,N_19006);
or UO_498 (O_498,N_19842,N_19874);
and UO_499 (O_499,N_19607,N_19882);
nor UO_500 (O_500,N_19244,N_19344);
xor UO_501 (O_501,N_19832,N_19784);
or UO_502 (O_502,N_19799,N_19506);
xnor UO_503 (O_503,N_19523,N_19361);
and UO_504 (O_504,N_19825,N_19452);
xor UO_505 (O_505,N_19634,N_19560);
nor UO_506 (O_506,N_19372,N_19543);
nor UO_507 (O_507,N_19940,N_19467);
xnor UO_508 (O_508,N_19517,N_19382);
or UO_509 (O_509,N_19428,N_19959);
nand UO_510 (O_510,N_19592,N_19784);
and UO_511 (O_511,N_19995,N_19492);
xnor UO_512 (O_512,N_19285,N_19427);
and UO_513 (O_513,N_19509,N_19428);
nand UO_514 (O_514,N_19027,N_19614);
nand UO_515 (O_515,N_19728,N_19417);
nor UO_516 (O_516,N_19437,N_19082);
and UO_517 (O_517,N_19824,N_19513);
and UO_518 (O_518,N_19966,N_19789);
xor UO_519 (O_519,N_19733,N_19407);
or UO_520 (O_520,N_19573,N_19767);
or UO_521 (O_521,N_19119,N_19541);
nor UO_522 (O_522,N_19080,N_19699);
and UO_523 (O_523,N_19744,N_19695);
or UO_524 (O_524,N_19587,N_19794);
nor UO_525 (O_525,N_19824,N_19121);
and UO_526 (O_526,N_19493,N_19697);
and UO_527 (O_527,N_19709,N_19251);
xor UO_528 (O_528,N_19267,N_19007);
nand UO_529 (O_529,N_19186,N_19345);
or UO_530 (O_530,N_19909,N_19320);
nor UO_531 (O_531,N_19646,N_19164);
xor UO_532 (O_532,N_19948,N_19687);
xnor UO_533 (O_533,N_19384,N_19288);
and UO_534 (O_534,N_19414,N_19380);
xnor UO_535 (O_535,N_19714,N_19573);
nor UO_536 (O_536,N_19368,N_19777);
xnor UO_537 (O_537,N_19490,N_19627);
nand UO_538 (O_538,N_19236,N_19182);
and UO_539 (O_539,N_19414,N_19400);
or UO_540 (O_540,N_19712,N_19800);
xor UO_541 (O_541,N_19675,N_19871);
nor UO_542 (O_542,N_19111,N_19204);
or UO_543 (O_543,N_19675,N_19251);
or UO_544 (O_544,N_19672,N_19760);
nor UO_545 (O_545,N_19579,N_19229);
and UO_546 (O_546,N_19719,N_19681);
and UO_547 (O_547,N_19932,N_19612);
nand UO_548 (O_548,N_19661,N_19844);
nand UO_549 (O_549,N_19761,N_19570);
nor UO_550 (O_550,N_19949,N_19131);
and UO_551 (O_551,N_19973,N_19444);
xor UO_552 (O_552,N_19708,N_19141);
nand UO_553 (O_553,N_19616,N_19506);
or UO_554 (O_554,N_19940,N_19996);
xnor UO_555 (O_555,N_19076,N_19426);
xnor UO_556 (O_556,N_19807,N_19670);
and UO_557 (O_557,N_19227,N_19703);
or UO_558 (O_558,N_19343,N_19023);
xor UO_559 (O_559,N_19119,N_19239);
nor UO_560 (O_560,N_19397,N_19372);
xor UO_561 (O_561,N_19293,N_19022);
nor UO_562 (O_562,N_19917,N_19411);
xor UO_563 (O_563,N_19979,N_19442);
xor UO_564 (O_564,N_19800,N_19396);
xnor UO_565 (O_565,N_19776,N_19911);
nand UO_566 (O_566,N_19649,N_19150);
xnor UO_567 (O_567,N_19634,N_19741);
xnor UO_568 (O_568,N_19248,N_19722);
nor UO_569 (O_569,N_19943,N_19118);
or UO_570 (O_570,N_19582,N_19162);
xnor UO_571 (O_571,N_19378,N_19976);
or UO_572 (O_572,N_19486,N_19778);
and UO_573 (O_573,N_19012,N_19339);
xnor UO_574 (O_574,N_19183,N_19002);
and UO_575 (O_575,N_19249,N_19062);
or UO_576 (O_576,N_19237,N_19760);
xor UO_577 (O_577,N_19565,N_19037);
or UO_578 (O_578,N_19641,N_19325);
or UO_579 (O_579,N_19597,N_19907);
nor UO_580 (O_580,N_19864,N_19350);
nand UO_581 (O_581,N_19363,N_19963);
nand UO_582 (O_582,N_19371,N_19373);
xor UO_583 (O_583,N_19309,N_19569);
xor UO_584 (O_584,N_19769,N_19093);
xor UO_585 (O_585,N_19781,N_19353);
nand UO_586 (O_586,N_19601,N_19592);
xnor UO_587 (O_587,N_19784,N_19618);
or UO_588 (O_588,N_19508,N_19831);
and UO_589 (O_589,N_19171,N_19808);
xor UO_590 (O_590,N_19512,N_19168);
nor UO_591 (O_591,N_19661,N_19928);
nand UO_592 (O_592,N_19445,N_19917);
and UO_593 (O_593,N_19428,N_19719);
nand UO_594 (O_594,N_19325,N_19820);
and UO_595 (O_595,N_19904,N_19884);
nor UO_596 (O_596,N_19108,N_19028);
and UO_597 (O_597,N_19928,N_19546);
xor UO_598 (O_598,N_19003,N_19458);
xor UO_599 (O_599,N_19087,N_19919);
xor UO_600 (O_600,N_19502,N_19916);
nor UO_601 (O_601,N_19105,N_19201);
xor UO_602 (O_602,N_19529,N_19493);
and UO_603 (O_603,N_19105,N_19748);
xor UO_604 (O_604,N_19724,N_19459);
or UO_605 (O_605,N_19110,N_19056);
or UO_606 (O_606,N_19529,N_19868);
nand UO_607 (O_607,N_19865,N_19412);
and UO_608 (O_608,N_19080,N_19598);
nor UO_609 (O_609,N_19912,N_19104);
or UO_610 (O_610,N_19495,N_19531);
nor UO_611 (O_611,N_19997,N_19571);
nand UO_612 (O_612,N_19968,N_19952);
nor UO_613 (O_613,N_19341,N_19531);
nand UO_614 (O_614,N_19634,N_19938);
or UO_615 (O_615,N_19827,N_19783);
and UO_616 (O_616,N_19830,N_19141);
xnor UO_617 (O_617,N_19644,N_19356);
xor UO_618 (O_618,N_19757,N_19714);
nand UO_619 (O_619,N_19798,N_19340);
or UO_620 (O_620,N_19316,N_19135);
nor UO_621 (O_621,N_19690,N_19639);
nor UO_622 (O_622,N_19688,N_19571);
nand UO_623 (O_623,N_19725,N_19002);
xor UO_624 (O_624,N_19366,N_19199);
nand UO_625 (O_625,N_19266,N_19815);
nand UO_626 (O_626,N_19169,N_19215);
or UO_627 (O_627,N_19619,N_19091);
xnor UO_628 (O_628,N_19493,N_19415);
nor UO_629 (O_629,N_19128,N_19381);
xor UO_630 (O_630,N_19689,N_19581);
or UO_631 (O_631,N_19985,N_19525);
nor UO_632 (O_632,N_19506,N_19092);
or UO_633 (O_633,N_19433,N_19172);
and UO_634 (O_634,N_19561,N_19763);
nor UO_635 (O_635,N_19743,N_19354);
nand UO_636 (O_636,N_19531,N_19083);
nand UO_637 (O_637,N_19165,N_19363);
and UO_638 (O_638,N_19855,N_19699);
and UO_639 (O_639,N_19175,N_19872);
nor UO_640 (O_640,N_19208,N_19129);
xnor UO_641 (O_641,N_19620,N_19265);
nor UO_642 (O_642,N_19475,N_19172);
and UO_643 (O_643,N_19651,N_19839);
and UO_644 (O_644,N_19410,N_19681);
xnor UO_645 (O_645,N_19608,N_19336);
or UO_646 (O_646,N_19606,N_19656);
xor UO_647 (O_647,N_19082,N_19279);
or UO_648 (O_648,N_19383,N_19427);
and UO_649 (O_649,N_19298,N_19337);
xor UO_650 (O_650,N_19172,N_19984);
nand UO_651 (O_651,N_19392,N_19971);
nor UO_652 (O_652,N_19041,N_19871);
xnor UO_653 (O_653,N_19180,N_19500);
xor UO_654 (O_654,N_19871,N_19809);
and UO_655 (O_655,N_19493,N_19681);
or UO_656 (O_656,N_19052,N_19261);
nor UO_657 (O_657,N_19181,N_19447);
xor UO_658 (O_658,N_19320,N_19400);
or UO_659 (O_659,N_19999,N_19809);
xnor UO_660 (O_660,N_19754,N_19530);
and UO_661 (O_661,N_19958,N_19010);
or UO_662 (O_662,N_19321,N_19130);
and UO_663 (O_663,N_19187,N_19503);
or UO_664 (O_664,N_19737,N_19521);
xnor UO_665 (O_665,N_19566,N_19109);
and UO_666 (O_666,N_19210,N_19541);
nand UO_667 (O_667,N_19176,N_19390);
xor UO_668 (O_668,N_19166,N_19891);
nor UO_669 (O_669,N_19252,N_19595);
and UO_670 (O_670,N_19509,N_19508);
xor UO_671 (O_671,N_19728,N_19378);
and UO_672 (O_672,N_19439,N_19512);
nand UO_673 (O_673,N_19451,N_19477);
or UO_674 (O_674,N_19750,N_19308);
nor UO_675 (O_675,N_19403,N_19636);
nand UO_676 (O_676,N_19371,N_19770);
and UO_677 (O_677,N_19815,N_19311);
xnor UO_678 (O_678,N_19883,N_19422);
xor UO_679 (O_679,N_19724,N_19836);
nor UO_680 (O_680,N_19197,N_19758);
and UO_681 (O_681,N_19681,N_19688);
nor UO_682 (O_682,N_19332,N_19661);
or UO_683 (O_683,N_19239,N_19447);
xor UO_684 (O_684,N_19835,N_19800);
or UO_685 (O_685,N_19646,N_19699);
xor UO_686 (O_686,N_19881,N_19928);
or UO_687 (O_687,N_19743,N_19431);
or UO_688 (O_688,N_19999,N_19396);
nor UO_689 (O_689,N_19176,N_19796);
or UO_690 (O_690,N_19475,N_19840);
nor UO_691 (O_691,N_19059,N_19029);
and UO_692 (O_692,N_19502,N_19689);
or UO_693 (O_693,N_19952,N_19732);
xnor UO_694 (O_694,N_19706,N_19197);
nor UO_695 (O_695,N_19917,N_19508);
nand UO_696 (O_696,N_19292,N_19085);
nand UO_697 (O_697,N_19836,N_19987);
nand UO_698 (O_698,N_19200,N_19920);
nor UO_699 (O_699,N_19484,N_19227);
xnor UO_700 (O_700,N_19580,N_19239);
xor UO_701 (O_701,N_19997,N_19760);
xnor UO_702 (O_702,N_19588,N_19188);
nand UO_703 (O_703,N_19208,N_19393);
xnor UO_704 (O_704,N_19826,N_19870);
nand UO_705 (O_705,N_19127,N_19179);
or UO_706 (O_706,N_19402,N_19508);
or UO_707 (O_707,N_19317,N_19380);
nand UO_708 (O_708,N_19397,N_19441);
nand UO_709 (O_709,N_19628,N_19831);
and UO_710 (O_710,N_19335,N_19087);
nand UO_711 (O_711,N_19530,N_19902);
or UO_712 (O_712,N_19418,N_19172);
and UO_713 (O_713,N_19880,N_19065);
nor UO_714 (O_714,N_19216,N_19336);
or UO_715 (O_715,N_19555,N_19217);
nand UO_716 (O_716,N_19068,N_19579);
xor UO_717 (O_717,N_19645,N_19308);
and UO_718 (O_718,N_19831,N_19938);
nor UO_719 (O_719,N_19867,N_19834);
nand UO_720 (O_720,N_19503,N_19500);
xor UO_721 (O_721,N_19963,N_19743);
nand UO_722 (O_722,N_19707,N_19228);
xor UO_723 (O_723,N_19161,N_19481);
xor UO_724 (O_724,N_19634,N_19080);
or UO_725 (O_725,N_19823,N_19338);
nor UO_726 (O_726,N_19840,N_19859);
nor UO_727 (O_727,N_19877,N_19360);
or UO_728 (O_728,N_19504,N_19088);
or UO_729 (O_729,N_19159,N_19368);
nand UO_730 (O_730,N_19897,N_19455);
xor UO_731 (O_731,N_19724,N_19608);
nand UO_732 (O_732,N_19685,N_19323);
and UO_733 (O_733,N_19163,N_19635);
xnor UO_734 (O_734,N_19307,N_19352);
xor UO_735 (O_735,N_19473,N_19939);
xor UO_736 (O_736,N_19850,N_19666);
xnor UO_737 (O_737,N_19784,N_19791);
nor UO_738 (O_738,N_19302,N_19732);
or UO_739 (O_739,N_19969,N_19615);
nand UO_740 (O_740,N_19271,N_19557);
or UO_741 (O_741,N_19587,N_19859);
nor UO_742 (O_742,N_19046,N_19177);
xnor UO_743 (O_743,N_19401,N_19018);
xnor UO_744 (O_744,N_19383,N_19925);
or UO_745 (O_745,N_19718,N_19427);
nor UO_746 (O_746,N_19853,N_19828);
or UO_747 (O_747,N_19218,N_19994);
xnor UO_748 (O_748,N_19458,N_19171);
nand UO_749 (O_749,N_19816,N_19858);
or UO_750 (O_750,N_19672,N_19859);
nor UO_751 (O_751,N_19829,N_19174);
xor UO_752 (O_752,N_19517,N_19666);
nor UO_753 (O_753,N_19369,N_19735);
nor UO_754 (O_754,N_19806,N_19353);
nand UO_755 (O_755,N_19049,N_19589);
and UO_756 (O_756,N_19033,N_19423);
nand UO_757 (O_757,N_19500,N_19829);
or UO_758 (O_758,N_19001,N_19641);
nor UO_759 (O_759,N_19199,N_19919);
and UO_760 (O_760,N_19205,N_19537);
nor UO_761 (O_761,N_19576,N_19459);
and UO_762 (O_762,N_19279,N_19496);
or UO_763 (O_763,N_19651,N_19431);
or UO_764 (O_764,N_19448,N_19071);
or UO_765 (O_765,N_19545,N_19028);
xnor UO_766 (O_766,N_19780,N_19469);
xnor UO_767 (O_767,N_19096,N_19380);
nand UO_768 (O_768,N_19469,N_19064);
nand UO_769 (O_769,N_19963,N_19817);
xor UO_770 (O_770,N_19584,N_19595);
and UO_771 (O_771,N_19932,N_19450);
xor UO_772 (O_772,N_19924,N_19807);
nor UO_773 (O_773,N_19682,N_19186);
or UO_774 (O_774,N_19753,N_19325);
nand UO_775 (O_775,N_19129,N_19724);
and UO_776 (O_776,N_19335,N_19791);
and UO_777 (O_777,N_19161,N_19745);
or UO_778 (O_778,N_19001,N_19261);
nand UO_779 (O_779,N_19038,N_19311);
nor UO_780 (O_780,N_19318,N_19524);
nor UO_781 (O_781,N_19695,N_19236);
nor UO_782 (O_782,N_19923,N_19369);
nand UO_783 (O_783,N_19220,N_19904);
nor UO_784 (O_784,N_19948,N_19707);
or UO_785 (O_785,N_19228,N_19770);
nand UO_786 (O_786,N_19908,N_19800);
or UO_787 (O_787,N_19824,N_19435);
nand UO_788 (O_788,N_19022,N_19788);
nor UO_789 (O_789,N_19184,N_19661);
or UO_790 (O_790,N_19654,N_19072);
xor UO_791 (O_791,N_19497,N_19395);
or UO_792 (O_792,N_19152,N_19086);
and UO_793 (O_793,N_19671,N_19282);
and UO_794 (O_794,N_19369,N_19414);
and UO_795 (O_795,N_19369,N_19273);
xnor UO_796 (O_796,N_19502,N_19965);
and UO_797 (O_797,N_19345,N_19247);
xor UO_798 (O_798,N_19079,N_19253);
xnor UO_799 (O_799,N_19831,N_19051);
nand UO_800 (O_800,N_19484,N_19632);
nor UO_801 (O_801,N_19721,N_19388);
or UO_802 (O_802,N_19998,N_19198);
xor UO_803 (O_803,N_19760,N_19865);
nor UO_804 (O_804,N_19730,N_19923);
xnor UO_805 (O_805,N_19007,N_19617);
xor UO_806 (O_806,N_19318,N_19910);
and UO_807 (O_807,N_19979,N_19222);
nand UO_808 (O_808,N_19933,N_19211);
nand UO_809 (O_809,N_19794,N_19106);
nand UO_810 (O_810,N_19330,N_19877);
xnor UO_811 (O_811,N_19308,N_19372);
or UO_812 (O_812,N_19749,N_19708);
nand UO_813 (O_813,N_19337,N_19727);
nor UO_814 (O_814,N_19983,N_19754);
and UO_815 (O_815,N_19227,N_19851);
xnor UO_816 (O_816,N_19099,N_19613);
and UO_817 (O_817,N_19263,N_19807);
nor UO_818 (O_818,N_19530,N_19955);
nand UO_819 (O_819,N_19723,N_19046);
nor UO_820 (O_820,N_19641,N_19012);
or UO_821 (O_821,N_19376,N_19452);
nor UO_822 (O_822,N_19557,N_19303);
or UO_823 (O_823,N_19214,N_19812);
and UO_824 (O_824,N_19662,N_19355);
xnor UO_825 (O_825,N_19503,N_19565);
nor UO_826 (O_826,N_19522,N_19509);
xnor UO_827 (O_827,N_19739,N_19460);
or UO_828 (O_828,N_19616,N_19952);
nand UO_829 (O_829,N_19892,N_19948);
or UO_830 (O_830,N_19522,N_19503);
xor UO_831 (O_831,N_19287,N_19193);
nor UO_832 (O_832,N_19160,N_19947);
nand UO_833 (O_833,N_19555,N_19773);
and UO_834 (O_834,N_19458,N_19577);
or UO_835 (O_835,N_19941,N_19140);
xor UO_836 (O_836,N_19970,N_19603);
nor UO_837 (O_837,N_19841,N_19751);
nor UO_838 (O_838,N_19006,N_19574);
xnor UO_839 (O_839,N_19023,N_19354);
xor UO_840 (O_840,N_19573,N_19296);
or UO_841 (O_841,N_19430,N_19875);
or UO_842 (O_842,N_19326,N_19793);
nand UO_843 (O_843,N_19277,N_19639);
nand UO_844 (O_844,N_19276,N_19699);
xor UO_845 (O_845,N_19777,N_19033);
and UO_846 (O_846,N_19904,N_19289);
or UO_847 (O_847,N_19851,N_19599);
nand UO_848 (O_848,N_19823,N_19954);
or UO_849 (O_849,N_19835,N_19936);
or UO_850 (O_850,N_19630,N_19883);
nand UO_851 (O_851,N_19790,N_19016);
and UO_852 (O_852,N_19711,N_19331);
nand UO_853 (O_853,N_19914,N_19704);
and UO_854 (O_854,N_19643,N_19407);
or UO_855 (O_855,N_19679,N_19265);
or UO_856 (O_856,N_19599,N_19942);
and UO_857 (O_857,N_19219,N_19725);
or UO_858 (O_858,N_19096,N_19377);
nor UO_859 (O_859,N_19573,N_19493);
xnor UO_860 (O_860,N_19155,N_19864);
nor UO_861 (O_861,N_19398,N_19973);
or UO_862 (O_862,N_19240,N_19200);
nand UO_863 (O_863,N_19311,N_19653);
nand UO_864 (O_864,N_19125,N_19331);
and UO_865 (O_865,N_19356,N_19560);
and UO_866 (O_866,N_19203,N_19495);
and UO_867 (O_867,N_19414,N_19172);
nand UO_868 (O_868,N_19292,N_19153);
nand UO_869 (O_869,N_19149,N_19040);
nor UO_870 (O_870,N_19459,N_19209);
nand UO_871 (O_871,N_19980,N_19109);
or UO_872 (O_872,N_19007,N_19462);
and UO_873 (O_873,N_19146,N_19573);
or UO_874 (O_874,N_19611,N_19110);
and UO_875 (O_875,N_19469,N_19443);
or UO_876 (O_876,N_19884,N_19938);
nor UO_877 (O_877,N_19041,N_19218);
or UO_878 (O_878,N_19727,N_19884);
or UO_879 (O_879,N_19060,N_19320);
xnor UO_880 (O_880,N_19105,N_19592);
xnor UO_881 (O_881,N_19063,N_19467);
or UO_882 (O_882,N_19452,N_19858);
and UO_883 (O_883,N_19884,N_19413);
and UO_884 (O_884,N_19918,N_19311);
nand UO_885 (O_885,N_19367,N_19885);
and UO_886 (O_886,N_19001,N_19550);
nor UO_887 (O_887,N_19998,N_19368);
nand UO_888 (O_888,N_19199,N_19530);
and UO_889 (O_889,N_19103,N_19809);
and UO_890 (O_890,N_19528,N_19573);
nor UO_891 (O_891,N_19241,N_19202);
nand UO_892 (O_892,N_19966,N_19072);
nor UO_893 (O_893,N_19812,N_19901);
and UO_894 (O_894,N_19844,N_19719);
nand UO_895 (O_895,N_19819,N_19844);
xor UO_896 (O_896,N_19390,N_19371);
nor UO_897 (O_897,N_19187,N_19868);
and UO_898 (O_898,N_19545,N_19903);
or UO_899 (O_899,N_19681,N_19783);
or UO_900 (O_900,N_19781,N_19193);
and UO_901 (O_901,N_19978,N_19221);
nand UO_902 (O_902,N_19346,N_19802);
or UO_903 (O_903,N_19804,N_19794);
nand UO_904 (O_904,N_19791,N_19312);
or UO_905 (O_905,N_19053,N_19645);
nand UO_906 (O_906,N_19834,N_19949);
nand UO_907 (O_907,N_19888,N_19666);
nand UO_908 (O_908,N_19387,N_19370);
or UO_909 (O_909,N_19365,N_19996);
and UO_910 (O_910,N_19949,N_19890);
nor UO_911 (O_911,N_19538,N_19542);
nand UO_912 (O_912,N_19066,N_19417);
nand UO_913 (O_913,N_19490,N_19726);
or UO_914 (O_914,N_19714,N_19637);
xor UO_915 (O_915,N_19855,N_19078);
and UO_916 (O_916,N_19157,N_19798);
nor UO_917 (O_917,N_19672,N_19362);
nor UO_918 (O_918,N_19120,N_19435);
nor UO_919 (O_919,N_19990,N_19102);
xor UO_920 (O_920,N_19729,N_19891);
xor UO_921 (O_921,N_19190,N_19324);
nor UO_922 (O_922,N_19931,N_19075);
nand UO_923 (O_923,N_19286,N_19528);
xor UO_924 (O_924,N_19067,N_19162);
nor UO_925 (O_925,N_19554,N_19402);
or UO_926 (O_926,N_19444,N_19332);
xnor UO_927 (O_927,N_19854,N_19676);
nand UO_928 (O_928,N_19490,N_19733);
and UO_929 (O_929,N_19520,N_19651);
nor UO_930 (O_930,N_19896,N_19307);
or UO_931 (O_931,N_19826,N_19017);
and UO_932 (O_932,N_19376,N_19306);
nand UO_933 (O_933,N_19058,N_19552);
and UO_934 (O_934,N_19912,N_19764);
or UO_935 (O_935,N_19071,N_19383);
nor UO_936 (O_936,N_19163,N_19413);
nand UO_937 (O_937,N_19958,N_19391);
and UO_938 (O_938,N_19520,N_19750);
nor UO_939 (O_939,N_19817,N_19387);
xor UO_940 (O_940,N_19209,N_19278);
nor UO_941 (O_941,N_19832,N_19292);
or UO_942 (O_942,N_19890,N_19344);
xor UO_943 (O_943,N_19506,N_19563);
nand UO_944 (O_944,N_19871,N_19527);
or UO_945 (O_945,N_19766,N_19814);
xnor UO_946 (O_946,N_19482,N_19806);
or UO_947 (O_947,N_19317,N_19261);
xor UO_948 (O_948,N_19679,N_19706);
and UO_949 (O_949,N_19525,N_19110);
xor UO_950 (O_950,N_19008,N_19268);
or UO_951 (O_951,N_19058,N_19127);
or UO_952 (O_952,N_19768,N_19681);
nor UO_953 (O_953,N_19409,N_19606);
or UO_954 (O_954,N_19886,N_19225);
nor UO_955 (O_955,N_19217,N_19866);
or UO_956 (O_956,N_19404,N_19462);
and UO_957 (O_957,N_19317,N_19838);
xnor UO_958 (O_958,N_19721,N_19252);
nand UO_959 (O_959,N_19745,N_19223);
and UO_960 (O_960,N_19906,N_19404);
nand UO_961 (O_961,N_19730,N_19564);
nand UO_962 (O_962,N_19772,N_19403);
xnor UO_963 (O_963,N_19854,N_19201);
nor UO_964 (O_964,N_19247,N_19755);
nand UO_965 (O_965,N_19417,N_19723);
and UO_966 (O_966,N_19719,N_19946);
or UO_967 (O_967,N_19656,N_19962);
or UO_968 (O_968,N_19850,N_19421);
nor UO_969 (O_969,N_19397,N_19030);
and UO_970 (O_970,N_19964,N_19196);
nand UO_971 (O_971,N_19352,N_19799);
xnor UO_972 (O_972,N_19613,N_19491);
or UO_973 (O_973,N_19613,N_19746);
or UO_974 (O_974,N_19290,N_19709);
xnor UO_975 (O_975,N_19291,N_19173);
nor UO_976 (O_976,N_19731,N_19344);
or UO_977 (O_977,N_19581,N_19115);
nor UO_978 (O_978,N_19135,N_19410);
or UO_979 (O_979,N_19123,N_19818);
nand UO_980 (O_980,N_19516,N_19166);
or UO_981 (O_981,N_19441,N_19479);
xnor UO_982 (O_982,N_19672,N_19355);
nor UO_983 (O_983,N_19027,N_19387);
or UO_984 (O_984,N_19326,N_19916);
and UO_985 (O_985,N_19372,N_19936);
nand UO_986 (O_986,N_19584,N_19898);
xor UO_987 (O_987,N_19116,N_19182);
xnor UO_988 (O_988,N_19385,N_19327);
and UO_989 (O_989,N_19960,N_19386);
and UO_990 (O_990,N_19016,N_19413);
xnor UO_991 (O_991,N_19132,N_19223);
and UO_992 (O_992,N_19687,N_19146);
nand UO_993 (O_993,N_19509,N_19279);
nor UO_994 (O_994,N_19699,N_19339);
nor UO_995 (O_995,N_19007,N_19746);
and UO_996 (O_996,N_19053,N_19203);
or UO_997 (O_997,N_19199,N_19283);
xnor UO_998 (O_998,N_19529,N_19100);
nand UO_999 (O_999,N_19967,N_19577);
or UO_1000 (O_1000,N_19084,N_19276);
xnor UO_1001 (O_1001,N_19207,N_19105);
nand UO_1002 (O_1002,N_19653,N_19480);
or UO_1003 (O_1003,N_19713,N_19149);
or UO_1004 (O_1004,N_19868,N_19601);
or UO_1005 (O_1005,N_19344,N_19604);
nand UO_1006 (O_1006,N_19197,N_19207);
or UO_1007 (O_1007,N_19489,N_19894);
or UO_1008 (O_1008,N_19745,N_19117);
nand UO_1009 (O_1009,N_19106,N_19499);
or UO_1010 (O_1010,N_19894,N_19239);
xor UO_1011 (O_1011,N_19484,N_19076);
nand UO_1012 (O_1012,N_19846,N_19449);
nand UO_1013 (O_1013,N_19021,N_19138);
nor UO_1014 (O_1014,N_19188,N_19032);
nor UO_1015 (O_1015,N_19029,N_19631);
nand UO_1016 (O_1016,N_19204,N_19094);
nor UO_1017 (O_1017,N_19429,N_19820);
and UO_1018 (O_1018,N_19118,N_19805);
or UO_1019 (O_1019,N_19627,N_19630);
nand UO_1020 (O_1020,N_19999,N_19819);
nand UO_1021 (O_1021,N_19120,N_19238);
nand UO_1022 (O_1022,N_19041,N_19158);
or UO_1023 (O_1023,N_19158,N_19600);
nor UO_1024 (O_1024,N_19813,N_19900);
nand UO_1025 (O_1025,N_19634,N_19520);
nand UO_1026 (O_1026,N_19489,N_19432);
xor UO_1027 (O_1027,N_19003,N_19370);
xor UO_1028 (O_1028,N_19889,N_19978);
nor UO_1029 (O_1029,N_19414,N_19841);
nor UO_1030 (O_1030,N_19516,N_19485);
nand UO_1031 (O_1031,N_19606,N_19591);
and UO_1032 (O_1032,N_19185,N_19179);
xnor UO_1033 (O_1033,N_19244,N_19210);
or UO_1034 (O_1034,N_19721,N_19297);
and UO_1035 (O_1035,N_19654,N_19880);
xor UO_1036 (O_1036,N_19973,N_19551);
or UO_1037 (O_1037,N_19785,N_19646);
or UO_1038 (O_1038,N_19547,N_19676);
or UO_1039 (O_1039,N_19349,N_19299);
or UO_1040 (O_1040,N_19316,N_19457);
and UO_1041 (O_1041,N_19029,N_19080);
xor UO_1042 (O_1042,N_19065,N_19723);
and UO_1043 (O_1043,N_19629,N_19015);
nor UO_1044 (O_1044,N_19750,N_19805);
and UO_1045 (O_1045,N_19585,N_19170);
or UO_1046 (O_1046,N_19407,N_19923);
and UO_1047 (O_1047,N_19355,N_19490);
nand UO_1048 (O_1048,N_19787,N_19149);
nor UO_1049 (O_1049,N_19620,N_19036);
nor UO_1050 (O_1050,N_19310,N_19891);
nor UO_1051 (O_1051,N_19982,N_19864);
or UO_1052 (O_1052,N_19633,N_19867);
xnor UO_1053 (O_1053,N_19564,N_19036);
nand UO_1054 (O_1054,N_19317,N_19939);
nand UO_1055 (O_1055,N_19514,N_19698);
xor UO_1056 (O_1056,N_19949,N_19217);
xnor UO_1057 (O_1057,N_19104,N_19102);
nand UO_1058 (O_1058,N_19738,N_19155);
and UO_1059 (O_1059,N_19305,N_19831);
xor UO_1060 (O_1060,N_19603,N_19501);
nand UO_1061 (O_1061,N_19973,N_19501);
nand UO_1062 (O_1062,N_19027,N_19277);
xor UO_1063 (O_1063,N_19752,N_19409);
xnor UO_1064 (O_1064,N_19535,N_19936);
or UO_1065 (O_1065,N_19656,N_19948);
xor UO_1066 (O_1066,N_19805,N_19516);
or UO_1067 (O_1067,N_19138,N_19135);
and UO_1068 (O_1068,N_19692,N_19975);
and UO_1069 (O_1069,N_19043,N_19639);
nor UO_1070 (O_1070,N_19014,N_19499);
or UO_1071 (O_1071,N_19979,N_19796);
or UO_1072 (O_1072,N_19543,N_19005);
nand UO_1073 (O_1073,N_19559,N_19220);
nand UO_1074 (O_1074,N_19136,N_19348);
xor UO_1075 (O_1075,N_19414,N_19283);
and UO_1076 (O_1076,N_19390,N_19480);
and UO_1077 (O_1077,N_19426,N_19117);
nor UO_1078 (O_1078,N_19703,N_19568);
xnor UO_1079 (O_1079,N_19974,N_19748);
nand UO_1080 (O_1080,N_19740,N_19340);
xor UO_1081 (O_1081,N_19154,N_19432);
nand UO_1082 (O_1082,N_19406,N_19906);
or UO_1083 (O_1083,N_19650,N_19938);
nor UO_1084 (O_1084,N_19812,N_19534);
nand UO_1085 (O_1085,N_19391,N_19401);
xor UO_1086 (O_1086,N_19500,N_19411);
and UO_1087 (O_1087,N_19982,N_19516);
or UO_1088 (O_1088,N_19918,N_19960);
xor UO_1089 (O_1089,N_19255,N_19636);
and UO_1090 (O_1090,N_19415,N_19852);
xnor UO_1091 (O_1091,N_19851,N_19385);
nor UO_1092 (O_1092,N_19766,N_19978);
and UO_1093 (O_1093,N_19179,N_19218);
nand UO_1094 (O_1094,N_19399,N_19255);
xnor UO_1095 (O_1095,N_19010,N_19893);
nand UO_1096 (O_1096,N_19860,N_19731);
and UO_1097 (O_1097,N_19361,N_19952);
and UO_1098 (O_1098,N_19857,N_19771);
and UO_1099 (O_1099,N_19983,N_19304);
xnor UO_1100 (O_1100,N_19283,N_19528);
nand UO_1101 (O_1101,N_19701,N_19310);
nand UO_1102 (O_1102,N_19655,N_19921);
xnor UO_1103 (O_1103,N_19439,N_19913);
nand UO_1104 (O_1104,N_19707,N_19030);
xor UO_1105 (O_1105,N_19285,N_19031);
or UO_1106 (O_1106,N_19927,N_19623);
and UO_1107 (O_1107,N_19773,N_19202);
xor UO_1108 (O_1108,N_19057,N_19909);
or UO_1109 (O_1109,N_19005,N_19434);
nand UO_1110 (O_1110,N_19178,N_19296);
nor UO_1111 (O_1111,N_19111,N_19494);
or UO_1112 (O_1112,N_19365,N_19849);
or UO_1113 (O_1113,N_19906,N_19737);
and UO_1114 (O_1114,N_19595,N_19816);
and UO_1115 (O_1115,N_19007,N_19594);
nand UO_1116 (O_1116,N_19705,N_19829);
xor UO_1117 (O_1117,N_19953,N_19844);
xor UO_1118 (O_1118,N_19452,N_19793);
nand UO_1119 (O_1119,N_19628,N_19895);
xor UO_1120 (O_1120,N_19422,N_19989);
xnor UO_1121 (O_1121,N_19497,N_19590);
nor UO_1122 (O_1122,N_19197,N_19060);
or UO_1123 (O_1123,N_19805,N_19194);
and UO_1124 (O_1124,N_19073,N_19326);
or UO_1125 (O_1125,N_19088,N_19920);
xnor UO_1126 (O_1126,N_19883,N_19318);
or UO_1127 (O_1127,N_19826,N_19752);
and UO_1128 (O_1128,N_19745,N_19087);
nand UO_1129 (O_1129,N_19243,N_19343);
xor UO_1130 (O_1130,N_19670,N_19669);
nor UO_1131 (O_1131,N_19024,N_19109);
nor UO_1132 (O_1132,N_19859,N_19057);
xnor UO_1133 (O_1133,N_19612,N_19346);
xor UO_1134 (O_1134,N_19252,N_19959);
xnor UO_1135 (O_1135,N_19741,N_19099);
or UO_1136 (O_1136,N_19040,N_19350);
nand UO_1137 (O_1137,N_19089,N_19814);
nand UO_1138 (O_1138,N_19315,N_19021);
xnor UO_1139 (O_1139,N_19181,N_19243);
nor UO_1140 (O_1140,N_19894,N_19393);
xor UO_1141 (O_1141,N_19942,N_19323);
xnor UO_1142 (O_1142,N_19362,N_19714);
and UO_1143 (O_1143,N_19592,N_19318);
or UO_1144 (O_1144,N_19819,N_19535);
and UO_1145 (O_1145,N_19133,N_19418);
and UO_1146 (O_1146,N_19299,N_19140);
nand UO_1147 (O_1147,N_19598,N_19661);
nor UO_1148 (O_1148,N_19425,N_19421);
nand UO_1149 (O_1149,N_19223,N_19267);
and UO_1150 (O_1150,N_19581,N_19802);
or UO_1151 (O_1151,N_19772,N_19445);
nor UO_1152 (O_1152,N_19790,N_19734);
or UO_1153 (O_1153,N_19725,N_19665);
nor UO_1154 (O_1154,N_19726,N_19921);
or UO_1155 (O_1155,N_19163,N_19013);
and UO_1156 (O_1156,N_19184,N_19980);
or UO_1157 (O_1157,N_19290,N_19317);
nand UO_1158 (O_1158,N_19851,N_19993);
and UO_1159 (O_1159,N_19726,N_19026);
or UO_1160 (O_1160,N_19856,N_19360);
or UO_1161 (O_1161,N_19628,N_19665);
nor UO_1162 (O_1162,N_19364,N_19940);
nor UO_1163 (O_1163,N_19441,N_19661);
or UO_1164 (O_1164,N_19214,N_19772);
nor UO_1165 (O_1165,N_19667,N_19305);
or UO_1166 (O_1166,N_19345,N_19492);
nand UO_1167 (O_1167,N_19004,N_19193);
nand UO_1168 (O_1168,N_19037,N_19361);
nand UO_1169 (O_1169,N_19427,N_19455);
xnor UO_1170 (O_1170,N_19970,N_19382);
nor UO_1171 (O_1171,N_19345,N_19125);
nor UO_1172 (O_1172,N_19582,N_19715);
nand UO_1173 (O_1173,N_19692,N_19869);
nor UO_1174 (O_1174,N_19117,N_19535);
nor UO_1175 (O_1175,N_19636,N_19031);
and UO_1176 (O_1176,N_19836,N_19736);
xnor UO_1177 (O_1177,N_19769,N_19652);
nor UO_1178 (O_1178,N_19358,N_19169);
or UO_1179 (O_1179,N_19197,N_19369);
or UO_1180 (O_1180,N_19640,N_19727);
xor UO_1181 (O_1181,N_19472,N_19929);
nand UO_1182 (O_1182,N_19539,N_19354);
or UO_1183 (O_1183,N_19029,N_19340);
nor UO_1184 (O_1184,N_19551,N_19614);
or UO_1185 (O_1185,N_19555,N_19505);
or UO_1186 (O_1186,N_19654,N_19260);
or UO_1187 (O_1187,N_19050,N_19751);
xnor UO_1188 (O_1188,N_19333,N_19053);
or UO_1189 (O_1189,N_19020,N_19631);
xor UO_1190 (O_1190,N_19960,N_19119);
nand UO_1191 (O_1191,N_19987,N_19249);
or UO_1192 (O_1192,N_19859,N_19287);
or UO_1193 (O_1193,N_19677,N_19069);
or UO_1194 (O_1194,N_19893,N_19124);
or UO_1195 (O_1195,N_19960,N_19742);
xnor UO_1196 (O_1196,N_19696,N_19587);
or UO_1197 (O_1197,N_19267,N_19403);
and UO_1198 (O_1198,N_19252,N_19633);
nor UO_1199 (O_1199,N_19430,N_19364);
and UO_1200 (O_1200,N_19119,N_19685);
nor UO_1201 (O_1201,N_19579,N_19504);
xnor UO_1202 (O_1202,N_19126,N_19295);
nand UO_1203 (O_1203,N_19685,N_19282);
and UO_1204 (O_1204,N_19818,N_19163);
and UO_1205 (O_1205,N_19354,N_19197);
xor UO_1206 (O_1206,N_19409,N_19848);
or UO_1207 (O_1207,N_19884,N_19675);
and UO_1208 (O_1208,N_19221,N_19507);
nor UO_1209 (O_1209,N_19739,N_19490);
xor UO_1210 (O_1210,N_19833,N_19623);
xnor UO_1211 (O_1211,N_19388,N_19897);
nor UO_1212 (O_1212,N_19090,N_19265);
or UO_1213 (O_1213,N_19783,N_19657);
nand UO_1214 (O_1214,N_19979,N_19803);
and UO_1215 (O_1215,N_19224,N_19653);
nand UO_1216 (O_1216,N_19371,N_19171);
or UO_1217 (O_1217,N_19918,N_19997);
and UO_1218 (O_1218,N_19008,N_19963);
and UO_1219 (O_1219,N_19411,N_19006);
and UO_1220 (O_1220,N_19798,N_19615);
xnor UO_1221 (O_1221,N_19981,N_19660);
and UO_1222 (O_1222,N_19544,N_19180);
xnor UO_1223 (O_1223,N_19886,N_19294);
xor UO_1224 (O_1224,N_19536,N_19114);
nor UO_1225 (O_1225,N_19053,N_19636);
xor UO_1226 (O_1226,N_19585,N_19951);
nand UO_1227 (O_1227,N_19099,N_19084);
or UO_1228 (O_1228,N_19506,N_19768);
or UO_1229 (O_1229,N_19079,N_19891);
xnor UO_1230 (O_1230,N_19588,N_19632);
nor UO_1231 (O_1231,N_19090,N_19936);
and UO_1232 (O_1232,N_19836,N_19603);
nor UO_1233 (O_1233,N_19210,N_19635);
or UO_1234 (O_1234,N_19275,N_19709);
nor UO_1235 (O_1235,N_19241,N_19328);
nor UO_1236 (O_1236,N_19289,N_19927);
nand UO_1237 (O_1237,N_19760,N_19196);
and UO_1238 (O_1238,N_19411,N_19746);
nand UO_1239 (O_1239,N_19946,N_19746);
nor UO_1240 (O_1240,N_19470,N_19643);
nand UO_1241 (O_1241,N_19219,N_19737);
and UO_1242 (O_1242,N_19864,N_19310);
and UO_1243 (O_1243,N_19226,N_19978);
and UO_1244 (O_1244,N_19526,N_19793);
or UO_1245 (O_1245,N_19302,N_19097);
nor UO_1246 (O_1246,N_19646,N_19276);
or UO_1247 (O_1247,N_19506,N_19496);
or UO_1248 (O_1248,N_19676,N_19224);
or UO_1249 (O_1249,N_19212,N_19057);
or UO_1250 (O_1250,N_19625,N_19796);
xnor UO_1251 (O_1251,N_19166,N_19854);
and UO_1252 (O_1252,N_19587,N_19642);
or UO_1253 (O_1253,N_19214,N_19337);
or UO_1254 (O_1254,N_19703,N_19771);
xor UO_1255 (O_1255,N_19608,N_19031);
xnor UO_1256 (O_1256,N_19633,N_19421);
nand UO_1257 (O_1257,N_19682,N_19648);
nor UO_1258 (O_1258,N_19268,N_19699);
and UO_1259 (O_1259,N_19867,N_19868);
nand UO_1260 (O_1260,N_19616,N_19682);
nand UO_1261 (O_1261,N_19878,N_19034);
xnor UO_1262 (O_1262,N_19166,N_19236);
nand UO_1263 (O_1263,N_19674,N_19013);
nand UO_1264 (O_1264,N_19412,N_19691);
or UO_1265 (O_1265,N_19218,N_19811);
xnor UO_1266 (O_1266,N_19571,N_19552);
nand UO_1267 (O_1267,N_19040,N_19640);
nor UO_1268 (O_1268,N_19099,N_19985);
nor UO_1269 (O_1269,N_19057,N_19221);
nand UO_1270 (O_1270,N_19938,N_19507);
xnor UO_1271 (O_1271,N_19848,N_19488);
or UO_1272 (O_1272,N_19650,N_19289);
nor UO_1273 (O_1273,N_19679,N_19983);
and UO_1274 (O_1274,N_19551,N_19088);
and UO_1275 (O_1275,N_19084,N_19634);
and UO_1276 (O_1276,N_19850,N_19689);
or UO_1277 (O_1277,N_19663,N_19757);
or UO_1278 (O_1278,N_19498,N_19875);
and UO_1279 (O_1279,N_19232,N_19173);
nand UO_1280 (O_1280,N_19666,N_19026);
or UO_1281 (O_1281,N_19820,N_19806);
and UO_1282 (O_1282,N_19518,N_19656);
xnor UO_1283 (O_1283,N_19181,N_19396);
nand UO_1284 (O_1284,N_19544,N_19252);
nor UO_1285 (O_1285,N_19775,N_19314);
nor UO_1286 (O_1286,N_19463,N_19174);
xor UO_1287 (O_1287,N_19465,N_19248);
xor UO_1288 (O_1288,N_19259,N_19463);
xor UO_1289 (O_1289,N_19159,N_19279);
or UO_1290 (O_1290,N_19986,N_19168);
or UO_1291 (O_1291,N_19622,N_19448);
nor UO_1292 (O_1292,N_19394,N_19030);
xor UO_1293 (O_1293,N_19566,N_19183);
nor UO_1294 (O_1294,N_19635,N_19023);
xnor UO_1295 (O_1295,N_19186,N_19092);
and UO_1296 (O_1296,N_19842,N_19706);
nand UO_1297 (O_1297,N_19257,N_19271);
and UO_1298 (O_1298,N_19542,N_19061);
or UO_1299 (O_1299,N_19984,N_19109);
nand UO_1300 (O_1300,N_19016,N_19859);
nor UO_1301 (O_1301,N_19197,N_19849);
and UO_1302 (O_1302,N_19114,N_19378);
and UO_1303 (O_1303,N_19352,N_19912);
or UO_1304 (O_1304,N_19709,N_19702);
nor UO_1305 (O_1305,N_19866,N_19358);
nor UO_1306 (O_1306,N_19138,N_19821);
nor UO_1307 (O_1307,N_19606,N_19414);
and UO_1308 (O_1308,N_19206,N_19018);
xnor UO_1309 (O_1309,N_19182,N_19552);
or UO_1310 (O_1310,N_19968,N_19375);
xnor UO_1311 (O_1311,N_19709,N_19838);
nor UO_1312 (O_1312,N_19360,N_19813);
nand UO_1313 (O_1313,N_19982,N_19506);
or UO_1314 (O_1314,N_19818,N_19312);
nor UO_1315 (O_1315,N_19771,N_19003);
xnor UO_1316 (O_1316,N_19022,N_19814);
nor UO_1317 (O_1317,N_19226,N_19544);
xor UO_1318 (O_1318,N_19387,N_19593);
nand UO_1319 (O_1319,N_19787,N_19052);
xor UO_1320 (O_1320,N_19727,N_19892);
and UO_1321 (O_1321,N_19932,N_19895);
xor UO_1322 (O_1322,N_19360,N_19047);
nand UO_1323 (O_1323,N_19372,N_19852);
nor UO_1324 (O_1324,N_19971,N_19342);
nor UO_1325 (O_1325,N_19505,N_19188);
xnor UO_1326 (O_1326,N_19520,N_19257);
nor UO_1327 (O_1327,N_19886,N_19743);
nor UO_1328 (O_1328,N_19352,N_19939);
xor UO_1329 (O_1329,N_19183,N_19956);
nand UO_1330 (O_1330,N_19272,N_19122);
xnor UO_1331 (O_1331,N_19236,N_19944);
xnor UO_1332 (O_1332,N_19817,N_19684);
and UO_1333 (O_1333,N_19179,N_19234);
xnor UO_1334 (O_1334,N_19801,N_19355);
and UO_1335 (O_1335,N_19103,N_19486);
and UO_1336 (O_1336,N_19133,N_19429);
xnor UO_1337 (O_1337,N_19792,N_19100);
nand UO_1338 (O_1338,N_19532,N_19859);
nor UO_1339 (O_1339,N_19562,N_19609);
or UO_1340 (O_1340,N_19005,N_19583);
xnor UO_1341 (O_1341,N_19012,N_19550);
or UO_1342 (O_1342,N_19452,N_19785);
nor UO_1343 (O_1343,N_19787,N_19561);
xnor UO_1344 (O_1344,N_19871,N_19496);
or UO_1345 (O_1345,N_19652,N_19566);
nor UO_1346 (O_1346,N_19766,N_19049);
xnor UO_1347 (O_1347,N_19824,N_19903);
nand UO_1348 (O_1348,N_19398,N_19423);
nor UO_1349 (O_1349,N_19421,N_19436);
nand UO_1350 (O_1350,N_19160,N_19033);
xor UO_1351 (O_1351,N_19137,N_19890);
xnor UO_1352 (O_1352,N_19257,N_19404);
and UO_1353 (O_1353,N_19801,N_19455);
nand UO_1354 (O_1354,N_19540,N_19329);
xnor UO_1355 (O_1355,N_19468,N_19547);
and UO_1356 (O_1356,N_19791,N_19114);
nor UO_1357 (O_1357,N_19821,N_19656);
or UO_1358 (O_1358,N_19295,N_19144);
or UO_1359 (O_1359,N_19650,N_19648);
nor UO_1360 (O_1360,N_19079,N_19658);
xor UO_1361 (O_1361,N_19331,N_19090);
and UO_1362 (O_1362,N_19693,N_19072);
or UO_1363 (O_1363,N_19129,N_19998);
nor UO_1364 (O_1364,N_19682,N_19094);
and UO_1365 (O_1365,N_19205,N_19080);
nor UO_1366 (O_1366,N_19168,N_19542);
nor UO_1367 (O_1367,N_19737,N_19070);
xor UO_1368 (O_1368,N_19539,N_19533);
nand UO_1369 (O_1369,N_19952,N_19437);
and UO_1370 (O_1370,N_19979,N_19350);
or UO_1371 (O_1371,N_19135,N_19133);
and UO_1372 (O_1372,N_19974,N_19328);
nor UO_1373 (O_1373,N_19988,N_19245);
and UO_1374 (O_1374,N_19175,N_19778);
and UO_1375 (O_1375,N_19309,N_19933);
and UO_1376 (O_1376,N_19044,N_19247);
or UO_1377 (O_1377,N_19209,N_19010);
nor UO_1378 (O_1378,N_19295,N_19296);
xnor UO_1379 (O_1379,N_19032,N_19688);
or UO_1380 (O_1380,N_19922,N_19889);
or UO_1381 (O_1381,N_19291,N_19044);
xnor UO_1382 (O_1382,N_19728,N_19032);
xor UO_1383 (O_1383,N_19641,N_19060);
nand UO_1384 (O_1384,N_19551,N_19595);
xnor UO_1385 (O_1385,N_19124,N_19676);
or UO_1386 (O_1386,N_19714,N_19835);
nand UO_1387 (O_1387,N_19986,N_19274);
xnor UO_1388 (O_1388,N_19549,N_19453);
or UO_1389 (O_1389,N_19644,N_19990);
or UO_1390 (O_1390,N_19790,N_19179);
and UO_1391 (O_1391,N_19846,N_19476);
nor UO_1392 (O_1392,N_19592,N_19748);
and UO_1393 (O_1393,N_19043,N_19366);
nand UO_1394 (O_1394,N_19032,N_19192);
or UO_1395 (O_1395,N_19060,N_19339);
nand UO_1396 (O_1396,N_19686,N_19640);
nor UO_1397 (O_1397,N_19662,N_19745);
nor UO_1398 (O_1398,N_19334,N_19946);
nor UO_1399 (O_1399,N_19473,N_19158);
nor UO_1400 (O_1400,N_19879,N_19594);
nand UO_1401 (O_1401,N_19337,N_19471);
xnor UO_1402 (O_1402,N_19869,N_19663);
nor UO_1403 (O_1403,N_19037,N_19717);
nand UO_1404 (O_1404,N_19122,N_19986);
xor UO_1405 (O_1405,N_19781,N_19115);
nor UO_1406 (O_1406,N_19520,N_19305);
nor UO_1407 (O_1407,N_19960,N_19431);
and UO_1408 (O_1408,N_19043,N_19243);
nor UO_1409 (O_1409,N_19573,N_19866);
nand UO_1410 (O_1410,N_19291,N_19607);
nor UO_1411 (O_1411,N_19811,N_19956);
and UO_1412 (O_1412,N_19744,N_19205);
or UO_1413 (O_1413,N_19541,N_19866);
nor UO_1414 (O_1414,N_19075,N_19612);
nor UO_1415 (O_1415,N_19994,N_19903);
nand UO_1416 (O_1416,N_19086,N_19718);
and UO_1417 (O_1417,N_19923,N_19832);
and UO_1418 (O_1418,N_19294,N_19408);
and UO_1419 (O_1419,N_19070,N_19263);
nand UO_1420 (O_1420,N_19564,N_19586);
and UO_1421 (O_1421,N_19107,N_19523);
and UO_1422 (O_1422,N_19015,N_19122);
nor UO_1423 (O_1423,N_19930,N_19592);
and UO_1424 (O_1424,N_19680,N_19783);
nand UO_1425 (O_1425,N_19040,N_19688);
nor UO_1426 (O_1426,N_19352,N_19843);
nand UO_1427 (O_1427,N_19864,N_19819);
and UO_1428 (O_1428,N_19110,N_19780);
xor UO_1429 (O_1429,N_19453,N_19391);
nand UO_1430 (O_1430,N_19513,N_19020);
nand UO_1431 (O_1431,N_19888,N_19760);
nand UO_1432 (O_1432,N_19451,N_19672);
nand UO_1433 (O_1433,N_19678,N_19094);
and UO_1434 (O_1434,N_19884,N_19610);
nand UO_1435 (O_1435,N_19081,N_19279);
xnor UO_1436 (O_1436,N_19934,N_19773);
or UO_1437 (O_1437,N_19790,N_19986);
and UO_1438 (O_1438,N_19443,N_19312);
and UO_1439 (O_1439,N_19555,N_19352);
xnor UO_1440 (O_1440,N_19372,N_19119);
xor UO_1441 (O_1441,N_19019,N_19003);
nand UO_1442 (O_1442,N_19007,N_19792);
nand UO_1443 (O_1443,N_19832,N_19273);
and UO_1444 (O_1444,N_19069,N_19984);
and UO_1445 (O_1445,N_19525,N_19299);
xnor UO_1446 (O_1446,N_19381,N_19233);
and UO_1447 (O_1447,N_19944,N_19307);
xor UO_1448 (O_1448,N_19418,N_19248);
nor UO_1449 (O_1449,N_19914,N_19437);
or UO_1450 (O_1450,N_19677,N_19872);
or UO_1451 (O_1451,N_19338,N_19749);
nand UO_1452 (O_1452,N_19098,N_19107);
and UO_1453 (O_1453,N_19633,N_19119);
and UO_1454 (O_1454,N_19907,N_19999);
nand UO_1455 (O_1455,N_19502,N_19339);
nand UO_1456 (O_1456,N_19252,N_19290);
and UO_1457 (O_1457,N_19701,N_19476);
nand UO_1458 (O_1458,N_19129,N_19147);
and UO_1459 (O_1459,N_19545,N_19128);
nor UO_1460 (O_1460,N_19863,N_19245);
or UO_1461 (O_1461,N_19935,N_19283);
nand UO_1462 (O_1462,N_19175,N_19566);
xor UO_1463 (O_1463,N_19856,N_19404);
nor UO_1464 (O_1464,N_19830,N_19890);
or UO_1465 (O_1465,N_19362,N_19058);
nand UO_1466 (O_1466,N_19569,N_19592);
nand UO_1467 (O_1467,N_19072,N_19188);
or UO_1468 (O_1468,N_19677,N_19339);
xnor UO_1469 (O_1469,N_19177,N_19234);
and UO_1470 (O_1470,N_19792,N_19150);
xnor UO_1471 (O_1471,N_19337,N_19966);
nor UO_1472 (O_1472,N_19285,N_19568);
xnor UO_1473 (O_1473,N_19680,N_19366);
and UO_1474 (O_1474,N_19782,N_19055);
nor UO_1475 (O_1475,N_19005,N_19689);
and UO_1476 (O_1476,N_19262,N_19035);
xor UO_1477 (O_1477,N_19605,N_19266);
nor UO_1478 (O_1478,N_19460,N_19977);
and UO_1479 (O_1479,N_19449,N_19412);
or UO_1480 (O_1480,N_19434,N_19138);
nand UO_1481 (O_1481,N_19835,N_19851);
xor UO_1482 (O_1482,N_19927,N_19823);
and UO_1483 (O_1483,N_19688,N_19375);
xor UO_1484 (O_1484,N_19965,N_19897);
nand UO_1485 (O_1485,N_19116,N_19436);
or UO_1486 (O_1486,N_19975,N_19721);
nand UO_1487 (O_1487,N_19230,N_19973);
nand UO_1488 (O_1488,N_19174,N_19699);
nor UO_1489 (O_1489,N_19522,N_19446);
nor UO_1490 (O_1490,N_19981,N_19067);
and UO_1491 (O_1491,N_19154,N_19082);
and UO_1492 (O_1492,N_19443,N_19602);
or UO_1493 (O_1493,N_19607,N_19494);
and UO_1494 (O_1494,N_19676,N_19435);
nand UO_1495 (O_1495,N_19561,N_19919);
xnor UO_1496 (O_1496,N_19285,N_19583);
nand UO_1497 (O_1497,N_19553,N_19407);
or UO_1498 (O_1498,N_19240,N_19208);
and UO_1499 (O_1499,N_19355,N_19471);
nand UO_1500 (O_1500,N_19652,N_19656);
nor UO_1501 (O_1501,N_19998,N_19880);
nor UO_1502 (O_1502,N_19100,N_19365);
or UO_1503 (O_1503,N_19042,N_19598);
nor UO_1504 (O_1504,N_19079,N_19504);
nand UO_1505 (O_1505,N_19711,N_19316);
nand UO_1506 (O_1506,N_19233,N_19049);
or UO_1507 (O_1507,N_19330,N_19436);
xor UO_1508 (O_1508,N_19437,N_19045);
xor UO_1509 (O_1509,N_19893,N_19298);
nor UO_1510 (O_1510,N_19997,N_19060);
nand UO_1511 (O_1511,N_19718,N_19372);
nor UO_1512 (O_1512,N_19717,N_19355);
and UO_1513 (O_1513,N_19211,N_19389);
xnor UO_1514 (O_1514,N_19887,N_19874);
nand UO_1515 (O_1515,N_19590,N_19406);
nor UO_1516 (O_1516,N_19268,N_19918);
nand UO_1517 (O_1517,N_19607,N_19589);
and UO_1518 (O_1518,N_19310,N_19810);
nor UO_1519 (O_1519,N_19576,N_19138);
xnor UO_1520 (O_1520,N_19832,N_19618);
xor UO_1521 (O_1521,N_19815,N_19254);
xor UO_1522 (O_1522,N_19554,N_19809);
or UO_1523 (O_1523,N_19557,N_19428);
nand UO_1524 (O_1524,N_19666,N_19743);
or UO_1525 (O_1525,N_19861,N_19124);
nand UO_1526 (O_1526,N_19836,N_19372);
nor UO_1527 (O_1527,N_19293,N_19192);
and UO_1528 (O_1528,N_19095,N_19914);
and UO_1529 (O_1529,N_19240,N_19858);
and UO_1530 (O_1530,N_19155,N_19825);
or UO_1531 (O_1531,N_19170,N_19901);
and UO_1532 (O_1532,N_19449,N_19193);
xnor UO_1533 (O_1533,N_19272,N_19005);
nor UO_1534 (O_1534,N_19977,N_19758);
xnor UO_1535 (O_1535,N_19787,N_19847);
xor UO_1536 (O_1536,N_19720,N_19976);
and UO_1537 (O_1537,N_19465,N_19479);
nand UO_1538 (O_1538,N_19868,N_19188);
nand UO_1539 (O_1539,N_19291,N_19557);
nand UO_1540 (O_1540,N_19984,N_19569);
or UO_1541 (O_1541,N_19053,N_19672);
nor UO_1542 (O_1542,N_19795,N_19490);
xor UO_1543 (O_1543,N_19713,N_19596);
nand UO_1544 (O_1544,N_19590,N_19291);
nand UO_1545 (O_1545,N_19615,N_19924);
xnor UO_1546 (O_1546,N_19723,N_19175);
nand UO_1547 (O_1547,N_19963,N_19841);
nor UO_1548 (O_1548,N_19382,N_19524);
nor UO_1549 (O_1549,N_19068,N_19503);
or UO_1550 (O_1550,N_19822,N_19281);
and UO_1551 (O_1551,N_19731,N_19939);
xnor UO_1552 (O_1552,N_19495,N_19906);
or UO_1553 (O_1553,N_19132,N_19553);
nor UO_1554 (O_1554,N_19128,N_19743);
nand UO_1555 (O_1555,N_19042,N_19507);
nand UO_1556 (O_1556,N_19076,N_19823);
and UO_1557 (O_1557,N_19162,N_19821);
xor UO_1558 (O_1558,N_19953,N_19849);
and UO_1559 (O_1559,N_19579,N_19091);
nor UO_1560 (O_1560,N_19846,N_19751);
xnor UO_1561 (O_1561,N_19887,N_19789);
and UO_1562 (O_1562,N_19359,N_19221);
nor UO_1563 (O_1563,N_19814,N_19672);
or UO_1564 (O_1564,N_19014,N_19307);
xor UO_1565 (O_1565,N_19061,N_19081);
nor UO_1566 (O_1566,N_19821,N_19953);
nor UO_1567 (O_1567,N_19606,N_19059);
or UO_1568 (O_1568,N_19982,N_19403);
and UO_1569 (O_1569,N_19050,N_19346);
nand UO_1570 (O_1570,N_19927,N_19728);
and UO_1571 (O_1571,N_19148,N_19426);
or UO_1572 (O_1572,N_19842,N_19156);
nand UO_1573 (O_1573,N_19133,N_19699);
or UO_1574 (O_1574,N_19773,N_19311);
and UO_1575 (O_1575,N_19161,N_19503);
nor UO_1576 (O_1576,N_19353,N_19129);
or UO_1577 (O_1577,N_19045,N_19933);
and UO_1578 (O_1578,N_19594,N_19219);
nand UO_1579 (O_1579,N_19071,N_19441);
and UO_1580 (O_1580,N_19348,N_19475);
or UO_1581 (O_1581,N_19944,N_19587);
or UO_1582 (O_1582,N_19226,N_19730);
xor UO_1583 (O_1583,N_19861,N_19021);
xor UO_1584 (O_1584,N_19198,N_19495);
nand UO_1585 (O_1585,N_19937,N_19677);
nand UO_1586 (O_1586,N_19733,N_19167);
xor UO_1587 (O_1587,N_19553,N_19902);
nand UO_1588 (O_1588,N_19077,N_19208);
or UO_1589 (O_1589,N_19258,N_19456);
xor UO_1590 (O_1590,N_19379,N_19920);
nor UO_1591 (O_1591,N_19395,N_19538);
or UO_1592 (O_1592,N_19018,N_19510);
nand UO_1593 (O_1593,N_19636,N_19850);
and UO_1594 (O_1594,N_19136,N_19867);
or UO_1595 (O_1595,N_19980,N_19926);
nor UO_1596 (O_1596,N_19870,N_19524);
or UO_1597 (O_1597,N_19321,N_19440);
or UO_1598 (O_1598,N_19122,N_19996);
and UO_1599 (O_1599,N_19866,N_19718);
and UO_1600 (O_1600,N_19493,N_19068);
or UO_1601 (O_1601,N_19827,N_19326);
or UO_1602 (O_1602,N_19320,N_19982);
or UO_1603 (O_1603,N_19972,N_19323);
nor UO_1604 (O_1604,N_19073,N_19082);
nand UO_1605 (O_1605,N_19878,N_19957);
xor UO_1606 (O_1606,N_19256,N_19133);
or UO_1607 (O_1607,N_19012,N_19174);
nor UO_1608 (O_1608,N_19429,N_19488);
xnor UO_1609 (O_1609,N_19032,N_19136);
nand UO_1610 (O_1610,N_19314,N_19229);
nor UO_1611 (O_1611,N_19270,N_19863);
nand UO_1612 (O_1612,N_19702,N_19407);
xor UO_1613 (O_1613,N_19493,N_19320);
or UO_1614 (O_1614,N_19199,N_19542);
or UO_1615 (O_1615,N_19454,N_19759);
nor UO_1616 (O_1616,N_19637,N_19298);
nor UO_1617 (O_1617,N_19685,N_19575);
nand UO_1618 (O_1618,N_19736,N_19768);
nand UO_1619 (O_1619,N_19057,N_19494);
or UO_1620 (O_1620,N_19739,N_19064);
or UO_1621 (O_1621,N_19355,N_19466);
xnor UO_1622 (O_1622,N_19580,N_19267);
and UO_1623 (O_1623,N_19896,N_19087);
or UO_1624 (O_1624,N_19471,N_19170);
nor UO_1625 (O_1625,N_19557,N_19789);
xor UO_1626 (O_1626,N_19023,N_19238);
nand UO_1627 (O_1627,N_19896,N_19868);
and UO_1628 (O_1628,N_19707,N_19843);
nand UO_1629 (O_1629,N_19597,N_19886);
xor UO_1630 (O_1630,N_19114,N_19247);
and UO_1631 (O_1631,N_19130,N_19444);
nor UO_1632 (O_1632,N_19202,N_19432);
or UO_1633 (O_1633,N_19285,N_19646);
nor UO_1634 (O_1634,N_19564,N_19005);
or UO_1635 (O_1635,N_19750,N_19187);
xnor UO_1636 (O_1636,N_19055,N_19340);
xor UO_1637 (O_1637,N_19490,N_19592);
nor UO_1638 (O_1638,N_19823,N_19670);
and UO_1639 (O_1639,N_19678,N_19783);
and UO_1640 (O_1640,N_19299,N_19689);
nand UO_1641 (O_1641,N_19743,N_19779);
or UO_1642 (O_1642,N_19298,N_19904);
xnor UO_1643 (O_1643,N_19818,N_19681);
or UO_1644 (O_1644,N_19013,N_19169);
or UO_1645 (O_1645,N_19441,N_19171);
nand UO_1646 (O_1646,N_19822,N_19830);
or UO_1647 (O_1647,N_19998,N_19647);
nor UO_1648 (O_1648,N_19580,N_19939);
and UO_1649 (O_1649,N_19171,N_19486);
nor UO_1650 (O_1650,N_19292,N_19754);
or UO_1651 (O_1651,N_19906,N_19907);
nor UO_1652 (O_1652,N_19273,N_19337);
nand UO_1653 (O_1653,N_19075,N_19659);
xnor UO_1654 (O_1654,N_19753,N_19657);
nor UO_1655 (O_1655,N_19833,N_19054);
nor UO_1656 (O_1656,N_19648,N_19074);
or UO_1657 (O_1657,N_19310,N_19302);
xnor UO_1658 (O_1658,N_19142,N_19656);
xor UO_1659 (O_1659,N_19195,N_19218);
nor UO_1660 (O_1660,N_19447,N_19555);
nor UO_1661 (O_1661,N_19442,N_19359);
nor UO_1662 (O_1662,N_19208,N_19024);
xnor UO_1663 (O_1663,N_19705,N_19587);
or UO_1664 (O_1664,N_19285,N_19965);
nor UO_1665 (O_1665,N_19726,N_19287);
and UO_1666 (O_1666,N_19869,N_19687);
xor UO_1667 (O_1667,N_19652,N_19518);
xor UO_1668 (O_1668,N_19315,N_19296);
or UO_1669 (O_1669,N_19995,N_19699);
nor UO_1670 (O_1670,N_19081,N_19881);
xor UO_1671 (O_1671,N_19940,N_19761);
and UO_1672 (O_1672,N_19607,N_19141);
xor UO_1673 (O_1673,N_19046,N_19358);
nor UO_1674 (O_1674,N_19727,N_19402);
nand UO_1675 (O_1675,N_19481,N_19345);
nor UO_1676 (O_1676,N_19476,N_19505);
xor UO_1677 (O_1677,N_19357,N_19235);
nor UO_1678 (O_1678,N_19747,N_19321);
nor UO_1679 (O_1679,N_19055,N_19831);
nor UO_1680 (O_1680,N_19674,N_19186);
nand UO_1681 (O_1681,N_19741,N_19476);
xor UO_1682 (O_1682,N_19017,N_19599);
or UO_1683 (O_1683,N_19833,N_19424);
nand UO_1684 (O_1684,N_19038,N_19450);
nand UO_1685 (O_1685,N_19092,N_19441);
or UO_1686 (O_1686,N_19141,N_19347);
or UO_1687 (O_1687,N_19138,N_19152);
nor UO_1688 (O_1688,N_19358,N_19347);
nor UO_1689 (O_1689,N_19180,N_19977);
xnor UO_1690 (O_1690,N_19060,N_19390);
nor UO_1691 (O_1691,N_19016,N_19737);
nand UO_1692 (O_1692,N_19419,N_19684);
or UO_1693 (O_1693,N_19820,N_19130);
or UO_1694 (O_1694,N_19655,N_19703);
nand UO_1695 (O_1695,N_19573,N_19209);
or UO_1696 (O_1696,N_19993,N_19842);
and UO_1697 (O_1697,N_19457,N_19918);
nand UO_1698 (O_1698,N_19503,N_19791);
and UO_1699 (O_1699,N_19794,N_19150);
xor UO_1700 (O_1700,N_19648,N_19474);
xor UO_1701 (O_1701,N_19087,N_19361);
nor UO_1702 (O_1702,N_19491,N_19445);
and UO_1703 (O_1703,N_19549,N_19682);
nand UO_1704 (O_1704,N_19798,N_19671);
and UO_1705 (O_1705,N_19820,N_19618);
nand UO_1706 (O_1706,N_19663,N_19391);
xnor UO_1707 (O_1707,N_19229,N_19776);
or UO_1708 (O_1708,N_19061,N_19648);
nand UO_1709 (O_1709,N_19877,N_19444);
nand UO_1710 (O_1710,N_19290,N_19781);
and UO_1711 (O_1711,N_19876,N_19550);
xnor UO_1712 (O_1712,N_19440,N_19239);
and UO_1713 (O_1713,N_19884,N_19633);
nor UO_1714 (O_1714,N_19909,N_19787);
xor UO_1715 (O_1715,N_19633,N_19770);
nor UO_1716 (O_1716,N_19179,N_19310);
nor UO_1717 (O_1717,N_19628,N_19382);
xnor UO_1718 (O_1718,N_19235,N_19362);
and UO_1719 (O_1719,N_19962,N_19138);
or UO_1720 (O_1720,N_19208,N_19468);
xnor UO_1721 (O_1721,N_19224,N_19779);
and UO_1722 (O_1722,N_19385,N_19473);
and UO_1723 (O_1723,N_19060,N_19603);
nor UO_1724 (O_1724,N_19032,N_19321);
and UO_1725 (O_1725,N_19074,N_19109);
xor UO_1726 (O_1726,N_19727,N_19961);
and UO_1727 (O_1727,N_19034,N_19704);
nand UO_1728 (O_1728,N_19443,N_19844);
nor UO_1729 (O_1729,N_19813,N_19228);
nand UO_1730 (O_1730,N_19875,N_19036);
nand UO_1731 (O_1731,N_19828,N_19663);
nand UO_1732 (O_1732,N_19485,N_19218);
and UO_1733 (O_1733,N_19866,N_19100);
nand UO_1734 (O_1734,N_19239,N_19069);
xor UO_1735 (O_1735,N_19342,N_19033);
nand UO_1736 (O_1736,N_19555,N_19875);
xor UO_1737 (O_1737,N_19387,N_19140);
or UO_1738 (O_1738,N_19777,N_19907);
and UO_1739 (O_1739,N_19113,N_19975);
or UO_1740 (O_1740,N_19933,N_19834);
or UO_1741 (O_1741,N_19035,N_19031);
xnor UO_1742 (O_1742,N_19785,N_19049);
nand UO_1743 (O_1743,N_19427,N_19871);
and UO_1744 (O_1744,N_19988,N_19361);
and UO_1745 (O_1745,N_19004,N_19444);
nor UO_1746 (O_1746,N_19486,N_19364);
nand UO_1747 (O_1747,N_19355,N_19958);
nor UO_1748 (O_1748,N_19910,N_19941);
nand UO_1749 (O_1749,N_19964,N_19130);
or UO_1750 (O_1750,N_19157,N_19230);
or UO_1751 (O_1751,N_19465,N_19481);
nand UO_1752 (O_1752,N_19926,N_19239);
nor UO_1753 (O_1753,N_19271,N_19135);
and UO_1754 (O_1754,N_19840,N_19468);
or UO_1755 (O_1755,N_19482,N_19219);
nand UO_1756 (O_1756,N_19900,N_19837);
and UO_1757 (O_1757,N_19007,N_19031);
or UO_1758 (O_1758,N_19786,N_19301);
xnor UO_1759 (O_1759,N_19103,N_19174);
xor UO_1760 (O_1760,N_19146,N_19389);
and UO_1761 (O_1761,N_19186,N_19838);
nor UO_1762 (O_1762,N_19016,N_19506);
nor UO_1763 (O_1763,N_19777,N_19922);
xnor UO_1764 (O_1764,N_19487,N_19296);
or UO_1765 (O_1765,N_19398,N_19937);
and UO_1766 (O_1766,N_19726,N_19069);
and UO_1767 (O_1767,N_19687,N_19116);
nand UO_1768 (O_1768,N_19235,N_19100);
and UO_1769 (O_1769,N_19678,N_19410);
nand UO_1770 (O_1770,N_19377,N_19179);
nand UO_1771 (O_1771,N_19392,N_19489);
and UO_1772 (O_1772,N_19815,N_19511);
nor UO_1773 (O_1773,N_19703,N_19352);
and UO_1774 (O_1774,N_19350,N_19844);
and UO_1775 (O_1775,N_19702,N_19810);
or UO_1776 (O_1776,N_19283,N_19978);
and UO_1777 (O_1777,N_19323,N_19260);
or UO_1778 (O_1778,N_19432,N_19429);
xor UO_1779 (O_1779,N_19222,N_19431);
nand UO_1780 (O_1780,N_19946,N_19718);
nor UO_1781 (O_1781,N_19343,N_19057);
or UO_1782 (O_1782,N_19598,N_19514);
and UO_1783 (O_1783,N_19195,N_19600);
xor UO_1784 (O_1784,N_19893,N_19047);
or UO_1785 (O_1785,N_19128,N_19744);
and UO_1786 (O_1786,N_19926,N_19423);
nor UO_1787 (O_1787,N_19940,N_19730);
xnor UO_1788 (O_1788,N_19724,N_19175);
or UO_1789 (O_1789,N_19196,N_19763);
or UO_1790 (O_1790,N_19863,N_19408);
nand UO_1791 (O_1791,N_19023,N_19114);
xnor UO_1792 (O_1792,N_19898,N_19980);
and UO_1793 (O_1793,N_19514,N_19390);
nor UO_1794 (O_1794,N_19050,N_19562);
nand UO_1795 (O_1795,N_19249,N_19615);
or UO_1796 (O_1796,N_19891,N_19615);
nand UO_1797 (O_1797,N_19852,N_19890);
or UO_1798 (O_1798,N_19532,N_19131);
nand UO_1799 (O_1799,N_19093,N_19670);
nand UO_1800 (O_1800,N_19034,N_19698);
xor UO_1801 (O_1801,N_19173,N_19799);
and UO_1802 (O_1802,N_19954,N_19773);
nor UO_1803 (O_1803,N_19388,N_19381);
and UO_1804 (O_1804,N_19158,N_19464);
or UO_1805 (O_1805,N_19867,N_19376);
nand UO_1806 (O_1806,N_19138,N_19664);
nand UO_1807 (O_1807,N_19217,N_19367);
nor UO_1808 (O_1808,N_19413,N_19473);
xor UO_1809 (O_1809,N_19010,N_19285);
and UO_1810 (O_1810,N_19429,N_19269);
nor UO_1811 (O_1811,N_19452,N_19621);
xor UO_1812 (O_1812,N_19809,N_19927);
xor UO_1813 (O_1813,N_19033,N_19887);
nand UO_1814 (O_1814,N_19197,N_19195);
nor UO_1815 (O_1815,N_19835,N_19159);
xnor UO_1816 (O_1816,N_19807,N_19586);
nand UO_1817 (O_1817,N_19680,N_19557);
or UO_1818 (O_1818,N_19865,N_19532);
and UO_1819 (O_1819,N_19347,N_19075);
nor UO_1820 (O_1820,N_19386,N_19379);
xor UO_1821 (O_1821,N_19573,N_19462);
and UO_1822 (O_1822,N_19956,N_19961);
or UO_1823 (O_1823,N_19506,N_19175);
xor UO_1824 (O_1824,N_19596,N_19733);
or UO_1825 (O_1825,N_19986,N_19688);
nor UO_1826 (O_1826,N_19581,N_19370);
nor UO_1827 (O_1827,N_19744,N_19068);
nor UO_1828 (O_1828,N_19591,N_19529);
xnor UO_1829 (O_1829,N_19325,N_19496);
nor UO_1830 (O_1830,N_19531,N_19365);
or UO_1831 (O_1831,N_19466,N_19502);
xor UO_1832 (O_1832,N_19309,N_19228);
or UO_1833 (O_1833,N_19840,N_19983);
or UO_1834 (O_1834,N_19326,N_19954);
xor UO_1835 (O_1835,N_19874,N_19419);
xnor UO_1836 (O_1836,N_19733,N_19230);
or UO_1837 (O_1837,N_19908,N_19038);
nor UO_1838 (O_1838,N_19852,N_19572);
and UO_1839 (O_1839,N_19901,N_19157);
nor UO_1840 (O_1840,N_19061,N_19552);
and UO_1841 (O_1841,N_19673,N_19084);
nor UO_1842 (O_1842,N_19936,N_19542);
nor UO_1843 (O_1843,N_19529,N_19239);
or UO_1844 (O_1844,N_19771,N_19685);
and UO_1845 (O_1845,N_19258,N_19962);
nand UO_1846 (O_1846,N_19460,N_19386);
nand UO_1847 (O_1847,N_19094,N_19715);
xor UO_1848 (O_1848,N_19387,N_19534);
xor UO_1849 (O_1849,N_19128,N_19997);
nand UO_1850 (O_1850,N_19432,N_19108);
nand UO_1851 (O_1851,N_19913,N_19138);
or UO_1852 (O_1852,N_19474,N_19745);
and UO_1853 (O_1853,N_19886,N_19676);
or UO_1854 (O_1854,N_19158,N_19693);
xnor UO_1855 (O_1855,N_19850,N_19668);
and UO_1856 (O_1856,N_19074,N_19955);
or UO_1857 (O_1857,N_19761,N_19450);
nand UO_1858 (O_1858,N_19693,N_19232);
nand UO_1859 (O_1859,N_19680,N_19537);
nor UO_1860 (O_1860,N_19109,N_19391);
xor UO_1861 (O_1861,N_19134,N_19360);
xnor UO_1862 (O_1862,N_19189,N_19991);
nand UO_1863 (O_1863,N_19762,N_19927);
nand UO_1864 (O_1864,N_19202,N_19069);
and UO_1865 (O_1865,N_19851,N_19136);
or UO_1866 (O_1866,N_19133,N_19795);
nand UO_1867 (O_1867,N_19601,N_19783);
or UO_1868 (O_1868,N_19770,N_19203);
and UO_1869 (O_1869,N_19554,N_19882);
nor UO_1870 (O_1870,N_19573,N_19771);
nand UO_1871 (O_1871,N_19816,N_19793);
xnor UO_1872 (O_1872,N_19538,N_19389);
and UO_1873 (O_1873,N_19453,N_19164);
nand UO_1874 (O_1874,N_19869,N_19742);
nand UO_1875 (O_1875,N_19469,N_19272);
nand UO_1876 (O_1876,N_19855,N_19126);
or UO_1877 (O_1877,N_19406,N_19503);
or UO_1878 (O_1878,N_19248,N_19635);
and UO_1879 (O_1879,N_19146,N_19087);
or UO_1880 (O_1880,N_19046,N_19896);
nor UO_1881 (O_1881,N_19621,N_19914);
and UO_1882 (O_1882,N_19550,N_19194);
and UO_1883 (O_1883,N_19058,N_19307);
nor UO_1884 (O_1884,N_19690,N_19417);
xor UO_1885 (O_1885,N_19983,N_19882);
or UO_1886 (O_1886,N_19368,N_19987);
or UO_1887 (O_1887,N_19593,N_19960);
and UO_1888 (O_1888,N_19253,N_19010);
nand UO_1889 (O_1889,N_19554,N_19545);
and UO_1890 (O_1890,N_19166,N_19612);
xor UO_1891 (O_1891,N_19966,N_19038);
and UO_1892 (O_1892,N_19252,N_19113);
nand UO_1893 (O_1893,N_19921,N_19616);
and UO_1894 (O_1894,N_19474,N_19037);
or UO_1895 (O_1895,N_19082,N_19144);
xor UO_1896 (O_1896,N_19324,N_19744);
nor UO_1897 (O_1897,N_19676,N_19280);
and UO_1898 (O_1898,N_19269,N_19508);
nand UO_1899 (O_1899,N_19588,N_19366);
xor UO_1900 (O_1900,N_19263,N_19007);
nand UO_1901 (O_1901,N_19361,N_19907);
and UO_1902 (O_1902,N_19869,N_19078);
or UO_1903 (O_1903,N_19177,N_19678);
nor UO_1904 (O_1904,N_19184,N_19640);
xnor UO_1905 (O_1905,N_19066,N_19306);
nor UO_1906 (O_1906,N_19669,N_19087);
nand UO_1907 (O_1907,N_19793,N_19564);
nor UO_1908 (O_1908,N_19562,N_19136);
nor UO_1909 (O_1909,N_19737,N_19863);
or UO_1910 (O_1910,N_19269,N_19923);
nor UO_1911 (O_1911,N_19965,N_19835);
nand UO_1912 (O_1912,N_19129,N_19241);
and UO_1913 (O_1913,N_19856,N_19290);
and UO_1914 (O_1914,N_19282,N_19218);
nand UO_1915 (O_1915,N_19070,N_19870);
nor UO_1916 (O_1916,N_19890,N_19600);
nand UO_1917 (O_1917,N_19052,N_19674);
or UO_1918 (O_1918,N_19002,N_19417);
and UO_1919 (O_1919,N_19001,N_19206);
nand UO_1920 (O_1920,N_19341,N_19865);
nand UO_1921 (O_1921,N_19514,N_19207);
nor UO_1922 (O_1922,N_19361,N_19532);
xor UO_1923 (O_1923,N_19398,N_19334);
nand UO_1924 (O_1924,N_19959,N_19484);
or UO_1925 (O_1925,N_19558,N_19012);
and UO_1926 (O_1926,N_19782,N_19771);
or UO_1927 (O_1927,N_19397,N_19613);
and UO_1928 (O_1928,N_19483,N_19424);
nand UO_1929 (O_1929,N_19432,N_19564);
and UO_1930 (O_1930,N_19645,N_19994);
nor UO_1931 (O_1931,N_19124,N_19396);
nor UO_1932 (O_1932,N_19014,N_19387);
or UO_1933 (O_1933,N_19793,N_19779);
nor UO_1934 (O_1934,N_19511,N_19585);
or UO_1935 (O_1935,N_19137,N_19139);
xor UO_1936 (O_1936,N_19838,N_19356);
or UO_1937 (O_1937,N_19694,N_19927);
xnor UO_1938 (O_1938,N_19883,N_19091);
nand UO_1939 (O_1939,N_19449,N_19602);
nor UO_1940 (O_1940,N_19910,N_19422);
nand UO_1941 (O_1941,N_19413,N_19400);
or UO_1942 (O_1942,N_19866,N_19856);
nand UO_1943 (O_1943,N_19547,N_19989);
xnor UO_1944 (O_1944,N_19854,N_19910);
xor UO_1945 (O_1945,N_19586,N_19290);
nor UO_1946 (O_1946,N_19106,N_19725);
nand UO_1947 (O_1947,N_19919,N_19126);
or UO_1948 (O_1948,N_19281,N_19677);
nor UO_1949 (O_1949,N_19093,N_19347);
xor UO_1950 (O_1950,N_19548,N_19883);
nand UO_1951 (O_1951,N_19906,N_19098);
nand UO_1952 (O_1952,N_19421,N_19696);
xor UO_1953 (O_1953,N_19198,N_19399);
or UO_1954 (O_1954,N_19454,N_19923);
xnor UO_1955 (O_1955,N_19566,N_19960);
nor UO_1956 (O_1956,N_19847,N_19413);
nor UO_1957 (O_1957,N_19989,N_19529);
nor UO_1958 (O_1958,N_19527,N_19874);
nor UO_1959 (O_1959,N_19003,N_19467);
and UO_1960 (O_1960,N_19288,N_19676);
xor UO_1961 (O_1961,N_19661,N_19588);
xnor UO_1962 (O_1962,N_19180,N_19996);
xor UO_1963 (O_1963,N_19286,N_19873);
or UO_1964 (O_1964,N_19871,N_19674);
or UO_1965 (O_1965,N_19268,N_19558);
and UO_1966 (O_1966,N_19820,N_19187);
and UO_1967 (O_1967,N_19793,N_19084);
xor UO_1968 (O_1968,N_19384,N_19117);
or UO_1969 (O_1969,N_19343,N_19075);
or UO_1970 (O_1970,N_19958,N_19080);
nand UO_1971 (O_1971,N_19629,N_19391);
xnor UO_1972 (O_1972,N_19118,N_19807);
and UO_1973 (O_1973,N_19384,N_19670);
and UO_1974 (O_1974,N_19712,N_19135);
and UO_1975 (O_1975,N_19354,N_19803);
or UO_1976 (O_1976,N_19257,N_19867);
nor UO_1977 (O_1977,N_19377,N_19549);
nand UO_1978 (O_1978,N_19777,N_19330);
nand UO_1979 (O_1979,N_19588,N_19451);
and UO_1980 (O_1980,N_19925,N_19589);
xnor UO_1981 (O_1981,N_19891,N_19766);
or UO_1982 (O_1982,N_19625,N_19096);
xor UO_1983 (O_1983,N_19902,N_19241);
xnor UO_1984 (O_1984,N_19689,N_19092);
and UO_1985 (O_1985,N_19021,N_19895);
nand UO_1986 (O_1986,N_19394,N_19084);
and UO_1987 (O_1987,N_19290,N_19971);
or UO_1988 (O_1988,N_19776,N_19026);
xor UO_1989 (O_1989,N_19552,N_19595);
xnor UO_1990 (O_1990,N_19320,N_19103);
or UO_1991 (O_1991,N_19801,N_19874);
xor UO_1992 (O_1992,N_19546,N_19788);
nor UO_1993 (O_1993,N_19462,N_19476);
and UO_1994 (O_1994,N_19187,N_19792);
nand UO_1995 (O_1995,N_19039,N_19390);
nor UO_1996 (O_1996,N_19631,N_19770);
nor UO_1997 (O_1997,N_19554,N_19963);
or UO_1998 (O_1998,N_19710,N_19047);
nand UO_1999 (O_1999,N_19306,N_19075);
or UO_2000 (O_2000,N_19012,N_19136);
nor UO_2001 (O_2001,N_19417,N_19433);
and UO_2002 (O_2002,N_19668,N_19129);
nor UO_2003 (O_2003,N_19005,N_19670);
nand UO_2004 (O_2004,N_19921,N_19810);
or UO_2005 (O_2005,N_19524,N_19081);
and UO_2006 (O_2006,N_19818,N_19159);
nor UO_2007 (O_2007,N_19538,N_19294);
xnor UO_2008 (O_2008,N_19376,N_19054);
nand UO_2009 (O_2009,N_19139,N_19758);
nand UO_2010 (O_2010,N_19456,N_19654);
or UO_2011 (O_2011,N_19628,N_19818);
nand UO_2012 (O_2012,N_19656,N_19292);
nor UO_2013 (O_2013,N_19928,N_19767);
and UO_2014 (O_2014,N_19126,N_19522);
and UO_2015 (O_2015,N_19642,N_19804);
or UO_2016 (O_2016,N_19215,N_19040);
xnor UO_2017 (O_2017,N_19084,N_19724);
xor UO_2018 (O_2018,N_19853,N_19563);
or UO_2019 (O_2019,N_19704,N_19577);
or UO_2020 (O_2020,N_19771,N_19044);
xnor UO_2021 (O_2021,N_19897,N_19887);
nor UO_2022 (O_2022,N_19720,N_19916);
nor UO_2023 (O_2023,N_19238,N_19473);
nand UO_2024 (O_2024,N_19598,N_19576);
and UO_2025 (O_2025,N_19983,N_19326);
nor UO_2026 (O_2026,N_19731,N_19804);
nand UO_2027 (O_2027,N_19444,N_19203);
xnor UO_2028 (O_2028,N_19037,N_19950);
or UO_2029 (O_2029,N_19765,N_19288);
or UO_2030 (O_2030,N_19532,N_19162);
nor UO_2031 (O_2031,N_19858,N_19497);
or UO_2032 (O_2032,N_19612,N_19297);
nor UO_2033 (O_2033,N_19528,N_19373);
nand UO_2034 (O_2034,N_19042,N_19945);
nand UO_2035 (O_2035,N_19194,N_19043);
nor UO_2036 (O_2036,N_19440,N_19387);
xnor UO_2037 (O_2037,N_19447,N_19840);
xnor UO_2038 (O_2038,N_19315,N_19094);
xor UO_2039 (O_2039,N_19146,N_19039);
or UO_2040 (O_2040,N_19146,N_19726);
xnor UO_2041 (O_2041,N_19100,N_19242);
and UO_2042 (O_2042,N_19082,N_19489);
or UO_2043 (O_2043,N_19813,N_19604);
and UO_2044 (O_2044,N_19737,N_19206);
or UO_2045 (O_2045,N_19227,N_19862);
nor UO_2046 (O_2046,N_19358,N_19254);
nand UO_2047 (O_2047,N_19819,N_19446);
nand UO_2048 (O_2048,N_19893,N_19157);
nor UO_2049 (O_2049,N_19446,N_19590);
xnor UO_2050 (O_2050,N_19652,N_19797);
or UO_2051 (O_2051,N_19001,N_19432);
xor UO_2052 (O_2052,N_19703,N_19734);
and UO_2053 (O_2053,N_19895,N_19514);
nor UO_2054 (O_2054,N_19263,N_19997);
nor UO_2055 (O_2055,N_19149,N_19136);
nand UO_2056 (O_2056,N_19277,N_19458);
or UO_2057 (O_2057,N_19546,N_19649);
nand UO_2058 (O_2058,N_19785,N_19153);
and UO_2059 (O_2059,N_19230,N_19618);
and UO_2060 (O_2060,N_19879,N_19240);
or UO_2061 (O_2061,N_19423,N_19891);
nor UO_2062 (O_2062,N_19185,N_19961);
or UO_2063 (O_2063,N_19115,N_19119);
and UO_2064 (O_2064,N_19855,N_19140);
nand UO_2065 (O_2065,N_19935,N_19168);
or UO_2066 (O_2066,N_19892,N_19634);
and UO_2067 (O_2067,N_19375,N_19969);
xnor UO_2068 (O_2068,N_19884,N_19715);
and UO_2069 (O_2069,N_19477,N_19549);
nand UO_2070 (O_2070,N_19894,N_19914);
xor UO_2071 (O_2071,N_19478,N_19718);
nand UO_2072 (O_2072,N_19987,N_19136);
nand UO_2073 (O_2073,N_19867,N_19719);
xor UO_2074 (O_2074,N_19050,N_19813);
nand UO_2075 (O_2075,N_19453,N_19535);
nor UO_2076 (O_2076,N_19429,N_19681);
xnor UO_2077 (O_2077,N_19896,N_19768);
or UO_2078 (O_2078,N_19172,N_19799);
and UO_2079 (O_2079,N_19650,N_19934);
xnor UO_2080 (O_2080,N_19691,N_19706);
xnor UO_2081 (O_2081,N_19295,N_19798);
xnor UO_2082 (O_2082,N_19664,N_19315);
or UO_2083 (O_2083,N_19116,N_19425);
xor UO_2084 (O_2084,N_19401,N_19122);
and UO_2085 (O_2085,N_19738,N_19056);
nor UO_2086 (O_2086,N_19844,N_19480);
xor UO_2087 (O_2087,N_19920,N_19252);
or UO_2088 (O_2088,N_19874,N_19798);
nand UO_2089 (O_2089,N_19035,N_19739);
nor UO_2090 (O_2090,N_19091,N_19940);
nand UO_2091 (O_2091,N_19496,N_19638);
nor UO_2092 (O_2092,N_19580,N_19787);
nand UO_2093 (O_2093,N_19857,N_19124);
nand UO_2094 (O_2094,N_19329,N_19069);
nor UO_2095 (O_2095,N_19534,N_19309);
and UO_2096 (O_2096,N_19846,N_19854);
nand UO_2097 (O_2097,N_19497,N_19772);
xnor UO_2098 (O_2098,N_19304,N_19654);
or UO_2099 (O_2099,N_19115,N_19586);
and UO_2100 (O_2100,N_19176,N_19531);
nor UO_2101 (O_2101,N_19755,N_19202);
nor UO_2102 (O_2102,N_19134,N_19371);
nand UO_2103 (O_2103,N_19144,N_19126);
nor UO_2104 (O_2104,N_19849,N_19783);
xnor UO_2105 (O_2105,N_19942,N_19293);
xnor UO_2106 (O_2106,N_19625,N_19875);
xor UO_2107 (O_2107,N_19990,N_19002);
nand UO_2108 (O_2108,N_19163,N_19745);
nand UO_2109 (O_2109,N_19758,N_19746);
xnor UO_2110 (O_2110,N_19609,N_19259);
or UO_2111 (O_2111,N_19133,N_19544);
nand UO_2112 (O_2112,N_19960,N_19422);
xor UO_2113 (O_2113,N_19602,N_19401);
and UO_2114 (O_2114,N_19450,N_19692);
nand UO_2115 (O_2115,N_19663,N_19580);
and UO_2116 (O_2116,N_19402,N_19407);
and UO_2117 (O_2117,N_19852,N_19562);
and UO_2118 (O_2118,N_19201,N_19856);
or UO_2119 (O_2119,N_19398,N_19032);
nand UO_2120 (O_2120,N_19584,N_19927);
nand UO_2121 (O_2121,N_19776,N_19672);
nor UO_2122 (O_2122,N_19084,N_19729);
nor UO_2123 (O_2123,N_19165,N_19607);
and UO_2124 (O_2124,N_19582,N_19386);
and UO_2125 (O_2125,N_19527,N_19545);
and UO_2126 (O_2126,N_19720,N_19545);
nand UO_2127 (O_2127,N_19581,N_19146);
or UO_2128 (O_2128,N_19552,N_19783);
xnor UO_2129 (O_2129,N_19465,N_19081);
and UO_2130 (O_2130,N_19250,N_19056);
or UO_2131 (O_2131,N_19359,N_19602);
and UO_2132 (O_2132,N_19899,N_19225);
xnor UO_2133 (O_2133,N_19749,N_19192);
xnor UO_2134 (O_2134,N_19990,N_19409);
nor UO_2135 (O_2135,N_19538,N_19321);
nand UO_2136 (O_2136,N_19613,N_19393);
xnor UO_2137 (O_2137,N_19690,N_19188);
or UO_2138 (O_2138,N_19294,N_19221);
xnor UO_2139 (O_2139,N_19962,N_19408);
nand UO_2140 (O_2140,N_19418,N_19713);
and UO_2141 (O_2141,N_19732,N_19602);
and UO_2142 (O_2142,N_19813,N_19082);
xnor UO_2143 (O_2143,N_19264,N_19430);
xnor UO_2144 (O_2144,N_19224,N_19482);
and UO_2145 (O_2145,N_19051,N_19805);
nand UO_2146 (O_2146,N_19683,N_19316);
xor UO_2147 (O_2147,N_19834,N_19848);
xnor UO_2148 (O_2148,N_19617,N_19234);
nor UO_2149 (O_2149,N_19391,N_19316);
xor UO_2150 (O_2150,N_19129,N_19747);
nand UO_2151 (O_2151,N_19580,N_19537);
or UO_2152 (O_2152,N_19856,N_19704);
xor UO_2153 (O_2153,N_19939,N_19913);
nor UO_2154 (O_2154,N_19665,N_19424);
nor UO_2155 (O_2155,N_19781,N_19682);
xnor UO_2156 (O_2156,N_19038,N_19755);
nor UO_2157 (O_2157,N_19748,N_19536);
xor UO_2158 (O_2158,N_19143,N_19025);
nor UO_2159 (O_2159,N_19695,N_19894);
nand UO_2160 (O_2160,N_19161,N_19730);
xnor UO_2161 (O_2161,N_19887,N_19945);
xnor UO_2162 (O_2162,N_19010,N_19552);
nand UO_2163 (O_2163,N_19994,N_19247);
or UO_2164 (O_2164,N_19717,N_19530);
xnor UO_2165 (O_2165,N_19098,N_19516);
nand UO_2166 (O_2166,N_19065,N_19272);
or UO_2167 (O_2167,N_19159,N_19077);
xor UO_2168 (O_2168,N_19875,N_19004);
xnor UO_2169 (O_2169,N_19452,N_19509);
and UO_2170 (O_2170,N_19886,N_19699);
nand UO_2171 (O_2171,N_19121,N_19802);
nor UO_2172 (O_2172,N_19405,N_19667);
nor UO_2173 (O_2173,N_19839,N_19177);
nor UO_2174 (O_2174,N_19342,N_19604);
or UO_2175 (O_2175,N_19472,N_19857);
nor UO_2176 (O_2176,N_19083,N_19036);
nand UO_2177 (O_2177,N_19895,N_19914);
and UO_2178 (O_2178,N_19402,N_19458);
or UO_2179 (O_2179,N_19507,N_19819);
nor UO_2180 (O_2180,N_19198,N_19595);
xnor UO_2181 (O_2181,N_19974,N_19912);
nand UO_2182 (O_2182,N_19917,N_19517);
nand UO_2183 (O_2183,N_19683,N_19639);
xor UO_2184 (O_2184,N_19933,N_19576);
and UO_2185 (O_2185,N_19279,N_19825);
nand UO_2186 (O_2186,N_19948,N_19913);
nor UO_2187 (O_2187,N_19390,N_19170);
or UO_2188 (O_2188,N_19634,N_19626);
or UO_2189 (O_2189,N_19181,N_19312);
and UO_2190 (O_2190,N_19973,N_19734);
and UO_2191 (O_2191,N_19551,N_19598);
xnor UO_2192 (O_2192,N_19360,N_19208);
and UO_2193 (O_2193,N_19807,N_19308);
nor UO_2194 (O_2194,N_19378,N_19539);
xor UO_2195 (O_2195,N_19697,N_19891);
and UO_2196 (O_2196,N_19136,N_19072);
and UO_2197 (O_2197,N_19541,N_19010);
nand UO_2198 (O_2198,N_19225,N_19005);
nand UO_2199 (O_2199,N_19929,N_19433);
xnor UO_2200 (O_2200,N_19379,N_19126);
xnor UO_2201 (O_2201,N_19298,N_19280);
and UO_2202 (O_2202,N_19317,N_19426);
nand UO_2203 (O_2203,N_19859,N_19879);
nor UO_2204 (O_2204,N_19101,N_19876);
nor UO_2205 (O_2205,N_19712,N_19599);
xnor UO_2206 (O_2206,N_19013,N_19228);
xnor UO_2207 (O_2207,N_19310,N_19868);
or UO_2208 (O_2208,N_19635,N_19261);
nand UO_2209 (O_2209,N_19399,N_19984);
nand UO_2210 (O_2210,N_19699,N_19814);
and UO_2211 (O_2211,N_19841,N_19732);
nand UO_2212 (O_2212,N_19827,N_19652);
nor UO_2213 (O_2213,N_19513,N_19361);
or UO_2214 (O_2214,N_19794,N_19534);
nand UO_2215 (O_2215,N_19602,N_19366);
nand UO_2216 (O_2216,N_19375,N_19458);
nor UO_2217 (O_2217,N_19024,N_19679);
nor UO_2218 (O_2218,N_19797,N_19618);
nand UO_2219 (O_2219,N_19033,N_19977);
nor UO_2220 (O_2220,N_19213,N_19185);
nand UO_2221 (O_2221,N_19045,N_19962);
and UO_2222 (O_2222,N_19906,N_19854);
or UO_2223 (O_2223,N_19914,N_19318);
nor UO_2224 (O_2224,N_19412,N_19878);
and UO_2225 (O_2225,N_19578,N_19211);
nor UO_2226 (O_2226,N_19347,N_19977);
xnor UO_2227 (O_2227,N_19389,N_19505);
xor UO_2228 (O_2228,N_19119,N_19608);
nor UO_2229 (O_2229,N_19160,N_19725);
or UO_2230 (O_2230,N_19653,N_19509);
or UO_2231 (O_2231,N_19758,N_19080);
and UO_2232 (O_2232,N_19640,N_19558);
or UO_2233 (O_2233,N_19110,N_19190);
or UO_2234 (O_2234,N_19172,N_19486);
and UO_2235 (O_2235,N_19011,N_19979);
or UO_2236 (O_2236,N_19833,N_19283);
and UO_2237 (O_2237,N_19241,N_19906);
and UO_2238 (O_2238,N_19151,N_19767);
and UO_2239 (O_2239,N_19700,N_19118);
nor UO_2240 (O_2240,N_19680,N_19806);
nor UO_2241 (O_2241,N_19953,N_19143);
nand UO_2242 (O_2242,N_19589,N_19879);
and UO_2243 (O_2243,N_19183,N_19030);
and UO_2244 (O_2244,N_19588,N_19441);
nand UO_2245 (O_2245,N_19587,N_19194);
nand UO_2246 (O_2246,N_19220,N_19213);
or UO_2247 (O_2247,N_19220,N_19926);
nand UO_2248 (O_2248,N_19812,N_19749);
nor UO_2249 (O_2249,N_19765,N_19651);
and UO_2250 (O_2250,N_19754,N_19323);
or UO_2251 (O_2251,N_19497,N_19195);
nand UO_2252 (O_2252,N_19002,N_19421);
xnor UO_2253 (O_2253,N_19230,N_19049);
and UO_2254 (O_2254,N_19189,N_19716);
or UO_2255 (O_2255,N_19142,N_19685);
and UO_2256 (O_2256,N_19700,N_19657);
or UO_2257 (O_2257,N_19873,N_19493);
nor UO_2258 (O_2258,N_19961,N_19771);
nand UO_2259 (O_2259,N_19482,N_19359);
xor UO_2260 (O_2260,N_19031,N_19937);
or UO_2261 (O_2261,N_19019,N_19521);
and UO_2262 (O_2262,N_19593,N_19380);
nor UO_2263 (O_2263,N_19326,N_19951);
xor UO_2264 (O_2264,N_19644,N_19858);
and UO_2265 (O_2265,N_19931,N_19755);
nor UO_2266 (O_2266,N_19120,N_19083);
nor UO_2267 (O_2267,N_19345,N_19925);
nand UO_2268 (O_2268,N_19949,N_19591);
or UO_2269 (O_2269,N_19275,N_19550);
nor UO_2270 (O_2270,N_19158,N_19629);
nor UO_2271 (O_2271,N_19608,N_19964);
or UO_2272 (O_2272,N_19254,N_19714);
and UO_2273 (O_2273,N_19460,N_19189);
nand UO_2274 (O_2274,N_19903,N_19374);
xor UO_2275 (O_2275,N_19725,N_19729);
or UO_2276 (O_2276,N_19661,N_19938);
or UO_2277 (O_2277,N_19714,N_19871);
nor UO_2278 (O_2278,N_19402,N_19642);
nand UO_2279 (O_2279,N_19769,N_19616);
nand UO_2280 (O_2280,N_19143,N_19986);
nand UO_2281 (O_2281,N_19765,N_19968);
or UO_2282 (O_2282,N_19458,N_19745);
or UO_2283 (O_2283,N_19690,N_19546);
and UO_2284 (O_2284,N_19132,N_19915);
and UO_2285 (O_2285,N_19226,N_19603);
nor UO_2286 (O_2286,N_19162,N_19763);
xor UO_2287 (O_2287,N_19942,N_19094);
nand UO_2288 (O_2288,N_19951,N_19220);
xor UO_2289 (O_2289,N_19838,N_19483);
xnor UO_2290 (O_2290,N_19507,N_19355);
or UO_2291 (O_2291,N_19337,N_19373);
xor UO_2292 (O_2292,N_19128,N_19257);
and UO_2293 (O_2293,N_19405,N_19520);
nand UO_2294 (O_2294,N_19192,N_19748);
nand UO_2295 (O_2295,N_19938,N_19352);
xor UO_2296 (O_2296,N_19442,N_19556);
and UO_2297 (O_2297,N_19196,N_19446);
nor UO_2298 (O_2298,N_19809,N_19193);
nor UO_2299 (O_2299,N_19054,N_19413);
or UO_2300 (O_2300,N_19004,N_19987);
nor UO_2301 (O_2301,N_19596,N_19921);
or UO_2302 (O_2302,N_19074,N_19950);
and UO_2303 (O_2303,N_19552,N_19598);
or UO_2304 (O_2304,N_19738,N_19662);
or UO_2305 (O_2305,N_19450,N_19760);
xnor UO_2306 (O_2306,N_19565,N_19252);
or UO_2307 (O_2307,N_19387,N_19610);
nand UO_2308 (O_2308,N_19003,N_19309);
or UO_2309 (O_2309,N_19447,N_19576);
nor UO_2310 (O_2310,N_19497,N_19385);
or UO_2311 (O_2311,N_19124,N_19767);
xor UO_2312 (O_2312,N_19362,N_19858);
xnor UO_2313 (O_2313,N_19155,N_19943);
and UO_2314 (O_2314,N_19317,N_19199);
or UO_2315 (O_2315,N_19296,N_19195);
and UO_2316 (O_2316,N_19194,N_19022);
nand UO_2317 (O_2317,N_19878,N_19975);
nor UO_2318 (O_2318,N_19809,N_19082);
xor UO_2319 (O_2319,N_19857,N_19271);
nor UO_2320 (O_2320,N_19664,N_19207);
nand UO_2321 (O_2321,N_19702,N_19552);
xor UO_2322 (O_2322,N_19244,N_19539);
nand UO_2323 (O_2323,N_19923,N_19498);
xnor UO_2324 (O_2324,N_19370,N_19763);
or UO_2325 (O_2325,N_19300,N_19527);
nor UO_2326 (O_2326,N_19657,N_19146);
or UO_2327 (O_2327,N_19825,N_19839);
nor UO_2328 (O_2328,N_19164,N_19035);
nand UO_2329 (O_2329,N_19225,N_19568);
nor UO_2330 (O_2330,N_19041,N_19778);
or UO_2331 (O_2331,N_19352,N_19227);
and UO_2332 (O_2332,N_19374,N_19299);
nor UO_2333 (O_2333,N_19946,N_19433);
nor UO_2334 (O_2334,N_19832,N_19905);
and UO_2335 (O_2335,N_19092,N_19483);
nand UO_2336 (O_2336,N_19471,N_19336);
nand UO_2337 (O_2337,N_19851,N_19710);
nand UO_2338 (O_2338,N_19976,N_19924);
nand UO_2339 (O_2339,N_19798,N_19479);
nand UO_2340 (O_2340,N_19941,N_19358);
xnor UO_2341 (O_2341,N_19894,N_19768);
or UO_2342 (O_2342,N_19487,N_19861);
xnor UO_2343 (O_2343,N_19037,N_19125);
nand UO_2344 (O_2344,N_19891,N_19829);
nand UO_2345 (O_2345,N_19502,N_19575);
xor UO_2346 (O_2346,N_19100,N_19423);
xor UO_2347 (O_2347,N_19486,N_19943);
and UO_2348 (O_2348,N_19021,N_19555);
or UO_2349 (O_2349,N_19388,N_19514);
nand UO_2350 (O_2350,N_19722,N_19759);
xnor UO_2351 (O_2351,N_19350,N_19614);
xnor UO_2352 (O_2352,N_19038,N_19096);
xor UO_2353 (O_2353,N_19542,N_19237);
nand UO_2354 (O_2354,N_19692,N_19972);
xnor UO_2355 (O_2355,N_19565,N_19354);
nor UO_2356 (O_2356,N_19516,N_19111);
nand UO_2357 (O_2357,N_19372,N_19105);
or UO_2358 (O_2358,N_19555,N_19459);
or UO_2359 (O_2359,N_19801,N_19144);
or UO_2360 (O_2360,N_19281,N_19776);
or UO_2361 (O_2361,N_19930,N_19077);
or UO_2362 (O_2362,N_19948,N_19535);
or UO_2363 (O_2363,N_19166,N_19269);
nor UO_2364 (O_2364,N_19258,N_19457);
and UO_2365 (O_2365,N_19798,N_19754);
nor UO_2366 (O_2366,N_19696,N_19941);
nor UO_2367 (O_2367,N_19117,N_19131);
nand UO_2368 (O_2368,N_19236,N_19443);
nor UO_2369 (O_2369,N_19139,N_19535);
nand UO_2370 (O_2370,N_19780,N_19725);
xor UO_2371 (O_2371,N_19876,N_19316);
nor UO_2372 (O_2372,N_19173,N_19422);
nor UO_2373 (O_2373,N_19529,N_19961);
nor UO_2374 (O_2374,N_19889,N_19233);
and UO_2375 (O_2375,N_19732,N_19024);
xnor UO_2376 (O_2376,N_19203,N_19687);
nor UO_2377 (O_2377,N_19268,N_19726);
nor UO_2378 (O_2378,N_19073,N_19021);
nand UO_2379 (O_2379,N_19617,N_19086);
or UO_2380 (O_2380,N_19388,N_19014);
xnor UO_2381 (O_2381,N_19934,N_19796);
nor UO_2382 (O_2382,N_19595,N_19800);
nand UO_2383 (O_2383,N_19522,N_19414);
xnor UO_2384 (O_2384,N_19747,N_19912);
nor UO_2385 (O_2385,N_19636,N_19852);
nor UO_2386 (O_2386,N_19631,N_19554);
and UO_2387 (O_2387,N_19140,N_19399);
nand UO_2388 (O_2388,N_19561,N_19736);
or UO_2389 (O_2389,N_19270,N_19508);
or UO_2390 (O_2390,N_19864,N_19020);
and UO_2391 (O_2391,N_19656,N_19859);
nand UO_2392 (O_2392,N_19973,N_19872);
and UO_2393 (O_2393,N_19774,N_19479);
and UO_2394 (O_2394,N_19155,N_19199);
nand UO_2395 (O_2395,N_19406,N_19068);
xor UO_2396 (O_2396,N_19043,N_19106);
xnor UO_2397 (O_2397,N_19816,N_19289);
and UO_2398 (O_2398,N_19251,N_19351);
xor UO_2399 (O_2399,N_19378,N_19897);
or UO_2400 (O_2400,N_19448,N_19962);
and UO_2401 (O_2401,N_19117,N_19003);
or UO_2402 (O_2402,N_19378,N_19075);
xor UO_2403 (O_2403,N_19233,N_19113);
nor UO_2404 (O_2404,N_19587,N_19135);
or UO_2405 (O_2405,N_19601,N_19086);
or UO_2406 (O_2406,N_19028,N_19301);
xor UO_2407 (O_2407,N_19862,N_19145);
and UO_2408 (O_2408,N_19879,N_19018);
or UO_2409 (O_2409,N_19449,N_19454);
xor UO_2410 (O_2410,N_19346,N_19937);
and UO_2411 (O_2411,N_19811,N_19528);
or UO_2412 (O_2412,N_19012,N_19785);
and UO_2413 (O_2413,N_19998,N_19853);
nand UO_2414 (O_2414,N_19672,N_19088);
or UO_2415 (O_2415,N_19026,N_19258);
or UO_2416 (O_2416,N_19716,N_19560);
xor UO_2417 (O_2417,N_19386,N_19442);
or UO_2418 (O_2418,N_19532,N_19889);
and UO_2419 (O_2419,N_19836,N_19389);
and UO_2420 (O_2420,N_19904,N_19471);
nand UO_2421 (O_2421,N_19931,N_19975);
nor UO_2422 (O_2422,N_19639,N_19950);
xnor UO_2423 (O_2423,N_19998,N_19658);
xor UO_2424 (O_2424,N_19013,N_19336);
nor UO_2425 (O_2425,N_19322,N_19701);
nand UO_2426 (O_2426,N_19699,N_19936);
and UO_2427 (O_2427,N_19429,N_19276);
nor UO_2428 (O_2428,N_19995,N_19782);
nor UO_2429 (O_2429,N_19741,N_19255);
nor UO_2430 (O_2430,N_19692,N_19754);
and UO_2431 (O_2431,N_19304,N_19442);
or UO_2432 (O_2432,N_19441,N_19431);
and UO_2433 (O_2433,N_19171,N_19274);
nand UO_2434 (O_2434,N_19076,N_19233);
and UO_2435 (O_2435,N_19208,N_19813);
and UO_2436 (O_2436,N_19895,N_19078);
or UO_2437 (O_2437,N_19845,N_19793);
and UO_2438 (O_2438,N_19530,N_19476);
xnor UO_2439 (O_2439,N_19059,N_19609);
and UO_2440 (O_2440,N_19036,N_19622);
nor UO_2441 (O_2441,N_19316,N_19814);
or UO_2442 (O_2442,N_19406,N_19889);
xnor UO_2443 (O_2443,N_19332,N_19667);
nand UO_2444 (O_2444,N_19723,N_19479);
and UO_2445 (O_2445,N_19172,N_19443);
or UO_2446 (O_2446,N_19370,N_19738);
or UO_2447 (O_2447,N_19181,N_19663);
or UO_2448 (O_2448,N_19450,N_19607);
nor UO_2449 (O_2449,N_19478,N_19293);
nand UO_2450 (O_2450,N_19567,N_19801);
and UO_2451 (O_2451,N_19893,N_19433);
nor UO_2452 (O_2452,N_19081,N_19543);
nand UO_2453 (O_2453,N_19235,N_19912);
and UO_2454 (O_2454,N_19709,N_19151);
or UO_2455 (O_2455,N_19098,N_19725);
nand UO_2456 (O_2456,N_19336,N_19317);
or UO_2457 (O_2457,N_19178,N_19715);
and UO_2458 (O_2458,N_19732,N_19267);
and UO_2459 (O_2459,N_19590,N_19177);
xnor UO_2460 (O_2460,N_19401,N_19788);
xnor UO_2461 (O_2461,N_19499,N_19349);
xor UO_2462 (O_2462,N_19925,N_19329);
nor UO_2463 (O_2463,N_19674,N_19930);
and UO_2464 (O_2464,N_19425,N_19221);
nand UO_2465 (O_2465,N_19298,N_19608);
or UO_2466 (O_2466,N_19506,N_19511);
or UO_2467 (O_2467,N_19060,N_19936);
or UO_2468 (O_2468,N_19447,N_19017);
or UO_2469 (O_2469,N_19868,N_19115);
xor UO_2470 (O_2470,N_19344,N_19729);
nor UO_2471 (O_2471,N_19694,N_19202);
nand UO_2472 (O_2472,N_19334,N_19993);
and UO_2473 (O_2473,N_19468,N_19131);
nor UO_2474 (O_2474,N_19634,N_19289);
nor UO_2475 (O_2475,N_19242,N_19720);
or UO_2476 (O_2476,N_19816,N_19478);
xnor UO_2477 (O_2477,N_19383,N_19149);
and UO_2478 (O_2478,N_19746,N_19041);
xnor UO_2479 (O_2479,N_19950,N_19566);
nor UO_2480 (O_2480,N_19980,N_19546);
or UO_2481 (O_2481,N_19144,N_19637);
xnor UO_2482 (O_2482,N_19422,N_19015);
xnor UO_2483 (O_2483,N_19252,N_19063);
xnor UO_2484 (O_2484,N_19350,N_19358);
and UO_2485 (O_2485,N_19621,N_19342);
nand UO_2486 (O_2486,N_19103,N_19153);
and UO_2487 (O_2487,N_19198,N_19693);
or UO_2488 (O_2488,N_19960,N_19948);
nor UO_2489 (O_2489,N_19306,N_19437);
nor UO_2490 (O_2490,N_19983,N_19460);
xor UO_2491 (O_2491,N_19265,N_19201);
xnor UO_2492 (O_2492,N_19883,N_19171);
xnor UO_2493 (O_2493,N_19052,N_19653);
or UO_2494 (O_2494,N_19216,N_19465);
nand UO_2495 (O_2495,N_19407,N_19398);
or UO_2496 (O_2496,N_19399,N_19250);
or UO_2497 (O_2497,N_19626,N_19426);
nor UO_2498 (O_2498,N_19464,N_19387);
or UO_2499 (O_2499,N_19721,N_19320);
endmodule