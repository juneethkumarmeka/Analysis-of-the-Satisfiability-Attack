module basic_500_3000_500_15_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_334,In_178);
xor U1 (N_1,In_216,In_346);
and U2 (N_2,In_390,In_348);
nand U3 (N_3,In_62,In_384);
and U4 (N_4,In_222,In_258);
nor U5 (N_5,In_380,In_399);
and U6 (N_6,In_61,In_293);
xor U7 (N_7,In_459,In_423);
or U8 (N_8,In_12,In_377);
nand U9 (N_9,In_96,In_357);
and U10 (N_10,In_137,In_217);
or U11 (N_11,In_259,In_197);
or U12 (N_12,In_337,In_44);
and U13 (N_13,In_382,In_246);
xnor U14 (N_14,In_243,In_455);
xnor U15 (N_15,In_34,In_430);
xor U16 (N_16,In_299,In_283);
and U17 (N_17,In_14,In_33);
and U18 (N_18,In_84,In_461);
xnor U19 (N_19,In_170,In_465);
nor U20 (N_20,In_129,In_195);
and U21 (N_21,In_238,In_172);
nand U22 (N_22,In_495,In_328);
or U23 (N_23,In_98,In_394);
nor U24 (N_24,In_302,In_231);
and U25 (N_25,In_429,In_119);
nor U26 (N_26,In_150,In_444);
nor U27 (N_27,In_60,In_58);
and U28 (N_28,In_426,In_57);
nand U29 (N_29,In_467,In_385);
nand U30 (N_30,In_28,In_145);
or U31 (N_31,In_166,In_341);
or U32 (N_32,In_305,In_225);
nand U33 (N_33,In_406,In_181);
nand U34 (N_34,In_374,In_250);
and U35 (N_35,In_412,In_144);
and U36 (N_36,In_351,In_474);
or U37 (N_37,In_221,In_26);
and U38 (N_38,In_48,In_453);
nor U39 (N_39,In_372,In_127);
nor U40 (N_40,In_173,In_1);
xnor U41 (N_41,In_497,In_253);
and U42 (N_42,In_239,In_236);
nand U43 (N_43,In_428,In_92);
xnor U44 (N_44,In_274,In_148);
nor U45 (N_45,In_440,In_151);
nand U46 (N_46,In_395,In_114);
and U47 (N_47,In_322,In_469);
nand U48 (N_48,In_248,In_138);
xnor U49 (N_49,In_358,In_121);
and U50 (N_50,In_229,In_392);
nor U51 (N_51,In_408,In_464);
xnor U52 (N_52,In_86,In_130);
nor U53 (N_53,In_403,In_280);
and U54 (N_54,In_198,In_165);
nand U55 (N_55,In_203,In_109);
xor U56 (N_56,In_163,In_23);
or U57 (N_57,In_20,In_366);
xor U58 (N_58,In_191,In_208);
nor U59 (N_59,In_164,In_344);
or U60 (N_60,In_95,In_448);
or U61 (N_61,In_100,In_261);
xor U62 (N_62,In_257,In_269);
and U63 (N_63,In_209,In_458);
or U64 (N_64,In_436,In_18);
and U65 (N_65,In_79,In_157);
nor U66 (N_66,In_364,In_370);
or U67 (N_67,In_213,In_468);
nand U68 (N_68,In_45,In_482);
nand U69 (N_69,In_398,In_146);
nor U70 (N_70,In_271,In_445);
nor U71 (N_71,In_402,In_397);
and U72 (N_72,In_111,In_211);
nand U73 (N_73,In_128,In_228);
nand U74 (N_74,In_36,In_386);
xnor U75 (N_75,In_381,In_207);
and U76 (N_76,In_296,In_49);
xor U77 (N_77,In_363,In_289);
and U78 (N_78,In_477,In_192);
nand U79 (N_79,In_53,In_347);
and U80 (N_80,In_488,In_227);
or U81 (N_81,In_407,In_319);
nand U82 (N_82,In_316,In_156);
xnor U83 (N_83,In_264,In_187);
or U84 (N_84,In_69,In_443);
nor U85 (N_85,In_471,In_354);
xor U86 (N_86,In_65,In_241);
or U87 (N_87,In_290,In_291);
or U88 (N_88,In_105,In_438);
and U89 (N_89,In_184,In_282);
nor U90 (N_90,In_244,In_484);
nand U91 (N_91,In_416,In_303);
nand U92 (N_92,In_162,In_94);
and U93 (N_93,In_204,In_133);
xnor U94 (N_94,In_159,In_498);
xor U95 (N_95,In_215,In_277);
xor U96 (N_96,In_55,In_169);
xor U97 (N_97,In_63,In_460);
xor U98 (N_98,In_186,In_107);
xnor U99 (N_99,In_410,In_494);
nor U100 (N_100,In_219,In_214);
and U101 (N_101,In_76,In_292);
nand U102 (N_102,In_155,In_233);
and U103 (N_103,In_249,In_450);
nand U104 (N_104,In_175,In_131);
and U105 (N_105,In_67,In_251);
nor U106 (N_106,In_147,In_330);
nor U107 (N_107,In_185,In_124);
nor U108 (N_108,In_457,In_353);
xnor U109 (N_109,In_19,In_311);
nor U110 (N_110,In_417,In_383);
nand U111 (N_111,In_401,In_281);
or U112 (N_112,In_273,In_476);
nor U113 (N_113,In_240,In_335);
or U114 (N_114,In_87,In_242);
xor U115 (N_115,In_441,In_327);
and U116 (N_116,In_409,In_182);
or U117 (N_117,In_224,In_349);
nor U118 (N_118,In_83,In_350);
nor U119 (N_119,In_85,In_356);
and U120 (N_120,In_89,In_266);
nand U121 (N_121,In_78,In_93);
nand U122 (N_122,In_134,In_325);
nor U123 (N_123,In_326,In_201);
nand U124 (N_124,In_110,In_15);
and U125 (N_125,In_493,In_125);
or U126 (N_126,In_359,In_309);
nand U127 (N_127,In_143,In_449);
nor U128 (N_128,In_345,In_489);
xnor U129 (N_129,In_220,In_252);
and U130 (N_130,In_480,In_499);
nor U131 (N_131,In_340,In_490);
nand U132 (N_132,In_71,In_177);
xor U133 (N_133,In_483,In_263);
nand U134 (N_134,In_6,In_415);
or U135 (N_135,In_492,In_140);
xor U136 (N_136,In_254,In_446);
nor U137 (N_137,In_210,In_22);
xor U138 (N_138,In_64,In_31);
or U139 (N_139,In_320,In_82);
and U140 (N_140,In_24,In_161);
and U141 (N_141,In_310,In_25);
or U142 (N_142,In_168,In_388);
and U143 (N_143,In_434,In_59);
nand U144 (N_144,In_142,In_400);
and U145 (N_145,In_424,In_314);
or U146 (N_146,In_27,In_376);
nand U147 (N_147,In_362,In_46);
xnor U148 (N_148,In_278,In_75);
or U149 (N_149,In_411,In_135);
and U150 (N_150,In_245,In_90);
nor U151 (N_151,In_331,In_152);
xnor U152 (N_152,In_387,In_132);
xnor U153 (N_153,In_315,In_432);
and U154 (N_154,In_452,In_112);
nor U155 (N_155,In_226,In_307);
nor U156 (N_156,In_43,In_439);
and U157 (N_157,In_37,In_300);
and U158 (N_158,In_42,In_205);
nand U159 (N_159,In_174,In_268);
xor U160 (N_160,In_389,In_115);
or U161 (N_161,In_478,In_0);
nor U162 (N_162,In_262,In_39);
nor U163 (N_163,In_295,In_223);
nor U164 (N_164,In_183,In_265);
nand U165 (N_165,In_88,In_312);
nand U166 (N_166,In_126,In_496);
and U167 (N_167,In_431,In_272);
or U168 (N_168,In_149,In_120);
nand U169 (N_169,In_237,In_102);
nand U170 (N_170,In_367,In_196);
or U171 (N_171,In_371,In_396);
and U172 (N_172,In_435,In_267);
nand U173 (N_173,In_103,In_433);
and U174 (N_174,In_454,In_206);
nand U175 (N_175,In_17,In_475);
and U176 (N_176,In_306,In_10);
nand U177 (N_177,In_301,In_297);
xor U178 (N_178,In_160,In_118);
nor U179 (N_179,In_180,In_355);
and U180 (N_180,In_72,In_442);
nor U181 (N_181,In_50,In_365);
and U182 (N_182,In_324,In_479);
xor U183 (N_183,In_232,In_481);
nand U184 (N_184,In_422,In_418);
nor U185 (N_185,In_9,In_329);
nor U186 (N_186,In_451,In_4);
nand U187 (N_187,In_286,In_97);
nand U188 (N_188,In_167,In_190);
nor U189 (N_189,In_323,In_285);
nand U190 (N_190,In_141,In_139);
nor U191 (N_191,In_466,In_360);
xnor U192 (N_192,In_279,In_379);
and U193 (N_193,In_470,In_101);
or U194 (N_194,In_38,In_485);
nand U195 (N_195,In_463,In_317);
nor U196 (N_196,In_2,In_373);
or U197 (N_197,In_113,In_73);
xor U198 (N_198,In_462,In_193);
and U199 (N_199,In_158,In_29);
and U200 (N_200,N_64,N_93);
or U201 (N_201,N_48,N_0);
and U202 (N_202,N_171,In_106);
or U203 (N_203,In_419,In_298);
and U204 (N_204,N_114,In_56);
nor U205 (N_205,N_174,In_393);
nor U206 (N_206,N_123,N_19);
xor U207 (N_207,N_41,In_66);
nand U208 (N_208,N_84,In_80);
nor U209 (N_209,N_58,N_185);
or U210 (N_210,In_3,In_425);
and U211 (N_211,N_148,N_132);
xnor U212 (N_212,In_342,In_234);
or U213 (N_213,In_321,In_437);
xnor U214 (N_214,N_79,N_140);
xnor U215 (N_215,N_97,N_29);
nand U216 (N_216,N_74,N_151);
and U217 (N_217,In_487,In_473);
xnor U218 (N_218,In_7,N_89);
or U219 (N_219,In_308,N_181);
and U220 (N_220,In_154,In_391);
nand U221 (N_221,In_343,N_178);
nor U222 (N_222,In_116,N_176);
or U223 (N_223,N_91,In_194);
or U224 (N_224,N_16,In_153);
nor U225 (N_225,N_38,In_47);
nand U226 (N_226,N_86,N_158);
xnor U227 (N_227,In_288,N_184);
xnor U228 (N_228,N_197,In_421);
nor U229 (N_229,N_157,In_54);
or U230 (N_230,N_12,N_83);
and U231 (N_231,In_447,In_200);
nand U232 (N_232,N_166,N_156);
xnor U233 (N_233,In_336,In_81);
or U234 (N_234,N_133,N_199);
or U235 (N_235,N_116,N_73);
or U236 (N_236,In_294,In_230);
nor U237 (N_237,N_179,N_60);
xor U238 (N_238,N_44,N_31);
or U239 (N_239,N_160,In_136);
xnor U240 (N_240,N_59,In_404);
xor U241 (N_241,N_105,In_270);
or U242 (N_242,N_106,N_126);
and U243 (N_243,In_5,In_212);
and U244 (N_244,N_152,N_71);
nand U245 (N_245,N_183,N_68);
or U246 (N_246,N_57,N_117);
xor U247 (N_247,N_78,In_104);
nand U248 (N_248,N_66,In_11);
and U249 (N_249,N_17,N_146);
and U250 (N_250,N_175,N_144);
and U251 (N_251,N_62,In_369);
and U252 (N_252,In_117,N_32);
xor U253 (N_253,N_121,In_472);
or U254 (N_254,N_145,In_99);
nand U255 (N_255,N_108,N_170);
or U256 (N_256,N_23,N_168);
and U257 (N_257,N_139,N_112);
xnor U258 (N_258,N_136,In_333);
or U259 (N_259,N_150,N_3);
or U260 (N_260,In_40,N_186);
or U261 (N_261,N_167,N_124);
and U262 (N_262,N_163,N_180);
xnor U263 (N_263,In_260,N_165);
or U264 (N_264,N_120,N_43);
and U265 (N_265,N_103,N_128);
or U266 (N_266,N_77,N_10);
nand U267 (N_267,N_76,N_143);
and U268 (N_268,N_72,N_21);
nor U269 (N_269,N_154,N_159);
nand U270 (N_270,N_22,N_53);
and U271 (N_271,N_4,In_199);
or U272 (N_272,N_70,In_332);
and U273 (N_273,N_194,N_26);
nand U274 (N_274,N_164,In_304);
or U275 (N_275,N_192,In_91);
and U276 (N_276,In_255,N_15);
nand U277 (N_277,N_107,N_118);
xor U278 (N_278,N_188,N_111);
or U279 (N_279,In_287,N_40);
and U280 (N_280,N_127,N_11);
or U281 (N_281,N_63,In_313);
and U282 (N_282,N_90,In_51);
xnor U283 (N_283,N_65,N_162);
nand U284 (N_284,N_135,N_96);
nor U285 (N_285,In_427,N_113);
and U286 (N_286,N_52,N_5);
nand U287 (N_287,In_35,N_45);
or U288 (N_288,In_420,N_2);
nand U289 (N_289,N_189,N_34);
and U290 (N_290,N_191,In_179);
and U291 (N_291,In_13,N_131);
nor U292 (N_292,N_39,In_284);
nand U293 (N_293,N_24,N_18);
nor U294 (N_294,In_202,N_155);
nor U295 (N_295,N_33,N_102);
nor U296 (N_296,In_171,In_77);
xor U297 (N_297,In_108,N_14);
nor U298 (N_298,N_30,N_94);
nor U299 (N_299,In_189,N_198);
xnor U300 (N_300,N_50,N_100);
xnor U301 (N_301,N_28,In_256);
nand U302 (N_302,In_375,N_85);
xnor U303 (N_303,N_6,In_235);
and U304 (N_304,In_247,N_149);
nand U305 (N_305,N_13,N_37);
nor U306 (N_306,N_187,In_123);
nand U307 (N_307,N_153,N_1);
and U308 (N_308,In_218,In_21);
or U309 (N_309,N_47,N_104);
xor U310 (N_310,N_177,In_70);
nand U311 (N_311,N_75,N_8);
or U312 (N_312,N_54,In_52);
nand U313 (N_313,N_49,N_98);
xnor U314 (N_314,N_25,N_69);
nand U315 (N_315,In_30,N_119);
and U316 (N_316,In_486,N_195);
and U317 (N_317,N_61,N_27);
and U318 (N_318,N_92,N_110);
or U319 (N_319,In_68,N_129);
nor U320 (N_320,In_352,N_138);
nor U321 (N_321,In_378,N_142);
nor U322 (N_322,In_276,N_87);
or U323 (N_323,In_405,N_196);
and U324 (N_324,N_169,N_80);
or U325 (N_325,N_122,N_125);
and U326 (N_326,N_46,N_101);
or U327 (N_327,N_99,In_16);
xnor U328 (N_328,In_491,In_368);
xor U329 (N_329,In_413,In_318);
or U330 (N_330,N_193,N_42);
or U331 (N_331,N_147,In_414);
or U332 (N_332,In_8,In_338);
xnor U333 (N_333,In_456,N_172);
xnor U334 (N_334,N_109,N_35);
and U335 (N_335,N_137,N_115);
nor U336 (N_336,N_9,N_55);
nand U337 (N_337,N_88,N_81);
xnor U338 (N_338,N_173,In_339);
nor U339 (N_339,N_134,N_182);
nor U340 (N_340,N_141,In_122);
nand U341 (N_341,In_32,In_275);
nor U342 (N_342,N_130,In_361);
nand U343 (N_343,In_176,In_74);
and U344 (N_344,N_67,N_56);
xor U345 (N_345,N_7,In_188);
nor U346 (N_346,N_190,In_41);
xnor U347 (N_347,N_95,N_20);
or U348 (N_348,N_161,N_36);
xor U349 (N_349,N_51,N_82);
or U350 (N_350,In_393,In_425);
xnor U351 (N_351,In_420,N_133);
and U352 (N_352,N_26,N_29);
xnor U353 (N_353,In_66,N_2);
nand U354 (N_354,In_375,In_104);
or U355 (N_355,N_74,N_47);
nor U356 (N_356,In_491,In_339);
and U357 (N_357,N_76,N_82);
and U358 (N_358,N_136,N_91);
or U359 (N_359,N_54,N_157);
nand U360 (N_360,N_102,N_93);
and U361 (N_361,N_42,N_176);
xnor U362 (N_362,In_212,In_276);
and U363 (N_363,N_126,In_104);
or U364 (N_364,N_142,In_352);
and U365 (N_365,N_32,N_79);
nor U366 (N_366,N_0,N_17);
and U367 (N_367,In_11,N_161);
nor U368 (N_368,In_421,N_62);
and U369 (N_369,In_375,In_136);
and U370 (N_370,In_472,N_35);
nor U371 (N_371,N_76,N_39);
nor U372 (N_372,N_101,N_68);
nor U373 (N_373,In_393,In_420);
xor U374 (N_374,N_144,N_75);
nor U375 (N_375,N_42,In_414);
nor U376 (N_376,N_137,N_23);
nand U377 (N_377,N_37,N_112);
or U378 (N_378,In_200,N_161);
or U379 (N_379,N_39,N_171);
nand U380 (N_380,N_26,In_425);
nand U381 (N_381,N_108,In_338);
nand U382 (N_382,In_333,N_101);
and U383 (N_383,In_419,N_11);
and U384 (N_384,N_59,N_198);
or U385 (N_385,In_313,N_7);
nand U386 (N_386,In_40,N_182);
or U387 (N_387,In_108,N_127);
nor U388 (N_388,N_4,In_136);
nor U389 (N_389,N_19,In_275);
or U390 (N_390,N_80,N_124);
or U391 (N_391,N_170,In_338);
xnor U392 (N_392,N_10,In_343);
nor U393 (N_393,N_46,N_164);
and U394 (N_394,In_154,In_473);
nor U395 (N_395,N_14,In_420);
nor U396 (N_396,N_63,In_342);
or U397 (N_397,In_276,In_32);
xor U398 (N_398,In_8,N_67);
xnor U399 (N_399,N_134,N_158);
nand U400 (N_400,N_206,N_328);
nand U401 (N_401,N_315,N_281);
xor U402 (N_402,N_360,N_336);
nand U403 (N_403,N_271,N_323);
nor U404 (N_404,N_361,N_290);
xor U405 (N_405,N_355,N_385);
and U406 (N_406,N_218,N_215);
or U407 (N_407,N_257,N_300);
and U408 (N_408,N_248,N_238);
or U409 (N_409,N_354,N_217);
or U410 (N_410,N_204,N_251);
or U411 (N_411,N_280,N_371);
nor U412 (N_412,N_203,N_283);
xnor U413 (N_413,N_298,N_252);
and U414 (N_414,N_369,N_239);
or U415 (N_415,N_229,N_324);
xnor U416 (N_416,N_382,N_249);
nand U417 (N_417,N_207,N_347);
and U418 (N_418,N_307,N_234);
xor U419 (N_419,N_295,N_380);
nand U420 (N_420,N_396,N_210);
or U421 (N_421,N_353,N_241);
xnor U422 (N_422,N_244,N_235);
xnor U423 (N_423,N_208,N_368);
xor U424 (N_424,N_224,N_306);
nor U425 (N_425,N_391,N_386);
nand U426 (N_426,N_263,N_351);
or U427 (N_427,N_225,N_376);
and U428 (N_428,N_265,N_329);
or U429 (N_429,N_387,N_284);
or U430 (N_430,N_213,N_335);
or U431 (N_431,N_250,N_350);
and U432 (N_432,N_321,N_322);
xor U433 (N_433,N_237,N_264);
xor U434 (N_434,N_358,N_375);
nor U435 (N_435,N_258,N_201);
nand U436 (N_436,N_236,N_344);
nand U437 (N_437,N_221,N_256);
nand U438 (N_438,N_342,N_395);
nor U439 (N_439,N_326,N_331);
nor U440 (N_440,N_373,N_392);
nor U441 (N_441,N_273,N_231);
nor U442 (N_442,N_319,N_318);
nand U443 (N_443,N_296,N_266);
or U444 (N_444,N_289,N_363);
xnor U445 (N_445,N_200,N_366);
or U446 (N_446,N_209,N_339);
nand U447 (N_447,N_245,N_294);
and U448 (N_448,N_383,N_381);
and U449 (N_449,N_352,N_243);
and U450 (N_450,N_349,N_356);
nand U451 (N_451,N_365,N_216);
or U452 (N_452,N_254,N_228);
nor U453 (N_453,N_338,N_230);
nor U454 (N_454,N_285,N_359);
nand U455 (N_455,N_379,N_345);
and U456 (N_456,N_212,N_222);
xor U457 (N_457,N_348,N_211);
xor U458 (N_458,N_388,N_279);
xnor U459 (N_459,N_316,N_370);
or U460 (N_460,N_275,N_374);
xnor U461 (N_461,N_292,N_327);
xor U462 (N_462,N_276,N_297);
or U463 (N_463,N_367,N_320);
nor U464 (N_464,N_260,N_202);
xor U465 (N_465,N_269,N_364);
nand U466 (N_466,N_384,N_310);
nand U467 (N_467,N_286,N_325);
xnor U468 (N_468,N_311,N_261);
nand U469 (N_469,N_233,N_301);
xor U470 (N_470,N_278,N_220);
or U471 (N_471,N_268,N_343);
nor U472 (N_472,N_226,N_274);
nand U473 (N_473,N_346,N_399);
xnor U474 (N_474,N_313,N_389);
nor U475 (N_475,N_272,N_255);
nor U476 (N_476,N_390,N_397);
or U477 (N_477,N_372,N_219);
nor U478 (N_478,N_393,N_314);
or U479 (N_479,N_253,N_240);
xor U480 (N_480,N_398,N_247);
or U481 (N_481,N_317,N_259);
nor U482 (N_482,N_357,N_232);
or U483 (N_483,N_333,N_277);
or U484 (N_484,N_341,N_246);
nand U485 (N_485,N_377,N_332);
nand U486 (N_486,N_205,N_288);
and U487 (N_487,N_291,N_302);
and U488 (N_488,N_227,N_312);
nand U489 (N_489,N_287,N_270);
xnor U490 (N_490,N_223,N_309);
or U491 (N_491,N_214,N_282);
nand U492 (N_492,N_308,N_267);
nor U493 (N_493,N_337,N_362);
nand U494 (N_494,N_340,N_293);
nor U495 (N_495,N_330,N_304);
and U496 (N_496,N_299,N_262);
or U497 (N_497,N_394,N_303);
or U498 (N_498,N_305,N_334);
and U499 (N_499,N_242,N_378);
or U500 (N_500,N_329,N_246);
nand U501 (N_501,N_328,N_393);
nand U502 (N_502,N_209,N_326);
xor U503 (N_503,N_268,N_222);
xnor U504 (N_504,N_239,N_262);
nand U505 (N_505,N_201,N_318);
nor U506 (N_506,N_301,N_261);
or U507 (N_507,N_221,N_288);
xnor U508 (N_508,N_236,N_377);
nor U509 (N_509,N_240,N_319);
or U510 (N_510,N_314,N_329);
nand U511 (N_511,N_332,N_334);
xnor U512 (N_512,N_210,N_355);
and U513 (N_513,N_207,N_213);
xnor U514 (N_514,N_220,N_398);
or U515 (N_515,N_209,N_213);
or U516 (N_516,N_365,N_346);
or U517 (N_517,N_342,N_283);
or U518 (N_518,N_359,N_244);
and U519 (N_519,N_271,N_233);
xnor U520 (N_520,N_287,N_341);
or U521 (N_521,N_223,N_287);
and U522 (N_522,N_246,N_322);
nor U523 (N_523,N_353,N_293);
nor U524 (N_524,N_348,N_385);
nand U525 (N_525,N_390,N_366);
xor U526 (N_526,N_218,N_327);
nor U527 (N_527,N_336,N_320);
and U528 (N_528,N_341,N_223);
xor U529 (N_529,N_265,N_392);
nand U530 (N_530,N_295,N_253);
xnor U531 (N_531,N_389,N_207);
nand U532 (N_532,N_245,N_212);
nor U533 (N_533,N_362,N_288);
xor U534 (N_534,N_260,N_282);
nand U535 (N_535,N_309,N_355);
xor U536 (N_536,N_281,N_218);
and U537 (N_537,N_269,N_215);
or U538 (N_538,N_313,N_332);
and U539 (N_539,N_365,N_280);
or U540 (N_540,N_276,N_323);
and U541 (N_541,N_231,N_368);
or U542 (N_542,N_253,N_382);
xor U543 (N_543,N_240,N_264);
and U544 (N_544,N_323,N_380);
xor U545 (N_545,N_293,N_266);
and U546 (N_546,N_218,N_283);
nand U547 (N_547,N_298,N_248);
nor U548 (N_548,N_274,N_346);
nor U549 (N_549,N_291,N_307);
or U550 (N_550,N_346,N_364);
nand U551 (N_551,N_339,N_203);
nand U552 (N_552,N_256,N_302);
nand U553 (N_553,N_240,N_392);
or U554 (N_554,N_380,N_275);
and U555 (N_555,N_345,N_304);
nand U556 (N_556,N_399,N_335);
or U557 (N_557,N_322,N_250);
xnor U558 (N_558,N_206,N_359);
nand U559 (N_559,N_315,N_267);
or U560 (N_560,N_314,N_237);
or U561 (N_561,N_235,N_207);
and U562 (N_562,N_220,N_207);
xor U563 (N_563,N_376,N_200);
nor U564 (N_564,N_256,N_388);
nor U565 (N_565,N_220,N_366);
or U566 (N_566,N_258,N_367);
xnor U567 (N_567,N_265,N_266);
nand U568 (N_568,N_283,N_303);
nand U569 (N_569,N_225,N_325);
nand U570 (N_570,N_362,N_248);
nand U571 (N_571,N_208,N_302);
nand U572 (N_572,N_343,N_240);
nand U573 (N_573,N_280,N_372);
xor U574 (N_574,N_375,N_267);
nor U575 (N_575,N_392,N_216);
nand U576 (N_576,N_343,N_229);
and U577 (N_577,N_286,N_274);
and U578 (N_578,N_255,N_372);
xor U579 (N_579,N_335,N_397);
or U580 (N_580,N_361,N_364);
nor U581 (N_581,N_247,N_305);
nor U582 (N_582,N_316,N_392);
nor U583 (N_583,N_299,N_276);
and U584 (N_584,N_224,N_343);
and U585 (N_585,N_314,N_339);
xnor U586 (N_586,N_399,N_343);
nand U587 (N_587,N_205,N_316);
or U588 (N_588,N_355,N_254);
nor U589 (N_589,N_208,N_304);
xnor U590 (N_590,N_200,N_257);
nor U591 (N_591,N_331,N_268);
nor U592 (N_592,N_221,N_273);
or U593 (N_593,N_258,N_371);
xor U594 (N_594,N_247,N_266);
nor U595 (N_595,N_321,N_320);
xor U596 (N_596,N_376,N_306);
and U597 (N_597,N_225,N_366);
and U598 (N_598,N_257,N_298);
nand U599 (N_599,N_255,N_300);
nand U600 (N_600,N_440,N_401);
nand U601 (N_601,N_489,N_424);
xnor U602 (N_602,N_455,N_415);
and U603 (N_603,N_533,N_487);
xor U604 (N_604,N_507,N_523);
nor U605 (N_605,N_594,N_555);
nand U606 (N_606,N_568,N_571);
xor U607 (N_607,N_579,N_536);
or U608 (N_608,N_505,N_532);
and U609 (N_609,N_477,N_509);
and U610 (N_610,N_495,N_491);
nand U611 (N_611,N_547,N_427);
and U612 (N_612,N_546,N_479);
nor U613 (N_613,N_451,N_432);
or U614 (N_614,N_552,N_482);
or U615 (N_615,N_410,N_591);
nor U616 (N_616,N_599,N_416);
and U617 (N_617,N_537,N_483);
and U618 (N_618,N_405,N_544);
or U619 (N_619,N_428,N_434);
and U620 (N_620,N_412,N_452);
nand U621 (N_621,N_459,N_450);
nand U622 (N_622,N_462,N_444);
xor U623 (N_623,N_549,N_504);
nand U624 (N_624,N_551,N_540);
and U625 (N_625,N_496,N_402);
nand U626 (N_626,N_562,N_461);
and U627 (N_627,N_525,N_473);
or U628 (N_628,N_511,N_460);
nand U629 (N_629,N_583,N_430);
xor U630 (N_630,N_590,N_560);
nand U631 (N_631,N_439,N_485);
xor U632 (N_632,N_519,N_570);
and U633 (N_633,N_500,N_408);
or U634 (N_634,N_472,N_515);
xor U635 (N_635,N_518,N_480);
xor U636 (N_636,N_573,N_466);
or U637 (N_637,N_596,N_403);
nor U638 (N_638,N_567,N_443);
xnor U639 (N_639,N_543,N_464);
nor U640 (N_640,N_513,N_565);
xor U641 (N_641,N_510,N_458);
xnor U642 (N_642,N_446,N_529);
nand U643 (N_643,N_490,N_463);
or U644 (N_644,N_413,N_441);
nand U645 (N_645,N_569,N_447);
nand U646 (N_646,N_431,N_512);
nor U647 (N_647,N_425,N_524);
xor U648 (N_648,N_556,N_531);
nor U649 (N_649,N_597,N_584);
or U650 (N_650,N_494,N_557);
and U651 (N_651,N_577,N_453);
nand U652 (N_652,N_488,N_474);
or U653 (N_653,N_582,N_575);
nor U654 (N_654,N_417,N_498);
and U655 (N_655,N_420,N_553);
and U656 (N_656,N_506,N_429);
and U657 (N_657,N_528,N_437);
nand U658 (N_658,N_574,N_442);
xor U659 (N_659,N_470,N_469);
xor U660 (N_660,N_542,N_419);
xnor U661 (N_661,N_404,N_433);
or U662 (N_662,N_559,N_400);
or U663 (N_663,N_576,N_465);
xnor U664 (N_664,N_521,N_445);
xor U665 (N_665,N_406,N_407);
or U666 (N_666,N_527,N_436);
nor U667 (N_667,N_508,N_592);
and U668 (N_668,N_486,N_564);
or U669 (N_669,N_554,N_548);
nand U670 (N_670,N_448,N_426);
nand U671 (N_671,N_438,N_520);
or U672 (N_672,N_539,N_499);
and U673 (N_673,N_456,N_421);
nand U674 (N_674,N_572,N_476);
xor U675 (N_675,N_538,N_481);
nor U676 (N_676,N_418,N_435);
or U677 (N_677,N_545,N_586);
xnor U678 (N_678,N_561,N_475);
nor U679 (N_679,N_535,N_422);
xor U680 (N_680,N_516,N_514);
nor U681 (N_681,N_468,N_457);
and U682 (N_682,N_580,N_409);
and U683 (N_683,N_526,N_522);
nor U684 (N_684,N_411,N_578);
or U685 (N_685,N_593,N_414);
or U686 (N_686,N_478,N_471);
and U687 (N_687,N_566,N_497);
nand U688 (N_688,N_587,N_595);
or U689 (N_689,N_588,N_467);
nand U690 (N_690,N_598,N_484);
nor U691 (N_691,N_541,N_530);
nand U692 (N_692,N_589,N_503);
or U693 (N_693,N_492,N_563);
nor U694 (N_694,N_585,N_501);
and U695 (N_695,N_493,N_550);
or U696 (N_696,N_454,N_534);
or U697 (N_697,N_558,N_581);
xor U698 (N_698,N_423,N_517);
nor U699 (N_699,N_502,N_449);
nand U700 (N_700,N_464,N_404);
nor U701 (N_701,N_564,N_573);
xor U702 (N_702,N_423,N_594);
nand U703 (N_703,N_452,N_560);
nor U704 (N_704,N_458,N_489);
or U705 (N_705,N_413,N_474);
nand U706 (N_706,N_449,N_585);
or U707 (N_707,N_484,N_563);
nand U708 (N_708,N_475,N_405);
xnor U709 (N_709,N_400,N_543);
and U710 (N_710,N_514,N_510);
xnor U711 (N_711,N_566,N_563);
and U712 (N_712,N_462,N_531);
or U713 (N_713,N_491,N_484);
and U714 (N_714,N_557,N_421);
nand U715 (N_715,N_562,N_496);
xnor U716 (N_716,N_497,N_599);
xnor U717 (N_717,N_548,N_514);
or U718 (N_718,N_435,N_447);
nand U719 (N_719,N_513,N_416);
nor U720 (N_720,N_533,N_523);
and U721 (N_721,N_414,N_518);
or U722 (N_722,N_410,N_570);
xnor U723 (N_723,N_428,N_551);
or U724 (N_724,N_447,N_514);
and U725 (N_725,N_502,N_554);
or U726 (N_726,N_407,N_573);
nor U727 (N_727,N_555,N_556);
nor U728 (N_728,N_587,N_596);
xor U729 (N_729,N_438,N_412);
or U730 (N_730,N_424,N_468);
nand U731 (N_731,N_529,N_516);
xor U732 (N_732,N_403,N_412);
or U733 (N_733,N_534,N_596);
or U734 (N_734,N_581,N_439);
or U735 (N_735,N_513,N_492);
nand U736 (N_736,N_470,N_467);
nand U737 (N_737,N_442,N_490);
and U738 (N_738,N_423,N_448);
or U739 (N_739,N_474,N_457);
nor U740 (N_740,N_498,N_489);
or U741 (N_741,N_420,N_518);
nand U742 (N_742,N_529,N_530);
nand U743 (N_743,N_457,N_592);
or U744 (N_744,N_467,N_595);
xor U745 (N_745,N_452,N_521);
or U746 (N_746,N_426,N_540);
nor U747 (N_747,N_439,N_440);
nand U748 (N_748,N_560,N_592);
nand U749 (N_749,N_503,N_442);
or U750 (N_750,N_407,N_548);
and U751 (N_751,N_482,N_550);
nand U752 (N_752,N_511,N_525);
or U753 (N_753,N_594,N_428);
or U754 (N_754,N_512,N_447);
nor U755 (N_755,N_409,N_475);
and U756 (N_756,N_588,N_553);
nand U757 (N_757,N_452,N_472);
and U758 (N_758,N_598,N_534);
nand U759 (N_759,N_443,N_551);
nor U760 (N_760,N_563,N_575);
xnor U761 (N_761,N_467,N_512);
nor U762 (N_762,N_547,N_490);
or U763 (N_763,N_481,N_401);
or U764 (N_764,N_464,N_489);
xnor U765 (N_765,N_442,N_543);
nand U766 (N_766,N_576,N_566);
or U767 (N_767,N_422,N_491);
xor U768 (N_768,N_468,N_428);
nand U769 (N_769,N_584,N_509);
xnor U770 (N_770,N_482,N_546);
xor U771 (N_771,N_481,N_465);
xnor U772 (N_772,N_490,N_505);
nor U773 (N_773,N_470,N_489);
xor U774 (N_774,N_468,N_524);
and U775 (N_775,N_449,N_536);
and U776 (N_776,N_492,N_566);
xor U777 (N_777,N_462,N_428);
xnor U778 (N_778,N_433,N_508);
xor U779 (N_779,N_519,N_596);
xor U780 (N_780,N_525,N_582);
or U781 (N_781,N_576,N_458);
and U782 (N_782,N_513,N_568);
and U783 (N_783,N_428,N_556);
nor U784 (N_784,N_497,N_440);
and U785 (N_785,N_436,N_544);
xnor U786 (N_786,N_473,N_574);
xnor U787 (N_787,N_442,N_483);
and U788 (N_788,N_498,N_466);
and U789 (N_789,N_504,N_548);
and U790 (N_790,N_567,N_588);
xnor U791 (N_791,N_547,N_418);
or U792 (N_792,N_534,N_405);
nand U793 (N_793,N_428,N_581);
and U794 (N_794,N_487,N_593);
nor U795 (N_795,N_532,N_450);
or U796 (N_796,N_463,N_533);
nor U797 (N_797,N_557,N_426);
nand U798 (N_798,N_419,N_573);
and U799 (N_799,N_510,N_452);
nor U800 (N_800,N_795,N_677);
xnor U801 (N_801,N_610,N_602);
nor U802 (N_802,N_609,N_741);
nand U803 (N_803,N_732,N_652);
nand U804 (N_804,N_751,N_711);
nor U805 (N_805,N_721,N_636);
nand U806 (N_806,N_716,N_611);
nand U807 (N_807,N_743,N_618);
nand U808 (N_808,N_726,N_753);
and U809 (N_809,N_798,N_695);
and U810 (N_810,N_737,N_633);
nand U811 (N_811,N_719,N_730);
and U812 (N_812,N_670,N_604);
or U813 (N_813,N_683,N_634);
nor U814 (N_814,N_693,N_665);
nand U815 (N_815,N_746,N_786);
and U816 (N_816,N_754,N_744);
xnor U817 (N_817,N_606,N_635);
nor U818 (N_818,N_789,N_714);
nand U819 (N_819,N_742,N_675);
and U820 (N_820,N_623,N_615);
nor U821 (N_821,N_662,N_740);
nor U822 (N_822,N_649,N_622);
nor U823 (N_823,N_768,N_766);
nor U824 (N_824,N_724,N_655);
nand U825 (N_825,N_619,N_647);
nand U826 (N_826,N_691,N_725);
or U827 (N_827,N_626,N_729);
nor U828 (N_828,N_661,N_648);
nand U829 (N_829,N_614,N_778);
nand U830 (N_830,N_687,N_660);
xor U831 (N_831,N_631,N_624);
xnor U832 (N_832,N_621,N_710);
and U833 (N_833,N_769,N_776);
xnor U834 (N_834,N_638,N_791);
nor U835 (N_835,N_669,N_722);
nor U836 (N_836,N_756,N_723);
nand U837 (N_837,N_612,N_603);
and U838 (N_838,N_651,N_748);
nor U839 (N_839,N_717,N_685);
nor U840 (N_840,N_787,N_765);
or U841 (N_841,N_601,N_715);
nand U842 (N_842,N_613,N_698);
or U843 (N_843,N_734,N_617);
nor U844 (N_844,N_678,N_681);
nand U845 (N_845,N_701,N_679);
xor U846 (N_846,N_656,N_600);
or U847 (N_847,N_699,N_666);
and U848 (N_848,N_720,N_674);
xor U849 (N_849,N_758,N_797);
nand U850 (N_850,N_779,N_780);
nor U851 (N_851,N_796,N_760);
or U852 (N_852,N_628,N_667);
and U853 (N_853,N_703,N_790);
xor U854 (N_854,N_625,N_735);
and U855 (N_855,N_620,N_728);
nor U856 (N_856,N_727,N_682);
or U857 (N_857,N_692,N_707);
or U858 (N_858,N_738,N_793);
xor U859 (N_859,N_777,N_657);
xnor U860 (N_860,N_772,N_739);
or U861 (N_861,N_627,N_694);
nor U862 (N_862,N_673,N_767);
xor U863 (N_863,N_646,N_771);
nor U864 (N_864,N_745,N_697);
and U865 (N_865,N_676,N_792);
nor U866 (N_866,N_664,N_650);
nor U867 (N_867,N_749,N_770);
and U868 (N_868,N_668,N_700);
nor U869 (N_869,N_689,N_653);
nor U870 (N_870,N_747,N_788);
nand U871 (N_871,N_607,N_764);
or U872 (N_872,N_718,N_690);
nor U873 (N_873,N_709,N_632);
and U874 (N_874,N_684,N_783);
and U875 (N_875,N_736,N_671);
nand U876 (N_876,N_696,N_645);
and U877 (N_877,N_781,N_688);
and U878 (N_878,N_616,N_629);
nor U879 (N_879,N_759,N_773);
and U880 (N_880,N_642,N_643);
or U881 (N_881,N_640,N_755);
nor U882 (N_882,N_672,N_639);
or U883 (N_883,N_608,N_750);
nor U884 (N_884,N_641,N_605);
nand U885 (N_885,N_757,N_712);
nor U886 (N_886,N_731,N_794);
nor U887 (N_887,N_775,N_680);
or U888 (N_888,N_713,N_704);
and U889 (N_889,N_708,N_663);
xor U890 (N_890,N_658,N_705);
and U891 (N_891,N_763,N_637);
or U892 (N_892,N_782,N_774);
nand U893 (N_893,N_654,N_644);
nor U894 (N_894,N_752,N_659);
and U895 (N_895,N_785,N_686);
and U896 (N_896,N_706,N_762);
nand U897 (N_897,N_784,N_799);
and U898 (N_898,N_761,N_733);
or U899 (N_899,N_702,N_630);
nand U900 (N_900,N_717,N_648);
nor U901 (N_901,N_655,N_733);
nor U902 (N_902,N_791,N_654);
xor U903 (N_903,N_691,N_712);
xor U904 (N_904,N_780,N_771);
nor U905 (N_905,N_666,N_602);
or U906 (N_906,N_610,N_628);
or U907 (N_907,N_705,N_634);
xnor U908 (N_908,N_654,N_799);
and U909 (N_909,N_798,N_700);
nor U910 (N_910,N_704,N_752);
and U911 (N_911,N_786,N_674);
xnor U912 (N_912,N_619,N_751);
nand U913 (N_913,N_764,N_751);
xnor U914 (N_914,N_779,N_706);
nand U915 (N_915,N_793,N_605);
or U916 (N_916,N_746,N_735);
nor U917 (N_917,N_776,N_668);
and U918 (N_918,N_773,N_754);
xor U919 (N_919,N_623,N_772);
nand U920 (N_920,N_672,N_601);
xnor U921 (N_921,N_791,N_705);
xor U922 (N_922,N_661,N_782);
nand U923 (N_923,N_688,N_754);
and U924 (N_924,N_603,N_663);
and U925 (N_925,N_640,N_623);
nand U926 (N_926,N_723,N_658);
xor U927 (N_927,N_684,N_678);
nor U928 (N_928,N_718,N_692);
xnor U929 (N_929,N_775,N_785);
and U930 (N_930,N_676,N_785);
and U931 (N_931,N_642,N_616);
and U932 (N_932,N_766,N_739);
and U933 (N_933,N_740,N_795);
nand U934 (N_934,N_721,N_652);
or U935 (N_935,N_608,N_690);
nor U936 (N_936,N_680,N_649);
xor U937 (N_937,N_755,N_708);
nor U938 (N_938,N_785,N_631);
and U939 (N_939,N_728,N_671);
nor U940 (N_940,N_772,N_611);
or U941 (N_941,N_793,N_659);
or U942 (N_942,N_693,N_641);
nand U943 (N_943,N_723,N_771);
nor U944 (N_944,N_662,N_769);
nand U945 (N_945,N_774,N_626);
xor U946 (N_946,N_643,N_621);
xnor U947 (N_947,N_619,N_700);
or U948 (N_948,N_659,N_725);
nor U949 (N_949,N_787,N_760);
nor U950 (N_950,N_633,N_787);
nor U951 (N_951,N_615,N_665);
xnor U952 (N_952,N_721,N_631);
or U953 (N_953,N_722,N_707);
nor U954 (N_954,N_720,N_752);
nor U955 (N_955,N_764,N_714);
and U956 (N_956,N_768,N_775);
or U957 (N_957,N_720,N_730);
and U958 (N_958,N_762,N_774);
and U959 (N_959,N_778,N_788);
nand U960 (N_960,N_684,N_742);
and U961 (N_961,N_721,N_715);
xor U962 (N_962,N_632,N_674);
nor U963 (N_963,N_703,N_644);
nor U964 (N_964,N_679,N_751);
xnor U965 (N_965,N_751,N_602);
and U966 (N_966,N_747,N_638);
xor U967 (N_967,N_696,N_702);
or U968 (N_968,N_695,N_726);
nand U969 (N_969,N_682,N_720);
nor U970 (N_970,N_777,N_678);
xor U971 (N_971,N_761,N_758);
xnor U972 (N_972,N_748,N_757);
nor U973 (N_973,N_720,N_619);
or U974 (N_974,N_644,N_641);
or U975 (N_975,N_628,N_747);
nand U976 (N_976,N_699,N_665);
and U977 (N_977,N_673,N_766);
and U978 (N_978,N_701,N_662);
xor U979 (N_979,N_747,N_605);
nor U980 (N_980,N_783,N_643);
xor U981 (N_981,N_694,N_686);
nand U982 (N_982,N_628,N_622);
nand U983 (N_983,N_655,N_603);
nand U984 (N_984,N_783,N_757);
or U985 (N_985,N_637,N_647);
and U986 (N_986,N_774,N_643);
or U987 (N_987,N_709,N_782);
or U988 (N_988,N_751,N_743);
and U989 (N_989,N_771,N_735);
nand U990 (N_990,N_736,N_624);
nand U991 (N_991,N_745,N_639);
nand U992 (N_992,N_764,N_717);
or U993 (N_993,N_603,N_649);
and U994 (N_994,N_677,N_753);
nand U995 (N_995,N_764,N_710);
and U996 (N_996,N_747,N_708);
nand U997 (N_997,N_644,N_726);
and U998 (N_998,N_779,N_624);
xnor U999 (N_999,N_773,N_624);
or U1000 (N_1000,N_977,N_873);
nand U1001 (N_1001,N_886,N_984);
nand U1002 (N_1002,N_927,N_898);
nand U1003 (N_1003,N_845,N_954);
nor U1004 (N_1004,N_816,N_917);
nand U1005 (N_1005,N_864,N_831);
or U1006 (N_1006,N_961,N_800);
nor U1007 (N_1007,N_807,N_987);
and U1008 (N_1008,N_853,N_993);
nand U1009 (N_1009,N_846,N_970);
or U1010 (N_1010,N_901,N_825);
nand U1011 (N_1011,N_885,N_809);
nor U1012 (N_1012,N_929,N_804);
and U1013 (N_1013,N_948,N_988);
nor U1014 (N_1014,N_887,N_960);
or U1015 (N_1015,N_995,N_969);
and U1016 (N_1016,N_973,N_888);
nor U1017 (N_1017,N_863,N_875);
xnor U1018 (N_1018,N_811,N_882);
and U1019 (N_1019,N_883,N_965);
nor U1020 (N_1020,N_994,N_981);
xnor U1021 (N_1021,N_904,N_830);
nor U1022 (N_1022,N_897,N_802);
xnor U1023 (N_1023,N_972,N_946);
nor U1024 (N_1024,N_998,N_935);
nand U1025 (N_1025,N_860,N_881);
or U1026 (N_1026,N_891,N_909);
nand U1027 (N_1027,N_928,N_952);
xor U1028 (N_1028,N_908,N_944);
xor U1029 (N_1029,N_843,N_953);
nor U1030 (N_1030,N_815,N_949);
nor U1031 (N_1031,N_925,N_962);
nand U1032 (N_1032,N_932,N_833);
and U1033 (N_1033,N_829,N_999);
or U1034 (N_1034,N_836,N_990);
xor U1035 (N_1035,N_936,N_895);
nor U1036 (N_1036,N_819,N_933);
nor U1037 (N_1037,N_905,N_892);
nand U1038 (N_1038,N_834,N_903);
nand U1039 (N_1039,N_850,N_934);
xor U1040 (N_1040,N_823,N_986);
nand U1041 (N_1041,N_907,N_992);
or U1042 (N_1042,N_912,N_982);
nor U1043 (N_1043,N_983,N_841);
xor U1044 (N_1044,N_827,N_810);
xor U1045 (N_1045,N_842,N_820);
and U1046 (N_1046,N_812,N_813);
nor U1047 (N_1047,N_900,N_978);
nor U1048 (N_1048,N_855,N_942);
nand U1049 (N_1049,N_920,N_910);
and U1050 (N_1050,N_902,N_997);
nand U1051 (N_1051,N_808,N_871);
and U1052 (N_1052,N_814,N_849);
nor U1053 (N_1053,N_824,N_865);
or U1054 (N_1054,N_966,N_958);
nor U1055 (N_1055,N_899,N_940);
nand U1056 (N_1056,N_918,N_877);
or U1057 (N_1057,N_818,N_950);
nand U1058 (N_1058,N_919,N_839);
nand U1059 (N_1059,N_822,N_957);
nor U1060 (N_1060,N_857,N_859);
xnor U1061 (N_1061,N_985,N_911);
nand U1062 (N_1062,N_867,N_941);
xnor U1063 (N_1063,N_894,N_832);
xor U1064 (N_1064,N_921,N_854);
nand U1065 (N_1065,N_996,N_989);
or U1066 (N_1066,N_852,N_971);
nor U1067 (N_1067,N_840,N_939);
nor U1068 (N_1068,N_976,N_844);
nand U1069 (N_1069,N_991,N_924);
and U1070 (N_1070,N_805,N_937);
xnor U1071 (N_1071,N_931,N_856);
and U1072 (N_1072,N_801,N_821);
and U1073 (N_1073,N_956,N_930);
nor U1074 (N_1074,N_923,N_893);
and U1075 (N_1075,N_913,N_838);
nand U1076 (N_1076,N_835,N_906);
nor U1077 (N_1077,N_926,N_858);
nand U1078 (N_1078,N_862,N_870);
and U1079 (N_1079,N_980,N_878);
xnor U1080 (N_1080,N_884,N_947);
xor U1081 (N_1081,N_964,N_943);
nand U1082 (N_1082,N_896,N_945);
and U1083 (N_1083,N_872,N_826);
and U1084 (N_1084,N_979,N_861);
nor U1085 (N_1085,N_874,N_847);
xnor U1086 (N_1086,N_868,N_967);
nand U1087 (N_1087,N_974,N_837);
and U1088 (N_1088,N_880,N_968);
xor U1089 (N_1089,N_975,N_959);
and U1090 (N_1090,N_963,N_869);
or U1091 (N_1091,N_915,N_889);
nand U1092 (N_1092,N_922,N_848);
nand U1093 (N_1093,N_803,N_914);
xor U1094 (N_1094,N_938,N_876);
nand U1095 (N_1095,N_866,N_879);
and U1096 (N_1096,N_817,N_955);
xnor U1097 (N_1097,N_916,N_828);
and U1098 (N_1098,N_890,N_851);
or U1099 (N_1099,N_806,N_951);
nand U1100 (N_1100,N_940,N_814);
xnor U1101 (N_1101,N_851,N_840);
or U1102 (N_1102,N_877,N_816);
or U1103 (N_1103,N_954,N_999);
xnor U1104 (N_1104,N_899,N_987);
xor U1105 (N_1105,N_819,N_964);
or U1106 (N_1106,N_880,N_977);
nor U1107 (N_1107,N_849,N_806);
nand U1108 (N_1108,N_860,N_997);
or U1109 (N_1109,N_808,N_963);
nand U1110 (N_1110,N_998,N_934);
or U1111 (N_1111,N_898,N_928);
or U1112 (N_1112,N_939,N_823);
and U1113 (N_1113,N_927,N_890);
nand U1114 (N_1114,N_918,N_916);
nor U1115 (N_1115,N_853,N_871);
nor U1116 (N_1116,N_892,N_882);
or U1117 (N_1117,N_944,N_811);
xnor U1118 (N_1118,N_882,N_995);
nor U1119 (N_1119,N_921,N_960);
and U1120 (N_1120,N_816,N_876);
or U1121 (N_1121,N_855,N_975);
xor U1122 (N_1122,N_892,N_870);
xnor U1123 (N_1123,N_970,N_839);
xnor U1124 (N_1124,N_976,N_928);
xor U1125 (N_1125,N_899,N_903);
nor U1126 (N_1126,N_867,N_923);
and U1127 (N_1127,N_980,N_993);
nand U1128 (N_1128,N_979,N_852);
xor U1129 (N_1129,N_818,N_816);
nand U1130 (N_1130,N_918,N_864);
nand U1131 (N_1131,N_828,N_958);
and U1132 (N_1132,N_928,N_818);
or U1133 (N_1133,N_928,N_951);
or U1134 (N_1134,N_890,N_907);
and U1135 (N_1135,N_963,N_961);
nand U1136 (N_1136,N_922,N_876);
and U1137 (N_1137,N_808,N_893);
nor U1138 (N_1138,N_939,N_819);
xnor U1139 (N_1139,N_832,N_997);
nor U1140 (N_1140,N_831,N_971);
and U1141 (N_1141,N_997,N_866);
and U1142 (N_1142,N_934,N_813);
xnor U1143 (N_1143,N_858,N_907);
and U1144 (N_1144,N_954,N_815);
xnor U1145 (N_1145,N_996,N_999);
or U1146 (N_1146,N_857,N_878);
xor U1147 (N_1147,N_932,N_964);
nor U1148 (N_1148,N_951,N_952);
xor U1149 (N_1149,N_803,N_955);
or U1150 (N_1150,N_957,N_956);
nand U1151 (N_1151,N_867,N_917);
nor U1152 (N_1152,N_812,N_970);
nor U1153 (N_1153,N_903,N_842);
xnor U1154 (N_1154,N_870,N_926);
or U1155 (N_1155,N_834,N_979);
or U1156 (N_1156,N_952,N_892);
and U1157 (N_1157,N_878,N_867);
xor U1158 (N_1158,N_987,N_985);
xnor U1159 (N_1159,N_984,N_814);
nand U1160 (N_1160,N_967,N_987);
xor U1161 (N_1161,N_903,N_851);
xnor U1162 (N_1162,N_932,N_820);
and U1163 (N_1163,N_956,N_991);
nor U1164 (N_1164,N_978,N_973);
nand U1165 (N_1165,N_857,N_905);
nor U1166 (N_1166,N_834,N_960);
and U1167 (N_1167,N_879,N_966);
or U1168 (N_1168,N_909,N_867);
or U1169 (N_1169,N_858,N_923);
xnor U1170 (N_1170,N_819,N_836);
xor U1171 (N_1171,N_862,N_863);
nand U1172 (N_1172,N_883,N_999);
nand U1173 (N_1173,N_912,N_914);
xnor U1174 (N_1174,N_963,N_941);
nor U1175 (N_1175,N_907,N_845);
nor U1176 (N_1176,N_845,N_962);
and U1177 (N_1177,N_903,N_803);
or U1178 (N_1178,N_813,N_976);
nand U1179 (N_1179,N_982,N_863);
nor U1180 (N_1180,N_888,N_914);
xor U1181 (N_1181,N_999,N_988);
nand U1182 (N_1182,N_995,N_996);
nand U1183 (N_1183,N_925,N_978);
and U1184 (N_1184,N_803,N_941);
xnor U1185 (N_1185,N_819,N_968);
nand U1186 (N_1186,N_900,N_986);
xnor U1187 (N_1187,N_857,N_895);
nand U1188 (N_1188,N_825,N_905);
and U1189 (N_1189,N_845,N_980);
and U1190 (N_1190,N_858,N_805);
nand U1191 (N_1191,N_817,N_900);
or U1192 (N_1192,N_886,N_812);
nand U1193 (N_1193,N_945,N_917);
xnor U1194 (N_1194,N_843,N_867);
nor U1195 (N_1195,N_999,N_880);
nand U1196 (N_1196,N_902,N_818);
or U1197 (N_1197,N_931,N_928);
or U1198 (N_1198,N_934,N_990);
and U1199 (N_1199,N_814,N_997);
nand U1200 (N_1200,N_1119,N_1106);
nor U1201 (N_1201,N_1064,N_1118);
and U1202 (N_1202,N_1163,N_1077);
nand U1203 (N_1203,N_1194,N_1051);
nand U1204 (N_1204,N_1083,N_1110);
and U1205 (N_1205,N_1127,N_1100);
nor U1206 (N_1206,N_1013,N_1136);
or U1207 (N_1207,N_1071,N_1022);
or U1208 (N_1208,N_1105,N_1183);
or U1209 (N_1209,N_1143,N_1153);
xor U1210 (N_1210,N_1081,N_1135);
nand U1211 (N_1211,N_1167,N_1180);
nor U1212 (N_1212,N_1054,N_1011);
or U1213 (N_1213,N_1010,N_1045);
or U1214 (N_1214,N_1079,N_1142);
xnor U1215 (N_1215,N_1103,N_1129);
xor U1216 (N_1216,N_1007,N_1168);
and U1217 (N_1217,N_1060,N_1154);
nor U1218 (N_1218,N_1092,N_1063);
or U1219 (N_1219,N_1000,N_1032);
or U1220 (N_1220,N_1021,N_1196);
or U1221 (N_1221,N_1102,N_1169);
nor U1222 (N_1222,N_1175,N_1004);
and U1223 (N_1223,N_1195,N_1041);
or U1224 (N_1224,N_1122,N_1098);
and U1225 (N_1225,N_1025,N_1101);
or U1226 (N_1226,N_1091,N_1146);
nor U1227 (N_1227,N_1087,N_1166);
nand U1228 (N_1228,N_1089,N_1026);
nor U1229 (N_1229,N_1162,N_1096);
nor U1230 (N_1230,N_1125,N_1027);
nand U1231 (N_1231,N_1057,N_1055);
xor U1232 (N_1232,N_1074,N_1171);
nor U1233 (N_1233,N_1151,N_1028);
nand U1234 (N_1234,N_1152,N_1117);
or U1235 (N_1235,N_1065,N_1040);
nand U1236 (N_1236,N_1123,N_1160);
nor U1237 (N_1237,N_1095,N_1053);
and U1238 (N_1238,N_1116,N_1198);
nand U1239 (N_1239,N_1003,N_1138);
xnor U1240 (N_1240,N_1085,N_1048);
nor U1241 (N_1241,N_1121,N_1037);
or U1242 (N_1242,N_1165,N_1097);
or U1243 (N_1243,N_1050,N_1178);
and U1244 (N_1244,N_1069,N_1139);
nand U1245 (N_1245,N_1161,N_1012);
or U1246 (N_1246,N_1197,N_1182);
or U1247 (N_1247,N_1009,N_1086);
nor U1248 (N_1248,N_1158,N_1187);
xor U1249 (N_1249,N_1190,N_1199);
nand U1250 (N_1250,N_1109,N_1020);
xor U1251 (N_1251,N_1059,N_1046);
or U1252 (N_1252,N_1067,N_1072);
nor U1253 (N_1253,N_1113,N_1130);
nand U1254 (N_1254,N_1164,N_1111);
or U1255 (N_1255,N_1185,N_1093);
and U1256 (N_1256,N_1140,N_1192);
nand U1257 (N_1257,N_1155,N_1145);
nand U1258 (N_1258,N_1172,N_1024);
or U1259 (N_1259,N_1137,N_1191);
nor U1260 (N_1260,N_1073,N_1141);
xor U1261 (N_1261,N_1128,N_1133);
xor U1262 (N_1262,N_1006,N_1005);
nand U1263 (N_1263,N_1039,N_1115);
and U1264 (N_1264,N_1108,N_1131);
or U1265 (N_1265,N_1148,N_1104);
nor U1266 (N_1266,N_1094,N_1159);
nand U1267 (N_1267,N_1157,N_1184);
nand U1268 (N_1268,N_1075,N_1035);
or U1269 (N_1269,N_1016,N_1181);
xnor U1270 (N_1270,N_1112,N_1070);
or U1271 (N_1271,N_1107,N_1132);
or U1272 (N_1272,N_1002,N_1008);
nand U1273 (N_1273,N_1170,N_1150);
nand U1274 (N_1274,N_1088,N_1031);
nor U1275 (N_1275,N_1126,N_1082);
nand U1276 (N_1276,N_1090,N_1134);
nor U1277 (N_1277,N_1173,N_1188);
and U1278 (N_1278,N_1018,N_1147);
xor U1279 (N_1279,N_1193,N_1177);
xnor U1280 (N_1280,N_1017,N_1061);
xor U1281 (N_1281,N_1144,N_1034);
nor U1282 (N_1282,N_1014,N_1001);
and U1283 (N_1283,N_1058,N_1099);
nand U1284 (N_1284,N_1114,N_1044);
and U1285 (N_1285,N_1078,N_1149);
and U1286 (N_1286,N_1062,N_1043);
or U1287 (N_1287,N_1030,N_1156);
or U1288 (N_1288,N_1047,N_1080);
nor U1289 (N_1289,N_1189,N_1179);
nor U1290 (N_1290,N_1038,N_1056);
and U1291 (N_1291,N_1029,N_1015);
nor U1292 (N_1292,N_1084,N_1019);
or U1293 (N_1293,N_1068,N_1124);
nand U1294 (N_1294,N_1186,N_1023);
xnor U1295 (N_1295,N_1066,N_1049);
and U1296 (N_1296,N_1036,N_1076);
nand U1297 (N_1297,N_1052,N_1176);
and U1298 (N_1298,N_1042,N_1174);
and U1299 (N_1299,N_1120,N_1033);
or U1300 (N_1300,N_1168,N_1033);
and U1301 (N_1301,N_1197,N_1109);
nor U1302 (N_1302,N_1071,N_1084);
nand U1303 (N_1303,N_1041,N_1089);
and U1304 (N_1304,N_1061,N_1031);
nor U1305 (N_1305,N_1009,N_1105);
nor U1306 (N_1306,N_1117,N_1155);
xor U1307 (N_1307,N_1033,N_1175);
and U1308 (N_1308,N_1135,N_1029);
xor U1309 (N_1309,N_1086,N_1101);
xnor U1310 (N_1310,N_1188,N_1149);
nand U1311 (N_1311,N_1013,N_1018);
nand U1312 (N_1312,N_1089,N_1154);
nand U1313 (N_1313,N_1167,N_1069);
xor U1314 (N_1314,N_1169,N_1010);
nor U1315 (N_1315,N_1105,N_1035);
xnor U1316 (N_1316,N_1000,N_1064);
nor U1317 (N_1317,N_1110,N_1144);
nor U1318 (N_1318,N_1158,N_1169);
nor U1319 (N_1319,N_1129,N_1123);
nand U1320 (N_1320,N_1054,N_1129);
or U1321 (N_1321,N_1116,N_1095);
or U1322 (N_1322,N_1152,N_1171);
nor U1323 (N_1323,N_1129,N_1015);
nor U1324 (N_1324,N_1168,N_1040);
and U1325 (N_1325,N_1095,N_1069);
or U1326 (N_1326,N_1184,N_1140);
nand U1327 (N_1327,N_1087,N_1052);
or U1328 (N_1328,N_1134,N_1089);
or U1329 (N_1329,N_1080,N_1025);
xor U1330 (N_1330,N_1002,N_1005);
xnor U1331 (N_1331,N_1138,N_1015);
xor U1332 (N_1332,N_1195,N_1039);
nor U1333 (N_1333,N_1087,N_1053);
nor U1334 (N_1334,N_1079,N_1110);
nor U1335 (N_1335,N_1104,N_1099);
nand U1336 (N_1336,N_1049,N_1108);
or U1337 (N_1337,N_1199,N_1105);
and U1338 (N_1338,N_1124,N_1063);
nand U1339 (N_1339,N_1029,N_1187);
nor U1340 (N_1340,N_1022,N_1076);
and U1341 (N_1341,N_1028,N_1084);
nor U1342 (N_1342,N_1088,N_1190);
and U1343 (N_1343,N_1086,N_1189);
xnor U1344 (N_1344,N_1044,N_1137);
and U1345 (N_1345,N_1143,N_1014);
and U1346 (N_1346,N_1025,N_1042);
and U1347 (N_1347,N_1193,N_1002);
or U1348 (N_1348,N_1091,N_1073);
xnor U1349 (N_1349,N_1147,N_1032);
nor U1350 (N_1350,N_1197,N_1171);
or U1351 (N_1351,N_1150,N_1020);
or U1352 (N_1352,N_1022,N_1157);
xnor U1353 (N_1353,N_1089,N_1058);
nor U1354 (N_1354,N_1012,N_1085);
or U1355 (N_1355,N_1181,N_1041);
and U1356 (N_1356,N_1120,N_1026);
nand U1357 (N_1357,N_1152,N_1170);
or U1358 (N_1358,N_1147,N_1015);
or U1359 (N_1359,N_1076,N_1120);
and U1360 (N_1360,N_1173,N_1032);
xor U1361 (N_1361,N_1001,N_1154);
nand U1362 (N_1362,N_1120,N_1039);
and U1363 (N_1363,N_1091,N_1057);
and U1364 (N_1364,N_1105,N_1167);
and U1365 (N_1365,N_1020,N_1058);
or U1366 (N_1366,N_1194,N_1185);
nor U1367 (N_1367,N_1007,N_1088);
xor U1368 (N_1368,N_1095,N_1038);
or U1369 (N_1369,N_1197,N_1090);
or U1370 (N_1370,N_1119,N_1148);
nor U1371 (N_1371,N_1043,N_1071);
or U1372 (N_1372,N_1183,N_1076);
or U1373 (N_1373,N_1126,N_1149);
xnor U1374 (N_1374,N_1137,N_1105);
nand U1375 (N_1375,N_1151,N_1052);
nand U1376 (N_1376,N_1161,N_1174);
or U1377 (N_1377,N_1183,N_1155);
and U1378 (N_1378,N_1023,N_1052);
and U1379 (N_1379,N_1099,N_1039);
nand U1380 (N_1380,N_1128,N_1151);
nand U1381 (N_1381,N_1040,N_1058);
nor U1382 (N_1382,N_1058,N_1053);
nand U1383 (N_1383,N_1167,N_1044);
nor U1384 (N_1384,N_1112,N_1109);
nor U1385 (N_1385,N_1037,N_1176);
xnor U1386 (N_1386,N_1005,N_1052);
nand U1387 (N_1387,N_1084,N_1150);
nand U1388 (N_1388,N_1113,N_1023);
nor U1389 (N_1389,N_1092,N_1184);
nand U1390 (N_1390,N_1039,N_1185);
nand U1391 (N_1391,N_1142,N_1013);
xnor U1392 (N_1392,N_1100,N_1163);
and U1393 (N_1393,N_1064,N_1072);
xnor U1394 (N_1394,N_1056,N_1177);
nand U1395 (N_1395,N_1069,N_1126);
or U1396 (N_1396,N_1080,N_1023);
xor U1397 (N_1397,N_1131,N_1144);
or U1398 (N_1398,N_1136,N_1009);
xnor U1399 (N_1399,N_1100,N_1123);
nor U1400 (N_1400,N_1226,N_1275);
nand U1401 (N_1401,N_1363,N_1277);
nor U1402 (N_1402,N_1379,N_1272);
nand U1403 (N_1403,N_1301,N_1358);
or U1404 (N_1404,N_1248,N_1278);
or U1405 (N_1405,N_1320,N_1221);
and U1406 (N_1406,N_1378,N_1218);
xor U1407 (N_1407,N_1213,N_1307);
nand U1408 (N_1408,N_1240,N_1343);
and U1409 (N_1409,N_1375,N_1341);
nand U1410 (N_1410,N_1286,N_1231);
nor U1411 (N_1411,N_1291,N_1207);
nor U1412 (N_1412,N_1298,N_1201);
and U1413 (N_1413,N_1266,N_1276);
nor U1414 (N_1414,N_1251,N_1233);
xor U1415 (N_1415,N_1263,N_1311);
and U1416 (N_1416,N_1377,N_1314);
nor U1417 (N_1417,N_1337,N_1317);
xnor U1418 (N_1418,N_1373,N_1295);
nand U1419 (N_1419,N_1388,N_1284);
nand U1420 (N_1420,N_1269,N_1366);
and U1421 (N_1421,N_1205,N_1394);
and U1422 (N_1422,N_1222,N_1217);
nor U1423 (N_1423,N_1398,N_1354);
and U1424 (N_1424,N_1374,N_1235);
xor U1425 (N_1425,N_1395,N_1345);
nor U1426 (N_1426,N_1316,N_1238);
and U1427 (N_1427,N_1326,N_1229);
and U1428 (N_1428,N_1302,N_1306);
and U1429 (N_1429,N_1247,N_1228);
xnor U1430 (N_1430,N_1250,N_1396);
nor U1431 (N_1431,N_1318,N_1342);
nor U1432 (N_1432,N_1350,N_1313);
and U1433 (N_1433,N_1360,N_1380);
or U1434 (N_1434,N_1293,N_1220);
or U1435 (N_1435,N_1265,N_1353);
or U1436 (N_1436,N_1219,N_1270);
and U1437 (N_1437,N_1339,N_1312);
or U1438 (N_1438,N_1232,N_1385);
xnor U1439 (N_1439,N_1204,N_1390);
nand U1440 (N_1440,N_1223,N_1210);
xor U1441 (N_1441,N_1212,N_1289);
nor U1442 (N_1442,N_1319,N_1281);
and U1443 (N_1443,N_1371,N_1288);
or U1444 (N_1444,N_1334,N_1338);
or U1445 (N_1445,N_1249,N_1308);
nand U1446 (N_1446,N_1389,N_1296);
nand U1447 (N_1447,N_1261,N_1333);
or U1448 (N_1448,N_1356,N_1340);
xor U1449 (N_1449,N_1310,N_1324);
nor U1450 (N_1450,N_1367,N_1268);
and U1451 (N_1451,N_1368,N_1351);
and U1452 (N_1452,N_1297,N_1225);
xnor U1453 (N_1453,N_1362,N_1391);
or U1454 (N_1454,N_1273,N_1393);
and U1455 (N_1455,N_1206,N_1256);
xor U1456 (N_1456,N_1234,N_1230);
and U1457 (N_1457,N_1399,N_1257);
nor U1458 (N_1458,N_1246,N_1372);
xnor U1459 (N_1459,N_1359,N_1322);
nor U1460 (N_1460,N_1203,N_1264);
xnor U1461 (N_1461,N_1357,N_1280);
nand U1462 (N_1462,N_1329,N_1323);
nor U1463 (N_1463,N_1325,N_1202);
and U1464 (N_1464,N_1237,N_1331);
and U1465 (N_1465,N_1255,N_1227);
xnor U1466 (N_1466,N_1344,N_1209);
or U1467 (N_1467,N_1347,N_1245);
nor U1468 (N_1468,N_1303,N_1332);
or U1469 (N_1469,N_1287,N_1387);
or U1470 (N_1470,N_1370,N_1244);
or U1471 (N_1471,N_1242,N_1282);
or U1472 (N_1472,N_1299,N_1241);
nor U1473 (N_1473,N_1267,N_1214);
nor U1474 (N_1474,N_1384,N_1382);
nor U1475 (N_1475,N_1336,N_1211);
or U1476 (N_1476,N_1383,N_1327);
nand U1477 (N_1477,N_1243,N_1305);
nand U1478 (N_1478,N_1200,N_1346);
and U1479 (N_1479,N_1304,N_1239);
xnor U1480 (N_1480,N_1271,N_1274);
nand U1481 (N_1481,N_1321,N_1355);
or U1482 (N_1482,N_1259,N_1292);
nand U1483 (N_1483,N_1283,N_1309);
and U1484 (N_1484,N_1315,N_1352);
nor U1485 (N_1485,N_1285,N_1262);
xor U1486 (N_1486,N_1361,N_1335);
nor U1487 (N_1487,N_1254,N_1330);
nand U1488 (N_1488,N_1224,N_1381);
and U1489 (N_1489,N_1369,N_1215);
and U1490 (N_1490,N_1392,N_1300);
or U1491 (N_1491,N_1376,N_1290);
and U1492 (N_1492,N_1328,N_1365);
nor U1493 (N_1493,N_1279,N_1216);
or U1494 (N_1494,N_1349,N_1252);
and U1495 (N_1495,N_1364,N_1260);
nor U1496 (N_1496,N_1386,N_1397);
nand U1497 (N_1497,N_1258,N_1236);
nand U1498 (N_1498,N_1294,N_1208);
nand U1499 (N_1499,N_1253,N_1348);
nor U1500 (N_1500,N_1358,N_1389);
nor U1501 (N_1501,N_1257,N_1203);
or U1502 (N_1502,N_1259,N_1208);
or U1503 (N_1503,N_1399,N_1365);
nand U1504 (N_1504,N_1313,N_1332);
and U1505 (N_1505,N_1244,N_1345);
or U1506 (N_1506,N_1223,N_1292);
nand U1507 (N_1507,N_1261,N_1344);
nor U1508 (N_1508,N_1234,N_1339);
xor U1509 (N_1509,N_1239,N_1312);
xnor U1510 (N_1510,N_1296,N_1318);
or U1511 (N_1511,N_1339,N_1265);
nor U1512 (N_1512,N_1302,N_1394);
nand U1513 (N_1513,N_1203,N_1385);
and U1514 (N_1514,N_1301,N_1225);
nor U1515 (N_1515,N_1270,N_1203);
nand U1516 (N_1516,N_1267,N_1306);
nand U1517 (N_1517,N_1253,N_1222);
xor U1518 (N_1518,N_1224,N_1266);
or U1519 (N_1519,N_1274,N_1367);
or U1520 (N_1520,N_1257,N_1303);
or U1521 (N_1521,N_1217,N_1372);
xor U1522 (N_1522,N_1294,N_1308);
nand U1523 (N_1523,N_1211,N_1370);
xnor U1524 (N_1524,N_1217,N_1338);
nand U1525 (N_1525,N_1294,N_1280);
nor U1526 (N_1526,N_1395,N_1231);
nor U1527 (N_1527,N_1317,N_1384);
xor U1528 (N_1528,N_1330,N_1342);
nand U1529 (N_1529,N_1237,N_1290);
nand U1530 (N_1530,N_1236,N_1308);
nand U1531 (N_1531,N_1222,N_1307);
or U1532 (N_1532,N_1336,N_1398);
and U1533 (N_1533,N_1221,N_1324);
or U1534 (N_1534,N_1397,N_1338);
xor U1535 (N_1535,N_1388,N_1245);
nand U1536 (N_1536,N_1218,N_1331);
xor U1537 (N_1537,N_1377,N_1208);
and U1538 (N_1538,N_1295,N_1267);
and U1539 (N_1539,N_1233,N_1245);
nand U1540 (N_1540,N_1220,N_1247);
nand U1541 (N_1541,N_1208,N_1311);
xnor U1542 (N_1542,N_1251,N_1337);
nand U1543 (N_1543,N_1214,N_1280);
and U1544 (N_1544,N_1317,N_1304);
or U1545 (N_1545,N_1206,N_1323);
nand U1546 (N_1546,N_1299,N_1368);
xnor U1547 (N_1547,N_1200,N_1227);
nor U1548 (N_1548,N_1247,N_1283);
or U1549 (N_1549,N_1383,N_1347);
nor U1550 (N_1550,N_1391,N_1280);
and U1551 (N_1551,N_1288,N_1205);
and U1552 (N_1552,N_1379,N_1307);
xnor U1553 (N_1553,N_1203,N_1302);
or U1554 (N_1554,N_1383,N_1372);
or U1555 (N_1555,N_1351,N_1324);
nand U1556 (N_1556,N_1276,N_1374);
nand U1557 (N_1557,N_1236,N_1263);
nand U1558 (N_1558,N_1258,N_1301);
and U1559 (N_1559,N_1391,N_1296);
nand U1560 (N_1560,N_1208,N_1382);
nand U1561 (N_1561,N_1230,N_1344);
or U1562 (N_1562,N_1219,N_1208);
or U1563 (N_1563,N_1365,N_1340);
xnor U1564 (N_1564,N_1360,N_1234);
xnor U1565 (N_1565,N_1353,N_1235);
xnor U1566 (N_1566,N_1256,N_1297);
nor U1567 (N_1567,N_1318,N_1242);
or U1568 (N_1568,N_1234,N_1231);
nor U1569 (N_1569,N_1345,N_1311);
xnor U1570 (N_1570,N_1389,N_1300);
and U1571 (N_1571,N_1274,N_1380);
or U1572 (N_1572,N_1323,N_1259);
or U1573 (N_1573,N_1372,N_1263);
nor U1574 (N_1574,N_1360,N_1351);
nand U1575 (N_1575,N_1236,N_1287);
or U1576 (N_1576,N_1317,N_1324);
nor U1577 (N_1577,N_1346,N_1316);
nand U1578 (N_1578,N_1285,N_1255);
and U1579 (N_1579,N_1322,N_1213);
or U1580 (N_1580,N_1218,N_1321);
nor U1581 (N_1581,N_1368,N_1241);
nand U1582 (N_1582,N_1285,N_1288);
nor U1583 (N_1583,N_1345,N_1300);
nor U1584 (N_1584,N_1285,N_1221);
nand U1585 (N_1585,N_1309,N_1336);
and U1586 (N_1586,N_1396,N_1230);
xnor U1587 (N_1587,N_1270,N_1267);
and U1588 (N_1588,N_1271,N_1373);
nor U1589 (N_1589,N_1232,N_1307);
and U1590 (N_1590,N_1270,N_1385);
nand U1591 (N_1591,N_1315,N_1368);
xnor U1592 (N_1592,N_1258,N_1317);
nor U1593 (N_1593,N_1243,N_1202);
or U1594 (N_1594,N_1288,N_1298);
and U1595 (N_1595,N_1274,N_1226);
xor U1596 (N_1596,N_1322,N_1367);
nand U1597 (N_1597,N_1341,N_1323);
nand U1598 (N_1598,N_1267,N_1253);
and U1599 (N_1599,N_1369,N_1332);
xor U1600 (N_1600,N_1516,N_1484);
nor U1601 (N_1601,N_1434,N_1496);
nor U1602 (N_1602,N_1460,N_1512);
or U1603 (N_1603,N_1574,N_1557);
nor U1604 (N_1604,N_1528,N_1442);
nor U1605 (N_1605,N_1451,N_1564);
xnor U1606 (N_1606,N_1549,N_1504);
xnor U1607 (N_1607,N_1492,N_1401);
nand U1608 (N_1608,N_1466,N_1413);
and U1609 (N_1609,N_1481,N_1506);
or U1610 (N_1610,N_1456,N_1432);
or U1611 (N_1611,N_1548,N_1527);
xor U1612 (N_1612,N_1446,N_1493);
nor U1613 (N_1613,N_1416,N_1536);
or U1614 (N_1614,N_1577,N_1480);
nand U1615 (N_1615,N_1579,N_1561);
nor U1616 (N_1616,N_1449,N_1403);
nor U1617 (N_1617,N_1558,N_1468);
nand U1618 (N_1618,N_1458,N_1587);
nor U1619 (N_1619,N_1569,N_1479);
nand U1620 (N_1620,N_1529,N_1483);
xnor U1621 (N_1621,N_1542,N_1552);
nor U1622 (N_1622,N_1475,N_1571);
xor U1623 (N_1623,N_1547,N_1515);
nand U1624 (N_1624,N_1538,N_1514);
nor U1625 (N_1625,N_1582,N_1505);
nor U1626 (N_1626,N_1533,N_1445);
xnor U1627 (N_1627,N_1502,N_1570);
xor U1628 (N_1628,N_1486,N_1510);
and U1629 (N_1629,N_1448,N_1584);
nand U1630 (N_1630,N_1411,N_1423);
or U1631 (N_1631,N_1556,N_1498);
or U1632 (N_1632,N_1581,N_1525);
nand U1633 (N_1633,N_1541,N_1566);
nor U1634 (N_1634,N_1440,N_1537);
and U1635 (N_1635,N_1490,N_1465);
and U1636 (N_1636,N_1439,N_1469);
nand U1637 (N_1637,N_1511,N_1425);
or U1638 (N_1638,N_1550,N_1489);
or U1639 (N_1639,N_1414,N_1450);
nor U1640 (N_1640,N_1530,N_1578);
xnor U1641 (N_1641,N_1501,N_1443);
nand U1642 (N_1642,N_1599,N_1539);
nor U1643 (N_1643,N_1453,N_1554);
nand U1644 (N_1644,N_1437,N_1565);
xor U1645 (N_1645,N_1412,N_1592);
nor U1646 (N_1646,N_1419,N_1474);
and U1647 (N_1647,N_1509,N_1424);
or U1648 (N_1648,N_1422,N_1477);
and U1649 (N_1649,N_1568,N_1467);
nor U1650 (N_1650,N_1596,N_1438);
nand U1651 (N_1651,N_1589,N_1531);
nand U1652 (N_1652,N_1462,N_1583);
or U1653 (N_1653,N_1518,N_1408);
nor U1654 (N_1654,N_1526,N_1573);
xnor U1655 (N_1655,N_1567,N_1420);
and U1656 (N_1656,N_1441,N_1435);
nor U1657 (N_1657,N_1591,N_1560);
nor U1658 (N_1658,N_1455,N_1430);
xor U1659 (N_1659,N_1508,N_1482);
or U1660 (N_1660,N_1551,N_1524);
or U1661 (N_1661,N_1595,N_1521);
and U1662 (N_1662,N_1494,N_1457);
and U1663 (N_1663,N_1546,N_1523);
xor U1664 (N_1664,N_1472,N_1459);
xnor U1665 (N_1665,N_1487,N_1405);
and U1666 (N_1666,N_1471,N_1562);
and U1667 (N_1667,N_1410,N_1559);
or U1668 (N_1668,N_1540,N_1491);
or U1669 (N_1669,N_1452,N_1431);
xor U1670 (N_1670,N_1500,N_1580);
nor U1671 (N_1671,N_1594,N_1586);
or U1672 (N_1672,N_1593,N_1545);
nand U1673 (N_1673,N_1454,N_1427);
or U1674 (N_1674,N_1436,N_1478);
xnor U1675 (N_1675,N_1585,N_1418);
nand U1676 (N_1676,N_1495,N_1473);
nand U1677 (N_1677,N_1499,N_1544);
and U1678 (N_1678,N_1555,N_1409);
xnor U1679 (N_1679,N_1461,N_1428);
and U1680 (N_1680,N_1517,N_1543);
xor U1681 (N_1681,N_1470,N_1415);
nor U1682 (N_1682,N_1404,N_1522);
and U1683 (N_1683,N_1519,N_1464);
nand U1684 (N_1684,N_1426,N_1576);
and U1685 (N_1685,N_1507,N_1598);
nor U1686 (N_1686,N_1476,N_1433);
nand U1687 (N_1687,N_1488,N_1535);
nand U1688 (N_1688,N_1429,N_1417);
nand U1689 (N_1689,N_1513,N_1497);
or U1690 (N_1690,N_1520,N_1588);
and U1691 (N_1691,N_1534,N_1575);
and U1692 (N_1692,N_1597,N_1421);
nor U1693 (N_1693,N_1563,N_1444);
xnor U1694 (N_1694,N_1406,N_1400);
and U1695 (N_1695,N_1553,N_1503);
xor U1696 (N_1696,N_1485,N_1463);
nor U1697 (N_1697,N_1572,N_1532);
nand U1698 (N_1698,N_1402,N_1407);
and U1699 (N_1699,N_1447,N_1590);
xnor U1700 (N_1700,N_1465,N_1525);
xnor U1701 (N_1701,N_1469,N_1585);
and U1702 (N_1702,N_1410,N_1472);
or U1703 (N_1703,N_1445,N_1522);
and U1704 (N_1704,N_1591,N_1513);
or U1705 (N_1705,N_1524,N_1480);
xnor U1706 (N_1706,N_1509,N_1531);
xor U1707 (N_1707,N_1459,N_1575);
and U1708 (N_1708,N_1563,N_1513);
nand U1709 (N_1709,N_1496,N_1493);
nor U1710 (N_1710,N_1459,N_1425);
nand U1711 (N_1711,N_1440,N_1486);
and U1712 (N_1712,N_1504,N_1401);
nor U1713 (N_1713,N_1444,N_1528);
xor U1714 (N_1714,N_1559,N_1571);
xnor U1715 (N_1715,N_1437,N_1449);
nand U1716 (N_1716,N_1581,N_1558);
nor U1717 (N_1717,N_1512,N_1406);
xor U1718 (N_1718,N_1588,N_1417);
and U1719 (N_1719,N_1478,N_1530);
or U1720 (N_1720,N_1421,N_1446);
or U1721 (N_1721,N_1514,N_1549);
or U1722 (N_1722,N_1534,N_1404);
or U1723 (N_1723,N_1486,N_1462);
nand U1724 (N_1724,N_1541,N_1438);
xnor U1725 (N_1725,N_1407,N_1453);
nor U1726 (N_1726,N_1569,N_1521);
nand U1727 (N_1727,N_1479,N_1599);
nor U1728 (N_1728,N_1427,N_1417);
or U1729 (N_1729,N_1521,N_1469);
nor U1730 (N_1730,N_1576,N_1503);
and U1731 (N_1731,N_1545,N_1464);
nand U1732 (N_1732,N_1516,N_1477);
or U1733 (N_1733,N_1487,N_1441);
nor U1734 (N_1734,N_1461,N_1598);
or U1735 (N_1735,N_1477,N_1585);
or U1736 (N_1736,N_1464,N_1475);
or U1737 (N_1737,N_1525,N_1455);
xnor U1738 (N_1738,N_1581,N_1403);
or U1739 (N_1739,N_1554,N_1425);
xnor U1740 (N_1740,N_1549,N_1529);
nor U1741 (N_1741,N_1490,N_1406);
nor U1742 (N_1742,N_1543,N_1513);
nor U1743 (N_1743,N_1530,N_1466);
xnor U1744 (N_1744,N_1515,N_1573);
and U1745 (N_1745,N_1481,N_1554);
nor U1746 (N_1746,N_1521,N_1478);
and U1747 (N_1747,N_1421,N_1585);
nor U1748 (N_1748,N_1582,N_1470);
xnor U1749 (N_1749,N_1493,N_1480);
or U1750 (N_1750,N_1524,N_1442);
xnor U1751 (N_1751,N_1476,N_1487);
or U1752 (N_1752,N_1483,N_1583);
and U1753 (N_1753,N_1531,N_1586);
and U1754 (N_1754,N_1452,N_1545);
nand U1755 (N_1755,N_1584,N_1563);
nor U1756 (N_1756,N_1409,N_1432);
or U1757 (N_1757,N_1554,N_1492);
and U1758 (N_1758,N_1475,N_1518);
or U1759 (N_1759,N_1438,N_1441);
xor U1760 (N_1760,N_1477,N_1471);
xor U1761 (N_1761,N_1527,N_1433);
xor U1762 (N_1762,N_1495,N_1599);
xor U1763 (N_1763,N_1470,N_1432);
nand U1764 (N_1764,N_1560,N_1441);
or U1765 (N_1765,N_1434,N_1545);
or U1766 (N_1766,N_1413,N_1537);
or U1767 (N_1767,N_1441,N_1483);
or U1768 (N_1768,N_1481,N_1493);
nand U1769 (N_1769,N_1499,N_1550);
and U1770 (N_1770,N_1442,N_1435);
and U1771 (N_1771,N_1427,N_1477);
xnor U1772 (N_1772,N_1410,N_1441);
or U1773 (N_1773,N_1445,N_1596);
nand U1774 (N_1774,N_1583,N_1498);
xnor U1775 (N_1775,N_1463,N_1589);
nor U1776 (N_1776,N_1566,N_1456);
nand U1777 (N_1777,N_1479,N_1503);
xnor U1778 (N_1778,N_1465,N_1454);
and U1779 (N_1779,N_1543,N_1404);
xor U1780 (N_1780,N_1545,N_1525);
and U1781 (N_1781,N_1526,N_1510);
or U1782 (N_1782,N_1505,N_1434);
or U1783 (N_1783,N_1542,N_1432);
nor U1784 (N_1784,N_1581,N_1401);
nor U1785 (N_1785,N_1484,N_1536);
nand U1786 (N_1786,N_1560,N_1563);
or U1787 (N_1787,N_1548,N_1572);
or U1788 (N_1788,N_1572,N_1593);
and U1789 (N_1789,N_1492,N_1487);
and U1790 (N_1790,N_1572,N_1595);
xnor U1791 (N_1791,N_1423,N_1421);
nor U1792 (N_1792,N_1589,N_1562);
nand U1793 (N_1793,N_1413,N_1548);
nor U1794 (N_1794,N_1536,N_1473);
xnor U1795 (N_1795,N_1460,N_1469);
and U1796 (N_1796,N_1590,N_1464);
nand U1797 (N_1797,N_1430,N_1440);
nand U1798 (N_1798,N_1511,N_1577);
and U1799 (N_1799,N_1506,N_1474);
nand U1800 (N_1800,N_1776,N_1770);
nor U1801 (N_1801,N_1661,N_1663);
nand U1802 (N_1802,N_1711,N_1612);
nor U1803 (N_1803,N_1790,N_1649);
nor U1804 (N_1804,N_1670,N_1730);
nand U1805 (N_1805,N_1746,N_1753);
or U1806 (N_1806,N_1761,N_1689);
nand U1807 (N_1807,N_1749,N_1762);
or U1808 (N_1808,N_1660,N_1675);
or U1809 (N_1809,N_1739,N_1691);
nand U1810 (N_1810,N_1760,N_1683);
xor U1811 (N_1811,N_1719,N_1605);
xor U1812 (N_1812,N_1635,N_1604);
nor U1813 (N_1813,N_1791,N_1772);
nand U1814 (N_1814,N_1621,N_1716);
and U1815 (N_1815,N_1743,N_1608);
and U1816 (N_1816,N_1742,N_1644);
and U1817 (N_1817,N_1633,N_1688);
or U1818 (N_1818,N_1609,N_1655);
and U1819 (N_1819,N_1636,N_1671);
xor U1820 (N_1820,N_1767,N_1678);
xor U1821 (N_1821,N_1773,N_1750);
nand U1822 (N_1822,N_1640,N_1641);
xor U1823 (N_1823,N_1706,N_1685);
and U1824 (N_1824,N_1657,N_1718);
or U1825 (N_1825,N_1673,N_1617);
and U1826 (N_1826,N_1793,N_1710);
or U1827 (N_1827,N_1796,N_1619);
nand U1828 (N_1828,N_1687,N_1727);
nor U1829 (N_1829,N_1734,N_1722);
nand U1830 (N_1830,N_1634,N_1638);
and U1831 (N_1831,N_1769,N_1603);
xnor U1832 (N_1832,N_1611,N_1795);
and U1833 (N_1833,N_1786,N_1668);
nor U1834 (N_1834,N_1610,N_1792);
nor U1835 (N_1835,N_1723,N_1709);
nor U1836 (N_1836,N_1616,N_1606);
nor U1837 (N_1837,N_1696,N_1724);
nor U1838 (N_1838,N_1680,N_1684);
nor U1839 (N_1839,N_1715,N_1628);
xnor U1840 (N_1840,N_1703,N_1741);
and U1841 (N_1841,N_1783,N_1720);
xnor U1842 (N_1842,N_1614,N_1707);
or U1843 (N_1843,N_1717,N_1702);
nand U1844 (N_1844,N_1699,N_1654);
nand U1845 (N_1845,N_1721,N_1764);
and U1846 (N_1846,N_1713,N_1697);
or U1847 (N_1847,N_1650,N_1704);
nor U1848 (N_1848,N_1625,N_1771);
nor U1849 (N_1849,N_1627,N_1690);
or U1850 (N_1850,N_1622,N_1639);
nand U1851 (N_1851,N_1701,N_1692);
or U1852 (N_1852,N_1726,N_1672);
xor U1853 (N_1853,N_1600,N_1787);
nor U1854 (N_1854,N_1781,N_1737);
nand U1855 (N_1855,N_1789,N_1666);
and U1856 (N_1856,N_1631,N_1662);
nand U1857 (N_1857,N_1758,N_1658);
or U1858 (N_1858,N_1731,N_1765);
xor U1859 (N_1859,N_1629,N_1775);
nand U1860 (N_1860,N_1752,N_1725);
and U1861 (N_1861,N_1756,N_1676);
and U1862 (N_1862,N_1618,N_1733);
nor U1863 (N_1863,N_1630,N_1607);
nor U1864 (N_1864,N_1754,N_1766);
xor U1865 (N_1865,N_1682,N_1708);
and U1866 (N_1866,N_1736,N_1744);
nor U1867 (N_1867,N_1788,N_1653);
nor U1868 (N_1868,N_1798,N_1664);
and U1869 (N_1869,N_1679,N_1651);
nand U1870 (N_1870,N_1785,N_1674);
nor U1871 (N_1871,N_1615,N_1768);
and U1872 (N_1872,N_1700,N_1613);
nor U1873 (N_1873,N_1686,N_1782);
nand U1874 (N_1874,N_1777,N_1714);
or U1875 (N_1875,N_1645,N_1735);
nor U1876 (N_1876,N_1643,N_1681);
or U1877 (N_1877,N_1748,N_1747);
nand U1878 (N_1878,N_1646,N_1751);
or U1879 (N_1879,N_1652,N_1694);
nand U1880 (N_1880,N_1778,N_1779);
and U1881 (N_1881,N_1659,N_1669);
or U1882 (N_1882,N_1759,N_1677);
or U1883 (N_1883,N_1784,N_1712);
nand U1884 (N_1884,N_1738,N_1647);
xnor U1885 (N_1885,N_1667,N_1693);
xor U1886 (N_1886,N_1705,N_1602);
or U1887 (N_1887,N_1732,N_1797);
or U1888 (N_1888,N_1656,N_1728);
nand U1889 (N_1889,N_1794,N_1624);
and U1890 (N_1890,N_1698,N_1601);
and U1891 (N_1891,N_1623,N_1799);
xnor U1892 (N_1892,N_1755,N_1757);
nor U1893 (N_1893,N_1695,N_1763);
and U1894 (N_1894,N_1642,N_1620);
or U1895 (N_1895,N_1774,N_1745);
nor U1896 (N_1896,N_1740,N_1780);
and U1897 (N_1897,N_1626,N_1665);
or U1898 (N_1898,N_1648,N_1637);
xor U1899 (N_1899,N_1632,N_1729);
or U1900 (N_1900,N_1609,N_1713);
nor U1901 (N_1901,N_1679,N_1706);
and U1902 (N_1902,N_1731,N_1622);
nor U1903 (N_1903,N_1610,N_1716);
xnor U1904 (N_1904,N_1736,N_1607);
nand U1905 (N_1905,N_1609,N_1641);
nand U1906 (N_1906,N_1737,N_1662);
xor U1907 (N_1907,N_1618,N_1775);
xnor U1908 (N_1908,N_1626,N_1721);
xnor U1909 (N_1909,N_1707,N_1749);
nor U1910 (N_1910,N_1622,N_1711);
nor U1911 (N_1911,N_1718,N_1717);
xor U1912 (N_1912,N_1791,N_1652);
and U1913 (N_1913,N_1787,N_1707);
nor U1914 (N_1914,N_1776,N_1698);
xnor U1915 (N_1915,N_1765,N_1708);
xnor U1916 (N_1916,N_1700,N_1687);
or U1917 (N_1917,N_1699,N_1650);
or U1918 (N_1918,N_1614,N_1600);
xor U1919 (N_1919,N_1653,N_1792);
and U1920 (N_1920,N_1623,N_1697);
xor U1921 (N_1921,N_1667,N_1674);
nor U1922 (N_1922,N_1698,N_1699);
nand U1923 (N_1923,N_1799,N_1703);
nand U1924 (N_1924,N_1732,N_1603);
or U1925 (N_1925,N_1669,N_1782);
nor U1926 (N_1926,N_1620,N_1772);
nor U1927 (N_1927,N_1650,N_1685);
and U1928 (N_1928,N_1622,N_1656);
nor U1929 (N_1929,N_1602,N_1759);
or U1930 (N_1930,N_1719,N_1797);
nor U1931 (N_1931,N_1761,N_1637);
nand U1932 (N_1932,N_1733,N_1749);
nand U1933 (N_1933,N_1730,N_1777);
nor U1934 (N_1934,N_1734,N_1615);
xor U1935 (N_1935,N_1741,N_1617);
and U1936 (N_1936,N_1718,N_1619);
xnor U1937 (N_1937,N_1719,N_1777);
or U1938 (N_1938,N_1739,N_1742);
nand U1939 (N_1939,N_1641,N_1654);
or U1940 (N_1940,N_1727,N_1747);
and U1941 (N_1941,N_1747,N_1774);
and U1942 (N_1942,N_1767,N_1611);
xnor U1943 (N_1943,N_1794,N_1789);
nand U1944 (N_1944,N_1781,N_1768);
or U1945 (N_1945,N_1715,N_1601);
or U1946 (N_1946,N_1782,N_1663);
and U1947 (N_1947,N_1718,N_1620);
nand U1948 (N_1948,N_1754,N_1778);
or U1949 (N_1949,N_1615,N_1738);
xnor U1950 (N_1950,N_1738,N_1644);
xnor U1951 (N_1951,N_1646,N_1658);
nor U1952 (N_1952,N_1779,N_1629);
xor U1953 (N_1953,N_1761,N_1714);
or U1954 (N_1954,N_1751,N_1726);
and U1955 (N_1955,N_1750,N_1740);
or U1956 (N_1956,N_1621,N_1763);
and U1957 (N_1957,N_1731,N_1715);
nand U1958 (N_1958,N_1695,N_1737);
xor U1959 (N_1959,N_1675,N_1656);
or U1960 (N_1960,N_1726,N_1783);
nand U1961 (N_1961,N_1705,N_1797);
or U1962 (N_1962,N_1699,N_1756);
nor U1963 (N_1963,N_1787,N_1711);
nand U1964 (N_1964,N_1652,N_1637);
xor U1965 (N_1965,N_1698,N_1608);
and U1966 (N_1966,N_1612,N_1703);
or U1967 (N_1967,N_1670,N_1739);
and U1968 (N_1968,N_1641,N_1759);
xnor U1969 (N_1969,N_1676,N_1790);
or U1970 (N_1970,N_1695,N_1663);
and U1971 (N_1971,N_1779,N_1683);
and U1972 (N_1972,N_1727,N_1792);
and U1973 (N_1973,N_1742,N_1743);
nor U1974 (N_1974,N_1617,N_1640);
nand U1975 (N_1975,N_1645,N_1744);
or U1976 (N_1976,N_1692,N_1628);
xnor U1977 (N_1977,N_1650,N_1661);
nor U1978 (N_1978,N_1782,N_1717);
or U1979 (N_1979,N_1732,N_1738);
or U1980 (N_1980,N_1613,N_1618);
nor U1981 (N_1981,N_1725,N_1759);
or U1982 (N_1982,N_1717,N_1642);
and U1983 (N_1983,N_1716,N_1623);
and U1984 (N_1984,N_1705,N_1634);
or U1985 (N_1985,N_1747,N_1640);
and U1986 (N_1986,N_1748,N_1616);
or U1987 (N_1987,N_1707,N_1751);
nand U1988 (N_1988,N_1797,N_1758);
xor U1989 (N_1989,N_1775,N_1734);
xor U1990 (N_1990,N_1689,N_1713);
nand U1991 (N_1991,N_1683,N_1730);
xnor U1992 (N_1992,N_1603,N_1604);
and U1993 (N_1993,N_1761,N_1795);
xnor U1994 (N_1994,N_1600,N_1635);
nor U1995 (N_1995,N_1612,N_1768);
xor U1996 (N_1996,N_1718,N_1644);
xor U1997 (N_1997,N_1713,N_1647);
or U1998 (N_1998,N_1751,N_1669);
and U1999 (N_1999,N_1702,N_1658);
or U2000 (N_2000,N_1969,N_1923);
and U2001 (N_2001,N_1983,N_1884);
nand U2002 (N_2002,N_1811,N_1854);
xor U2003 (N_2003,N_1926,N_1894);
xnor U2004 (N_2004,N_1818,N_1945);
nand U2005 (N_2005,N_1816,N_1905);
xnor U2006 (N_2006,N_1862,N_1840);
and U2007 (N_2007,N_1901,N_1868);
nand U2008 (N_2008,N_1910,N_1833);
or U2009 (N_2009,N_1971,N_1907);
nor U2010 (N_2010,N_1891,N_1902);
nor U2011 (N_2011,N_1878,N_1917);
or U2012 (N_2012,N_1898,N_1890);
and U2013 (N_2013,N_1807,N_1974);
and U2014 (N_2014,N_1880,N_1994);
nand U2015 (N_2015,N_1920,N_1822);
and U2016 (N_2016,N_1951,N_1936);
nor U2017 (N_2017,N_1808,N_1848);
nand U2018 (N_2018,N_1801,N_1900);
and U2019 (N_2019,N_1837,N_1961);
and U2020 (N_2020,N_1999,N_1869);
nand U2021 (N_2021,N_1815,N_1872);
nor U2022 (N_2022,N_1873,N_1934);
and U2023 (N_2023,N_1942,N_1863);
and U2024 (N_2024,N_1913,N_1829);
nor U2025 (N_2025,N_1877,N_1897);
nand U2026 (N_2026,N_1982,N_1813);
nor U2027 (N_2027,N_1879,N_1827);
and U2028 (N_2028,N_1941,N_1979);
xnor U2029 (N_2029,N_1928,N_1978);
and U2030 (N_2030,N_1859,N_1949);
or U2031 (N_2031,N_1881,N_1975);
nor U2032 (N_2032,N_1903,N_1857);
nand U2033 (N_2033,N_1933,N_1866);
or U2034 (N_2034,N_1855,N_1943);
and U2035 (N_2035,N_1956,N_1885);
nor U2036 (N_2036,N_1906,N_1952);
xor U2037 (N_2037,N_1981,N_1925);
nor U2038 (N_2038,N_1939,N_1856);
xor U2039 (N_2039,N_1957,N_1966);
or U2040 (N_2040,N_1865,N_1842);
xor U2041 (N_2041,N_1944,N_1990);
or U2042 (N_2042,N_1893,N_1882);
or U2043 (N_2043,N_1812,N_1922);
nor U2044 (N_2044,N_1962,N_1932);
nand U2045 (N_2045,N_1916,N_1846);
nand U2046 (N_2046,N_1993,N_1914);
nand U2047 (N_2047,N_1940,N_1947);
xor U2048 (N_2048,N_1921,N_1870);
and U2049 (N_2049,N_1953,N_1985);
nor U2050 (N_2050,N_1844,N_1858);
or U2051 (N_2051,N_1876,N_1988);
or U2052 (N_2052,N_1805,N_1828);
or U2053 (N_2053,N_1826,N_1960);
nand U2054 (N_2054,N_1834,N_1852);
and U2055 (N_2055,N_1888,N_1970);
xnor U2056 (N_2056,N_1883,N_1929);
nand U2057 (N_2057,N_1806,N_1927);
nor U2058 (N_2058,N_1867,N_1959);
nor U2059 (N_2059,N_1976,N_1937);
nor U2060 (N_2060,N_1850,N_1972);
nor U2061 (N_2061,N_1935,N_1909);
xor U2062 (N_2062,N_1845,N_1924);
or U2063 (N_2063,N_1820,N_1823);
xnor U2064 (N_2064,N_1958,N_1892);
nand U2065 (N_2065,N_1802,N_1887);
and U2066 (N_2066,N_1817,N_1835);
or U2067 (N_2067,N_1896,N_1995);
and U2068 (N_2068,N_1998,N_1821);
nand U2069 (N_2069,N_1973,N_1819);
and U2070 (N_2070,N_1946,N_1874);
nor U2071 (N_2071,N_1830,N_1851);
nand U2072 (N_2072,N_1860,N_1997);
or U2073 (N_2073,N_1809,N_1930);
nand U2074 (N_2074,N_1841,N_1987);
or U2075 (N_2075,N_1899,N_1871);
nor U2076 (N_2076,N_1967,N_1992);
nand U2077 (N_2077,N_1918,N_1875);
nor U2078 (N_2078,N_1886,N_1810);
and U2079 (N_2079,N_1991,N_1853);
xnor U2080 (N_2080,N_1904,N_1996);
nor U2081 (N_2081,N_1838,N_1912);
nor U2082 (N_2082,N_1843,N_1955);
or U2083 (N_2083,N_1963,N_1977);
xor U2084 (N_2084,N_1984,N_1965);
xnor U2085 (N_2085,N_1911,N_1832);
xor U2086 (N_2086,N_1804,N_1847);
or U2087 (N_2087,N_1831,N_1964);
nand U2088 (N_2088,N_1986,N_1948);
and U2089 (N_2089,N_1864,N_1989);
xnor U2090 (N_2090,N_1895,N_1861);
nand U2091 (N_2091,N_1814,N_1980);
and U2092 (N_2092,N_1889,N_1938);
nand U2093 (N_2093,N_1915,N_1954);
or U2094 (N_2094,N_1803,N_1836);
or U2095 (N_2095,N_1825,N_1908);
and U2096 (N_2096,N_1950,N_1968);
or U2097 (N_2097,N_1800,N_1919);
xnor U2098 (N_2098,N_1824,N_1849);
nand U2099 (N_2099,N_1931,N_1839);
xnor U2100 (N_2100,N_1919,N_1964);
xnor U2101 (N_2101,N_1837,N_1832);
xnor U2102 (N_2102,N_1971,N_1972);
or U2103 (N_2103,N_1869,N_1828);
and U2104 (N_2104,N_1845,N_1807);
xor U2105 (N_2105,N_1846,N_1950);
nor U2106 (N_2106,N_1972,N_1913);
nor U2107 (N_2107,N_1801,N_1847);
or U2108 (N_2108,N_1869,N_1911);
or U2109 (N_2109,N_1986,N_1876);
nand U2110 (N_2110,N_1915,N_1968);
nor U2111 (N_2111,N_1920,N_1898);
or U2112 (N_2112,N_1831,N_1868);
xnor U2113 (N_2113,N_1842,N_1803);
nor U2114 (N_2114,N_1869,N_1804);
xnor U2115 (N_2115,N_1918,N_1850);
xor U2116 (N_2116,N_1913,N_1986);
xnor U2117 (N_2117,N_1848,N_1914);
or U2118 (N_2118,N_1876,N_1975);
and U2119 (N_2119,N_1807,N_1871);
nor U2120 (N_2120,N_1861,N_1838);
and U2121 (N_2121,N_1829,N_1855);
or U2122 (N_2122,N_1818,N_1809);
nor U2123 (N_2123,N_1803,N_1848);
nor U2124 (N_2124,N_1839,N_1831);
nor U2125 (N_2125,N_1896,N_1920);
xor U2126 (N_2126,N_1907,N_1877);
or U2127 (N_2127,N_1802,N_1835);
or U2128 (N_2128,N_1868,N_1943);
nor U2129 (N_2129,N_1926,N_1900);
nor U2130 (N_2130,N_1880,N_1935);
or U2131 (N_2131,N_1821,N_1968);
or U2132 (N_2132,N_1807,N_1824);
nor U2133 (N_2133,N_1878,N_1967);
or U2134 (N_2134,N_1865,N_1853);
nor U2135 (N_2135,N_1853,N_1806);
xor U2136 (N_2136,N_1862,N_1842);
or U2137 (N_2137,N_1922,N_1870);
or U2138 (N_2138,N_1968,N_1911);
or U2139 (N_2139,N_1833,N_1928);
xnor U2140 (N_2140,N_1875,N_1915);
xnor U2141 (N_2141,N_1907,N_1951);
nand U2142 (N_2142,N_1978,N_1825);
or U2143 (N_2143,N_1909,N_1821);
nand U2144 (N_2144,N_1814,N_1926);
nand U2145 (N_2145,N_1982,N_1947);
and U2146 (N_2146,N_1926,N_1843);
xnor U2147 (N_2147,N_1872,N_1810);
nand U2148 (N_2148,N_1906,N_1884);
xnor U2149 (N_2149,N_1849,N_1882);
nor U2150 (N_2150,N_1855,N_1828);
nand U2151 (N_2151,N_1880,N_1892);
nand U2152 (N_2152,N_1951,N_1821);
xor U2153 (N_2153,N_1925,N_1861);
nor U2154 (N_2154,N_1805,N_1859);
and U2155 (N_2155,N_1818,N_1821);
nor U2156 (N_2156,N_1892,N_1877);
and U2157 (N_2157,N_1910,N_1847);
nand U2158 (N_2158,N_1855,N_1887);
nand U2159 (N_2159,N_1822,N_1809);
or U2160 (N_2160,N_1824,N_1867);
nor U2161 (N_2161,N_1906,N_1849);
xnor U2162 (N_2162,N_1840,N_1940);
nand U2163 (N_2163,N_1875,N_1835);
xnor U2164 (N_2164,N_1901,N_1994);
nor U2165 (N_2165,N_1810,N_1809);
nand U2166 (N_2166,N_1804,N_1832);
nor U2167 (N_2167,N_1835,N_1966);
and U2168 (N_2168,N_1908,N_1886);
nand U2169 (N_2169,N_1900,N_1869);
xnor U2170 (N_2170,N_1851,N_1820);
and U2171 (N_2171,N_1904,N_1960);
xnor U2172 (N_2172,N_1884,N_1887);
xnor U2173 (N_2173,N_1873,N_1848);
nand U2174 (N_2174,N_1902,N_1815);
xor U2175 (N_2175,N_1856,N_1895);
nand U2176 (N_2176,N_1873,N_1912);
nand U2177 (N_2177,N_1868,N_1830);
or U2178 (N_2178,N_1845,N_1851);
and U2179 (N_2179,N_1840,N_1970);
xor U2180 (N_2180,N_1885,N_1802);
nor U2181 (N_2181,N_1903,N_1970);
and U2182 (N_2182,N_1980,N_1944);
and U2183 (N_2183,N_1897,N_1986);
xor U2184 (N_2184,N_1856,N_1855);
nor U2185 (N_2185,N_1998,N_1878);
or U2186 (N_2186,N_1935,N_1806);
and U2187 (N_2187,N_1808,N_1850);
nand U2188 (N_2188,N_1910,N_1915);
nand U2189 (N_2189,N_1837,N_1980);
or U2190 (N_2190,N_1872,N_1882);
xor U2191 (N_2191,N_1907,N_1803);
nor U2192 (N_2192,N_1822,N_1817);
or U2193 (N_2193,N_1974,N_1803);
or U2194 (N_2194,N_1983,N_1841);
nand U2195 (N_2195,N_1835,N_1969);
xor U2196 (N_2196,N_1908,N_1855);
and U2197 (N_2197,N_1870,N_1817);
or U2198 (N_2198,N_1981,N_1936);
or U2199 (N_2199,N_1885,N_1892);
and U2200 (N_2200,N_2107,N_2043);
nand U2201 (N_2201,N_2193,N_2170);
and U2202 (N_2202,N_2182,N_2060);
nor U2203 (N_2203,N_2097,N_2013);
nor U2204 (N_2204,N_2184,N_2111);
xor U2205 (N_2205,N_2118,N_2100);
and U2206 (N_2206,N_2044,N_2092);
nand U2207 (N_2207,N_2134,N_2183);
nand U2208 (N_2208,N_2081,N_2130);
and U2209 (N_2209,N_2075,N_2171);
or U2210 (N_2210,N_2147,N_2047);
or U2211 (N_2211,N_2098,N_2051);
nor U2212 (N_2212,N_2096,N_2008);
xor U2213 (N_2213,N_2122,N_2073);
nor U2214 (N_2214,N_2142,N_2007);
and U2215 (N_2215,N_2151,N_2089);
or U2216 (N_2216,N_2058,N_2066);
and U2217 (N_2217,N_2024,N_2093);
xor U2218 (N_2218,N_2131,N_2002);
and U2219 (N_2219,N_2196,N_2037);
nor U2220 (N_2220,N_2119,N_2186);
or U2221 (N_2221,N_2031,N_2138);
and U2222 (N_2222,N_2121,N_2102);
nor U2223 (N_2223,N_2152,N_2115);
xnor U2224 (N_2224,N_2000,N_2195);
nand U2225 (N_2225,N_2156,N_2129);
nor U2226 (N_2226,N_2125,N_2103);
xor U2227 (N_2227,N_2192,N_2133);
nand U2228 (N_2228,N_2128,N_2150);
xor U2229 (N_2229,N_2003,N_2139);
or U2230 (N_2230,N_2021,N_2176);
or U2231 (N_2231,N_2140,N_2114);
nor U2232 (N_2232,N_2095,N_2042);
or U2233 (N_2233,N_2101,N_2076);
or U2234 (N_2234,N_2175,N_2053);
xnor U2235 (N_2235,N_2046,N_2143);
xor U2236 (N_2236,N_2009,N_2070);
xnor U2237 (N_2237,N_2025,N_2030);
xor U2238 (N_2238,N_2079,N_2035);
or U2239 (N_2239,N_2168,N_2157);
and U2240 (N_2240,N_2069,N_2149);
nor U2241 (N_2241,N_2054,N_2127);
nand U2242 (N_2242,N_2136,N_2078);
nor U2243 (N_2243,N_2099,N_2194);
and U2244 (N_2244,N_2029,N_2012);
nand U2245 (N_2245,N_2166,N_2014);
nand U2246 (N_2246,N_2036,N_2191);
and U2247 (N_2247,N_2085,N_2145);
nor U2248 (N_2248,N_2019,N_2006);
or U2249 (N_2249,N_2050,N_2088);
or U2250 (N_2250,N_2023,N_2039);
and U2251 (N_2251,N_2165,N_2056);
nor U2252 (N_2252,N_2072,N_2005);
nand U2253 (N_2253,N_2173,N_2124);
nand U2254 (N_2254,N_2055,N_2162);
nor U2255 (N_2255,N_2155,N_2190);
or U2256 (N_2256,N_2015,N_2163);
or U2257 (N_2257,N_2052,N_2188);
or U2258 (N_2258,N_2179,N_2180);
or U2259 (N_2259,N_2057,N_2197);
and U2260 (N_2260,N_2109,N_2001);
and U2261 (N_2261,N_2068,N_2177);
nor U2262 (N_2262,N_2199,N_2027);
nor U2263 (N_2263,N_2040,N_2105);
nand U2264 (N_2264,N_2126,N_2153);
nor U2265 (N_2265,N_2198,N_2074);
nor U2266 (N_2266,N_2181,N_2032);
nor U2267 (N_2267,N_2110,N_2091);
and U2268 (N_2268,N_2038,N_2067);
and U2269 (N_2269,N_2082,N_2164);
nand U2270 (N_2270,N_2148,N_2059);
nand U2271 (N_2271,N_2094,N_2185);
xnor U2272 (N_2272,N_2049,N_2154);
and U2273 (N_2273,N_2116,N_2187);
or U2274 (N_2274,N_2161,N_2064);
or U2275 (N_2275,N_2087,N_2090);
and U2276 (N_2276,N_2033,N_2004);
nand U2277 (N_2277,N_2174,N_2132);
and U2278 (N_2278,N_2034,N_2062);
xor U2279 (N_2279,N_2144,N_2160);
or U2280 (N_2280,N_2041,N_2084);
or U2281 (N_2281,N_2045,N_2158);
nor U2282 (N_2282,N_2117,N_2086);
nor U2283 (N_2283,N_2071,N_2022);
nand U2284 (N_2284,N_2028,N_2048);
nand U2285 (N_2285,N_2061,N_2167);
nand U2286 (N_2286,N_2113,N_2141);
or U2287 (N_2287,N_2010,N_2172);
and U2288 (N_2288,N_2065,N_2146);
or U2289 (N_2289,N_2063,N_2026);
nor U2290 (N_2290,N_2077,N_2120);
nand U2291 (N_2291,N_2018,N_2016);
nand U2292 (N_2292,N_2169,N_2020);
nor U2293 (N_2293,N_2108,N_2017);
nor U2294 (N_2294,N_2159,N_2178);
nand U2295 (N_2295,N_2011,N_2112);
xnor U2296 (N_2296,N_2104,N_2135);
and U2297 (N_2297,N_2189,N_2106);
nor U2298 (N_2298,N_2123,N_2083);
nor U2299 (N_2299,N_2137,N_2080);
or U2300 (N_2300,N_2189,N_2063);
or U2301 (N_2301,N_2153,N_2103);
nand U2302 (N_2302,N_2098,N_2050);
nand U2303 (N_2303,N_2049,N_2079);
or U2304 (N_2304,N_2122,N_2118);
or U2305 (N_2305,N_2026,N_2155);
nor U2306 (N_2306,N_2042,N_2190);
or U2307 (N_2307,N_2189,N_2179);
and U2308 (N_2308,N_2036,N_2019);
xor U2309 (N_2309,N_2088,N_2123);
xor U2310 (N_2310,N_2180,N_2182);
xor U2311 (N_2311,N_2070,N_2130);
nor U2312 (N_2312,N_2097,N_2087);
xnor U2313 (N_2313,N_2170,N_2027);
nand U2314 (N_2314,N_2166,N_2003);
or U2315 (N_2315,N_2095,N_2165);
and U2316 (N_2316,N_2007,N_2163);
nand U2317 (N_2317,N_2063,N_2049);
and U2318 (N_2318,N_2093,N_2168);
and U2319 (N_2319,N_2189,N_2147);
xor U2320 (N_2320,N_2127,N_2191);
or U2321 (N_2321,N_2079,N_2039);
and U2322 (N_2322,N_2073,N_2113);
nand U2323 (N_2323,N_2133,N_2089);
and U2324 (N_2324,N_2142,N_2092);
nand U2325 (N_2325,N_2080,N_2036);
or U2326 (N_2326,N_2081,N_2083);
and U2327 (N_2327,N_2130,N_2109);
nand U2328 (N_2328,N_2175,N_2121);
nor U2329 (N_2329,N_2063,N_2123);
nand U2330 (N_2330,N_2042,N_2038);
or U2331 (N_2331,N_2098,N_2003);
and U2332 (N_2332,N_2100,N_2119);
xnor U2333 (N_2333,N_2048,N_2176);
nor U2334 (N_2334,N_2126,N_2023);
xnor U2335 (N_2335,N_2000,N_2056);
xnor U2336 (N_2336,N_2086,N_2112);
or U2337 (N_2337,N_2032,N_2005);
and U2338 (N_2338,N_2163,N_2194);
nand U2339 (N_2339,N_2161,N_2008);
and U2340 (N_2340,N_2136,N_2073);
and U2341 (N_2341,N_2122,N_2026);
or U2342 (N_2342,N_2175,N_2090);
or U2343 (N_2343,N_2127,N_2153);
xor U2344 (N_2344,N_2166,N_2174);
nor U2345 (N_2345,N_2161,N_2013);
xor U2346 (N_2346,N_2056,N_2052);
or U2347 (N_2347,N_2069,N_2030);
nand U2348 (N_2348,N_2065,N_2098);
xor U2349 (N_2349,N_2115,N_2082);
nand U2350 (N_2350,N_2060,N_2107);
and U2351 (N_2351,N_2163,N_2051);
xnor U2352 (N_2352,N_2027,N_2030);
nand U2353 (N_2353,N_2195,N_2030);
nand U2354 (N_2354,N_2102,N_2035);
xnor U2355 (N_2355,N_2091,N_2114);
or U2356 (N_2356,N_2111,N_2082);
xor U2357 (N_2357,N_2059,N_2161);
nor U2358 (N_2358,N_2092,N_2089);
and U2359 (N_2359,N_2146,N_2086);
and U2360 (N_2360,N_2013,N_2131);
nor U2361 (N_2361,N_2135,N_2011);
or U2362 (N_2362,N_2023,N_2137);
xnor U2363 (N_2363,N_2142,N_2058);
nand U2364 (N_2364,N_2012,N_2103);
and U2365 (N_2365,N_2072,N_2006);
nor U2366 (N_2366,N_2119,N_2135);
xor U2367 (N_2367,N_2162,N_2053);
nand U2368 (N_2368,N_2070,N_2083);
nor U2369 (N_2369,N_2153,N_2145);
nor U2370 (N_2370,N_2075,N_2009);
xnor U2371 (N_2371,N_2002,N_2096);
and U2372 (N_2372,N_2173,N_2022);
xor U2373 (N_2373,N_2061,N_2005);
nor U2374 (N_2374,N_2018,N_2019);
and U2375 (N_2375,N_2009,N_2151);
nor U2376 (N_2376,N_2128,N_2101);
nand U2377 (N_2377,N_2172,N_2070);
and U2378 (N_2378,N_2157,N_2131);
nor U2379 (N_2379,N_2084,N_2191);
nand U2380 (N_2380,N_2070,N_2164);
nor U2381 (N_2381,N_2087,N_2049);
nor U2382 (N_2382,N_2188,N_2085);
and U2383 (N_2383,N_2035,N_2052);
or U2384 (N_2384,N_2169,N_2007);
nor U2385 (N_2385,N_2107,N_2042);
or U2386 (N_2386,N_2036,N_2114);
xnor U2387 (N_2387,N_2152,N_2126);
and U2388 (N_2388,N_2058,N_2018);
xnor U2389 (N_2389,N_2024,N_2030);
nor U2390 (N_2390,N_2003,N_2063);
xor U2391 (N_2391,N_2086,N_2158);
and U2392 (N_2392,N_2017,N_2157);
and U2393 (N_2393,N_2130,N_2047);
xnor U2394 (N_2394,N_2168,N_2086);
nor U2395 (N_2395,N_2047,N_2104);
or U2396 (N_2396,N_2125,N_2194);
nand U2397 (N_2397,N_2062,N_2074);
xor U2398 (N_2398,N_2110,N_2033);
nand U2399 (N_2399,N_2131,N_2034);
nor U2400 (N_2400,N_2334,N_2286);
xnor U2401 (N_2401,N_2277,N_2318);
and U2402 (N_2402,N_2364,N_2230);
and U2403 (N_2403,N_2288,N_2280);
or U2404 (N_2404,N_2217,N_2293);
xnor U2405 (N_2405,N_2335,N_2250);
nor U2406 (N_2406,N_2300,N_2238);
nor U2407 (N_2407,N_2313,N_2207);
or U2408 (N_2408,N_2257,N_2330);
and U2409 (N_2409,N_2392,N_2348);
nor U2410 (N_2410,N_2247,N_2393);
and U2411 (N_2411,N_2235,N_2315);
xnor U2412 (N_2412,N_2360,N_2397);
xnor U2413 (N_2413,N_2345,N_2273);
xnor U2414 (N_2414,N_2203,N_2279);
xnor U2415 (N_2415,N_2284,N_2375);
nand U2416 (N_2416,N_2222,N_2248);
nor U2417 (N_2417,N_2385,N_2371);
or U2418 (N_2418,N_2256,N_2304);
xor U2419 (N_2419,N_2218,N_2295);
or U2420 (N_2420,N_2359,N_2326);
or U2421 (N_2421,N_2249,N_2339);
and U2422 (N_2422,N_2316,N_2261);
xnor U2423 (N_2423,N_2283,N_2213);
nand U2424 (N_2424,N_2387,N_2240);
xnor U2425 (N_2425,N_2351,N_2308);
and U2426 (N_2426,N_2281,N_2252);
or U2427 (N_2427,N_2206,N_2390);
nand U2428 (N_2428,N_2357,N_2366);
xor U2429 (N_2429,N_2242,N_2377);
nor U2430 (N_2430,N_2205,N_2299);
or U2431 (N_2431,N_2241,N_2204);
or U2432 (N_2432,N_2341,N_2297);
or U2433 (N_2433,N_2228,N_2278);
and U2434 (N_2434,N_2368,N_2322);
nand U2435 (N_2435,N_2285,N_2232);
xor U2436 (N_2436,N_2225,N_2275);
xnor U2437 (N_2437,N_2337,N_2216);
nand U2438 (N_2438,N_2386,N_2263);
xor U2439 (N_2439,N_2374,N_2290);
xnor U2440 (N_2440,N_2255,N_2201);
or U2441 (N_2441,N_2219,N_2254);
xnor U2442 (N_2442,N_2226,N_2289);
nand U2443 (N_2443,N_2271,N_2258);
xor U2444 (N_2444,N_2323,N_2391);
nand U2445 (N_2445,N_2269,N_2296);
xor U2446 (N_2446,N_2233,N_2331);
and U2447 (N_2447,N_2298,N_2262);
nor U2448 (N_2448,N_2378,N_2311);
xnor U2449 (N_2449,N_2245,N_2350);
xor U2450 (N_2450,N_2363,N_2381);
xor U2451 (N_2451,N_2354,N_2200);
or U2452 (N_2452,N_2314,N_2212);
nand U2453 (N_2453,N_2367,N_2399);
and U2454 (N_2454,N_2382,N_2292);
nand U2455 (N_2455,N_2265,N_2383);
nor U2456 (N_2456,N_2264,N_2272);
nand U2457 (N_2457,N_2353,N_2352);
nand U2458 (N_2458,N_2342,N_2398);
and U2459 (N_2459,N_2343,N_2224);
xor U2460 (N_2460,N_2389,N_2356);
or U2461 (N_2461,N_2302,N_2324);
and U2462 (N_2462,N_2347,N_2332);
and U2463 (N_2463,N_2303,N_2291);
xor U2464 (N_2464,N_2319,N_2394);
nand U2465 (N_2465,N_2236,N_2346);
nor U2466 (N_2466,N_2294,N_2325);
nand U2467 (N_2467,N_2307,N_2376);
nor U2468 (N_2468,N_2395,N_2305);
nand U2469 (N_2469,N_2333,N_2329);
nand U2470 (N_2470,N_2361,N_2251);
nand U2471 (N_2471,N_2287,N_2220);
nand U2472 (N_2472,N_2349,N_2202);
and U2473 (N_2473,N_2328,N_2301);
xor U2474 (N_2474,N_2253,N_2215);
and U2475 (N_2475,N_2210,N_2384);
and U2476 (N_2476,N_2372,N_2380);
xor U2477 (N_2477,N_2358,N_2336);
nor U2478 (N_2478,N_2355,N_2246);
xnor U2479 (N_2479,N_2327,N_2365);
nand U2480 (N_2480,N_2211,N_2270);
nor U2481 (N_2481,N_2369,N_2309);
nor U2482 (N_2482,N_2306,N_2231);
xnor U2483 (N_2483,N_2370,N_2320);
or U2484 (N_2484,N_2379,N_2234);
nand U2485 (N_2485,N_2243,N_2338);
xnor U2486 (N_2486,N_2310,N_2396);
nand U2487 (N_2487,N_2340,N_2260);
nor U2488 (N_2488,N_2282,N_2237);
nand U2489 (N_2489,N_2317,N_2266);
nand U2490 (N_2490,N_2208,N_2373);
xnor U2491 (N_2491,N_2388,N_2362);
and U2492 (N_2492,N_2227,N_2214);
xor U2493 (N_2493,N_2267,N_2321);
or U2494 (N_2494,N_2244,N_2223);
xnor U2495 (N_2495,N_2259,N_2239);
xnor U2496 (N_2496,N_2229,N_2344);
nand U2497 (N_2497,N_2276,N_2312);
or U2498 (N_2498,N_2274,N_2221);
or U2499 (N_2499,N_2268,N_2209);
and U2500 (N_2500,N_2254,N_2210);
or U2501 (N_2501,N_2280,N_2334);
nand U2502 (N_2502,N_2354,N_2253);
xnor U2503 (N_2503,N_2318,N_2289);
or U2504 (N_2504,N_2224,N_2220);
nor U2505 (N_2505,N_2202,N_2311);
or U2506 (N_2506,N_2389,N_2238);
and U2507 (N_2507,N_2285,N_2336);
nor U2508 (N_2508,N_2258,N_2355);
and U2509 (N_2509,N_2359,N_2242);
or U2510 (N_2510,N_2289,N_2326);
nor U2511 (N_2511,N_2204,N_2244);
nor U2512 (N_2512,N_2322,N_2307);
xor U2513 (N_2513,N_2233,N_2392);
nor U2514 (N_2514,N_2240,N_2216);
nand U2515 (N_2515,N_2212,N_2275);
nand U2516 (N_2516,N_2365,N_2342);
xnor U2517 (N_2517,N_2289,N_2393);
nor U2518 (N_2518,N_2237,N_2248);
xnor U2519 (N_2519,N_2357,N_2258);
nor U2520 (N_2520,N_2311,N_2201);
or U2521 (N_2521,N_2287,N_2339);
xor U2522 (N_2522,N_2288,N_2204);
nor U2523 (N_2523,N_2274,N_2257);
and U2524 (N_2524,N_2365,N_2241);
or U2525 (N_2525,N_2322,N_2293);
xor U2526 (N_2526,N_2265,N_2385);
xnor U2527 (N_2527,N_2336,N_2315);
xnor U2528 (N_2528,N_2329,N_2221);
or U2529 (N_2529,N_2371,N_2279);
xnor U2530 (N_2530,N_2399,N_2236);
xnor U2531 (N_2531,N_2202,N_2203);
xnor U2532 (N_2532,N_2220,N_2382);
and U2533 (N_2533,N_2342,N_2253);
nand U2534 (N_2534,N_2348,N_2230);
xor U2535 (N_2535,N_2331,N_2215);
and U2536 (N_2536,N_2394,N_2376);
xor U2537 (N_2537,N_2279,N_2398);
xor U2538 (N_2538,N_2384,N_2223);
nand U2539 (N_2539,N_2392,N_2365);
nor U2540 (N_2540,N_2367,N_2215);
nand U2541 (N_2541,N_2311,N_2277);
nand U2542 (N_2542,N_2337,N_2275);
nor U2543 (N_2543,N_2281,N_2208);
xor U2544 (N_2544,N_2356,N_2304);
or U2545 (N_2545,N_2326,N_2261);
nor U2546 (N_2546,N_2377,N_2294);
and U2547 (N_2547,N_2375,N_2334);
nand U2548 (N_2548,N_2335,N_2279);
or U2549 (N_2549,N_2340,N_2221);
and U2550 (N_2550,N_2308,N_2273);
xor U2551 (N_2551,N_2207,N_2324);
or U2552 (N_2552,N_2379,N_2323);
and U2553 (N_2553,N_2397,N_2253);
xor U2554 (N_2554,N_2257,N_2346);
and U2555 (N_2555,N_2318,N_2216);
and U2556 (N_2556,N_2222,N_2206);
or U2557 (N_2557,N_2304,N_2353);
xor U2558 (N_2558,N_2348,N_2382);
or U2559 (N_2559,N_2338,N_2284);
and U2560 (N_2560,N_2353,N_2323);
and U2561 (N_2561,N_2285,N_2299);
xor U2562 (N_2562,N_2292,N_2377);
nand U2563 (N_2563,N_2347,N_2363);
nand U2564 (N_2564,N_2272,N_2284);
or U2565 (N_2565,N_2244,N_2356);
xnor U2566 (N_2566,N_2306,N_2364);
and U2567 (N_2567,N_2299,N_2275);
and U2568 (N_2568,N_2399,N_2294);
and U2569 (N_2569,N_2243,N_2317);
nor U2570 (N_2570,N_2373,N_2237);
nand U2571 (N_2571,N_2227,N_2317);
nand U2572 (N_2572,N_2304,N_2334);
and U2573 (N_2573,N_2341,N_2210);
nand U2574 (N_2574,N_2269,N_2276);
xnor U2575 (N_2575,N_2359,N_2383);
and U2576 (N_2576,N_2364,N_2332);
or U2577 (N_2577,N_2266,N_2298);
nand U2578 (N_2578,N_2248,N_2262);
nand U2579 (N_2579,N_2217,N_2221);
or U2580 (N_2580,N_2361,N_2348);
xnor U2581 (N_2581,N_2305,N_2269);
and U2582 (N_2582,N_2214,N_2255);
nor U2583 (N_2583,N_2392,N_2236);
nor U2584 (N_2584,N_2399,N_2391);
or U2585 (N_2585,N_2306,N_2382);
or U2586 (N_2586,N_2396,N_2240);
nand U2587 (N_2587,N_2308,N_2286);
nor U2588 (N_2588,N_2369,N_2264);
nand U2589 (N_2589,N_2237,N_2358);
nor U2590 (N_2590,N_2219,N_2362);
nand U2591 (N_2591,N_2234,N_2239);
nand U2592 (N_2592,N_2360,N_2296);
nor U2593 (N_2593,N_2329,N_2313);
nand U2594 (N_2594,N_2313,N_2288);
nand U2595 (N_2595,N_2265,N_2380);
nor U2596 (N_2596,N_2229,N_2202);
xnor U2597 (N_2597,N_2200,N_2206);
nand U2598 (N_2598,N_2316,N_2236);
nor U2599 (N_2599,N_2273,N_2347);
and U2600 (N_2600,N_2461,N_2580);
nor U2601 (N_2601,N_2459,N_2447);
or U2602 (N_2602,N_2508,N_2587);
nor U2603 (N_2603,N_2460,N_2564);
nand U2604 (N_2604,N_2500,N_2475);
or U2605 (N_2605,N_2555,N_2551);
xor U2606 (N_2606,N_2462,N_2540);
and U2607 (N_2607,N_2570,N_2517);
xor U2608 (N_2608,N_2549,N_2449);
nor U2609 (N_2609,N_2576,N_2512);
and U2610 (N_2610,N_2552,N_2547);
or U2611 (N_2611,N_2582,N_2424);
xnor U2612 (N_2612,N_2569,N_2521);
nor U2613 (N_2613,N_2450,N_2565);
or U2614 (N_2614,N_2478,N_2581);
or U2615 (N_2615,N_2445,N_2593);
or U2616 (N_2616,N_2527,N_2511);
or U2617 (N_2617,N_2529,N_2488);
nand U2618 (N_2618,N_2453,N_2448);
xor U2619 (N_2619,N_2573,N_2400);
nor U2620 (N_2620,N_2544,N_2413);
nor U2621 (N_2621,N_2480,N_2531);
nor U2622 (N_2622,N_2458,N_2572);
xnor U2623 (N_2623,N_2454,N_2416);
and U2624 (N_2624,N_2430,N_2410);
or U2625 (N_2625,N_2437,N_2492);
xnor U2626 (N_2626,N_2466,N_2423);
nand U2627 (N_2627,N_2446,N_2510);
nand U2628 (N_2628,N_2441,N_2487);
nand U2629 (N_2629,N_2420,N_2477);
and U2630 (N_2630,N_2401,N_2473);
nand U2631 (N_2631,N_2496,N_2451);
or U2632 (N_2632,N_2495,N_2405);
nand U2633 (N_2633,N_2426,N_2556);
and U2634 (N_2634,N_2403,N_2548);
and U2635 (N_2635,N_2428,N_2502);
or U2636 (N_2636,N_2546,N_2474);
or U2637 (N_2637,N_2559,N_2452);
or U2638 (N_2638,N_2463,N_2408);
nand U2639 (N_2639,N_2493,N_2585);
nand U2640 (N_2640,N_2439,N_2586);
nand U2641 (N_2641,N_2505,N_2524);
and U2642 (N_2642,N_2592,N_2421);
nor U2643 (N_2643,N_2516,N_2434);
or U2644 (N_2644,N_2571,N_2519);
nand U2645 (N_2645,N_2543,N_2507);
xor U2646 (N_2646,N_2566,N_2553);
nand U2647 (N_2647,N_2432,N_2407);
nor U2648 (N_2648,N_2442,N_2535);
nor U2649 (N_2649,N_2528,N_2561);
or U2650 (N_2650,N_2594,N_2577);
nor U2651 (N_2651,N_2455,N_2568);
xnor U2652 (N_2652,N_2418,N_2435);
xor U2653 (N_2653,N_2545,N_2412);
or U2654 (N_2654,N_2415,N_2406);
or U2655 (N_2655,N_2563,N_2562);
nand U2656 (N_2656,N_2498,N_2575);
or U2657 (N_2657,N_2425,N_2438);
and U2658 (N_2658,N_2431,N_2444);
nand U2659 (N_2659,N_2479,N_2596);
nor U2660 (N_2660,N_2494,N_2523);
and U2661 (N_2661,N_2491,N_2595);
nand U2662 (N_2662,N_2558,N_2536);
xnor U2663 (N_2663,N_2469,N_2489);
nor U2664 (N_2664,N_2482,N_2530);
and U2665 (N_2665,N_2574,N_2486);
and U2666 (N_2666,N_2579,N_2467);
nand U2667 (N_2667,N_2578,N_2506);
xor U2668 (N_2668,N_2567,N_2541);
and U2669 (N_2669,N_2501,N_2533);
and U2670 (N_2670,N_2422,N_2597);
nand U2671 (N_2671,N_2514,N_2509);
or U2672 (N_2672,N_2537,N_2526);
xnor U2673 (N_2673,N_2542,N_2472);
nor U2674 (N_2674,N_2518,N_2468);
and U2675 (N_2675,N_2598,N_2550);
nor U2676 (N_2676,N_2476,N_2499);
or U2677 (N_2677,N_2554,N_2414);
nand U2678 (N_2678,N_2515,N_2456);
or U2679 (N_2679,N_2470,N_2525);
or U2680 (N_2680,N_2534,N_2590);
xor U2681 (N_2681,N_2539,N_2497);
nor U2682 (N_2682,N_2588,N_2522);
and U2683 (N_2683,N_2599,N_2481);
nor U2684 (N_2684,N_2411,N_2429);
nor U2685 (N_2685,N_2591,N_2584);
or U2686 (N_2686,N_2433,N_2490);
nand U2687 (N_2687,N_2513,N_2538);
xnor U2688 (N_2688,N_2404,N_2484);
or U2689 (N_2689,N_2483,N_2464);
or U2690 (N_2690,N_2504,N_2583);
and U2691 (N_2691,N_2443,N_2457);
and U2692 (N_2692,N_2503,N_2465);
xor U2693 (N_2693,N_2520,N_2532);
nand U2694 (N_2694,N_2409,N_2471);
nand U2695 (N_2695,N_2485,N_2557);
or U2696 (N_2696,N_2417,N_2440);
xnor U2697 (N_2697,N_2427,N_2436);
and U2698 (N_2698,N_2589,N_2402);
xor U2699 (N_2699,N_2419,N_2560);
or U2700 (N_2700,N_2464,N_2573);
and U2701 (N_2701,N_2596,N_2562);
xor U2702 (N_2702,N_2474,N_2425);
nor U2703 (N_2703,N_2485,N_2443);
and U2704 (N_2704,N_2432,N_2446);
or U2705 (N_2705,N_2476,N_2555);
or U2706 (N_2706,N_2594,N_2414);
xor U2707 (N_2707,N_2481,N_2545);
xnor U2708 (N_2708,N_2460,N_2557);
or U2709 (N_2709,N_2592,N_2594);
or U2710 (N_2710,N_2559,N_2494);
nor U2711 (N_2711,N_2510,N_2410);
nor U2712 (N_2712,N_2555,N_2597);
nand U2713 (N_2713,N_2490,N_2417);
or U2714 (N_2714,N_2442,N_2552);
xor U2715 (N_2715,N_2545,N_2532);
nor U2716 (N_2716,N_2562,N_2457);
nand U2717 (N_2717,N_2417,N_2430);
nor U2718 (N_2718,N_2511,N_2504);
nor U2719 (N_2719,N_2522,N_2518);
xnor U2720 (N_2720,N_2412,N_2506);
nand U2721 (N_2721,N_2406,N_2577);
or U2722 (N_2722,N_2585,N_2522);
xor U2723 (N_2723,N_2432,N_2455);
nor U2724 (N_2724,N_2412,N_2467);
and U2725 (N_2725,N_2425,N_2436);
nor U2726 (N_2726,N_2565,N_2558);
nor U2727 (N_2727,N_2401,N_2547);
nor U2728 (N_2728,N_2465,N_2511);
nand U2729 (N_2729,N_2415,N_2536);
xor U2730 (N_2730,N_2570,N_2494);
and U2731 (N_2731,N_2423,N_2519);
nand U2732 (N_2732,N_2588,N_2548);
nor U2733 (N_2733,N_2459,N_2594);
and U2734 (N_2734,N_2490,N_2584);
and U2735 (N_2735,N_2515,N_2431);
and U2736 (N_2736,N_2493,N_2575);
nand U2737 (N_2737,N_2519,N_2425);
and U2738 (N_2738,N_2591,N_2567);
xor U2739 (N_2739,N_2461,N_2435);
nor U2740 (N_2740,N_2471,N_2519);
xnor U2741 (N_2741,N_2470,N_2435);
nor U2742 (N_2742,N_2490,N_2547);
nand U2743 (N_2743,N_2494,N_2485);
nor U2744 (N_2744,N_2566,N_2534);
xnor U2745 (N_2745,N_2551,N_2498);
and U2746 (N_2746,N_2441,N_2423);
xnor U2747 (N_2747,N_2437,N_2418);
nand U2748 (N_2748,N_2577,N_2547);
nor U2749 (N_2749,N_2573,N_2416);
or U2750 (N_2750,N_2538,N_2439);
nor U2751 (N_2751,N_2505,N_2568);
xnor U2752 (N_2752,N_2482,N_2598);
nand U2753 (N_2753,N_2599,N_2578);
nand U2754 (N_2754,N_2480,N_2563);
nor U2755 (N_2755,N_2529,N_2531);
and U2756 (N_2756,N_2400,N_2592);
nor U2757 (N_2757,N_2516,N_2491);
xnor U2758 (N_2758,N_2597,N_2414);
nand U2759 (N_2759,N_2589,N_2472);
or U2760 (N_2760,N_2443,N_2553);
nor U2761 (N_2761,N_2592,N_2587);
nand U2762 (N_2762,N_2461,N_2558);
xor U2763 (N_2763,N_2585,N_2423);
nand U2764 (N_2764,N_2558,N_2515);
or U2765 (N_2765,N_2415,N_2407);
xor U2766 (N_2766,N_2493,N_2582);
and U2767 (N_2767,N_2592,N_2578);
nand U2768 (N_2768,N_2448,N_2451);
and U2769 (N_2769,N_2546,N_2431);
nand U2770 (N_2770,N_2597,N_2424);
nor U2771 (N_2771,N_2436,N_2523);
xor U2772 (N_2772,N_2488,N_2541);
or U2773 (N_2773,N_2535,N_2541);
nor U2774 (N_2774,N_2417,N_2507);
or U2775 (N_2775,N_2562,N_2597);
nand U2776 (N_2776,N_2564,N_2585);
and U2777 (N_2777,N_2423,N_2421);
nand U2778 (N_2778,N_2573,N_2598);
or U2779 (N_2779,N_2435,N_2414);
nor U2780 (N_2780,N_2558,N_2414);
or U2781 (N_2781,N_2481,N_2408);
and U2782 (N_2782,N_2564,N_2545);
nand U2783 (N_2783,N_2478,N_2493);
nor U2784 (N_2784,N_2438,N_2596);
and U2785 (N_2785,N_2543,N_2546);
nand U2786 (N_2786,N_2495,N_2545);
nor U2787 (N_2787,N_2579,N_2555);
nor U2788 (N_2788,N_2535,N_2544);
nor U2789 (N_2789,N_2497,N_2476);
and U2790 (N_2790,N_2477,N_2527);
nor U2791 (N_2791,N_2405,N_2515);
xor U2792 (N_2792,N_2434,N_2415);
or U2793 (N_2793,N_2496,N_2460);
or U2794 (N_2794,N_2545,N_2538);
nand U2795 (N_2795,N_2474,N_2506);
nor U2796 (N_2796,N_2465,N_2538);
xnor U2797 (N_2797,N_2405,N_2513);
xor U2798 (N_2798,N_2566,N_2512);
and U2799 (N_2799,N_2475,N_2562);
and U2800 (N_2800,N_2665,N_2711);
nand U2801 (N_2801,N_2638,N_2734);
nand U2802 (N_2802,N_2781,N_2780);
nor U2803 (N_2803,N_2691,N_2758);
and U2804 (N_2804,N_2614,N_2624);
or U2805 (N_2805,N_2799,N_2688);
xnor U2806 (N_2806,N_2735,N_2702);
xor U2807 (N_2807,N_2701,N_2766);
or U2808 (N_2808,N_2733,N_2689);
xnor U2809 (N_2809,N_2725,N_2694);
nor U2810 (N_2810,N_2661,N_2706);
and U2811 (N_2811,N_2654,N_2723);
or U2812 (N_2812,N_2622,N_2667);
xnor U2813 (N_2813,N_2732,N_2659);
nand U2814 (N_2814,N_2672,N_2728);
and U2815 (N_2815,N_2745,N_2684);
or U2816 (N_2816,N_2737,N_2721);
and U2817 (N_2817,N_2643,N_2777);
or U2818 (N_2818,N_2754,N_2696);
and U2819 (N_2819,N_2794,N_2646);
and U2820 (N_2820,N_2633,N_2603);
xnor U2821 (N_2821,N_2731,N_2724);
and U2822 (N_2822,N_2783,N_2620);
nor U2823 (N_2823,N_2755,N_2623);
or U2824 (N_2824,N_2615,N_2703);
nand U2825 (N_2825,N_2631,N_2788);
nand U2826 (N_2826,N_2670,N_2768);
xnor U2827 (N_2827,N_2632,N_2704);
nand U2828 (N_2828,N_2769,N_2787);
nand U2829 (N_2829,N_2695,N_2668);
or U2830 (N_2830,N_2729,N_2759);
nand U2831 (N_2831,N_2651,N_2625);
xor U2832 (N_2832,N_2647,N_2678);
xor U2833 (N_2833,N_2714,N_2687);
and U2834 (N_2834,N_2621,N_2772);
or U2835 (N_2835,N_2606,N_2677);
nor U2836 (N_2836,N_2674,N_2685);
or U2837 (N_2837,N_2719,N_2686);
xor U2838 (N_2838,N_2756,N_2792);
nor U2839 (N_2839,N_2717,N_2660);
or U2840 (N_2840,N_2607,N_2690);
nor U2841 (N_2841,N_2644,N_2791);
nand U2842 (N_2842,N_2765,N_2797);
or U2843 (N_2843,N_2736,N_2708);
nor U2844 (N_2844,N_2793,N_2770);
or U2845 (N_2845,N_2753,N_2648);
xnor U2846 (N_2846,N_2602,N_2611);
or U2847 (N_2847,N_2730,N_2612);
and U2848 (N_2848,N_2649,N_2634);
or U2849 (N_2849,N_2776,N_2785);
nor U2850 (N_2850,N_2675,N_2626);
nor U2851 (N_2851,N_2764,N_2786);
nor U2852 (N_2852,N_2739,N_2617);
or U2853 (N_2853,N_2682,N_2742);
and U2854 (N_2854,N_2750,N_2700);
and U2855 (N_2855,N_2662,N_2639);
xor U2856 (N_2856,N_2681,N_2747);
xnor U2857 (N_2857,N_2669,N_2763);
or U2858 (N_2858,N_2705,N_2710);
xor U2859 (N_2859,N_2699,N_2778);
and U2860 (N_2860,N_2743,N_2722);
nand U2861 (N_2861,N_2608,N_2697);
nor U2862 (N_2862,N_2738,N_2746);
xnor U2863 (N_2863,N_2618,N_2653);
xor U2864 (N_2864,N_2679,N_2771);
nor U2865 (N_2865,N_2616,N_2761);
and U2866 (N_2866,N_2671,N_2628);
nand U2867 (N_2867,N_2749,N_2609);
and U2868 (N_2868,N_2605,N_2640);
or U2869 (N_2869,N_2707,N_2666);
nor U2870 (N_2870,N_2664,N_2741);
xor U2871 (N_2871,N_2795,N_2613);
xnor U2872 (N_2872,N_2720,N_2740);
or U2873 (N_2873,N_2782,N_2637);
nand U2874 (N_2874,N_2713,N_2619);
or U2875 (N_2875,N_2709,N_2796);
or U2876 (N_2876,N_2676,N_2757);
and U2877 (N_2877,N_2798,N_2642);
xor U2878 (N_2878,N_2600,N_2760);
and U2879 (N_2879,N_2716,N_2774);
xnor U2880 (N_2880,N_2627,N_2752);
xor U2881 (N_2881,N_2726,N_2784);
nand U2882 (N_2882,N_2635,N_2767);
nor U2883 (N_2883,N_2641,N_2650);
nand U2884 (N_2884,N_2601,N_2673);
or U2885 (N_2885,N_2629,N_2727);
xnor U2886 (N_2886,N_2655,N_2604);
xor U2887 (N_2887,N_2773,N_2658);
and U2888 (N_2888,N_2718,N_2680);
and U2889 (N_2889,N_2610,N_2712);
nor U2890 (N_2890,N_2636,N_2715);
nand U2891 (N_2891,N_2692,N_2656);
nor U2892 (N_2892,N_2657,N_2779);
and U2893 (N_2893,N_2693,N_2645);
or U2894 (N_2894,N_2744,N_2748);
nor U2895 (N_2895,N_2789,N_2652);
and U2896 (N_2896,N_2790,N_2775);
or U2897 (N_2897,N_2698,N_2751);
or U2898 (N_2898,N_2630,N_2663);
or U2899 (N_2899,N_2683,N_2762);
and U2900 (N_2900,N_2664,N_2711);
nand U2901 (N_2901,N_2643,N_2721);
or U2902 (N_2902,N_2614,N_2671);
xor U2903 (N_2903,N_2601,N_2635);
and U2904 (N_2904,N_2645,N_2657);
xnor U2905 (N_2905,N_2640,N_2756);
nand U2906 (N_2906,N_2682,N_2740);
nor U2907 (N_2907,N_2669,N_2758);
xnor U2908 (N_2908,N_2748,N_2781);
or U2909 (N_2909,N_2796,N_2710);
and U2910 (N_2910,N_2633,N_2646);
and U2911 (N_2911,N_2688,N_2609);
or U2912 (N_2912,N_2616,N_2791);
or U2913 (N_2913,N_2654,N_2733);
nor U2914 (N_2914,N_2699,N_2644);
and U2915 (N_2915,N_2789,N_2644);
or U2916 (N_2916,N_2601,N_2756);
and U2917 (N_2917,N_2772,N_2791);
or U2918 (N_2918,N_2785,N_2700);
nor U2919 (N_2919,N_2616,N_2717);
xor U2920 (N_2920,N_2679,N_2742);
and U2921 (N_2921,N_2788,N_2738);
or U2922 (N_2922,N_2714,N_2664);
nor U2923 (N_2923,N_2756,N_2646);
or U2924 (N_2924,N_2795,N_2797);
nand U2925 (N_2925,N_2713,N_2709);
or U2926 (N_2926,N_2682,N_2649);
xnor U2927 (N_2927,N_2700,N_2789);
nor U2928 (N_2928,N_2693,N_2748);
xnor U2929 (N_2929,N_2747,N_2645);
nand U2930 (N_2930,N_2797,N_2675);
nor U2931 (N_2931,N_2780,N_2633);
xor U2932 (N_2932,N_2661,N_2738);
xnor U2933 (N_2933,N_2624,N_2668);
nor U2934 (N_2934,N_2673,N_2647);
and U2935 (N_2935,N_2656,N_2672);
nand U2936 (N_2936,N_2710,N_2628);
nand U2937 (N_2937,N_2721,N_2619);
or U2938 (N_2938,N_2658,N_2673);
xnor U2939 (N_2939,N_2764,N_2674);
and U2940 (N_2940,N_2744,N_2761);
or U2941 (N_2941,N_2637,N_2683);
xor U2942 (N_2942,N_2768,N_2767);
xor U2943 (N_2943,N_2606,N_2612);
nor U2944 (N_2944,N_2778,N_2620);
or U2945 (N_2945,N_2739,N_2713);
nand U2946 (N_2946,N_2763,N_2759);
xor U2947 (N_2947,N_2746,N_2635);
and U2948 (N_2948,N_2619,N_2719);
and U2949 (N_2949,N_2696,N_2690);
nand U2950 (N_2950,N_2749,N_2643);
and U2951 (N_2951,N_2683,N_2712);
xor U2952 (N_2952,N_2739,N_2658);
xor U2953 (N_2953,N_2788,N_2647);
and U2954 (N_2954,N_2722,N_2602);
xnor U2955 (N_2955,N_2668,N_2602);
xor U2956 (N_2956,N_2652,N_2694);
nand U2957 (N_2957,N_2785,N_2730);
nor U2958 (N_2958,N_2689,N_2750);
nor U2959 (N_2959,N_2783,N_2788);
nor U2960 (N_2960,N_2732,N_2655);
or U2961 (N_2961,N_2775,N_2681);
nand U2962 (N_2962,N_2608,N_2667);
and U2963 (N_2963,N_2609,N_2724);
and U2964 (N_2964,N_2767,N_2769);
nand U2965 (N_2965,N_2684,N_2622);
nand U2966 (N_2966,N_2708,N_2707);
and U2967 (N_2967,N_2659,N_2612);
nor U2968 (N_2968,N_2712,N_2600);
xnor U2969 (N_2969,N_2769,N_2750);
or U2970 (N_2970,N_2643,N_2722);
nor U2971 (N_2971,N_2700,N_2677);
and U2972 (N_2972,N_2777,N_2776);
xnor U2973 (N_2973,N_2720,N_2677);
nor U2974 (N_2974,N_2720,N_2797);
nor U2975 (N_2975,N_2781,N_2614);
nor U2976 (N_2976,N_2684,N_2771);
nor U2977 (N_2977,N_2601,N_2662);
and U2978 (N_2978,N_2720,N_2717);
or U2979 (N_2979,N_2629,N_2700);
nand U2980 (N_2980,N_2708,N_2668);
xnor U2981 (N_2981,N_2657,N_2730);
or U2982 (N_2982,N_2790,N_2619);
nor U2983 (N_2983,N_2648,N_2758);
nand U2984 (N_2984,N_2769,N_2707);
xnor U2985 (N_2985,N_2637,N_2605);
and U2986 (N_2986,N_2660,N_2731);
nand U2987 (N_2987,N_2751,N_2679);
nand U2988 (N_2988,N_2713,N_2674);
nor U2989 (N_2989,N_2697,N_2675);
nand U2990 (N_2990,N_2725,N_2652);
or U2991 (N_2991,N_2684,N_2760);
nor U2992 (N_2992,N_2688,N_2794);
xnor U2993 (N_2993,N_2736,N_2608);
and U2994 (N_2994,N_2662,N_2678);
and U2995 (N_2995,N_2634,N_2681);
and U2996 (N_2996,N_2757,N_2619);
nand U2997 (N_2997,N_2733,N_2709);
or U2998 (N_2998,N_2694,N_2763);
xor U2999 (N_2999,N_2794,N_2735);
nand UO_0 (O_0,N_2869,N_2822);
nor UO_1 (O_1,N_2828,N_2809);
and UO_2 (O_2,N_2815,N_2852);
or UO_3 (O_3,N_2948,N_2859);
and UO_4 (O_4,N_2875,N_2977);
nand UO_5 (O_5,N_2965,N_2889);
nor UO_6 (O_6,N_2997,N_2892);
and UO_7 (O_7,N_2934,N_2865);
or UO_8 (O_8,N_2813,N_2998);
xor UO_9 (O_9,N_2970,N_2855);
nand UO_10 (O_10,N_2808,N_2844);
xnor UO_11 (O_11,N_2983,N_2959);
xnor UO_12 (O_12,N_2823,N_2899);
nand UO_13 (O_13,N_2963,N_2898);
nor UO_14 (O_14,N_2818,N_2928);
nand UO_15 (O_15,N_2827,N_2907);
and UO_16 (O_16,N_2924,N_2964);
xor UO_17 (O_17,N_2890,N_2851);
xnor UO_18 (O_18,N_2936,N_2858);
nand UO_19 (O_19,N_2806,N_2939);
or UO_20 (O_20,N_2803,N_2881);
or UO_21 (O_21,N_2863,N_2968);
nand UO_22 (O_22,N_2876,N_2984);
nor UO_23 (O_23,N_2980,N_2807);
or UO_24 (O_24,N_2825,N_2961);
nor UO_25 (O_25,N_2975,N_2868);
and UO_26 (O_26,N_2935,N_2897);
nor UO_27 (O_27,N_2919,N_2882);
and UO_28 (O_28,N_2923,N_2840);
nand UO_29 (O_29,N_2991,N_2916);
nor UO_30 (O_30,N_2930,N_2942);
nor UO_31 (O_31,N_2801,N_2973);
or UO_32 (O_32,N_2888,N_2914);
xnor UO_33 (O_33,N_2837,N_2860);
nand UO_34 (O_34,N_2954,N_2857);
nor UO_35 (O_35,N_2925,N_2812);
nand UO_36 (O_36,N_2960,N_2816);
and UO_37 (O_37,N_2992,N_2943);
and UO_38 (O_38,N_2893,N_2871);
nand UO_39 (O_39,N_2874,N_2901);
or UO_40 (O_40,N_2996,N_2802);
nor UO_41 (O_41,N_2873,N_2955);
nor UO_42 (O_42,N_2938,N_2979);
or UO_43 (O_43,N_2982,N_2969);
or UO_44 (O_44,N_2845,N_2826);
nand UO_45 (O_45,N_2829,N_2995);
nand UO_46 (O_46,N_2946,N_2966);
nor UO_47 (O_47,N_2940,N_2931);
and UO_48 (O_48,N_2832,N_2976);
xnor UO_49 (O_49,N_2842,N_2817);
or UO_50 (O_50,N_2821,N_2841);
nor UO_51 (O_51,N_2985,N_2945);
xnor UO_52 (O_52,N_2835,N_2952);
xnor UO_53 (O_53,N_2911,N_2904);
nor UO_54 (O_54,N_2921,N_2885);
and UO_55 (O_55,N_2953,N_2804);
or UO_56 (O_56,N_2972,N_2879);
or UO_57 (O_57,N_2993,N_2847);
and UO_58 (O_58,N_2917,N_2978);
and UO_59 (O_59,N_2870,N_2974);
xnor UO_60 (O_60,N_2856,N_2805);
and UO_61 (O_61,N_2958,N_2944);
or UO_62 (O_62,N_2932,N_2900);
nand UO_63 (O_63,N_2918,N_2877);
nand UO_64 (O_64,N_2913,N_2849);
nor UO_65 (O_65,N_2846,N_2908);
and UO_66 (O_66,N_2988,N_2800);
nand UO_67 (O_67,N_2867,N_2947);
nor UO_68 (O_68,N_2994,N_2926);
and UO_69 (O_69,N_2937,N_2962);
xor UO_70 (O_70,N_2990,N_2811);
and UO_71 (O_71,N_2912,N_2824);
nor UO_72 (O_72,N_2902,N_2971);
nor UO_73 (O_73,N_2929,N_2820);
and UO_74 (O_74,N_2883,N_2951);
nand UO_75 (O_75,N_2814,N_2895);
nand UO_76 (O_76,N_2880,N_2967);
xor UO_77 (O_77,N_2987,N_2878);
and UO_78 (O_78,N_2862,N_2839);
nand UO_79 (O_79,N_2920,N_2861);
and UO_80 (O_80,N_2941,N_2884);
and UO_81 (O_81,N_2838,N_2886);
nand UO_82 (O_82,N_2887,N_2896);
and UO_83 (O_83,N_2949,N_2866);
nand UO_84 (O_84,N_2905,N_2810);
and UO_85 (O_85,N_2927,N_2872);
and UO_86 (O_86,N_2830,N_2894);
nor UO_87 (O_87,N_2864,N_2909);
nand UO_88 (O_88,N_2956,N_2922);
xor UO_89 (O_89,N_2981,N_2891);
and UO_90 (O_90,N_2834,N_2989);
or UO_91 (O_91,N_2933,N_2906);
and UO_92 (O_92,N_2957,N_2850);
or UO_93 (O_93,N_2819,N_2999);
nor UO_94 (O_94,N_2836,N_2903);
or UO_95 (O_95,N_2833,N_2915);
and UO_96 (O_96,N_2986,N_2910);
nor UO_97 (O_97,N_2848,N_2854);
nand UO_98 (O_98,N_2853,N_2950);
or UO_99 (O_99,N_2843,N_2831);
nand UO_100 (O_100,N_2870,N_2885);
nand UO_101 (O_101,N_2997,N_2879);
or UO_102 (O_102,N_2872,N_2861);
xor UO_103 (O_103,N_2867,N_2989);
nor UO_104 (O_104,N_2891,N_2954);
nor UO_105 (O_105,N_2902,N_2860);
or UO_106 (O_106,N_2909,N_2956);
and UO_107 (O_107,N_2843,N_2801);
or UO_108 (O_108,N_2858,N_2811);
nand UO_109 (O_109,N_2851,N_2961);
nand UO_110 (O_110,N_2876,N_2901);
xnor UO_111 (O_111,N_2979,N_2993);
nand UO_112 (O_112,N_2851,N_2852);
or UO_113 (O_113,N_2920,N_2840);
or UO_114 (O_114,N_2855,N_2933);
and UO_115 (O_115,N_2856,N_2831);
and UO_116 (O_116,N_2871,N_2868);
or UO_117 (O_117,N_2900,N_2916);
nand UO_118 (O_118,N_2803,N_2958);
xnor UO_119 (O_119,N_2938,N_2804);
nor UO_120 (O_120,N_2966,N_2856);
and UO_121 (O_121,N_2933,N_2834);
xor UO_122 (O_122,N_2839,N_2887);
nand UO_123 (O_123,N_2810,N_2935);
xor UO_124 (O_124,N_2859,N_2945);
xnor UO_125 (O_125,N_2949,N_2902);
xor UO_126 (O_126,N_2847,N_2937);
nor UO_127 (O_127,N_2984,N_2964);
xnor UO_128 (O_128,N_2938,N_2994);
or UO_129 (O_129,N_2962,N_2821);
and UO_130 (O_130,N_2826,N_2930);
and UO_131 (O_131,N_2822,N_2809);
or UO_132 (O_132,N_2815,N_2857);
nand UO_133 (O_133,N_2843,N_2841);
nand UO_134 (O_134,N_2903,N_2895);
nand UO_135 (O_135,N_2958,N_2919);
and UO_136 (O_136,N_2907,N_2857);
or UO_137 (O_137,N_2858,N_2826);
xor UO_138 (O_138,N_2827,N_2941);
nor UO_139 (O_139,N_2983,N_2967);
xor UO_140 (O_140,N_2810,N_2840);
xor UO_141 (O_141,N_2802,N_2905);
and UO_142 (O_142,N_2807,N_2837);
xor UO_143 (O_143,N_2986,N_2817);
nand UO_144 (O_144,N_2813,N_2811);
nor UO_145 (O_145,N_2851,N_2892);
nor UO_146 (O_146,N_2970,N_2988);
nand UO_147 (O_147,N_2893,N_2884);
or UO_148 (O_148,N_2864,N_2951);
and UO_149 (O_149,N_2974,N_2841);
xnor UO_150 (O_150,N_2869,N_2968);
xnor UO_151 (O_151,N_2916,N_2896);
nor UO_152 (O_152,N_2923,N_2950);
nor UO_153 (O_153,N_2971,N_2884);
or UO_154 (O_154,N_2839,N_2969);
nand UO_155 (O_155,N_2927,N_2815);
nand UO_156 (O_156,N_2804,N_2961);
or UO_157 (O_157,N_2866,N_2846);
nand UO_158 (O_158,N_2876,N_2856);
and UO_159 (O_159,N_2958,N_2878);
or UO_160 (O_160,N_2811,N_2851);
nor UO_161 (O_161,N_2801,N_2847);
and UO_162 (O_162,N_2930,N_2882);
or UO_163 (O_163,N_2940,N_2863);
and UO_164 (O_164,N_2954,N_2956);
or UO_165 (O_165,N_2984,N_2902);
and UO_166 (O_166,N_2858,N_2925);
nand UO_167 (O_167,N_2927,N_2806);
or UO_168 (O_168,N_2916,N_2985);
nor UO_169 (O_169,N_2864,N_2902);
nand UO_170 (O_170,N_2850,N_2930);
xor UO_171 (O_171,N_2858,N_2971);
nand UO_172 (O_172,N_2894,N_2880);
nand UO_173 (O_173,N_2982,N_2806);
nor UO_174 (O_174,N_2859,N_2977);
nor UO_175 (O_175,N_2892,N_2825);
or UO_176 (O_176,N_2908,N_2902);
or UO_177 (O_177,N_2974,N_2978);
or UO_178 (O_178,N_2975,N_2849);
nor UO_179 (O_179,N_2815,N_2972);
and UO_180 (O_180,N_2886,N_2854);
and UO_181 (O_181,N_2959,N_2925);
or UO_182 (O_182,N_2906,N_2904);
xnor UO_183 (O_183,N_2987,N_2814);
or UO_184 (O_184,N_2813,N_2912);
nor UO_185 (O_185,N_2870,N_2846);
nand UO_186 (O_186,N_2941,N_2950);
xnor UO_187 (O_187,N_2997,N_2880);
or UO_188 (O_188,N_2985,N_2995);
xor UO_189 (O_189,N_2916,N_2827);
or UO_190 (O_190,N_2912,N_2883);
xor UO_191 (O_191,N_2985,N_2934);
nand UO_192 (O_192,N_2807,N_2905);
or UO_193 (O_193,N_2845,N_2974);
or UO_194 (O_194,N_2858,N_2952);
nor UO_195 (O_195,N_2853,N_2841);
xor UO_196 (O_196,N_2931,N_2809);
nand UO_197 (O_197,N_2885,N_2984);
nand UO_198 (O_198,N_2802,N_2920);
and UO_199 (O_199,N_2929,N_2903);
nand UO_200 (O_200,N_2907,N_2957);
nor UO_201 (O_201,N_2823,N_2972);
nor UO_202 (O_202,N_2966,N_2895);
and UO_203 (O_203,N_2889,N_2884);
and UO_204 (O_204,N_2817,N_2947);
nor UO_205 (O_205,N_2873,N_2864);
nand UO_206 (O_206,N_2826,N_2819);
and UO_207 (O_207,N_2903,N_2862);
xor UO_208 (O_208,N_2892,N_2931);
xnor UO_209 (O_209,N_2955,N_2899);
or UO_210 (O_210,N_2808,N_2871);
nor UO_211 (O_211,N_2897,N_2803);
or UO_212 (O_212,N_2928,N_2960);
nand UO_213 (O_213,N_2867,N_2934);
xnor UO_214 (O_214,N_2859,N_2802);
and UO_215 (O_215,N_2805,N_2812);
and UO_216 (O_216,N_2869,N_2818);
nor UO_217 (O_217,N_2801,N_2872);
or UO_218 (O_218,N_2910,N_2931);
and UO_219 (O_219,N_2930,N_2810);
nand UO_220 (O_220,N_2871,N_2823);
nand UO_221 (O_221,N_2953,N_2946);
nand UO_222 (O_222,N_2983,N_2856);
or UO_223 (O_223,N_2892,N_2932);
nor UO_224 (O_224,N_2986,N_2889);
nor UO_225 (O_225,N_2852,N_2920);
xnor UO_226 (O_226,N_2853,N_2953);
nand UO_227 (O_227,N_2990,N_2826);
nand UO_228 (O_228,N_2856,N_2830);
or UO_229 (O_229,N_2920,N_2896);
nor UO_230 (O_230,N_2891,N_2992);
xor UO_231 (O_231,N_2924,N_2828);
nor UO_232 (O_232,N_2866,N_2933);
or UO_233 (O_233,N_2841,N_2973);
nand UO_234 (O_234,N_2850,N_2958);
nor UO_235 (O_235,N_2826,N_2836);
or UO_236 (O_236,N_2920,N_2956);
and UO_237 (O_237,N_2977,N_2966);
and UO_238 (O_238,N_2922,N_2857);
or UO_239 (O_239,N_2894,N_2937);
nand UO_240 (O_240,N_2980,N_2877);
or UO_241 (O_241,N_2841,N_2872);
or UO_242 (O_242,N_2883,N_2974);
nand UO_243 (O_243,N_2852,N_2802);
xnor UO_244 (O_244,N_2941,N_2857);
nand UO_245 (O_245,N_2937,N_2872);
or UO_246 (O_246,N_2864,N_2863);
or UO_247 (O_247,N_2925,N_2951);
or UO_248 (O_248,N_2815,N_2969);
nor UO_249 (O_249,N_2969,N_2800);
xnor UO_250 (O_250,N_2821,N_2900);
nand UO_251 (O_251,N_2969,N_2931);
and UO_252 (O_252,N_2967,N_2900);
xor UO_253 (O_253,N_2819,N_2937);
or UO_254 (O_254,N_2992,N_2980);
nor UO_255 (O_255,N_2881,N_2998);
and UO_256 (O_256,N_2869,N_2998);
xnor UO_257 (O_257,N_2947,N_2987);
or UO_258 (O_258,N_2825,N_2882);
nor UO_259 (O_259,N_2833,N_2871);
xnor UO_260 (O_260,N_2843,N_2952);
and UO_261 (O_261,N_2832,N_2967);
nor UO_262 (O_262,N_2896,N_2985);
xor UO_263 (O_263,N_2824,N_2809);
and UO_264 (O_264,N_2950,N_2846);
and UO_265 (O_265,N_2941,N_2930);
or UO_266 (O_266,N_2982,N_2999);
nand UO_267 (O_267,N_2990,N_2926);
or UO_268 (O_268,N_2802,N_2882);
nor UO_269 (O_269,N_2950,N_2891);
nand UO_270 (O_270,N_2997,N_2946);
nand UO_271 (O_271,N_2855,N_2995);
and UO_272 (O_272,N_2808,N_2946);
nand UO_273 (O_273,N_2969,N_2947);
nand UO_274 (O_274,N_2883,N_2815);
xnor UO_275 (O_275,N_2866,N_2821);
or UO_276 (O_276,N_2842,N_2924);
or UO_277 (O_277,N_2843,N_2826);
xor UO_278 (O_278,N_2909,N_2994);
or UO_279 (O_279,N_2872,N_2855);
nor UO_280 (O_280,N_2805,N_2981);
or UO_281 (O_281,N_2821,N_2992);
nor UO_282 (O_282,N_2863,N_2820);
xnor UO_283 (O_283,N_2855,N_2993);
and UO_284 (O_284,N_2940,N_2913);
or UO_285 (O_285,N_2884,N_2802);
and UO_286 (O_286,N_2941,N_2902);
or UO_287 (O_287,N_2984,N_2992);
nor UO_288 (O_288,N_2820,N_2806);
and UO_289 (O_289,N_2803,N_2864);
or UO_290 (O_290,N_2985,N_2888);
nor UO_291 (O_291,N_2880,N_2810);
or UO_292 (O_292,N_2845,N_2980);
nand UO_293 (O_293,N_2997,N_2840);
nor UO_294 (O_294,N_2981,N_2957);
or UO_295 (O_295,N_2838,N_2937);
or UO_296 (O_296,N_2891,N_2837);
xnor UO_297 (O_297,N_2858,N_2889);
or UO_298 (O_298,N_2953,N_2975);
nor UO_299 (O_299,N_2894,N_2893);
nor UO_300 (O_300,N_2827,N_2894);
or UO_301 (O_301,N_2985,N_2847);
nand UO_302 (O_302,N_2933,N_2909);
or UO_303 (O_303,N_2881,N_2817);
xnor UO_304 (O_304,N_2831,N_2936);
and UO_305 (O_305,N_2973,N_2810);
nand UO_306 (O_306,N_2977,N_2931);
and UO_307 (O_307,N_2882,N_2891);
xor UO_308 (O_308,N_2914,N_2810);
nor UO_309 (O_309,N_2938,N_2829);
nand UO_310 (O_310,N_2986,N_2812);
nor UO_311 (O_311,N_2944,N_2917);
or UO_312 (O_312,N_2913,N_2827);
or UO_313 (O_313,N_2849,N_2888);
and UO_314 (O_314,N_2855,N_2852);
nand UO_315 (O_315,N_2838,N_2826);
nand UO_316 (O_316,N_2975,N_2902);
or UO_317 (O_317,N_2846,N_2860);
xnor UO_318 (O_318,N_2923,N_2954);
and UO_319 (O_319,N_2962,N_2842);
xor UO_320 (O_320,N_2942,N_2940);
and UO_321 (O_321,N_2804,N_2806);
xor UO_322 (O_322,N_2852,N_2894);
and UO_323 (O_323,N_2869,N_2957);
nand UO_324 (O_324,N_2992,N_2844);
xnor UO_325 (O_325,N_2990,N_2855);
nor UO_326 (O_326,N_2954,N_2806);
xnor UO_327 (O_327,N_2996,N_2815);
nand UO_328 (O_328,N_2993,N_2833);
and UO_329 (O_329,N_2866,N_2850);
and UO_330 (O_330,N_2829,N_2813);
nand UO_331 (O_331,N_2817,N_2877);
xnor UO_332 (O_332,N_2961,N_2891);
or UO_333 (O_333,N_2900,N_2857);
xnor UO_334 (O_334,N_2805,N_2914);
or UO_335 (O_335,N_2961,N_2809);
or UO_336 (O_336,N_2906,N_2845);
and UO_337 (O_337,N_2817,N_2882);
and UO_338 (O_338,N_2920,N_2898);
nand UO_339 (O_339,N_2931,N_2831);
nor UO_340 (O_340,N_2849,N_2988);
or UO_341 (O_341,N_2937,N_2903);
nand UO_342 (O_342,N_2848,N_2872);
nor UO_343 (O_343,N_2946,N_2802);
or UO_344 (O_344,N_2981,N_2848);
nor UO_345 (O_345,N_2990,N_2909);
nor UO_346 (O_346,N_2966,N_2876);
nor UO_347 (O_347,N_2894,N_2828);
nand UO_348 (O_348,N_2912,N_2875);
or UO_349 (O_349,N_2863,N_2949);
nor UO_350 (O_350,N_2842,N_2923);
or UO_351 (O_351,N_2872,N_2943);
xor UO_352 (O_352,N_2919,N_2902);
nor UO_353 (O_353,N_2852,N_2864);
or UO_354 (O_354,N_2848,N_2957);
nor UO_355 (O_355,N_2938,N_2902);
nor UO_356 (O_356,N_2899,N_2849);
nand UO_357 (O_357,N_2875,N_2902);
and UO_358 (O_358,N_2818,N_2857);
and UO_359 (O_359,N_2843,N_2943);
xnor UO_360 (O_360,N_2982,N_2836);
xor UO_361 (O_361,N_2896,N_2974);
or UO_362 (O_362,N_2803,N_2911);
nand UO_363 (O_363,N_2982,N_2960);
nand UO_364 (O_364,N_2931,N_2980);
nor UO_365 (O_365,N_2803,N_2984);
nand UO_366 (O_366,N_2881,N_2807);
nor UO_367 (O_367,N_2882,N_2929);
or UO_368 (O_368,N_2840,N_2996);
and UO_369 (O_369,N_2928,N_2863);
xnor UO_370 (O_370,N_2871,N_2932);
nor UO_371 (O_371,N_2985,N_2981);
or UO_372 (O_372,N_2960,N_2891);
xor UO_373 (O_373,N_2869,N_2933);
nor UO_374 (O_374,N_2913,N_2944);
nor UO_375 (O_375,N_2821,N_2869);
xor UO_376 (O_376,N_2829,N_2942);
nand UO_377 (O_377,N_2872,N_2858);
xor UO_378 (O_378,N_2926,N_2813);
xor UO_379 (O_379,N_2925,N_2841);
and UO_380 (O_380,N_2965,N_2903);
nand UO_381 (O_381,N_2906,N_2920);
or UO_382 (O_382,N_2957,N_2949);
nor UO_383 (O_383,N_2841,N_2929);
xnor UO_384 (O_384,N_2987,N_2929);
and UO_385 (O_385,N_2893,N_2827);
nand UO_386 (O_386,N_2865,N_2933);
nor UO_387 (O_387,N_2990,N_2907);
nor UO_388 (O_388,N_2996,N_2909);
xor UO_389 (O_389,N_2896,N_2907);
nor UO_390 (O_390,N_2916,N_2978);
xnor UO_391 (O_391,N_2949,N_2950);
nand UO_392 (O_392,N_2948,N_2938);
nor UO_393 (O_393,N_2825,N_2939);
nand UO_394 (O_394,N_2992,N_2956);
nor UO_395 (O_395,N_2821,N_2879);
xor UO_396 (O_396,N_2988,N_2976);
nand UO_397 (O_397,N_2960,N_2815);
nor UO_398 (O_398,N_2843,N_2852);
and UO_399 (O_399,N_2954,N_2820);
or UO_400 (O_400,N_2944,N_2994);
xnor UO_401 (O_401,N_2921,N_2816);
xnor UO_402 (O_402,N_2924,N_2876);
xnor UO_403 (O_403,N_2986,N_2953);
nand UO_404 (O_404,N_2992,N_2853);
nand UO_405 (O_405,N_2809,N_2976);
xor UO_406 (O_406,N_2906,N_2883);
xor UO_407 (O_407,N_2952,N_2819);
nor UO_408 (O_408,N_2943,N_2965);
and UO_409 (O_409,N_2881,N_2851);
or UO_410 (O_410,N_2938,N_2876);
xnor UO_411 (O_411,N_2957,N_2822);
nor UO_412 (O_412,N_2929,N_2857);
nand UO_413 (O_413,N_2812,N_2905);
xnor UO_414 (O_414,N_2843,N_2913);
and UO_415 (O_415,N_2969,N_2875);
nand UO_416 (O_416,N_2914,N_2847);
or UO_417 (O_417,N_2818,N_2805);
and UO_418 (O_418,N_2942,N_2837);
and UO_419 (O_419,N_2990,N_2891);
nand UO_420 (O_420,N_2873,N_2889);
or UO_421 (O_421,N_2929,N_2931);
nor UO_422 (O_422,N_2899,N_2931);
or UO_423 (O_423,N_2861,N_2895);
or UO_424 (O_424,N_2914,N_2843);
nor UO_425 (O_425,N_2955,N_2816);
xor UO_426 (O_426,N_2882,N_2986);
and UO_427 (O_427,N_2842,N_2833);
nor UO_428 (O_428,N_2921,N_2981);
or UO_429 (O_429,N_2882,N_2844);
xor UO_430 (O_430,N_2810,N_2981);
and UO_431 (O_431,N_2969,N_2963);
nor UO_432 (O_432,N_2890,N_2814);
and UO_433 (O_433,N_2983,N_2867);
xnor UO_434 (O_434,N_2820,N_2969);
or UO_435 (O_435,N_2925,N_2806);
nor UO_436 (O_436,N_2809,N_2950);
or UO_437 (O_437,N_2852,N_2916);
or UO_438 (O_438,N_2875,N_2854);
nor UO_439 (O_439,N_2905,N_2805);
and UO_440 (O_440,N_2912,N_2907);
xnor UO_441 (O_441,N_2910,N_2892);
or UO_442 (O_442,N_2855,N_2897);
xnor UO_443 (O_443,N_2914,N_2961);
and UO_444 (O_444,N_2815,N_2806);
nand UO_445 (O_445,N_2970,N_2858);
nand UO_446 (O_446,N_2850,N_2959);
xnor UO_447 (O_447,N_2872,N_2916);
nand UO_448 (O_448,N_2992,N_2807);
xor UO_449 (O_449,N_2800,N_2868);
nor UO_450 (O_450,N_2857,N_2968);
and UO_451 (O_451,N_2972,N_2813);
nand UO_452 (O_452,N_2849,N_2937);
nand UO_453 (O_453,N_2833,N_2921);
xnor UO_454 (O_454,N_2820,N_2831);
xor UO_455 (O_455,N_2933,N_2985);
nand UO_456 (O_456,N_2842,N_2875);
nor UO_457 (O_457,N_2891,N_2804);
nand UO_458 (O_458,N_2827,N_2859);
nand UO_459 (O_459,N_2940,N_2807);
nand UO_460 (O_460,N_2999,N_2817);
nand UO_461 (O_461,N_2809,N_2881);
and UO_462 (O_462,N_2910,N_2974);
nand UO_463 (O_463,N_2993,N_2885);
or UO_464 (O_464,N_2819,N_2912);
nand UO_465 (O_465,N_2818,N_2971);
nor UO_466 (O_466,N_2821,N_2985);
nand UO_467 (O_467,N_2981,N_2858);
nand UO_468 (O_468,N_2818,N_2945);
nand UO_469 (O_469,N_2866,N_2894);
xnor UO_470 (O_470,N_2989,N_2984);
nand UO_471 (O_471,N_2874,N_2852);
nand UO_472 (O_472,N_2837,N_2828);
nand UO_473 (O_473,N_2932,N_2814);
nand UO_474 (O_474,N_2826,N_2938);
xnor UO_475 (O_475,N_2945,N_2965);
or UO_476 (O_476,N_2933,N_2986);
and UO_477 (O_477,N_2984,N_2806);
xnor UO_478 (O_478,N_2870,N_2949);
nand UO_479 (O_479,N_2922,N_2816);
and UO_480 (O_480,N_2970,N_2831);
and UO_481 (O_481,N_2917,N_2956);
xnor UO_482 (O_482,N_2867,N_2848);
nand UO_483 (O_483,N_2841,N_2986);
or UO_484 (O_484,N_2997,N_2902);
or UO_485 (O_485,N_2870,N_2930);
and UO_486 (O_486,N_2941,N_2901);
nand UO_487 (O_487,N_2988,N_2953);
nor UO_488 (O_488,N_2936,N_2886);
nand UO_489 (O_489,N_2882,N_2890);
or UO_490 (O_490,N_2978,N_2989);
and UO_491 (O_491,N_2895,N_2949);
xnor UO_492 (O_492,N_2973,N_2915);
or UO_493 (O_493,N_2839,N_2919);
xor UO_494 (O_494,N_2993,N_2843);
xnor UO_495 (O_495,N_2859,N_2923);
and UO_496 (O_496,N_2860,N_2810);
or UO_497 (O_497,N_2946,N_2831);
or UO_498 (O_498,N_2800,N_2952);
or UO_499 (O_499,N_2947,N_2877);
endmodule