module basic_500_3000_500_60_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_282,In_228);
or U1 (N_1,In_247,In_489);
nor U2 (N_2,In_288,In_405);
nand U3 (N_3,In_2,In_137);
nor U4 (N_4,In_11,In_145);
or U5 (N_5,In_472,In_172);
and U6 (N_6,In_236,In_360);
and U7 (N_7,In_243,In_264);
nand U8 (N_8,In_469,In_178);
or U9 (N_9,In_182,In_224);
xnor U10 (N_10,In_492,In_81);
nor U11 (N_11,In_412,In_316);
and U12 (N_12,In_50,In_402);
and U13 (N_13,In_349,In_306);
nor U14 (N_14,In_488,In_302);
or U15 (N_15,In_348,In_152);
or U16 (N_16,In_35,In_193);
nor U17 (N_17,In_231,In_209);
and U18 (N_18,In_363,In_387);
or U19 (N_19,In_106,In_205);
nand U20 (N_20,In_221,In_40);
xnor U21 (N_21,In_391,In_68);
and U22 (N_22,In_304,In_338);
or U23 (N_23,In_109,In_263);
or U24 (N_24,In_163,In_21);
nand U25 (N_25,In_173,In_14);
or U26 (N_26,In_158,In_371);
or U27 (N_27,In_426,In_200);
or U28 (N_28,In_162,In_12);
nand U29 (N_29,In_181,In_234);
and U30 (N_30,In_120,In_199);
xnor U31 (N_31,In_83,In_186);
and U32 (N_32,In_429,In_286);
nand U33 (N_33,In_273,In_215);
nand U34 (N_34,In_259,In_127);
or U35 (N_35,In_313,In_317);
nor U36 (N_36,In_277,In_115);
nand U37 (N_37,In_444,In_237);
or U38 (N_38,In_458,In_353);
nand U39 (N_39,In_111,In_157);
or U40 (N_40,In_296,In_93);
or U41 (N_41,In_323,In_256);
or U42 (N_42,In_44,In_250);
and U43 (N_43,In_8,In_98);
or U44 (N_44,In_239,In_122);
or U45 (N_45,In_356,In_188);
or U46 (N_46,In_153,In_142);
or U47 (N_47,In_107,In_89);
nor U48 (N_48,In_419,In_386);
nor U49 (N_49,In_244,In_407);
and U50 (N_50,In_167,In_326);
xor U51 (N_51,In_384,In_150);
nand U52 (N_52,In_357,In_431);
nand U53 (N_53,In_265,In_380);
xnor U54 (N_54,In_97,In_34);
and U55 (N_55,In_342,In_362);
nand U56 (N_56,In_123,In_438);
nand U57 (N_57,In_432,In_379);
or U58 (N_58,In_445,In_132);
or U59 (N_59,In_148,In_245);
nor U60 (N_60,In_38,In_169);
nand U61 (N_61,In_451,In_143);
and U62 (N_62,N_15,In_87);
and U63 (N_63,In_427,In_269);
or U64 (N_64,In_457,In_393);
or U65 (N_65,N_7,In_185);
nor U66 (N_66,In_179,In_227);
nand U67 (N_67,In_77,In_423);
and U68 (N_68,In_26,In_147);
nand U69 (N_69,In_43,In_206);
and U70 (N_70,In_170,In_345);
nor U71 (N_71,In_18,In_389);
nand U72 (N_72,In_203,In_294);
or U73 (N_73,In_494,In_482);
nor U74 (N_74,In_298,In_329);
nor U75 (N_75,In_33,In_71);
or U76 (N_76,In_320,In_351);
nand U77 (N_77,In_110,In_315);
or U78 (N_78,In_411,In_80);
or U79 (N_79,In_382,In_418);
or U80 (N_80,In_156,In_76);
nor U81 (N_81,In_401,In_7);
nor U82 (N_82,In_390,In_108);
nand U83 (N_83,In_271,In_74);
nor U84 (N_84,In_394,In_90);
or U85 (N_85,In_184,In_295);
nor U86 (N_86,In_493,In_210);
and U87 (N_87,In_434,In_254);
and U88 (N_88,N_31,In_216);
xnor U89 (N_89,In_456,In_103);
and U90 (N_90,In_318,In_39);
nor U91 (N_91,In_177,In_481);
xnor U92 (N_92,In_281,In_42);
nor U93 (N_93,In_435,In_60);
nor U94 (N_94,In_129,In_314);
nand U95 (N_95,In_327,In_330);
nand U96 (N_96,In_372,In_113);
or U97 (N_97,In_119,In_450);
nand U98 (N_98,N_30,In_187);
nor U99 (N_99,In_171,In_428);
and U100 (N_100,In_136,In_149);
nand U101 (N_101,In_61,N_79);
or U102 (N_102,In_430,N_88);
nand U103 (N_103,In_219,In_366);
or U104 (N_104,In_91,N_85);
nand U105 (N_105,In_354,In_344);
and U106 (N_106,In_58,N_33);
and U107 (N_107,In_460,In_347);
nand U108 (N_108,In_341,In_220);
and U109 (N_109,In_131,In_297);
or U110 (N_110,In_41,In_232);
and U111 (N_111,In_217,In_112);
nand U112 (N_112,In_138,In_346);
nor U113 (N_113,In_57,In_300);
and U114 (N_114,In_241,In_84);
and U115 (N_115,In_0,In_252);
nand U116 (N_116,In_262,In_499);
nor U117 (N_117,In_102,In_126);
and U118 (N_118,N_98,N_63);
or U119 (N_119,In_4,N_66);
nand U120 (N_120,In_238,In_278);
or U121 (N_121,In_465,In_397);
and U122 (N_122,N_56,In_75);
nor U123 (N_123,N_27,In_161);
or U124 (N_124,In_274,N_47);
nand U125 (N_125,In_332,N_6);
nor U126 (N_126,N_38,N_71);
or U127 (N_127,In_424,N_72);
nand U128 (N_128,In_62,In_287);
and U129 (N_129,In_339,In_358);
and U130 (N_130,In_246,N_24);
nor U131 (N_131,In_459,In_462);
nand U132 (N_132,In_19,In_409);
nor U133 (N_133,N_90,In_155);
nor U134 (N_134,In_420,In_257);
nand U135 (N_135,N_37,In_1);
or U136 (N_136,In_414,N_20);
and U137 (N_137,In_66,In_324);
nand U138 (N_138,N_52,In_73);
nor U139 (N_139,In_248,N_53);
and U140 (N_140,N_42,In_168);
nand U141 (N_141,In_470,N_83);
nand U142 (N_142,In_214,N_95);
or U143 (N_143,In_495,In_10);
or U144 (N_144,N_26,In_201);
nand U145 (N_145,In_189,N_51);
and U146 (N_146,N_81,N_13);
nand U147 (N_147,In_303,In_388);
or U148 (N_148,In_352,In_308);
nand U149 (N_149,N_67,In_198);
nor U150 (N_150,In_9,N_17);
and U151 (N_151,In_194,In_174);
or U152 (N_152,In_133,In_355);
or U153 (N_153,N_50,N_133);
nand U154 (N_154,N_128,N_22);
nand U155 (N_155,N_44,In_82);
nand U156 (N_156,In_395,N_64);
and U157 (N_157,N_57,N_59);
nand U158 (N_158,N_58,In_31);
nand U159 (N_159,N_110,In_29);
and U160 (N_160,In_27,N_11);
xnor U161 (N_161,In_180,N_139);
nor U162 (N_162,In_159,N_35);
nor U163 (N_163,In_392,N_40);
nand U164 (N_164,In_125,In_464);
or U165 (N_165,In_416,In_72);
or U166 (N_166,N_131,In_211);
and U167 (N_167,In_485,N_104);
nand U168 (N_168,In_183,N_136);
or U169 (N_169,In_367,N_122);
nand U170 (N_170,N_75,N_68);
nand U171 (N_171,In_311,N_84);
or U172 (N_172,In_48,N_74);
nor U173 (N_173,In_455,N_134);
and U174 (N_174,In_54,In_279);
and U175 (N_175,In_233,In_307);
nor U176 (N_176,In_94,N_130);
and U177 (N_177,In_249,N_60);
and U178 (N_178,N_93,N_39);
nor U179 (N_179,N_146,N_119);
nor U180 (N_180,In_283,In_291);
or U181 (N_181,In_266,In_160);
nand U182 (N_182,In_13,In_253);
nand U183 (N_183,In_410,In_101);
nor U184 (N_184,In_486,In_114);
or U185 (N_185,In_473,In_222);
or U186 (N_186,In_70,In_400);
nand U187 (N_187,In_116,In_196);
or U188 (N_188,N_114,In_299);
or U189 (N_189,N_28,In_447);
nor U190 (N_190,N_124,N_132);
nand U191 (N_191,In_359,N_121);
and U192 (N_192,In_439,N_142);
nor U193 (N_193,In_292,In_5);
and U194 (N_194,N_120,In_130);
nand U195 (N_195,In_377,In_467);
nor U196 (N_196,N_101,In_24);
nor U197 (N_197,N_143,In_452);
and U198 (N_198,N_96,In_289);
nor U199 (N_199,In_16,In_334);
and U200 (N_200,In_197,In_364);
and U201 (N_201,In_208,N_70);
nor U202 (N_202,N_193,N_55);
and U203 (N_203,In_280,N_105);
or U204 (N_204,N_155,In_370);
nor U205 (N_205,N_3,In_207);
or U206 (N_206,In_374,N_168);
nand U207 (N_207,In_309,N_99);
and U208 (N_208,N_18,N_144);
nand U209 (N_209,In_325,In_403);
and U210 (N_210,In_23,N_129);
and U211 (N_211,In_333,N_135);
or U212 (N_212,N_103,In_335);
or U213 (N_213,In_497,In_421);
nand U214 (N_214,In_56,In_22);
nor U215 (N_215,In_37,N_86);
nor U216 (N_216,N_76,In_30);
and U217 (N_217,In_117,In_272);
and U218 (N_218,N_171,N_150);
or U219 (N_219,N_152,N_1);
or U220 (N_220,In_484,N_140);
and U221 (N_221,In_496,In_165);
nor U222 (N_222,In_202,N_69);
or U223 (N_223,In_79,In_340);
nand U224 (N_224,In_396,In_312);
nand U225 (N_225,In_375,N_156);
and U226 (N_226,N_141,In_310);
nand U227 (N_227,In_99,N_157);
nor U228 (N_228,N_117,In_261);
nor U229 (N_229,In_490,In_78);
and U230 (N_230,N_160,In_229);
nand U231 (N_231,In_223,In_276);
or U232 (N_232,N_147,In_285);
or U233 (N_233,N_137,N_148);
and U234 (N_234,N_34,N_16);
or U235 (N_235,In_65,N_159);
and U236 (N_236,In_46,N_170);
nand U237 (N_237,N_153,In_383);
nor U238 (N_238,N_196,In_154);
or U239 (N_239,N_194,N_192);
or U240 (N_240,In_475,In_213);
nor U241 (N_241,In_251,In_240);
nand U242 (N_242,In_218,N_107);
nor U243 (N_243,N_174,In_487);
nor U244 (N_244,N_108,In_437);
and U245 (N_245,In_381,N_125);
nor U246 (N_246,N_25,In_166);
nand U247 (N_247,N_43,In_100);
or U248 (N_248,In_192,In_275);
or U249 (N_249,In_164,In_6);
nor U250 (N_250,N_239,N_5);
nor U251 (N_251,N_176,N_166);
and U252 (N_252,In_449,In_190);
nor U253 (N_253,N_91,In_373);
and U254 (N_254,In_284,In_378);
nand U255 (N_255,In_144,In_343);
or U256 (N_256,N_45,In_96);
or U257 (N_257,N_199,N_138);
or U258 (N_258,N_187,N_242);
and U259 (N_259,In_448,N_115);
nand U260 (N_260,N_46,In_336);
nand U261 (N_261,N_220,N_211);
nor U262 (N_262,In_36,N_94);
nor U263 (N_263,N_201,In_88);
nor U264 (N_264,In_404,In_350);
nor U265 (N_265,N_188,N_145);
and U266 (N_266,In_463,In_365);
and U267 (N_267,In_461,In_151);
and U268 (N_268,N_237,N_197);
xor U269 (N_269,N_233,N_212);
nor U270 (N_270,N_116,N_169);
nor U271 (N_271,N_218,N_14);
nand U272 (N_272,In_175,N_113);
or U273 (N_273,N_221,N_163);
nand U274 (N_274,In_69,N_246);
nand U275 (N_275,N_207,N_21);
or U276 (N_276,N_161,In_121);
or U277 (N_277,In_105,N_216);
nor U278 (N_278,N_189,N_48);
nor U279 (N_279,N_9,N_185);
nor U280 (N_280,In_204,In_422);
nor U281 (N_281,N_202,In_293);
nor U282 (N_282,N_245,N_92);
or U283 (N_283,N_182,In_466);
xor U284 (N_284,N_173,N_151);
or U285 (N_285,N_181,In_399);
nand U286 (N_286,In_408,N_204);
and U287 (N_287,N_200,N_12);
and U288 (N_288,N_230,In_376);
nand U289 (N_289,In_52,N_248);
nand U290 (N_290,N_183,N_82);
or U291 (N_291,In_433,In_45);
or U292 (N_292,In_361,In_385);
nand U293 (N_293,N_54,In_478);
and U294 (N_294,N_89,N_111);
nand U295 (N_295,N_78,N_167);
or U296 (N_296,N_36,N_178);
or U297 (N_297,In_368,N_203);
nor U298 (N_298,In_454,N_234);
and U299 (N_299,N_77,N_240);
or U300 (N_300,In_191,N_206);
nor U301 (N_301,In_268,N_263);
nor U302 (N_302,N_205,In_135);
nand U303 (N_303,In_479,N_243);
nor U304 (N_304,In_474,N_294);
xnor U305 (N_305,N_123,N_224);
nand U306 (N_306,N_165,N_232);
nor U307 (N_307,N_299,N_231);
or U308 (N_308,N_223,N_162);
nand U309 (N_309,N_257,N_158);
or U310 (N_310,N_102,N_61);
or U311 (N_311,N_228,In_413);
nor U312 (N_312,N_215,N_154);
nor U313 (N_313,N_184,N_270);
or U314 (N_314,N_254,In_483);
nand U315 (N_315,In_337,N_250);
nor U316 (N_316,N_2,N_247);
xor U317 (N_317,In_17,In_235);
nand U318 (N_318,N_29,In_225);
and U319 (N_319,N_112,In_146);
or U320 (N_320,N_274,In_118);
and U321 (N_321,In_47,N_244);
nand U322 (N_322,In_20,N_87);
or U323 (N_323,N_219,N_269);
nor U324 (N_324,N_296,In_398);
nor U325 (N_325,N_177,N_268);
nand U326 (N_326,N_41,N_172);
nand U327 (N_327,In_480,In_260);
xor U328 (N_328,In_305,In_417);
and U329 (N_329,N_73,N_23);
nand U330 (N_330,In_255,In_369);
nor U331 (N_331,N_229,N_287);
nor U332 (N_332,In_95,N_8);
nor U333 (N_333,In_436,N_285);
or U334 (N_334,In_270,N_271);
and U335 (N_335,N_295,In_59);
nand U336 (N_336,N_265,N_175);
and U337 (N_337,N_118,N_259);
or U338 (N_338,N_255,N_191);
nand U339 (N_339,In_498,In_140);
nor U340 (N_340,N_279,N_179);
and U341 (N_341,In_49,N_266);
nor U342 (N_342,In_86,In_441);
or U343 (N_343,N_258,In_468);
nand U344 (N_344,N_238,In_319);
nor U345 (N_345,In_446,In_443);
nand U346 (N_346,In_53,N_214);
nand U347 (N_347,N_208,In_64);
and U348 (N_348,In_290,N_19);
nand U349 (N_349,N_62,N_80);
and U350 (N_350,N_278,In_442);
and U351 (N_351,In_212,N_251);
and U352 (N_352,N_323,N_317);
and U353 (N_353,In_134,N_304);
and U354 (N_354,N_276,N_126);
nand U355 (N_355,N_0,In_471);
nand U356 (N_356,N_267,N_32);
nand U357 (N_357,N_327,N_65);
and U358 (N_358,N_332,N_325);
and U359 (N_359,N_322,N_180);
nand U360 (N_360,N_333,N_195);
or U361 (N_361,N_253,N_292);
or U362 (N_362,N_260,N_273);
or U363 (N_363,N_227,N_340);
xor U364 (N_364,In_25,In_92);
nor U365 (N_365,N_249,N_337);
nand U366 (N_366,N_198,In_32);
or U367 (N_367,N_213,N_275);
and U368 (N_368,N_336,N_302);
or U369 (N_369,N_261,N_288);
nor U370 (N_370,In_477,In_124);
nand U371 (N_371,N_298,N_225);
and U372 (N_372,N_226,N_344);
and U373 (N_373,In_476,N_109);
nand U374 (N_374,N_286,N_303);
nor U375 (N_375,N_300,N_186);
xor U376 (N_376,N_349,N_330);
nor U377 (N_377,N_346,N_342);
nand U378 (N_378,N_282,N_328);
nor U379 (N_379,N_217,In_63);
or U380 (N_380,N_326,N_209);
or U381 (N_381,In_28,In_415);
nand U382 (N_382,N_320,In_51);
and U383 (N_383,N_301,N_293);
nor U384 (N_384,In_85,N_100);
xnor U385 (N_385,In_258,N_252);
nor U386 (N_386,N_190,N_321);
or U387 (N_387,N_97,N_309);
and U388 (N_388,N_305,N_334);
and U389 (N_389,N_315,N_210);
and U390 (N_390,N_281,N_308);
nand U391 (N_391,In_15,N_280);
nor U392 (N_392,N_262,In_321);
xnor U393 (N_393,N_338,N_283);
or U394 (N_394,N_306,In_230);
or U395 (N_395,N_222,N_127);
nor U396 (N_396,N_345,N_49);
or U397 (N_397,N_311,N_307);
nand U398 (N_398,N_4,N_343);
and U399 (N_399,N_310,In_453);
and U400 (N_400,In_104,N_397);
nor U401 (N_401,N_364,N_149);
nand U402 (N_402,N_367,N_354);
nor U403 (N_403,N_290,N_391);
xor U404 (N_404,N_352,N_351);
or U405 (N_405,N_399,N_291);
and U406 (N_406,N_362,N_393);
nor U407 (N_407,N_387,N_331);
and U408 (N_408,N_374,N_264);
or U409 (N_409,In_67,N_341);
nand U410 (N_410,N_388,N_353);
or U411 (N_411,N_379,N_313);
and U412 (N_412,N_370,In_141);
nand U413 (N_413,N_272,N_372);
and U414 (N_414,In_440,N_335);
nor U415 (N_415,N_381,N_329);
nand U416 (N_416,N_355,In_267);
and U417 (N_417,In_139,In_55);
nor U418 (N_418,N_236,In_3);
or U419 (N_419,N_394,In_406);
and U420 (N_420,N_348,In_322);
and U421 (N_421,In_425,N_389);
and U422 (N_422,N_235,N_360);
or U423 (N_423,N_324,N_384);
or U424 (N_424,N_363,N_316);
and U425 (N_425,N_395,N_256);
nor U426 (N_426,N_350,N_375);
and U427 (N_427,In_331,N_312);
and U428 (N_428,N_289,N_382);
or U429 (N_429,N_385,N_241);
nor U430 (N_430,N_378,In_226);
nor U431 (N_431,N_359,In_301);
and U432 (N_432,N_365,N_356);
nand U433 (N_433,N_383,N_297);
or U434 (N_434,In_491,N_277);
nor U435 (N_435,N_371,N_392);
and U436 (N_436,In_176,N_369);
nand U437 (N_437,N_396,N_386);
nor U438 (N_438,In_242,N_318);
nor U439 (N_439,N_284,In_195);
and U440 (N_440,N_377,N_106);
and U441 (N_441,N_347,N_373);
nand U442 (N_442,N_339,N_366);
and U443 (N_443,N_376,In_328);
nand U444 (N_444,N_398,N_357);
and U445 (N_445,N_361,N_380);
nor U446 (N_446,N_368,N_390);
or U447 (N_447,N_10,N_314);
and U448 (N_448,In_128,N_319);
nor U449 (N_449,N_358,N_164);
or U450 (N_450,N_434,N_447);
nor U451 (N_451,N_441,N_406);
and U452 (N_452,N_420,N_442);
and U453 (N_453,N_431,N_421);
nand U454 (N_454,N_449,N_404);
and U455 (N_455,N_419,N_415);
and U456 (N_456,N_430,N_409);
nor U457 (N_457,N_410,N_444);
or U458 (N_458,N_448,N_424);
nor U459 (N_459,N_416,N_402);
nand U460 (N_460,N_426,N_427);
nand U461 (N_461,N_443,N_412);
nor U462 (N_462,N_432,N_411);
nor U463 (N_463,N_446,N_418);
nand U464 (N_464,N_445,N_438);
nor U465 (N_465,N_429,N_425);
or U466 (N_466,N_407,N_422);
nor U467 (N_467,N_401,N_417);
and U468 (N_468,N_423,N_437);
and U469 (N_469,N_414,N_436);
and U470 (N_470,N_433,N_405);
or U471 (N_471,N_428,N_400);
and U472 (N_472,N_439,N_440);
or U473 (N_473,N_403,N_413);
nor U474 (N_474,N_435,N_408);
nand U475 (N_475,N_444,N_401);
and U476 (N_476,N_434,N_422);
and U477 (N_477,N_404,N_433);
nand U478 (N_478,N_442,N_412);
nor U479 (N_479,N_431,N_427);
or U480 (N_480,N_425,N_416);
or U481 (N_481,N_440,N_408);
nand U482 (N_482,N_404,N_415);
nand U483 (N_483,N_440,N_431);
or U484 (N_484,N_409,N_407);
or U485 (N_485,N_404,N_408);
nand U486 (N_486,N_406,N_419);
nand U487 (N_487,N_434,N_433);
and U488 (N_488,N_433,N_418);
or U489 (N_489,N_428,N_427);
or U490 (N_490,N_414,N_437);
nand U491 (N_491,N_443,N_409);
and U492 (N_492,N_435,N_416);
or U493 (N_493,N_400,N_404);
nand U494 (N_494,N_403,N_416);
nor U495 (N_495,N_422,N_417);
nand U496 (N_496,N_434,N_442);
nor U497 (N_497,N_401,N_410);
and U498 (N_498,N_447,N_412);
and U499 (N_499,N_426,N_415);
nand U500 (N_500,N_455,N_493);
xor U501 (N_501,N_488,N_477);
and U502 (N_502,N_495,N_451);
nor U503 (N_503,N_466,N_474);
and U504 (N_504,N_464,N_473);
or U505 (N_505,N_478,N_468);
xor U506 (N_506,N_491,N_484);
or U507 (N_507,N_499,N_457);
nor U508 (N_508,N_454,N_460);
and U509 (N_509,N_475,N_487);
nand U510 (N_510,N_492,N_485);
or U511 (N_511,N_496,N_472);
or U512 (N_512,N_489,N_458);
nand U513 (N_513,N_450,N_453);
nor U514 (N_514,N_459,N_498);
nor U515 (N_515,N_463,N_462);
nor U516 (N_516,N_456,N_480);
and U517 (N_517,N_452,N_481);
nand U518 (N_518,N_476,N_490);
or U519 (N_519,N_471,N_482);
or U520 (N_520,N_470,N_483);
nor U521 (N_521,N_494,N_465);
and U522 (N_522,N_467,N_486);
nand U523 (N_523,N_461,N_469);
nand U524 (N_524,N_479,N_497);
and U525 (N_525,N_473,N_491);
nand U526 (N_526,N_496,N_469);
nand U527 (N_527,N_469,N_492);
nor U528 (N_528,N_495,N_460);
and U529 (N_529,N_467,N_450);
xnor U530 (N_530,N_475,N_473);
or U531 (N_531,N_460,N_486);
and U532 (N_532,N_454,N_484);
nand U533 (N_533,N_455,N_472);
and U534 (N_534,N_479,N_474);
or U535 (N_535,N_457,N_460);
and U536 (N_536,N_467,N_461);
or U537 (N_537,N_486,N_465);
and U538 (N_538,N_499,N_451);
or U539 (N_539,N_465,N_476);
and U540 (N_540,N_453,N_462);
nand U541 (N_541,N_468,N_463);
nand U542 (N_542,N_451,N_484);
and U543 (N_543,N_475,N_497);
nor U544 (N_544,N_466,N_463);
or U545 (N_545,N_470,N_494);
or U546 (N_546,N_475,N_491);
nor U547 (N_547,N_455,N_470);
nand U548 (N_548,N_497,N_487);
or U549 (N_549,N_468,N_467);
nand U550 (N_550,N_517,N_530);
and U551 (N_551,N_509,N_533);
nand U552 (N_552,N_532,N_513);
or U553 (N_553,N_541,N_529);
or U554 (N_554,N_524,N_501);
nor U555 (N_555,N_512,N_516);
or U556 (N_556,N_522,N_508);
and U557 (N_557,N_506,N_520);
or U558 (N_558,N_500,N_518);
nand U559 (N_559,N_503,N_538);
nand U560 (N_560,N_528,N_519);
or U561 (N_561,N_526,N_544);
nand U562 (N_562,N_545,N_546);
xnor U563 (N_563,N_539,N_523);
nand U564 (N_564,N_511,N_525);
and U565 (N_565,N_514,N_535);
or U566 (N_566,N_543,N_502);
nand U567 (N_567,N_548,N_537);
or U568 (N_568,N_540,N_505);
or U569 (N_569,N_547,N_531);
and U570 (N_570,N_534,N_549);
nand U571 (N_571,N_542,N_510);
nor U572 (N_572,N_507,N_504);
nor U573 (N_573,N_536,N_515);
or U574 (N_574,N_521,N_527);
nand U575 (N_575,N_545,N_504);
and U576 (N_576,N_543,N_523);
nor U577 (N_577,N_504,N_508);
and U578 (N_578,N_518,N_540);
nand U579 (N_579,N_505,N_535);
nand U580 (N_580,N_501,N_531);
nor U581 (N_581,N_541,N_527);
nor U582 (N_582,N_512,N_531);
and U583 (N_583,N_515,N_527);
nand U584 (N_584,N_525,N_500);
or U585 (N_585,N_540,N_519);
nand U586 (N_586,N_506,N_521);
or U587 (N_587,N_523,N_534);
or U588 (N_588,N_521,N_518);
nor U589 (N_589,N_523,N_546);
xnor U590 (N_590,N_502,N_528);
and U591 (N_591,N_539,N_546);
and U592 (N_592,N_543,N_511);
nand U593 (N_593,N_529,N_540);
nand U594 (N_594,N_524,N_538);
nand U595 (N_595,N_504,N_502);
nand U596 (N_596,N_506,N_522);
xor U597 (N_597,N_522,N_521);
nor U598 (N_598,N_500,N_543);
nor U599 (N_599,N_518,N_511);
nand U600 (N_600,N_562,N_557);
nand U601 (N_601,N_599,N_568);
nand U602 (N_602,N_564,N_559);
nand U603 (N_603,N_582,N_550);
nor U604 (N_604,N_578,N_589);
nor U605 (N_605,N_590,N_591);
nand U606 (N_606,N_558,N_575);
and U607 (N_607,N_581,N_565);
and U608 (N_608,N_585,N_584);
nor U609 (N_609,N_592,N_553);
nor U610 (N_610,N_567,N_569);
and U611 (N_611,N_574,N_560);
or U612 (N_612,N_580,N_587);
or U613 (N_613,N_551,N_576);
and U614 (N_614,N_556,N_552);
or U615 (N_615,N_598,N_566);
or U616 (N_616,N_579,N_554);
or U617 (N_617,N_571,N_596);
nand U618 (N_618,N_573,N_561);
and U619 (N_619,N_563,N_583);
nor U620 (N_620,N_593,N_594);
or U621 (N_621,N_588,N_555);
nand U622 (N_622,N_597,N_572);
nor U623 (N_623,N_570,N_577);
nor U624 (N_624,N_586,N_595);
nand U625 (N_625,N_597,N_569);
nand U626 (N_626,N_556,N_553);
or U627 (N_627,N_593,N_582);
or U628 (N_628,N_589,N_593);
nand U629 (N_629,N_586,N_592);
or U630 (N_630,N_577,N_590);
nand U631 (N_631,N_594,N_554);
or U632 (N_632,N_577,N_586);
nand U633 (N_633,N_553,N_577);
nor U634 (N_634,N_554,N_591);
nand U635 (N_635,N_552,N_571);
and U636 (N_636,N_590,N_596);
or U637 (N_637,N_591,N_571);
and U638 (N_638,N_598,N_557);
and U639 (N_639,N_569,N_591);
and U640 (N_640,N_562,N_597);
or U641 (N_641,N_578,N_599);
nor U642 (N_642,N_555,N_589);
nand U643 (N_643,N_572,N_568);
nand U644 (N_644,N_572,N_589);
and U645 (N_645,N_554,N_550);
and U646 (N_646,N_561,N_592);
and U647 (N_647,N_563,N_580);
or U648 (N_648,N_599,N_555);
or U649 (N_649,N_575,N_577);
or U650 (N_650,N_646,N_633);
and U651 (N_651,N_610,N_627);
nor U652 (N_652,N_625,N_634);
and U653 (N_653,N_643,N_614);
nor U654 (N_654,N_639,N_631);
nor U655 (N_655,N_611,N_618);
nand U656 (N_656,N_612,N_608);
xor U657 (N_657,N_626,N_617);
nor U658 (N_658,N_605,N_624);
or U659 (N_659,N_616,N_630);
nor U660 (N_660,N_636,N_602);
nor U661 (N_661,N_601,N_613);
and U662 (N_662,N_647,N_603);
or U663 (N_663,N_604,N_649);
or U664 (N_664,N_615,N_620);
and U665 (N_665,N_619,N_648);
nor U666 (N_666,N_621,N_600);
and U667 (N_667,N_607,N_623);
or U668 (N_668,N_628,N_629);
or U669 (N_669,N_609,N_642);
and U670 (N_670,N_645,N_622);
and U671 (N_671,N_641,N_637);
nand U672 (N_672,N_635,N_632);
nand U673 (N_673,N_640,N_644);
nand U674 (N_674,N_638,N_606);
nand U675 (N_675,N_613,N_612);
nor U676 (N_676,N_603,N_616);
nor U677 (N_677,N_622,N_647);
nand U678 (N_678,N_634,N_638);
and U679 (N_679,N_631,N_633);
nand U680 (N_680,N_605,N_644);
or U681 (N_681,N_627,N_639);
and U682 (N_682,N_647,N_602);
and U683 (N_683,N_600,N_646);
and U684 (N_684,N_614,N_605);
nand U685 (N_685,N_614,N_634);
nand U686 (N_686,N_634,N_605);
nor U687 (N_687,N_630,N_643);
and U688 (N_688,N_648,N_600);
nor U689 (N_689,N_619,N_634);
or U690 (N_690,N_644,N_607);
and U691 (N_691,N_603,N_624);
and U692 (N_692,N_620,N_641);
and U693 (N_693,N_621,N_608);
nor U694 (N_694,N_649,N_629);
and U695 (N_695,N_632,N_627);
or U696 (N_696,N_605,N_648);
or U697 (N_697,N_625,N_610);
and U698 (N_698,N_600,N_608);
nand U699 (N_699,N_642,N_633);
nor U700 (N_700,N_688,N_654);
nor U701 (N_701,N_680,N_667);
or U702 (N_702,N_674,N_655);
or U703 (N_703,N_692,N_691);
xor U704 (N_704,N_676,N_698);
nor U705 (N_705,N_687,N_675);
nand U706 (N_706,N_660,N_685);
nand U707 (N_707,N_677,N_694);
or U708 (N_708,N_669,N_662);
nand U709 (N_709,N_699,N_650);
or U710 (N_710,N_697,N_681);
and U711 (N_711,N_672,N_689);
or U712 (N_712,N_656,N_683);
or U713 (N_713,N_658,N_666);
nor U714 (N_714,N_679,N_671);
and U715 (N_715,N_690,N_652);
nor U716 (N_716,N_695,N_673);
nor U717 (N_717,N_684,N_657);
nor U718 (N_718,N_663,N_682);
xor U719 (N_719,N_686,N_693);
nor U720 (N_720,N_678,N_661);
nor U721 (N_721,N_670,N_665);
and U722 (N_722,N_653,N_664);
nand U723 (N_723,N_696,N_659);
or U724 (N_724,N_668,N_651);
nand U725 (N_725,N_650,N_678);
nand U726 (N_726,N_675,N_654);
xor U727 (N_727,N_692,N_664);
or U728 (N_728,N_691,N_688);
nor U729 (N_729,N_678,N_674);
or U730 (N_730,N_692,N_662);
nand U731 (N_731,N_668,N_670);
nor U732 (N_732,N_653,N_679);
nor U733 (N_733,N_671,N_689);
nor U734 (N_734,N_664,N_698);
or U735 (N_735,N_696,N_695);
nand U736 (N_736,N_665,N_689);
nor U737 (N_737,N_670,N_674);
nand U738 (N_738,N_668,N_687);
and U739 (N_739,N_668,N_657);
and U740 (N_740,N_684,N_650);
or U741 (N_741,N_677,N_668);
nor U742 (N_742,N_672,N_652);
nand U743 (N_743,N_656,N_695);
and U744 (N_744,N_663,N_671);
nand U745 (N_745,N_654,N_694);
nor U746 (N_746,N_682,N_697);
nand U747 (N_747,N_652,N_698);
or U748 (N_748,N_653,N_699);
nand U749 (N_749,N_670,N_650);
xnor U750 (N_750,N_704,N_740);
nor U751 (N_751,N_712,N_747);
or U752 (N_752,N_705,N_703);
and U753 (N_753,N_729,N_744);
or U754 (N_754,N_718,N_745);
nor U755 (N_755,N_702,N_713);
nor U756 (N_756,N_730,N_707);
or U757 (N_757,N_737,N_726);
nand U758 (N_758,N_722,N_743);
nor U759 (N_759,N_736,N_731);
and U760 (N_760,N_734,N_711);
xor U761 (N_761,N_706,N_710);
nand U762 (N_762,N_742,N_738);
or U763 (N_763,N_727,N_701);
or U764 (N_764,N_733,N_717);
or U765 (N_765,N_716,N_748);
and U766 (N_766,N_739,N_725);
or U767 (N_767,N_709,N_708);
nand U768 (N_768,N_746,N_720);
or U769 (N_769,N_700,N_728);
or U770 (N_770,N_719,N_723);
nand U771 (N_771,N_735,N_724);
nand U772 (N_772,N_732,N_714);
nor U773 (N_773,N_749,N_715);
nor U774 (N_774,N_721,N_741);
nor U775 (N_775,N_714,N_747);
nor U776 (N_776,N_725,N_738);
and U777 (N_777,N_731,N_748);
and U778 (N_778,N_703,N_748);
or U779 (N_779,N_728,N_711);
and U780 (N_780,N_730,N_704);
and U781 (N_781,N_745,N_727);
nor U782 (N_782,N_727,N_707);
or U783 (N_783,N_728,N_722);
nor U784 (N_784,N_726,N_721);
or U785 (N_785,N_749,N_709);
nor U786 (N_786,N_710,N_747);
nand U787 (N_787,N_710,N_722);
or U788 (N_788,N_726,N_708);
nand U789 (N_789,N_731,N_704);
and U790 (N_790,N_739,N_722);
or U791 (N_791,N_722,N_737);
nand U792 (N_792,N_745,N_723);
and U793 (N_793,N_716,N_701);
or U794 (N_794,N_716,N_724);
or U795 (N_795,N_709,N_711);
nor U796 (N_796,N_745,N_703);
and U797 (N_797,N_733,N_740);
or U798 (N_798,N_735,N_737);
nand U799 (N_799,N_730,N_705);
nand U800 (N_800,N_771,N_764);
nand U801 (N_801,N_787,N_753);
nand U802 (N_802,N_794,N_754);
nor U803 (N_803,N_759,N_758);
or U804 (N_804,N_772,N_798);
and U805 (N_805,N_768,N_775);
and U806 (N_806,N_790,N_767);
nor U807 (N_807,N_799,N_792);
and U808 (N_808,N_756,N_762);
or U809 (N_809,N_793,N_752);
xnor U810 (N_810,N_755,N_795);
or U811 (N_811,N_789,N_779);
nor U812 (N_812,N_765,N_777);
or U813 (N_813,N_791,N_783);
nor U814 (N_814,N_788,N_778);
and U815 (N_815,N_761,N_774);
nor U816 (N_816,N_763,N_782);
and U817 (N_817,N_780,N_766);
and U818 (N_818,N_797,N_751);
nand U819 (N_819,N_784,N_750);
nor U820 (N_820,N_781,N_757);
or U821 (N_821,N_769,N_773);
nor U822 (N_822,N_776,N_786);
and U823 (N_823,N_785,N_770);
and U824 (N_824,N_760,N_796);
or U825 (N_825,N_771,N_782);
or U826 (N_826,N_797,N_763);
nor U827 (N_827,N_797,N_772);
and U828 (N_828,N_764,N_793);
nor U829 (N_829,N_779,N_798);
and U830 (N_830,N_778,N_773);
and U831 (N_831,N_750,N_796);
or U832 (N_832,N_759,N_754);
or U833 (N_833,N_751,N_796);
nor U834 (N_834,N_755,N_777);
nor U835 (N_835,N_789,N_753);
nor U836 (N_836,N_752,N_782);
or U837 (N_837,N_774,N_773);
nor U838 (N_838,N_780,N_755);
and U839 (N_839,N_784,N_796);
or U840 (N_840,N_779,N_795);
and U841 (N_841,N_761,N_763);
nand U842 (N_842,N_760,N_781);
nor U843 (N_843,N_786,N_787);
nor U844 (N_844,N_759,N_771);
or U845 (N_845,N_754,N_783);
and U846 (N_846,N_797,N_774);
nand U847 (N_847,N_779,N_796);
or U848 (N_848,N_779,N_775);
or U849 (N_849,N_761,N_789);
nor U850 (N_850,N_832,N_821);
or U851 (N_851,N_834,N_815);
nor U852 (N_852,N_800,N_819);
nor U853 (N_853,N_838,N_812);
nor U854 (N_854,N_816,N_817);
and U855 (N_855,N_839,N_846);
nand U856 (N_856,N_833,N_849);
nand U857 (N_857,N_810,N_814);
and U858 (N_858,N_802,N_808);
nand U859 (N_859,N_811,N_809);
nor U860 (N_860,N_807,N_844);
nor U861 (N_861,N_824,N_836);
and U862 (N_862,N_837,N_827);
and U863 (N_863,N_804,N_803);
and U864 (N_864,N_829,N_823);
and U865 (N_865,N_841,N_805);
or U866 (N_866,N_813,N_845);
and U867 (N_867,N_822,N_840);
nor U868 (N_868,N_848,N_826);
nor U869 (N_869,N_801,N_842);
nand U870 (N_870,N_830,N_843);
nand U871 (N_871,N_820,N_831);
nor U872 (N_872,N_825,N_818);
nor U873 (N_873,N_806,N_835);
or U874 (N_874,N_847,N_828);
or U875 (N_875,N_849,N_828);
nand U876 (N_876,N_840,N_807);
nand U877 (N_877,N_816,N_846);
and U878 (N_878,N_818,N_820);
nand U879 (N_879,N_834,N_836);
nand U880 (N_880,N_818,N_846);
nor U881 (N_881,N_836,N_809);
and U882 (N_882,N_818,N_829);
or U883 (N_883,N_814,N_815);
or U884 (N_884,N_814,N_842);
and U885 (N_885,N_823,N_846);
xor U886 (N_886,N_838,N_805);
or U887 (N_887,N_841,N_808);
nor U888 (N_888,N_817,N_840);
and U889 (N_889,N_806,N_823);
xor U890 (N_890,N_835,N_831);
nand U891 (N_891,N_833,N_809);
or U892 (N_892,N_803,N_849);
and U893 (N_893,N_800,N_834);
nand U894 (N_894,N_814,N_837);
nand U895 (N_895,N_815,N_849);
nor U896 (N_896,N_816,N_830);
nor U897 (N_897,N_847,N_808);
nor U898 (N_898,N_849,N_802);
and U899 (N_899,N_846,N_833);
and U900 (N_900,N_888,N_880);
or U901 (N_901,N_851,N_881);
or U902 (N_902,N_865,N_877);
nor U903 (N_903,N_868,N_882);
and U904 (N_904,N_885,N_879);
nand U905 (N_905,N_892,N_864);
nor U906 (N_906,N_890,N_894);
and U907 (N_907,N_862,N_876);
or U908 (N_908,N_857,N_889);
nor U909 (N_909,N_872,N_861);
nor U910 (N_910,N_858,N_863);
or U911 (N_911,N_850,N_883);
and U912 (N_912,N_870,N_855);
and U913 (N_913,N_871,N_869);
or U914 (N_914,N_859,N_867);
nand U915 (N_915,N_874,N_878);
and U916 (N_916,N_899,N_875);
xnor U917 (N_917,N_896,N_895);
and U918 (N_918,N_893,N_886);
nor U919 (N_919,N_873,N_852);
nor U920 (N_920,N_856,N_891);
or U921 (N_921,N_854,N_866);
or U922 (N_922,N_898,N_853);
or U923 (N_923,N_884,N_897);
or U924 (N_924,N_887,N_860);
or U925 (N_925,N_893,N_872);
nor U926 (N_926,N_890,N_860);
xnor U927 (N_927,N_855,N_865);
nor U928 (N_928,N_852,N_882);
nand U929 (N_929,N_857,N_855);
nand U930 (N_930,N_883,N_899);
or U931 (N_931,N_881,N_887);
or U932 (N_932,N_882,N_894);
and U933 (N_933,N_884,N_856);
and U934 (N_934,N_897,N_875);
nand U935 (N_935,N_862,N_866);
nor U936 (N_936,N_885,N_894);
and U937 (N_937,N_876,N_859);
or U938 (N_938,N_858,N_865);
nor U939 (N_939,N_894,N_892);
or U940 (N_940,N_868,N_899);
and U941 (N_941,N_867,N_895);
or U942 (N_942,N_885,N_888);
nor U943 (N_943,N_854,N_879);
nand U944 (N_944,N_874,N_853);
and U945 (N_945,N_892,N_862);
or U946 (N_946,N_885,N_858);
nor U947 (N_947,N_869,N_853);
or U948 (N_948,N_867,N_871);
nand U949 (N_949,N_890,N_861);
nand U950 (N_950,N_919,N_948);
nor U951 (N_951,N_938,N_939);
and U952 (N_952,N_932,N_946);
nand U953 (N_953,N_944,N_906);
or U954 (N_954,N_901,N_918);
and U955 (N_955,N_937,N_942);
nor U956 (N_956,N_949,N_912);
nor U957 (N_957,N_945,N_902);
nand U958 (N_958,N_921,N_947);
and U959 (N_959,N_935,N_941);
xnor U960 (N_960,N_924,N_940);
and U961 (N_961,N_927,N_928);
and U962 (N_962,N_903,N_920);
or U963 (N_963,N_915,N_922);
nand U964 (N_964,N_943,N_909);
nor U965 (N_965,N_900,N_931);
or U966 (N_966,N_905,N_911);
nor U967 (N_967,N_908,N_929);
or U968 (N_968,N_930,N_925);
nand U969 (N_969,N_913,N_936);
nand U970 (N_970,N_934,N_933);
nand U971 (N_971,N_926,N_904);
or U972 (N_972,N_917,N_910);
nand U973 (N_973,N_923,N_907);
nand U974 (N_974,N_914,N_916);
and U975 (N_975,N_925,N_948);
and U976 (N_976,N_923,N_938);
and U977 (N_977,N_902,N_935);
and U978 (N_978,N_900,N_908);
or U979 (N_979,N_907,N_912);
nor U980 (N_980,N_918,N_919);
nand U981 (N_981,N_924,N_907);
or U982 (N_982,N_927,N_913);
xor U983 (N_983,N_908,N_949);
and U984 (N_984,N_933,N_923);
nand U985 (N_985,N_938,N_943);
and U986 (N_986,N_947,N_941);
and U987 (N_987,N_904,N_948);
nand U988 (N_988,N_946,N_949);
nand U989 (N_989,N_937,N_904);
nand U990 (N_990,N_932,N_919);
and U991 (N_991,N_940,N_930);
nor U992 (N_992,N_912,N_947);
or U993 (N_993,N_917,N_934);
and U994 (N_994,N_943,N_929);
and U995 (N_995,N_944,N_909);
nand U996 (N_996,N_944,N_934);
nor U997 (N_997,N_920,N_947);
or U998 (N_998,N_913,N_924);
xnor U999 (N_999,N_908,N_935);
nor U1000 (N_1000,N_957,N_962);
nor U1001 (N_1001,N_993,N_998);
and U1002 (N_1002,N_958,N_968);
nand U1003 (N_1003,N_986,N_991);
nand U1004 (N_1004,N_996,N_965);
nand U1005 (N_1005,N_997,N_956);
or U1006 (N_1006,N_951,N_999);
nand U1007 (N_1007,N_961,N_995);
or U1008 (N_1008,N_981,N_953);
nor U1009 (N_1009,N_960,N_972);
and U1010 (N_1010,N_989,N_971);
nand U1011 (N_1011,N_967,N_973);
nand U1012 (N_1012,N_954,N_950);
nand U1013 (N_1013,N_987,N_988);
and U1014 (N_1014,N_979,N_966);
or U1015 (N_1015,N_970,N_983);
nand U1016 (N_1016,N_980,N_994);
nor U1017 (N_1017,N_955,N_984);
and U1018 (N_1018,N_992,N_975);
nand U1019 (N_1019,N_963,N_964);
nand U1020 (N_1020,N_985,N_977);
nor U1021 (N_1021,N_982,N_974);
or U1022 (N_1022,N_990,N_976);
nand U1023 (N_1023,N_978,N_959);
nor U1024 (N_1024,N_969,N_952);
or U1025 (N_1025,N_988,N_983);
xor U1026 (N_1026,N_963,N_951);
nor U1027 (N_1027,N_954,N_957);
nand U1028 (N_1028,N_950,N_960);
nor U1029 (N_1029,N_984,N_983);
or U1030 (N_1030,N_987,N_999);
or U1031 (N_1031,N_967,N_958);
nand U1032 (N_1032,N_965,N_983);
nand U1033 (N_1033,N_955,N_969);
or U1034 (N_1034,N_959,N_968);
nor U1035 (N_1035,N_952,N_995);
nor U1036 (N_1036,N_963,N_972);
or U1037 (N_1037,N_958,N_971);
and U1038 (N_1038,N_952,N_954);
or U1039 (N_1039,N_972,N_971);
or U1040 (N_1040,N_964,N_973);
or U1041 (N_1041,N_983,N_976);
nand U1042 (N_1042,N_963,N_953);
nand U1043 (N_1043,N_963,N_976);
or U1044 (N_1044,N_977,N_993);
nor U1045 (N_1045,N_998,N_980);
nor U1046 (N_1046,N_950,N_973);
and U1047 (N_1047,N_985,N_986);
and U1048 (N_1048,N_995,N_959);
nor U1049 (N_1049,N_998,N_978);
and U1050 (N_1050,N_1027,N_1006);
nor U1051 (N_1051,N_1014,N_1046);
nor U1052 (N_1052,N_1007,N_1047);
nor U1053 (N_1053,N_1035,N_1033);
or U1054 (N_1054,N_1019,N_1036);
nor U1055 (N_1055,N_1045,N_1043);
or U1056 (N_1056,N_1012,N_1013);
nor U1057 (N_1057,N_1042,N_1049);
nand U1058 (N_1058,N_1044,N_1032);
and U1059 (N_1059,N_1030,N_1018);
and U1060 (N_1060,N_1040,N_1016);
or U1061 (N_1061,N_1028,N_1010);
nor U1062 (N_1062,N_1029,N_1039);
and U1063 (N_1063,N_1000,N_1020);
nor U1064 (N_1064,N_1034,N_1023);
or U1065 (N_1065,N_1038,N_1015);
or U1066 (N_1066,N_1048,N_1025);
or U1067 (N_1067,N_1005,N_1037);
nor U1068 (N_1068,N_1026,N_1004);
nand U1069 (N_1069,N_1001,N_1002);
and U1070 (N_1070,N_1031,N_1021);
nor U1071 (N_1071,N_1003,N_1009);
nor U1072 (N_1072,N_1022,N_1017);
nor U1073 (N_1073,N_1024,N_1041);
nand U1074 (N_1074,N_1011,N_1008);
nand U1075 (N_1075,N_1008,N_1049);
nand U1076 (N_1076,N_1029,N_1022);
nor U1077 (N_1077,N_1048,N_1028);
and U1078 (N_1078,N_1011,N_1026);
or U1079 (N_1079,N_1010,N_1042);
nand U1080 (N_1080,N_1040,N_1000);
and U1081 (N_1081,N_1010,N_1049);
and U1082 (N_1082,N_1048,N_1023);
nand U1083 (N_1083,N_1040,N_1018);
and U1084 (N_1084,N_1013,N_1041);
or U1085 (N_1085,N_1019,N_1000);
nand U1086 (N_1086,N_1040,N_1043);
nand U1087 (N_1087,N_1034,N_1001);
nand U1088 (N_1088,N_1038,N_1037);
nor U1089 (N_1089,N_1007,N_1001);
xor U1090 (N_1090,N_1014,N_1038);
or U1091 (N_1091,N_1032,N_1038);
and U1092 (N_1092,N_1039,N_1016);
and U1093 (N_1093,N_1019,N_1045);
and U1094 (N_1094,N_1041,N_1029);
and U1095 (N_1095,N_1030,N_1040);
nor U1096 (N_1096,N_1025,N_1002);
nor U1097 (N_1097,N_1009,N_1004);
nand U1098 (N_1098,N_1008,N_1002);
and U1099 (N_1099,N_1008,N_1003);
or U1100 (N_1100,N_1088,N_1054);
nor U1101 (N_1101,N_1082,N_1081);
nor U1102 (N_1102,N_1069,N_1061);
or U1103 (N_1103,N_1072,N_1083);
nor U1104 (N_1104,N_1080,N_1076);
and U1105 (N_1105,N_1055,N_1098);
nand U1106 (N_1106,N_1089,N_1091);
or U1107 (N_1107,N_1085,N_1090);
nor U1108 (N_1108,N_1092,N_1093);
nor U1109 (N_1109,N_1096,N_1095);
nand U1110 (N_1110,N_1063,N_1079);
nor U1111 (N_1111,N_1075,N_1077);
nand U1112 (N_1112,N_1099,N_1062);
nand U1113 (N_1113,N_1087,N_1073);
or U1114 (N_1114,N_1052,N_1071);
or U1115 (N_1115,N_1084,N_1074);
or U1116 (N_1116,N_1057,N_1097);
nor U1117 (N_1117,N_1056,N_1051);
nand U1118 (N_1118,N_1060,N_1086);
nor U1119 (N_1119,N_1050,N_1094);
nor U1120 (N_1120,N_1064,N_1059);
nand U1121 (N_1121,N_1068,N_1067);
and U1122 (N_1122,N_1065,N_1066);
nand U1123 (N_1123,N_1053,N_1078);
or U1124 (N_1124,N_1058,N_1070);
and U1125 (N_1125,N_1071,N_1061);
and U1126 (N_1126,N_1056,N_1099);
or U1127 (N_1127,N_1064,N_1085);
and U1128 (N_1128,N_1096,N_1097);
nor U1129 (N_1129,N_1083,N_1051);
or U1130 (N_1130,N_1068,N_1087);
or U1131 (N_1131,N_1082,N_1070);
and U1132 (N_1132,N_1058,N_1085);
or U1133 (N_1133,N_1050,N_1051);
or U1134 (N_1134,N_1077,N_1052);
nor U1135 (N_1135,N_1050,N_1080);
nor U1136 (N_1136,N_1069,N_1085);
or U1137 (N_1137,N_1073,N_1053);
or U1138 (N_1138,N_1097,N_1076);
and U1139 (N_1139,N_1085,N_1056);
or U1140 (N_1140,N_1087,N_1061);
or U1141 (N_1141,N_1098,N_1069);
or U1142 (N_1142,N_1095,N_1054);
or U1143 (N_1143,N_1084,N_1080);
nor U1144 (N_1144,N_1064,N_1061);
or U1145 (N_1145,N_1098,N_1079);
and U1146 (N_1146,N_1071,N_1051);
and U1147 (N_1147,N_1090,N_1084);
and U1148 (N_1148,N_1061,N_1053);
or U1149 (N_1149,N_1097,N_1075);
nor U1150 (N_1150,N_1122,N_1119);
nor U1151 (N_1151,N_1112,N_1113);
and U1152 (N_1152,N_1148,N_1107);
or U1153 (N_1153,N_1108,N_1149);
or U1154 (N_1154,N_1106,N_1104);
xor U1155 (N_1155,N_1134,N_1147);
or U1156 (N_1156,N_1111,N_1141);
nand U1157 (N_1157,N_1133,N_1144);
nand U1158 (N_1158,N_1136,N_1138);
and U1159 (N_1159,N_1130,N_1115);
nor U1160 (N_1160,N_1121,N_1123);
and U1161 (N_1161,N_1110,N_1135);
or U1162 (N_1162,N_1145,N_1125);
nand U1163 (N_1163,N_1100,N_1127);
nor U1164 (N_1164,N_1140,N_1146);
nand U1165 (N_1165,N_1102,N_1116);
and U1166 (N_1166,N_1114,N_1131);
nand U1167 (N_1167,N_1128,N_1101);
nor U1168 (N_1168,N_1105,N_1142);
and U1169 (N_1169,N_1139,N_1132);
nor U1170 (N_1170,N_1129,N_1103);
or U1171 (N_1171,N_1137,N_1124);
nand U1172 (N_1172,N_1117,N_1109);
or U1173 (N_1173,N_1126,N_1118);
nor U1174 (N_1174,N_1143,N_1120);
nand U1175 (N_1175,N_1122,N_1100);
nand U1176 (N_1176,N_1126,N_1117);
and U1177 (N_1177,N_1106,N_1103);
or U1178 (N_1178,N_1149,N_1145);
and U1179 (N_1179,N_1109,N_1133);
nand U1180 (N_1180,N_1149,N_1139);
or U1181 (N_1181,N_1142,N_1139);
or U1182 (N_1182,N_1133,N_1146);
nor U1183 (N_1183,N_1106,N_1134);
and U1184 (N_1184,N_1124,N_1138);
nor U1185 (N_1185,N_1133,N_1129);
and U1186 (N_1186,N_1126,N_1108);
and U1187 (N_1187,N_1119,N_1111);
nor U1188 (N_1188,N_1113,N_1145);
nor U1189 (N_1189,N_1103,N_1119);
nor U1190 (N_1190,N_1104,N_1112);
nand U1191 (N_1191,N_1130,N_1146);
xor U1192 (N_1192,N_1112,N_1101);
or U1193 (N_1193,N_1137,N_1112);
nand U1194 (N_1194,N_1140,N_1117);
xnor U1195 (N_1195,N_1140,N_1105);
nand U1196 (N_1196,N_1100,N_1112);
nand U1197 (N_1197,N_1103,N_1136);
nor U1198 (N_1198,N_1101,N_1130);
nor U1199 (N_1199,N_1110,N_1123);
nor U1200 (N_1200,N_1150,N_1195);
nand U1201 (N_1201,N_1162,N_1156);
nor U1202 (N_1202,N_1193,N_1175);
and U1203 (N_1203,N_1164,N_1171);
and U1204 (N_1204,N_1158,N_1184);
nand U1205 (N_1205,N_1152,N_1157);
nand U1206 (N_1206,N_1154,N_1166);
nand U1207 (N_1207,N_1168,N_1165);
xnor U1208 (N_1208,N_1182,N_1151);
nand U1209 (N_1209,N_1174,N_1181);
and U1210 (N_1210,N_1159,N_1178);
nor U1211 (N_1211,N_1155,N_1194);
nor U1212 (N_1212,N_1187,N_1186);
or U1213 (N_1213,N_1160,N_1173);
nor U1214 (N_1214,N_1172,N_1190);
and U1215 (N_1215,N_1163,N_1179);
xor U1216 (N_1216,N_1197,N_1191);
and U1217 (N_1217,N_1188,N_1196);
and U1218 (N_1218,N_1198,N_1167);
or U1219 (N_1219,N_1170,N_1192);
nor U1220 (N_1220,N_1180,N_1176);
nand U1221 (N_1221,N_1189,N_1183);
or U1222 (N_1222,N_1177,N_1185);
and U1223 (N_1223,N_1169,N_1199);
and U1224 (N_1224,N_1161,N_1153);
or U1225 (N_1225,N_1164,N_1188);
xnor U1226 (N_1226,N_1160,N_1165);
nand U1227 (N_1227,N_1163,N_1193);
and U1228 (N_1228,N_1194,N_1171);
nor U1229 (N_1229,N_1168,N_1154);
nor U1230 (N_1230,N_1185,N_1155);
xor U1231 (N_1231,N_1194,N_1198);
nor U1232 (N_1232,N_1189,N_1191);
nor U1233 (N_1233,N_1160,N_1170);
and U1234 (N_1234,N_1163,N_1172);
and U1235 (N_1235,N_1152,N_1189);
and U1236 (N_1236,N_1163,N_1152);
nor U1237 (N_1237,N_1177,N_1156);
and U1238 (N_1238,N_1189,N_1185);
or U1239 (N_1239,N_1176,N_1160);
nand U1240 (N_1240,N_1185,N_1152);
nand U1241 (N_1241,N_1164,N_1163);
nor U1242 (N_1242,N_1161,N_1174);
nand U1243 (N_1243,N_1180,N_1154);
nor U1244 (N_1244,N_1185,N_1191);
or U1245 (N_1245,N_1178,N_1195);
and U1246 (N_1246,N_1191,N_1167);
nor U1247 (N_1247,N_1183,N_1198);
or U1248 (N_1248,N_1170,N_1163);
nor U1249 (N_1249,N_1173,N_1163);
nor U1250 (N_1250,N_1234,N_1222);
and U1251 (N_1251,N_1241,N_1244);
or U1252 (N_1252,N_1231,N_1245);
or U1253 (N_1253,N_1225,N_1237);
nor U1254 (N_1254,N_1243,N_1219);
nand U1255 (N_1255,N_1235,N_1240);
or U1256 (N_1256,N_1248,N_1223);
nand U1257 (N_1257,N_1249,N_1209);
nor U1258 (N_1258,N_1228,N_1229);
and U1259 (N_1259,N_1238,N_1205);
or U1260 (N_1260,N_1201,N_1210);
or U1261 (N_1261,N_1224,N_1206);
or U1262 (N_1262,N_1246,N_1217);
and U1263 (N_1263,N_1226,N_1242);
and U1264 (N_1264,N_1230,N_1214);
nor U1265 (N_1265,N_1200,N_1215);
or U1266 (N_1266,N_1213,N_1221);
or U1267 (N_1267,N_1212,N_1202);
nand U1268 (N_1268,N_1227,N_1211);
or U1269 (N_1269,N_1208,N_1216);
or U1270 (N_1270,N_1239,N_1203);
nor U1271 (N_1271,N_1220,N_1236);
nand U1272 (N_1272,N_1232,N_1218);
and U1273 (N_1273,N_1207,N_1247);
or U1274 (N_1274,N_1233,N_1204);
nor U1275 (N_1275,N_1220,N_1200);
nor U1276 (N_1276,N_1212,N_1243);
or U1277 (N_1277,N_1225,N_1248);
nor U1278 (N_1278,N_1244,N_1223);
nor U1279 (N_1279,N_1249,N_1223);
or U1280 (N_1280,N_1233,N_1229);
or U1281 (N_1281,N_1230,N_1238);
nand U1282 (N_1282,N_1204,N_1207);
nand U1283 (N_1283,N_1246,N_1203);
or U1284 (N_1284,N_1203,N_1248);
nor U1285 (N_1285,N_1212,N_1213);
or U1286 (N_1286,N_1239,N_1246);
or U1287 (N_1287,N_1225,N_1243);
and U1288 (N_1288,N_1223,N_1202);
and U1289 (N_1289,N_1206,N_1233);
or U1290 (N_1290,N_1207,N_1224);
or U1291 (N_1291,N_1220,N_1248);
nor U1292 (N_1292,N_1237,N_1207);
or U1293 (N_1293,N_1235,N_1245);
and U1294 (N_1294,N_1247,N_1233);
nand U1295 (N_1295,N_1232,N_1245);
or U1296 (N_1296,N_1203,N_1222);
nand U1297 (N_1297,N_1216,N_1210);
nand U1298 (N_1298,N_1203,N_1237);
or U1299 (N_1299,N_1207,N_1200);
or U1300 (N_1300,N_1250,N_1255);
and U1301 (N_1301,N_1256,N_1260);
and U1302 (N_1302,N_1266,N_1258);
nand U1303 (N_1303,N_1295,N_1262);
nand U1304 (N_1304,N_1288,N_1297);
nor U1305 (N_1305,N_1289,N_1292);
or U1306 (N_1306,N_1276,N_1286);
nand U1307 (N_1307,N_1271,N_1280);
nor U1308 (N_1308,N_1299,N_1252);
and U1309 (N_1309,N_1296,N_1283);
and U1310 (N_1310,N_1263,N_1282);
nor U1311 (N_1311,N_1287,N_1264);
nand U1312 (N_1312,N_1270,N_1261);
and U1313 (N_1313,N_1254,N_1267);
or U1314 (N_1314,N_1275,N_1298);
nand U1315 (N_1315,N_1293,N_1294);
nor U1316 (N_1316,N_1268,N_1272);
and U1317 (N_1317,N_1274,N_1277);
or U1318 (N_1318,N_1273,N_1284);
and U1319 (N_1319,N_1265,N_1285);
and U1320 (N_1320,N_1291,N_1259);
nor U1321 (N_1321,N_1278,N_1251);
nand U1322 (N_1322,N_1279,N_1281);
nor U1323 (N_1323,N_1290,N_1257);
nand U1324 (N_1324,N_1253,N_1269);
or U1325 (N_1325,N_1259,N_1268);
and U1326 (N_1326,N_1289,N_1293);
nand U1327 (N_1327,N_1294,N_1257);
and U1328 (N_1328,N_1266,N_1274);
xor U1329 (N_1329,N_1289,N_1287);
and U1330 (N_1330,N_1271,N_1265);
nand U1331 (N_1331,N_1290,N_1264);
nand U1332 (N_1332,N_1275,N_1269);
nand U1333 (N_1333,N_1269,N_1252);
and U1334 (N_1334,N_1296,N_1251);
nand U1335 (N_1335,N_1282,N_1283);
nor U1336 (N_1336,N_1269,N_1284);
nand U1337 (N_1337,N_1295,N_1266);
nor U1338 (N_1338,N_1287,N_1257);
nand U1339 (N_1339,N_1276,N_1278);
and U1340 (N_1340,N_1279,N_1298);
nand U1341 (N_1341,N_1283,N_1257);
and U1342 (N_1342,N_1272,N_1278);
nor U1343 (N_1343,N_1269,N_1288);
and U1344 (N_1344,N_1255,N_1268);
nor U1345 (N_1345,N_1251,N_1289);
and U1346 (N_1346,N_1286,N_1253);
nand U1347 (N_1347,N_1295,N_1257);
xor U1348 (N_1348,N_1269,N_1295);
and U1349 (N_1349,N_1297,N_1296);
and U1350 (N_1350,N_1341,N_1336);
or U1351 (N_1351,N_1307,N_1317);
and U1352 (N_1352,N_1323,N_1318);
nand U1353 (N_1353,N_1308,N_1340);
nand U1354 (N_1354,N_1339,N_1343);
xor U1355 (N_1355,N_1347,N_1344);
nor U1356 (N_1356,N_1345,N_1342);
or U1357 (N_1357,N_1302,N_1335);
and U1358 (N_1358,N_1334,N_1346);
nand U1359 (N_1359,N_1305,N_1300);
or U1360 (N_1360,N_1321,N_1304);
nand U1361 (N_1361,N_1326,N_1301);
or U1362 (N_1362,N_1310,N_1316);
nor U1363 (N_1363,N_1324,N_1331);
and U1364 (N_1364,N_1325,N_1306);
nand U1365 (N_1365,N_1338,N_1320);
nor U1366 (N_1366,N_1332,N_1309);
nor U1367 (N_1367,N_1327,N_1333);
nor U1368 (N_1368,N_1328,N_1337);
nor U1369 (N_1369,N_1303,N_1312);
nor U1370 (N_1370,N_1319,N_1313);
nor U1371 (N_1371,N_1330,N_1348);
or U1372 (N_1372,N_1314,N_1315);
nor U1373 (N_1373,N_1349,N_1322);
nor U1374 (N_1374,N_1311,N_1329);
and U1375 (N_1375,N_1313,N_1323);
nor U1376 (N_1376,N_1334,N_1324);
and U1377 (N_1377,N_1336,N_1311);
nor U1378 (N_1378,N_1300,N_1336);
and U1379 (N_1379,N_1309,N_1329);
or U1380 (N_1380,N_1324,N_1314);
and U1381 (N_1381,N_1333,N_1324);
or U1382 (N_1382,N_1328,N_1318);
xor U1383 (N_1383,N_1330,N_1339);
and U1384 (N_1384,N_1303,N_1327);
nor U1385 (N_1385,N_1304,N_1340);
nand U1386 (N_1386,N_1313,N_1320);
and U1387 (N_1387,N_1336,N_1305);
and U1388 (N_1388,N_1316,N_1337);
nor U1389 (N_1389,N_1329,N_1318);
and U1390 (N_1390,N_1328,N_1316);
and U1391 (N_1391,N_1317,N_1346);
or U1392 (N_1392,N_1311,N_1349);
and U1393 (N_1393,N_1320,N_1343);
nor U1394 (N_1394,N_1328,N_1313);
nor U1395 (N_1395,N_1320,N_1319);
or U1396 (N_1396,N_1319,N_1305);
and U1397 (N_1397,N_1300,N_1328);
or U1398 (N_1398,N_1322,N_1301);
nor U1399 (N_1399,N_1344,N_1336);
nor U1400 (N_1400,N_1378,N_1369);
and U1401 (N_1401,N_1359,N_1350);
nor U1402 (N_1402,N_1391,N_1360);
and U1403 (N_1403,N_1352,N_1393);
or U1404 (N_1404,N_1377,N_1396);
and U1405 (N_1405,N_1384,N_1353);
or U1406 (N_1406,N_1390,N_1372);
nor U1407 (N_1407,N_1398,N_1351);
or U1408 (N_1408,N_1367,N_1376);
and U1409 (N_1409,N_1379,N_1382);
nand U1410 (N_1410,N_1361,N_1399);
nor U1411 (N_1411,N_1392,N_1386);
and U1412 (N_1412,N_1387,N_1381);
or U1413 (N_1413,N_1366,N_1373);
nor U1414 (N_1414,N_1365,N_1395);
nand U1415 (N_1415,N_1380,N_1383);
nand U1416 (N_1416,N_1374,N_1364);
nor U1417 (N_1417,N_1388,N_1363);
or U1418 (N_1418,N_1355,N_1358);
and U1419 (N_1419,N_1371,N_1362);
nor U1420 (N_1420,N_1368,N_1354);
nor U1421 (N_1421,N_1385,N_1370);
and U1422 (N_1422,N_1394,N_1397);
nor U1423 (N_1423,N_1356,N_1389);
nor U1424 (N_1424,N_1375,N_1357);
nor U1425 (N_1425,N_1387,N_1360);
nand U1426 (N_1426,N_1362,N_1388);
nor U1427 (N_1427,N_1394,N_1398);
and U1428 (N_1428,N_1379,N_1386);
and U1429 (N_1429,N_1375,N_1371);
and U1430 (N_1430,N_1355,N_1365);
or U1431 (N_1431,N_1387,N_1374);
or U1432 (N_1432,N_1359,N_1381);
nor U1433 (N_1433,N_1363,N_1355);
or U1434 (N_1434,N_1369,N_1356);
and U1435 (N_1435,N_1354,N_1396);
or U1436 (N_1436,N_1373,N_1392);
or U1437 (N_1437,N_1390,N_1366);
and U1438 (N_1438,N_1375,N_1385);
and U1439 (N_1439,N_1364,N_1361);
nand U1440 (N_1440,N_1351,N_1354);
or U1441 (N_1441,N_1394,N_1362);
and U1442 (N_1442,N_1375,N_1388);
nand U1443 (N_1443,N_1392,N_1355);
nor U1444 (N_1444,N_1381,N_1386);
xnor U1445 (N_1445,N_1387,N_1395);
or U1446 (N_1446,N_1397,N_1361);
or U1447 (N_1447,N_1367,N_1380);
or U1448 (N_1448,N_1395,N_1397);
or U1449 (N_1449,N_1361,N_1389);
nand U1450 (N_1450,N_1425,N_1423);
and U1451 (N_1451,N_1417,N_1428);
or U1452 (N_1452,N_1444,N_1433);
or U1453 (N_1453,N_1411,N_1404);
or U1454 (N_1454,N_1424,N_1419);
and U1455 (N_1455,N_1405,N_1446);
and U1456 (N_1456,N_1418,N_1440);
and U1457 (N_1457,N_1420,N_1410);
nand U1458 (N_1458,N_1426,N_1422);
or U1459 (N_1459,N_1416,N_1438);
or U1460 (N_1460,N_1427,N_1429);
nor U1461 (N_1461,N_1412,N_1435);
nor U1462 (N_1462,N_1415,N_1448);
and U1463 (N_1463,N_1442,N_1413);
and U1464 (N_1464,N_1407,N_1401);
nor U1465 (N_1465,N_1434,N_1445);
or U1466 (N_1466,N_1409,N_1447);
or U1467 (N_1467,N_1408,N_1443);
nor U1468 (N_1468,N_1403,N_1437);
and U1469 (N_1469,N_1432,N_1414);
nand U1470 (N_1470,N_1441,N_1406);
or U1471 (N_1471,N_1436,N_1449);
nand U1472 (N_1472,N_1421,N_1402);
nand U1473 (N_1473,N_1400,N_1431);
nor U1474 (N_1474,N_1439,N_1430);
nand U1475 (N_1475,N_1426,N_1423);
nor U1476 (N_1476,N_1436,N_1402);
nand U1477 (N_1477,N_1437,N_1430);
nor U1478 (N_1478,N_1413,N_1409);
nor U1479 (N_1479,N_1426,N_1438);
nor U1480 (N_1480,N_1408,N_1420);
nand U1481 (N_1481,N_1418,N_1421);
nand U1482 (N_1482,N_1445,N_1429);
or U1483 (N_1483,N_1405,N_1406);
nor U1484 (N_1484,N_1415,N_1431);
or U1485 (N_1485,N_1448,N_1449);
nor U1486 (N_1486,N_1431,N_1435);
or U1487 (N_1487,N_1419,N_1426);
nor U1488 (N_1488,N_1419,N_1434);
nand U1489 (N_1489,N_1439,N_1428);
nor U1490 (N_1490,N_1420,N_1416);
and U1491 (N_1491,N_1418,N_1425);
nand U1492 (N_1492,N_1408,N_1415);
and U1493 (N_1493,N_1401,N_1433);
and U1494 (N_1494,N_1416,N_1421);
nand U1495 (N_1495,N_1417,N_1434);
and U1496 (N_1496,N_1428,N_1423);
and U1497 (N_1497,N_1405,N_1432);
or U1498 (N_1498,N_1429,N_1418);
nor U1499 (N_1499,N_1429,N_1412);
nor U1500 (N_1500,N_1469,N_1465);
nor U1501 (N_1501,N_1455,N_1495);
or U1502 (N_1502,N_1471,N_1496);
nand U1503 (N_1503,N_1459,N_1467);
nand U1504 (N_1504,N_1475,N_1499);
nand U1505 (N_1505,N_1492,N_1452);
and U1506 (N_1506,N_1498,N_1478);
or U1507 (N_1507,N_1482,N_1472);
nand U1508 (N_1508,N_1487,N_1462);
nand U1509 (N_1509,N_1476,N_1457);
nor U1510 (N_1510,N_1485,N_1490);
nand U1511 (N_1511,N_1464,N_1460);
nand U1512 (N_1512,N_1451,N_1488);
or U1513 (N_1513,N_1470,N_1483);
nand U1514 (N_1514,N_1491,N_1484);
nand U1515 (N_1515,N_1453,N_1454);
or U1516 (N_1516,N_1466,N_1456);
or U1517 (N_1517,N_1477,N_1461);
nand U1518 (N_1518,N_1497,N_1489);
nand U1519 (N_1519,N_1479,N_1493);
nand U1520 (N_1520,N_1480,N_1468);
xor U1521 (N_1521,N_1458,N_1474);
nand U1522 (N_1522,N_1473,N_1463);
nor U1523 (N_1523,N_1494,N_1450);
nand U1524 (N_1524,N_1481,N_1486);
nand U1525 (N_1525,N_1472,N_1474);
and U1526 (N_1526,N_1452,N_1457);
nand U1527 (N_1527,N_1454,N_1483);
or U1528 (N_1528,N_1487,N_1499);
or U1529 (N_1529,N_1464,N_1452);
or U1530 (N_1530,N_1482,N_1484);
nand U1531 (N_1531,N_1478,N_1459);
nor U1532 (N_1532,N_1457,N_1461);
or U1533 (N_1533,N_1492,N_1456);
or U1534 (N_1534,N_1492,N_1465);
or U1535 (N_1535,N_1492,N_1464);
or U1536 (N_1536,N_1456,N_1477);
or U1537 (N_1537,N_1482,N_1457);
or U1538 (N_1538,N_1464,N_1493);
and U1539 (N_1539,N_1461,N_1454);
nand U1540 (N_1540,N_1468,N_1492);
and U1541 (N_1541,N_1454,N_1499);
or U1542 (N_1542,N_1471,N_1478);
nand U1543 (N_1543,N_1484,N_1464);
nor U1544 (N_1544,N_1450,N_1496);
nor U1545 (N_1545,N_1473,N_1476);
nor U1546 (N_1546,N_1480,N_1487);
and U1547 (N_1547,N_1485,N_1453);
nand U1548 (N_1548,N_1453,N_1489);
and U1549 (N_1549,N_1491,N_1488);
and U1550 (N_1550,N_1510,N_1543);
and U1551 (N_1551,N_1516,N_1524);
xnor U1552 (N_1552,N_1507,N_1512);
and U1553 (N_1553,N_1506,N_1535);
nand U1554 (N_1554,N_1541,N_1518);
nor U1555 (N_1555,N_1547,N_1504);
or U1556 (N_1556,N_1533,N_1540);
or U1557 (N_1557,N_1530,N_1542);
nor U1558 (N_1558,N_1513,N_1529);
nand U1559 (N_1559,N_1503,N_1546);
or U1560 (N_1560,N_1511,N_1520);
xnor U1561 (N_1561,N_1537,N_1505);
nor U1562 (N_1562,N_1517,N_1527);
nand U1563 (N_1563,N_1534,N_1514);
or U1564 (N_1564,N_1544,N_1521);
xnor U1565 (N_1565,N_1515,N_1531);
and U1566 (N_1566,N_1548,N_1502);
nor U1567 (N_1567,N_1523,N_1500);
or U1568 (N_1568,N_1532,N_1522);
xor U1569 (N_1569,N_1549,N_1525);
and U1570 (N_1570,N_1526,N_1519);
or U1571 (N_1571,N_1509,N_1539);
nand U1572 (N_1572,N_1545,N_1528);
and U1573 (N_1573,N_1501,N_1538);
or U1574 (N_1574,N_1536,N_1508);
or U1575 (N_1575,N_1538,N_1529);
and U1576 (N_1576,N_1500,N_1507);
and U1577 (N_1577,N_1508,N_1510);
nor U1578 (N_1578,N_1545,N_1526);
and U1579 (N_1579,N_1523,N_1530);
nand U1580 (N_1580,N_1521,N_1539);
or U1581 (N_1581,N_1505,N_1541);
nor U1582 (N_1582,N_1543,N_1513);
nor U1583 (N_1583,N_1517,N_1523);
nor U1584 (N_1584,N_1535,N_1508);
and U1585 (N_1585,N_1540,N_1504);
nand U1586 (N_1586,N_1536,N_1548);
nor U1587 (N_1587,N_1509,N_1520);
nor U1588 (N_1588,N_1535,N_1548);
nand U1589 (N_1589,N_1534,N_1505);
and U1590 (N_1590,N_1500,N_1542);
nor U1591 (N_1591,N_1525,N_1533);
xnor U1592 (N_1592,N_1534,N_1528);
nor U1593 (N_1593,N_1532,N_1516);
and U1594 (N_1594,N_1511,N_1505);
nor U1595 (N_1595,N_1500,N_1503);
and U1596 (N_1596,N_1518,N_1519);
or U1597 (N_1597,N_1548,N_1529);
nand U1598 (N_1598,N_1522,N_1511);
nand U1599 (N_1599,N_1512,N_1522);
nand U1600 (N_1600,N_1586,N_1588);
or U1601 (N_1601,N_1593,N_1579);
and U1602 (N_1602,N_1583,N_1599);
or U1603 (N_1603,N_1585,N_1596);
nor U1604 (N_1604,N_1566,N_1561);
nand U1605 (N_1605,N_1598,N_1572);
or U1606 (N_1606,N_1589,N_1551);
nand U1607 (N_1607,N_1577,N_1574);
or U1608 (N_1608,N_1590,N_1595);
or U1609 (N_1609,N_1557,N_1555);
and U1610 (N_1610,N_1562,N_1563);
nor U1611 (N_1611,N_1556,N_1554);
or U1612 (N_1612,N_1584,N_1567);
or U1613 (N_1613,N_1581,N_1570);
or U1614 (N_1614,N_1576,N_1568);
nor U1615 (N_1615,N_1560,N_1553);
and U1616 (N_1616,N_1575,N_1552);
and U1617 (N_1617,N_1597,N_1573);
and U1618 (N_1618,N_1571,N_1580);
and U1619 (N_1619,N_1564,N_1550);
nor U1620 (N_1620,N_1558,N_1587);
and U1621 (N_1621,N_1559,N_1569);
nor U1622 (N_1622,N_1582,N_1592);
xor U1623 (N_1623,N_1591,N_1565);
nand U1624 (N_1624,N_1594,N_1578);
nand U1625 (N_1625,N_1593,N_1565);
nand U1626 (N_1626,N_1555,N_1574);
nor U1627 (N_1627,N_1553,N_1559);
and U1628 (N_1628,N_1596,N_1568);
and U1629 (N_1629,N_1569,N_1580);
nor U1630 (N_1630,N_1597,N_1581);
nand U1631 (N_1631,N_1594,N_1554);
nor U1632 (N_1632,N_1557,N_1585);
nand U1633 (N_1633,N_1597,N_1590);
nor U1634 (N_1634,N_1553,N_1579);
or U1635 (N_1635,N_1595,N_1587);
nand U1636 (N_1636,N_1565,N_1586);
and U1637 (N_1637,N_1572,N_1581);
nor U1638 (N_1638,N_1580,N_1581);
or U1639 (N_1639,N_1562,N_1568);
nand U1640 (N_1640,N_1563,N_1597);
nand U1641 (N_1641,N_1575,N_1569);
nand U1642 (N_1642,N_1583,N_1593);
and U1643 (N_1643,N_1570,N_1566);
and U1644 (N_1644,N_1593,N_1598);
nand U1645 (N_1645,N_1573,N_1596);
xnor U1646 (N_1646,N_1597,N_1588);
and U1647 (N_1647,N_1564,N_1582);
or U1648 (N_1648,N_1581,N_1577);
nor U1649 (N_1649,N_1560,N_1583);
nand U1650 (N_1650,N_1637,N_1634);
or U1651 (N_1651,N_1605,N_1624);
and U1652 (N_1652,N_1636,N_1613);
or U1653 (N_1653,N_1627,N_1641);
nor U1654 (N_1654,N_1647,N_1619);
nor U1655 (N_1655,N_1607,N_1618);
or U1656 (N_1656,N_1640,N_1626);
or U1657 (N_1657,N_1604,N_1645);
nor U1658 (N_1658,N_1629,N_1649);
and U1659 (N_1659,N_1602,N_1628);
nand U1660 (N_1660,N_1615,N_1616);
nand U1661 (N_1661,N_1633,N_1606);
nor U1662 (N_1662,N_1614,N_1623);
and U1663 (N_1663,N_1631,N_1638);
nand U1664 (N_1664,N_1646,N_1603);
nand U1665 (N_1665,N_1635,N_1642);
nor U1666 (N_1666,N_1617,N_1643);
or U1667 (N_1667,N_1608,N_1648);
nor U1668 (N_1668,N_1620,N_1644);
nand U1669 (N_1669,N_1621,N_1610);
and U1670 (N_1670,N_1639,N_1612);
nand U1671 (N_1671,N_1611,N_1601);
or U1672 (N_1672,N_1625,N_1609);
and U1673 (N_1673,N_1632,N_1600);
nor U1674 (N_1674,N_1622,N_1630);
nand U1675 (N_1675,N_1620,N_1612);
and U1676 (N_1676,N_1629,N_1614);
or U1677 (N_1677,N_1649,N_1630);
nand U1678 (N_1678,N_1619,N_1636);
nand U1679 (N_1679,N_1613,N_1638);
or U1680 (N_1680,N_1602,N_1601);
or U1681 (N_1681,N_1638,N_1649);
nand U1682 (N_1682,N_1620,N_1633);
or U1683 (N_1683,N_1647,N_1646);
nor U1684 (N_1684,N_1630,N_1644);
or U1685 (N_1685,N_1631,N_1644);
or U1686 (N_1686,N_1615,N_1634);
nor U1687 (N_1687,N_1616,N_1639);
nor U1688 (N_1688,N_1614,N_1622);
and U1689 (N_1689,N_1601,N_1630);
nand U1690 (N_1690,N_1606,N_1627);
and U1691 (N_1691,N_1609,N_1622);
nor U1692 (N_1692,N_1641,N_1637);
or U1693 (N_1693,N_1613,N_1617);
nor U1694 (N_1694,N_1647,N_1622);
nor U1695 (N_1695,N_1622,N_1624);
or U1696 (N_1696,N_1628,N_1634);
nand U1697 (N_1697,N_1605,N_1647);
nor U1698 (N_1698,N_1638,N_1648);
or U1699 (N_1699,N_1614,N_1645);
and U1700 (N_1700,N_1657,N_1675);
nand U1701 (N_1701,N_1680,N_1690);
and U1702 (N_1702,N_1662,N_1674);
and U1703 (N_1703,N_1667,N_1696);
nor U1704 (N_1704,N_1689,N_1652);
nand U1705 (N_1705,N_1698,N_1655);
nor U1706 (N_1706,N_1682,N_1695);
nand U1707 (N_1707,N_1681,N_1651);
nand U1708 (N_1708,N_1656,N_1659);
nor U1709 (N_1709,N_1676,N_1686);
and U1710 (N_1710,N_1692,N_1671);
or U1711 (N_1711,N_1699,N_1678);
or U1712 (N_1712,N_1666,N_1653);
and U1713 (N_1713,N_1687,N_1669);
and U1714 (N_1714,N_1685,N_1679);
nand U1715 (N_1715,N_1663,N_1660);
or U1716 (N_1716,N_1668,N_1677);
or U1717 (N_1717,N_1683,N_1691);
xor U1718 (N_1718,N_1650,N_1694);
or U1719 (N_1719,N_1658,N_1688);
or U1720 (N_1720,N_1665,N_1693);
xor U1721 (N_1721,N_1661,N_1684);
and U1722 (N_1722,N_1673,N_1697);
or U1723 (N_1723,N_1672,N_1654);
nand U1724 (N_1724,N_1670,N_1664);
nor U1725 (N_1725,N_1699,N_1670);
nor U1726 (N_1726,N_1669,N_1654);
or U1727 (N_1727,N_1678,N_1658);
nor U1728 (N_1728,N_1658,N_1657);
nand U1729 (N_1729,N_1652,N_1691);
nor U1730 (N_1730,N_1681,N_1657);
or U1731 (N_1731,N_1699,N_1651);
nand U1732 (N_1732,N_1670,N_1668);
nor U1733 (N_1733,N_1659,N_1699);
nand U1734 (N_1734,N_1673,N_1681);
and U1735 (N_1735,N_1679,N_1692);
nor U1736 (N_1736,N_1671,N_1678);
or U1737 (N_1737,N_1686,N_1653);
and U1738 (N_1738,N_1655,N_1660);
nor U1739 (N_1739,N_1652,N_1665);
nor U1740 (N_1740,N_1674,N_1690);
or U1741 (N_1741,N_1686,N_1673);
or U1742 (N_1742,N_1686,N_1671);
nor U1743 (N_1743,N_1663,N_1698);
and U1744 (N_1744,N_1673,N_1693);
nand U1745 (N_1745,N_1660,N_1671);
xor U1746 (N_1746,N_1699,N_1656);
and U1747 (N_1747,N_1675,N_1666);
or U1748 (N_1748,N_1664,N_1675);
nor U1749 (N_1749,N_1662,N_1679);
nor U1750 (N_1750,N_1734,N_1725);
nor U1751 (N_1751,N_1744,N_1714);
nor U1752 (N_1752,N_1748,N_1715);
or U1753 (N_1753,N_1730,N_1749);
and U1754 (N_1754,N_1706,N_1717);
nor U1755 (N_1755,N_1703,N_1713);
or U1756 (N_1756,N_1728,N_1737);
nand U1757 (N_1757,N_1736,N_1708);
xor U1758 (N_1758,N_1712,N_1739);
xor U1759 (N_1759,N_1727,N_1711);
or U1760 (N_1760,N_1731,N_1741);
nand U1761 (N_1761,N_1743,N_1704);
nand U1762 (N_1762,N_1700,N_1723);
or U1763 (N_1763,N_1746,N_1720);
and U1764 (N_1764,N_1732,N_1729);
xnor U1765 (N_1765,N_1722,N_1716);
nor U1766 (N_1766,N_1705,N_1745);
nand U1767 (N_1767,N_1726,N_1740);
nor U1768 (N_1768,N_1721,N_1718);
and U1769 (N_1769,N_1742,N_1702);
or U1770 (N_1770,N_1733,N_1710);
and U1771 (N_1771,N_1709,N_1707);
nand U1772 (N_1772,N_1701,N_1719);
and U1773 (N_1773,N_1738,N_1724);
nand U1774 (N_1774,N_1735,N_1747);
and U1775 (N_1775,N_1747,N_1748);
or U1776 (N_1776,N_1740,N_1725);
nor U1777 (N_1777,N_1721,N_1748);
nand U1778 (N_1778,N_1714,N_1711);
nand U1779 (N_1779,N_1735,N_1725);
or U1780 (N_1780,N_1707,N_1725);
xnor U1781 (N_1781,N_1726,N_1705);
or U1782 (N_1782,N_1717,N_1734);
nor U1783 (N_1783,N_1741,N_1715);
or U1784 (N_1784,N_1704,N_1719);
or U1785 (N_1785,N_1729,N_1721);
or U1786 (N_1786,N_1719,N_1729);
or U1787 (N_1787,N_1716,N_1747);
or U1788 (N_1788,N_1711,N_1739);
or U1789 (N_1789,N_1707,N_1713);
xnor U1790 (N_1790,N_1721,N_1743);
nor U1791 (N_1791,N_1701,N_1735);
or U1792 (N_1792,N_1704,N_1723);
and U1793 (N_1793,N_1731,N_1710);
nand U1794 (N_1794,N_1726,N_1714);
nand U1795 (N_1795,N_1730,N_1703);
and U1796 (N_1796,N_1732,N_1748);
or U1797 (N_1797,N_1702,N_1715);
or U1798 (N_1798,N_1719,N_1721);
and U1799 (N_1799,N_1712,N_1744);
nor U1800 (N_1800,N_1785,N_1774);
nand U1801 (N_1801,N_1760,N_1759);
and U1802 (N_1802,N_1781,N_1787);
nand U1803 (N_1803,N_1766,N_1768);
or U1804 (N_1804,N_1765,N_1755);
and U1805 (N_1805,N_1792,N_1751);
or U1806 (N_1806,N_1775,N_1779);
and U1807 (N_1807,N_1763,N_1761);
and U1808 (N_1808,N_1750,N_1798);
or U1809 (N_1809,N_1796,N_1772);
nor U1810 (N_1810,N_1762,N_1754);
xnor U1811 (N_1811,N_1776,N_1793);
nand U1812 (N_1812,N_1758,N_1784);
or U1813 (N_1813,N_1764,N_1757);
or U1814 (N_1814,N_1756,N_1777);
and U1815 (N_1815,N_1767,N_1786);
nor U1816 (N_1816,N_1753,N_1773);
nand U1817 (N_1817,N_1771,N_1752);
nor U1818 (N_1818,N_1791,N_1799);
nand U1819 (N_1819,N_1789,N_1790);
or U1820 (N_1820,N_1770,N_1769);
nand U1821 (N_1821,N_1778,N_1788);
or U1822 (N_1822,N_1783,N_1797);
and U1823 (N_1823,N_1782,N_1794);
nand U1824 (N_1824,N_1795,N_1780);
and U1825 (N_1825,N_1778,N_1759);
and U1826 (N_1826,N_1775,N_1773);
nand U1827 (N_1827,N_1799,N_1798);
or U1828 (N_1828,N_1783,N_1776);
and U1829 (N_1829,N_1761,N_1793);
nand U1830 (N_1830,N_1751,N_1789);
nand U1831 (N_1831,N_1753,N_1784);
and U1832 (N_1832,N_1757,N_1775);
nor U1833 (N_1833,N_1775,N_1759);
nand U1834 (N_1834,N_1752,N_1762);
or U1835 (N_1835,N_1761,N_1794);
and U1836 (N_1836,N_1788,N_1765);
nor U1837 (N_1837,N_1772,N_1778);
nor U1838 (N_1838,N_1756,N_1784);
nor U1839 (N_1839,N_1791,N_1752);
nor U1840 (N_1840,N_1781,N_1797);
nand U1841 (N_1841,N_1756,N_1755);
and U1842 (N_1842,N_1769,N_1776);
or U1843 (N_1843,N_1789,N_1755);
nor U1844 (N_1844,N_1794,N_1758);
and U1845 (N_1845,N_1751,N_1762);
nand U1846 (N_1846,N_1774,N_1784);
and U1847 (N_1847,N_1792,N_1750);
or U1848 (N_1848,N_1770,N_1775);
nand U1849 (N_1849,N_1789,N_1763);
or U1850 (N_1850,N_1809,N_1830);
and U1851 (N_1851,N_1824,N_1823);
nor U1852 (N_1852,N_1833,N_1820);
xor U1853 (N_1853,N_1828,N_1806);
and U1854 (N_1854,N_1846,N_1829);
or U1855 (N_1855,N_1849,N_1839);
nor U1856 (N_1856,N_1808,N_1807);
and U1857 (N_1857,N_1844,N_1805);
nand U1858 (N_1858,N_1802,N_1834);
xnor U1859 (N_1859,N_1812,N_1847);
or U1860 (N_1860,N_1821,N_1838);
nor U1861 (N_1861,N_1845,N_1826);
or U1862 (N_1862,N_1804,N_1810);
nand U1863 (N_1863,N_1817,N_1825);
nor U1864 (N_1864,N_1800,N_1803);
or U1865 (N_1865,N_1840,N_1822);
xnor U1866 (N_1866,N_1814,N_1815);
or U1867 (N_1867,N_1801,N_1811);
nand U1868 (N_1868,N_1832,N_1835);
nor U1869 (N_1869,N_1841,N_1831);
and U1870 (N_1870,N_1813,N_1819);
nor U1871 (N_1871,N_1843,N_1827);
nand U1872 (N_1872,N_1842,N_1818);
nand U1873 (N_1873,N_1848,N_1816);
or U1874 (N_1874,N_1837,N_1836);
and U1875 (N_1875,N_1801,N_1824);
or U1876 (N_1876,N_1824,N_1831);
nor U1877 (N_1877,N_1843,N_1816);
and U1878 (N_1878,N_1829,N_1831);
nor U1879 (N_1879,N_1815,N_1840);
or U1880 (N_1880,N_1825,N_1821);
nor U1881 (N_1881,N_1808,N_1849);
nor U1882 (N_1882,N_1800,N_1824);
and U1883 (N_1883,N_1834,N_1805);
nor U1884 (N_1884,N_1843,N_1832);
nor U1885 (N_1885,N_1835,N_1807);
or U1886 (N_1886,N_1815,N_1836);
and U1887 (N_1887,N_1825,N_1820);
or U1888 (N_1888,N_1845,N_1807);
and U1889 (N_1889,N_1841,N_1804);
and U1890 (N_1890,N_1839,N_1832);
nand U1891 (N_1891,N_1827,N_1847);
or U1892 (N_1892,N_1827,N_1835);
nand U1893 (N_1893,N_1812,N_1809);
or U1894 (N_1894,N_1800,N_1823);
nand U1895 (N_1895,N_1827,N_1848);
nand U1896 (N_1896,N_1839,N_1820);
or U1897 (N_1897,N_1804,N_1845);
nand U1898 (N_1898,N_1836,N_1824);
and U1899 (N_1899,N_1809,N_1813);
nand U1900 (N_1900,N_1879,N_1883);
nand U1901 (N_1901,N_1861,N_1887);
nor U1902 (N_1902,N_1858,N_1865);
or U1903 (N_1903,N_1896,N_1863);
nor U1904 (N_1904,N_1851,N_1864);
nand U1905 (N_1905,N_1869,N_1873);
or U1906 (N_1906,N_1890,N_1888);
nand U1907 (N_1907,N_1859,N_1898);
nand U1908 (N_1908,N_1872,N_1881);
or U1909 (N_1909,N_1899,N_1854);
nand U1910 (N_1910,N_1852,N_1886);
nand U1911 (N_1911,N_1877,N_1878);
and U1912 (N_1912,N_1857,N_1894);
nor U1913 (N_1913,N_1860,N_1889);
nor U1914 (N_1914,N_1871,N_1855);
or U1915 (N_1915,N_1882,N_1876);
xnor U1916 (N_1916,N_1892,N_1870);
or U1917 (N_1917,N_1853,N_1884);
and U1918 (N_1918,N_1895,N_1867);
nor U1919 (N_1919,N_1880,N_1862);
nand U1920 (N_1920,N_1875,N_1868);
or U1921 (N_1921,N_1897,N_1893);
or U1922 (N_1922,N_1850,N_1866);
and U1923 (N_1923,N_1885,N_1856);
and U1924 (N_1924,N_1874,N_1891);
and U1925 (N_1925,N_1881,N_1863);
nor U1926 (N_1926,N_1858,N_1850);
or U1927 (N_1927,N_1868,N_1863);
xnor U1928 (N_1928,N_1867,N_1878);
nor U1929 (N_1929,N_1889,N_1875);
nand U1930 (N_1930,N_1895,N_1865);
and U1931 (N_1931,N_1888,N_1889);
nand U1932 (N_1932,N_1896,N_1852);
nand U1933 (N_1933,N_1855,N_1864);
and U1934 (N_1934,N_1889,N_1859);
nand U1935 (N_1935,N_1897,N_1858);
or U1936 (N_1936,N_1856,N_1870);
nor U1937 (N_1937,N_1887,N_1871);
nand U1938 (N_1938,N_1882,N_1867);
and U1939 (N_1939,N_1887,N_1854);
or U1940 (N_1940,N_1883,N_1878);
nor U1941 (N_1941,N_1888,N_1885);
nand U1942 (N_1942,N_1874,N_1861);
nand U1943 (N_1943,N_1859,N_1857);
nor U1944 (N_1944,N_1879,N_1859);
or U1945 (N_1945,N_1856,N_1875);
nand U1946 (N_1946,N_1858,N_1880);
or U1947 (N_1947,N_1895,N_1875);
xnor U1948 (N_1948,N_1868,N_1861);
and U1949 (N_1949,N_1851,N_1887);
or U1950 (N_1950,N_1909,N_1932);
nor U1951 (N_1951,N_1929,N_1941);
nand U1952 (N_1952,N_1945,N_1906);
nand U1953 (N_1953,N_1904,N_1940);
and U1954 (N_1954,N_1914,N_1938);
and U1955 (N_1955,N_1918,N_1942);
nand U1956 (N_1956,N_1913,N_1920);
nor U1957 (N_1957,N_1924,N_1933);
nor U1958 (N_1958,N_1939,N_1907);
xnor U1959 (N_1959,N_1912,N_1916);
or U1960 (N_1960,N_1917,N_1923);
or U1961 (N_1961,N_1949,N_1931);
and U1962 (N_1962,N_1901,N_1903);
nand U1963 (N_1963,N_1928,N_1926);
and U1964 (N_1964,N_1905,N_1934);
or U1965 (N_1965,N_1946,N_1925);
nand U1966 (N_1966,N_1935,N_1915);
nor U1967 (N_1967,N_1910,N_1911);
nor U1968 (N_1968,N_1937,N_1948);
nand U1969 (N_1969,N_1921,N_1922);
or U1970 (N_1970,N_1919,N_1947);
nor U1971 (N_1971,N_1900,N_1930);
or U1972 (N_1972,N_1908,N_1902);
xnor U1973 (N_1973,N_1936,N_1943);
nor U1974 (N_1974,N_1944,N_1927);
or U1975 (N_1975,N_1900,N_1948);
nand U1976 (N_1976,N_1946,N_1910);
or U1977 (N_1977,N_1947,N_1946);
or U1978 (N_1978,N_1949,N_1932);
nand U1979 (N_1979,N_1944,N_1921);
or U1980 (N_1980,N_1947,N_1935);
xnor U1981 (N_1981,N_1915,N_1936);
nor U1982 (N_1982,N_1910,N_1919);
or U1983 (N_1983,N_1933,N_1937);
nor U1984 (N_1984,N_1941,N_1931);
nor U1985 (N_1985,N_1945,N_1928);
nor U1986 (N_1986,N_1930,N_1929);
or U1987 (N_1987,N_1946,N_1908);
nand U1988 (N_1988,N_1902,N_1921);
xor U1989 (N_1989,N_1943,N_1914);
xnor U1990 (N_1990,N_1939,N_1918);
and U1991 (N_1991,N_1907,N_1903);
or U1992 (N_1992,N_1900,N_1945);
and U1993 (N_1993,N_1916,N_1902);
and U1994 (N_1994,N_1933,N_1916);
nand U1995 (N_1995,N_1928,N_1918);
nand U1996 (N_1996,N_1927,N_1943);
nand U1997 (N_1997,N_1941,N_1905);
or U1998 (N_1998,N_1905,N_1943);
or U1999 (N_1999,N_1934,N_1911);
nand U2000 (N_2000,N_1966,N_1967);
nor U2001 (N_2001,N_1989,N_1973);
or U2002 (N_2002,N_1986,N_1995);
nand U2003 (N_2003,N_1954,N_1971);
or U2004 (N_2004,N_1968,N_1957);
and U2005 (N_2005,N_1970,N_1975);
xnor U2006 (N_2006,N_1983,N_1956);
or U2007 (N_2007,N_1976,N_1965);
or U2008 (N_2008,N_1960,N_1996);
nand U2009 (N_2009,N_1979,N_1992);
nand U2010 (N_2010,N_1981,N_1969);
nor U2011 (N_2011,N_1964,N_1980);
nand U2012 (N_2012,N_1998,N_1984);
nor U2013 (N_2013,N_1963,N_1974);
and U2014 (N_2014,N_1959,N_1990);
nor U2015 (N_2015,N_1999,N_1987);
or U2016 (N_2016,N_1993,N_1985);
nor U2017 (N_2017,N_1994,N_1950);
nor U2018 (N_2018,N_1991,N_1962);
nor U2019 (N_2019,N_1982,N_1953);
or U2020 (N_2020,N_1988,N_1997);
and U2021 (N_2021,N_1978,N_1955);
or U2022 (N_2022,N_1972,N_1952);
and U2023 (N_2023,N_1977,N_1958);
or U2024 (N_2024,N_1951,N_1961);
nand U2025 (N_2025,N_1950,N_1980);
or U2026 (N_2026,N_1990,N_1997);
nand U2027 (N_2027,N_1987,N_1966);
nor U2028 (N_2028,N_1970,N_1973);
and U2029 (N_2029,N_1961,N_1972);
nor U2030 (N_2030,N_1971,N_1969);
nand U2031 (N_2031,N_1982,N_1975);
and U2032 (N_2032,N_1985,N_1956);
or U2033 (N_2033,N_1994,N_1957);
or U2034 (N_2034,N_1977,N_1960);
and U2035 (N_2035,N_1985,N_1952);
nor U2036 (N_2036,N_1957,N_1989);
nand U2037 (N_2037,N_1987,N_1963);
nor U2038 (N_2038,N_1958,N_1974);
nor U2039 (N_2039,N_1973,N_1998);
nor U2040 (N_2040,N_1992,N_1978);
xor U2041 (N_2041,N_1987,N_1998);
or U2042 (N_2042,N_1971,N_1957);
and U2043 (N_2043,N_1974,N_1952);
nand U2044 (N_2044,N_1999,N_1997);
nand U2045 (N_2045,N_1970,N_1994);
nor U2046 (N_2046,N_1954,N_1972);
nor U2047 (N_2047,N_1958,N_1984);
nor U2048 (N_2048,N_1998,N_1957);
or U2049 (N_2049,N_1980,N_1985);
nor U2050 (N_2050,N_2013,N_2044);
or U2051 (N_2051,N_2000,N_2003);
nand U2052 (N_2052,N_2041,N_2039);
nor U2053 (N_2053,N_2015,N_2020);
nand U2054 (N_2054,N_2035,N_2004);
and U2055 (N_2055,N_2008,N_2022);
and U2056 (N_2056,N_2027,N_2006);
or U2057 (N_2057,N_2001,N_2014);
or U2058 (N_2058,N_2025,N_2033);
nor U2059 (N_2059,N_2046,N_2031);
nand U2060 (N_2060,N_2034,N_2032);
or U2061 (N_2061,N_2021,N_2002);
or U2062 (N_2062,N_2010,N_2017);
nor U2063 (N_2063,N_2038,N_2023);
nand U2064 (N_2064,N_2036,N_2029);
nand U2065 (N_2065,N_2048,N_2042);
and U2066 (N_2066,N_2026,N_2011);
and U2067 (N_2067,N_2005,N_2049);
nand U2068 (N_2068,N_2018,N_2030);
and U2069 (N_2069,N_2007,N_2009);
and U2070 (N_2070,N_2043,N_2028);
or U2071 (N_2071,N_2012,N_2047);
and U2072 (N_2072,N_2016,N_2019);
or U2073 (N_2073,N_2040,N_2037);
or U2074 (N_2074,N_2045,N_2024);
nor U2075 (N_2075,N_2003,N_2046);
or U2076 (N_2076,N_2011,N_2014);
nand U2077 (N_2077,N_2037,N_2012);
nand U2078 (N_2078,N_2009,N_2036);
nor U2079 (N_2079,N_2007,N_2017);
or U2080 (N_2080,N_2037,N_2006);
or U2081 (N_2081,N_2043,N_2046);
nand U2082 (N_2082,N_2021,N_2028);
and U2083 (N_2083,N_2009,N_2013);
and U2084 (N_2084,N_2044,N_2028);
and U2085 (N_2085,N_2016,N_2011);
nor U2086 (N_2086,N_2038,N_2001);
nand U2087 (N_2087,N_2020,N_2013);
nand U2088 (N_2088,N_2031,N_2024);
nor U2089 (N_2089,N_2046,N_2033);
and U2090 (N_2090,N_2008,N_2046);
xor U2091 (N_2091,N_2039,N_2004);
or U2092 (N_2092,N_2029,N_2004);
nand U2093 (N_2093,N_2028,N_2035);
nor U2094 (N_2094,N_2024,N_2047);
nand U2095 (N_2095,N_2021,N_2044);
nor U2096 (N_2096,N_2032,N_2046);
nand U2097 (N_2097,N_2034,N_2000);
nand U2098 (N_2098,N_2014,N_2047);
or U2099 (N_2099,N_2026,N_2015);
and U2100 (N_2100,N_2091,N_2051);
and U2101 (N_2101,N_2077,N_2068);
nand U2102 (N_2102,N_2089,N_2066);
nand U2103 (N_2103,N_2098,N_2082);
and U2104 (N_2104,N_2074,N_2079);
nor U2105 (N_2105,N_2083,N_2096);
xor U2106 (N_2106,N_2072,N_2058);
nor U2107 (N_2107,N_2055,N_2071);
and U2108 (N_2108,N_2086,N_2060);
or U2109 (N_2109,N_2062,N_2061);
nand U2110 (N_2110,N_2088,N_2054);
or U2111 (N_2111,N_2097,N_2076);
nand U2112 (N_2112,N_2087,N_2075);
nor U2113 (N_2113,N_2059,N_2090);
nor U2114 (N_2114,N_2095,N_2052);
nand U2115 (N_2115,N_2092,N_2080);
or U2116 (N_2116,N_2084,N_2069);
or U2117 (N_2117,N_2099,N_2065);
or U2118 (N_2118,N_2057,N_2078);
and U2119 (N_2119,N_2070,N_2073);
nand U2120 (N_2120,N_2063,N_2094);
nor U2121 (N_2121,N_2056,N_2050);
nor U2122 (N_2122,N_2067,N_2085);
or U2123 (N_2123,N_2064,N_2081);
or U2124 (N_2124,N_2093,N_2053);
or U2125 (N_2125,N_2067,N_2060);
nand U2126 (N_2126,N_2051,N_2054);
and U2127 (N_2127,N_2065,N_2058);
nor U2128 (N_2128,N_2081,N_2093);
and U2129 (N_2129,N_2051,N_2080);
nand U2130 (N_2130,N_2071,N_2074);
nand U2131 (N_2131,N_2096,N_2077);
nor U2132 (N_2132,N_2087,N_2074);
and U2133 (N_2133,N_2093,N_2066);
nor U2134 (N_2134,N_2098,N_2065);
nand U2135 (N_2135,N_2094,N_2090);
nor U2136 (N_2136,N_2056,N_2067);
and U2137 (N_2137,N_2097,N_2083);
nor U2138 (N_2138,N_2055,N_2066);
or U2139 (N_2139,N_2073,N_2063);
nor U2140 (N_2140,N_2062,N_2054);
nor U2141 (N_2141,N_2089,N_2076);
xnor U2142 (N_2142,N_2073,N_2087);
nor U2143 (N_2143,N_2075,N_2077);
and U2144 (N_2144,N_2056,N_2066);
or U2145 (N_2145,N_2095,N_2093);
nor U2146 (N_2146,N_2072,N_2087);
or U2147 (N_2147,N_2072,N_2079);
nand U2148 (N_2148,N_2076,N_2050);
nand U2149 (N_2149,N_2074,N_2094);
and U2150 (N_2150,N_2132,N_2101);
and U2151 (N_2151,N_2109,N_2145);
nor U2152 (N_2152,N_2125,N_2128);
nor U2153 (N_2153,N_2119,N_2118);
or U2154 (N_2154,N_2146,N_2105);
and U2155 (N_2155,N_2100,N_2130);
or U2156 (N_2156,N_2103,N_2140);
nand U2157 (N_2157,N_2116,N_2144);
or U2158 (N_2158,N_2115,N_2108);
and U2159 (N_2159,N_2148,N_2117);
or U2160 (N_2160,N_2135,N_2123);
nand U2161 (N_2161,N_2102,N_2126);
nor U2162 (N_2162,N_2142,N_2139);
or U2163 (N_2163,N_2136,N_2131);
and U2164 (N_2164,N_2111,N_2110);
nand U2165 (N_2165,N_2141,N_2112);
nand U2166 (N_2166,N_2149,N_2124);
and U2167 (N_2167,N_2143,N_2114);
nor U2168 (N_2168,N_2127,N_2104);
nor U2169 (N_2169,N_2138,N_2121);
and U2170 (N_2170,N_2122,N_2106);
and U2171 (N_2171,N_2113,N_2120);
and U2172 (N_2172,N_2137,N_2147);
nand U2173 (N_2173,N_2107,N_2129);
nor U2174 (N_2174,N_2133,N_2134);
nand U2175 (N_2175,N_2105,N_2149);
or U2176 (N_2176,N_2144,N_2100);
and U2177 (N_2177,N_2146,N_2135);
or U2178 (N_2178,N_2119,N_2108);
or U2179 (N_2179,N_2133,N_2117);
and U2180 (N_2180,N_2135,N_2140);
or U2181 (N_2181,N_2101,N_2115);
and U2182 (N_2182,N_2106,N_2141);
or U2183 (N_2183,N_2116,N_2145);
nor U2184 (N_2184,N_2121,N_2145);
and U2185 (N_2185,N_2124,N_2123);
nand U2186 (N_2186,N_2138,N_2123);
nand U2187 (N_2187,N_2141,N_2124);
and U2188 (N_2188,N_2133,N_2108);
and U2189 (N_2189,N_2120,N_2102);
nor U2190 (N_2190,N_2102,N_2128);
or U2191 (N_2191,N_2101,N_2139);
nor U2192 (N_2192,N_2102,N_2136);
nand U2193 (N_2193,N_2109,N_2127);
and U2194 (N_2194,N_2131,N_2123);
or U2195 (N_2195,N_2125,N_2127);
nor U2196 (N_2196,N_2137,N_2140);
nor U2197 (N_2197,N_2141,N_2102);
and U2198 (N_2198,N_2116,N_2131);
nor U2199 (N_2199,N_2137,N_2110);
nor U2200 (N_2200,N_2170,N_2174);
nor U2201 (N_2201,N_2156,N_2159);
or U2202 (N_2202,N_2167,N_2198);
and U2203 (N_2203,N_2197,N_2195);
nand U2204 (N_2204,N_2152,N_2183);
nand U2205 (N_2205,N_2192,N_2176);
nand U2206 (N_2206,N_2158,N_2187);
or U2207 (N_2207,N_2161,N_2178);
nor U2208 (N_2208,N_2194,N_2199);
nor U2209 (N_2209,N_2185,N_2196);
and U2210 (N_2210,N_2190,N_2155);
or U2211 (N_2211,N_2157,N_2162);
and U2212 (N_2212,N_2151,N_2154);
nand U2213 (N_2213,N_2177,N_2150);
and U2214 (N_2214,N_2179,N_2164);
nor U2215 (N_2215,N_2153,N_2181);
or U2216 (N_2216,N_2166,N_2186);
nor U2217 (N_2217,N_2165,N_2193);
or U2218 (N_2218,N_2175,N_2184);
nand U2219 (N_2219,N_2182,N_2191);
and U2220 (N_2220,N_2160,N_2173);
and U2221 (N_2221,N_2189,N_2172);
nand U2222 (N_2222,N_2180,N_2168);
nor U2223 (N_2223,N_2171,N_2188);
and U2224 (N_2224,N_2163,N_2169);
nand U2225 (N_2225,N_2191,N_2183);
nor U2226 (N_2226,N_2169,N_2196);
nand U2227 (N_2227,N_2168,N_2193);
or U2228 (N_2228,N_2155,N_2198);
nand U2229 (N_2229,N_2192,N_2153);
nor U2230 (N_2230,N_2171,N_2172);
nand U2231 (N_2231,N_2188,N_2178);
or U2232 (N_2232,N_2162,N_2169);
and U2233 (N_2233,N_2184,N_2181);
nand U2234 (N_2234,N_2191,N_2195);
nand U2235 (N_2235,N_2172,N_2198);
nor U2236 (N_2236,N_2156,N_2197);
nor U2237 (N_2237,N_2196,N_2192);
or U2238 (N_2238,N_2180,N_2153);
and U2239 (N_2239,N_2197,N_2168);
or U2240 (N_2240,N_2178,N_2199);
nor U2241 (N_2241,N_2184,N_2198);
and U2242 (N_2242,N_2165,N_2179);
nand U2243 (N_2243,N_2183,N_2190);
or U2244 (N_2244,N_2185,N_2157);
or U2245 (N_2245,N_2168,N_2199);
nand U2246 (N_2246,N_2180,N_2187);
and U2247 (N_2247,N_2178,N_2177);
nor U2248 (N_2248,N_2199,N_2155);
nand U2249 (N_2249,N_2163,N_2196);
nand U2250 (N_2250,N_2209,N_2215);
and U2251 (N_2251,N_2228,N_2211);
nor U2252 (N_2252,N_2248,N_2214);
nor U2253 (N_2253,N_2226,N_2229);
nor U2254 (N_2254,N_2233,N_2249);
nand U2255 (N_2255,N_2224,N_2241);
nand U2256 (N_2256,N_2204,N_2243);
or U2257 (N_2257,N_2216,N_2231);
nor U2258 (N_2258,N_2235,N_2200);
nor U2259 (N_2259,N_2237,N_2219);
nand U2260 (N_2260,N_2223,N_2242);
and U2261 (N_2261,N_2207,N_2203);
nor U2262 (N_2262,N_2205,N_2220);
nor U2263 (N_2263,N_2222,N_2202);
or U2264 (N_2264,N_2238,N_2232);
nor U2265 (N_2265,N_2244,N_2236);
nand U2266 (N_2266,N_2208,N_2227);
and U2267 (N_2267,N_2240,N_2230);
and U2268 (N_2268,N_2245,N_2225);
and U2269 (N_2269,N_2206,N_2239);
and U2270 (N_2270,N_2212,N_2217);
nand U2271 (N_2271,N_2247,N_2218);
nand U2272 (N_2272,N_2221,N_2210);
and U2273 (N_2273,N_2213,N_2246);
xor U2274 (N_2274,N_2234,N_2201);
nor U2275 (N_2275,N_2213,N_2230);
nor U2276 (N_2276,N_2249,N_2240);
or U2277 (N_2277,N_2228,N_2246);
and U2278 (N_2278,N_2222,N_2209);
or U2279 (N_2279,N_2234,N_2200);
and U2280 (N_2280,N_2237,N_2248);
or U2281 (N_2281,N_2231,N_2215);
nor U2282 (N_2282,N_2216,N_2200);
nand U2283 (N_2283,N_2234,N_2206);
nand U2284 (N_2284,N_2236,N_2237);
nor U2285 (N_2285,N_2246,N_2230);
nand U2286 (N_2286,N_2234,N_2211);
and U2287 (N_2287,N_2247,N_2243);
nand U2288 (N_2288,N_2218,N_2209);
and U2289 (N_2289,N_2208,N_2215);
xnor U2290 (N_2290,N_2227,N_2229);
nor U2291 (N_2291,N_2206,N_2228);
nor U2292 (N_2292,N_2203,N_2227);
nor U2293 (N_2293,N_2224,N_2213);
nor U2294 (N_2294,N_2240,N_2216);
or U2295 (N_2295,N_2225,N_2219);
and U2296 (N_2296,N_2240,N_2210);
nand U2297 (N_2297,N_2225,N_2239);
nor U2298 (N_2298,N_2249,N_2213);
or U2299 (N_2299,N_2217,N_2231);
or U2300 (N_2300,N_2285,N_2276);
nand U2301 (N_2301,N_2279,N_2294);
or U2302 (N_2302,N_2252,N_2277);
nor U2303 (N_2303,N_2288,N_2269);
and U2304 (N_2304,N_2257,N_2295);
nor U2305 (N_2305,N_2273,N_2263);
nor U2306 (N_2306,N_2290,N_2272);
and U2307 (N_2307,N_2274,N_2268);
or U2308 (N_2308,N_2253,N_2283);
nor U2309 (N_2309,N_2264,N_2284);
nand U2310 (N_2310,N_2251,N_2292);
and U2311 (N_2311,N_2250,N_2281);
nand U2312 (N_2312,N_2266,N_2265);
and U2313 (N_2313,N_2270,N_2296);
or U2314 (N_2314,N_2289,N_2267);
and U2315 (N_2315,N_2291,N_2256);
or U2316 (N_2316,N_2280,N_2297);
and U2317 (N_2317,N_2255,N_2298);
or U2318 (N_2318,N_2262,N_2275);
or U2319 (N_2319,N_2282,N_2271);
nor U2320 (N_2320,N_2258,N_2299);
and U2321 (N_2321,N_2278,N_2261);
and U2322 (N_2322,N_2260,N_2287);
and U2323 (N_2323,N_2259,N_2286);
nor U2324 (N_2324,N_2293,N_2254);
and U2325 (N_2325,N_2258,N_2296);
or U2326 (N_2326,N_2295,N_2289);
and U2327 (N_2327,N_2250,N_2269);
nand U2328 (N_2328,N_2267,N_2276);
or U2329 (N_2329,N_2288,N_2255);
and U2330 (N_2330,N_2261,N_2268);
nand U2331 (N_2331,N_2268,N_2275);
and U2332 (N_2332,N_2262,N_2282);
xor U2333 (N_2333,N_2269,N_2257);
and U2334 (N_2334,N_2269,N_2259);
nor U2335 (N_2335,N_2276,N_2268);
and U2336 (N_2336,N_2294,N_2297);
nor U2337 (N_2337,N_2298,N_2276);
or U2338 (N_2338,N_2295,N_2281);
nor U2339 (N_2339,N_2278,N_2250);
nand U2340 (N_2340,N_2285,N_2268);
and U2341 (N_2341,N_2267,N_2298);
nor U2342 (N_2342,N_2279,N_2250);
or U2343 (N_2343,N_2257,N_2274);
nor U2344 (N_2344,N_2268,N_2250);
nand U2345 (N_2345,N_2286,N_2262);
or U2346 (N_2346,N_2251,N_2264);
or U2347 (N_2347,N_2250,N_2261);
and U2348 (N_2348,N_2278,N_2283);
nand U2349 (N_2349,N_2251,N_2297);
nand U2350 (N_2350,N_2303,N_2335);
nand U2351 (N_2351,N_2317,N_2319);
and U2352 (N_2352,N_2348,N_2347);
or U2353 (N_2353,N_2314,N_2323);
nand U2354 (N_2354,N_2334,N_2327);
or U2355 (N_2355,N_2330,N_2304);
and U2356 (N_2356,N_2324,N_2332);
or U2357 (N_2357,N_2336,N_2302);
or U2358 (N_2358,N_2326,N_2313);
nand U2359 (N_2359,N_2309,N_2341);
nand U2360 (N_2360,N_2343,N_2318);
or U2361 (N_2361,N_2321,N_2339);
or U2362 (N_2362,N_2316,N_2306);
nand U2363 (N_2363,N_2301,N_2346);
or U2364 (N_2364,N_2331,N_2300);
nand U2365 (N_2365,N_2338,N_2315);
nor U2366 (N_2366,N_2305,N_2325);
and U2367 (N_2367,N_2344,N_2310);
or U2368 (N_2368,N_2320,N_2342);
or U2369 (N_2369,N_2308,N_2322);
and U2370 (N_2370,N_2333,N_2345);
and U2371 (N_2371,N_2340,N_2328);
or U2372 (N_2372,N_2337,N_2307);
nand U2373 (N_2373,N_2312,N_2349);
or U2374 (N_2374,N_2329,N_2311);
or U2375 (N_2375,N_2300,N_2316);
or U2376 (N_2376,N_2320,N_2328);
or U2377 (N_2377,N_2334,N_2333);
nor U2378 (N_2378,N_2324,N_2335);
and U2379 (N_2379,N_2328,N_2310);
nor U2380 (N_2380,N_2344,N_2341);
nand U2381 (N_2381,N_2339,N_2315);
or U2382 (N_2382,N_2316,N_2338);
nor U2383 (N_2383,N_2313,N_2332);
nor U2384 (N_2384,N_2316,N_2311);
nor U2385 (N_2385,N_2308,N_2302);
and U2386 (N_2386,N_2338,N_2326);
or U2387 (N_2387,N_2338,N_2348);
or U2388 (N_2388,N_2315,N_2308);
nor U2389 (N_2389,N_2311,N_2309);
nor U2390 (N_2390,N_2327,N_2313);
nand U2391 (N_2391,N_2322,N_2319);
nand U2392 (N_2392,N_2329,N_2304);
nor U2393 (N_2393,N_2344,N_2312);
or U2394 (N_2394,N_2334,N_2307);
and U2395 (N_2395,N_2323,N_2322);
or U2396 (N_2396,N_2338,N_2344);
and U2397 (N_2397,N_2305,N_2324);
xnor U2398 (N_2398,N_2338,N_2320);
nor U2399 (N_2399,N_2347,N_2320);
nand U2400 (N_2400,N_2380,N_2366);
nand U2401 (N_2401,N_2361,N_2351);
nand U2402 (N_2402,N_2368,N_2386);
nor U2403 (N_2403,N_2371,N_2365);
nand U2404 (N_2404,N_2391,N_2394);
nor U2405 (N_2405,N_2387,N_2374);
or U2406 (N_2406,N_2355,N_2358);
xor U2407 (N_2407,N_2369,N_2398);
or U2408 (N_2408,N_2353,N_2388);
or U2409 (N_2409,N_2396,N_2377);
nand U2410 (N_2410,N_2378,N_2367);
and U2411 (N_2411,N_2382,N_2362);
nand U2412 (N_2412,N_2350,N_2376);
nor U2413 (N_2413,N_2357,N_2392);
nor U2414 (N_2414,N_2360,N_2399);
nor U2415 (N_2415,N_2372,N_2375);
and U2416 (N_2416,N_2363,N_2379);
or U2417 (N_2417,N_2381,N_2356);
or U2418 (N_2418,N_2393,N_2373);
and U2419 (N_2419,N_2383,N_2370);
and U2420 (N_2420,N_2352,N_2384);
xnor U2421 (N_2421,N_2397,N_2385);
and U2422 (N_2422,N_2395,N_2389);
and U2423 (N_2423,N_2359,N_2364);
and U2424 (N_2424,N_2390,N_2354);
nand U2425 (N_2425,N_2354,N_2357);
and U2426 (N_2426,N_2392,N_2382);
nand U2427 (N_2427,N_2384,N_2391);
nand U2428 (N_2428,N_2375,N_2351);
nor U2429 (N_2429,N_2364,N_2355);
or U2430 (N_2430,N_2375,N_2388);
and U2431 (N_2431,N_2364,N_2378);
or U2432 (N_2432,N_2357,N_2368);
and U2433 (N_2433,N_2375,N_2368);
and U2434 (N_2434,N_2365,N_2352);
nor U2435 (N_2435,N_2368,N_2387);
or U2436 (N_2436,N_2386,N_2363);
and U2437 (N_2437,N_2353,N_2395);
nand U2438 (N_2438,N_2392,N_2395);
nand U2439 (N_2439,N_2350,N_2372);
nand U2440 (N_2440,N_2356,N_2390);
nand U2441 (N_2441,N_2381,N_2350);
nor U2442 (N_2442,N_2354,N_2360);
and U2443 (N_2443,N_2398,N_2395);
and U2444 (N_2444,N_2374,N_2361);
nor U2445 (N_2445,N_2387,N_2371);
and U2446 (N_2446,N_2360,N_2386);
and U2447 (N_2447,N_2377,N_2385);
and U2448 (N_2448,N_2382,N_2394);
nand U2449 (N_2449,N_2375,N_2359);
nand U2450 (N_2450,N_2443,N_2409);
nand U2451 (N_2451,N_2444,N_2438);
or U2452 (N_2452,N_2429,N_2431);
and U2453 (N_2453,N_2404,N_2436);
or U2454 (N_2454,N_2410,N_2440);
nand U2455 (N_2455,N_2427,N_2406);
nor U2456 (N_2456,N_2435,N_2407);
nand U2457 (N_2457,N_2419,N_2437);
nand U2458 (N_2458,N_2402,N_2441);
and U2459 (N_2459,N_2434,N_2405);
nand U2460 (N_2460,N_2422,N_2401);
or U2461 (N_2461,N_2421,N_2420);
or U2462 (N_2462,N_2447,N_2412);
nand U2463 (N_2463,N_2433,N_2400);
and U2464 (N_2464,N_2445,N_2424);
nor U2465 (N_2465,N_2432,N_2426);
and U2466 (N_2466,N_2413,N_2428);
nand U2467 (N_2467,N_2417,N_2442);
nand U2468 (N_2468,N_2448,N_2403);
and U2469 (N_2469,N_2423,N_2430);
or U2470 (N_2470,N_2418,N_2411);
nand U2471 (N_2471,N_2415,N_2449);
nand U2472 (N_2472,N_2414,N_2439);
nand U2473 (N_2473,N_2425,N_2446);
and U2474 (N_2474,N_2416,N_2408);
or U2475 (N_2475,N_2447,N_2427);
and U2476 (N_2476,N_2445,N_2448);
nor U2477 (N_2477,N_2420,N_2406);
nor U2478 (N_2478,N_2407,N_2427);
nor U2479 (N_2479,N_2405,N_2406);
and U2480 (N_2480,N_2429,N_2425);
nor U2481 (N_2481,N_2412,N_2416);
or U2482 (N_2482,N_2427,N_2403);
and U2483 (N_2483,N_2430,N_2400);
or U2484 (N_2484,N_2422,N_2445);
nor U2485 (N_2485,N_2417,N_2421);
nor U2486 (N_2486,N_2410,N_2414);
and U2487 (N_2487,N_2439,N_2406);
nor U2488 (N_2488,N_2442,N_2443);
and U2489 (N_2489,N_2424,N_2440);
nand U2490 (N_2490,N_2445,N_2436);
and U2491 (N_2491,N_2404,N_2417);
and U2492 (N_2492,N_2434,N_2402);
nor U2493 (N_2493,N_2408,N_2423);
nor U2494 (N_2494,N_2416,N_2406);
nor U2495 (N_2495,N_2435,N_2437);
nor U2496 (N_2496,N_2408,N_2417);
and U2497 (N_2497,N_2446,N_2407);
nand U2498 (N_2498,N_2449,N_2410);
nand U2499 (N_2499,N_2434,N_2435);
nor U2500 (N_2500,N_2457,N_2464);
nand U2501 (N_2501,N_2482,N_2486);
and U2502 (N_2502,N_2470,N_2487);
xor U2503 (N_2503,N_2491,N_2497);
nor U2504 (N_2504,N_2469,N_2463);
and U2505 (N_2505,N_2452,N_2461);
nor U2506 (N_2506,N_2485,N_2471);
nand U2507 (N_2507,N_2476,N_2488);
and U2508 (N_2508,N_2474,N_2465);
and U2509 (N_2509,N_2455,N_2493);
and U2510 (N_2510,N_2462,N_2450);
and U2511 (N_2511,N_2495,N_2460);
and U2512 (N_2512,N_2484,N_2480);
and U2513 (N_2513,N_2451,N_2489);
or U2514 (N_2514,N_2492,N_2483);
nor U2515 (N_2515,N_2475,N_2479);
and U2516 (N_2516,N_2458,N_2454);
xor U2517 (N_2517,N_2498,N_2478);
nand U2518 (N_2518,N_2473,N_2490);
nor U2519 (N_2519,N_2496,N_2467);
xnor U2520 (N_2520,N_2466,N_2459);
nor U2521 (N_2521,N_2468,N_2494);
nor U2522 (N_2522,N_2499,N_2472);
or U2523 (N_2523,N_2456,N_2453);
or U2524 (N_2524,N_2477,N_2481);
and U2525 (N_2525,N_2493,N_2456);
and U2526 (N_2526,N_2490,N_2458);
or U2527 (N_2527,N_2469,N_2465);
nor U2528 (N_2528,N_2475,N_2461);
nor U2529 (N_2529,N_2480,N_2463);
nor U2530 (N_2530,N_2470,N_2489);
and U2531 (N_2531,N_2456,N_2466);
and U2532 (N_2532,N_2478,N_2491);
and U2533 (N_2533,N_2479,N_2451);
or U2534 (N_2534,N_2498,N_2494);
nand U2535 (N_2535,N_2499,N_2483);
nor U2536 (N_2536,N_2486,N_2471);
or U2537 (N_2537,N_2463,N_2489);
nor U2538 (N_2538,N_2479,N_2494);
nand U2539 (N_2539,N_2453,N_2460);
nand U2540 (N_2540,N_2458,N_2496);
or U2541 (N_2541,N_2464,N_2476);
nor U2542 (N_2542,N_2492,N_2480);
or U2543 (N_2543,N_2493,N_2465);
nor U2544 (N_2544,N_2497,N_2456);
and U2545 (N_2545,N_2487,N_2467);
nand U2546 (N_2546,N_2458,N_2455);
nand U2547 (N_2547,N_2490,N_2476);
or U2548 (N_2548,N_2466,N_2486);
nor U2549 (N_2549,N_2455,N_2462);
nand U2550 (N_2550,N_2514,N_2522);
and U2551 (N_2551,N_2538,N_2516);
nand U2552 (N_2552,N_2546,N_2520);
nand U2553 (N_2553,N_2536,N_2519);
nor U2554 (N_2554,N_2507,N_2532);
nor U2555 (N_2555,N_2542,N_2500);
and U2556 (N_2556,N_2528,N_2512);
nor U2557 (N_2557,N_2511,N_2513);
nand U2558 (N_2558,N_2541,N_2535);
and U2559 (N_2559,N_2502,N_2534);
or U2560 (N_2560,N_2545,N_2518);
and U2561 (N_2561,N_2517,N_2526);
nand U2562 (N_2562,N_2537,N_2530);
nor U2563 (N_2563,N_2533,N_2515);
xor U2564 (N_2564,N_2505,N_2529);
or U2565 (N_2565,N_2523,N_2540);
or U2566 (N_2566,N_2527,N_2544);
and U2567 (N_2567,N_2543,N_2547);
or U2568 (N_2568,N_2521,N_2504);
nand U2569 (N_2569,N_2548,N_2531);
nor U2570 (N_2570,N_2539,N_2508);
and U2571 (N_2571,N_2509,N_2549);
xor U2572 (N_2572,N_2501,N_2524);
nand U2573 (N_2573,N_2510,N_2525);
or U2574 (N_2574,N_2506,N_2503);
nand U2575 (N_2575,N_2543,N_2516);
nand U2576 (N_2576,N_2504,N_2533);
and U2577 (N_2577,N_2521,N_2503);
nor U2578 (N_2578,N_2539,N_2534);
and U2579 (N_2579,N_2525,N_2543);
and U2580 (N_2580,N_2539,N_2524);
nor U2581 (N_2581,N_2513,N_2545);
nor U2582 (N_2582,N_2545,N_2521);
nand U2583 (N_2583,N_2531,N_2500);
and U2584 (N_2584,N_2506,N_2520);
nand U2585 (N_2585,N_2525,N_2537);
nor U2586 (N_2586,N_2501,N_2538);
and U2587 (N_2587,N_2523,N_2510);
nand U2588 (N_2588,N_2539,N_2549);
and U2589 (N_2589,N_2534,N_2501);
or U2590 (N_2590,N_2518,N_2512);
nor U2591 (N_2591,N_2521,N_2522);
nand U2592 (N_2592,N_2511,N_2526);
or U2593 (N_2593,N_2520,N_2528);
and U2594 (N_2594,N_2522,N_2543);
nor U2595 (N_2595,N_2524,N_2525);
nand U2596 (N_2596,N_2546,N_2548);
and U2597 (N_2597,N_2522,N_2502);
nor U2598 (N_2598,N_2515,N_2506);
and U2599 (N_2599,N_2523,N_2500);
and U2600 (N_2600,N_2575,N_2560);
nor U2601 (N_2601,N_2593,N_2557);
xor U2602 (N_2602,N_2589,N_2577);
nor U2603 (N_2603,N_2588,N_2586);
and U2604 (N_2604,N_2562,N_2552);
and U2605 (N_2605,N_2554,N_2596);
or U2606 (N_2606,N_2578,N_2567);
and U2607 (N_2607,N_2598,N_2566);
and U2608 (N_2608,N_2574,N_2565);
and U2609 (N_2609,N_2582,N_2592);
nor U2610 (N_2610,N_2556,N_2561);
and U2611 (N_2611,N_2558,N_2584);
nand U2612 (N_2612,N_2597,N_2573);
and U2613 (N_2613,N_2595,N_2568);
and U2614 (N_2614,N_2580,N_2559);
xnor U2615 (N_2615,N_2583,N_2551);
nand U2616 (N_2616,N_2564,N_2571);
and U2617 (N_2617,N_2590,N_2594);
and U2618 (N_2618,N_2555,N_2581);
nor U2619 (N_2619,N_2572,N_2599);
nand U2620 (N_2620,N_2570,N_2550);
or U2621 (N_2621,N_2569,N_2553);
xnor U2622 (N_2622,N_2576,N_2587);
and U2623 (N_2623,N_2579,N_2585);
and U2624 (N_2624,N_2591,N_2563);
nor U2625 (N_2625,N_2574,N_2566);
nand U2626 (N_2626,N_2577,N_2571);
and U2627 (N_2627,N_2570,N_2555);
nand U2628 (N_2628,N_2573,N_2583);
and U2629 (N_2629,N_2591,N_2565);
nor U2630 (N_2630,N_2573,N_2596);
nor U2631 (N_2631,N_2552,N_2569);
nand U2632 (N_2632,N_2566,N_2562);
xnor U2633 (N_2633,N_2584,N_2597);
nor U2634 (N_2634,N_2554,N_2595);
nand U2635 (N_2635,N_2596,N_2556);
nor U2636 (N_2636,N_2574,N_2569);
or U2637 (N_2637,N_2582,N_2577);
and U2638 (N_2638,N_2572,N_2569);
nor U2639 (N_2639,N_2591,N_2581);
and U2640 (N_2640,N_2564,N_2570);
or U2641 (N_2641,N_2568,N_2593);
and U2642 (N_2642,N_2561,N_2551);
and U2643 (N_2643,N_2555,N_2595);
nor U2644 (N_2644,N_2566,N_2581);
or U2645 (N_2645,N_2584,N_2573);
or U2646 (N_2646,N_2575,N_2561);
or U2647 (N_2647,N_2550,N_2567);
nand U2648 (N_2648,N_2561,N_2564);
nand U2649 (N_2649,N_2564,N_2572);
or U2650 (N_2650,N_2608,N_2620);
or U2651 (N_2651,N_2613,N_2619);
and U2652 (N_2652,N_2645,N_2617);
nand U2653 (N_2653,N_2614,N_2629);
nor U2654 (N_2654,N_2648,N_2649);
nor U2655 (N_2655,N_2607,N_2628);
xnor U2656 (N_2656,N_2611,N_2636);
or U2657 (N_2657,N_2603,N_2612);
and U2658 (N_2658,N_2601,N_2621);
and U2659 (N_2659,N_2618,N_2643);
nor U2660 (N_2660,N_2647,N_2602);
nor U2661 (N_2661,N_2635,N_2616);
nor U2662 (N_2662,N_2600,N_2627);
nand U2663 (N_2663,N_2630,N_2646);
or U2664 (N_2664,N_2637,N_2644);
or U2665 (N_2665,N_2638,N_2639);
nor U2666 (N_2666,N_2606,N_2631);
or U2667 (N_2667,N_2605,N_2633);
and U2668 (N_2668,N_2642,N_2624);
and U2669 (N_2669,N_2641,N_2626);
nand U2670 (N_2670,N_2640,N_2632);
and U2671 (N_2671,N_2622,N_2609);
nand U2672 (N_2672,N_2604,N_2634);
or U2673 (N_2673,N_2625,N_2610);
and U2674 (N_2674,N_2623,N_2615);
or U2675 (N_2675,N_2602,N_2626);
and U2676 (N_2676,N_2645,N_2621);
nand U2677 (N_2677,N_2617,N_2639);
or U2678 (N_2678,N_2625,N_2607);
nor U2679 (N_2679,N_2603,N_2604);
and U2680 (N_2680,N_2620,N_2625);
xnor U2681 (N_2681,N_2620,N_2612);
and U2682 (N_2682,N_2614,N_2625);
or U2683 (N_2683,N_2616,N_2632);
nor U2684 (N_2684,N_2604,N_2623);
or U2685 (N_2685,N_2648,N_2614);
or U2686 (N_2686,N_2602,N_2640);
or U2687 (N_2687,N_2606,N_2643);
nor U2688 (N_2688,N_2641,N_2640);
and U2689 (N_2689,N_2609,N_2602);
nor U2690 (N_2690,N_2603,N_2602);
nand U2691 (N_2691,N_2628,N_2627);
nand U2692 (N_2692,N_2639,N_2640);
nor U2693 (N_2693,N_2618,N_2627);
nor U2694 (N_2694,N_2633,N_2648);
or U2695 (N_2695,N_2607,N_2624);
nor U2696 (N_2696,N_2609,N_2615);
or U2697 (N_2697,N_2601,N_2623);
and U2698 (N_2698,N_2628,N_2622);
nand U2699 (N_2699,N_2610,N_2649);
or U2700 (N_2700,N_2678,N_2691);
nand U2701 (N_2701,N_2681,N_2661);
or U2702 (N_2702,N_2654,N_2693);
or U2703 (N_2703,N_2672,N_2688);
nor U2704 (N_2704,N_2666,N_2686);
or U2705 (N_2705,N_2656,N_2684);
nor U2706 (N_2706,N_2669,N_2650);
nor U2707 (N_2707,N_2673,N_2683);
nand U2708 (N_2708,N_2663,N_2692);
and U2709 (N_2709,N_2677,N_2652);
and U2710 (N_2710,N_2653,N_2689);
or U2711 (N_2711,N_2665,N_2664);
and U2712 (N_2712,N_2694,N_2657);
nand U2713 (N_2713,N_2667,N_2687);
nand U2714 (N_2714,N_2658,N_2659);
and U2715 (N_2715,N_2699,N_2698);
or U2716 (N_2716,N_2670,N_2682);
nor U2717 (N_2717,N_2679,N_2668);
nand U2718 (N_2718,N_2697,N_2674);
and U2719 (N_2719,N_2696,N_2695);
nor U2720 (N_2720,N_2675,N_2690);
nor U2721 (N_2721,N_2662,N_2685);
nor U2722 (N_2722,N_2671,N_2660);
nor U2723 (N_2723,N_2680,N_2676);
nor U2724 (N_2724,N_2655,N_2651);
and U2725 (N_2725,N_2650,N_2653);
nand U2726 (N_2726,N_2673,N_2699);
and U2727 (N_2727,N_2692,N_2673);
or U2728 (N_2728,N_2653,N_2696);
nor U2729 (N_2729,N_2651,N_2653);
nand U2730 (N_2730,N_2650,N_2673);
or U2731 (N_2731,N_2666,N_2683);
and U2732 (N_2732,N_2689,N_2687);
nor U2733 (N_2733,N_2665,N_2653);
and U2734 (N_2734,N_2665,N_2674);
nand U2735 (N_2735,N_2659,N_2657);
nor U2736 (N_2736,N_2676,N_2665);
and U2737 (N_2737,N_2691,N_2666);
nor U2738 (N_2738,N_2697,N_2685);
and U2739 (N_2739,N_2681,N_2677);
or U2740 (N_2740,N_2680,N_2682);
nand U2741 (N_2741,N_2662,N_2694);
or U2742 (N_2742,N_2681,N_2693);
or U2743 (N_2743,N_2679,N_2660);
or U2744 (N_2744,N_2679,N_2696);
nand U2745 (N_2745,N_2660,N_2694);
or U2746 (N_2746,N_2650,N_2679);
nor U2747 (N_2747,N_2664,N_2663);
nor U2748 (N_2748,N_2699,N_2667);
nor U2749 (N_2749,N_2670,N_2688);
or U2750 (N_2750,N_2744,N_2747);
or U2751 (N_2751,N_2706,N_2746);
or U2752 (N_2752,N_2711,N_2742);
nand U2753 (N_2753,N_2740,N_2716);
nor U2754 (N_2754,N_2729,N_2739);
nand U2755 (N_2755,N_2743,N_2737);
and U2756 (N_2756,N_2710,N_2707);
and U2757 (N_2757,N_2701,N_2705);
nand U2758 (N_2758,N_2726,N_2718);
and U2759 (N_2759,N_2703,N_2736);
or U2760 (N_2760,N_2700,N_2722);
xnor U2761 (N_2761,N_2709,N_2721);
nand U2762 (N_2762,N_2708,N_2748);
or U2763 (N_2763,N_2732,N_2713);
nand U2764 (N_2764,N_2725,N_2714);
or U2765 (N_2765,N_2741,N_2723);
and U2766 (N_2766,N_2704,N_2727);
nand U2767 (N_2767,N_2717,N_2728);
or U2768 (N_2768,N_2724,N_2733);
xnor U2769 (N_2769,N_2715,N_2745);
or U2770 (N_2770,N_2719,N_2734);
nand U2771 (N_2771,N_2702,N_2720);
nor U2772 (N_2772,N_2731,N_2730);
nand U2773 (N_2773,N_2735,N_2738);
or U2774 (N_2774,N_2749,N_2712);
nor U2775 (N_2775,N_2733,N_2732);
and U2776 (N_2776,N_2725,N_2716);
nand U2777 (N_2777,N_2717,N_2729);
nor U2778 (N_2778,N_2730,N_2708);
nand U2779 (N_2779,N_2706,N_2733);
xnor U2780 (N_2780,N_2704,N_2716);
and U2781 (N_2781,N_2722,N_2703);
or U2782 (N_2782,N_2717,N_2706);
and U2783 (N_2783,N_2706,N_2708);
or U2784 (N_2784,N_2704,N_2718);
and U2785 (N_2785,N_2729,N_2711);
and U2786 (N_2786,N_2748,N_2738);
and U2787 (N_2787,N_2703,N_2725);
and U2788 (N_2788,N_2748,N_2736);
nor U2789 (N_2789,N_2748,N_2714);
or U2790 (N_2790,N_2729,N_2718);
nand U2791 (N_2791,N_2727,N_2745);
and U2792 (N_2792,N_2749,N_2733);
nand U2793 (N_2793,N_2708,N_2721);
and U2794 (N_2794,N_2722,N_2738);
nand U2795 (N_2795,N_2727,N_2743);
or U2796 (N_2796,N_2740,N_2727);
nand U2797 (N_2797,N_2719,N_2749);
nor U2798 (N_2798,N_2720,N_2727);
nand U2799 (N_2799,N_2742,N_2706);
xnor U2800 (N_2800,N_2779,N_2758);
and U2801 (N_2801,N_2753,N_2751);
and U2802 (N_2802,N_2795,N_2768);
or U2803 (N_2803,N_2790,N_2770);
nand U2804 (N_2804,N_2789,N_2776);
and U2805 (N_2805,N_2754,N_2761);
nor U2806 (N_2806,N_2766,N_2778);
or U2807 (N_2807,N_2785,N_2796);
nand U2808 (N_2808,N_2760,N_2786);
and U2809 (N_2809,N_2788,N_2771);
nand U2810 (N_2810,N_2777,N_2764);
nand U2811 (N_2811,N_2780,N_2755);
or U2812 (N_2812,N_2783,N_2799);
nand U2813 (N_2813,N_2767,N_2798);
nand U2814 (N_2814,N_2782,N_2787);
and U2815 (N_2815,N_2794,N_2792);
nor U2816 (N_2816,N_2765,N_2793);
nor U2817 (N_2817,N_2791,N_2757);
nor U2818 (N_2818,N_2775,N_2784);
or U2819 (N_2819,N_2769,N_2772);
nand U2820 (N_2820,N_2781,N_2756);
nor U2821 (N_2821,N_2763,N_2797);
and U2822 (N_2822,N_2750,N_2773);
or U2823 (N_2823,N_2774,N_2759);
xnor U2824 (N_2824,N_2762,N_2752);
and U2825 (N_2825,N_2757,N_2783);
nand U2826 (N_2826,N_2794,N_2791);
nand U2827 (N_2827,N_2769,N_2758);
nand U2828 (N_2828,N_2756,N_2776);
and U2829 (N_2829,N_2769,N_2755);
nand U2830 (N_2830,N_2753,N_2750);
nand U2831 (N_2831,N_2784,N_2786);
and U2832 (N_2832,N_2760,N_2770);
nor U2833 (N_2833,N_2777,N_2793);
or U2834 (N_2834,N_2776,N_2783);
nand U2835 (N_2835,N_2773,N_2760);
nand U2836 (N_2836,N_2776,N_2766);
nor U2837 (N_2837,N_2773,N_2771);
nor U2838 (N_2838,N_2774,N_2785);
or U2839 (N_2839,N_2762,N_2768);
nand U2840 (N_2840,N_2770,N_2797);
nand U2841 (N_2841,N_2775,N_2751);
nand U2842 (N_2842,N_2761,N_2787);
nor U2843 (N_2843,N_2764,N_2761);
and U2844 (N_2844,N_2752,N_2751);
nor U2845 (N_2845,N_2798,N_2795);
and U2846 (N_2846,N_2753,N_2754);
nor U2847 (N_2847,N_2767,N_2784);
nor U2848 (N_2848,N_2786,N_2764);
and U2849 (N_2849,N_2756,N_2799);
or U2850 (N_2850,N_2843,N_2824);
nor U2851 (N_2851,N_2828,N_2837);
and U2852 (N_2852,N_2823,N_2833);
or U2853 (N_2853,N_2825,N_2819);
nand U2854 (N_2854,N_2846,N_2812);
nand U2855 (N_2855,N_2827,N_2818);
and U2856 (N_2856,N_2832,N_2849);
nor U2857 (N_2857,N_2807,N_2805);
nor U2858 (N_2858,N_2841,N_2810);
and U2859 (N_2859,N_2809,N_2826);
and U2860 (N_2860,N_2811,N_2808);
or U2861 (N_2861,N_2845,N_2815);
xor U2862 (N_2862,N_2802,N_2806);
and U2863 (N_2863,N_2847,N_2842);
nand U2864 (N_2864,N_2816,N_2836);
xor U2865 (N_2865,N_2800,N_2831);
or U2866 (N_2866,N_2817,N_2801);
or U2867 (N_2867,N_2829,N_2848);
and U2868 (N_2868,N_2804,N_2830);
nand U2869 (N_2869,N_2803,N_2840);
or U2870 (N_2870,N_2835,N_2820);
and U2871 (N_2871,N_2813,N_2822);
xnor U2872 (N_2872,N_2844,N_2839);
and U2873 (N_2873,N_2838,N_2814);
nor U2874 (N_2874,N_2834,N_2821);
and U2875 (N_2875,N_2833,N_2839);
nor U2876 (N_2876,N_2839,N_2847);
nor U2877 (N_2877,N_2831,N_2848);
and U2878 (N_2878,N_2801,N_2826);
or U2879 (N_2879,N_2835,N_2838);
and U2880 (N_2880,N_2835,N_2837);
or U2881 (N_2881,N_2846,N_2845);
and U2882 (N_2882,N_2800,N_2825);
or U2883 (N_2883,N_2840,N_2836);
nor U2884 (N_2884,N_2811,N_2844);
nor U2885 (N_2885,N_2819,N_2828);
and U2886 (N_2886,N_2837,N_2826);
and U2887 (N_2887,N_2834,N_2836);
and U2888 (N_2888,N_2843,N_2800);
nor U2889 (N_2889,N_2822,N_2815);
nand U2890 (N_2890,N_2846,N_2848);
or U2891 (N_2891,N_2813,N_2839);
nand U2892 (N_2892,N_2830,N_2837);
nand U2893 (N_2893,N_2842,N_2809);
or U2894 (N_2894,N_2845,N_2844);
and U2895 (N_2895,N_2800,N_2815);
nand U2896 (N_2896,N_2830,N_2821);
nor U2897 (N_2897,N_2819,N_2841);
and U2898 (N_2898,N_2845,N_2839);
nand U2899 (N_2899,N_2808,N_2803);
nand U2900 (N_2900,N_2859,N_2881);
nor U2901 (N_2901,N_2891,N_2872);
and U2902 (N_2902,N_2875,N_2893);
nor U2903 (N_2903,N_2889,N_2890);
nand U2904 (N_2904,N_2850,N_2853);
nor U2905 (N_2905,N_2880,N_2864);
and U2906 (N_2906,N_2892,N_2861);
nand U2907 (N_2907,N_2855,N_2854);
nand U2908 (N_2908,N_2896,N_2888);
nor U2909 (N_2909,N_2856,N_2871);
xnor U2910 (N_2910,N_2851,N_2866);
and U2911 (N_2911,N_2877,N_2883);
nand U2912 (N_2912,N_2863,N_2882);
and U2913 (N_2913,N_2894,N_2897);
nand U2914 (N_2914,N_2865,N_2878);
or U2915 (N_2915,N_2860,N_2895);
or U2916 (N_2916,N_2884,N_2885);
or U2917 (N_2917,N_2887,N_2874);
or U2918 (N_2918,N_2876,N_2898);
and U2919 (N_2919,N_2869,N_2868);
or U2920 (N_2920,N_2899,N_2852);
and U2921 (N_2921,N_2870,N_2862);
nand U2922 (N_2922,N_2879,N_2857);
nand U2923 (N_2923,N_2867,N_2873);
nand U2924 (N_2924,N_2858,N_2886);
xnor U2925 (N_2925,N_2893,N_2854);
nand U2926 (N_2926,N_2882,N_2898);
nand U2927 (N_2927,N_2880,N_2857);
and U2928 (N_2928,N_2883,N_2893);
nand U2929 (N_2929,N_2866,N_2870);
nor U2930 (N_2930,N_2896,N_2876);
and U2931 (N_2931,N_2866,N_2858);
and U2932 (N_2932,N_2899,N_2853);
xor U2933 (N_2933,N_2850,N_2867);
nand U2934 (N_2934,N_2862,N_2850);
nand U2935 (N_2935,N_2863,N_2850);
nand U2936 (N_2936,N_2882,N_2894);
or U2937 (N_2937,N_2897,N_2898);
nor U2938 (N_2938,N_2859,N_2893);
and U2939 (N_2939,N_2876,N_2879);
nand U2940 (N_2940,N_2874,N_2873);
nand U2941 (N_2941,N_2878,N_2898);
nor U2942 (N_2942,N_2875,N_2866);
nand U2943 (N_2943,N_2893,N_2853);
and U2944 (N_2944,N_2861,N_2897);
nand U2945 (N_2945,N_2853,N_2873);
nand U2946 (N_2946,N_2860,N_2882);
nor U2947 (N_2947,N_2880,N_2856);
or U2948 (N_2948,N_2855,N_2886);
or U2949 (N_2949,N_2874,N_2870);
and U2950 (N_2950,N_2926,N_2947);
nand U2951 (N_2951,N_2932,N_2914);
and U2952 (N_2952,N_2944,N_2915);
nand U2953 (N_2953,N_2920,N_2937);
nor U2954 (N_2954,N_2931,N_2948);
nor U2955 (N_2955,N_2940,N_2903);
nand U2956 (N_2956,N_2930,N_2922);
xnor U2957 (N_2957,N_2943,N_2902);
and U2958 (N_2958,N_2919,N_2941);
nor U2959 (N_2959,N_2901,N_2933);
nor U2960 (N_2960,N_2912,N_2929);
or U2961 (N_2961,N_2935,N_2949);
nor U2962 (N_2962,N_2938,N_2924);
nor U2963 (N_2963,N_2908,N_2906);
and U2964 (N_2964,N_2909,N_2921);
nand U2965 (N_2965,N_2910,N_2934);
and U2966 (N_2966,N_2946,N_2936);
or U2967 (N_2967,N_2939,N_2911);
and U2968 (N_2968,N_2928,N_2916);
or U2969 (N_2969,N_2942,N_2945);
nor U2970 (N_2970,N_2917,N_2923);
or U2971 (N_2971,N_2925,N_2927);
nand U2972 (N_2972,N_2918,N_2907);
nor U2973 (N_2973,N_2900,N_2904);
nand U2974 (N_2974,N_2913,N_2905);
nand U2975 (N_2975,N_2929,N_2909);
nand U2976 (N_2976,N_2941,N_2934);
and U2977 (N_2977,N_2907,N_2905);
or U2978 (N_2978,N_2924,N_2933);
and U2979 (N_2979,N_2941,N_2921);
or U2980 (N_2980,N_2904,N_2916);
and U2981 (N_2981,N_2945,N_2919);
nor U2982 (N_2982,N_2949,N_2922);
or U2983 (N_2983,N_2930,N_2904);
or U2984 (N_2984,N_2931,N_2908);
nor U2985 (N_2985,N_2926,N_2908);
and U2986 (N_2986,N_2925,N_2944);
nor U2987 (N_2987,N_2930,N_2940);
and U2988 (N_2988,N_2940,N_2904);
nor U2989 (N_2989,N_2904,N_2909);
or U2990 (N_2990,N_2913,N_2921);
nor U2991 (N_2991,N_2915,N_2927);
xor U2992 (N_2992,N_2937,N_2930);
and U2993 (N_2993,N_2928,N_2902);
or U2994 (N_2994,N_2931,N_2928);
nand U2995 (N_2995,N_2937,N_2928);
nand U2996 (N_2996,N_2924,N_2918);
and U2997 (N_2997,N_2913,N_2907);
or U2998 (N_2998,N_2918,N_2913);
nand U2999 (N_2999,N_2908,N_2927);
and UO_0 (O_0,N_2992,N_2962);
nand UO_1 (O_1,N_2979,N_2973);
or UO_2 (O_2,N_2958,N_2968);
and UO_3 (O_3,N_2999,N_2964);
or UO_4 (O_4,N_2972,N_2988);
nor UO_5 (O_5,N_2980,N_2983);
and UO_6 (O_6,N_2997,N_2985);
and UO_7 (O_7,N_2971,N_2981);
nand UO_8 (O_8,N_2956,N_2974);
nor UO_9 (O_9,N_2951,N_2986);
nor UO_10 (O_10,N_2967,N_2987);
nor UO_11 (O_11,N_2977,N_2953);
nor UO_12 (O_12,N_2996,N_2952);
and UO_13 (O_13,N_2991,N_2998);
nand UO_14 (O_14,N_2960,N_2966);
and UO_15 (O_15,N_2978,N_2969);
nor UO_16 (O_16,N_2993,N_2982);
nand UO_17 (O_17,N_2970,N_2963);
and UO_18 (O_18,N_2989,N_2957);
nand UO_19 (O_19,N_2975,N_2955);
and UO_20 (O_20,N_2965,N_2954);
and UO_21 (O_21,N_2994,N_2961);
xnor UO_22 (O_22,N_2990,N_2984);
and UO_23 (O_23,N_2950,N_2995);
nor UO_24 (O_24,N_2959,N_2976);
nand UO_25 (O_25,N_2950,N_2968);
nand UO_26 (O_26,N_2996,N_2974);
nor UO_27 (O_27,N_2996,N_2990);
or UO_28 (O_28,N_2986,N_2996);
nand UO_29 (O_29,N_2995,N_2968);
or UO_30 (O_30,N_2994,N_2999);
or UO_31 (O_31,N_2968,N_2952);
and UO_32 (O_32,N_2984,N_2958);
nand UO_33 (O_33,N_2954,N_2971);
or UO_34 (O_34,N_2999,N_2966);
or UO_35 (O_35,N_2954,N_2970);
nor UO_36 (O_36,N_2953,N_2975);
or UO_37 (O_37,N_2963,N_2988);
nor UO_38 (O_38,N_2997,N_2955);
nand UO_39 (O_39,N_2988,N_2991);
or UO_40 (O_40,N_2986,N_2970);
and UO_41 (O_41,N_2954,N_2993);
or UO_42 (O_42,N_2958,N_2996);
and UO_43 (O_43,N_2965,N_2974);
and UO_44 (O_44,N_2993,N_2979);
nor UO_45 (O_45,N_2978,N_2974);
or UO_46 (O_46,N_2951,N_2974);
nor UO_47 (O_47,N_2965,N_2968);
nor UO_48 (O_48,N_2976,N_2963);
nor UO_49 (O_49,N_2955,N_2959);
nor UO_50 (O_50,N_2987,N_2963);
or UO_51 (O_51,N_2952,N_2956);
nor UO_52 (O_52,N_2986,N_2964);
nand UO_53 (O_53,N_2982,N_2975);
xor UO_54 (O_54,N_2994,N_2964);
and UO_55 (O_55,N_2962,N_2952);
nor UO_56 (O_56,N_2970,N_2956);
nor UO_57 (O_57,N_2959,N_2971);
or UO_58 (O_58,N_2986,N_2965);
nand UO_59 (O_59,N_2972,N_2999);
nor UO_60 (O_60,N_2956,N_2955);
and UO_61 (O_61,N_2965,N_2993);
and UO_62 (O_62,N_2976,N_2980);
or UO_63 (O_63,N_2960,N_2988);
or UO_64 (O_64,N_2970,N_2990);
or UO_65 (O_65,N_2982,N_2990);
or UO_66 (O_66,N_2998,N_2981);
nand UO_67 (O_67,N_2960,N_2974);
or UO_68 (O_68,N_2953,N_2951);
and UO_69 (O_69,N_2959,N_2990);
and UO_70 (O_70,N_2977,N_2983);
nand UO_71 (O_71,N_2952,N_2954);
or UO_72 (O_72,N_2984,N_2963);
or UO_73 (O_73,N_2964,N_2980);
and UO_74 (O_74,N_2956,N_2985);
and UO_75 (O_75,N_2957,N_2956);
nor UO_76 (O_76,N_2957,N_2950);
or UO_77 (O_77,N_2978,N_2983);
or UO_78 (O_78,N_2993,N_2997);
and UO_79 (O_79,N_2982,N_2956);
nand UO_80 (O_80,N_2998,N_2950);
nand UO_81 (O_81,N_2954,N_2956);
or UO_82 (O_82,N_2965,N_2971);
and UO_83 (O_83,N_2960,N_2952);
and UO_84 (O_84,N_2956,N_2987);
or UO_85 (O_85,N_2965,N_2959);
and UO_86 (O_86,N_2955,N_2968);
nor UO_87 (O_87,N_2959,N_2961);
nor UO_88 (O_88,N_2966,N_2987);
and UO_89 (O_89,N_2956,N_2969);
and UO_90 (O_90,N_2964,N_2952);
nor UO_91 (O_91,N_2952,N_2993);
nor UO_92 (O_92,N_2991,N_2981);
and UO_93 (O_93,N_2971,N_2963);
nand UO_94 (O_94,N_2964,N_2988);
nor UO_95 (O_95,N_2986,N_2969);
and UO_96 (O_96,N_2992,N_2983);
and UO_97 (O_97,N_2956,N_2992);
or UO_98 (O_98,N_2966,N_2963);
nand UO_99 (O_99,N_2962,N_2988);
nand UO_100 (O_100,N_2993,N_2957);
nand UO_101 (O_101,N_2967,N_2994);
nand UO_102 (O_102,N_2973,N_2966);
and UO_103 (O_103,N_2976,N_2962);
nor UO_104 (O_104,N_2978,N_2967);
or UO_105 (O_105,N_2959,N_2970);
or UO_106 (O_106,N_2976,N_2969);
and UO_107 (O_107,N_2958,N_2994);
nand UO_108 (O_108,N_2953,N_2996);
or UO_109 (O_109,N_2973,N_2951);
or UO_110 (O_110,N_2969,N_2961);
nand UO_111 (O_111,N_2975,N_2964);
nand UO_112 (O_112,N_2998,N_2977);
and UO_113 (O_113,N_2993,N_2959);
and UO_114 (O_114,N_2968,N_2964);
or UO_115 (O_115,N_2978,N_2976);
or UO_116 (O_116,N_2959,N_2966);
nor UO_117 (O_117,N_2983,N_2970);
or UO_118 (O_118,N_2972,N_2994);
or UO_119 (O_119,N_2982,N_2989);
nor UO_120 (O_120,N_2985,N_2959);
or UO_121 (O_121,N_2986,N_2991);
nor UO_122 (O_122,N_2954,N_2950);
nor UO_123 (O_123,N_2957,N_2955);
nand UO_124 (O_124,N_2972,N_2959);
nand UO_125 (O_125,N_2951,N_2996);
nand UO_126 (O_126,N_2957,N_2962);
nor UO_127 (O_127,N_2968,N_2963);
and UO_128 (O_128,N_2984,N_2972);
and UO_129 (O_129,N_2992,N_2959);
and UO_130 (O_130,N_2980,N_2974);
nand UO_131 (O_131,N_2971,N_2956);
or UO_132 (O_132,N_2986,N_2984);
nor UO_133 (O_133,N_2981,N_2980);
or UO_134 (O_134,N_2995,N_2951);
nand UO_135 (O_135,N_2951,N_2969);
and UO_136 (O_136,N_2975,N_2992);
nor UO_137 (O_137,N_2996,N_2975);
or UO_138 (O_138,N_2950,N_2999);
nor UO_139 (O_139,N_2989,N_2973);
and UO_140 (O_140,N_2984,N_2983);
nor UO_141 (O_141,N_2969,N_2982);
or UO_142 (O_142,N_2959,N_2986);
or UO_143 (O_143,N_2957,N_2976);
nor UO_144 (O_144,N_2986,N_2985);
or UO_145 (O_145,N_2956,N_2994);
nand UO_146 (O_146,N_2978,N_2972);
nor UO_147 (O_147,N_2987,N_2951);
nand UO_148 (O_148,N_2951,N_2988);
and UO_149 (O_149,N_2995,N_2972);
nand UO_150 (O_150,N_2969,N_2987);
and UO_151 (O_151,N_2977,N_2956);
or UO_152 (O_152,N_2979,N_2969);
and UO_153 (O_153,N_2962,N_2981);
nor UO_154 (O_154,N_2958,N_2980);
and UO_155 (O_155,N_2983,N_2999);
nor UO_156 (O_156,N_2988,N_2997);
or UO_157 (O_157,N_2974,N_2979);
and UO_158 (O_158,N_2988,N_2967);
nor UO_159 (O_159,N_2961,N_2950);
nand UO_160 (O_160,N_2964,N_2966);
nand UO_161 (O_161,N_2965,N_2973);
nand UO_162 (O_162,N_2961,N_2983);
nand UO_163 (O_163,N_2979,N_2953);
and UO_164 (O_164,N_2982,N_2966);
or UO_165 (O_165,N_2998,N_2996);
or UO_166 (O_166,N_2990,N_2956);
or UO_167 (O_167,N_2952,N_2970);
nand UO_168 (O_168,N_2966,N_2975);
and UO_169 (O_169,N_2968,N_2969);
nand UO_170 (O_170,N_2971,N_2990);
nand UO_171 (O_171,N_2970,N_2964);
and UO_172 (O_172,N_2972,N_2970);
xnor UO_173 (O_173,N_2978,N_2958);
nand UO_174 (O_174,N_2974,N_2990);
nor UO_175 (O_175,N_2956,N_2993);
nor UO_176 (O_176,N_2990,N_2985);
nor UO_177 (O_177,N_2951,N_2963);
or UO_178 (O_178,N_2966,N_2950);
and UO_179 (O_179,N_2995,N_2973);
and UO_180 (O_180,N_2997,N_2979);
and UO_181 (O_181,N_2965,N_2998);
and UO_182 (O_182,N_2960,N_2977);
and UO_183 (O_183,N_2992,N_2986);
nor UO_184 (O_184,N_2994,N_2984);
nand UO_185 (O_185,N_2995,N_2954);
or UO_186 (O_186,N_2986,N_2980);
nand UO_187 (O_187,N_2968,N_2953);
or UO_188 (O_188,N_2969,N_2957);
and UO_189 (O_189,N_2994,N_2986);
and UO_190 (O_190,N_2955,N_2967);
nand UO_191 (O_191,N_2963,N_2990);
nand UO_192 (O_192,N_2979,N_2998);
and UO_193 (O_193,N_2962,N_2985);
nand UO_194 (O_194,N_2993,N_2980);
nor UO_195 (O_195,N_2961,N_2964);
nor UO_196 (O_196,N_2989,N_2966);
nand UO_197 (O_197,N_2965,N_2999);
or UO_198 (O_198,N_2964,N_2974);
nand UO_199 (O_199,N_2986,N_2995);
or UO_200 (O_200,N_2992,N_2957);
nor UO_201 (O_201,N_2958,N_2956);
nor UO_202 (O_202,N_2982,N_2951);
nand UO_203 (O_203,N_2950,N_2990);
nand UO_204 (O_204,N_2965,N_2952);
nand UO_205 (O_205,N_2954,N_2961);
nand UO_206 (O_206,N_2966,N_2970);
nor UO_207 (O_207,N_2993,N_2976);
and UO_208 (O_208,N_2990,N_2976);
and UO_209 (O_209,N_2995,N_2990);
nand UO_210 (O_210,N_2980,N_2984);
or UO_211 (O_211,N_2989,N_2951);
and UO_212 (O_212,N_2967,N_2986);
nor UO_213 (O_213,N_2981,N_2997);
nor UO_214 (O_214,N_2960,N_2983);
or UO_215 (O_215,N_2955,N_2991);
nand UO_216 (O_216,N_2963,N_2954);
nand UO_217 (O_217,N_2997,N_2992);
nand UO_218 (O_218,N_2969,N_2955);
nor UO_219 (O_219,N_2985,N_2961);
xor UO_220 (O_220,N_2985,N_2964);
or UO_221 (O_221,N_2955,N_2964);
nand UO_222 (O_222,N_2987,N_2986);
or UO_223 (O_223,N_2962,N_2967);
nor UO_224 (O_224,N_2972,N_2951);
or UO_225 (O_225,N_2975,N_2963);
nor UO_226 (O_226,N_2999,N_2985);
nand UO_227 (O_227,N_2958,N_2955);
or UO_228 (O_228,N_2983,N_2968);
nor UO_229 (O_229,N_2957,N_2970);
or UO_230 (O_230,N_2988,N_2998);
or UO_231 (O_231,N_2989,N_2972);
nor UO_232 (O_232,N_2954,N_2999);
and UO_233 (O_233,N_2956,N_2998);
and UO_234 (O_234,N_2997,N_2968);
xnor UO_235 (O_235,N_2996,N_2961);
and UO_236 (O_236,N_2956,N_2976);
nand UO_237 (O_237,N_2977,N_2989);
nor UO_238 (O_238,N_2991,N_2952);
nor UO_239 (O_239,N_2982,N_2997);
nand UO_240 (O_240,N_2964,N_2950);
nor UO_241 (O_241,N_2952,N_2992);
nand UO_242 (O_242,N_2964,N_2971);
and UO_243 (O_243,N_2976,N_2986);
nand UO_244 (O_244,N_2960,N_2978);
and UO_245 (O_245,N_2988,N_2968);
nor UO_246 (O_246,N_2987,N_2989);
nor UO_247 (O_247,N_2984,N_2997);
and UO_248 (O_248,N_2964,N_2977);
or UO_249 (O_249,N_2981,N_2987);
nor UO_250 (O_250,N_2951,N_2950);
nor UO_251 (O_251,N_2977,N_2976);
nor UO_252 (O_252,N_2950,N_2982);
nor UO_253 (O_253,N_2992,N_2993);
and UO_254 (O_254,N_2983,N_2991);
nand UO_255 (O_255,N_2982,N_2984);
nand UO_256 (O_256,N_2989,N_2969);
and UO_257 (O_257,N_2957,N_2974);
nor UO_258 (O_258,N_2985,N_2966);
nor UO_259 (O_259,N_2989,N_2958);
nor UO_260 (O_260,N_2991,N_2958);
xor UO_261 (O_261,N_2956,N_2997);
nand UO_262 (O_262,N_2956,N_2986);
nand UO_263 (O_263,N_2983,N_2982);
nand UO_264 (O_264,N_2998,N_2989);
nor UO_265 (O_265,N_2958,N_2995);
or UO_266 (O_266,N_2954,N_2989);
nand UO_267 (O_267,N_2951,N_2998);
nor UO_268 (O_268,N_2964,N_2978);
or UO_269 (O_269,N_2951,N_2957);
and UO_270 (O_270,N_2996,N_2969);
nor UO_271 (O_271,N_2960,N_2950);
and UO_272 (O_272,N_2981,N_2952);
or UO_273 (O_273,N_2987,N_2974);
and UO_274 (O_274,N_2968,N_2971);
and UO_275 (O_275,N_2978,N_2955);
nor UO_276 (O_276,N_2990,N_2966);
or UO_277 (O_277,N_2953,N_2998);
and UO_278 (O_278,N_2983,N_2988);
nor UO_279 (O_279,N_2984,N_2976);
xnor UO_280 (O_280,N_2992,N_2971);
and UO_281 (O_281,N_2951,N_2959);
nor UO_282 (O_282,N_2979,N_2955);
and UO_283 (O_283,N_2962,N_2989);
or UO_284 (O_284,N_2982,N_2962);
nor UO_285 (O_285,N_2982,N_2972);
nand UO_286 (O_286,N_2959,N_2988);
or UO_287 (O_287,N_2970,N_2985);
and UO_288 (O_288,N_2963,N_2986);
or UO_289 (O_289,N_2995,N_2969);
and UO_290 (O_290,N_2993,N_2986);
or UO_291 (O_291,N_2975,N_2971);
and UO_292 (O_292,N_2996,N_2967);
nand UO_293 (O_293,N_2998,N_2976);
and UO_294 (O_294,N_2958,N_2974);
or UO_295 (O_295,N_2962,N_2958);
nor UO_296 (O_296,N_2952,N_2979);
or UO_297 (O_297,N_2973,N_2957);
nor UO_298 (O_298,N_2964,N_2954);
and UO_299 (O_299,N_2971,N_2957);
nand UO_300 (O_300,N_2968,N_2991);
or UO_301 (O_301,N_2961,N_2984);
and UO_302 (O_302,N_2992,N_2950);
or UO_303 (O_303,N_2970,N_2978);
and UO_304 (O_304,N_2997,N_2974);
or UO_305 (O_305,N_2988,N_2996);
and UO_306 (O_306,N_2977,N_2987);
and UO_307 (O_307,N_2989,N_2985);
or UO_308 (O_308,N_2981,N_2953);
and UO_309 (O_309,N_2977,N_2963);
nor UO_310 (O_310,N_2970,N_2993);
nand UO_311 (O_311,N_2961,N_2962);
or UO_312 (O_312,N_2971,N_2973);
and UO_313 (O_313,N_2978,N_2979);
and UO_314 (O_314,N_2992,N_2958);
nor UO_315 (O_315,N_2972,N_2967);
and UO_316 (O_316,N_2972,N_2960);
nor UO_317 (O_317,N_2961,N_2998);
nand UO_318 (O_318,N_2996,N_2957);
nand UO_319 (O_319,N_2992,N_2988);
nand UO_320 (O_320,N_2976,N_2994);
nor UO_321 (O_321,N_2957,N_2979);
nand UO_322 (O_322,N_2952,N_2978);
or UO_323 (O_323,N_2953,N_2976);
or UO_324 (O_324,N_2952,N_2986);
and UO_325 (O_325,N_2984,N_2960);
or UO_326 (O_326,N_2983,N_2957);
nor UO_327 (O_327,N_2976,N_2954);
and UO_328 (O_328,N_2969,N_2965);
or UO_329 (O_329,N_2986,N_2955);
or UO_330 (O_330,N_2997,N_2951);
nand UO_331 (O_331,N_2958,N_2983);
and UO_332 (O_332,N_2978,N_2965);
and UO_333 (O_333,N_2955,N_2974);
nand UO_334 (O_334,N_2985,N_2971);
nand UO_335 (O_335,N_2968,N_2999);
or UO_336 (O_336,N_2995,N_2970);
and UO_337 (O_337,N_2974,N_2992);
or UO_338 (O_338,N_2953,N_2987);
nor UO_339 (O_339,N_2972,N_2987);
and UO_340 (O_340,N_2998,N_2986);
nor UO_341 (O_341,N_2973,N_2950);
xor UO_342 (O_342,N_2974,N_2961);
or UO_343 (O_343,N_2996,N_2966);
nand UO_344 (O_344,N_2971,N_2980);
and UO_345 (O_345,N_2968,N_2966);
nand UO_346 (O_346,N_2958,N_2971);
and UO_347 (O_347,N_2992,N_2990);
or UO_348 (O_348,N_2954,N_2981);
and UO_349 (O_349,N_2983,N_2994);
or UO_350 (O_350,N_2984,N_2988);
or UO_351 (O_351,N_2981,N_2964);
nor UO_352 (O_352,N_2987,N_2991);
nor UO_353 (O_353,N_2967,N_2995);
nor UO_354 (O_354,N_2987,N_2960);
nand UO_355 (O_355,N_2999,N_2998);
and UO_356 (O_356,N_2994,N_2990);
nor UO_357 (O_357,N_2961,N_2991);
nor UO_358 (O_358,N_2985,N_2973);
nand UO_359 (O_359,N_2956,N_2999);
and UO_360 (O_360,N_2957,N_2987);
or UO_361 (O_361,N_2978,N_2999);
or UO_362 (O_362,N_2957,N_2966);
or UO_363 (O_363,N_2968,N_2993);
nand UO_364 (O_364,N_2985,N_2993);
nand UO_365 (O_365,N_2954,N_2960);
nor UO_366 (O_366,N_2982,N_2981);
or UO_367 (O_367,N_2958,N_2998);
or UO_368 (O_368,N_2964,N_2957);
xor UO_369 (O_369,N_2967,N_2979);
nand UO_370 (O_370,N_2992,N_2981);
or UO_371 (O_371,N_2983,N_2975);
nand UO_372 (O_372,N_2954,N_2986);
or UO_373 (O_373,N_2974,N_2989);
and UO_374 (O_374,N_2991,N_2956);
nor UO_375 (O_375,N_2988,N_2985);
nand UO_376 (O_376,N_2981,N_2995);
nor UO_377 (O_377,N_2978,N_2995);
or UO_378 (O_378,N_2970,N_2950);
and UO_379 (O_379,N_2996,N_2991);
or UO_380 (O_380,N_2984,N_2995);
or UO_381 (O_381,N_2994,N_2993);
xnor UO_382 (O_382,N_2960,N_2996);
and UO_383 (O_383,N_2957,N_2982);
nor UO_384 (O_384,N_2999,N_2984);
nor UO_385 (O_385,N_2958,N_2950);
nand UO_386 (O_386,N_2992,N_2966);
nor UO_387 (O_387,N_2967,N_2999);
nand UO_388 (O_388,N_2976,N_2955);
and UO_389 (O_389,N_2996,N_2993);
nand UO_390 (O_390,N_2976,N_2967);
or UO_391 (O_391,N_2992,N_2999);
and UO_392 (O_392,N_2989,N_2996);
nor UO_393 (O_393,N_2955,N_2998);
or UO_394 (O_394,N_2991,N_2960);
nand UO_395 (O_395,N_2999,N_2975);
and UO_396 (O_396,N_2969,N_2970);
nor UO_397 (O_397,N_2981,N_2990);
and UO_398 (O_398,N_2994,N_2980);
or UO_399 (O_399,N_2982,N_2968);
nor UO_400 (O_400,N_2997,N_2962);
nor UO_401 (O_401,N_2998,N_2987);
and UO_402 (O_402,N_2973,N_2977);
xnor UO_403 (O_403,N_2994,N_2995);
nand UO_404 (O_404,N_2962,N_2969);
and UO_405 (O_405,N_2955,N_2950);
or UO_406 (O_406,N_2991,N_2992);
and UO_407 (O_407,N_2966,N_2984);
or UO_408 (O_408,N_2957,N_2972);
or UO_409 (O_409,N_2965,N_2982);
and UO_410 (O_410,N_2988,N_2975);
and UO_411 (O_411,N_2955,N_2966);
xor UO_412 (O_412,N_2965,N_2990);
or UO_413 (O_413,N_2975,N_2968);
and UO_414 (O_414,N_2971,N_2961);
nand UO_415 (O_415,N_2973,N_2987);
nand UO_416 (O_416,N_2983,N_2981);
nand UO_417 (O_417,N_2952,N_2966);
and UO_418 (O_418,N_2952,N_2984);
and UO_419 (O_419,N_2985,N_2950);
nand UO_420 (O_420,N_2958,N_2953);
nand UO_421 (O_421,N_2972,N_2979);
or UO_422 (O_422,N_2970,N_2991);
or UO_423 (O_423,N_2973,N_2968);
nor UO_424 (O_424,N_2990,N_2979);
xnor UO_425 (O_425,N_2961,N_2972);
and UO_426 (O_426,N_2959,N_2977);
or UO_427 (O_427,N_2975,N_2952);
nor UO_428 (O_428,N_2999,N_2963);
and UO_429 (O_429,N_2953,N_2982);
or UO_430 (O_430,N_2957,N_2985);
xnor UO_431 (O_431,N_2982,N_2961);
nand UO_432 (O_432,N_2967,N_2963);
nor UO_433 (O_433,N_2956,N_2996);
nor UO_434 (O_434,N_2973,N_2964);
and UO_435 (O_435,N_2996,N_2982);
and UO_436 (O_436,N_2980,N_2970);
or UO_437 (O_437,N_2990,N_2986);
or UO_438 (O_438,N_2992,N_2984);
and UO_439 (O_439,N_2969,N_2960);
nor UO_440 (O_440,N_2969,N_2985);
and UO_441 (O_441,N_2955,N_2992);
nor UO_442 (O_442,N_2978,N_2996);
or UO_443 (O_443,N_2968,N_2954);
nor UO_444 (O_444,N_2964,N_2953);
nand UO_445 (O_445,N_2982,N_2980);
or UO_446 (O_446,N_2984,N_2950);
and UO_447 (O_447,N_2966,N_2983);
nand UO_448 (O_448,N_2994,N_2982);
and UO_449 (O_449,N_2998,N_2975);
and UO_450 (O_450,N_2988,N_2977);
nor UO_451 (O_451,N_2973,N_2975);
nand UO_452 (O_452,N_2979,N_2954);
and UO_453 (O_453,N_2979,N_2965);
and UO_454 (O_454,N_2950,N_2997);
or UO_455 (O_455,N_2994,N_2969);
nor UO_456 (O_456,N_2956,N_2966);
or UO_457 (O_457,N_2973,N_2961);
nor UO_458 (O_458,N_2995,N_2971);
nand UO_459 (O_459,N_2983,N_2965);
or UO_460 (O_460,N_2973,N_2963);
or UO_461 (O_461,N_2987,N_2971);
nor UO_462 (O_462,N_2961,N_2997);
and UO_463 (O_463,N_2952,N_2963);
nor UO_464 (O_464,N_2959,N_2950);
and UO_465 (O_465,N_2963,N_2981);
or UO_466 (O_466,N_2964,N_2960);
and UO_467 (O_467,N_2975,N_2957);
and UO_468 (O_468,N_2958,N_2961);
nor UO_469 (O_469,N_2965,N_2960);
nor UO_470 (O_470,N_2984,N_2971);
or UO_471 (O_471,N_2961,N_2965);
nand UO_472 (O_472,N_2967,N_2981);
nand UO_473 (O_473,N_2954,N_2990);
and UO_474 (O_474,N_2979,N_2985);
nor UO_475 (O_475,N_2988,N_2955);
and UO_476 (O_476,N_2977,N_2991);
nand UO_477 (O_477,N_2998,N_2997);
or UO_478 (O_478,N_2959,N_2964);
nand UO_479 (O_479,N_2996,N_2964);
nand UO_480 (O_480,N_2964,N_2951);
xnor UO_481 (O_481,N_2979,N_2980);
and UO_482 (O_482,N_2997,N_2987);
or UO_483 (O_483,N_2976,N_2968);
and UO_484 (O_484,N_2967,N_2980);
nand UO_485 (O_485,N_2974,N_2971);
nor UO_486 (O_486,N_2964,N_2956);
and UO_487 (O_487,N_2997,N_2983);
nand UO_488 (O_488,N_2986,N_2982);
and UO_489 (O_489,N_2978,N_2957);
nor UO_490 (O_490,N_2952,N_2973);
nand UO_491 (O_491,N_2965,N_2964);
nand UO_492 (O_492,N_2971,N_2978);
nand UO_493 (O_493,N_2987,N_2964);
and UO_494 (O_494,N_2977,N_2955);
and UO_495 (O_495,N_2990,N_2993);
nand UO_496 (O_496,N_2977,N_2990);
nor UO_497 (O_497,N_2997,N_2966);
and UO_498 (O_498,N_2964,N_2958);
nor UO_499 (O_499,N_2996,N_2972);
endmodule