module basic_2000_20000_2500_40_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1561,In_1360);
xor U1 (N_1,In_321,In_310);
xnor U2 (N_2,In_37,In_1684);
xor U3 (N_3,In_1349,In_290);
nand U4 (N_4,In_1955,In_627);
xnor U5 (N_5,In_1789,In_1695);
nand U6 (N_6,In_212,In_860);
nand U7 (N_7,In_840,In_2);
and U8 (N_8,In_36,In_945);
and U9 (N_9,In_560,In_691);
xnor U10 (N_10,In_721,In_1138);
nor U11 (N_11,In_1599,In_1831);
nor U12 (N_12,In_1612,In_81);
xor U13 (N_13,In_984,In_548);
nand U14 (N_14,In_423,In_1072);
nand U15 (N_15,In_314,In_16);
nor U16 (N_16,In_1067,In_1980);
and U17 (N_17,In_1914,In_131);
and U18 (N_18,In_20,In_1832);
nand U19 (N_19,In_800,In_857);
and U20 (N_20,In_694,In_1711);
nor U21 (N_21,In_951,In_146);
nand U22 (N_22,In_1492,In_1194);
nand U23 (N_23,In_514,In_655);
nor U24 (N_24,In_1763,In_718);
or U25 (N_25,In_1025,In_1503);
xor U26 (N_26,In_26,In_1127);
or U27 (N_27,In_1402,In_1493);
and U28 (N_28,In_1873,In_923);
and U29 (N_29,In_412,In_1875);
and U30 (N_30,In_111,In_1165);
nand U31 (N_31,In_1741,In_1309);
nor U32 (N_32,In_159,In_1097);
or U33 (N_33,In_1911,In_303);
and U34 (N_34,In_316,In_1488);
or U35 (N_35,In_1233,In_824);
nand U36 (N_36,In_1334,In_736);
or U37 (N_37,In_397,In_877);
nand U38 (N_38,In_209,In_830);
nand U39 (N_39,In_93,In_1180);
and U40 (N_40,In_917,In_1634);
or U41 (N_41,In_664,In_1191);
xnor U42 (N_42,In_1927,In_1463);
xor U43 (N_43,In_5,In_165);
xor U44 (N_44,In_1753,In_661);
nor U45 (N_45,In_138,In_1514);
or U46 (N_46,In_1703,In_167);
or U47 (N_47,In_1778,In_1727);
nand U48 (N_48,In_1132,In_1827);
or U49 (N_49,In_734,In_1659);
xor U50 (N_50,In_818,In_1251);
and U51 (N_51,In_853,In_1845);
and U52 (N_52,In_304,In_1237);
or U53 (N_53,In_704,In_1800);
and U54 (N_54,In_1079,In_1013);
xor U55 (N_55,In_660,In_1143);
xnor U56 (N_56,In_1805,In_119);
and U57 (N_57,In_953,In_667);
nor U58 (N_58,In_267,In_1175);
nor U59 (N_59,In_7,In_297);
nand U60 (N_60,In_162,In_774);
nor U61 (N_61,In_1031,In_1618);
nor U62 (N_62,In_21,In_298);
xor U63 (N_63,In_935,In_1972);
nor U64 (N_64,In_1449,In_139);
and U65 (N_65,In_849,In_963);
nand U66 (N_66,In_404,In_1699);
xnor U67 (N_67,In_1498,In_788);
nor U68 (N_68,In_508,In_1395);
xor U69 (N_69,In_1048,In_712);
and U70 (N_70,In_1663,In_1055);
xnor U71 (N_71,In_442,In_1584);
nor U72 (N_72,In_253,In_772);
nor U73 (N_73,In_1565,In_1650);
nor U74 (N_74,In_907,In_931);
nor U75 (N_75,In_1316,In_556);
or U76 (N_76,In_1234,In_1253);
and U77 (N_77,In_176,In_595);
xnor U78 (N_78,In_601,In_597);
xor U79 (N_79,In_66,In_1276);
nand U80 (N_80,In_1003,In_129);
and U81 (N_81,In_549,In_965);
or U82 (N_82,In_605,In_743);
nand U83 (N_83,In_491,In_1485);
or U84 (N_84,In_1456,In_1796);
nor U85 (N_85,In_1706,In_161);
xnor U86 (N_86,In_588,In_859);
nand U87 (N_87,In_783,In_1883);
xor U88 (N_88,In_1662,In_1523);
nor U89 (N_89,In_551,In_753);
nor U90 (N_90,In_1720,In_637);
nand U91 (N_91,In_1280,In_152);
and U92 (N_92,In_1962,In_465);
nor U93 (N_93,In_1836,In_1841);
nand U94 (N_94,In_1902,In_1405);
and U95 (N_95,In_1022,In_1975);
xnor U96 (N_96,In_1500,In_172);
nor U97 (N_97,In_416,In_1495);
nand U98 (N_98,In_103,In_1869);
nand U99 (N_99,In_1231,In_424);
nand U100 (N_100,In_510,In_532);
xnor U101 (N_101,In_1023,In_911);
xnor U102 (N_102,In_1169,In_1390);
and U103 (N_103,In_594,In_977);
xor U104 (N_104,In_775,In_1772);
or U105 (N_105,In_14,In_1524);
nor U106 (N_106,In_150,In_750);
or U107 (N_107,In_1757,In_1118);
and U108 (N_108,In_1707,In_1243);
xor U109 (N_109,In_83,In_194);
xnor U110 (N_110,In_1462,In_130);
and U111 (N_111,In_1846,In_794);
or U112 (N_112,In_418,In_242);
or U113 (N_113,In_1196,In_1440);
or U114 (N_114,In_1080,In_102);
nor U115 (N_115,In_805,In_67);
and U116 (N_116,In_1547,In_156);
nand U117 (N_117,In_1855,In_99);
xor U118 (N_118,In_522,In_703);
and U119 (N_119,In_1105,In_1822);
nor U120 (N_120,In_558,In_887);
nand U121 (N_121,In_1446,In_199);
nand U122 (N_122,In_1812,In_1859);
and U123 (N_123,In_912,In_1054);
or U124 (N_124,In_1035,In_1701);
nor U125 (N_125,In_1550,In_419);
nand U126 (N_126,In_1636,In_1630);
nor U127 (N_127,In_612,In_447);
and U128 (N_128,In_1956,In_1521);
and U129 (N_129,In_389,In_732);
nor U130 (N_130,In_1810,In_92);
xor U131 (N_131,In_838,In_1781);
or U132 (N_132,In_1502,In_757);
xnor U133 (N_133,In_229,In_1037);
nand U134 (N_134,In_1867,In_680);
nand U135 (N_135,In_407,In_482);
nor U136 (N_136,In_968,In_399);
nor U137 (N_137,In_969,In_751);
xnor U138 (N_138,In_1329,In_127);
nand U139 (N_139,In_972,In_237);
xor U140 (N_140,In_647,In_1549);
nand U141 (N_141,In_1490,In_1623);
nor U142 (N_142,In_1677,In_1724);
or U143 (N_143,In_1043,In_1120);
nand U144 (N_144,In_262,In_436);
or U145 (N_145,In_967,In_1219);
xor U146 (N_146,In_120,In_433);
xnor U147 (N_147,In_1217,In_367);
nand U148 (N_148,In_484,In_1819);
nor U149 (N_149,In_3,In_1399);
nand U150 (N_150,In_1115,In_1526);
xor U151 (N_151,In_1155,In_1259);
nor U152 (N_152,In_188,In_631);
or U153 (N_153,In_185,In_485);
or U154 (N_154,In_844,In_51);
nor U155 (N_155,In_1814,In_638);
nand U156 (N_156,In_1984,In_198);
nand U157 (N_157,In_35,In_468);
or U158 (N_158,In_994,In_1445);
nor U159 (N_159,In_983,In_1570);
xnor U160 (N_160,In_1858,In_1793);
or U161 (N_161,In_1751,In_1953);
nor U162 (N_162,In_1900,In_1575);
nor U163 (N_163,In_155,In_797);
and U164 (N_164,In_1664,In_697);
or U165 (N_165,In_625,In_1702);
xor U166 (N_166,In_1389,In_1158);
nand U167 (N_167,In_219,In_1596);
nor U168 (N_168,In_707,In_1327);
nor U169 (N_169,In_490,In_1014);
or U170 (N_170,In_1690,In_939);
or U171 (N_171,In_1294,In_1070);
nor U172 (N_172,In_279,In_1947);
nor U173 (N_173,In_1693,In_24);
nor U174 (N_174,In_1685,In_1619);
nand U175 (N_175,In_1000,In_975);
and U176 (N_176,In_184,In_1254);
nand U177 (N_177,In_1649,In_1917);
and U178 (N_178,In_1366,In_265);
nor U179 (N_179,In_791,In_591);
xor U180 (N_180,In_1718,In_1834);
or U181 (N_181,In_144,In_101);
nor U182 (N_182,In_620,In_294);
and U183 (N_183,In_1053,In_415);
nor U184 (N_184,In_825,In_344);
xnor U185 (N_185,In_1675,In_763);
xnor U186 (N_186,In_1150,In_1933);
or U187 (N_187,In_1744,In_879);
and U188 (N_188,In_133,In_1313);
xnor U189 (N_189,In_782,In_534);
nand U190 (N_190,In_1046,In_1183);
nor U191 (N_191,In_1430,In_677);
or U192 (N_192,In_828,In_280);
xnor U193 (N_193,In_910,In_1246);
nor U194 (N_194,In_47,In_1790);
nand U195 (N_195,In_200,In_890);
or U196 (N_196,In_1944,In_1729);
and U197 (N_197,In_706,In_1347);
nor U198 (N_198,In_545,In_1588);
or U199 (N_199,In_1333,In_1019);
and U200 (N_200,In_44,In_1892);
or U201 (N_201,In_322,In_220);
nor U202 (N_202,In_635,In_11);
xnor U203 (N_203,In_1177,In_143);
nor U204 (N_204,In_1226,In_475);
or U205 (N_205,In_312,In_479);
or U206 (N_206,In_296,In_1129);
or U207 (N_207,In_1296,In_640);
xnor U208 (N_208,In_868,In_110);
xor U209 (N_209,In_674,In_1350);
nor U210 (N_210,In_405,In_429);
nand U211 (N_211,In_538,In_4);
nand U212 (N_212,In_642,In_271);
and U213 (N_213,In_1197,In_1843);
nand U214 (N_214,In_875,In_192);
or U215 (N_215,In_976,In_1726);
xor U216 (N_216,In_1406,In_223);
and U217 (N_217,In_684,In_1218);
or U218 (N_218,In_1027,In_1378);
and U219 (N_219,In_173,In_896);
or U220 (N_220,In_1899,In_793);
xnor U221 (N_221,In_1365,In_1563);
or U222 (N_222,In_347,In_1416);
and U223 (N_223,In_957,In_1799);
xor U224 (N_224,In_858,In_1420);
xor U225 (N_225,In_1239,In_996);
nand U226 (N_226,In_96,In_1908);
nand U227 (N_227,In_1172,In_1638);
nor U228 (N_228,In_100,In_537);
nor U229 (N_229,In_472,In_1182);
xor U230 (N_230,In_600,In_1890);
or U231 (N_231,In_1973,In_1766);
and U232 (N_232,In_1787,In_1431);
xnor U233 (N_233,In_523,In_134);
nor U234 (N_234,In_752,In_61);
nand U235 (N_235,In_1056,In_460);
and U236 (N_236,In_1939,In_1881);
xnor U237 (N_237,In_123,In_593);
and U238 (N_238,In_1759,In_668);
nand U239 (N_239,In_478,In_819);
nand U240 (N_240,In_1093,In_767);
and U241 (N_241,In_1278,In_43);
and U242 (N_242,In_852,In_1489);
nand U243 (N_243,In_390,In_724);
xnor U244 (N_244,In_1530,In_1216);
and U245 (N_245,In_621,In_941);
xnor U246 (N_246,In_284,In_1696);
nand U247 (N_247,In_837,In_784);
and U248 (N_248,In_1994,In_1011);
nand U249 (N_249,In_1756,In_289);
xor U250 (N_250,In_876,In_1566);
or U251 (N_251,In_1142,In_1971);
or U252 (N_252,In_1808,In_731);
or U253 (N_253,In_1016,In_533);
or U254 (N_254,In_1464,In_609);
nor U255 (N_255,In_1008,In_973);
or U256 (N_256,In_688,In_74);
and U257 (N_257,In_1300,In_1587);
xor U258 (N_258,In_934,In_228);
nand U259 (N_259,In_392,In_1354);
nand U260 (N_260,In_745,In_550);
nor U261 (N_261,In_1725,In_417);
nand U262 (N_262,In_1614,In_581);
and U263 (N_263,In_903,In_1106);
nand U264 (N_264,In_1052,In_1247);
or U265 (N_265,In_603,In_1797);
and U266 (N_266,In_216,In_1136);
nor U267 (N_267,In_248,In_1862);
and U268 (N_268,In_1730,In_831);
xnor U269 (N_269,In_1765,In_1714);
xnor U270 (N_270,In_1660,In_956);
or U271 (N_271,In_554,In_1768);
or U272 (N_272,In_933,In_98);
xnor U273 (N_273,In_1291,In_1077);
xor U274 (N_274,In_596,In_68);
or U275 (N_275,In_323,In_1227);
or U276 (N_276,In_572,In_374);
and U277 (N_277,In_473,In_300);
xor U278 (N_278,In_1,In_1211);
nor U279 (N_279,In_1511,In_608);
and U280 (N_280,In_94,In_1328);
and U281 (N_281,In_512,In_1471);
xor U282 (N_282,In_1673,In_1117);
nand U283 (N_283,In_273,In_1382);
nor U284 (N_284,In_702,In_1178);
xor U285 (N_285,In_1905,In_249);
and U286 (N_286,In_1857,In_204);
nand U287 (N_287,In_1128,In_1020);
nand U288 (N_288,In_1779,In_1880);
nand U289 (N_289,In_1400,In_201);
or U290 (N_290,In_1746,In_1861);
nand U291 (N_291,In_1769,In_808);
or U292 (N_292,In_489,In_1361);
xnor U293 (N_293,In_1422,In_370);
or U294 (N_294,In_483,In_1397);
and U295 (N_295,In_206,In_886);
nor U296 (N_296,In_1181,In_974);
nand U297 (N_297,In_1784,In_78);
nor U298 (N_298,In_387,In_1308);
nor U299 (N_299,In_1341,In_1223);
and U300 (N_300,In_1731,In_1174);
nand U301 (N_301,In_1222,In_1686);
xnor U302 (N_302,In_1583,In_364);
and U303 (N_303,In_1543,In_922);
and U304 (N_304,In_1921,In_286);
and U305 (N_305,In_1340,In_1412);
or U306 (N_306,In_1713,In_1894);
nand U307 (N_307,In_1209,In_187);
and U308 (N_308,In_464,In_717);
and U309 (N_309,In_1670,In_1557);
or U310 (N_310,In_451,In_1930);
xor U311 (N_311,In_234,In_881);
or U312 (N_312,In_613,In_1356);
nor U313 (N_313,In_589,In_1267);
nand U314 (N_314,In_1041,In_1210);
and U315 (N_315,In_1315,In_1998);
and U316 (N_316,In_1518,In_30);
nand U317 (N_317,In_1922,In_1184);
and U318 (N_318,In_1337,In_336);
xnor U319 (N_319,In_1667,In_1376);
or U320 (N_320,In_820,In_145);
nor U321 (N_321,In_1585,In_1133);
and U322 (N_322,In_672,In_126);
or U323 (N_323,In_1479,In_1644);
and U324 (N_324,In_564,In_832);
and U325 (N_325,In_573,In_1418);
xnor U326 (N_326,In_1042,In_1652);
nor U327 (N_327,In_1324,In_811);
or U328 (N_328,In_88,In_870);
and U329 (N_329,In_1472,In_1373);
nand U330 (N_330,In_463,In_15);
and U331 (N_331,In_924,In_946);
xnor U332 (N_332,In_64,In_319);
nand U333 (N_333,In_1934,In_1611);
xnor U334 (N_334,In_1487,In_263);
xnor U335 (N_335,In_737,In_710);
xor U336 (N_336,In_714,In_656);
nor U337 (N_337,In_227,In_1438);
nor U338 (N_338,In_1582,In_644);
and U339 (N_339,In_1275,In_1051);
or U340 (N_340,In_378,In_458);
or U341 (N_341,In_563,In_1249);
nor U342 (N_342,In_1950,In_892);
xor U343 (N_343,In_353,In_1806);
xnor U344 (N_344,In_1739,In_85);
nand U345 (N_345,In_108,In_1461);
or U346 (N_346,In_444,In_799);
or U347 (N_347,In_217,In_170);
and U348 (N_348,In_252,In_1568);
nand U349 (N_349,In_1504,In_708);
nor U350 (N_350,In_1826,In_1606);
nand U351 (N_351,In_1958,In_769);
nor U352 (N_352,In_520,In_1352);
xor U353 (N_353,In_1413,In_295);
nor U354 (N_354,In_1964,In_401);
and U355 (N_355,In_1656,In_1874);
and U356 (N_356,In_1468,In_542);
xor U357 (N_357,In_1617,In_1928);
xnor U358 (N_358,In_1310,In_1853);
nor U359 (N_359,In_735,In_238);
nand U360 (N_360,In_1141,In_1126);
and U361 (N_361,In_115,In_106);
xnor U362 (N_362,In_1532,In_1111);
nand U363 (N_363,In_606,In_873);
nand U364 (N_364,In_954,In_231);
or U365 (N_365,In_1920,In_59);
nor U366 (N_366,In_1122,In_1533);
nor U367 (N_367,In_1512,In_1095);
xor U368 (N_368,In_157,In_1897);
nand U369 (N_369,In_553,In_42);
or U370 (N_370,In_362,In_69);
nor U371 (N_371,In_823,In_1103);
or U372 (N_372,In_104,In_1546);
or U373 (N_373,In_1989,In_1666);
nor U374 (N_374,In_676,In_789);
or U375 (N_375,In_1909,In_1379);
nor U376 (N_376,In_1336,In_1137);
or U377 (N_377,In_363,In_1669);
nand U378 (N_378,In_584,In_1392);
and U379 (N_379,In_938,In_125);
xnor U380 (N_380,In_889,In_440);
nor U381 (N_381,In_128,In_1081);
and U382 (N_382,In_1534,In_1633);
and U383 (N_383,In_1467,In_1854);
nor U384 (N_384,In_1363,In_1483);
nand U385 (N_385,In_778,In_1435);
nand U386 (N_386,In_632,In_1362);
or U387 (N_387,In_1168,In_693);
nor U388 (N_388,In_1820,In_1491);
nor U389 (N_389,In_926,In_663);
and U390 (N_390,In_835,In_1966);
and U391 (N_391,In_1576,In_1065);
nor U392 (N_392,In_862,In_1952);
or U393 (N_393,In_1864,In_41);
or U394 (N_394,In_1268,In_222);
and U395 (N_395,In_1086,In_31);
and U396 (N_396,In_985,In_864);
xor U397 (N_397,In_1213,In_1108);
xnor U398 (N_398,In_1396,In_998);
nand U399 (N_399,In_86,In_777);
and U400 (N_400,In_48,In_654);
nand U401 (N_401,In_1629,In_536);
and U402 (N_402,In_507,In_515);
nor U403 (N_403,In_662,In_254);
xor U404 (N_404,In_908,In_383);
xor U405 (N_405,In_1551,In_180);
nand U406 (N_406,In_1214,In_1015);
and U407 (N_407,In_1740,In_1887);
or U408 (N_408,In_193,In_1076);
nor U409 (N_409,In_225,In_1424);
and U410 (N_410,In_50,In_181);
nor U411 (N_411,In_19,In_1654);
xor U412 (N_412,In_277,In_1466);
nor U413 (N_413,In_1750,In_571);
nor U414 (N_414,In_919,In_274);
nand U415 (N_415,In_1320,In_275);
and U416 (N_416,In_1256,In_1426);
or U417 (N_417,In_80,In_1087);
nor U418 (N_418,In_264,In_689);
or U419 (N_419,In_871,In_513);
and U420 (N_420,In_409,In_333);
and U421 (N_421,In_1645,In_1199);
xnor U422 (N_422,In_1453,In_117);
or U423 (N_423,In_1647,In_1786);
and U424 (N_424,In_1804,In_995);
and U425 (N_425,In_645,In_906);
nor U426 (N_426,In_798,In_1559);
and U427 (N_427,In_1680,In_1536);
or U428 (N_428,In_679,In_324);
and U429 (N_429,In_982,In_1553);
nor U430 (N_430,In_1538,In_1288);
xor U431 (N_431,In_255,In_178);
nand U432 (N_432,In_1865,In_1469);
or U433 (N_433,In_1539,In_334);
xnor U434 (N_434,In_1620,In_239);
xor U435 (N_435,In_400,In_1032);
nand U436 (N_436,In_1509,In_813);
nor U437 (N_437,In_1807,In_135);
or U438 (N_438,In_205,In_773);
or U439 (N_439,In_1613,In_1476);
nand U440 (N_440,In_1135,In_659);
nor U441 (N_441,In_1595,In_719);
nor U442 (N_442,In_1096,In_337);
xor U443 (N_443,In_208,In_1295);
nor U444 (N_444,In_874,In_1977);
nor U445 (N_445,In_46,In_1066);
nand U446 (N_446,In_1358,In_1732);
or U447 (N_447,In_1242,In_1432);
and U448 (N_448,In_1357,In_163);
and U449 (N_449,In_854,In_1527);
xnor U450 (N_450,In_283,In_1372);
nor U451 (N_451,In_577,In_505);
or U452 (N_452,In_1991,In_1157);
nor U453 (N_453,In_516,In_1683);
nand U454 (N_454,In_1282,In_1788);
nand U455 (N_455,In_950,In_320);
and U456 (N_456,In_244,In_82);
nor U457 (N_457,In_1038,In_1215);
xor U458 (N_458,In_1529,In_1228);
and U459 (N_459,In_1326,In_827);
nand U460 (N_460,In_1236,In_1889);
nand U461 (N_461,In_299,In_755);
or U462 (N_462,In_1036,In_1837);
xor U463 (N_463,In_1995,In_268);
nand U464 (N_464,In_413,In_1640);
or U465 (N_465,In_1069,In_1303);
and U466 (N_466,In_1156,In_1331);
nor U467 (N_467,In_459,In_87);
or U468 (N_468,In_118,In_602);
xnor U469 (N_469,In_1009,In_1496);
and U470 (N_470,In_372,In_107);
nor U471 (N_471,In_1260,In_937);
and U472 (N_472,In_151,In_326);
nor U473 (N_473,In_278,In_301);
nor U474 (N_474,In_1580,In_803);
xnor U475 (N_475,In_214,In_1153);
nand U476 (N_476,In_1754,In_1562);
nor U477 (N_477,In_709,In_865);
xor U478 (N_478,In_1879,In_1104);
and U479 (N_479,In_618,In_1969);
xnor U480 (N_480,In_492,In_1383);
xor U481 (N_481,In_1411,In_959);
nor U482 (N_482,In_23,In_1764);
or U483 (N_483,In_1965,In_1205);
nand U484 (N_484,In_1474,In_701);
xor U485 (N_485,In_1311,In_361);
nor U486 (N_486,In_179,In_1747);
xnor U487 (N_487,In_1918,In_1335);
xor U488 (N_488,In_1007,In_113);
xnor U489 (N_489,In_756,In_421);
nor U490 (N_490,In_1948,In_742);
or U491 (N_491,In_1925,In_302);
nand U492 (N_492,In_1044,In_1099);
and U493 (N_493,In_1915,In_943);
or U494 (N_494,In_1075,In_1497);
and U495 (N_495,In_928,In_681);
nand U496 (N_496,In_1398,In_705);
nor U497 (N_497,In_431,In_95);
nor U498 (N_498,In_952,In_1004);
xnor U499 (N_499,In_1791,In_257);
or U500 (N_500,In_929,In_958);
xnor U501 (N_501,N_21,In_884);
and U502 (N_502,In_1970,In_1144);
nor U503 (N_503,In_1263,In_738);
and U504 (N_504,In_575,In_970);
and U505 (N_505,In_1064,In_1798);
nor U506 (N_506,In_883,In_746);
or U507 (N_507,In_1101,In_455);
and U508 (N_508,N_345,In_1368);
or U509 (N_509,N_486,In_1317);
or U510 (N_510,In_1151,In_369);
nand U511 (N_511,In_368,N_377);
nor U512 (N_512,In_358,N_67);
xor U513 (N_513,In_1710,In_845);
nor U514 (N_514,In_683,In_1513);
nand U515 (N_515,N_494,In_899);
and U516 (N_516,In_1269,In_1114);
nor U517 (N_517,In_535,N_7);
and U518 (N_518,In_927,N_406);
or U519 (N_519,In_1480,In_1868);
or U520 (N_520,In_1351,N_94);
and U521 (N_521,In_1201,N_299);
or U522 (N_522,In_1113,N_147);
nand U523 (N_523,N_317,In_685);
nand U524 (N_524,N_2,In_759);
nor U525 (N_525,In_453,In_498);
nand U526 (N_526,In_1499,In_1615);
xnor U527 (N_527,In_1342,In_944);
nor U528 (N_528,In_1451,In_467);
nor U529 (N_529,In_771,In_1802);
nand U530 (N_530,N_87,In_916);
nor U531 (N_531,In_1084,In_411);
nand U532 (N_532,N_327,In_169);
nand U533 (N_533,N_123,In_812);
nor U534 (N_534,In_307,In_1851);
and U535 (N_535,In_197,In_586);
xor U536 (N_536,In_1045,In_1162);
and U537 (N_537,N_476,N_106);
xnor U538 (N_538,In_790,In_241);
xor U539 (N_539,In_670,N_71);
xnor U540 (N_540,In_897,In_1220);
nand U541 (N_541,In_1318,N_222);
nand U542 (N_542,In_191,N_474);
or U543 (N_543,N_463,In_1678);
xnor U544 (N_544,In_28,In_1258);
and U545 (N_545,In_1439,N_75);
nand U546 (N_546,In_1203,N_172);
xor U547 (N_547,N_173,In_91);
nand U548 (N_548,In_1062,In_1367);
nand U549 (N_549,In_999,In_1364);
nor U550 (N_550,N_42,N_111);
xor U551 (N_551,N_200,N_235);
and U552 (N_552,In_1888,In_885);
xnor U553 (N_553,In_733,In_166);
xnor U554 (N_554,In_377,N_52);
or U555 (N_555,In_1185,N_467);
and U556 (N_556,In_1658,N_359);
xor U557 (N_557,In_822,In_1555);
and U558 (N_558,N_294,In_250);
nand U559 (N_559,In_948,In_531);
nor U560 (N_560,In_1444,In_1255);
and U561 (N_561,N_128,N_49);
nand U562 (N_562,In_1830,N_321);
nor U563 (N_563,In_1829,N_229);
xnor U564 (N_564,In_408,In_1906);
xor U565 (N_565,In_1261,In_315);
xor U566 (N_566,In_1895,In_240);
and U567 (N_567,N_447,In_1094);
nor U568 (N_568,In_1592,N_399);
nand U569 (N_569,In_470,N_74);
nand U570 (N_570,In_1083,In_1370);
xor U571 (N_571,N_247,In_1154);
and U572 (N_572,In_1293,N_325);
or U573 (N_573,N_356,In_700);
or U574 (N_574,In_1385,In_77);
nand U575 (N_575,In_1943,In_391);
xor U576 (N_576,In_658,In_848);
or U577 (N_577,In_340,N_369);
and U578 (N_578,N_141,In_1737);
and U579 (N_579,In_1605,N_307);
and U580 (N_580,N_459,In_149);
or U581 (N_581,N_300,In_1591);
nor U582 (N_582,In_1441,N_471);
and U583 (N_583,N_304,In_611);
xor U584 (N_584,N_113,In_1520);
xor U585 (N_585,In_282,In_814);
xor U586 (N_586,In_1782,In_726);
xnor U587 (N_587,N_152,N_298);
nand U588 (N_588,N_216,N_446);
nand U589 (N_589,N_202,In_1494);
xor U590 (N_590,In_1651,N_341);
or U591 (N_591,In_1200,N_140);
or U592 (N_592,In_687,N_100);
nor U593 (N_593,In_306,In_915);
and U594 (N_594,In_33,In_1119);
nand U595 (N_595,In_530,N_358);
or U596 (N_596,In_947,In_1882);
or U597 (N_597,In_1579,In_1281);
nand U598 (N_598,N_297,In_1381);
or U599 (N_599,In_1507,N_167);
nand U600 (N_600,N_381,N_50);
or U601 (N_601,N_38,In_1192);
nand U602 (N_602,In_1558,N_20);
xnor U603 (N_603,N_194,In_396);
or U604 (N_604,In_566,In_504);
nor U605 (N_605,In_801,In_1728);
nor U606 (N_606,In_1743,N_461);
nand U607 (N_607,N_378,In_1795);
xnor U608 (N_608,In_428,In_880);
xor U609 (N_609,In_1371,In_1377);
and U610 (N_610,N_495,N_204);
or U611 (N_611,In_1265,In_1149);
xor U612 (N_612,In_1353,In_582);
nand U613 (N_613,N_316,N_45);
xnor U614 (N_614,In_607,In_45);
or U615 (N_615,In_587,N_419);
or U616 (N_616,In_359,In_1560);
nand U617 (N_617,In_1427,In_754);
xor U618 (N_618,In_381,In_1332);
nor U619 (N_619,In_331,In_1626);
or U620 (N_620,N_282,N_412);
or U621 (N_621,In_1026,In_1809);
nand U622 (N_622,In_1131,N_363);
nand U623 (N_623,In_1465,In_1608);
xor U624 (N_624,In_1001,In_259);
or U625 (N_625,In_1248,In_1635);
or U626 (N_626,In_1679,N_335);
nor U627 (N_627,In_1091,N_273);
xnor U628 (N_628,In_713,N_291);
or U629 (N_629,In_1709,In_1839);
nor U630 (N_630,In_653,In_1676);
and U631 (N_631,N_295,N_256);
xor U632 (N_632,N_370,In_426);
or U633 (N_633,In_1508,In_38);
or U634 (N_634,In_765,N_488);
nand U635 (N_635,N_360,In_1123);
nor U636 (N_636,In_1976,N_234);
and U637 (N_637,N_92,In_1924);
and U638 (N_638,N_466,In_1590);
xnor U639 (N_639,N_232,In_1452);
nand U640 (N_640,In_511,In_1688);
nand U641 (N_641,In_675,In_1848);
xnor U642 (N_642,In_287,In_1161);
or U643 (N_643,In_1721,In_730);
nor U644 (N_644,In_1904,N_110);
and U645 (N_645,In_872,In_955);
and U646 (N_646,In_1621,In_992);
nor U647 (N_647,In_1668,In_624);
nor U648 (N_648,N_133,N_404);
xnor U649 (N_649,In_1188,N_371);
and U650 (N_650,In_1531,In_1945);
or U651 (N_651,N_483,N_258);
nor U652 (N_652,In_821,In_1871);
nand U653 (N_653,In_1705,In_855);
and U654 (N_654,N_109,In_666);
nand U655 (N_655,In_1940,N_444);
nor U656 (N_656,In_1193,In_174);
or U657 (N_657,In_63,In_648);
and U658 (N_658,In_1903,In_1159);
nand U659 (N_659,In_1545,In_867);
nor U660 (N_660,In_1107,In_445);
or U661 (N_661,In_1033,In_604);
and U662 (N_662,In_1102,N_55);
nand U663 (N_663,N_440,In_75);
or U664 (N_664,In_493,N_153);
nor U665 (N_665,N_445,N_271);
nand U666 (N_666,N_242,In_1999);
and U667 (N_667,In_846,In_1164);
and U668 (N_668,N_190,In_497);
or U669 (N_669,N_171,In_183);
xor U670 (N_670,In_1780,N_398);
or U671 (N_671,In_1816,N_468);
xor U672 (N_672,N_10,In_1985);
and U673 (N_673,In_895,N_238);
and U674 (N_674,N_254,N_246);
or U675 (N_675,In_592,In_964);
and U676 (N_676,In_1322,In_1811);
and U677 (N_677,N_77,In_1946);
and U678 (N_678,In_441,In_70);
nor U679 (N_679,N_449,In_97);
nor U680 (N_680,In_195,In_981);
and U681 (N_681,N_385,N_479);
nor U682 (N_682,In_626,In_1145);
nor U683 (N_683,In_1224,In_1541);
and U684 (N_684,In_1567,N_99);
nand U685 (N_685,N_396,N_146);
xnor U686 (N_686,In_346,N_184);
nand U687 (N_687,In_1116,In_1306);
nand U688 (N_688,In_1996,In_1866);
nand U689 (N_689,In_84,N_187);
nor U690 (N_690,In_1872,In_1574);
and U691 (N_691,In_1535,In_914);
xnor U692 (N_692,In_39,In_501);
xnor U693 (N_693,In_1813,N_186);
or U694 (N_694,In_1773,In_124);
nor U695 (N_695,In_8,N_364);
and U696 (N_696,In_650,N_287);
xor U697 (N_697,In_1134,N_118);
and U698 (N_698,In_1653,In_1957);
or U699 (N_699,In_1604,N_59);
or U700 (N_700,In_1098,In_317);
and U701 (N_701,In_1896,N_251);
xor U702 (N_702,In_9,In_559);
xor U703 (N_703,N_64,In_942);
xnor U704 (N_704,N_414,In_529);
and U705 (N_705,N_95,In_639);
nand U706 (N_706,In_1665,In_1907);
xnor U707 (N_707,N_394,In_1204);
xor U708 (N_708,In_235,N_32);
xor U709 (N_709,In_1671,In_1160);
nand U710 (N_710,In_1936,In_1733);
or U711 (N_711,N_124,In_1586);
xnor U712 (N_712,N_320,In_1029);
xor U713 (N_713,In_1244,In_786);
or U714 (N_714,In_6,In_215);
xnor U715 (N_715,In_1992,N_333);
nor U716 (N_716,In_652,N_272);
and U717 (N_717,N_18,N_410);
nand U718 (N_718,N_154,N_284);
and U719 (N_719,In_1639,In_232);
nor U720 (N_720,N_454,N_125);
nor U721 (N_721,In_1325,In_1844);
xor U722 (N_722,In_555,N_233);
or U723 (N_723,In_863,In_395);
nand U724 (N_724,In_918,N_314);
and U725 (N_725,In_153,In_1556);
xnor U726 (N_726,In_494,In_1384);
nor U727 (N_727,N_155,N_383);
or U728 (N_728,In_539,In_673);
xor U729 (N_729,In_565,In_1012);
nand U730 (N_730,In_1404,N_46);
nand U731 (N_731,N_105,N_386);
nor U732 (N_732,In_1803,In_690);
xor U733 (N_733,In_246,In_1409);
nand U734 (N_734,In_1073,In_1624);
nor U735 (N_735,N_228,In_646);
and U736 (N_736,N_422,In_623);
nor U737 (N_737,In_1825,N_470);
nand U738 (N_738,In_1312,N_192);
and U739 (N_739,In_1522,In_1852);
xnor U740 (N_740,N_16,N_122);
and U741 (N_741,In_506,N_145);
xnor U742 (N_742,In_1021,In_260);
xnor U743 (N_743,N_326,N_208);
or U744 (N_744,In_457,N_337);
nand U745 (N_745,In_1935,N_117);
nor U746 (N_746,N_14,N_17);
nor U747 (N_747,In_682,In_1425);
nor U748 (N_748,In_292,In_839);
and U749 (N_749,In_617,In_1287);
or U750 (N_750,In_1460,In_1092);
nor U751 (N_751,In_452,N_31);
and U752 (N_752,In_1609,N_441);
nand U753 (N_753,N_130,In_990);
nor U754 (N_754,N_243,N_413);
xnor U755 (N_755,In_1993,In_1388);
nand U756 (N_756,In_861,In_1847);
or U757 (N_757,N_478,In_1961);
xnor U758 (N_758,In_1594,In_160);
and U759 (N_759,In_1783,In_393);
and U760 (N_760,N_168,In_761);
xor U761 (N_761,In_1655,In_804);
and U762 (N_762,In_1284,N_306);
and U763 (N_763,N_388,In_1028);
and U764 (N_764,In_1124,N_54);
or U765 (N_765,N_475,In_90);
nand U766 (N_766,N_33,In_1997);
and U767 (N_767,In_816,N_217);
nor U768 (N_768,N_313,In_462);
or U769 (N_769,In_1631,In_1742);
and U770 (N_770,N_1,In_196);
xnor U771 (N_771,In_388,In_925);
nor U772 (N_772,N_451,N_131);
and U773 (N_773,In_671,In_519);
and U774 (N_774,N_357,N_331);
and U775 (N_775,In_481,N_3);
and U776 (N_776,N_149,In_1147);
nor U777 (N_777,In_1661,In_936);
and U778 (N_778,In_308,In_569);
and U779 (N_779,N_91,In_986);
nor U780 (N_780,N_181,In_1171);
nand U781 (N_781,In_1625,In_1304);
or U782 (N_782,In_1774,In_836);
nor U783 (N_783,N_281,N_252);
nand U784 (N_784,In_780,In_1330);
nand U785 (N_785,In_1289,In_1885);
nand U786 (N_786,N_83,In_815);
xnor U787 (N_787,In_1407,N_257);
and U788 (N_788,In_272,In_330);
nand U789 (N_789,N_448,In_1010);
nand U790 (N_790,In_32,In_1482);
xnor U791 (N_791,In_776,N_79);
or U792 (N_792,In_1082,In_1186);
and U793 (N_793,In_1057,In_1931);
nand U794 (N_794,N_23,In_132);
nand U795 (N_795,N_43,N_387);
nor U796 (N_796,N_97,N_85);
nand U797 (N_797,N_215,In_318);
or U798 (N_798,In_1979,N_24);
and U799 (N_799,In_711,N_221);
or U800 (N_800,In_1516,N_457);
nor U801 (N_801,In_1229,N_462);
xnor U802 (N_802,N_157,In_1146);
and U803 (N_803,In_1238,In_991);
or U804 (N_804,N_6,In_1386);
nor U805 (N_805,N_395,N_9);
or U806 (N_806,N_250,In_980);
or U807 (N_807,In_528,In_779);
or U808 (N_808,In_1712,In_795);
or U809 (N_809,In_590,In_949);
nor U810 (N_810,In_438,In_1375);
and U811 (N_811,In_350,In_1893);
or U812 (N_812,In_1849,N_57);
and U813 (N_813,In_500,In_1824);
nor U814 (N_814,In_1305,In_357);
nand U815 (N_815,In_1968,In_379);
nor U816 (N_816,In_1458,In_1190);
nor U817 (N_817,In_1241,In_425);
or U818 (N_818,In_384,In_810);
nor U819 (N_819,N_104,In_723);
xnor U820 (N_820,In_826,N_211);
nor U821 (N_821,In_54,In_1572);
or U822 (N_822,In_1457,N_212);
and U823 (N_823,In_495,N_275);
or U824 (N_824,In_435,N_76);
nor U825 (N_825,N_236,In_562);
nor U826 (N_826,In_1987,In_1682);
nand U827 (N_827,N_391,N_142);
xor U828 (N_828,N_189,In_1719);
nand U829 (N_829,In_1818,N_350);
and U830 (N_830,N_185,In_1273);
nand U831 (N_831,N_39,In_930);
xor U832 (N_832,In_385,N_80);
nor U833 (N_833,In_1459,N_35);
xnor U834 (N_834,N_279,In_437);
nand U835 (N_835,In_557,In_715);
nor U836 (N_836,N_176,In_993);
or U837 (N_837,N_70,N_107);
and U838 (N_838,N_334,N_241);
nor U839 (N_839,In_1090,In_1005);
nor U840 (N_840,N_324,In_747);
xor U841 (N_841,N_311,In_1886);
and U842 (N_842,N_368,N_443);
nand U843 (N_843,In_1913,In_1277);
xor U844 (N_844,N_318,In_190);
and U845 (N_845,In_1109,In_1481);
xor U846 (N_846,N_156,In_1510);
nand U847 (N_847,In_1232,N_159);
nor U848 (N_848,In_1581,In_1369);
xor U849 (N_849,N_151,N_116);
nand U850 (N_850,In_1770,N_48);
nand U851 (N_851,In_741,N_72);
nor U852 (N_852,N_397,N_366);
and U853 (N_853,N_169,In_1923);
nor U854 (N_854,In_233,In_978);
or U855 (N_855,N_480,In_619);
xnor U856 (N_856,In_1736,In_610);
xnor U857 (N_857,In_686,N_180);
and U858 (N_858,In_17,In_291);
nand U859 (N_859,N_438,In_809);
or U860 (N_860,N_90,N_453);
xor U861 (N_861,N_464,In_1982);
or U862 (N_862,N_58,In_1187);
nor U863 (N_863,N_439,N_389);
nand U864 (N_864,In_1433,In_189);
xor U865 (N_865,In_1691,In_1250);
nor U866 (N_866,N_305,N_485);
or U867 (N_867,In_1603,In_833);
xnor U868 (N_868,N_429,N_408);
and U869 (N_869,In_371,N_218);
nor U870 (N_870,In_729,N_96);
and U871 (N_871,In_1775,In_1597);
nand U872 (N_872,In_207,N_426);
and U873 (N_873,N_143,N_259);
or U874 (N_874,In_1910,In_1932);
nor U875 (N_875,In_665,In_1348);
and U876 (N_876,In_882,In_807);
or U877 (N_877,N_68,N_497);
xnor U878 (N_878,In_1173,In_966);
nor U879 (N_879,In_12,In_599);
nand U880 (N_880,In_720,N_384);
nor U881 (N_881,In_524,N_465);
and U882 (N_882,N_231,N_30);
nor U883 (N_883,In_987,In_669);
nand U884 (N_884,N_62,N_409);
xor U885 (N_885,In_1071,In_1024);
or U886 (N_886,N_428,N_417);
xor U887 (N_887,N_424,In_1401);
xnor U888 (N_888,In_829,In_1986);
or U889 (N_889,N_379,In_893);
xor U890 (N_890,In_430,In_1578);
and U891 (N_891,N_8,In_345);
nor U892 (N_892,N_239,In_802);
nor U893 (N_893,In_1298,In_521);
and U894 (N_894,In_725,In_332);
and U895 (N_895,In_434,N_119);
and U896 (N_896,N_205,In_1919);
and U897 (N_897,In_122,N_353);
and U898 (N_898,In_1387,In_456);
or U899 (N_899,N_206,N_73);
and U900 (N_900,In_1285,In_1148);
xor U901 (N_901,In_448,N_245);
nor U902 (N_902,In_394,In_1761);
nand U903 (N_903,In_1642,In_1163);
xor U904 (N_904,In_1271,In_1030);
nor U905 (N_905,In_496,N_193);
or U906 (N_906,In_1898,In_1657);
or U907 (N_907,In_1423,In_247);
and U908 (N_908,In_1410,In_841);
xnor U909 (N_909,In_1794,In_580);
nand U910 (N_910,In_909,In_1593);
nand U911 (N_911,In_1735,In_1486);
xnor U912 (N_912,N_492,In_1959);
nor U913 (N_913,N_88,N_436);
and U914 (N_914,In_1525,In_1941);
xnor U915 (N_915,N_199,In_1152);
nor U916 (N_916,N_489,N_392);
nor U917 (N_917,In_1264,In_1359);
xor U918 (N_918,N_263,In_137);
nand U919 (N_919,N_415,N_351);
nor U920 (N_920,In_1981,In_698);
and U921 (N_921,N_161,N_223);
xor U922 (N_922,N_498,In_1189);
nor U923 (N_923,In_851,N_342);
nand U924 (N_924,In_477,In_450);
and U925 (N_925,In_1600,In_1687);
or U926 (N_926,In_1419,In_141);
or U927 (N_927,In_695,In_888);
nor U928 (N_928,In_932,N_4);
and U929 (N_929,N_127,N_278);
xnor U930 (N_930,N_458,In_1314);
nor U931 (N_931,In_526,In_850);
and U932 (N_932,In_1758,N_213);
nand U933 (N_933,In_1752,In_1415);
or U934 (N_934,In_1002,N_493);
and U935 (N_935,N_121,In_140);
xnor U936 (N_936,In_276,In_1018);
or U937 (N_937,N_13,In_1167);
nor U938 (N_938,In_89,In_1938);
nand U939 (N_939,In_116,In_1876);
or U940 (N_940,N_487,In_1121);
and U941 (N_941,N_214,In_1225);
nand U942 (N_942,In_1506,In_1537);
nor U943 (N_943,In_1681,In_503);
nor U944 (N_944,In_921,In_1715);
and U945 (N_945,In_305,N_244);
nand U946 (N_946,In_920,N_60);
nand U947 (N_947,In_1823,In_1130);
nor U948 (N_948,In_1252,In_1112);
or U949 (N_949,In_1776,In_657);
or U950 (N_950,N_65,N_491);
and U951 (N_951,N_115,In_1540);
xor U952 (N_952,In_643,N_416);
and U953 (N_953,In_834,In_1436);
nor U954 (N_954,In_1179,N_390);
nor U955 (N_955,In_1515,In_335);
nand U956 (N_956,N_219,N_308);
xor U957 (N_957,In_171,N_112);
xnor U958 (N_958,N_139,N_280);
xor U959 (N_959,In_56,In_1878);
nor U960 (N_960,N_303,N_163);
and U961 (N_961,In_1286,N_203);
nor U962 (N_962,In_432,In_1863);
and U963 (N_963,N_290,N_166);
or U964 (N_964,In_474,In_1230);
nor U965 (N_965,In_1891,N_237);
or U966 (N_966,In_71,N_472);
or U967 (N_967,N_477,N_420);
xor U968 (N_968,N_332,In_842);
or U969 (N_969,N_473,N_36);
nand U970 (N_970,In_1085,N_158);
or U971 (N_971,In_1648,N_283);
and U972 (N_972,N_53,In_1916);
nand U973 (N_973,In_22,In_518);
xnor U974 (N_974,In_1937,In_309);
nor U975 (N_975,N_44,In_148);
xor U976 (N_976,N_349,N_136);
and U977 (N_977,In_1272,In_1573);
nor U978 (N_978,In_1745,In_1391);
nand U979 (N_979,In_843,In_1437);
xor U980 (N_980,N_103,N_393);
and U981 (N_981,In_175,In_1674);
nand U982 (N_982,In_1475,N_268);
or U983 (N_983,N_210,In_1929);
and U984 (N_984,N_362,N_11);
or U985 (N_985,N_89,N_255);
nor U986 (N_986,N_336,N_248);
nand U987 (N_987,In_722,In_427);
or U988 (N_988,N_81,In_1589);
or U989 (N_989,N_253,In_1454);
nand U990 (N_990,In_356,In_57);
xor U991 (N_991,N_348,In_1470);
nor U992 (N_992,In_636,In_781);
and U993 (N_993,N_138,N_361);
or U994 (N_994,N_309,In_1176);
xor U995 (N_995,In_509,In_76);
or U996 (N_996,In_1505,In_342);
or U997 (N_997,In_988,In_1345);
nor U998 (N_998,In_1017,In_1061);
or U999 (N_999,In_1125,In_243);
and U1000 (N_1000,N_871,In_1988);
or U1001 (N_1001,In_62,N_867);
nand U1002 (N_1002,N_673,N_702);
and U1003 (N_1003,N_730,In_1616);
nand U1004 (N_1004,N_160,In_365);
and U1005 (N_1005,N_554,In_1738);
nand U1006 (N_1006,N_938,In_598);
and U1007 (N_1007,In_1414,In_678);
nor U1008 (N_1008,N_547,In_410);
nand U1009 (N_1009,In_486,N_963);
nand U1010 (N_1010,N_767,In_406);
nor U1011 (N_1011,N_999,In_869);
and U1012 (N_1012,In_1960,In_1517);
xnor U1013 (N_1013,N_931,N_870);
and U1014 (N_1014,In_1637,N_897);
nand U1015 (N_1015,In_177,In_1235);
nand U1016 (N_1016,In_360,In_1266);
nand U1017 (N_1017,In_1749,N_148);
and U1018 (N_1018,N_879,N_874);
xor U1019 (N_1019,In_1974,N_579);
nand U1020 (N_1020,N_338,In_1835);
or U1021 (N_1021,In_112,In_574);
nand U1022 (N_1022,N_937,N_126);
or U1023 (N_1023,In_114,N_817);
and U1024 (N_1024,In_651,N_319);
or U1025 (N_1025,N_545,In_1564);
nor U1026 (N_1026,N_896,In_1601);
or U1027 (N_1027,N_556,N_323);
nor U1028 (N_1028,In_226,In_1717);
nor U1029 (N_1029,N_909,N_129);
nand U1030 (N_1030,N_716,In_256);
and U1031 (N_1031,N_41,N_700);
nand U1032 (N_1032,In_1297,In_901);
and U1033 (N_1033,In_517,N_812);
nor U1034 (N_1034,In_961,N_536);
nand U1035 (N_1035,N_818,In_328);
or U1036 (N_1036,N_590,In_1059);
and U1037 (N_1037,N_581,N_828);
nand U1038 (N_1038,N_580,N_520);
nand U1039 (N_1039,N_738,N_588);
or U1040 (N_1040,In_1047,N_144);
nand U1041 (N_1041,In_1060,N_552);
or U1042 (N_1042,N_744,N_865);
xnor U1043 (N_1043,N_310,N_854);
and U1044 (N_1044,N_904,In_758);
xor U1045 (N_1045,N_946,N_714);
nor U1046 (N_1046,N_427,In_1068);
nand U1047 (N_1047,In_962,In_142);
nor U1048 (N_1048,N_945,N_407);
or U1049 (N_1049,N_780,N_773);
xor U1050 (N_1050,N_432,N_882);
or U1051 (N_1051,N_919,N_722);
and U1052 (N_1052,N_800,N_548);
nor U1053 (N_1053,In_541,In_52);
and U1054 (N_1054,In_629,N_765);
or U1055 (N_1055,In_218,N_921);
xor U1056 (N_1056,In_1195,N_991);
xor U1057 (N_1057,N_343,N_433);
and U1058 (N_1058,N_659,N_733);
xnor U1059 (N_1059,In_785,N_549);
and U1060 (N_1060,In_147,N_811);
or U1061 (N_1061,In_1355,N_132);
xnor U1062 (N_1062,In_1704,N_354);
and U1063 (N_1063,In_73,N_881);
nor U1064 (N_1064,N_689,N_748);
xnor U1065 (N_1065,In_480,In_1842);
nand U1066 (N_1066,In_552,N_725);
nand U1067 (N_1067,N_857,N_777);
xnor U1068 (N_1068,N_849,N_989);
nor U1069 (N_1069,N_423,In_634);
nor U1070 (N_1070,N_831,In_1926);
and U1071 (N_1071,In_1760,In_311);
nand U1072 (N_1072,N_532,N_286);
nor U1073 (N_1073,N_610,N_834);
nor U1074 (N_1074,In_900,N_920);
nand U1075 (N_1075,N_365,In_1100);
nand U1076 (N_1076,N_935,N_134);
and U1077 (N_1077,N_972,N_511);
xnor U1078 (N_1078,N_789,N_374);
or U1079 (N_1079,In_578,In_1801);
or U1080 (N_1080,N_966,N_0);
and U1081 (N_1081,N_847,In_1627);
nor U1082 (N_1082,In_281,N_992);
nand U1083 (N_1083,In_1270,In_1777);
nand U1084 (N_1084,N_82,N_675);
or U1085 (N_1085,In_373,N_928);
and U1086 (N_1086,In_1274,In_1078);
and U1087 (N_1087,N_681,In_740);
nand U1088 (N_1088,N_569,In_1443);
or U1089 (N_1089,In_898,N_885);
xnor U1090 (N_1090,In_1110,In_1299);
or U1091 (N_1091,N_652,In_261);
xnor U1092 (N_1092,In_285,In_1448);
nor U1093 (N_1093,N_93,In_1393);
nor U1094 (N_1094,N_860,In_1901);
nor U1095 (N_1095,N_537,N_625);
or U1096 (N_1096,N_616,N_614);
nor U1097 (N_1097,N_763,N_499);
nor U1098 (N_1098,N_913,In_1343);
nand U1099 (N_1099,N_968,In_258);
nor U1100 (N_1100,In_439,In_402);
nand U1101 (N_1101,N_732,In_1963);
or U1102 (N_1102,N_612,In_971);
nand U1103 (N_1103,N_496,N_661);
nor U1104 (N_1104,In_1212,In_58);
xnor U1105 (N_1105,In_1484,N_731);
and U1106 (N_1106,N_724,In_633);
xnor U1107 (N_1107,N_69,N_509);
and U1108 (N_1108,In_1817,N_576);
xor U1109 (N_1109,N_810,N_276);
nor U1110 (N_1110,In_121,N_979);
nand U1111 (N_1111,In_792,In_1049);
nor U1112 (N_1112,N_718,In_692);
nand U1113 (N_1113,In_728,N_982);
nand U1114 (N_1114,N_823,In_866);
nor U1115 (N_1115,N_521,N_289);
nand U1116 (N_1116,In_502,N_795);
or U1117 (N_1117,In_1428,N_633);
or U1118 (N_1118,N_188,In_1339);
nand U1119 (N_1119,In_269,In_1767);
and U1120 (N_1120,In_65,In_1240);
nor U1121 (N_1121,N_709,N_667);
nand U1122 (N_1122,N_842,N_608);
xor U1123 (N_1123,In_1884,In_1528);
or U1124 (N_1124,N_183,In_1856);
nand U1125 (N_1125,In_105,N_749);
and U1126 (N_1126,N_609,In_164);
and U1127 (N_1127,N_905,N_887);
or U1128 (N_1128,In_1628,N_745);
nand U1129 (N_1129,In_1571,N_941);
or U1130 (N_1130,N_740,N_801);
nand U1131 (N_1131,N_692,N_915);
and U1132 (N_1132,In_29,N_840);
nor U1133 (N_1133,In_1140,N_562);
or U1134 (N_1134,N_910,N_403);
or U1135 (N_1135,N_835,N_685);
nand U1136 (N_1136,N_312,In_1006);
and U1137 (N_1137,N_170,N_672);
or U1138 (N_1138,N_568,In_251);
and U1139 (N_1139,In_1840,N_523);
nand U1140 (N_1140,In_1723,N_51);
xor U1141 (N_1141,N_174,N_676);
xnor U1142 (N_1142,N_502,In_1700);
and U1143 (N_1143,N_656,N_515);
nor U1144 (N_1144,In_744,N_197);
nor U1145 (N_1145,N_934,N_756);
and U1146 (N_1146,N_758,N_984);
nor U1147 (N_1147,In_699,N_956);
xor U1148 (N_1148,N_191,In_1821);
nor U1149 (N_1149,N_640,N_655);
nand U1150 (N_1150,In_34,N_890);
nand U1151 (N_1151,N_802,N_240);
xor U1152 (N_1152,N_878,N_844);
nand U1153 (N_1153,N_665,N_622);
or U1154 (N_1154,N_431,In_325);
xor U1155 (N_1155,N_78,In_940);
nand U1156 (N_1156,N_582,N_601);
xnor U1157 (N_1157,N_628,In_1058);
nand U1158 (N_1158,N_892,N_769);
nor U1159 (N_1159,N_737,N_534);
xnor U1160 (N_1160,N_816,N_435);
xnor U1161 (N_1161,In_1734,In_414);
nor U1162 (N_1162,In_136,In_213);
nor U1163 (N_1163,N_691,N_37);
and U1164 (N_1164,N_687,N_807);
nand U1165 (N_1165,In_355,N_944);
or U1166 (N_1166,N_848,In_878);
xor U1167 (N_1167,N_646,N_484);
nor U1168 (N_1168,In_1403,N_629);
nand U1169 (N_1169,N_274,N_997);
and U1170 (N_1170,N_739,N_546);
or U1171 (N_1171,N_843,N_923);
xnor U1172 (N_1172,In_446,N_711);
or U1173 (N_1173,N_803,In_561);
or U1174 (N_1174,N_712,N_522);
nand U1175 (N_1175,In_245,N_619);
nor U1176 (N_1176,N_670,N_933);
or U1177 (N_1177,N_994,In_570);
xor U1178 (N_1178,In_567,N_605);
xnor U1179 (N_1179,N_352,N_539);
nor U1180 (N_1180,In_1374,N_788);
xnor U1181 (N_1181,N_561,In_1542);
xnor U1182 (N_1182,In_1762,N_734);
and U1183 (N_1183,In_1290,In_1323);
or U1184 (N_1184,In_1394,In_1450);
or U1185 (N_1185,In_894,In_1602);
and U1186 (N_1186,In_1912,In_348);
xor U1187 (N_1187,N_551,In_540);
or U1188 (N_1188,N_830,N_5);
nand U1189 (N_1189,N_611,In_1434);
and U1190 (N_1190,In_787,N_804);
xnor U1191 (N_1191,N_296,N_747);
or U1192 (N_1192,N_198,N_367);
nor U1193 (N_1193,In_210,N_859);
or U1194 (N_1194,N_805,N_631);
nor U1195 (N_1195,N_855,In_1577);
nor U1196 (N_1196,N_694,N_851);
nor U1197 (N_1197,N_292,N_821);
and U1198 (N_1198,N_265,N_293);
and U1199 (N_1199,N_861,N_671);
xnor U1200 (N_1200,In_1050,N_372);
xor U1201 (N_1201,In_905,In_904);
nand U1202 (N_1202,N_586,N_482);
xnor U1203 (N_1203,In_1755,In_403);
and U1204 (N_1204,N_544,N_686);
nor U1205 (N_1205,N_627,N_533);
or U1206 (N_1206,In_1170,In_615);
nor U1207 (N_1207,N_602,N_697);
and U1208 (N_1208,N_645,N_706);
nand U1209 (N_1209,In_109,In_1221);
nand U1210 (N_1210,N_693,N_668);
and U1211 (N_1211,N_642,N_653);
xnor U1212 (N_1212,N_952,N_735);
and U1213 (N_1213,In_351,In_1421);
and U1214 (N_1214,N_678,N_512);
nand U1215 (N_1215,N_927,N_922);
xnor U1216 (N_1216,N_641,In_1442);
nor U1217 (N_1217,In_1877,In_168);
xnor U1218 (N_1218,N_723,In_544);
nand U1219 (N_1219,In_1501,N_995);
nand U1220 (N_1220,N_742,In_1279);
or U1221 (N_1221,N_538,N_567);
and U1222 (N_1222,N_541,In_1206);
or U1223 (N_1223,N_376,N_876);
xor U1224 (N_1224,N_637,N_797);
xnor U1225 (N_1225,N_791,N_727);
xor U1226 (N_1226,N_699,N_380);
xor U1227 (N_1227,N_690,N_527);
and U1228 (N_1228,In_1321,N_779);
nor U1229 (N_1229,N_677,N_768);
nor U1230 (N_1230,N_566,In_224);
xor U1231 (N_1231,N_530,N_647);
or U1232 (N_1232,N_707,In_1455);
nand U1233 (N_1233,In_422,In_1207);
xor U1234 (N_1234,N_858,N_964);
xnor U1235 (N_1235,In_1771,N_720);
or U1236 (N_1236,N_974,N_778);
or U1237 (N_1237,N_650,N_965);
xor U1238 (N_1238,In_1063,N_120);
and U1239 (N_1239,N_901,N_674);
and U1240 (N_1240,N_604,N_679);
or U1241 (N_1241,N_418,N_826);
xnor U1242 (N_1242,N_598,N_220);
and U1243 (N_1243,In_1697,N_880);
xnor U1244 (N_1244,N_531,N_618);
xor U1245 (N_1245,N_595,In_25);
or U1246 (N_1246,In_583,In_293);
nand U1247 (N_1247,In_313,N_469);
or U1248 (N_1248,In_547,In_55);
or U1249 (N_1249,In_1978,In_270);
nor U1250 (N_1250,N_102,N_781);
nor U1251 (N_1251,N_759,In_211);
or U1252 (N_1252,N_517,N_943);
xnor U1253 (N_1253,N_939,N_829);
and U1254 (N_1254,N_261,N_315);
or U1255 (N_1255,In_398,N_630);
or U1256 (N_1256,N_907,In_1301);
nand U1257 (N_1257,In_1166,N_277);
or U1258 (N_1258,N_135,N_838);
nand U1259 (N_1259,N_402,In_1622);
or U1260 (N_1260,N_267,N_434);
xnor U1261 (N_1261,In_1672,In_488);
nor U1262 (N_1262,N_755,In_1554);
nor U1263 (N_1263,N_565,N_302);
xor U1264 (N_1264,N_108,N_524);
nor U1265 (N_1265,N_573,N_98);
and U1266 (N_1266,N_721,In_696);
xor U1267 (N_1267,In_1039,N_813);
xor U1268 (N_1268,In_1257,N_620);
or U1269 (N_1269,In_18,N_912);
or U1270 (N_1270,N_908,In_382);
xnor U1271 (N_1271,In_0,N_572);
xor U1272 (N_1272,N_25,N_883);
and U1273 (N_1273,N_195,N_455);
or U1274 (N_1274,In_1408,N_864);
and U1275 (N_1275,N_866,N_285);
nor U1276 (N_1276,In_202,N_682);
and U1277 (N_1277,N_836,In_461);
nand U1278 (N_1278,N_508,N_442);
and U1279 (N_1279,N_959,N_696);
and U1280 (N_1280,N_750,N_636);
and U1281 (N_1281,In_1598,N_953);
nor U1282 (N_1282,In_1716,In_616);
nor U1283 (N_1283,N_814,In_1983);
xor U1284 (N_1284,N_688,In_1302);
nand U1285 (N_1285,N_893,N_762);
xnor U1286 (N_1286,N_996,N_899);
xnor U1287 (N_1287,N_249,N_998);
xor U1288 (N_1288,In_1473,In_1954);
nor U1289 (N_1289,In_186,In_768);
and U1290 (N_1290,N_375,N_555);
xor U1291 (N_1291,N_819,N_101);
nand U1292 (N_1292,In_1380,N_751);
and U1293 (N_1293,In_40,N_929);
nor U1294 (N_1294,N_884,N_264);
and U1295 (N_1295,N_550,N_500);
xnor U1296 (N_1296,N_501,In_1074);
or U1297 (N_1297,In_329,N_644);
nand U1298 (N_1298,N_987,N_782);
and U1299 (N_1299,In_568,N_61);
xor U1300 (N_1300,N_540,N_510);
or U1301 (N_1301,In_1785,N_664);
xnor U1302 (N_1302,N_757,N_613);
nor U1303 (N_1303,N_761,N_930);
and U1304 (N_1304,N_783,N_658);
or U1305 (N_1305,In_1607,N_178);
nor U1306 (N_1306,N_950,N_84);
or U1307 (N_1307,N_230,N_985);
and U1308 (N_1308,N_322,In_979);
nand U1309 (N_1309,N_868,N_201);
and U1310 (N_1310,N_898,N_980);
nor U1311 (N_1311,In_817,N_852);
xor U1312 (N_1312,N_863,N_820);
or U1313 (N_1313,N_86,N_599);
xnor U1314 (N_1314,N_634,N_660);
nand U1315 (N_1315,N_571,N_894);
nand U1316 (N_1316,N_962,N_638);
and U1317 (N_1317,N_585,N_339);
nand U1318 (N_1318,In_576,N_746);
and U1319 (N_1319,N_662,In_622);
nor U1320 (N_1320,N_961,In_525);
nand U1321 (N_1321,N_535,In_716);
xnor U1322 (N_1322,N_889,N_954);
and U1323 (N_1323,N_875,In_614);
nor U1324 (N_1324,In_1344,In_343);
xnor U1325 (N_1325,N_975,In_1346);
or U1326 (N_1326,N_570,In_1646);
nor U1327 (N_1327,N_796,N_506);
xnor U1328 (N_1328,N_760,N_639);
or U1329 (N_1329,N_617,N_850);
nor U1330 (N_1330,N_26,In_236);
nor U1331 (N_1331,N_648,In_796);
nor U1332 (N_1332,N_421,N_574);
nor U1333 (N_1333,N_976,N_705);
nor U1334 (N_1334,In_579,N_649);
or U1335 (N_1335,N_764,N_400);
xnor U1336 (N_1336,N_164,In_466);
nor U1337 (N_1337,In_341,N_137);
nor U1338 (N_1338,N_832,In_1202);
or U1339 (N_1339,In_1610,In_546);
or U1340 (N_1340,N_822,N_862);
or U1341 (N_1341,N_853,N_373);
or U1342 (N_1342,In_1262,N_340);
nand U1343 (N_1343,N_643,In_1951);
nand U1344 (N_1344,N_951,N_726);
nand U1345 (N_1345,N_917,N_695);
nand U1346 (N_1346,N_717,In_376);
xnor U1347 (N_1347,N_663,N_772);
and U1348 (N_1348,N_606,N_507);
and U1349 (N_1349,In_1692,In_476);
xor U1350 (N_1350,N_771,N_808);
nand U1351 (N_1351,In_1088,N_266);
and U1352 (N_1352,In_471,N_22);
nor U1353 (N_1353,N_177,N_209);
nand U1354 (N_1354,N_743,In_764);
nor U1355 (N_1355,In_1708,N_873);
xor U1356 (N_1356,N_703,In_327);
nand U1357 (N_1357,N_990,In_1139);
nand U1358 (N_1358,N_729,N_651);
nor U1359 (N_1359,N_301,In_1860);
or U1360 (N_1360,In_352,N_845);
nor U1361 (N_1361,N_564,In_1034);
and U1362 (N_1362,In_1689,N_635);
nand U1363 (N_1363,In_1833,In_630);
xor U1364 (N_1364,In_72,N_798);
or U1365 (N_1365,In_1815,In_749);
nor U1366 (N_1366,In_1417,N_578);
nand U1367 (N_1367,In_727,N_425);
xor U1368 (N_1368,N_270,N_615);
or U1369 (N_1369,N_563,In_1519);
nor U1370 (N_1370,N_824,In_527);
or U1371 (N_1371,N_809,In_770);
xnor U1372 (N_1372,In_1283,N_895);
and U1373 (N_1373,In_1208,N_63);
nand U1374 (N_1374,In_1643,N_969);
and U1375 (N_1375,N_513,N_926);
and U1376 (N_1376,N_207,N_698);
or U1377 (N_1377,N_940,N_607);
nor U1378 (N_1378,N_355,N_162);
nand U1379 (N_1379,N_481,N_981);
or U1380 (N_1380,In_1828,N_328);
nor U1381 (N_1381,N_932,In_891);
xnor U1382 (N_1382,N_906,N_704);
nor U1383 (N_1383,N_787,N_600);
and U1384 (N_1384,In_53,N_710);
nor U1385 (N_1385,In_766,N_988);
nand U1386 (N_1386,N_970,N_752);
and U1387 (N_1387,N_680,In_628);
or U1388 (N_1388,N_925,N_401);
nand U1389 (N_1389,N_150,N_986);
nand U1390 (N_1390,In_762,In_806);
nor U1391 (N_1391,N_888,In_856);
xor U1392 (N_1392,In_10,N_793);
or U1393 (N_1393,In_487,In_469);
nand U1394 (N_1394,N_902,In_1949);
xnor U1395 (N_1395,N_503,In_443);
xor U1396 (N_1396,N_799,N_877);
nand U1397 (N_1397,In_158,N_583);
nor U1398 (N_1398,N_753,N_175);
nand U1399 (N_1399,N_741,In_1990);
and U1400 (N_1400,In_49,In_203);
and U1401 (N_1401,N_983,In_543);
nand U1402 (N_1402,N_872,In_1967);
and U1403 (N_1403,In_1850,N_654);
nor U1404 (N_1404,N_587,N_591);
or U1405 (N_1405,N_19,N_40);
nand U1406 (N_1406,In_339,N_774);
nor U1407 (N_1407,N_182,In_997);
or U1408 (N_1408,In_449,N_825);
or U1409 (N_1409,N_225,N_514);
nor U1410 (N_1410,N_557,N_669);
or U1411 (N_1411,In_154,N_770);
or U1412 (N_1412,N_942,N_196);
and U1413 (N_1413,N_542,N_504);
or U1414 (N_1414,N_973,N_452);
xor U1415 (N_1415,N_437,N_784);
nor U1416 (N_1416,In_1694,N_456);
and U1417 (N_1417,N_66,N_165);
nand U1418 (N_1418,In_1792,N_330);
nand U1419 (N_1419,N_593,In_454);
nand U1420 (N_1420,N_262,In_420);
and U1421 (N_1421,N_450,N_869);
and U1422 (N_1422,N_15,N_827);
nor U1423 (N_1423,N_948,In_338);
xor U1424 (N_1424,In_1429,N_775);
or U1425 (N_1425,N_914,N_344);
or U1426 (N_1426,In_902,N_288);
nor U1427 (N_1427,In_266,In_1292);
or U1428 (N_1428,In_1641,N_28);
nand U1429 (N_1429,N_490,In_1040);
nor U1430 (N_1430,In_1569,N_846);
xnor U1431 (N_1431,In_354,N_558);
xnor U1432 (N_1432,N_815,N_978);
nor U1433 (N_1433,N_833,In_641);
xor U1434 (N_1434,N_226,N_594);
nor U1435 (N_1435,N_227,N_592);
or U1436 (N_1436,N_430,N_411);
nor U1437 (N_1437,In_1748,N_589);
nand U1438 (N_1438,N_346,N_728);
nand U1439 (N_1439,N_786,N_903);
xor U1440 (N_1440,N_347,In_288);
xnor U1441 (N_1441,N_960,In_1722);
or U1442 (N_1442,In_60,N_736);
or U1443 (N_1443,N_916,In_649);
nand U1444 (N_1444,In_1552,N_34);
and U1445 (N_1445,N_575,In_1548);
nor U1446 (N_1446,In_79,N_584);
and U1447 (N_1447,N_505,N_856);
nand U1448 (N_1448,N_955,N_806);
xor U1449 (N_1449,N_519,In_1870);
nor U1450 (N_1450,N_657,N_460);
and U1451 (N_1451,In_847,In_1245);
and U1452 (N_1452,In_960,N_56);
xor U1453 (N_1453,N_790,N_114);
xor U1454 (N_1454,In_760,N_47);
nor U1455 (N_1455,N_708,N_526);
nor U1456 (N_1456,N_715,In_221);
or U1457 (N_1457,N_766,N_911);
xnor U1458 (N_1458,In_1478,In_27);
or U1459 (N_1459,In_739,In_386);
nor U1460 (N_1460,In_1477,N_958);
or U1461 (N_1461,N_936,In_1338);
nor U1462 (N_1462,N_701,N_624);
and U1463 (N_1463,In_1447,In_989);
and U1464 (N_1464,In_585,N_957);
nand U1465 (N_1465,In_748,In_1632);
nand U1466 (N_1466,N_543,N_528);
or U1467 (N_1467,In_182,In_1198);
nor U1468 (N_1468,N_886,N_577);
or U1469 (N_1469,In_13,In_1544);
xnor U1470 (N_1470,N_529,N_382);
xnor U1471 (N_1471,N_596,N_792);
nor U1472 (N_1472,In_1089,In_366);
xnor U1473 (N_1473,N_683,N_621);
nor U1474 (N_1474,N_924,N_947);
nor U1475 (N_1475,N_993,N_29);
and U1476 (N_1476,In_1319,N_525);
xnor U1477 (N_1477,N_27,N_949);
and U1478 (N_1478,In_230,N_785);
nand U1479 (N_1479,In_375,In_1698);
xnor U1480 (N_1480,N_837,N_269);
nand U1481 (N_1481,In_1307,N_841);
xor U1482 (N_1482,N_12,N_179);
xor U1483 (N_1483,N_891,In_913);
or U1484 (N_1484,In_349,N_623);
nor U1485 (N_1485,N_559,N_684);
nor U1486 (N_1486,N_967,N_603);
nand U1487 (N_1487,N_719,In_1838);
nor U1488 (N_1488,N_516,N_632);
and U1489 (N_1489,N_918,N_839);
nand U1490 (N_1490,N_900,In_1942);
nor U1491 (N_1491,N_666,N_553);
nand U1492 (N_1492,In_499,N_560);
xor U1493 (N_1493,N_776,N_518);
or U1494 (N_1494,N_794,In_380);
xnor U1495 (N_1495,N_405,N_626);
and U1496 (N_1496,N_977,N_224);
and U1497 (N_1497,N_971,N_329);
xor U1498 (N_1498,N_754,N_713);
xnor U1499 (N_1499,N_260,N_597);
or U1500 (N_1500,N_1440,N_1358);
xor U1501 (N_1501,N_1063,N_1033);
nand U1502 (N_1502,N_1324,N_1010);
xor U1503 (N_1503,N_1349,N_1342);
xnor U1504 (N_1504,N_1370,N_1187);
nor U1505 (N_1505,N_1415,N_1079);
xor U1506 (N_1506,N_1020,N_1316);
or U1507 (N_1507,N_1400,N_1326);
nand U1508 (N_1508,N_1015,N_1492);
or U1509 (N_1509,N_1080,N_1110);
nand U1510 (N_1510,N_1484,N_1188);
xnor U1511 (N_1511,N_1221,N_1149);
or U1512 (N_1512,N_1351,N_1359);
nor U1513 (N_1513,N_1023,N_1158);
or U1514 (N_1514,N_1241,N_1369);
xnor U1515 (N_1515,N_1470,N_1275);
xor U1516 (N_1516,N_1165,N_1488);
nor U1517 (N_1517,N_1215,N_1452);
or U1518 (N_1518,N_1138,N_1334);
and U1519 (N_1519,N_1049,N_1024);
nor U1520 (N_1520,N_1398,N_1421);
nand U1521 (N_1521,N_1106,N_1093);
xor U1522 (N_1522,N_1205,N_1461);
nand U1523 (N_1523,N_1307,N_1203);
nor U1524 (N_1524,N_1026,N_1222);
and U1525 (N_1525,N_1410,N_1424);
nor U1526 (N_1526,N_1150,N_1227);
xor U1527 (N_1527,N_1490,N_1425);
nor U1528 (N_1528,N_1076,N_1048);
xor U1529 (N_1529,N_1035,N_1261);
or U1530 (N_1530,N_1312,N_1185);
and U1531 (N_1531,N_1419,N_1135);
xor U1532 (N_1532,N_1041,N_1084);
and U1533 (N_1533,N_1384,N_1070);
nand U1534 (N_1534,N_1281,N_1357);
xor U1535 (N_1535,N_1371,N_1255);
nand U1536 (N_1536,N_1477,N_1305);
xnor U1537 (N_1537,N_1061,N_1417);
xor U1538 (N_1538,N_1038,N_1167);
nor U1539 (N_1539,N_1163,N_1345);
and U1540 (N_1540,N_1431,N_1082);
xor U1541 (N_1541,N_1314,N_1169);
nor U1542 (N_1542,N_1223,N_1242);
xor U1543 (N_1543,N_1204,N_1181);
xnor U1544 (N_1544,N_1375,N_1438);
nand U1545 (N_1545,N_1253,N_1174);
nand U1546 (N_1546,N_1233,N_1091);
and U1547 (N_1547,N_1145,N_1360);
nand U1548 (N_1548,N_1140,N_1354);
xnor U1549 (N_1549,N_1151,N_1126);
or U1550 (N_1550,N_1347,N_1245);
nor U1551 (N_1551,N_1146,N_1496);
or U1552 (N_1552,N_1389,N_1131);
nor U1553 (N_1553,N_1178,N_1240);
and U1554 (N_1554,N_1113,N_1086);
nand U1555 (N_1555,N_1430,N_1045);
or U1556 (N_1556,N_1271,N_1372);
xor U1557 (N_1557,N_1030,N_1052);
nand U1558 (N_1558,N_1405,N_1081);
nor U1559 (N_1559,N_1047,N_1467);
or U1560 (N_1560,N_1127,N_1441);
nand U1561 (N_1561,N_1460,N_1473);
nand U1562 (N_1562,N_1154,N_1497);
xor U1563 (N_1563,N_1128,N_1306);
or U1564 (N_1564,N_1414,N_1226);
nor U1565 (N_1565,N_1427,N_1277);
nand U1566 (N_1566,N_1008,N_1406);
and U1567 (N_1567,N_1160,N_1159);
or U1568 (N_1568,N_1054,N_1013);
nor U1569 (N_1569,N_1195,N_1348);
or U1570 (N_1570,N_1311,N_1249);
xnor U1571 (N_1571,N_1474,N_1259);
nor U1572 (N_1572,N_1476,N_1144);
or U1573 (N_1573,N_1239,N_1450);
or U1574 (N_1574,N_1141,N_1225);
nand U1575 (N_1575,N_1236,N_1394);
xnor U1576 (N_1576,N_1278,N_1403);
nor U1577 (N_1577,N_1022,N_1433);
nand U1578 (N_1578,N_1214,N_1464);
nand U1579 (N_1579,N_1270,N_1437);
xor U1580 (N_1580,N_1420,N_1279);
and U1581 (N_1581,N_1285,N_1028);
or U1582 (N_1582,N_1147,N_1393);
and U1583 (N_1583,N_1292,N_1290);
or U1584 (N_1584,N_1273,N_1186);
and U1585 (N_1585,N_1029,N_1265);
or U1586 (N_1586,N_1336,N_1331);
nor U1587 (N_1587,N_1243,N_1300);
and U1588 (N_1588,N_1274,N_1392);
xnor U1589 (N_1589,N_1107,N_1442);
nand U1590 (N_1590,N_1044,N_1459);
nand U1591 (N_1591,N_1129,N_1269);
nor U1592 (N_1592,N_1206,N_1489);
and U1593 (N_1593,N_1175,N_1021);
and U1594 (N_1594,N_1304,N_1077);
and U1595 (N_1595,N_1379,N_1355);
nor U1596 (N_1596,N_1040,N_1257);
nand U1597 (N_1597,N_1465,N_1260);
or U1598 (N_1598,N_1017,N_1447);
and U1599 (N_1599,N_1014,N_1193);
nand U1600 (N_1600,N_1267,N_1209);
nor U1601 (N_1601,N_1212,N_1254);
nand U1602 (N_1602,N_1137,N_1074);
nor U1603 (N_1603,N_1182,N_1058);
and U1604 (N_1604,N_1196,N_1027);
xor U1605 (N_1605,N_1055,N_1344);
nor U1606 (N_1606,N_1383,N_1401);
and U1607 (N_1607,N_1287,N_1157);
and U1608 (N_1608,N_1031,N_1121);
nor U1609 (N_1609,N_1266,N_1457);
or U1610 (N_1610,N_1262,N_1268);
and U1611 (N_1611,N_1320,N_1216);
nand U1612 (N_1612,N_1059,N_1374);
nand U1613 (N_1613,N_1072,N_1130);
nor U1614 (N_1614,N_1382,N_1485);
nor U1615 (N_1615,N_1328,N_1337);
nor U1616 (N_1616,N_1201,N_1495);
and U1617 (N_1617,N_1002,N_1184);
and U1618 (N_1618,N_1179,N_1011);
or U1619 (N_1619,N_1264,N_1362);
nand U1620 (N_1620,N_1321,N_1211);
or U1621 (N_1621,N_1381,N_1418);
nand U1622 (N_1622,N_1258,N_1340);
xnor U1623 (N_1623,N_1180,N_1455);
xor U1624 (N_1624,N_1164,N_1053);
nand U1625 (N_1625,N_1098,N_1170);
nor U1626 (N_1626,N_1475,N_1089);
nor U1627 (N_1627,N_1119,N_1397);
or U1628 (N_1628,N_1118,N_1272);
xor U1629 (N_1629,N_1202,N_1120);
nor U1630 (N_1630,N_1218,N_1310);
nor U1631 (N_1631,N_1325,N_1162);
and U1632 (N_1632,N_1469,N_1487);
nand U1633 (N_1633,N_1036,N_1067);
nor U1634 (N_1634,N_1399,N_1057);
and U1635 (N_1635,N_1112,N_1220);
nor U1636 (N_1636,N_1308,N_1256);
xnor U1637 (N_1637,N_1208,N_1376);
nand U1638 (N_1638,N_1352,N_1166);
and U1639 (N_1639,N_1483,N_1378);
nand U1640 (N_1640,N_1032,N_1050);
nand U1641 (N_1641,N_1005,N_1343);
nor U1642 (N_1642,N_1230,N_1143);
and U1643 (N_1643,N_1039,N_1046);
nand U1644 (N_1644,N_1037,N_1361);
nand U1645 (N_1645,N_1191,N_1213);
and U1646 (N_1646,N_1244,N_1016);
nand U1647 (N_1647,N_1231,N_1094);
or U1648 (N_1648,N_1391,N_1333);
nand U1649 (N_1649,N_1377,N_1248);
or U1650 (N_1650,N_1114,N_1283);
nand U1651 (N_1651,N_1228,N_1282);
and U1652 (N_1652,N_1001,N_1303);
and U1653 (N_1653,N_1246,N_1408);
nor U1654 (N_1654,N_1172,N_1482);
xnor U1655 (N_1655,N_1198,N_1042);
nand U1656 (N_1656,N_1341,N_1122);
nand U1657 (N_1657,N_1060,N_1451);
xnor U1658 (N_1658,N_1066,N_1319);
nor U1659 (N_1659,N_1432,N_1125);
and U1660 (N_1660,N_1177,N_1090);
xor U1661 (N_1661,N_1004,N_1356);
or U1662 (N_1662,N_1478,N_1136);
xor U1663 (N_1663,N_1329,N_1315);
nand U1664 (N_1664,N_1051,N_1224);
or U1665 (N_1665,N_1139,N_1263);
or U1666 (N_1666,N_1353,N_1006);
nand U1667 (N_1667,N_1373,N_1366);
xor U1668 (N_1668,N_1207,N_1109);
xnor U1669 (N_1669,N_1498,N_1429);
and U1670 (N_1670,N_1439,N_1462);
or U1671 (N_1671,N_1176,N_1083);
xor U1672 (N_1672,N_1402,N_1380);
xnor U1673 (N_1673,N_1096,N_1364);
and U1674 (N_1674,N_1087,N_1108);
or U1675 (N_1675,N_1105,N_1018);
xnor U1676 (N_1676,N_1289,N_1073);
or U1677 (N_1677,N_1493,N_1449);
or U1678 (N_1678,N_1156,N_1189);
nand U1679 (N_1679,N_1210,N_1445);
or U1680 (N_1680,N_1064,N_1409);
nor U1681 (N_1681,N_1322,N_1075);
or U1682 (N_1682,N_1238,N_1390);
or U1683 (N_1683,N_1332,N_1152);
xnor U1684 (N_1684,N_1155,N_1171);
nor U1685 (N_1685,N_1363,N_1099);
nor U1686 (N_1686,N_1297,N_1251);
or U1687 (N_1687,N_1472,N_1368);
nor U1688 (N_1688,N_1346,N_1388);
nand U1689 (N_1689,N_1330,N_1088);
nor U1690 (N_1690,N_1471,N_1078);
nor U1691 (N_1691,N_1062,N_1115);
nand U1692 (N_1692,N_1302,N_1480);
nor U1693 (N_1693,N_1097,N_1291);
and U1694 (N_1694,N_1416,N_1434);
nor U1695 (N_1695,N_1365,N_1298);
or U1696 (N_1696,N_1069,N_1486);
or U1697 (N_1697,N_1288,N_1428);
or U1698 (N_1698,N_1000,N_1327);
xor U1699 (N_1699,N_1446,N_1318);
nand U1700 (N_1700,N_1499,N_1313);
xor U1701 (N_1701,N_1423,N_1200);
nand U1702 (N_1702,N_1436,N_1103);
nor U1703 (N_1703,N_1468,N_1190);
nor U1704 (N_1704,N_1095,N_1250);
or U1705 (N_1705,N_1142,N_1194);
xor U1706 (N_1706,N_1068,N_1395);
nand U1707 (N_1707,N_1229,N_1301);
and U1708 (N_1708,N_1168,N_1153);
nor U1709 (N_1709,N_1007,N_1217);
and U1710 (N_1710,N_1280,N_1435);
nor U1711 (N_1711,N_1411,N_1056);
nor U1712 (N_1712,N_1219,N_1309);
or U1713 (N_1713,N_1133,N_1386);
or U1714 (N_1714,N_1456,N_1183);
nand U1715 (N_1715,N_1479,N_1286);
nand U1716 (N_1716,N_1161,N_1123);
nor U1717 (N_1717,N_1197,N_1323);
nor U1718 (N_1718,N_1117,N_1092);
and U1719 (N_1719,N_1296,N_1339);
nor U1720 (N_1720,N_1422,N_1335);
and U1721 (N_1721,N_1148,N_1350);
nand U1722 (N_1722,N_1012,N_1111);
xor U1723 (N_1723,N_1071,N_1019);
nor U1724 (N_1724,N_1367,N_1124);
or U1725 (N_1725,N_1101,N_1116);
nor U1726 (N_1726,N_1293,N_1294);
nor U1727 (N_1727,N_1003,N_1134);
and U1728 (N_1728,N_1043,N_1235);
nand U1729 (N_1729,N_1299,N_1199);
and U1730 (N_1730,N_1284,N_1454);
xor U1731 (N_1731,N_1338,N_1412);
and U1732 (N_1732,N_1173,N_1065);
and U1733 (N_1733,N_1466,N_1443);
xnor U1734 (N_1734,N_1102,N_1407);
nand U1735 (N_1735,N_1295,N_1276);
xnor U1736 (N_1736,N_1237,N_1491);
or U1737 (N_1737,N_1234,N_1034);
and U1738 (N_1738,N_1404,N_1247);
nand U1739 (N_1739,N_1252,N_1494);
xnor U1740 (N_1740,N_1317,N_1009);
and U1741 (N_1741,N_1448,N_1192);
nor U1742 (N_1742,N_1085,N_1413);
xnor U1743 (N_1743,N_1396,N_1481);
nand U1744 (N_1744,N_1232,N_1385);
xor U1745 (N_1745,N_1025,N_1426);
xnor U1746 (N_1746,N_1444,N_1463);
xnor U1747 (N_1747,N_1453,N_1100);
nor U1748 (N_1748,N_1387,N_1104);
xnor U1749 (N_1749,N_1132,N_1458);
nand U1750 (N_1750,N_1465,N_1255);
and U1751 (N_1751,N_1050,N_1072);
or U1752 (N_1752,N_1201,N_1309);
and U1753 (N_1753,N_1420,N_1393);
xnor U1754 (N_1754,N_1328,N_1284);
xor U1755 (N_1755,N_1462,N_1423);
nand U1756 (N_1756,N_1187,N_1293);
nor U1757 (N_1757,N_1124,N_1238);
nand U1758 (N_1758,N_1321,N_1278);
and U1759 (N_1759,N_1299,N_1292);
nand U1760 (N_1760,N_1405,N_1084);
xor U1761 (N_1761,N_1204,N_1198);
or U1762 (N_1762,N_1197,N_1252);
nor U1763 (N_1763,N_1262,N_1453);
and U1764 (N_1764,N_1237,N_1206);
xor U1765 (N_1765,N_1232,N_1126);
and U1766 (N_1766,N_1087,N_1302);
nor U1767 (N_1767,N_1170,N_1174);
nor U1768 (N_1768,N_1443,N_1318);
and U1769 (N_1769,N_1170,N_1077);
nor U1770 (N_1770,N_1103,N_1256);
and U1771 (N_1771,N_1478,N_1416);
nor U1772 (N_1772,N_1161,N_1392);
or U1773 (N_1773,N_1171,N_1093);
nor U1774 (N_1774,N_1128,N_1379);
and U1775 (N_1775,N_1145,N_1343);
nor U1776 (N_1776,N_1218,N_1459);
nor U1777 (N_1777,N_1131,N_1002);
and U1778 (N_1778,N_1400,N_1170);
nor U1779 (N_1779,N_1286,N_1290);
nor U1780 (N_1780,N_1191,N_1469);
nand U1781 (N_1781,N_1311,N_1116);
nand U1782 (N_1782,N_1050,N_1383);
nor U1783 (N_1783,N_1269,N_1430);
or U1784 (N_1784,N_1462,N_1127);
and U1785 (N_1785,N_1497,N_1151);
nor U1786 (N_1786,N_1098,N_1162);
or U1787 (N_1787,N_1439,N_1392);
or U1788 (N_1788,N_1071,N_1409);
xnor U1789 (N_1789,N_1100,N_1304);
or U1790 (N_1790,N_1345,N_1119);
nand U1791 (N_1791,N_1061,N_1489);
and U1792 (N_1792,N_1103,N_1106);
nand U1793 (N_1793,N_1169,N_1349);
xnor U1794 (N_1794,N_1378,N_1079);
nand U1795 (N_1795,N_1285,N_1168);
nor U1796 (N_1796,N_1162,N_1054);
or U1797 (N_1797,N_1352,N_1120);
or U1798 (N_1798,N_1393,N_1339);
nand U1799 (N_1799,N_1115,N_1038);
nand U1800 (N_1800,N_1210,N_1230);
nand U1801 (N_1801,N_1088,N_1092);
and U1802 (N_1802,N_1142,N_1149);
nand U1803 (N_1803,N_1004,N_1318);
and U1804 (N_1804,N_1274,N_1052);
xor U1805 (N_1805,N_1420,N_1486);
xnor U1806 (N_1806,N_1442,N_1167);
and U1807 (N_1807,N_1186,N_1238);
or U1808 (N_1808,N_1088,N_1446);
xnor U1809 (N_1809,N_1442,N_1216);
and U1810 (N_1810,N_1097,N_1293);
xnor U1811 (N_1811,N_1376,N_1193);
nor U1812 (N_1812,N_1190,N_1093);
or U1813 (N_1813,N_1125,N_1341);
xnor U1814 (N_1814,N_1109,N_1378);
and U1815 (N_1815,N_1404,N_1097);
xor U1816 (N_1816,N_1338,N_1006);
xor U1817 (N_1817,N_1126,N_1491);
nor U1818 (N_1818,N_1025,N_1244);
xor U1819 (N_1819,N_1224,N_1042);
and U1820 (N_1820,N_1493,N_1115);
and U1821 (N_1821,N_1334,N_1181);
and U1822 (N_1822,N_1043,N_1485);
nand U1823 (N_1823,N_1471,N_1416);
xor U1824 (N_1824,N_1055,N_1033);
nand U1825 (N_1825,N_1298,N_1045);
and U1826 (N_1826,N_1451,N_1053);
nand U1827 (N_1827,N_1279,N_1153);
or U1828 (N_1828,N_1048,N_1388);
nand U1829 (N_1829,N_1322,N_1195);
and U1830 (N_1830,N_1307,N_1375);
nor U1831 (N_1831,N_1244,N_1310);
xnor U1832 (N_1832,N_1313,N_1464);
nor U1833 (N_1833,N_1297,N_1361);
and U1834 (N_1834,N_1329,N_1000);
nand U1835 (N_1835,N_1073,N_1014);
and U1836 (N_1836,N_1465,N_1297);
or U1837 (N_1837,N_1086,N_1192);
and U1838 (N_1838,N_1360,N_1333);
or U1839 (N_1839,N_1309,N_1126);
or U1840 (N_1840,N_1350,N_1052);
nand U1841 (N_1841,N_1407,N_1207);
nor U1842 (N_1842,N_1282,N_1330);
nand U1843 (N_1843,N_1349,N_1172);
and U1844 (N_1844,N_1425,N_1421);
or U1845 (N_1845,N_1343,N_1214);
xnor U1846 (N_1846,N_1223,N_1079);
nor U1847 (N_1847,N_1220,N_1284);
nand U1848 (N_1848,N_1240,N_1045);
and U1849 (N_1849,N_1439,N_1351);
or U1850 (N_1850,N_1277,N_1487);
or U1851 (N_1851,N_1367,N_1425);
or U1852 (N_1852,N_1484,N_1178);
or U1853 (N_1853,N_1216,N_1324);
or U1854 (N_1854,N_1134,N_1226);
and U1855 (N_1855,N_1229,N_1390);
xnor U1856 (N_1856,N_1106,N_1146);
and U1857 (N_1857,N_1452,N_1027);
nand U1858 (N_1858,N_1209,N_1327);
nor U1859 (N_1859,N_1282,N_1028);
or U1860 (N_1860,N_1384,N_1256);
nand U1861 (N_1861,N_1037,N_1241);
xnor U1862 (N_1862,N_1068,N_1467);
and U1863 (N_1863,N_1331,N_1318);
and U1864 (N_1864,N_1327,N_1314);
or U1865 (N_1865,N_1192,N_1019);
nand U1866 (N_1866,N_1337,N_1309);
or U1867 (N_1867,N_1118,N_1368);
or U1868 (N_1868,N_1482,N_1165);
or U1869 (N_1869,N_1312,N_1139);
and U1870 (N_1870,N_1404,N_1285);
nor U1871 (N_1871,N_1330,N_1229);
nor U1872 (N_1872,N_1307,N_1354);
xnor U1873 (N_1873,N_1403,N_1154);
xor U1874 (N_1874,N_1316,N_1450);
nand U1875 (N_1875,N_1027,N_1335);
nand U1876 (N_1876,N_1215,N_1223);
xnor U1877 (N_1877,N_1149,N_1315);
or U1878 (N_1878,N_1358,N_1352);
nand U1879 (N_1879,N_1065,N_1138);
or U1880 (N_1880,N_1099,N_1196);
nor U1881 (N_1881,N_1147,N_1287);
nand U1882 (N_1882,N_1471,N_1192);
nand U1883 (N_1883,N_1344,N_1317);
and U1884 (N_1884,N_1019,N_1488);
xor U1885 (N_1885,N_1499,N_1201);
nand U1886 (N_1886,N_1470,N_1465);
nand U1887 (N_1887,N_1202,N_1171);
nand U1888 (N_1888,N_1399,N_1409);
or U1889 (N_1889,N_1374,N_1109);
nand U1890 (N_1890,N_1191,N_1489);
or U1891 (N_1891,N_1463,N_1073);
nand U1892 (N_1892,N_1347,N_1477);
and U1893 (N_1893,N_1307,N_1154);
and U1894 (N_1894,N_1465,N_1374);
nand U1895 (N_1895,N_1239,N_1467);
nand U1896 (N_1896,N_1198,N_1373);
nor U1897 (N_1897,N_1233,N_1411);
and U1898 (N_1898,N_1168,N_1061);
nand U1899 (N_1899,N_1074,N_1353);
xnor U1900 (N_1900,N_1414,N_1393);
or U1901 (N_1901,N_1169,N_1184);
nand U1902 (N_1902,N_1487,N_1427);
and U1903 (N_1903,N_1040,N_1269);
nand U1904 (N_1904,N_1172,N_1366);
xor U1905 (N_1905,N_1485,N_1413);
nand U1906 (N_1906,N_1471,N_1244);
nor U1907 (N_1907,N_1005,N_1406);
nand U1908 (N_1908,N_1082,N_1274);
xnor U1909 (N_1909,N_1110,N_1061);
or U1910 (N_1910,N_1457,N_1117);
or U1911 (N_1911,N_1428,N_1063);
xnor U1912 (N_1912,N_1403,N_1416);
or U1913 (N_1913,N_1408,N_1155);
nor U1914 (N_1914,N_1373,N_1355);
xnor U1915 (N_1915,N_1058,N_1238);
and U1916 (N_1916,N_1494,N_1218);
or U1917 (N_1917,N_1158,N_1032);
nor U1918 (N_1918,N_1435,N_1476);
xnor U1919 (N_1919,N_1442,N_1225);
xor U1920 (N_1920,N_1237,N_1379);
or U1921 (N_1921,N_1306,N_1072);
and U1922 (N_1922,N_1113,N_1432);
and U1923 (N_1923,N_1300,N_1184);
nand U1924 (N_1924,N_1087,N_1152);
and U1925 (N_1925,N_1083,N_1091);
xnor U1926 (N_1926,N_1229,N_1016);
xnor U1927 (N_1927,N_1474,N_1455);
and U1928 (N_1928,N_1168,N_1385);
xor U1929 (N_1929,N_1435,N_1042);
or U1930 (N_1930,N_1357,N_1388);
nor U1931 (N_1931,N_1022,N_1180);
and U1932 (N_1932,N_1439,N_1269);
and U1933 (N_1933,N_1321,N_1393);
or U1934 (N_1934,N_1363,N_1338);
or U1935 (N_1935,N_1375,N_1355);
nor U1936 (N_1936,N_1072,N_1308);
and U1937 (N_1937,N_1449,N_1450);
nand U1938 (N_1938,N_1395,N_1080);
and U1939 (N_1939,N_1359,N_1239);
and U1940 (N_1940,N_1210,N_1255);
and U1941 (N_1941,N_1181,N_1339);
nor U1942 (N_1942,N_1138,N_1152);
xor U1943 (N_1943,N_1278,N_1002);
nor U1944 (N_1944,N_1468,N_1065);
nand U1945 (N_1945,N_1369,N_1197);
nor U1946 (N_1946,N_1158,N_1410);
xor U1947 (N_1947,N_1014,N_1424);
nand U1948 (N_1948,N_1312,N_1234);
xnor U1949 (N_1949,N_1204,N_1352);
xor U1950 (N_1950,N_1026,N_1249);
or U1951 (N_1951,N_1069,N_1439);
nor U1952 (N_1952,N_1397,N_1223);
nor U1953 (N_1953,N_1241,N_1443);
nand U1954 (N_1954,N_1430,N_1497);
or U1955 (N_1955,N_1122,N_1087);
nor U1956 (N_1956,N_1058,N_1467);
and U1957 (N_1957,N_1062,N_1019);
nand U1958 (N_1958,N_1247,N_1213);
or U1959 (N_1959,N_1150,N_1068);
or U1960 (N_1960,N_1213,N_1229);
and U1961 (N_1961,N_1389,N_1275);
and U1962 (N_1962,N_1428,N_1426);
nand U1963 (N_1963,N_1483,N_1466);
nand U1964 (N_1964,N_1352,N_1287);
or U1965 (N_1965,N_1176,N_1294);
or U1966 (N_1966,N_1210,N_1439);
and U1967 (N_1967,N_1182,N_1324);
and U1968 (N_1968,N_1394,N_1139);
xor U1969 (N_1969,N_1402,N_1465);
and U1970 (N_1970,N_1440,N_1093);
and U1971 (N_1971,N_1039,N_1146);
and U1972 (N_1972,N_1353,N_1033);
or U1973 (N_1973,N_1326,N_1024);
xnor U1974 (N_1974,N_1167,N_1096);
nand U1975 (N_1975,N_1468,N_1312);
xnor U1976 (N_1976,N_1118,N_1205);
nand U1977 (N_1977,N_1210,N_1471);
and U1978 (N_1978,N_1142,N_1170);
nor U1979 (N_1979,N_1175,N_1279);
and U1980 (N_1980,N_1452,N_1305);
nand U1981 (N_1981,N_1422,N_1072);
nand U1982 (N_1982,N_1152,N_1437);
xnor U1983 (N_1983,N_1225,N_1091);
and U1984 (N_1984,N_1261,N_1298);
nor U1985 (N_1985,N_1201,N_1422);
and U1986 (N_1986,N_1099,N_1326);
and U1987 (N_1987,N_1251,N_1258);
nand U1988 (N_1988,N_1327,N_1358);
xnor U1989 (N_1989,N_1060,N_1174);
xor U1990 (N_1990,N_1126,N_1459);
or U1991 (N_1991,N_1173,N_1319);
nand U1992 (N_1992,N_1240,N_1055);
or U1993 (N_1993,N_1041,N_1037);
xor U1994 (N_1994,N_1402,N_1028);
nor U1995 (N_1995,N_1167,N_1428);
or U1996 (N_1996,N_1340,N_1079);
nand U1997 (N_1997,N_1115,N_1196);
nor U1998 (N_1998,N_1207,N_1461);
nor U1999 (N_1999,N_1470,N_1293);
nand U2000 (N_2000,N_1599,N_1765);
nand U2001 (N_2001,N_1965,N_1829);
or U2002 (N_2002,N_1523,N_1676);
nor U2003 (N_2003,N_1884,N_1846);
or U2004 (N_2004,N_1951,N_1998);
nand U2005 (N_2005,N_1573,N_1686);
or U2006 (N_2006,N_1997,N_1612);
xor U2007 (N_2007,N_1794,N_1899);
nor U2008 (N_2008,N_1742,N_1943);
nor U2009 (N_2009,N_1613,N_1597);
xnor U2010 (N_2010,N_1946,N_1865);
and U2011 (N_2011,N_1770,N_1890);
nor U2012 (N_2012,N_1838,N_1729);
and U2013 (N_2013,N_1807,N_1837);
nor U2014 (N_2014,N_1856,N_1505);
nor U2015 (N_2015,N_1702,N_1559);
xnor U2016 (N_2016,N_1691,N_1693);
and U2017 (N_2017,N_1840,N_1562);
nand U2018 (N_2018,N_1969,N_1642);
xnor U2019 (N_2019,N_1787,N_1883);
nand U2020 (N_2020,N_1684,N_1879);
nor U2021 (N_2021,N_1836,N_1720);
xnor U2022 (N_2022,N_1581,N_1761);
nand U2023 (N_2023,N_1726,N_1782);
nand U2024 (N_2024,N_1985,N_1803);
nand U2025 (N_2025,N_1610,N_1519);
nor U2026 (N_2026,N_1930,N_1931);
xnor U2027 (N_2027,N_1821,N_1949);
nor U2028 (N_2028,N_1815,N_1939);
nor U2029 (N_2029,N_1587,N_1988);
nand U2030 (N_2030,N_1517,N_1711);
nor U2031 (N_2031,N_1744,N_1816);
and U2032 (N_2032,N_1525,N_1889);
nor U2033 (N_2033,N_1666,N_1870);
or U2034 (N_2034,N_1574,N_1800);
and U2035 (N_2035,N_1506,N_1905);
nor U2036 (N_2036,N_1772,N_1937);
nand U2037 (N_2037,N_1601,N_1593);
or U2038 (N_2038,N_1552,N_1826);
or U2039 (N_2039,N_1755,N_1877);
xor U2040 (N_2040,N_1553,N_1687);
and U2041 (N_2041,N_1814,N_1618);
or U2042 (N_2042,N_1619,N_1888);
or U2043 (N_2043,N_1564,N_1764);
nor U2044 (N_2044,N_1876,N_1784);
nand U2045 (N_2045,N_1802,N_1674);
nor U2046 (N_2046,N_1945,N_1911);
and U2047 (N_2047,N_1694,N_1961);
nor U2048 (N_2048,N_1842,N_1844);
and U2049 (N_2049,N_1653,N_1766);
and U2050 (N_2050,N_1735,N_1572);
nor U2051 (N_2051,N_1960,N_1586);
xnor U2052 (N_2052,N_1973,N_1896);
xor U2053 (N_2053,N_1692,N_1790);
nor U2054 (N_2054,N_1512,N_1547);
nand U2055 (N_2055,N_1660,N_1806);
and U2056 (N_2056,N_1500,N_1809);
or U2057 (N_2057,N_1866,N_1994);
or U2058 (N_2058,N_1835,N_1665);
or U2059 (N_2059,N_1914,N_1753);
or U2060 (N_2060,N_1743,N_1585);
nor U2061 (N_2061,N_1626,N_1526);
xnor U2062 (N_2062,N_1857,N_1947);
nand U2063 (N_2063,N_1819,N_1875);
nand U2064 (N_2064,N_1780,N_1749);
xor U2065 (N_2065,N_1594,N_1541);
nand U2066 (N_2066,N_1569,N_1959);
xnor U2067 (N_2067,N_1705,N_1941);
nor U2068 (N_2068,N_1556,N_1680);
nor U2069 (N_2069,N_1813,N_1577);
or U2070 (N_2070,N_1623,N_1774);
or U2071 (N_2071,N_1799,N_1608);
or U2072 (N_2072,N_1980,N_1964);
and U2073 (N_2073,N_1810,N_1703);
nor U2074 (N_2074,N_1617,N_1528);
nand U2075 (N_2075,N_1622,N_1918);
nand U2076 (N_2076,N_1841,N_1935);
nand U2077 (N_2077,N_1565,N_1558);
nand U2078 (N_2078,N_1536,N_1696);
xor U2079 (N_2079,N_1724,N_1737);
nor U2080 (N_2080,N_1631,N_1926);
xnor U2081 (N_2081,N_1797,N_1812);
xor U2082 (N_2082,N_1741,N_1853);
nand U2083 (N_2083,N_1944,N_1887);
or U2084 (N_2084,N_1561,N_1527);
nand U2085 (N_2085,N_1637,N_1791);
nand U2086 (N_2086,N_1940,N_1854);
or U2087 (N_2087,N_1751,N_1700);
nor U2088 (N_2088,N_1921,N_1954);
xor U2089 (N_2089,N_1628,N_1717);
xnor U2090 (N_2090,N_1646,N_1859);
and U2091 (N_2091,N_1509,N_1834);
and U2092 (N_2092,N_1828,N_1847);
and U2093 (N_2093,N_1669,N_1993);
nand U2094 (N_2094,N_1734,N_1952);
or U2095 (N_2095,N_1625,N_1897);
nor U2096 (N_2096,N_1578,N_1502);
nor U2097 (N_2097,N_1658,N_1670);
nand U2098 (N_2098,N_1977,N_1732);
nand U2099 (N_2099,N_1706,N_1663);
xnor U2100 (N_2100,N_1793,N_1839);
nand U2101 (N_2101,N_1685,N_1886);
xnor U2102 (N_2102,N_1563,N_1583);
nand U2103 (N_2103,N_1754,N_1624);
xnor U2104 (N_2104,N_1615,N_1867);
xnor U2105 (N_2105,N_1704,N_1823);
nand U2106 (N_2106,N_1588,N_1598);
and U2107 (N_2107,N_1745,N_1648);
xor U2108 (N_2108,N_1683,N_1970);
nor U2109 (N_2109,N_1881,N_1928);
xnor U2110 (N_2110,N_1851,N_1657);
and U2111 (N_2111,N_1689,N_1983);
nor U2112 (N_2112,N_1645,N_1664);
or U2113 (N_2113,N_1701,N_1773);
and U2114 (N_2114,N_1752,N_1638);
and U2115 (N_2115,N_1589,N_1739);
or U2116 (N_2116,N_1592,N_1820);
nand U2117 (N_2117,N_1798,N_1833);
xor U2118 (N_2118,N_1762,N_1900);
xnor U2119 (N_2119,N_1609,N_1759);
or U2120 (N_2120,N_1981,N_1882);
or U2121 (N_2121,N_1655,N_1603);
xor U2122 (N_2122,N_1554,N_1989);
and U2123 (N_2123,N_1605,N_1920);
and U2124 (N_2124,N_1795,N_1571);
xor U2125 (N_2125,N_1864,N_1709);
nor U2126 (N_2126,N_1874,N_1781);
or U2127 (N_2127,N_1768,N_1650);
nand U2128 (N_2128,N_1649,N_1933);
and U2129 (N_2129,N_1986,N_1942);
and U2130 (N_2130,N_1999,N_1629);
or U2131 (N_2131,N_1818,N_1555);
nand U2132 (N_2132,N_1919,N_1777);
nor U2133 (N_2133,N_1643,N_1641);
nor U2134 (N_2134,N_1962,N_1904);
nor U2135 (N_2135,N_1721,N_1630);
and U2136 (N_2136,N_1733,N_1544);
nor U2137 (N_2137,N_1785,N_1934);
and U2138 (N_2138,N_1968,N_1927);
xor U2139 (N_2139,N_1640,N_1746);
nand U2140 (N_2140,N_1974,N_1542);
nand U2141 (N_2141,N_1673,N_1923);
nor U2142 (N_2142,N_1659,N_1667);
xnor U2143 (N_2143,N_1539,N_1924);
or U2144 (N_2144,N_1596,N_1675);
or U2145 (N_2145,N_1730,N_1860);
or U2146 (N_2146,N_1540,N_1995);
and U2147 (N_2147,N_1932,N_1632);
and U2148 (N_2148,N_1568,N_1894);
xor U2149 (N_2149,N_1783,N_1710);
or U2150 (N_2150,N_1727,N_1796);
and U2151 (N_2151,N_1567,N_1906);
nand U2152 (N_2152,N_1551,N_1672);
and U2153 (N_2153,N_1644,N_1576);
nand U2154 (N_2154,N_1714,N_1908);
xnor U2155 (N_2155,N_1849,N_1805);
nor U2156 (N_2156,N_1843,N_1695);
and U2157 (N_2157,N_1756,N_1991);
nor U2158 (N_2158,N_1775,N_1521);
and U2159 (N_2159,N_1907,N_1736);
or U2160 (N_2160,N_1917,N_1582);
nand U2161 (N_2161,N_1858,N_1716);
or U2162 (N_2162,N_1713,N_1822);
or U2163 (N_2163,N_1824,N_1501);
nor U2164 (N_2164,N_1901,N_1925);
nor U2165 (N_2165,N_1671,N_1808);
or U2166 (N_2166,N_1878,N_1845);
nand U2167 (N_2167,N_1715,N_1992);
nor U2168 (N_2168,N_1915,N_1682);
and U2169 (N_2169,N_1507,N_1862);
nand U2170 (N_2170,N_1910,N_1913);
or U2171 (N_2171,N_1872,N_1712);
nand U2172 (N_2172,N_1690,N_1535);
or U2173 (N_2173,N_1662,N_1902);
xnor U2174 (N_2174,N_1855,N_1634);
and U2175 (N_2175,N_1955,N_1725);
nand U2176 (N_2176,N_1976,N_1757);
nor U2177 (N_2177,N_1817,N_1533);
nand U2178 (N_2178,N_1922,N_1750);
nand U2179 (N_2179,N_1990,N_1731);
or U2180 (N_2180,N_1560,N_1909);
or U2181 (N_2181,N_1788,N_1548);
xor U2182 (N_2182,N_1825,N_1779);
and U2183 (N_2183,N_1723,N_1957);
nor U2184 (N_2184,N_1831,N_1863);
and U2185 (N_2185,N_1604,N_1880);
and U2186 (N_2186,N_1679,N_1530);
nand U2187 (N_2187,N_1982,N_1979);
nor U2188 (N_2188,N_1852,N_1570);
nor U2189 (N_2189,N_1871,N_1892);
xor U2190 (N_2190,N_1748,N_1738);
xnor U2191 (N_2191,N_1963,N_1929);
nor U2192 (N_2192,N_1621,N_1504);
or U2193 (N_2193,N_1639,N_1967);
and U2194 (N_2194,N_1869,N_1545);
and U2195 (N_2195,N_1938,N_1614);
or U2196 (N_2196,N_1789,N_1543);
nand U2197 (N_2197,N_1956,N_1698);
or U2198 (N_2198,N_1699,N_1513);
or U2199 (N_2199,N_1747,N_1776);
and U2200 (N_2200,N_1978,N_1972);
nor U2201 (N_2201,N_1778,N_1678);
xnor U2202 (N_2202,N_1635,N_1531);
nor U2203 (N_2203,N_1893,N_1868);
nor U2204 (N_2204,N_1651,N_1936);
nor U2205 (N_2205,N_1616,N_1861);
nor U2206 (N_2206,N_1804,N_1903);
or U2207 (N_2207,N_1654,N_1885);
xnor U2208 (N_2208,N_1811,N_1950);
and U2209 (N_2209,N_1740,N_1719);
nand U2210 (N_2210,N_1830,N_1546);
nand U2211 (N_2211,N_1850,N_1771);
or U2212 (N_2212,N_1827,N_1677);
or U2213 (N_2213,N_1516,N_1891);
nor U2214 (N_2214,N_1832,N_1873);
and U2215 (N_2215,N_1550,N_1848);
nor U2216 (N_2216,N_1707,N_1514);
nand U2217 (N_2217,N_1579,N_1984);
or U2218 (N_2218,N_1515,N_1996);
xnor U2219 (N_2219,N_1600,N_1681);
xnor U2220 (N_2220,N_1607,N_1549);
and U2221 (N_2221,N_1627,N_1520);
nand U2222 (N_2222,N_1503,N_1538);
or U2223 (N_2223,N_1580,N_1524);
xnor U2224 (N_2224,N_1786,N_1590);
or U2225 (N_2225,N_1760,N_1611);
nor U2226 (N_2226,N_1566,N_1895);
nand U2227 (N_2227,N_1602,N_1975);
and U2228 (N_2228,N_1591,N_1511);
and U2229 (N_2229,N_1584,N_1529);
and U2230 (N_2230,N_1718,N_1953);
nand U2231 (N_2231,N_1971,N_1661);
and U2232 (N_2232,N_1688,N_1508);
or U2233 (N_2233,N_1633,N_1534);
or U2234 (N_2234,N_1697,N_1758);
xnor U2235 (N_2235,N_1763,N_1575);
and U2236 (N_2236,N_1537,N_1652);
xor U2237 (N_2237,N_1966,N_1916);
nor U2238 (N_2238,N_1801,N_1728);
nor U2239 (N_2239,N_1636,N_1647);
or U2240 (N_2240,N_1606,N_1769);
xnor U2241 (N_2241,N_1708,N_1522);
or U2242 (N_2242,N_1656,N_1532);
or U2243 (N_2243,N_1948,N_1620);
and U2244 (N_2244,N_1898,N_1668);
or U2245 (N_2245,N_1518,N_1792);
nor U2246 (N_2246,N_1595,N_1510);
and U2247 (N_2247,N_1722,N_1958);
nor U2248 (N_2248,N_1912,N_1557);
xor U2249 (N_2249,N_1767,N_1987);
nand U2250 (N_2250,N_1876,N_1817);
nor U2251 (N_2251,N_1751,N_1516);
and U2252 (N_2252,N_1679,N_1536);
nand U2253 (N_2253,N_1794,N_1617);
and U2254 (N_2254,N_1822,N_1670);
nor U2255 (N_2255,N_1956,N_1743);
nand U2256 (N_2256,N_1784,N_1938);
or U2257 (N_2257,N_1887,N_1878);
xnor U2258 (N_2258,N_1529,N_1950);
or U2259 (N_2259,N_1635,N_1668);
and U2260 (N_2260,N_1509,N_1827);
or U2261 (N_2261,N_1948,N_1601);
and U2262 (N_2262,N_1940,N_1828);
and U2263 (N_2263,N_1924,N_1617);
nor U2264 (N_2264,N_1954,N_1761);
nand U2265 (N_2265,N_1907,N_1775);
or U2266 (N_2266,N_1637,N_1541);
xor U2267 (N_2267,N_1814,N_1750);
and U2268 (N_2268,N_1506,N_1880);
nand U2269 (N_2269,N_1561,N_1535);
nand U2270 (N_2270,N_1622,N_1985);
nand U2271 (N_2271,N_1985,N_1786);
or U2272 (N_2272,N_1868,N_1889);
nor U2273 (N_2273,N_1835,N_1917);
nor U2274 (N_2274,N_1521,N_1793);
or U2275 (N_2275,N_1625,N_1816);
xnor U2276 (N_2276,N_1731,N_1930);
and U2277 (N_2277,N_1917,N_1837);
and U2278 (N_2278,N_1646,N_1940);
or U2279 (N_2279,N_1911,N_1899);
and U2280 (N_2280,N_1732,N_1962);
xnor U2281 (N_2281,N_1795,N_1858);
xnor U2282 (N_2282,N_1973,N_1982);
or U2283 (N_2283,N_1945,N_1516);
nor U2284 (N_2284,N_1946,N_1810);
and U2285 (N_2285,N_1679,N_1629);
nand U2286 (N_2286,N_1576,N_1548);
or U2287 (N_2287,N_1776,N_1929);
and U2288 (N_2288,N_1512,N_1862);
nand U2289 (N_2289,N_1643,N_1947);
and U2290 (N_2290,N_1554,N_1632);
nand U2291 (N_2291,N_1571,N_1662);
xor U2292 (N_2292,N_1705,N_1708);
nor U2293 (N_2293,N_1840,N_1852);
and U2294 (N_2294,N_1775,N_1840);
and U2295 (N_2295,N_1663,N_1911);
xor U2296 (N_2296,N_1638,N_1645);
and U2297 (N_2297,N_1520,N_1694);
nor U2298 (N_2298,N_1510,N_1628);
and U2299 (N_2299,N_1569,N_1667);
and U2300 (N_2300,N_1911,N_1664);
or U2301 (N_2301,N_1637,N_1742);
xor U2302 (N_2302,N_1891,N_1701);
and U2303 (N_2303,N_1952,N_1758);
nor U2304 (N_2304,N_1523,N_1793);
nor U2305 (N_2305,N_1860,N_1553);
nor U2306 (N_2306,N_1600,N_1952);
and U2307 (N_2307,N_1889,N_1596);
or U2308 (N_2308,N_1884,N_1803);
or U2309 (N_2309,N_1925,N_1711);
nand U2310 (N_2310,N_1894,N_1704);
nand U2311 (N_2311,N_1554,N_1576);
nand U2312 (N_2312,N_1711,N_1505);
nand U2313 (N_2313,N_1680,N_1638);
and U2314 (N_2314,N_1877,N_1739);
nor U2315 (N_2315,N_1876,N_1923);
nor U2316 (N_2316,N_1692,N_1658);
or U2317 (N_2317,N_1657,N_1986);
or U2318 (N_2318,N_1777,N_1906);
nand U2319 (N_2319,N_1590,N_1951);
or U2320 (N_2320,N_1656,N_1902);
nor U2321 (N_2321,N_1759,N_1705);
nand U2322 (N_2322,N_1881,N_1966);
or U2323 (N_2323,N_1910,N_1862);
and U2324 (N_2324,N_1995,N_1506);
and U2325 (N_2325,N_1714,N_1798);
xnor U2326 (N_2326,N_1593,N_1594);
nand U2327 (N_2327,N_1531,N_1954);
nand U2328 (N_2328,N_1866,N_1981);
and U2329 (N_2329,N_1556,N_1706);
nor U2330 (N_2330,N_1792,N_1597);
and U2331 (N_2331,N_1777,N_1731);
and U2332 (N_2332,N_1951,N_1734);
nand U2333 (N_2333,N_1802,N_1889);
or U2334 (N_2334,N_1807,N_1979);
nor U2335 (N_2335,N_1897,N_1559);
xor U2336 (N_2336,N_1970,N_1655);
xnor U2337 (N_2337,N_1598,N_1866);
xnor U2338 (N_2338,N_1799,N_1996);
or U2339 (N_2339,N_1711,N_1834);
nor U2340 (N_2340,N_1878,N_1988);
xnor U2341 (N_2341,N_1675,N_1814);
or U2342 (N_2342,N_1508,N_1633);
nor U2343 (N_2343,N_1828,N_1928);
nor U2344 (N_2344,N_1639,N_1857);
nor U2345 (N_2345,N_1960,N_1578);
nand U2346 (N_2346,N_1923,N_1886);
and U2347 (N_2347,N_1797,N_1816);
nor U2348 (N_2348,N_1767,N_1974);
or U2349 (N_2349,N_1820,N_1951);
and U2350 (N_2350,N_1784,N_1971);
or U2351 (N_2351,N_1854,N_1810);
xnor U2352 (N_2352,N_1520,N_1622);
nand U2353 (N_2353,N_1963,N_1866);
or U2354 (N_2354,N_1875,N_1729);
xnor U2355 (N_2355,N_1777,N_1597);
or U2356 (N_2356,N_1793,N_1833);
xnor U2357 (N_2357,N_1875,N_1876);
xor U2358 (N_2358,N_1686,N_1898);
nor U2359 (N_2359,N_1538,N_1715);
and U2360 (N_2360,N_1658,N_1717);
and U2361 (N_2361,N_1691,N_1544);
nor U2362 (N_2362,N_1779,N_1549);
nand U2363 (N_2363,N_1837,N_1572);
xor U2364 (N_2364,N_1890,N_1959);
nor U2365 (N_2365,N_1843,N_1792);
nand U2366 (N_2366,N_1679,N_1711);
or U2367 (N_2367,N_1674,N_1962);
or U2368 (N_2368,N_1929,N_1807);
or U2369 (N_2369,N_1624,N_1776);
or U2370 (N_2370,N_1696,N_1601);
and U2371 (N_2371,N_1992,N_1638);
xnor U2372 (N_2372,N_1570,N_1999);
nor U2373 (N_2373,N_1737,N_1640);
or U2374 (N_2374,N_1689,N_1929);
and U2375 (N_2375,N_1600,N_1535);
and U2376 (N_2376,N_1553,N_1633);
and U2377 (N_2377,N_1645,N_1784);
xor U2378 (N_2378,N_1546,N_1961);
or U2379 (N_2379,N_1971,N_1907);
or U2380 (N_2380,N_1809,N_1823);
nand U2381 (N_2381,N_1574,N_1940);
xnor U2382 (N_2382,N_1532,N_1802);
nor U2383 (N_2383,N_1609,N_1809);
nand U2384 (N_2384,N_1864,N_1663);
and U2385 (N_2385,N_1994,N_1576);
nor U2386 (N_2386,N_1850,N_1845);
or U2387 (N_2387,N_1609,N_1554);
or U2388 (N_2388,N_1937,N_1928);
nand U2389 (N_2389,N_1560,N_1638);
nor U2390 (N_2390,N_1937,N_1892);
xnor U2391 (N_2391,N_1861,N_1969);
or U2392 (N_2392,N_1963,N_1905);
nor U2393 (N_2393,N_1950,N_1919);
or U2394 (N_2394,N_1823,N_1758);
nor U2395 (N_2395,N_1701,N_1684);
or U2396 (N_2396,N_1858,N_1668);
and U2397 (N_2397,N_1753,N_1568);
nor U2398 (N_2398,N_1563,N_1710);
nor U2399 (N_2399,N_1703,N_1974);
and U2400 (N_2400,N_1577,N_1996);
and U2401 (N_2401,N_1978,N_1849);
nand U2402 (N_2402,N_1652,N_1623);
nor U2403 (N_2403,N_1980,N_1539);
xor U2404 (N_2404,N_1591,N_1547);
xnor U2405 (N_2405,N_1751,N_1690);
nor U2406 (N_2406,N_1659,N_1518);
or U2407 (N_2407,N_1890,N_1579);
nor U2408 (N_2408,N_1525,N_1815);
and U2409 (N_2409,N_1598,N_1996);
and U2410 (N_2410,N_1656,N_1970);
and U2411 (N_2411,N_1983,N_1634);
and U2412 (N_2412,N_1751,N_1534);
nor U2413 (N_2413,N_1999,N_1601);
or U2414 (N_2414,N_1744,N_1889);
nor U2415 (N_2415,N_1639,N_1590);
and U2416 (N_2416,N_1986,N_1533);
and U2417 (N_2417,N_1697,N_1724);
and U2418 (N_2418,N_1909,N_1664);
nand U2419 (N_2419,N_1553,N_1672);
or U2420 (N_2420,N_1998,N_1627);
or U2421 (N_2421,N_1534,N_1924);
nand U2422 (N_2422,N_1647,N_1714);
nand U2423 (N_2423,N_1846,N_1995);
or U2424 (N_2424,N_1711,N_1976);
nand U2425 (N_2425,N_1531,N_1713);
and U2426 (N_2426,N_1668,N_1516);
or U2427 (N_2427,N_1645,N_1801);
xor U2428 (N_2428,N_1869,N_1613);
and U2429 (N_2429,N_1948,N_1541);
nor U2430 (N_2430,N_1859,N_1919);
or U2431 (N_2431,N_1662,N_1632);
or U2432 (N_2432,N_1777,N_1799);
nor U2433 (N_2433,N_1881,N_1629);
nand U2434 (N_2434,N_1584,N_1582);
and U2435 (N_2435,N_1603,N_1587);
nor U2436 (N_2436,N_1516,N_1901);
nand U2437 (N_2437,N_1764,N_1655);
nand U2438 (N_2438,N_1791,N_1894);
or U2439 (N_2439,N_1546,N_1549);
and U2440 (N_2440,N_1849,N_1598);
and U2441 (N_2441,N_1847,N_1827);
xnor U2442 (N_2442,N_1750,N_1673);
or U2443 (N_2443,N_1960,N_1558);
and U2444 (N_2444,N_1900,N_1730);
xor U2445 (N_2445,N_1995,N_1978);
and U2446 (N_2446,N_1591,N_1957);
nand U2447 (N_2447,N_1786,N_1559);
nor U2448 (N_2448,N_1599,N_1754);
nand U2449 (N_2449,N_1931,N_1784);
nand U2450 (N_2450,N_1558,N_1527);
xnor U2451 (N_2451,N_1714,N_1985);
nand U2452 (N_2452,N_1629,N_1685);
and U2453 (N_2453,N_1544,N_1618);
and U2454 (N_2454,N_1593,N_1830);
nand U2455 (N_2455,N_1568,N_1791);
nor U2456 (N_2456,N_1791,N_1989);
nor U2457 (N_2457,N_1724,N_1749);
xnor U2458 (N_2458,N_1950,N_1676);
or U2459 (N_2459,N_1904,N_1967);
or U2460 (N_2460,N_1899,N_1578);
nand U2461 (N_2461,N_1967,N_1875);
nor U2462 (N_2462,N_1818,N_1962);
or U2463 (N_2463,N_1803,N_1892);
and U2464 (N_2464,N_1584,N_1580);
nand U2465 (N_2465,N_1815,N_1874);
nor U2466 (N_2466,N_1645,N_1877);
nor U2467 (N_2467,N_1892,N_1908);
xnor U2468 (N_2468,N_1701,N_1636);
and U2469 (N_2469,N_1525,N_1556);
nor U2470 (N_2470,N_1998,N_1565);
xnor U2471 (N_2471,N_1609,N_1595);
nand U2472 (N_2472,N_1712,N_1628);
or U2473 (N_2473,N_1966,N_1550);
and U2474 (N_2474,N_1512,N_1761);
nor U2475 (N_2475,N_1516,N_1698);
and U2476 (N_2476,N_1910,N_1964);
nor U2477 (N_2477,N_1546,N_1728);
nor U2478 (N_2478,N_1757,N_1723);
or U2479 (N_2479,N_1603,N_1558);
and U2480 (N_2480,N_1879,N_1829);
xor U2481 (N_2481,N_1985,N_1706);
nor U2482 (N_2482,N_1755,N_1684);
nand U2483 (N_2483,N_1875,N_1859);
and U2484 (N_2484,N_1841,N_1908);
xnor U2485 (N_2485,N_1967,N_1760);
xnor U2486 (N_2486,N_1600,N_1626);
nand U2487 (N_2487,N_1562,N_1984);
xor U2488 (N_2488,N_1934,N_1521);
xnor U2489 (N_2489,N_1843,N_1730);
nor U2490 (N_2490,N_1855,N_1768);
nor U2491 (N_2491,N_1655,N_1528);
and U2492 (N_2492,N_1969,N_1718);
xor U2493 (N_2493,N_1558,N_1982);
nand U2494 (N_2494,N_1954,N_1996);
nor U2495 (N_2495,N_1872,N_1632);
nand U2496 (N_2496,N_1845,N_1612);
and U2497 (N_2497,N_1899,N_1524);
nand U2498 (N_2498,N_1709,N_1745);
nand U2499 (N_2499,N_1517,N_1944);
xnor U2500 (N_2500,N_2262,N_2358);
nor U2501 (N_2501,N_2454,N_2410);
nand U2502 (N_2502,N_2020,N_2433);
and U2503 (N_2503,N_2055,N_2189);
nand U2504 (N_2504,N_2060,N_2079);
nor U2505 (N_2505,N_2125,N_2013);
nor U2506 (N_2506,N_2472,N_2187);
or U2507 (N_2507,N_2217,N_2077);
or U2508 (N_2508,N_2123,N_2219);
or U2509 (N_2509,N_2407,N_2299);
nand U2510 (N_2510,N_2283,N_2387);
and U2511 (N_2511,N_2302,N_2260);
nor U2512 (N_2512,N_2459,N_2203);
nand U2513 (N_2513,N_2300,N_2360);
nor U2514 (N_2514,N_2434,N_2478);
xor U2515 (N_2515,N_2267,N_2150);
xor U2516 (N_2516,N_2206,N_2422);
or U2517 (N_2517,N_2221,N_2258);
and U2518 (N_2518,N_2448,N_2265);
xnor U2519 (N_2519,N_2092,N_2313);
and U2520 (N_2520,N_2450,N_2185);
nor U2521 (N_2521,N_2320,N_2363);
xnor U2522 (N_2522,N_2132,N_2438);
nor U2523 (N_2523,N_2345,N_2366);
xor U2524 (N_2524,N_2172,N_2093);
or U2525 (N_2525,N_2115,N_2065);
nand U2526 (N_2526,N_2164,N_2034);
nor U2527 (N_2527,N_2086,N_2056);
or U2528 (N_2528,N_2044,N_2463);
xor U2529 (N_2529,N_2067,N_2229);
xnor U2530 (N_2530,N_2102,N_2310);
and U2531 (N_2531,N_2008,N_2073);
or U2532 (N_2532,N_2257,N_2404);
or U2533 (N_2533,N_2235,N_2452);
xor U2534 (N_2534,N_2242,N_2182);
and U2535 (N_2535,N_2490,N_2054);
nor U2536 (N_2536,N_2402,N_2100);
nor U2537 (N_2537,N_2499,N_2066);
nor U2538 (N_2538,N_2352,N_2351);
nand U2539 (N_2539,N_2367,N_2427);
and U2540 (N_2540,N_2290,N_2280);
nand U2541 (N_2541,N_2117,N_2035);
nor U2542 (N_2542,N_2089,N_2443);
nand U2543 (N_2543,N_2070,N_2451);
or U2544 (N_2544,N_2471,N_2425);
and U2545 (N_2545,N_2482,N_2250);
nand U2546 (N_2546,N_2080,N_2133);
nand U2547 (N_2547,N_2043,N_2173);
or U2548 (N_2548,N_2446,N_2480);
and U2549 (N_2549,N_2096,N_2292);
and U2550 (N_2550,N_2322,N_2042);
and U2551 (N_2551,N_2255,N_2460);
nor U2552 (N_2552,N_2435,N_2406);
or U2553 (N_2553,N_2312,N_2160);
or U2554 (N_2554,N_2445,N_2147);
nand U2555 (N_2555,N_2101,N_2266);
xor U2556 (N_2556,N_2447,N_2362);
nand U2557 (N_2557,N_2186,N_2168);
nand U2558 (N_2558,N_2212,N_2201);
or U2559 (N_2559,N_2076,N_2138);
and U2560 (N_2560,N_2315,N_2276);
or U2561 (N_2561,N_2491,N_2364);
nand U2562 (N_2562,N_2475,N_2399);
and U2563 (N_2563,N_2074,N_2423);
xor U2564 (N_2564,N_2375,N_2090);
nand U2565 (N_2565,N_2036,N_2294);
xor U2566 (N_2566,N_2129,N_2325);
nor U2567 (N_2567,N_2139,N_2296);
or U2568 (N_2568,N_2208,N_2327);
and U2569 (N_2569,N_2304,N_2154);
nand U2570 (N_2570,N_2050,N_2205);
nor U2571 (N_2571,N_2347,N_2157);
nand U2572 (N_2572,N_2025,N_2441);
or U2573 (N_2573,N_2116,N_2062);
xnor U2574 (N_2574,N_2226,N_2316);
nor U2575 (N_2575,N_2314,N_2383);
and U2576 (N_2576,N_2477,N_2069);
xnor U2577 (N_2577,N_2377,N_2061);
nor U2578 (N_2578,N_2468,N_2330);
nor U2579 (N_2579,N_2493,N_2151);
nor U2580 (N_2580,N_2017,N_2419);
nor U2581 (N_2581,N_2455,N_2112);
or U2582 (N_2582,N_2376,N_2024);
xnor U2583 (N_2583,N_2097,N_2128);
or U2584 (N_2584,N_2122,N_2002);
and U2585 (N_2585,N_2174,N_2071);
and U2586 (N_2586,N_2251,N_2195);
and U2587 (N_2587,N_2344,N_2170);
and U2588 (N_2588,N_2457,N_2489);
xor U2589 (N_2589,N_2119,N_2078);
or U2590 (N_2590,N_2428,N_2289);
nand U2591 (N_2591,N_2403,N_2485);
nand U2592 (N_2592,N_2130,N_2311);
nand U2593 (N_2593,N_2113,N_2405);
nor U2594 (N_2594,N_2094,N_2033);
or U2595 (N_2595,N_2487,N_2194);
nand U2596 (N_2596,N_2385,N_2297);
or U2597 (N_2597,N_2210,N_2177);
xor U2598 (N_2598,N_2335,N_2496);
or U2599 (N_2599,N_2497,N_2264);
and U2600 (N_2600,N_2368,N_2343);
or U2601 (N_2601,N_2396,N_2091);
or U2602 (N_2602,N_2253,N_2437);
nor U2603 (N_2603,N_2488,N_2254);
or U2604 (N_2604,N_2243,N_2340);
or U2605 (N_2605,N_2167,N_2301);
nor U2606 (N_2606,N_2287,N_2007);
xor U2607 (N_2607,N_2395,N_2233);
or U2608 (N_2608,N_2326,N_2436);
nor U2609 (N_2609,N_2373,N_2381);
nand U2610 (N_2610,N_2412,N_2269);
or U2611 (N_2611,N_2430,N_2191);
nand U2612 (N_2612,N_2021,N_2059);
xor U2613 (N_2613,N_2222,N_2409);
nor U2614 (N_2614,N_2286,N_2214);
nand U2615 (N_2615,N_2088,N_2004);
and U2616 (N_2616,N_2440,N_2204);
and U2617 (N_2617,N_2388,N_2481);
nand U2618 (N_2618,N_2279,N_2458);
and U2619 (N_2619,N_2126,N_2483);
xor U2620 (N_2620,N_2275,N_2389);
nor U2621 (N_2621,N_2291,N_2051);
nor U2622 (N_2622,N_2328,N_2228);
nand U2623 (N_2623,N_2336,N_2426);
and U2624 (N_2624,N_2188,N_2317);
and U2625 (N_2625,N_2259,N_2469);
or U2626 (N_2626,N_2161,N_2215);
or U2627 (N_2627,N_2282,N_2393);
and U2628 (N_2628,N_2365,N_2107);
xnor U2629 (N_2629,N_2324,N_2057);
and U2630 (N_2630,N_2152,N_2048);
xnor U2631 (N_2631,N_2005,N_2019);
nor U2632 (N_2632,N_2361,N_2156);
and U2633 (N_2633,N_2305,N_2099);
and U2634 (N_2634,N_2010,N_2196);
xnor U2635 (N_2635,N_2081,N_2342);
and U2636 (N_2636,N_2415,N_2391);
xnor U2637 (N_2637,N_2307,N_2431);
nor U2638 (N_2638,N_2084,N_2369);
nor U2639 (N_2639,N_2323,N_2199);
and U2640 (N_2640,N_2319,N_2207);
and U2641 (N_2641,N_2232,N_2417);
xor U2642 (N_2642,N_2338,N_2023);
or U2643 (N_2643,N_2163,N_2392);
or U2644 (N_2644,N_2353,N_2153);
nor U2645 (N_2645,N_2142,N_2348);
nor U2646 (N_2646,N_2148,N_2394);
nor U2647 (N_2647,N_2047,N_2244);
nand U2648 (N_2648,N_2137,N_2144);
or U2649 (N_2649,N_2141,N_2041);
nand U2650 (N_2650,N_2341,N_2045);
and U2651 (N_2651,N_2379,N_2064);
xnor U2652 (N_2652,N_2072,N_2155);
and U2653 (N_2653,N_2176,N_2237);
or U2654 (N_2654,N_2408,N_2009);
or U2655 (N_2655,N_2098,N_2183);
or U2656 (N_2656,N_2052,N_2498);
xnor U2657 (N_2657,N_2135,N_2223);
xnor U2658 (N_2658,N_2018,N_2241);
nor U2659 (N_2659,N_2295,N_2046);
nor U2660 (N_2660,N_2334,N_2467);
and U2661 (N_2661,N_2382,N_2053);
nor U2662 (N_2662,N_2306,N_2256);
or U2663 (N_2663,N_2439,N_2236);
xor U2664 (N_2664,N_2166,N_2416);
nand U2665 (N_2665,N_2397,N_2401);
and U2666 (N_2666,N_2372,N_2424);
nand U2667 (N_2667,N_2145,N_2285);
nor U2668 (N_2668,N_2281,N_2022);
or U2669 (N_2669,N_2238,N_2095);
or U2670 (N_2670,N_2308,N_2003);
xor U2671 (N_2671,N_2121,N_2371);
and U2672 (N_2672,N_2085,N_2252);
and U2673 (N_2673,N_2421,N_2227);
or U2674 (N_2674,N_2209,N_2037);
xnor U2675 (N_2675,N_2271,N_2136);
nand U2676 (N_2676,N_2058,N_2380);
nor U2677 (N_2677,N_2465,N_2225);
nor U2678 (N_2678,N_2479,N_2159);
xor U2679 (N_2679,N_2026,N_2240);
or U2680 (N_2680,N_2261,N_2087);
xor U2681 (N_2681,N_2106,N_2231);
and U2682 (N_2682,N_2200,N_2202);
nor U2683 (N_2683,N_2143,N_2337);
xor U2684 (N_2684,N_2263,N_2198);
nor U2685 (N_2685,N_2246,N_2211);
xnor U2686 (N_2686,N_2103,N_2321);
nand U2687 (N_2687,N_2378,N_2179);
nor U2688 (N_2688,N_2027,N_2015);
or U2689 (N_2689,N_2175,N_2278);
xnor U2690 (N_2690,N_2429,N_2118);
nand U2691 (N_2691,N_2068,N_2356);
nand U2692 (N_2692,N_2350,N_2268);
nand U2693 (N_2693,N_2014,N_2359);
and U2694 (N_2694,N_2354,N_2171);
xnor U2695 (N_2695,N_2470,N_2131);
nand U2696 (N_2696,N_2104,N_2462);
nor U2697 (N_2697,N_2111,N_2213);
nand U2698 (N_2698,N_2032,N_2384);
nand U2699 (N_2699,N_2184,N_2190);
nand U2700 (N_2700,N_2464,N_2030);
nor U2701 (N_2701,N_2247,N_2414);
and U2702 (N_2702,N_2218,N_2432);
nand U2703 (N_2703,N_2109,N_2331);
nor U2704 (N_2704,N_2110,N_2355);
and U2705 (N_2705,N_2063,N_2105);
or U2706 (N_2706,N_2273,N_2230);
nand U2707 (N_2707,N_2333,N_2473);
xnor U2708 (N_2708,N_2245,N_2220);
or U2709 (N_2709,N_2083,N_2474);
nor U2710 (N_2710,N_2461,N_2332);
xor U2711 (N_2711,N_2274,N_2000);
or U2712 (N_2712,N_2249,N_2040);
and U2713 (N_2713,N_2012,N_2492);
or U2714 (N_2714,N_2288,N_2272);
or U2715 (N_2715,N_2400,N_2169);
or U2716 (N_2716,N_2016,N_2277);
and U2717 (N_2717,N_2039,N_2495);
xor U2718 (N_2718,N_2456,N_2049);
or U2719 (N_2719,N_2270,N_2357);
and U2720 (N_2720,N_2162,N_2134);
or U2721 (N_2721,N_2309,N_2216);
and U2722 (N_2722,N_2390,N_2158);
nor U2723 (N_2723,N_2284,N_2192);
nand U2724 (N_2724,N_2413,N_2370);
xor U2725 (N_2725,N_2120,N_2075);
or U2726 (N_2726,N_2082,N_2476);
xor U2727 (N_2727,N_2453,N_2165);
or U2728 (N_2728,N_2374,N_2146);
nor U2729 (N_2729,N_2418,N_2114);
or U2730 (N_2730,N_2124,N_2346);
and U2731 (N_2731,N_2180,N_2140);
xor U2732 (N_2732,N_2149,N_2293);
nor U2733 (N_2733,N_2442,N_2127);
xor U2734 (N_2734,N_2494,N_2486);
xor U2735 (N_2735,N_2349,N_2318);
and U2736 (N_2736,N_2234,N_2239);
nand U2737 (N_2737,N_2444,N_2484);
and U2738 (N_2738,N_2466,N_2181);
and U2739 (N_2739,N_2178,N_2031);
nor U2740 (N_2740,N_2029,N_2197);
or U2741 (N_2741,N_2303,N_2011);
nand U2742 (N_2742,N_2006,N_2398);
nand U2743 (N_2743,N_2329,N_2224);
nand U2744 (N_2744,N_2339,N_2449);
or U2745 (N_2745,N_2386,N_2001);
nor U2746 (N_2746,N_2193,N_2248);
xnor U2747 (N_2747,N_2038,N_2411);
nand U2748 (N_2748,N_2108,N_2298);
nand U2749 (N_2749,N_2420,N_2028);
xor U2750 (N_2750,N_2311,N_2083);
or U2751 (N_2751,N_2420,N_2075);
nor U2752 (N_2752,N_2435,N_2245);
or U2753 (N_2753,N_2409,N_2396);
xnor U2754 (N_2754,N_2160,N_2451);
and U2755 (N_2755,N_2386,N_2037);
and U2756 (N_2756,N_2399,N_2410);
nor U2757 (N_2757,N_2371,N_2066);
nor U2758 (N_2758,N_2199,N_2427);
xnor U2759 (N_2759,N_2239,N_2462);
xnor U2760 (N_2760,N_2344,N_2354);
nor U2761 (N_2761,N_2487,N_2132);
xor U2762 (N_2762,N_2121,N_2264);
or U2763 (N_2763,N_2307,N_2347);
and U2764 (N_2764,N_2195,N_2167);
xnor U2765 (N_2765,N_2305,N_2116);
xor U2766 (N_2766,N_2200,N_2019);
nand U2767 (N_2767,N_2265,N_2100);
xor U2768 (N_2768,N_2280,N_2010);
and U2769 (N_2769,N_2051,N_2146);
nand U2770 (N_2770,N_2369,N_2119);
or U2771 (N_2771,N_2321,N_2094);
nor U2772 (N_2772,N_2058,N_2228);
xnor U2773 (N_2773,N_2151,N_2023);
xor U2774 (N_2774,N_2289,N_2370);
or U2775 (N_2775,N_2105,N_2239);
or U2776 (N_2776,N_2423,N_2475);
and U2777 (N_2777,N_2347,N_2356);
xnor U2778 (N_2778,N_2222,N_2075);
nand U2779 (N_2779,N_2044,N_2279);
nand U2780 (N_2780,N_2315,N_2022);
or U2781 (N_2781,N_2351,N_2179);
and U2782 (N_2782,N_2369,N_2163);
and U2783 (N_2783,N_2474,N_2027);
and U2784 (N_2784,N_2286,N_2469);
and U2785 (N_2785,N_2256,N_2112);
or U2786 (N_2786,N_2327,N_2226);
or U2787 (N_2787,N_2114,N_2134);
xnor U2788 (N_2788,N_2429,N_2201);
xnor U2789 (N_2789,N_2185,N_2215);
xnor U2790 (N_2790,N_2132,N_2320);
nor U2791 (N_2791,N_2139,N_2149);
xnor U2792 (N_2792,N_2039,N_2151);
or U2793 (N_2793,N_2421,N_2171);
nor U2794 (N_2794,N_2094,N_2036);
nor U2795 (N_2795,N_2138,N_2033);
xnor U2796 (N_2796,N_2474,N_2330);
xnor U2797 (N_2797,N_2018,N_2199);
or U2798 (N_2798,N_2329,N_2165);
xnor U2799 (N_2799,N_2290,N_2446);
nand U2800 (N_2800,N_2492,N_2270);
and U2801 (N_2801,N_2003,N_2436);
and U2802 (N_2802,N_2091,N_2293);
xnor U2803 (N_2803,N_2229,N_2460);
xnor U2804 (N_2804,N_2396,N_2323);
xor U2805 (N_2805,N_2115,N_2477);
xor U2806 (N_2806,N_2100,N_2070);
nor U2807 (N_2807,N_2465,N_2383);
or U2808 (N_2808,N_2325,N_2348);
xnor U2809 (N_2809,N_2172,N_2443);
nand U2810 (N_2810,N_2463,N_2223);
nor U2811 (N_2811,N_2375,N_2236);
nand U2812 (N_2812,N_2190,N_2043);
nor U2813 (N_2813,N_2214,N_2213);
or U2814 (N_2814,N_2177,N_2034);
xnor U2815 (N_2815,N_2207,N_2270);
or U2816 (N_2816,N_2458,N_2120);
or U2817 (N_2817,N_2461,N_2477);
nor U2818 (N_2818,N_2494,N_2241);
xor U2819 (N_2819,N_2360,N_2482);
nor U2820 (N_2820,N_2390,N_2296);
and U2821 (N_2821,N_2439,N_2271);
nor U2822 (N_2822,N_2219,N_2380);
nor U2823 (N_2823,N_2444,N_2421);
nand U2824 (N_2824,N_2350,N_2057);
xnor U2825 (N_2825,N_2217,N_2254);
xnor U2826 (N_2826,N_2413,N_2081);
or U2827 (N_2827,N_2445,N_2066);
and U2828 (N_2828,N_2187,N_2434);
and U2829 (N_2829,N_2013,N_2051);
or U2830 (N_2830,N_2234,N_2208);
and U2831 (N_2831,N_2141,N_2200);
nand U2832 (N_2832,N_2217,N_2387);
and U2833 (N_2833,N_2200,N_2216);
nor U2834 (N_2834,N_2092,N_2134);
nor U2835 (N_2835,N_2475,N_2323);
xnor U2836 (N_2836,N_2343,N_2108);
nand U2837 (N_2837,N_2017,N_2391);
or U2838 (N_2838,N_2140,N_2079);
xor U2839 (N_2839,N_2426,N_2313);
xor U2840 (N_2840,N_2245,N_2338);
nand U2841 (N_2841,N_2268,N_2053);
and U2842 (N_2842,N_2213,N_2339);
and U2843 (N_2843,N_2261,N_2310);
and U2844 (N_2844,N_2415,N_2063);
and U2845 (N_2845,N_2172,N_2438);
or U2846 (N_2846,N_2443,N_2138);
nand U2847 (N_2847,N_2472,N_2274);
xor U2848 (N_2848,N_2343,N_2100);
nand U2849 (N_2849,N_2228,N_2104);
or U2850 (N_2850,N_2403,N_2057);
xnor U2851 (N_2851,N_2459,N_2463);
xor U2852 (N_2852,N_2423,N_2033);
nor U2853 (N_2853,N_2170,N_2192);
xnor U2854 (N_2854,N_2177,N_2347);
and U2855 (N_2855,N_2141,N_2284);
nor U2856 (N_2856,N_2230,N_2041);
and U2857 (N_2857,N_2310,N_2469);
and U2858 (N_2858,N_2442,N_2426);
xor U2859 (N_2859,N_2301,N_2169);
nor U2860 (N_2860,N_2150,N_2368);
nor U2861 (N_2861,N_2067,N_2469);
nand U2862 (N_2862,N_2111,N_2253);
and U2863 (N_2863,N_2155,N_2224);
and U2864 (N_2864,N_2297,N_2387);
and U2865 (N_2865,N_2097,N_2261);
or U2866 (N_2866,N_2323,N_2316);
xnor U2867 (N_2867,N_2309,N_2008);
xnor U2868 (N_2868,N_2426,N_2063);
nor U2869 (N_2869,N_2181,N_2035);
or U2870 (N_2870,N_2351,N_2435);
and U2871 (N_2871,N_2412,N_2205);
and U2872 (N_2872,N_2085,N_2144);
xor U2873 (N_2873,N_2124,N_2181);
nor U2874 (N_2874,N_2246,N_2488);
nor U2875 (N_2875,N_2142,N_2264);
and U2876 (N_2876,N_2440,N_2292);
xor U2877 (N_2877,N_2294,N_2095);
nor U2878 (N_2878,N_2394,N_2426);
and U2879 (N_2879,N_2019,N_2376);
or U2880 (N_2880,N_2194,N_2163);
or U2881 (N_2881,N_2004,N_2209);
nor U2882 (N_2882,N_2107,N_2233);
xor U2883 (N_2883,N_2247,N_2098);
nor U2884 (N_2884,N_2251,N_2269);
or U2885 (N_2885,N_2084,N_2208);
and U2886 (N_2886,N_2210,N_2230);
or U2887 (N_2887,N_2170,N_2117);
nand U2888 (N_2888,N_2002,N_2227);
or U2889 (N_2889,N_2301,N_2353);
and U2890 (N_2890,N_2282,N_2016);
nand U2891 (N_2891,N_2134,N_2481);
nor U2892 (N_2892,N_2252,N_2134);
or U2893 (N_2893,N_2006,N_2141);
xor U2894 (N_2894,N_2036,N_2483);
or U2895 (N_2895,N_2020,N_2280);
nand U2896 (N_2896,N_2465,N_2174);
nand U2897 (N_2897,N_2294,N_2428);
nor U2898 (N_2898,N_2264,N_2356);
and U2899 (N_2899,N_2084,N_2370);
nand U2900 (N_2900,N_2478,N_2344);
or U2901 (N_2901,N_2074,N_2139);
nand U2902 (N_2902,N_2435,N_2434);
and U2903 (N_2903,N_2186,N_2167);
xnor U2904 (N_2904,N_2383,N_2071);
and U2905 (N_2905,N_2460,N_2083);
and U2906 (N_2906,N_2069,N_2377);
or U2907 (N_2907,N_2379,N_2305);
xor U2908 (N_2908,N_2278,N_2126);
and U2909 (N_2909,N_2474,N_2128);
or U2910 (N_2910,N_2268,N_2153);
or U2911 (N_2911,N_2205,N_2383);
and U2912 (N_2912,N_2177,N_2455);
xor U2913 (N_2913,N_2330,N_2197);
nor U2914 (N_2914,N_2215,N_2239);
and U2915 (N_2915,N_2485,N_2323);
nor U2916 (N_2916,N_2179,N_2358);
nand U2917 (N_2917,N_2433,N_2432);
nand U2918 (N_2918,N_2398,N_2498);
or U2919 (N_2919,N_2053,N_2380);
xnor U2920 (N_2920,N_2148,N_2009);
xor U2921 (N_2921,N_2283,N_2459);
xor U2922 (N_2922,N_2358,N_2456);
xor U2923 (N_2923,N_2410,N_2204);
nand U2924 (N_2924,N_2478,N_2018);
and U2925 (N_2925,N_2056,N_2352);
nand U2926 (N_2926,N_2369,N_2223);
nand U2927 (N_2927,N_2413,N_2270);
xnor U2928 (N_2928,N_2200,N_2468);
nor U2929 (N_2929,N_2017,N_2491);
and U2930 (N_2930,N_2380,N_2479);
and U2931 (N_2931,N_2452,N_2271);
xor U2932 (N_2932,N_2117,N_2230);
nor U2933 (N_2933,N_2210,N_2204);
or U2934 (N_2934,N_2023,N_2207);
nand U2935 (N_2935,N_2018,N_2438);
xnor U2936 (N_2936,N_2210,N_2187);
xor U2937 (N_2937,N_2176,N_2345);
nand U2938 (N_2938,N_2175,N_2131);
xor U2939 (N_2939,N_2382,N_2156);
xor U2940 (N_2940,N_2383,N_2069);
nor U2941 (N_2941,N_2158,N_2012);
or U2942 (N_2942,N_2021,N_2010);
xnor U2943 (N_2943,N_2222,N_2362);
xor U2944 (N_2944,N_2395,N_2446);
and U2945 (N_2945,N_2405,N_2186);
xor U2946 (N_2946,N_2141,N_2153);
or U2947 (N_2947,N_2341,N_2307);
xnor U2948 (N_2948,N_2372,N_2405);
and U2949 (N_2949,N_2092,N_2475);
xor U2950 (N_2950,N_2084,N_2336);
xor U2951 (N_2951,N_2498,N_2486);
xor U2952 (N_2952,N_2335,N_2155);
and U2953 (N_2953,N_2116,N_2012);
nand U2954 (N_2954,N_2110,N_2242);
or U2955 (N_2955,N_2103,N_2457);
nand U2956 (N_2956,N_2262,N_2016);
or U2957 (N_2957,N_2001,N_2236);
or U2958 (N_2958,N_2136,N_2216);
or U2959 (N_2959,N_2181,N_2162);
or U2960 (N_2960,N_2276,N_2491);
nor U2961 (N_2961,N_2453,N_2413);
and U2962 (N_2962,N_2448,N_2032);
or U2963 (N_2963,N_2245,N_2349);
and U2964 (N_2964,N_2378,N_2224);
and U2965 (N_2965,N_2277,N_2261);
and U2966 (N_2966,N_2358,N_2193);
or U2967 (N_2967,N_2216,N_2363);
xnor U2968 (N_2968,N_2240,N_2379);
or U2969 (N_2969,N_2207,N_2329);
or U2970 (N_2970,N_2084,N_2186);
nor U2971 (N_2971,N_2268,N_2023);
nand U2972 (N_2972,N_2210,N_2147);
nor U2973 (N_2973,N_2124,N_2057);
nand U2974 (N_2974,N_2481,N_2092);
or U2975 (N_2975,N_2439,N_2111);
xnor U2976 (N_2976,N_2403,N_2494);
or U2977 (N_2977,N_2360,N_2218);
or U2978 (N_2978,N_2028,N_2022);
and U2979 (N_2979,N_2065,N_2489);
or U2980 (N_2980,N_2154,N_2415);
or U2981 (N_2981,N_2118,N_2386);
nor U2982 (N_2982,N_2376,N_2364);
and U2983 (N_2983,N_2007,N_2381);
nand U2984 (N_2984,N_2148,N_2390);
or U2985 (N_2985,N_2292,N_2107);
xor U2986 (N_2986,N_2334,N_2122);
nor U2987 (N_2987,N_2195,N_2033);
nand U2988 (N_2988,N_2340,N_2165);
nor U2989 (N_2989,N_2197,N_2282);
or U2990 (N_2990,N_2402,N_2369);
or U2991 (N_2991,N_2177,N_2375);
xnor U2992 (N_2992,N_2292,N_2275);
nor U2993 (N_2993,N_2240,N_2325);
nand U2994 (N_2994,N_2253,N_2376);
nor U2995 (N_2995,N_2429,N_2217);
or U2996 (N_2996,N_2180,N_2002);
and U2997 (N_2997,N_2002,N_2319);
xnor U2998 (N_2998,N_2032,N_2295);
xnor U2999 (N_2999,N_2215,N_2269);
and U3000 (N_3000,N_2939,N_2770);
and U3001 (N_3001,N_2993,N_2568);
nor U3002 (N_3002,N_2859,N_2681);
and U3003 (N_3003,N_2744,N_2669);
xor U3004 (N_3004,N_2827,N_2591);
or U3005 (N_3005,N_2559,N_2773);
and U3006 (N_3006,N_2960,N_2605);
xnor U3007 (N_3007,N_2961,N_2587);
nor U3008 (N_3008,N_2600,N_2740);
and U3009 (N_3009,N_2851,N_2572);
or U3010 (N_3010,N_2588,N_2604);
nand U3011 (N_3011,N_2837,N_2517);
xor U3012 (N_3012,N_2713,N_2875);
nand U3013 (N_3013,N_2627,N_2545);
nor U3014 (N_3014,N_2916,N_2644);
nor U3015 (N_3015,N_2509,N_2979);
nand U3016 (N_3016,N_2535,N_2743);
and U3017 (N_3017,N_2716,N_2776);
xor U3018 (N_3018,N_2641,N_2595);
nand U3019 (N_3019,N_2552,N_2758);
or U3020 (N_3020,N_2786,N_2684);
nor U3021 (N_3021,N_2699,N_2735);
nand U3022 (N_3022,N_2694,N_2696);
xor U3023 (N_3023,N_2935,N_2668);
nor U3024 (N_3024,N_2645,N_2687);
nand U3025 (N_3025,N_2823,N_2557);
xnor U3026 (N_3026,N_2998,N_2531);
or U3027 (N_3027,N_2819,N_2755);
or U3028 (N_3028,N_2825,N_2788);
nor U3029 (N_3029,N_2880,N_2522);
nand U3030 (N_3030,N_2863,N_2529);
xor U3031 (N_3031,N_2843,N_2726);
and U3032 (N_3032,N_2822,N_2629);
xor U3033 (N_3033,N_2594,N_2611);
xor U3034 (N_3034,N_2577,N_2897);
xor U3035 (N_3035,N_2760,N_2962);
and U3036 (N_3036,N_2796,N_2781);
and U3037 (N_3037,N_2723,N_2797);
nor U3038 (N_3038,N_2861,N_2942);
xor U3039 (N_3039,N_2907,N_2849);
nor U3040 (N_3040,N_2757,N_2515);
nand U3041 (N_3041,N_2651,N_2637);
nand U3042 (N_3042,N_2632,N_2976);
or U3043 (N_3043,N_2834,N_2556);
nor U3044 (N_3044,N_2769,N_2959);
nor U3045 (N_3045,N_2938,N_2877);
nand U3046 (N_3046,N_2724,N_2874);
and U3047 (N_3047,N_2670,N_2663);
and U3048 (N_3048,N_2898,N_2840);
nor U3049 (N_3049,N_2656,N_2904);
nand U3050 (N_3050,N_2816,N_2900);
nor U3051 (N_3051,N_2538,N_2844);
xor U3052 (N_3052,N_2860,N_2682);
nor U3053 (N_3053,N_2782,N_2934);
nor U3054 (N_3054,N_2799,N_2737);
xnor U3055 (N_3055,N_2858,N_2665);
or U3056 (N_3056,N_2583,N_2746);
nor U3057 (N_3057,N_2566,N_2905);
or U3058 (N_3058,N_2547,N_2745);
and U3059 (N_3059,N_2866,N_2933);
and U3060 (N_3060,N_2650,N_2625);
nand U3061 (N_3061,N_2853,N_2731);
nor U3062 (N_3062,N_2734,N_2852);
nand U3063 (N_3063,N_2946,N_2766);
xor U3064 (N_3064,N_2884,N_2977);
or U3065 (N_3065,N_2544,N_2995);
nor U3066 (N_3066,N_2765,N_2963);
and U3067 (N_3067,N_2764,N_2541);
or U3068 (N_3068,N_2865,N_2653);
or U3069 (N_3069,N_2831,N_2708);
or U3070 (N_3070,N_2753,N_2623);
and U3071 (N_3071,N_2862,N_2599);
nor U3072 (N_3072,N_2619,N_2864);
or U3073 (N_3073,N_2748,N_2752);
or U3074 (N_3074,N_2972,N_2542);
nand U3075 (N_3075,N_2771,N_2525);
xnor U3076 (N_3076,N_2881,N_2915);
nand U3077 (N_3077,N_2514,N_2536);
nor U3078 (N_3078,N_2673,N_2603);
and U3079 (N_3079,N_2879,N_2891);
or U3080 (N_3080,N_2922,N_2917);
or U3081 (N_3081,N_2944,N_2574);
nand U3082 (N_3082,N_2551,N_2826);
and U3083 (N_3083,N_2793,N_2503);
nor U3084 (N_3084,N_2507,N_2919);
nand U3085 (N_3085,N_2792,N_2582);
or U3086 (N_3086,N_2839,N_2794);
nor U3087 (N_3087,N_2947,N_2948);
xnor U3088 (N_3088,N_2675,N_2848);
or U3089 (N_3089,N_2523,N_2689);
and U3090 (N_3090,N_2589,N_2506);
xor U3091 (N_3091,N_2512,N_2520);
and U3092 (N_3092,N_2980,N_2911);
xnor U3093 (N_3093,N_2832,N_2667);
nor U3094 (N_3094,N_2649,N_2931);
nor U3095 (N_3095,N_2672,N_2607);
or U3096 (N_3096,N_2937,N_2890);
and U3097 (N_3097,N_2612,N_2569);
and U3098 (N_3098,N_2913,N_2666);
and U3099 (N_3099,N_2883,N_2690);
and U3100 (N_3100,N_2876,N_2870);
nor U3101 (N_3101,N_2856,N_2996);
xor U3102 (N_3102,N_2558,N_2842);
xnor U3103 (N_3103,N_2854,N_2957);
xor U3104 (N_3104,N_2534,N_2945);
nand U3105 (N_3105,N_2759,N_2941);
and U3106 (N_3106,N_2953,N_2721);
nor U3107 (N_3107,N_2710,N_2973);
nand U3108 (N_3108,N_2969,N_2958);
xnor U3109 (N_3109,N_2789,N_2887);
and U3110 (N_3110,N_2553,N_2648);
nor U3111 (N_3111,N_2732,N_2562);
or U3112 (N_3112,N_2626,N_2555);
xor U3113 (N_3113,N_2817,N_2994);
nor U3114 (N_3114,N_2927,N_2560);
xnor U3115 (N_3115,N_2809,N_2728);
and U3116 (N_3116,N_2787,N_2571);
or U3117 (N_3117,N_2711,N_2833);
nor U3118 (N_3118,N_2992,N_2878);
xor U3119 (N_3119,N_2808,N_2775);
or U3120 (N_3120,N_2655,N_2680);
xnor U3121 (N_3121,N_2585,N_2803);
and U3122 (N_3122,N_2873,N_2688);
nor U3123 (N_3123,N_2700,N_2754);
nand U3124 (N_3124,N_2633,N_2530);
and U3125 (N_3125,N_2780,N_2621);
nor U3126 (N_3126,N_2750,N_2950);
nor U3127 (N_3127,N_2986,N_2722);
and U3128 (N_3128,N_2642,N_2964);
nor U3129 (N_3129,N_2624,N_2872);
nand U3130 (N_3130,N_2657,N_2918);
or U3131 (N_3131,N_2504,N_2906);
nor U3132 (N_3132,N_2970,N_2593);
nand U3133 (N_3133,N_2967,N_2747);
nand U3134 (N_3134,N_2838,N_2899);
or U3135 (N_3135,N_2749,N_2845);
xnor U3136 (N_3136,N_2867,N_2889);
nand U3137 (N_3137,N_2615,N_2762);
nand U3138 (N_3138,N_2617,N_2791);
or U3139 (N_3139,N_2524,N_2982);
nand U3140 (N_3140,N_2988,N_2691);
nor U3141 (N_3141,N_2850,N_2736);
nor U3142 (N_3142,N_2720,N_2955);
nor U3143 (N_3143,N_2609,N_2614);
nor U3144 (N_3144,N_2903,N_2601);
and U3145 (N_3145,N_2698,N_2701);
xnor U3146 (N_3146,N_2725,N_2990);
nor U3147 (N_3147,N_2705,N_2800);
or U3148 (N_3148,N_2802,N_2868);
or U3149 (N_3149,N_2706,N_2886);
nand U3150 (N_3150,N_2991,N_2707);
xnor U3151 (N_3151,N_2608,N_2613);
xor U3152 (N_3152,N_2968,N_2533);
nor U3153 (N_3153,N_2638,N_2719);
xor U3154 (N_3154,N_2679,N_2767);
and U3155 (N_3155,N_2703,N_2954);
nor U3156 (N_3156,N_2636,N_2510);
nand U3157 (N_3157,N_2590,N_2567);
nand U3158 (N_3158,N_2674,N_2661);
nor U3159 (N_3159,N_2527,N_2761);
xor U3160 (N_3160,N_2902,N_2981);
nor U3161 (N_3161,N_2561,N_2662);
xnor U3162 (N_3162,N_2597,N_2932);
xnor U3163 (N_3163,N_2717,N_2565);
nand U3164 (N_3164,N_2584,N_2885);
nor U3165 (N_3165,N_2807,N_2974);
xnor U3166 (N_3166,N_2810,N_2631);
nand U3167 (N_3167,N_2686,N_2622);
nor U3168 (N_3168,N_2936,N_2778);
or U3169 (N_3169,N_2965,N_2580);
nand U3170 (N_3170,N_2829,N_2537);
nand U3171 (N_3171,N_2596,N_2824);
nor U3172 (N_3172,N_2804,N_2893);
nor U3173 (N_3173,N_2949,N_2820);
xor U3174 (N_3174,N_2573,N_2830);
or U3175 (N_3175,N_2846,N_2501);
nand U3176 (N_3176,N_2579,N_2575);
xor U3177 (N_3177,N_2664,N_2586);
or U3178 (N_3178,N_2628,N_2930);
or U3179 (N_3179,N_2733,N_2805);
or U3180 (N_3180,N_2882,N_2634);
or U3181 (N_3181,N_2521,N_2836);
nor U3182 (N_3182,N_2801,N_2772);
or U3183 (N_3183,N_2598,N_2928);
nand U3184 (N_3184,N_2659,N_2654);
and U3185 (N_3185,N_2847,N_2639);
xor U3186 (N_3186,N_2540,N_2790);
or U3187 (N_3187,N_2564,N_2539);
or U3188 (N_3188,N_2971,N_2806);
nor U3189 (N_3189,N_2896,N_2606);
nor U3190 (N_3190,N_2989,N_2795);
nor U3191 (N_3191,N_2502,N_2923);
xnor U3192 (N_3192,N_2841,N_2618);
xor U3193 (N_3193,N_2563,N_2500);
or U3194 (N_3194,N_2511,N_2813);
nor U3195 (N_3195,N_2695,N_2652);
xor U3196 (N_3196,N_2951,N_2643);
or U3197 (N_3197,N_2742,N_2718);
nand U3198 (N_3198,N_2818,N_2901);
and U3199 (N_3199,N_2578,N_2678);
nand U3200 (N_3200,N_2894,N_2798);
xnor U3201 (N_3201,N_2895,N_2549);
nor U3202 (N_3202,N_2784,N_2943);
nor U3203 (N_3203,N_2985,N_2821);
nor U3204 (N_3204,N_2581,N_2756);
and U3205 (N_3205,N_2676,N_2857);
xor U3206 (N_3206,N_2871,N_2739);
or U3207 (N_3207,N_2774,N_2620);
xor U3208 (N_3208,N_2925,N_2812);
nand U3209 (N_3209,N_2909,N_2546);
xor U3210 (N_3210,N_2912,N_2592);
or U3211 (N_3211,N_2671,N_2727);
or U3212 (N_3212,N_2602,N_2630);
or U3213 (N_3213,N_2814,N_2978);
xnor U3214 (N_3214,N_2576,N_2997);
nor U3215 (N_3215,N_2677,N_2526);
and U3216 (N_3216,N_2516,N_2888);
or U3217 (N_3217,N_2685,N_2712);
nand U3218 (N_3218,N_2751,N_2983);
or U3219 (N_3219,N_2697,N_2892);
nand U3220 (N_3220,N_2730,N_2646);
and U3221 (N_3221,N_2785,N_2738);
or U3222 (N_3222,N_2702,N_2570);
nor U3223 (N_3223,N_2777,N_2956);
nand U3224 (N_3224,N_2543,N_2924);
nor U3225 (N_3225,N_2518,N_2815);
xor U3226 (N_3226,N_2714,N_2528);
xor U3227 (N_3227,N_2554,N_2908);
nor U3228 (N_3228,N_2984,N_2966);
and U3229 (N_3229,N_2811,N_2729);
or U3230 (N_3230,N_2704,N_2715);
and U3231 (N_3231,N_2914,N_2741);
and U3232 (N_3232,N_2975,N_2635);
nand U3233 (N_3233,N_2987,N_2940);
or U3234 (N_3234,N_2610,N_2855);
nand U3235 (N_3235,N_2828,N_2519);
and U3236 (N_3236,N_2779,N_2999);
and U3237 (N_3237,N_2921,N_2926);
and U3238 (N_3238,N_2513,N_2505);
xnor U3239 (N_3239,N_2869,N_2692);
and U3240 (N_3240,N_2920,N_2683);
nor U3241 (N_3241,N_2835,N_2616);
and U3242 (N_3242,N_2693,N_2763);
nor U3243 (N_3243,N_2640,N_2660);
or U3244 (N_3244,N_2550,N_2709);
and U3245 (N_3245,N_2508,N_2532);
xnor U3246 (N_3246,N_2929,N_2952);
or U3247 (N_3247,N_2768,N_2658);
nand U3248 (N_3248,N_2910,N_2783);
nor U3249 (N_3249,N_2647,N_2548);
nand U3250 (N_3250,N_2879,N_2702);
nor U3251 (N_3251,N_2761,N_2872);
nor U3252 (N_3252,N_2557,N_2585);
nor U3253 (N_3253,N_2962,N_2621);
nor U3254 (N_3254,N_2755,N_2665);
xnor U3255 (N_3255,N_2841,N_2743);
xnor U3256 (N_3256,N_2501,N_2702);
xor U3257 (N_3257,N_2892,N_2542);
or U3258 (N_3258,N_2857,N_2947);
and U3259 (N_3259,N_2993,N_2941);
nand U3260 (N_3260,N_2597,N_2718);
nand U3261 (N_3261,N_2708,N_2571);
xnor U3262 (N_3262,N_2796,N_2769);
xor U3263 (N_3263,N_2713,N_2882);
nor U3264 (N_3264,N_2550,N_2906);
or U3265 (N_3265,N_2503,N_2557);
nand U3266 (N_3266,N_2568,N_2599);
and U3267 (N_3267,N_2848,N_2596);
nor U3268 (N_3268,N_2609,N_2989);
nor U3269 (N_3269,N_2843,N_2590);
nand U3270 (N_3270,N_2990,N_2876);
nand U3271 (N_3271,N_2562,N_2718);
and U3272 (N_3272,N_2810,N_2738);
xor U3273 (N_3273,N_2538,N_2508);
xor U3274 (N_3274,N_2840,N_2733);
nand U3275 (N_3275,N_2723,N_2950);
nand U3276 (N_3276,N_2731,N_2979);
nor U3277 (N_3277,N_2587,N_2936);
or U3278 (N_3278,N_2722,N_2535);
nor U3279 (N_3279,N_2841,N_2959);
or U3280 (N_3280,N_2545,N_2656);
nand U3281 (N_3281,N_2798,N_2672);
or U3282 (N_3282,N_2913,N_2839);
or U3283 (N_3283,N_2589,N_2628);
and U3284 (N_3284,N_2599,N_2635);
nand U3285 (N_3285,N_2954,N_2909);
nor U3286 (N_3286,N_2965,N_2983);
or U3287 (N_3287,N_2541,N_2911);
nand U3288 (N_3288,N_2920,N_2685);
or U3289 (N_3289,N_2742,N_2938);
nand U3290 (N_3290,N_2613,N_2943);
and U3291 (N_3291,N_2670,N_2979);
or U3292 (N_3292,N_2798,N_2515);
xnor U3293 (N_3293,N_2810,N_2831);
xor U3294 (N_3294,N_2986,N_2869);
nor U3295 (N_3295,N_2710,N_2599);
xnor U3296 (N_3296,N_2618,N_2569);
and U3297 (N_3297,N_2803,N_2591);
or U3298 (N_3298,N_2813,N_2966);
nor U3299 (N_3299,N_2965,N_2730);
nor U3300 (N_3300,N_2745,N_2723);
nand U3301 (N_3301,N_2513,N_2766);
nand U3302 (N_3302,N_2958,N_2874);
or U3303 (N_3303,N_2517,N_2600);
xnor U3304 (N_3304,N_2895,N_2611);
and U3305 (N_3305,N_2787,N_2573);
xor U3306 (N_3306,N_2733,N_2722);
nand U3307 (N_3307,N_2500,N_2920);
nand U3308 (N_3308,N_2806,N_2641);
nand U3309 (N_3309,N_2778,N_2868);
xnor U3310 (N_3310,N_2953,N_2864);
or U3311 (N_3311,N_2502,N_2977);
and U3312 (N_3312,N_2509,N_2909);
xor U3313 (N_3313,N_2884,N_2582);
nand U3314 (N_3314,N_2709,N_2907);
nor U3315 (N_3315,N_2521,N_2636);
nor U3316 (N_3316,N_2695,N_2772);
xnor U3317 (N_3317,N_2598,N_2601);
or U3318 (N_3318,N_2600,N_2908);
or U3319 (N_3319,N_2554,N_2830);
xnor U3320 (N_3320,N_2747,N_2814);
nor U3321 (N_3321,N_2663,N_2871);
xor U3322 (N_3322,N_2511,N_2702);
nor U3323 (N_3323,N_2752,N_2509);
and U3324 (N_3324,N_2896,N_2900);
and U3325 (N_3325,N_2986,N_2795);
and U3326 (N_3326,N_2721,N_2731);
or U3327 (N_3327,N_2913,N_2574);
nand U3328 (N_3328,N_2870,N_2559);
and U3329 (N_3329,N_2982,N_2634);
nor U3330 (N_3330,N_2697,N_2670);
nand U3331 (N_3331,N_2948,N_2867);
nor U3332 (N_3332,N_2630,N_2582);
xor U3333 (N_3333,N_2713,N_2929);
nor U3334 (N_3334,N_2999,N_2602);
nor U3335 (N_3335,N_2636,N_2627);
nand U3336 (N_3336,N_2505,N_2881);
or U3337 (N_3337,N_2910,N_2954);
nor U3338 (N_3338,N_2879,N_2929);
nand U3339 (N_3339,N_2784,N_2664);
xor U3340 (N_3340,N_2955,N_2832);
xor U3341 (N_3341,N_2652,N_2907);
xor U3342 (N_3342,N_2758,N_2533);
and U3343 (N_3343,N_2638,N_2948);
and U3344 (N_3344,N_2535,N_2522);
nand U3345 (N_3345,N_2906,N_2634);
nand U3346 (N_3346,N_2567,N_2733);
nand U3347 (N_3347,N_2688,N_2730);
or U3348 (N_3348,N_2753,N_2510);
nor U3349 (N_3349,N_2668,N_2958);
xor U3350 (N_3350,N_2673,N_2832);
nor U3351 (N_3351,N_2918,N_2822);
nand U3352 (N_3352,N_2682,N_2885);
and U3353 (N_3353,N_2538,N_2951);
or U3354 (N_3354,N_2634,N_2598);
and U3355 (N_3355,N_2520,N_2738);
and U3356 (N_3356,N_2644,N_2919);
nor U3357 (N_3357,N_2911,N_2531);
or U3358 (N_3358,N_2537,N_2523);
nor U3359 (N_3359,N_2598,N_2582);
nor U3360 (N_3360,N_2763,N_2612);
or U3361 (N_3361,N_2880,N_2835);
xor U3362 (N_3362,N_2912,N_2690);
and U3363 (N_3363,N_2722,N_2575);
nor U3364 (N_3364,N_2995,N_2872);
and U3365 (N_3365,N_2627,N_2817);
or U3366 (N_3366,N_2516,N_2783);
nand U3367 (N_3367,N_2676,N_2946);
and U3368 (N_3368,N_2582,N_2594);
nor U3369 (N_3369,N_2609,N_2667);
xor U3370 (N_3370,N_2650,N_2622);
xor U3371 (N_3371,N_2826,N_2506);
nor U3372 (N_3372,N_2864,N_2996);
xor U3373 (N_3373,N_2909,N_2840);
nor U3374 (N_3374,N_2857,N_2830);
and U3375 (N_3375,N_2968,N_2660);
and U3376 (N_3376,N_2534,N_2716);
xnor U3377 (N_3377,N_2924,N_2973);
nand U3378 (N_3378,N_2554,N_2911);
or U3379 (N_3379,N_2772,N_2968);
and U3380 (N_3380,N_2895,N_2561);
xor U3381 (N_3381,N_2646,N_2543);
nor U3382 (N_3382,N_2566,N_2512);
and U3383 (N_3383,N_2794,N_2733);
nor U3384 (N_3384,N_2986,N_2651);
or U3385 (N_3385,N_2594,N_2916);
nor U3386 (N_3386,N_2753,N_2617);
xor U3387 (N_3387,N_2972,N_2690);
nand U3388 (N_3388,N_2740,N_2760);
nor U3389 (N_3389,N_2624,N_2829);
nand U3390 (N_3390,N_2662,N_2879);
or U3391 (N_3391,N_2685,N_2759);
nor U3392 (N_3392,N_2785,N_2558);
and U3393 (N_3393,N_2891,N_2898);
nor U3394 (N_3394,N_2813,N_2844);
xnor U3395 (N_3395,N_2903,N_2801);
xor U3396 (N_3396,N_2726,N_2553);
xor U3397 (N_3397,N_2826,N_2503);
or U3398 (N_3398,N_2729,N_2979);
xnor U3399 (N_3399,N_2744,N_2613);
and U3400 (N_3400,N_2714,N_2720);
nor U3401 (N_3401,N_2510,N_2935);
and U3402 (N_3402,N_2616,N_2900);
nor U3403 (N_3403,N_2562,N_2888);
or U3404 (N_3404,N_2940,N_2823);
and U3405 (N_3405,N_2857,N_2705);
or U3406 (N_3406,N_2944,N_2703);
xnor U3407 (N_3407,N_2705,N_2958);
and U3408 (N_3408,N_2505,N_2955);
nand U3409 (N_3409,N_2616,N_2988);
nand U3410 (N_3410,N_2514,N_2871);
xor U3411 (N_3411,N_2744,N_2850);
xnor U3412 (N_3412,N_2942,N_2827);
or U3413 (N_3413,N_2561,N_2695);
nor U3414 (N_3414,N_2846,N_2747);
nand U3415 (N_3415,N_2984,N_2633);
xnor U3416 (N_3416,N_2837,N_2523);
nand U3417 (N_3417,N_2601,N_2854);
nand U3418 (N_3418,N_2929,N_2602);
or U3419 (N_3419,N_2952,N_2528);
and U3420 (N_3420,N_2981,N_2649);
nor U3421 (N_3421,N_2585,N_2708);
nor U3422 (N_3422,N_2598,N_2873);
xor U3423 (N_3423,N_2536,N_2718);
or U3424 (N_3424,N_2696,N_2671);
nor U3425 (N_3425,N_2688,N_2980);
xor U3426 (N_3426,N_2944,N_2550);
nand U3427 (N_3427,N_2636,N_2872);
and U3428 (N_3428,N_2664,N_2523);
nand U3429 (N_3429,N_2705,N_2866);
xnor U3430 (N_3430,N_2844,N_2599);
xnor U3431 (N_3431,N_2645,N_2905);
nand U3432 (N_3432,N_2713,N_2546);
xnor U3433 (N_3433,N_2868,N_2765);
nand U3434 (N_3434,N_2892,N_2822);
and U3435 (N_3435,N_2822,N_2582);
nor U3436 (N_3436,N_2524,N_2506);
nor U3437 (N_3437,N_2643,N_2566);
xnor U3438 (N_3438,N_2777,N_2605);
and U3439 (N_3439,N_2503,N_2889);
xor U3440 (N_3440,N_2617,N_2643);
or U3441 (N_3441,N_2762,N_2713);
xnor U3442 (N_3442,N_2630,N_2965);
xnor U3443 (N_3443,N_2627,N_2729);
or U3444 (N_3444,N_2993,N_2942);
nor U3445 (N_3445,N_2806,N_2804);
xor U3446 (N_3446,N_2935,N_2658);
nor U3447 (N_3447,N_2587,N_2579);
nand U3448 (N_3448,N_2838,N_2563);
xnor U3449 (N_3449,N_2781,N_2898);
or U3450 (N_3450,N_2786,N_2634);
xor U3451 (N_3451,N_2891,N_2950);
xnor U3452 (N_3452,N_2876,N_2815);
nand U3453 (N_3453,N_2525,N_2863);
xor U3454 (N_3454,N_2877,N_2878);
and U3455 (N_3455,N_2502,N_2848);
xnor U3456 (N_3456,N_2982,N_2603);
nand U3457 (N_3457,N_2890,N_2888);
xor U3458 (N_3458,N_2998,N_2559);
nor U3459 (N_3459,N_2896,N_2799);
nor U3460 (N_3460,N_2928,N_2636);
or U3461 (N_3461,N_2932,N_2911);
or U3462 (N_3462,N_2962,N_2708);
and U3463 (N_3463,N_2911,N_2948);
xnor U3464 (N_3464,N_2940,N_2886);
nand U3465 (N_3465,N_2693,N_2969);
xnor U3466 (N_3466,N_2810,N_2673);
xnor U3467 (N_3467,N_2821,N_2980);
nor U3468 (N_3468,N_2803,N_2637);
xor U3469 (N_3469,N_2677,N_2996);
or U3470 (N_3470,N_2501,N_2537);
xnor U3471 (N_3471,N_2878,N_2982);
nor U3472 (N_3472,N_2790,N_2728);
nor U3473 (N_3473,N_2984,N_2869);
nand U3474 (N_3474,N_2652,N_2610);
or U3475 (N_3475,N_2720,N_2586);
or U3476 (N_3476,N_2908,N_2794);
or U3477 (N_3477,N_2689,N_2627);
and U3478 (N_3478,N_2967,N_2549);
nor U3479 (N_3479,N_2871,N_2603);
nand U3480 (N_3480,N_2922,N_2646);
nand U3481 (N_3481,N_2530,N_2796);
nor U3482 (N_3482,N_2682,N_2697);
or U3483 (N_3483,N_2804,N_2964);
xor U3484 (N_3484,N_2787,N_2885);
or U3485 (N_3485,N_2681,N_2926);
xor U3486 (N_3486,N_2852,N_2506);
and U3487 (N_3487,N_2553,N_2791);
nand U3488 (N_3488,N_2586,N_2570);
nand U3489 (N_3489,N_2983,N_2957);
and U3490 (N_3490,N_2827,N_2867);
xnor U3491 (N_3491,N_2651,N_2863);
nor U3492 (N_3492,N_2887,N_2983);
xnor U3493 (N_3493,N_2763,N_2863);
and U3494 (N_3494,N_2971,N_2550);
nor U3495 (N_3495,N_2765,N_2874);
xnor U3496 (N_3496,N_2918,N_2699);
nor U3497 (N_3497,N_2574,N_2963);
and U3498 (N_3498,N_2896,N_2851);
or U3499 (N_3499,N_2925,N_2534);
or U3500 (N_3500,N_3496,N_3166);
and U3501 (N_3501,N_3067,N_3441);
and U3502 (N_3502,N_3319,N_3420);
nand U3503 (N_3503,N_3235,N_3105);
or U3504 (N_3504,N_3238,N_3134);
or U3505 (N_3505,N_3186,N_3359);
nor U3506 (N_3506,N_3495,N_3203);
or U3507 (N_3507,N_3361,N_3239);
or U3508 (N_3508,N_3453,N_3040);
nor U3509 (N_3509,N_3336,N_3430);
nand U3510 (N_3510,N_3218,N_3277);
nand U3511 (N_3511,N_3225,N_3059);
and U3512 (N_3512,N_3443,N_3199);
xor U3513 (N_3513,N_3070,N_3398);
nor U3514 (N_3514,N_3012,N_3342);
nor U3515 (N_3515,N_3088,N_3139);
xor U3516 (N_3516,N_3330,N_3331);
nand U3517 (N_3517,N_3071,N_3208);
and U3518 (N_3518,N_3432,N_3138);
nand U3519 (N_3519,N_3178,N_3376);
xnor U3520 (N_3520,N_3488,N_3050);
or U3521 (N_3521,N_3475,N_3299);
xnor U3522 (N_3522,N_3037,N_3324);
or U3523 (N_3523,N_3397,N_3018);
and U3524 (N_3524,N_3415,N_3472);
and U3525 (N_3525,N_3051,N_3272);
xor U3526 (N_3526,N_3349,N_3157);
nand U3527 (N_3527,N_3011,N_3114);
nand U3528 (N_3528,N_3303,N_3090);
and U3529 (N_3529,N_3484,N_3285);
nand U3530 (N_3530,N_3222,N_3276);
and U3531 (N_3531,N_3392,N_3162);
or U3532 (N_3532,N_3262,N_3395);
and U3533 (N_3533,N_3164,N_3409);
nor U3534 (N_3534,N_3217,N_3085);
xnor U3535 (N_3535,N_3391,N_3099);
and U3536 (N_3536,N_3448,N_3419);
nor U3537 (N_3537,N_3403,N_3060);
nand U3538 (N_3538,N_3388,N_3323);
or U3539 (N_3539,N_3023,N_3389);
and U3540 (N_3540,N_3030,N_3038);
and U3541 (N_3541,N_3130,N_3043);
or U3542 (N_3542,N_3245,N_3132);
and U3543 (N_3543,N_3160,N_3205);
or U3544 (N_3544,N_3461,N_3032);
xor U3545 (N_3545,N_3007,N_3044);
or U3546 (N_3546,N_3252,N_3219);
xor U3547 (N_3547,N_3268,N_3109);
or U3548 (N_3548,N_3026,N_3412);
nor U3549 (N_3549,N_3321,N_3387);
nor U3550 (N_3550,N_3146,N_3015);
nand U3551 (N_3551,N_3363,N_3092);
nor U3552 (N_3552,N_3131,N_3347);
nand U3553 (N_3553,N_3156,N_3192);
xnor U3554 (N_3554,N_3489,N_3234);
and U3555 (N_3555,N_3485,N_3444);
nor U3556 (N_3556,N_3343,N_3263);
nand U3557 (N_3557,N_3104,N_3127);
xor U3558 (N_3558,N_3357,N_3125);
or U3559 (N_3559,N_3456,N_3355);
xor U3560 (N_3560,N_3214,N_3490);
xnor U3561 (N_3561,N_3077,N_3098);
or U3562 (N_3562,N_3399,N_3035);
and U3563 (N_3563,N_3325,N_3020);
or U3564 (N_3564,N_3280,N_3148);
or U3565 (N_3565,N_3300,N_3297);
nor U3566 (N_3566,N_3188,N_3149);
nor U3567 (N_3567,N_3338,N_3438);
nand U3568 (N_3568,N_3337,N_3224);
nor U3569 (N_3569,N_3074,N_3163);
or U3570 (N_3570,N_3422,N_3406);
xnor U3571 (N_3571,N_3101,N_3463);
and U3572 (N_3572,N_3147,N_3108);
nor U3573 (N_3573,N_3264,N_3401);
and U3574 (N_3574,N_3426,N_3243);
and U3575 (N_3575,N_3492,N_3253);
nand U3576 (N_3576,N_3190,N_3402);
xor U3577 (N_3577,N_3143,N_3052);
or U3578 (N_3578,N_3258,N_3478);
nand U3579 (N_3579,N_3145,N_3182);
and U3580 (N_3580,N_3408,N_3123);
and U3581 (N_3581,N_3309,N_3251);
nor U3582 (N_3582,N_3332,N_3000);
xor U3583 (N_3583,N_3294,N_3194);
nor U3584 (N_3584,N_3446,N_3209);
nand U3585 (N_3585,N_3340,N_3317);
nor U3586 (N_3586,N_3047,N_3107);
nor U3587 (N_3587,N_3170,N_3291);
nor U3588 (N_3588,N_3173,N_3082);
nand U3589 (N_3589,N_3168,N_3322);
or U3590 (N_3590,N_3121,N_3236);
or U3591 (N_3591,N_3110,N_3117);
and U3592 (N_3592,N_3418,N_3255);
or U3593 (N_3593,N_3024,N_3482);
nor U3594 (N_3594,N_3233,N_3341);
and U3595 (N_3595,N_3008,N_3068);
nor U3596 (N_3596,N_3187,N_3137);
nor U3597 (N_3597,N_3036,N_3346);
xor U3598 (N_3598,N_3474,N_3014);
xnor U3599 (N_3599,N_3487,N_3435);
or U3600 (N_3600,N_3307,N_3028);
and U3601 (N_3601,N_3230,N_3304);
or U3602 (N_3602,N_3259,N_3126);
nor U3603 (N_3603,N_3053,N_3046);
or U3604 (N_3604,N_3016,N_3334);
xnor U3605 (N_3605,N_3013,N_3200);
and U3606 (N_3606,N_3031,N_3249);
nand U3607 (N_3607,N_3039,N_3494);
nor U3608 (N_3608,N_3497,N_3017);
and U3609 (N_3609,N_3498,N_3486);
xnor U3610 (N_3610,N_3351,N_3278);
and U3611 (N_3611,N_3370,N_3371);
or U3612 (N_3612,N_3298,N_3318);
and U3613 (N_3613,N_3350,N_3223);
and U3614 (N_3614,N_3310,N_3124);
and U3615 (N_3615,N_3177,N_3081);
or U3616 (N_3616,N_3119,N_3248);
nor U3617 (N_3617,N_3111,N_3083);
nor U3618 (N_3618,N_3103,N_3073);
and U3619 (N_3619,N_3042,N_3010);
xnor U3620 (N_3620,N_3381,N_3179);
or U3621 (N_3621,N_3279,N_3476);
nor U3622 (N_3622,N_3049,N_3167);
xor U3623 (N_3623,N_3410,N_3150);
or U3624 (N_3624,N_3369,N_3069);
nand U3625 (N_3625,N_3057,N_3404);
or U3626 (N_3626,N_3172,N_3006);
or U3627 (N_3627,N_3033,N_3451);
or U3628 (N_3628,N_3483,N_3189);
nand U3629 (N_3629,N_3380,N_3048);
and U3630 (N_3630,N_3440,N_3247);
nor U3631 (N_3631,N_3019,N_3241);
xor U3632 (N_3632,N_3362,N_3457);
nor U3633 (N_3633,N_3384,N_3458);
xor U3634 (N_3634,N_3154,N_3301);
or U3635 (N_3635,N_3064,N_3153);
xor U3636 (N_3636,N_3159,N_3091);
nor U3637 (N_3637,N_3282,N_3352);
or U3638 (N_3638,N_3424,N_3425);
or U3639 (N_3639,N_3118,N_3407);
xor U3640 (N_3640,N_3447,N_3335);
xnor U3641 (N_3641,N_3206,N_3436);
xnor U3642 (N_3642,N_3289,N_3454);
and U3643 (N_3643,N_3464,N_3041);
and U3644 (N_3644,N_3029,N_3393);
or U3645 (N_3645,N_3411,N_3326);
nand U3646 (N_3646,N_3140,N_3229);
and U3647 (N_3647,N_3356,N_3396);
or U3648 (N_3648,N_3433,N_3377);
xnor U3649 (N_3649,N_3292,N_3093);
nor U3650 (N_3650,N_3078,N_3311);
or U3651 (N_3651,N_3450,N_3261);
or U3652 (N_3652,N_3320,N_3204);
nand U3653 (N_3653,N_3169,N_3316);
xor U3654 (N_3654,N_3231,N_3021);
nor U3655 (N_3655,N_3378,N_3034);
nand U3656 (N_3656,N_3372,N_3174);
and U3657 (N_3657,N_3094,N_3246);
nor U3658 (N_3658,N_3287,N_3345);
xnor U3659 (N_3659,N_3305,N_3191);
and U3660 (N_3660,N_3465,N_3417);
and U3661 (N_3661,N_3133,N_3455);
nand U3662 (N_3662,N_3314,N_3469);
nor U3663 (N_3663,N_3423,N_3001);
and U3664 (N_3664,N_3221,N_3437);
nor U3665 (N_3665,N_3184,N_3212);
or U3666 (N_3666,N_3065,N_3273);
and U3667 (N_3667,N_3227,N_3267);
nor U3668 (N_3668,N_3055,N_3256);
or U3669 (N_3669,N_3009,N_3144);
and U3670 (N_3670,N_3244,N_3075);
nand U3671 (N_3671,N_3328,N_3327);
nor U3672 (N_3672,N_3152,N_3274);
xnor U3673 (N_3673,N_3480,N_3353);
xor U3674 (N_3674,N_3479,N_3281);
or U3675 (N_3675,N_3201,N_3066);
and U3676 (N_3676,N_3079,N_3383);
and U3677 (N_3677,N_3116,N_3265);
or U3678 (N_3678,N_3220,N_3493);
nor U3679 (N_3679,N_3100,N_3286);
nand U3680 (N_3680,N_3242,N_3106);
nor U3681 (N_3681,N_3364,N_3061);
or U3682 (N_3682,N_3471,N_3344);
nor U3683 (N_3683,N_3386,N_3385);
xor U3684 (N_3684,N_3115,N_3449);
nor U3685 (N_3685,N_3468,N_3076);
and U3686 (N_3686,N_3405,N_3462);
nor U3687 (N_3687,N_3266,N_3271);
or U3688 (N_3688,N_3491,N_3459);
or U3689 (N_3689,N_3431,N_3390);
or U3690 (N_3690,N_3312,N_3382);
xor U3691 (N_3691,N_3202,N_3445);
and U3692 (N_3692,N_3354,N_3270);
nor U3693 (N_3693,N_3004,N_3439);
nand U3694 (N_3694,N_3084,N_3113);
xor U3695 (N_3695,N_3141,N_3466);
or U3696 (N_3696,N_3250,N_3087);
nand U3697 (N_3697,N_3136,N_3413);
nor U3698 (N_3698,N_3228,N_3308);
nor U3699 (N_3699,N_3373,N_3195);
xor U3700 (N_3700,N_3213,N_3151);
nand U3701 (N_3701,N_3302,N_3002);
xnor U3702 (N_3702,N_3470,N_3368);
or U3703 (N_3703,N_3089,N_3460);
or U3704 (N_3704,N_3207,N_3348);
nand U3705 (N_3705,N_3176,N_3414);
nand U3706 (N_3706,N_3128,N_3269);
xnor U3707 (N_3707,N_3215,N_3211);
nand U3708 (N_3708,N_3056,N_3333);
or U3709 (N_3709,N_3315,N_3185);
and U3710 (N_3710,N_3275,N_3260);
nand U3711 (N_3711,N_3421,N_3197);
xnor U3712 (N_3712,N_3313,N_3063);
xnor U3713 (N_3713,N_3254,N_3232);
nor U3714 (N_3714,N_3142,N_3473);
xnor U3715 (N_3715,N_3155,N_3072);
nor U3716 (N_3716,N_3025,N_3120);
nor U3717 (N_3717,N_3096,N_3257);
nand U3718 (N_3718,N_3122,N_3358);
xor U3719 (N_3719,N_3434,N_3210);
and U3720 (N_3720,N_3027,N_3295);
and U3721 (N_3721,N_3296,N_3161);
nor U3722 (N_3722,N_3366,N_3102);
or U3723 (N_3723,N_3481,N_3339);
xnor U3724 (N_3724,N_3442,N_3400);
nor U3725 (N_3725,N_3135,N_3005);
xnor U3726 (N_3726,N_3290,N_3181);
nor U3727 (N_3727,N_3158,N_3198);
and U3728 (N_3728,N_3045,N_3427);
xnor U3729 (N_3729,N_3360,N_3054);
or U3730 (N_3730,N_3329,N_3086);
and U3731 (N_3731,N_3193,N_3080);
nor U3732 (N_3732,N_3058,N_3375);
or U3733 (N_3733,N_3129,N_3429);
or U3734 (N_3734,N_3097,N_3112);
and U3735 (N_3735,N_3288,N_3226);
nor U3736 (N_3736,N_3416,N_3171);
or U3737 (N_3737,N_3284,N_3477);
nor U3738 (N_3738,N_3095,N_3467);
nand U3739 (N_3739,N_3394,N_3379);
nor U3740 (N_3740,N_3293,N_3183);
nand U3741 (N_3741,N_3003,N_3499);
and U3742 (N_3742,N_3237,N_3365);
or U3743 (N_3743,N_3062,N_3240);
and U3744 (N_3744,N_3306,N_3196);
and U3745 (N_3745,N_3022,N_3452);
or U3746 (N_3746,N_3367,N_3180);
nor U3747 (N_3747,N_3165,N_3283);
or U3748 (N_3748,N_3216,N_3428);
nand U3749 (N_3749,N_3175,N_3374);
or U3750 (N_3750,N_3484,N_3128);
or U3751 (N_3751,N_3178,N_3277);
xor U3752 (N_3752,N_3412,N_3340);
nor U3753 (N_3753,N_3124,N_3088);
or U3754 (N_3754,N_3395,N_3243);
and U3755 (N_3755,N_3150,N_3313);
xnor U3756 (N_3756,N_3296,N_3038);
and U3757 (N_3757,N_3088,N_3236);
and U3758 (N_3758,N_3341,N_3368);
and U3759 (N_3759,N_3431,N_3025);
and U3760 (N_3760,N_3418,N_3112);
nor U3761 (N_3761,N_3200,N_3175);
or U3762 (N_3762,N_3153,N_3379);
nor U3763 (N_3763,N_3137,N_3159);
and U3764 (N_3764,N_3453,N_3405);
nand U3765 (N_3765,N_3117,N_3073);
nand U3766 (N_3766,N_3036,N_3027);
or U3767 (N_3767,N_3222,N_3007);
nor U3768 (N_3768,N_3001,N_3147);
or U3769 (N_3769,N_3368,N_3201);
nand U3770 (N_3770,N_3385,N_3446);
or U3771 (N_3771,N_3251,N_3267);
and U3772 (N_3772,N_3156,N_3054);
or U3773 (N_3773,N_3130,N_3237);
xnor U3774 (N_3774,N_3204,N_3181);
and U3775 (N_3775,N_3462,N_3386);
nor U3776 (N_3776,N_3146,N_3288);
and U3777 (N_3777,N_3033,N_3124);
nor U3778 (N_3778,N_3445,N_3121);
or U3779 (N_3779,N_3179,N_3393);
nand U3780 (N_3780,N_3125,N_3388);
nand U3781 (N_3781,N_3233,N_3496);
xor U3782 (N_3782,N_3476,N_3357);
nor U3783 (N_3783,N_3255,N_3411);
xnor U3784 (N_3784,N_3287,N_3330);
nand U3785 (N_3785,N_3109,N_3010);
nand U3786 (N_3786,N_3099,N_3260);
or U3787 (N_3787,N_3200,N_3071);
and U3788 (N_3788,N_3378,N_3447);
nor U3789 (N_3789,N_3175,N_3149);
xor U3790 (N_3790,N_3100,N_3258);
and U3791 (N_3791,N_3032,N_3101);
xnor U3792 (N_3792,N_3159,N_3327);
nor U3793 (N_3793,N_3374,N_3457);
xor U3794 (N_3794,N_3443,N_3389);
and U3795 (N_3795,N_3350,N_3401);
and U3796 (N_3796,N_3240,N_3451);
nand U3797 (N_3797,N_3188,N_3299);
or U3798 (N_3798,N_3185,N_3192);
nor U3799 (N_3799,N_3244,N_3299);
and U3800 (N_3800,N_3196,N_3166);
or U3801 (N_3801,N_3271,N_3169);
or U3802 (N_3802,N_3138,N_3458);
nand U3803 (N_3803,N_3465,N_3493);
or U3804 (N_3804,N_3377,N_3351);
and U3805 (N_3805,N_3281,N_3484);
xnor U3806 (N_3806,N_3432,N_3356);
xor U3807 (N_3807,N_3165,N_3247);
and U3808 (N_3808,N_3284,N_3481);
and U3809 (N_3809,N_3314,N_3112);
xor U3810 (N_3810,N_3242,N_3360);
or U3811 (N_3811,N_3051,N_3312);
or U3812 (N_3812,N_3021,N_3246);
or U3813 (N_3813,N_3111,N_3047);
or U3814 (N_3814,N_3474,N_3037);
nand U3815 (N_3815,N_3150,N_3272);
nor U3816 (N_3816,N_3354,N_3343);
nand U3817 (N_3817,N_3330,N_3055);
and U3818 (N_3818,N_3024,N_3166);
nand U3819 (N_3819,N_3092,N_3009);
xor U3820 (N_3820,N_3352,N_3055);
and U3821 (N_3821,N_3155,N_3023);
xor U3822 (N_3822,N_3262,N_3111);
nand U3823 (N_3823,N_3296,N_3077);
or U3824 (N_3824,N_3020,N_3449);
and U3825 (N_3825,N_3178,N_3037);
xor U3826 (N_3826,N_3096,N_3059);
nand U3827 (N_3827,N_3438,N_3159);
and U3828 (N_3828,N_3261,N_3047);
nor U3829 (N_3829,N_3201,N_3311);
or U3830 (N_3830,N_3035,N_3362);
xor U3831 (N_3831,N_3471,N_3374);
nand U3832 (N_3832,N_3115,N_3416);
xor U3833 (N_3833,N_3275,N_3160);
nor U3834 (N_3834,N_3234,N_3273);
or U3835 (N_3835,N_3477,N_3280);
and U3836 (N_3836,N_3343,N_3318);
and U3837 (N_3837,N_3105,N_3266);
xnor U3838 (N_3838,N_3309,N_3001);
nand U3839 (N_3839,N_3130,N_3387);
or U3840 (N_3840,N_3471,N_3180);
xnor U3841 (N_3841,N_3419,N_3313);
nand U3842 (N_3842,N_3449,N_3209);
nand U3843 (N_3843,N_3051,N_3391);
nand U3844 (N_3844,N_3201,N_3339);
or U3845 (N_3845,N_3432,N_3233);
nor U3846 (N_3846,N_3173,N_3477);
nand U3847 (N_3847,N_3261,N_3381);
and U3848 (N_3848,N_3234,N_3053);
nand U3849 (N_3849,N_3038,N_3418);
nand U3850 (N_3850,N_3488,N_3393);
nor U3851 (N_3851,N_3051,N_3480);
and U3852 (N_3852,N_3142,N_3117);
and U3853 (N_3853,N_3252,N_3474);
nor U3854 (N_3854,N_3194,N_3141);
and U3855 (N_3855,N_3126,N_3147);
nor U3856 (N_3856,N_3378,N_3107);
nand U3857 (N_3857,N_3373,N_3012);
nand U3858 (N_3858,N_3434,N_3328);
nor U3859 (N_3859,N_3091,N_3004);
or U3860 (N_3860,N_3275,N_3003);
or U3861 (N_3861,N_3141,N_3170);
nand U3862 (N_3862,N_3012,N_3204);
nor U3863 (N_3863,N_3133,N_3072);
nand U3864 (N_3864,N_3164,N_3469);
and U3865 (N_3865,N_3318,N_3065);
or U3866 (N_3866,N_3493,N_3432);
nand U3867 (N_3867,N_3492,N_3090);
and U3868 (N_3868,N_3220,N_3495);
and U3869 (N_3869,N_3213,N_3487);
and U3870 (N_3870,N_3307,N_3431);
nor U3871 (N_3871,N_3437,N_3002);
xor U3872 (N_3872,N_3011,N_3338);
and U3873 (N_3873,N_3270,N_3014);
nor U3874 (N_3874,N_3154,N_3481);
xnor U3875 (N_3875,N_3181,N_3309);
or U3876 (N_3876,N_3322,N_3328);
or U3877 (N_3877,N_3186,N_3017);
and U3878 (N_3878,N_3437,N_3083);
nor U3879 (N_3879,N_3101,N_3398);
or U3880 (N_3880,N_3408,N_3469);
nor U3881 (N_3881,N_3066,N_3050);
nor U3882 (N_3882,N_3377,N_3091);
or U3883 (N_3883,N_3449,N_3170);
and U3884 (N_3884,N_3491,N_3076);
xor U3885 (N_3885,N_3086,N_3431);
and U3886 (N_3886,N_3014,N_3342);
xnor U3887 (N_3887,N_3427,N_3171);
or U3888 (N_3888,N_3453,N_3299);
nand U3889 (N_3889,N_3180,N_3292);
xnor U3890 (N_3890,N_3358,N_3407);
and U3891 (N_3891,N_3212,N_3170);
or U3892 (N_3892,N_3393,N_3360);
and U3893 (N_3893,N_3421,N_3387);
and U3894 (N_3894,N_3017,N_3094);
nor U3895 (N_3895,N_3018,N_3031);
and U3896 (N_3896,N_3437,N_3335);
xnor U3897 (N_3897,N_3344,N_3466);
and U3898 (N_3898,N_3362,N_3220);
and U3899 (N_3899,N_3360,N_3213);
nor U3900 (N_3900,N_3360,N_3060);
nor U3901 (N_3901,N_3402,N_3282);
nor U3902 (N_3902,N_3416,N_3292);
and U3903 (N_3903,N_3128,N_3181);
or U3904 (N_3904,N_3083,N_3065);
or U3905 (N_3905,N_3400,N_3491);
nor U3906 (N_3906,N_3393,N_3356);
or U3907 (N_3907,N_3010,N_3065);
xnor U3908 (N_3908,N_3029,N_3250);
nand U3909 (N_3909,N_3285,N_3003);
xnor U3910 (N_3910,N_3263,N_3335);
and U3911 (N_3911,N_3053,N_3347);
nand U3912 (N_3912,N_3235,N_3288);
xor U3913 (N_3913,N_3000,N_3295);
nand U3914 (N_3914,N_3171,N_3222);
nand U3915 (N_3915,N_3169,N_3119);
nor U3916 (N_3916,N_3444,N_3357);
nand U3917 (N_3917,N_3440,N_3124);
nand U3918 (N_3918,N_3447,N_3199);
xor U3919 (N_3919,N_3315,N_3089);
nor U3920 (N_3920,N_3083,N_3092);
xor U3921 (N_3921,N_3174,N_3240);
or U3922 (N_3922,N_3358,N_3487);
xor U3923 (N_3923,N_3238,N_3199);
nand U3924 (N_3924,N_3481,N_3014);
nor U3925 (N_3925,N_3143,N_3063);
and U3926 (N_3926,N_3277,N_3259);
nor U3927 (N_3927,N_3429,N_3290);
and U3928 (N_3928,N_3414,N_3345);
nand U3929 (N_3929,N_3361,N_3067);
or U3930 (N_3930,N_3115,N_3291);
xor U3931 (N_3931,N_3055,N_3494);
nand U3932 (N_3932,N_3083,N_3471);
xnor U3933 (N_3933,N_3265,N_3307);
nor U3934 (N_3934,N_3141,N_3186);
or U3935 (N_3935,N_3313,N_3472);
nor U3936 (N_3936,N_3195,N_3065);
nor U3937 (N_3937,N_3326,N_3131);
and U3938 (N_3938,N_3374,N_3470);
nor U3939 (N_3939,N_3130,N_3054);
xnor U3940 (N_3940,N_3465,N_3171);
nand U3941 (N_3941,N_3151,N_3072);
and U3942 (N_3942,N_3272,N_3401);
nand U3943 (N_3943,N_3123,N_3351);
nor U3944 (N_3944,N_3042,N_3105);
xor U3945 (N_3945,N_3159,N_3463);
and U3946 (N_3946,N_3010,N_3001);
xnor U3947 (N_3947,N_3267,N_3041);
or U3948 (N_3948,N_3257,N_3254);
nor U3949 (N_3949,N_3314,N_3313);
xor U3950 (N_3950,N_3062,N_3292);
and U3951 (N_3951,N_3463,N_3164);
nor U3952 (N_3952,N_3100,N_3289);
nand U3953 (N_3953,N_3142,N_3130);
and U3954 (N_3954,N_3244,N_3228);
nand U3955 (N_3955,N_3492,N_3296);
nand U3956 (N_3956,N_3442,N_3237);
nand U3957 (N_3957,N_3111,N_3484);
and U3958 (N_3958,N_3162,N_3035);
nand U3959 (N_3959,N_3313,N_3337);
nor U3960 (N_3960,N_3445,N_3383);
nor U3961 (N_3961,N_3112,N_3288);
or U3962 (N_3962,N_3395,N_3175);
nor U3963 (N_3963,N_3306,N_3398);
nor U3964 (N_3964,N_3350,N_3046);
nand U3965 (N_3965,N_3181,N_3263);
xor U3966 (N_3966,N_3421,N_3159);
or U3967 (N_3967,N_3199,N_3283);
xor U3968 (N_3968,N_3237,N_3126);
nand U3969 (N_3969,N_3041,N_3350);
or U3970 (N_3970,N_3073,N_3316);
or U3971 (N_3971,N_3311,N_3412);
and U3972 (N_3972,N_3353,N_3389);
xor U3973 (N_3973,N_3054,N_3382);
nand U3974 (N_3974,N_3142,N_3357);
and U3975 (N_3975,N_3075,N_3213);
and U3976 (N_3976,N_3011,N_3239);
and U3977 (N_3977,N_3325,N_3163);
nor U3978 (N_3978,N_3451,N_3198);
and U3979 (N_3979,N_3413,N_3206);
nand U3980 (N_3980,N_3209,N_3248);
xnor U3981 (N_3981,N_3215,N_3377);
xor U3982 (N_3982,N_3274,N_3388);
and U3983 (N_3983,N_3067,N_3404);
nand U3984 (N_3984,N_3361,N_3376);
nand U3985 (N_3985,N_3165,N_3443);
nand U3986 (N_3986,N_3383,N_3015);
nand U3987 (N_3987,N_3255,N_3278);
and U3988 (N_3988,N_3278,N_3002);
and U3989 (N_3989,N_3112,N_3159);
or U3990 (N_3990,N_3423,N_3440);
xnor U3991 (N_3991,N_3343,N_3046);
nor U3992 (N_3992,N_3190,N_3137);
and U3993 (N_3993,N_3497,N_3094);
xor U3994 (N_3994,N_3085,N_3355);
xor U3995 (N_3995,N_3356,N_3235);
and U3996 (N_3996,N_3027,N_3421);
and U3997 (N_3997,N_3082,N_3054);
nor U3998 (N_3998,N_3473,N_3391);
xnor U3999 (N_3999,N_3045,N_3407);
or U4000 (N_4000,N_3769,N_3986);
xor U4001 (N_4001,N_3990,N_3975);
and U4002 (N_4002,N_3669,N_3994);
nand U4003 (N_4003,N_3979,N_3968);
xnor U4004 (N_4004,N_3629,N_3795);
nor U4005 (N_4005,N_3964,N_3650);
and U4006 (N_4006,N_3544,N_3542);
nor U4007 (N_4007,N_3703,N_3872);
or U4008 (N_4008,N_3779,N_3783);
nand U4009 (N_4009,N_3527,N_3899);
xor U4010 (N_4010,N_3992,N_3880);
and U4011 (N_4011,N_3746,N_3826);
nand U4012 (N_4012,N_3583,N_3891);
and U4013 (N_4013,N_3988,N_3612);
nand U4014 (N_4014,N_3755,N_3858);
and U4015 (N_4015,N_3649,N_3913);
nor U4016 (N_4016,N_3907,N_3934);
nand U4017 (N_4017,N_3809,N_3545);
nand U4018 (N_4018,N_3712,N_3705);
or U4019 (N_4019,N_3831,N_3620);
nand U4020 (N_4020,N_3663,N_3726);
nor U4021 (N_4021,N_3509,N_3697);
nor U4022 (N_4022,N_3626,N_3757);
or U4023 (N_4023,N_3977,N_3548);
nor U4024 (N_4024,N_3958,N_3512);
nand U4025 (N_4025,N_3846,N_3694);
and U4026 (N_4026,N_3800,N_3867);
xor U4027 (N_4027,N_3517,N_3941);
xor U4028 (N_4028,N_3801,N_3980);
nand U4029 (N_4029,N_3943,N_3895);
xor U4030 (N_4030,N_3804,N_3947);
xnor U4031 (N_4031,N_3820,N_3824);
and U4032 (N_4032,N_3675,N_3734);
nand U4033 (N_4033,N_3571,N_3728);
nand U4034 (N_4034,N_3580,N_3767);
or U4035 (N_4035,N_3744,N_3984);
or U4036 (N_4036,N_3614,N_3752);
xnor U4037 (N_4037,N_3729,N_3554);
nand U4038 (N_4038,N_3569,N_3641);
nand U4039 (N_4039,N_3791,N_3922);
nand U4040 (N_4040,N_3806,N_3938);
xor U4041 (N_4041,N_3701,N_3516);
or U4042 (N_4042,N_3508,N_3910);
or U4043 (N_4043,N_3631,N_3605);
nor U4044 (N_4044,N_3736,N_3957);
nand U4045 (N_4045,N_3985,N_3682);
nand U4046 (N_4046,N_3638,N_3608);
nor U4047 (N_4047,N_3514,N_3999);
nand U4048 (N_4048,N_3749,N_3533);
nand U4049 (N_4049,N_3901,N_3772);
nand U4050 (N_4050,N_3504,N_3616);
or U4051 (N_4051,N_3507,N_3933);
nand U4052 (N_4052,N_3646,N_3923);
nor U4053 (N_4053,N_3596,N_3573);
and U4054 (N_4054,N_3978,N_3671);
or U4055 (N_4055,N_3720,N_3925);
and U4056 (N_4056,N_3929,N_3528);
nand U4057 (N_4057,N_3763,N_3642);
or U4058 (N_4058,N_3883,N_3981);
nand U4059 (N_4059,N_3607,N_3799);
nor U4060 (N_4060,N_3756,N_3843);
nor U4061 (N_4061,N_3724,N_3802);
nor U4062 (N_4062,N_3515,N_3661);
nand U4063 (N_4063,N_3568,N_3719);
xor U4064 (N_4064,N_3559,N_3630);
xnor U4065 (N_4065,N_3645,N_3759);
nor U4066 (N_4066,N_3892,N_3911);
xnor U4067 (N_4067,N_3590,N_3625);
xnor U4068 (N_4068,N_3885,N_3893);
nor U4069 (N_4069,N_3534,N_3577);
and U4070 (N_4070,N_3730,N_3776);
xor U4071 (N_4071,N_3648,N_3857);
nor U4072 (N_4072,N_3853,N_3627);
nand U4073 (N_4073,N_3737,N_3502);
nand U4074 (N_4074,N_3793,N_3819);
nor U4075 (N_4075,N_3942,N_3537);
xnor U4076 (N_4076,N_3969,N_3635);
nor U4077 (N_4077,N_3844,N_3636);
nor U4078 (N_4078,N_3796,N_3982);
and U4079 (N_4079,N_3556,N_3774);
nand U4080 (N_4080,N_3618,N_3816);
nor U4081 (N_4081,N_3909,N_3830);
xor U4082 (N_4082,N_3570,N_3996);
nor U4083 (N_4083,N_3722,N_3547);
and U4084 (N_4084,N_3597,N_3731);
and U4085 (N_4085,N_3829,N_3550);
or U4086 (N_4086,N_3790,N_3866);
and U4087 (N_4087,N_3860,N_3887);
and U4088 (N_4088,N_3777,N_3739);
and U4089 (N_4089,N_3924,N_3558);
or U4090 (N_4090,N_3588,N_3567);
nand U4091 (N_4091,N_3871,N_3935);
xor U4092 (N_4092,N_3666,N_3639);
nand U4093 (N_4093,N_3691,N_3662);
xor U4094 (N_4094,N_3735,N_3751);
nor U4095 (N_4095,N_3535,N_3561);
or U4096 (N_4096,N_3989,N_3825);
or U4097 (N_4097,N_3747,N_3681);
and U4098 (N_4098,N_3814,N_3797);
or U4099 (N_4099,N_3927,N_3594);
xnor U4100 (N_4100,N_3584,N_3503);
xor U4101 (N_4101,N_3847,N_3762);
xor U4102 (N_4102,N_3531,N_3785);
and U4103 (N_4103,N_3678,N_3741);
xor U4104 (N_4104,N_3604,N_3684);
nand U4105 (N_4105,N_3837,N_3578);
nor U4106 (N_4106,N_3715,N_3953);
nor U4107 (N_4107,N_3812,N_3794);
xnor U4108 (N_4108,N_3881,N_3764);
and U4109 (N_4109,N_3889,N_3928);
xnor U4110 (N_4110,N_3900,N_3738);
nor U4111 (N_4111,N_3810,N_3813);
xor U4112 (N_4112,N_3840,N_3939);
and U4113 (N_4113,N_3827,N_3742);
or U4114 (N_4114,N_3564,N_3699);
xor U4115 (N_4115,N_3771,N_3654);
nand U4116 (N_4116,N_3864,N_3619);
nand U4117 (N_4117,N_3949,N_3637);
nor U4118 (N_4118,N_3879,N_3613);
and U4119 (N_4119,N_3601,N_3760);
xor U4120 (N_4120,N_3510,N_3842);
nand U4121 (N_4121,N_3593,N_3700);
and U4122 (N_4122,N_3963,N_3833);
nand U4123 (N_4123,N_3967,N_3713);
or U4124 (N_4124,N_3782,N_3983);
nand U4125 (N_4125,N_3972,N_3665);
xor U4126 (N_4126,N_3587,N_3773);
xor U4127 (N_4127,N_3716,N_3575);
nand U4128 (N_4128,N_3960,N_3894);
xnor U4129 (N_4129,N_3965,N_3740);
xnor U4130 (N_4130,N_3634,N_3946);
nor U4131 (N_4131,N_3788,N_3818);
and U4132 (N_4132,N_3815,N_3803);
nand U4133 (N_4133,N_3997,N_3640);
or U4134 (N_4134,N_3657,N_3538);
nand U4135 (N_4135,N_3898,N_3930);
xor U4136 (N_4136,N_3768,N_3750);
nor U4137 (N_4137,N_3539,N_3674);
nand U4138 (N_4138,N_3706,N_3655);
nor U4139 (N_4139,N_3991,N_3805);
or U4140 (N_4140,N_3617,N_3621);
xnor U4141 (N_4141,N_3652,N_3600);
xor U4142 (N_4142,N_3670,N_3529);
nand U4143 (N_4143,N_3656,N_3526);
nand U4144 (N_4144,N_3623,N_3970);
nand U4145 (N_4145,N_3677,N_3693);
nand U4146 (N_4146,N_3851,N_3521);
xnor U4147 (N_4147,N_3672,N_3505);
and U4148 (N_4148,N_3552,N_3973);
and U4149 (N_4149,N_3676,N_3565);
xnor U4150 (N_4150,N_3823,N_3828);
nand U4151 (N_4151,N_3723,N_3950);
nand U4152 (N_4152,N_3944,N_3778);
nor U4153 (N_4153,N_3589,N_3849);
and U4154 (N_4154,N_3501,N_3838);
nand U4155 (N_4155,N_3572,N_3566);
nand U4156 (N_4156,N_3955,N_3884);
nor U4157 (N_4157,N_3956,N_3850);
nor U4158 (N_4158,N_3836,N_3822);
nor U4159 (N_4159,N_3733,N_3852);
nand U4160 (N_4160,N_3518,N_3915);
or U4161 (N_4161,N_3974,N_3886);
xor U4162 (N_4162,N_3993,N_3921);
nand U4163 (N_4163,N_3954,N_3692);
and U4164 (N_4164,N_3543,N_3717);
nand U4165 (N_4165,N_3951,N_3859);
xnor U4166 (N_4166,N_3848,N_3835);
nor U4167 (N_4167,N_3781,N_3586);
and U4168 (N_4168,N_3916,N_3668);
or U4169 (N_4169,N_3856,N_3520);
xnor U4170 (N_4170,N_3709,N_3702);
nor U4171 (N_4171,N_3667,N_3714);
nand U4172 (N_4172,N_3727,N_3904);
and U4173 (N_4173,N_3917,N_3875);
nand U4174 (N_4174,N_3732,N_3890);
and U4175 (N_4175,N_3937,N_3761);
xnor U4176 (N_4176,N_3873,N_3609);
and U4177 (N_4177,N_3841,N_3780);
xor U4178 (N_4178,N_3753,N_3585);
or U4179 (N_4179,N_3952,N_3659);
xnor U4180 (N_4180,N_3811,N_3821);
nor U4181 (N_4181,N_3513,N_3863);
and U4182 (N_4182,N_3932,N_3708);
nor U4183 (N_4183,N_3754,N_3987);
nor U4184 (N_4184,N_3870,N_3511);
xnor U4185 (N_4185,N_3786,N_3882);
xor U4186 (N_4186,N_3817,N_3926);
nor U4187 (N_4187,N_3563,N_3976);
and U4188 (N_4188,N_3660,N_3673);
and U4189 (N_4189,N_3845,N_3888);
and U4190 (N_4190,N_3748,N_3683);
xnor U4191 (N_4191,N_3710,N_3628);
or U4192 (N_4192,N_3834,N_3553);
nor U4193 (N_4193,N_3591,N_3903);
and U4194 (N_4194,N_3798,N_3592);
nor U4195 (N_4195,N_3546,N_3966);
nor U4196 (N_4196,N_3653,N_3962);
xor U4197 (N_4197,N_3536,N_3862);
xor U4198 (N_4198,N_3868,N_3765);
nand U4199 (N_4199,N_3602,N_3555);
or U4200 (N_4200,N_3721,N_3869);
nor U4201 (N_4201,N_3599,N_3971);
nand U4202 (N_4202,N_3787,N_3680);
nor U4203 (N_4203,N_3995,N_3745);
and U4204 (N_4204,N_3549,N_3579);
nor U4205 (N_4205,N_3743,N_3876);
and U4206 (N_4206,N_3598,N_3689);
xor U4207 (N_4207,N_3908,N_3919);
xnor U4208 (N_4208,N_3861,N_3865);
and U4209 (N_4209,N_3603,N_3948);
and U4210 (N_4210,N_3914,N_3688);
nor U4211 (N_4211,N_3664,N_3897);
and U4212 (N_4212,N_3615,N_3506);
nor U4213 (N_4213,N_3920,N_3690);
xnor U4214 (N_4214,N_3912,N_3540);
and U4215 (N_4215,N_3839,N_3582);
nor U4216 (N_4216,N_3695,N_3905);
or U4217 (N_4217,N_3931,N_3647);
or U4218 (N_4218,N_3562,N_3576);
xor U4219 (N_4219,N_3595,N_3644);
nand U4220 (N_4220,N_3522,N_3808);
nand U4221 (N_4221,N_3686,N_3633);
nand U4222 (N_4222,N_3718,N_3581);
nand U4223 (N_4223,N_3854,N_3789);
and U4224 (N_4224,N_3698,N_3832);
and U4225 (N_4225,N_3918,N_3961);
or U4226 (N_4226,N_3519,N_3766);
nand U4227 (N_4227,N_3998,N_3792);
and U4228 (N_4228,N_3896,N_3685);
or U4229 (N_4229,N_3524,N_3679);
xnor U4230 (N_4230,N_3725,N_3622);
and U4231 (N_4231,N_3687,N_3807);
xnor U4232 (N_4232,N_3770,N_3560);
and U4233 (N_4233,N_3624,N_3940);
nor U4234 (N_4234,N_3611,N_3855);
and U4235 (N_4235,N_3704,N_3784);
xnor U4236 (N_4236,N_3610,N_3500);
nor U4237 (N_4237,N_3658,N_3874);
xor U4238 (N_4238,N_3632,N_3959);
nor U4239 (N_4239,N_3525,N_3711);
or U4240 (N_4240,N_3758,N_3877);
xor U4241 (N_4241,N_3775,N_3878);
and U4242 (N_4242,N_3945,N_3557);
nor U4243 (N_4243,N_3643,N_3902);
nand U4244 (N_4244,N_3574,N_3651);
xnor U4245 (N_4245,N_3532,N_3530);
nand U4246 (N_4246,N_3906,N_3936);
or U4247 (N_4247,N_3523,N_3541);
or U4248 (N_4248,N_3551,N_3707);
xnor U4249 (N_4249,N_3606,N_3696);
xnor U4250 (N_4250,N_3859,N_3687);
or U4251 (N_4251,N_3888,N_3734);
or U4252 (N_4252,N_3934,N_3856);
xnor U4253 (N_4253,N_3835,N_3859);
nor U4254 (N_4254,N_3962,N_3968);
nand U4255 (N_4255,N_3898,N_3675);
nand U4256 (N_4256,N_3994,N_3915);
nor U4257 (N_4257,N_3528,N_3543);
or U4258 (N_4258,N_3510,N_3681);
or U4259 (N_4259,N_3956,N_3940);
and U4260 (N_4260,N_3860,N_3556);
xor U4261 (N_4261,N_3905,N_3827);
and U4262 (N_4262,N_3866,N_3710);
nand U4263 (N_4263,N_3598,N_3618);
or U4264 (N_4264,N_3572,N_3506);
nand U4265 (N_4265,N_3907,N_3992);
nand U4266 (N_4266,N_3869,N_3579);
nor U4267 (N_4267,N_3936,N_3988);
nand U4268 (N_4268,N_3816,N_3501);
xnor U4269 (N_4269,N_3928,N_3582);
nand U4270 (N_4270,N_3893,N_3811);
xnor U4271 (N_4271,N_3827,N_3649);
nand U4272 (N_4272,N_3734,N_3916);
nand U4273 (N_4273,N_3509,N_3868);
nand U4274 (N_4274,N_3566,N_3500);
nor U4275 (N_4275,N_3726,N_3932);
and U4276 (N_4276,N_3752,N_3667);
nor U4277 (N_4277,N_3999,N_3585);
xnor U4278 (N_4278,N_3627,N_3509);
xnor U4279 (N_4279,N_3907,N_3679);
xnor U4280 (N_4280,N_3507,N_3846);
and U4281 (N_4281,N_3981,N_3833);
or U4282 (N_4282,N_3589,N_3657);
nor U4283 (N_4283,N_3833,N_3970);
nand U4284 (N_4284,N_3722,N_3555);
nand U4285 (N_4285,N_3506,N_3797);
nand U4286 (N_4286,N_3899,N_3810);
nor U4287 (N_4287,N_3929,N_3767);
nor U4288 (N_4288,N_3909,N_3594);
xnor U4289 (N_4289,N_3727,N_3819);
and U4290 (N_4290,N_3510,N_3641);
nand U4291 (N_4291,N_3997,N_3728);
nor U4292 (N_4292,N_3508,N_3823);
xnor U4293 (N_4293,N_3902,N_3958);
xnor U4294 (N_4294,N_3861,N_3809);
xor U4295 (N_4295,N_3594,N_3617);
xnor U4296 (N_4296,N_3764,N_3511);
nor U4297 (N_4297,N_3506,N_3736);
nand U4298 (N_4298,N_3913,N_3675);
or U4299 (N_4299,N_3551,N_3695);
and U4300 (N_4300,N_3669,N_3660);
or U4301 (N_4301,N_3558,N_3920);
xor U4302 (N_4302,N_3827,N_3946);
nand U4303 (N_4303,N_3895,N_3605);
or U4304 (N_4304,N_3936,N_3935);
nand U4305 (N_4305,N_3514,N_3881);
xor U4306 (N_4306,N_3915,N_3888);
xnor U4307 (N_4307,N_3859,N_3786);
and U4308 (N_4308,N_3944,N_3500);
nand U4309 (N_4309,N_3814,N_3568);
or U4310 (N_4310,N_3982,N_3504);
xor U4311 (N_4311,N_3594,N_3614);
and U4312 (N_4312,N_3953,N_3517);
and U4313 (N_4313,N_3832,N_3613);
and U4314 (N_4314,N_3736,N_3566);
or U4315 (N_4315,N_3706,N_3976);
nor U4316 (N_4316,N_3748,N_3501);
or U4317 (N_4317,N_3919,N_3566);
or U4318 (N_4318,N_3913,N_3882);
nor U4319 (N_4319,N_3798,N_3927);
xnor U4320 (N_4320,N_3744,N_3592);
xor U4321 (N_4321,N_3801,N_3663);
and U4322 (N_4322,N_3679,N_3652);
nand U4323 (N_4323,N_3940,N_3867);
nand U4324 (N_4324,N_3537,N_3693);
xor U4325 (N_4325,N_3903,N_3679);
xor U4326 (N_4326,N_3929,N_3660);
or U4327 (N_4327,N_3585,N_3938);
nor U4328 (N_4328,N_3954,N_3907);
xor U4329 (N_4329,N_3506,N_3891);
nor U4330 (N_4330,N_3949,N_3775);
nand U4331 (N_4331,N_3890,N_3903);
or U4332 (N_4332,N_3516,N_3645);
nand U4333 (N_4333,N_3841,N_3857);
xnor U4334 (N_4334,N_3599,N_3787);
and U4335 (N_4335,N_3934,N_3835);
and U4336 (N_4336,N_3826,N_3944);
and U4337 (N_4337,N_3927,N_3611);
and U4338 (N_4338,N_3792,N_3674);
nand U4339 (N_4339,N_3615,N_3669);
nor U4340 (N_4340,N_3928,N_3709);
xnor U4341 (N_4341,N_3583,N_3631);
xor U4342 (N_4342,N_3708,N_3662);
xnor U4343 (N_4343,N_3802,N_3607);
or U4344 (N_4344,N_3789,N_3617);
nand U4345 (N_4345,N_3684,N_3810);
xor U4346 (N_4346,N_3712,N_3673);
or U4347 (N_4347,N_3570,N_3960);
nor U4348 (N_4348,N_3592,N_3750);
nor U4349 (N_4349,N_3596,N_3695);
nor U4350 (N_4350,N_3549,N_3828);
xnor U4351 (N_4351,N_3946,N_3612);
xnor U4352 (N_4352,N_3676,N_3761);
nor U4353 (N_4353,N_3948,N_3857);
or U4354 (N_4354,N_3962,N_3923);
and U4355 (N_4355,N_3767,N_3779);
or U4356 (N_4356,N_3616,N_3925);
nor U4357 (N_4357,N_3570,N_3758);
and U4358 (N_4358,N_3942,N_3929);
nor U4359 (N_4359,N_3710,N_3678);
or U4360 (N_4360,N_3809,N_3793);
and U4361 (N_4361,N_3819,N_3774);
nand U4362 (N_4362,N_3781,N_3715);
xor U4363 (N_4363,N_3745,N_3818);
nand U4364 (N_4364,N_3766,N_3658);
and U4365 (N_4365,N_3501,N_3882);
and U4366 (N_4366,N_3853,N_3656);
nand U4367 (N_4367,N_3955,N_3586);
xor U4368 (N_4368,N_3853,N_3950);
nand U4369 (N_4369,N_3699,N_3688);
or U4370 (N_4370,N_3965,N_3847);
xnor U4371 (N_4371,N_3669,N_3550);
or U4372 (N_4372,N_3544,N_3742);
and U4373 (N_4373,N_3677,N_3539);
xnor U4374 (N_4374,N_3605,N_3544);
or U4375 (N_4375,N_3941,N_3907);
nand U4376 (N_4376,N_3554,N_3560);
nand U4377 (N_4377,N_3647,N_3638);
and U4378 (N_4378,N_3559,N_3648);
xor U4379 (N_4379,N_3762,N_3837);
xor U4380 (N_4380,N_3764,N_3728);
or U4381 (N_4381,N_3570,N_3994);
and U4382 (N_4382,N_3951,N_3949);
nand U4383 (N_4383,N_3653,N_3846);
nand U4384 (N_4384,N_3969,N_3786);
xnor U4385 (N_4385,N_3505,N_3785);
nor U4386 (N_4386,N_3694,N_3993);
or U4387 (N_4387,N_3893,N_3798);
nor U4388 (N_4388,N_3994,N_3677);
nor U4389 (N_4389,N_3559,N_3831);
and U4390 (N_4390,N_3777,N_3715);
nor U4391 (N_4391,N_3939,N_3774);
and U4392 (N_4392,N_3938,N_3846);
xnor U4393 (N_4393,N_3747,N_3566);
and U4394 (N_4394,N_3862,N_3899);
or U4395 (N_4395,N_3653,N_3978);
or U4396 (N_4396,N_3503,N_3817);
xor U4397 (N_4397,N_3624,N_3657);
and U4398 (N_4398,N_3977,N_3651);
and U4399 (N_4399,N_3553,N_3753);
and U4400 (N_4400,N_3808,N_3553);
nor U4401 (N_4401,N_3982,N_3983);
nor U4402 (N_4402,N_3824,N_3660);
or U4403 (N_4403,N_3695,N_3565);
xor U4404 (N_4404,N_3972,N_3517);
and U4405 (N_4405,N_3525,N_3610);
or U4406 (N_4406,N_3579,N_3643);
nor U4407 (N_4407,N_3979,N_3649);
or U4408 (N_4408,N_3697,N_3733);
and U4409 (N_4409,N_3696,N_3839);
xor U4410 (N_4410,N_3575,N_3570);
and U4411 (N_4411,N_3782,N_3806);
nand U4412 (N_4412,N_3959,N_3568);
and U4413 (N_4413,N_3894,N_3848);
nand U4414 (N_4414,N_3741,N_3753);
xnor U4415 (N_4415,N_3604,N_3842);
xnor U4416 (N_4416,N_3768,N_3785);
nor U4417 (N_4417,N_3815,N_3730);
nor U4418 (N_4418,N_3588,N_3532);
nand U4419 (N_4419,N_3852,N_3570);
nor U4420 (N_4420,N_3757,N_3719);
xnor U4421 (N_4421,N_3950,N_3903);
and U4422 (N_4422,N_3826,N_3628);
nand U4423 (N_4423,N_3534,N_3551);
or U4424 (N_4424,N_3817,N_3994);
nor U4425 (N_4425,N_3898,N_3850);
nor U4426 (N_4426,N_3765,N_3674);
and U4427 (N_4427,N_3987,N_3937);
nand U4428 (N_4428,N_3774,N_3776);
nor U4429 (N_4429,N_3969,N_3936);
and U4430 (N_4430,N_3792,N_3543);
or U4431 (N_4431,N_3814,N_3919);
xor U4432 (N_4432,N_3793,N_3912);
xnor U4433 (N_4433,N_3684,N_3527);
xor U4434 (N_4434,N_3555,N_3615);
xnor U4435 (N_4435,N_3555,N_3845);
nor U4436 (N_4436,N_3571,N_3557);
or U4437 (N_4437,N_3830,N_3614);
or U4438 (N_4438,N_3971,N_3671);
xnor U4439 (N_4439,N_3693,N_3641);
and U4440 (N_4440,N_3524,N_3741);
nor U4441 (N_4441,N_3616,N_3627);
or U4442 (N_4442,N_3774,N_3550);
nor U4443 (N_4443,N_3900,N_3642);
and U4444 (N_4444,N_3893,N_3698);
or U4445 (N_4445,N_3936,N_3842);
xor U4446 (N_4446,N_3681,N_3752);
or U4447 (N_4447,N_3647,N_3605);
nor U4448 (N_4448,N_3893,N_3503);
nor U4449 (N_4449,N_3947,N_3589);
nor U4450 (N_4450,N_3622,N_3826);
xnor U4451 (N_4451,N_3500,N_3540);
xor U4452 (N_4452,N_3596,N_3863);
xnor U4453 (N_4453,N_3961,N_3726);
nand U4454 (N_4454,N_3526,N_3683);
xnor U4455 (N_4455,N_3964,N_3634);
nand U4456 (N_4456,N_3714,N_3542);
nor U4457 (N_4457,N_3590,N_3684);
or U4458 (N_4458,N_3595,N_3521);
or U4459 (N_4459,N_3814,N_3854);
or U4460 (N_4460,N_3631,N_3570);
and U4461 (N_4461,N_3843,N_3742);
nand U4462 (N_4462,N_3674,N_3895);
nor U4463 (N_4463,N_3998,N_3666);
or U4464 (N_4464,N_3575,N_3773);
or U4465 (N_4465,N_3512,N_3756);
nor U4466 (N_4466,N_3707,N_3524);
nor U4467 (N_4467,N_3682,N_3879);
nor U4468 (N_4468,N_3802,N_3818);
nor U4469 (N_4469,N_3982,N_3726);
nor U4470 (N_4470,N_3655,N_3986);
and U4471 (N_4471,N_3914,N_3862);
and U4472 (N_4472,N_3532,N_3628);
nand U4473 (N_4473,N_3765,N_3753);
nor U4474 (N_4474,N_3789,N_3859);
and U4475 (N_4475,N_3617,N_3832);
xor U4476 (N_4476,N_3793,N_3546);
and U4477 (N_4477,N_3943,N_3838);
xnor U4478 (N_4478,N_3922,N_3519);
or U4479 (N_4479,N_3702,N_3567);
and U4480 (N_4480,N_3541,N_3712);
nand U4481 (N_4481,N_3964,N_3947);
and U4482 (N_4482,N_3685,N_3662);
nor U4483 (N_4483,N_3555,N_3737);
or U4484 (N_4484,N_3617,N_3873);
and U4485 (N_4485,N_3605,N_3776);
xnor U4486 (N_4486,N_3744,N_3678);
nor U4487 (N_4487,N_3859,N_3828);
nand U4488 (N_4488,N_3746,N_3676);
nor U4489 (N_4489,N_3956,N_3659);
or U4490 (N_4490,N_3750,N_3637);
nor U4491 (N_4491,N_3515,N_3832);
xor U4492 (N_4492,N_3889,N_3616);
and U4493 (N_4493,N_3587,N_3671);
or U4494 (N_4494,N_3707,N_3519);
nor U4495 (N_4495,N_3829,N_3960);
xnor U4496 (N_4496,N_3888,N_3650);
nand U4497 (N_4497,N_3984,N_3888);
and U4498 (N_4498,N_3544,N_3879);
nand U4499 (N_4499,N_3682,N_3851);
or U4500 (N_4500,N_4125,N_4144);
nand U4501 (N_4501,N_4283,N_4419);
xor U4502 (N_4502,N_4442,N_4090);
xor U4503 (N_4503,N_4321,N_4402);
xor U4504 (N_4504,N_4295,N_4223);
xor U4505 (N_4505,N_4207,N_4369);
xor U4506 (N_4506,N_4334,N_4398);
nor U4507 (N_4507,N_4226,N_4490);
nor U4508 (N_4508,N_4263,N_4439);
xor U4509 (N_4509,N_4141,N_4359);
nor U4510 (N_4510,N_4327,N_4497);
or U4511 (N_4511,N_4237,N_4469);
nand U4512 (N_4512,N_4244,N_4395);
nor U4513 (N_4513,N_4296,N_4115);
or U4514 (N_4514,N_4029,N_4139);
nand U4515 (N_4515,N_4026,N_4384);
nand U4516 (N_4516,N_4488,N_4265);
nand U4517 (N_4517,N_4380,N_4448);
or U4518 (N_4518,N_4375,N_4153);
or U4519 (N_4519,N_4192,N_4072);
or U4520 (N_4520,N_4007,N_4466);
and U4521 (N_4521,N_4053,N_4453);
nor U4522 (N_4522,N_4459,N_4008);
nor U4523 (N_4523,N_4270,N_4203);
and U4524 (N_4524,N_4422,N_4160);
and U4525 (N_4525,N_4087,N_4432);
nand U4526 (N_4526,N_4070,N_4117);
and U4527 (N_4527,N_4409,N_4037);
and U4528 (N_4528,N_4478,N_4483);
xor U4529 (N_4529,N_4039,N_4079);
and U4530 (N_4530,N_4062,N_4132);
nand U4531 (N_4531,N_4162,N_4371);
nand U4532 (N_4532,N_4475,N_4012);
xor U4533 (N_4533,N_4116,N_4157);
and U4534 (N_4534,N_4175,N_4074);
nor U4535 (N_4535,N_4433,N_4462);
or U4536 (N_4536,N_4282,N_4388);
xor U4537 (N_4537,N_4417,N_4121);
xor U4538 (N_4538,N_4251,N_4155);
or U4539 (N_4539,N_4047,N_4108);
xor U4540 (N_4540,N_4418,N_4260);
xor U4541 (N_4541,N_4014,N_4254);
nor U4542 (N_4542,N_4159,N_4069);
and U4543 (N_4543,N_4122,N_4022);
nor U4544 (N_4544,N_4335,N_4147);
nor U4545 (N_4545,N_4452,N_4127);
xnor U4546 (N_4546,N_4058,N_4236);
nand U4547 (N_4547,N_4294,N_4373);
or U4548 (N_4548,N_4305,N_4205);
and U4549 (N_4549,N_4013,N_4474);
xnor U4550 (N_4550,N_4403,N_4044);
nor U4551 (N_4551,N_4392,N_4233);
xor U4552 (N_4552,N_4183,N_4315);
and U4553 (N_4553,N_4225,N_4298);
nand U4554 (N_4554,N_4286,N_4397);
xor U4555 (N_4555,N_4146,N_4138);
xor U4556 (N_4556,N_4428,N_4168);
nand U4557 (N_4557,N_4293,N_4420);
or U4558 (N_4558,N_4498,N_4038);
or U4559 (N_4559,N_4342,N_4017);
and U4560 (N_4560,N_4479,N_4083);
xor U4561 (N_4561,N_4326,N_4274);
nand U4562 (N_4562,N_4352,N_4118);
xor U4563 (N_4563,N_4387,N_4345);
and U4564 (N_4564,N_4219,N_4246);
xnor U4565 (N_4565,N_4280,N_4241);
xor U4566 (N_4566,N_4336,N_4101);
or U4567 (N_4567,N_4458,N_4048);
xor U4568 (N_4568,N_4091,N_4455);
nand U4569 (N_4569,N_4361,N_4393);
nor U4570 (N_4570,N_4036,N_4487);
xnor U4571 (N_4571,N_4339,N_4094);
nor U4572 (N_4572,N_4229,N_4224);
or U4573 (N_4573,N_4316,N_4340);
and U4574 (N_4574,N_4003,N_4164);
or U4575 (N_4575,N_4399,N_4357);
nand U4576 (N_4576,N_4436,N_4285);
nor U4577 (N_4577,N_4093,N_4178);
nor U4578 (N_4578,N_4252,N_4460);
nor U4579 (N_4579,N_4346,N_4016);
nand U4580 (N_4580,N_4173,N_4319);
nor U4581 (N_4581,N_4234,N_4218);
xor U4582 (N_4582,N_4067,N_4322);
or U4583 (N_4583,N_4194,N_4080);
or U4584 (N_4584,N_4096,N_4228);
or U4585 (N_4585,N_4098,N_4005);
xnor U4586 (N_4586,N_4201,N_4112);
and U4587 (N_4587,N_4105,N_4377);
nand U4588 (N_4588,N_4411,N_4054);
and U4589 (N_4589,N_4120,N_4430);
or U4590 (N_4590,N_4358,N_4413);
and U4591 (N_4591,N_4231,N_4104);
nor U4592 (N_4592,N_4481,N_4347);
xor U4593 (N_4593,N_4291,N_4495);
xnor U4594 (N_4594,N_4063,N_4243);
or U4595 (N_4595,N_4140,N_4196);
nand U4596 (N_4596,N_4142,N_4467);
nor U4597 (N_4597,N_4214,N_4043);
xor U4598 (N_4598,N_4372,N_4208);
nand U4599 (N_4599,N_4440,N_4177);
xnor U4600 (N_4600,N_4416,N_4189);
xor U4601 (N_4601,N_4221,N_4386);
xor U4602 (N_4602,N_4126,N_4354);
nor U4603 (N_4603,N_4331,N_4249);
and U4604 (N_4604,N_4099,N_4493);
nand U4605 (N_4605,N_4077,N_4449);
nor U4606 (N_4606,N_4057,N_4222);
nor U4607 (N_4607,N_4206,N_4451);
xnor U4608 (N_4608,N_4482,N_4181);
xor U4609 (N_4609,N_4176,N_4367);
xor U4610 (N_4610,N_4353,N_4134);
nand U4611 (N_4611,N_4021,N_4020);
nor U4612 (N_4612,N_4006,N_4064);
and U4613 (N_4613,N_4267,N_4195);
or U4614 (N_4614,N_4076,N_4100);
xor U4615 (N_4615,N_4253,N_4349);
or U4616 (N_4616,N_4211,N_4033);
or U4617 (N_4617,N_4485,N_4425);
and U4618 (N_4618,N_4438,N_4097);
nor U4619 (N_4619,N_4227,N_4174);
nor U4620 (N_4620,N_4360,N_4133);
nand U4621 (N_4621,N_4281,N_4423);
nand U4622 (N_4622,N_4198,N_4001);
or U4623 (N_4623,N_4089,N_4102);
and U4624 (N_4624,N_4257,N_4179);
nor U4625 (N_4625,N_4341,N_4071);
xor U4626 (N_4626,N_4035,N_4250);
and U4627 (N_4627,N_4171,N_4492);
xnor U4628 (N_4628,N_4239,N_4051);
nand U4629 (N_4629,N_4193,N_4461);
and U4630 (N_4630,N_4473,N_4078);
or U4631 (N_4631,N_4052,N_4275);
or U4632 (N_4632,N_4400,N_4303);
nor U4633 (N_4633,N_4050,N_4318);
nand U4634 (N_4634,N_4042,N_4027);
nand U4635 (N_4635,N_4300,N_4216);
nor U4636 (N_4636,N_4385,N_4313);
or U4637 (N_4637,N_4412,N_4023);
xnor U4638 (N_4638,N_4103,N_4230);
nor U4639 (N_4639,N_4031,N_4232);
and U4640 (N_4640,N_4376,N_4289);
or U4641 (N_4641,N_4476,N_4025);
and U4642 (N_4642,N_4355,N_4145);
or U4643 (N_4643,N_4009,N_4030);
or U4644 (N_4644,N_4187,N_4032);
and U4645 (N_4645,N_4329,N_4266);
nand U4646 (N_4646,N_4041,N_4129);
xnor U4647 (N_4647,N_4435,N_4024);
nand U4648 (N_4648,N_4421,N_4337);
and U4649 (N_4649,N_4317,N_4150);
nand U4650 (N_4650,N_4163,N_4169);
xnor U4651 (N_4651,N_4499,N_4434);
nor U4652 (N_4652,N_4463,N_4262);
nand U4653 (N_4653,N_4068,N_4278);
nand U4654 (N_4654,N_4445,N_4055);
xnor U4655 (N_4655,N_4242,N_4310);
and U4656 (N_4656,N_4456,N_4004);
xnor U4657 (N_4657,N_4156,N_4287);
nor U4658 (N_4658,N_4343,N_4279);
nand U4659 (N_4659,N_4113,N_4363);
nand U4660 (N_4660,N_4111,N_4441);
and U4661 (N_4661,N_4396,N_4061);
xor U4662 (N_4662,N_4213,N_4084);
and U4663 (N_4663,N_4366,N_4060);
nor U4664 (N_4664,N_4209,N_4390);
and U4665 (N_4665,N_4269,N_4256);
or U4666 (N_4666,N_4086,N_4307);
nand U4667 (N_4667,N_4344,N_4191);
or U4668 (N_4668,N_4019,N_4365);
or U4669 (N_4669,N_4472,N_4235);
or U4670 (N_4670,N_4464,N_4370);
nand U4671 (N_4671,N_4161,N_4410);
and U4672 (N_4672,N_4381,N_4148);
or U4673 (N_4673,N_4407,N_4426);
xor U4674 (N_4674,N_4212,N_4268);
xor U4675 (N_4675,N_4301,N_4496);
and U4676 (N_4676,N_4220,N_4356);
xor U4677 (N_4677,N_4348,N_4477);
or U4678 (N_4678,N_4284,N_4170);
or U4679 (N_4679,N_4489,N_4325);
xnor U4680 (N_4680,N_4065,N_4180);
or U4681 (N_4681,N_4049,N_4172);
and U4682 (N_4682,N_4378,N_4314);
and U4683 (N_4683,N_4082,N_4130);
xnor U4684 (N_4684,N_4109,N_4202);
or U4685 (N_4685,N_4010,N_4107);
and U4686 (N_4686,N_4364,N_4018);
xor U4687 (N_4687,N_4081,N_4034);
nor U4688 (N_4688,N_4131,N_4288);
and U4689 (N_4689,N_4292,N_4330);
nand U4690 (N_4690,N_4471,N_4255);
and U4691 (N_4691,N_4092,N_4324);
xor U4692 (N_4692,N_4309,N_4190);
nor U4693 (N_4693,N_4088,N_4491);
nand U4694 (N_4694,N_4110,N_4240);
nor U4695 (N_4695,N_4320,N_4106);
xor U4696 (N_4696,N_4158,N_4167);
and U4697 (N_4697,N_4028,N_4323);
and U4698 (N_4698,N_4429,N_4186);
or U4699 (N_4699,N_4379,N_4272);
nor U4700 (N_4700,N_4200,N_4165);
nand U4701 (N_4701,N_4484,N_4450);
nand U4702 (N_4702,N_4182,N_4338);
or U4703 (N_4703,N_4188,N_4394);
xor U4704 (N_4704,N_4391,N_4304);
nand U4705 (N_4705,N_4143,N_4245);
nor U4706 (N_4706,N_4277,N_4470);
and U4707 (N_4707,N_4152,N_4351);
xor U4708 (N_4708,N_4415,N_4184);
nor U4709 (N_4709,N_4166,N_4261);
nand U4710 (N_4710,N_4271,N_4302);
nor U4711 (N_4711,N_4437,N_4238);
nand U4712 (N_4712,N_4408,N_4328);
and U4713 (N_4713,N_4486,N_4215);
nor U4714 (N_4714,N_4149,N_4414);
or U4715 (N_4715,N_4123,N_4075);
nor U4716 (N_4716,N_4114,N_4406);
nor U4717 (N_4717,N_4197,N_4154);
nand U4718 (N_4718,N_4312,N_4045);
nand U4719 (N_4719,N_4443,N_4002);
nand U4720 (N_4720,N_4446,N_4362);
xor U4721 (N_4721,N_4056,N_4494);
nor U4722 (N_4722,N_4468,N_4217);
or U4723 (N_4723,N_4066,N_4405);
or U4724 (N_4724,N_4308,N_4185);
and U4725 (N_4725,N_4306,N_4389);
or U4726 (N_4726,N_4444,N_4311);
nand U4727 (N_4727,N_4457,N_4136);
nand U4728 (N_4728,N_4258,N_4424);
and U4729 (N_4729,N_4374,N_4059);
and U4730 (N_4730,N_4137,N_4119);
and U4731 (N_4731,N_4383,N_4480);
and U4732 (N_4732,N_4259,N_4350);
nor U4733 (N_4733,N_4046,N_4015);
nand U4734 (N_4734,N_4427,N_4431);
xnor U4735 (N_4735,N_4095,N_4368);
xor U4736 (N_4736,N_4273,N_4247);
and U4737 (N_4737,N_4199,N_4382);
nor U4738 (N_4738,N_4297,N_4299);
nor U4739 (N_4739,N_4333,N_4135);
or U4740 (N_4740,N_4332,N_4085);
nand U4741 (N_4741,N_4404,N_4465);
xor U4742 (N_4742,N_4454,N_4447);
and U4743 (N_4743,N_4204,N_4264);
xor U4744 (N_4744,N_4011,N_4151);
and U4745 (N_4745,N_4040,N_4290);
or U4746 (N_4746,N_4248,N_4073);
xnor U4747 (N_4747,N_4124,N_4401);
or U4748 (N_4748,N_4276,N_4128);
xor U4749 (N_4749,N_4000,N_4210);
xor U4750 (N_4750,N_4212,N_4164);
nor U4751 (N_4751,N_4160,N_4390);
nand U4752 (N_4752,N_4186,N_4041);
nor U4753 (N_4753,N_4012,N_4018);
nor U4754 (N_4754,N_4071,N_4050);
and U4755 (N_4755,N_4001,N_4325);
and U4756 (N_4756,N_4440,N_4007);
or U4757 (N_4757,N_4172,N_4193);
or U4758 (N_4758,N_4363,N_4411);
nand U4759 (N_4759,N_4021,N_4009);
xor U4760 (N_4760,N_4370,N_4379);
or U4761 (N_4761,N_4314,N_4230);
nand U4762 (N_4762,N_4093,N_4157);
xor U4763 (N_4763,N_4174,N_4208);
or U4764 (N_4764,N_4225,N_4451);
xor U4765 (N_4765,N_4369,N_4459);
xor U4766 (N_4766,N_4409,N_4173);
nand U4767 (N_4767,N_4474,N_4304);
and U4768 (N_4768,N_4148,N_4225);
or U4769 (N_4769,N_4475,N_4468);
or U4770 (N_4770,N_4042,N_4176);
or U4771 (N_4771,N_4307,N_4152);
or U4772 (N_4772,N_4317,N_4430);
xnor U4773 (N_4773,N_4377,N_4115);
or U4774 (N_4774,N_4390,N_4311);
nand U4775 (N_4775,N_4397,N_4207);
and U4776 (N_4776,N_4406,N_4461);
nand U4777 (N_4777,N_4191,N_4384);
or U4778 (N_4778,N_4139,N_4468);
nor U4779 (N_4779,N_4131,N_4107);
nor U4780 (N_4780,N_4355,N_4054);
or U4781 (N_4781,N_4040,N_4411);
or U4782 (N_4782,N_4292,N_4428);
xnor U4783 (N_4783,N_4395,N_4455);
or U4784 (N_4784,N_4356,N_4187);
xor U4785 (N_4785,N_4147,N_4009);
nor U4786 (N_4786,N_4330,N_4063);
xnor U4787 (N_4787,N_4383,N_4264);
nor U4788 (N_4788,N_4396,N_4294);
nor U4789 (N_4789,N_4149,N_4358);
and U4790 (N_4790,N_4147,N_4314);
nand U4791 (N_4791,N_4257,N_4135);
or U4792 (N_4792,N_4147,N_4127);
nand U4793 (N_4793,N_4085,N_4123);
or U4794 (N_4794,N_4373,N_4422);
nand U4795 (N_4795,N_4260,N_4381);
nand U4796 (N_4796,N_4387,N_4239);
or U4797 (N_4797,N_4252,N_4136);
and U4798 (N_4798,N_4409,N_4376);
nand U4799 (N_4799,N_4075,N_4282);
xor U4800 (N_4800,N_4318,N_4119);
and U4801 (N_4801,N_4059,N_4130);
or U4802 (N_4802,N_4443,N_4132);
nand U4803 (N_4803,N_4209,N_4204);
nor U4804 (N_4804,N_4462,N_4104);
or U4805 (N_4805,N_4411,N_4190);
nor U4806 (N_4806,N_4095,N_4458);
nor U4807 (N_4807,N_4324,N_4179);
xnor U4808 (N_4808,N_4124,N_4339);
nor U4809 (N_4809,N_4195,N_4302);
or U4810 (N_4810,N_4314,N_4263);
nor U4811 (N_4811,N_4249,N_4351);
xor U4812 (N_4812,N_4144,N_4404);
xnor U4813 (N_4813,N_4466,N_4163);
nor U4814 (N_4814,N_4270,N_4324);
nor U4815 (N_4815,N_4245,N_4002);
nor U4816 (N_4816,N_4005,N_4111);
xnor U4817 (N_4817,N_4486,N_4169);
xnor U4818 (N_4818,N_4063,N_4385);
nor U4819 (N_4819,N_4147,N_4179);
or U4820 (N_4820,N_4417,N_4146);
nor U4821 (N_4821,N_4317,N_4425);
nor U4822 (N_4822,N_4099,N_4447);
and U4823 (N_4823,N_4041,N_4258);
and U4824 (N_4824,N_4381,N_4287);
and U4825 (N_4825,N_4390,N_4426);
xor U4826 (N_4826,N_4358,N_4006);
nand U4827 (N_4827,N_4093,N_4134);
and U4828 (N_4828,N_4019,N_4253);
nand U4829 (N_4829,N_4319,N_4242);
and U4830 (N_4830,N_4066,N_4059);
nand U4831 (N_4831,N_4122,N_4109);
and U4832 (N_4832,N_4314,N_4088);
nand U4833 (N_4833,N_4185,N_4123);
nor U4834 (N_4834,N_4039,N_4212);
xor U4835 (N_4835,N_4225,N_4460);
or U4836 (N_4836,N_4485,N_4089);
and U4837 (N_4837,N_4183,N_4373);
nor U4838 (N_4838,N_4065,N_4162);
xor U4839 (N_4839,N_4165,N_4072);
xor U4840 (N_4840,N_4139,N_4477);
or U4841 (N_4841,N_4060,N_4134);
nor U4842 (N_4842,N_4183,N_4094);
nand U4843 (N_4843,N_4436,N_4073);
nor U4844 (N_4844,N_4052,N_4449);
or U4845 (N_4845,N_4482,N_4465);
xor U4846 (N_4846,N_4261,N_4008);
xor U4847 (N_4847,N_4448,N_4400);
or U4848 (N_4848,N_4086,N_4199);
nand U4849 (N_4849,N_4042,N_4360);
nor U4850 (N_4850,N_4356,N_4218);
or U4851 (N_4851,N_4159,N_4441);
xnor U4852 (N_4852,N_4481,N_4134);
xor U4853 (N_4853,N_4416,N_4365);
xor U4854 (N_4854,N_4390,N_4178);
nor U4855 (N_4855,N_4249,N_4373);
nor U4856 (N_4856,N_4046,N_4401);
xor U4857 (N_4857,N_4262,N_4117);
nor U4858 (N_4858,N_4222,N_4234);
nor U4859 (N_4859,N_4468,N_4347);
or U4860 (N_4860,N_4339,N_4345);
xor U4861 (N_4861,N_4185,N_4206);
and U4862 (N_4862,N_4447,N_4104);
nor U4863 (N_4863,N_4196,N_4169);
or U4864 (N_4864,N_4166,N_4244);
and U4865 (N_4865,N_4421,N_4251);
xnor U4866 (N_4866,N_4189,N_4444);
xor U4867 (N_4867,N_4365,N_4398);
and U4868 (N_4868,N_4413,N_4077);
nand U4869 (N_4869,N_4467,N_4165);
nor U4870 (N_4870,N_4039,N_4151);
nor U4871 (N_4871,N_4478,N_4258);
xor U4872 (N_4872,N_4374,N_4350);
xnor U4873 (N_4873,N_4117,N_4316);
xor U4874 (N_4874,N_4487,N_4462);
and U4875 (N_4875,N_4368,N_4184);
and U4876 (N_4876,N_4393,N_4078);
and U4877 (N_4877,N_4154,N_4333);
and U4878 (N_4878,N_4184,N_4478);
nor U4879 (N_4879,N_4148,N_4271);
xor U4880 (N_4880,N_4043,N_4475);
and U4881 (N_4881,N_4136,N_4138);
and U4882 (N_4882,N_4215,N_4366);
xnor U4883 (N_4883,N_4358,N_4143);
nor U4884 (N_4884,N_4465,N_4334);
and U4885 (N_4885,N_4206,N_4169);
and U4886 (N_4886,N_4435,N_4236);
or U4887 (N_4887,N_4310,N_4327);
and U4888 (N_4888,N_4174,N_4455);
xor U4889 (N_4889,N_4319,N_4453);
nor U4890 (N_4890,N_4254,N_4366);
or U4891 (N_4891,N_4252,N_4348);
and U4892 (N_4892,N_4277,N_4463);
xnor U4893 (N_4893,N_4127,N_4076);
nand U4894 (N_4894,N_4132,N_4227);
xnor U4895 (N_4895,N_4331,N_4382);
and U4896 (N_4896,N_4490,N_4296);
nor U4897 (N_4897,N_4299,N_4029);
xor U4898 (N_4898,N_4302,N_4176);
nand U4899 (N_4899,N_4127,N_4237);
nand U4900 (N_4900,N_4107,N_4475);
or U4901 (N_4901,N_4229,N_4425);
and U4902 (N_4902,N_4426,N_4235);
xor U4903 (N_4903,N_4098,N_4010);
nor U4904 (N_4904,N_4131,N_4287);
xor U4905 (N_4905,N_4433,N_4380);
xor U4906 (N_4906,N_4157,N_4453);
xor U4907 (N_4907,N_4416,N_4053);
or U4908 (N_4908,N_4222,N_4325);
and U4909 (N_4909,N_4494,N_4382);
or U4910 (N_4910,N_4320,N_4034);
nand U4911 (N_4911,N_4316,N_4246);
xnor U4912 (N_4912,N_4440,N_4078);
or U4913 (N_4913,N_4209,N_4478);
nand U4914 (N_4914,N_4185,N_4255);
xor U4915 (N_4915,N_4273,N_4287);
nand U4916 (N_4916,N_4095,N_4069);
or U4917 (N_4917,N_4074,N_4251);
or U4918 (N_4918,N_4109,N_4421);
or U4919 (N_4919,N_4351,N_4469);
or U4920 (N_4920,N_4399,N_4293);
xnor U4921 (N_4921,N_4408,N_4219);
xnor U4922 (N_4922,N_4369,N_4024);
xor U4923 (N_4923,N_4144,N_4120);
nand U4924 (N_4924,N_4460,N_4058);
or U4925 (N_4925,N_4459,N_4142);
xnor U4926 (N_4926,N_4132,N_4105);
xnor U4927 (N_4927,N_4282,N_4112);
nor U4928 (N_4928,N_4253,N_4230);
nand U4929 (N_4929,N_4450,N_4378);
xnor U4930 (N_4930,N_4179,N_4331);
nand U4931 (N_4931,N_4377,N_4148);
nor U4932 (N_4932,N_4072,N_4019);
nand U4933 (N_4933,N_4325,N_4349);
and U4934 (N_4934,N_4268,N_4155);
nor U4935 (N_4935,N_4323,N_4061);
xnor U4936 (N_4936,N_4272,N_4360);
nand U4937 (N_4937,N_4099,N_4426);
nand U4938 (N_4938,N_4376,N_4238);
nand U4939 (N_4939,N_4025,N_4313);
xnor U4940 (N_4940,N_4037,N_4396);
or U4941 (N_4941,N_4084,N_4089);
xnor U4942 (N_4942,N_4312,N_4457);
nor U4943 (N_4943,N_4376,N_4021);
or U4944 (N_4944,N_4043,N_4136);
nor U4945 (N_4945,N_4183,N_4469);
or U4946 (N_4946,N_4446,N_4374);
or U4947 (N_4947,N_4394,N_4197);
nor U4948 (N_4948,N_4476,N_4197);
xor U4949 (N_4949,N_4256,N_4078);
or U4950 (N_4950,N_4347,N_4320);
nand U4951 (N_4951,N_4097,N_4141);
nor U4952 (N_4952,N_4279,N_4482);
and U4953 (N_4953,N_4344,N_4255);
nand U4954 (N_4954,N_4130,N_4091);
nand U4955 (N_4955,N_4432,N_4139);
nand U4956 (N_4956,N_4231,N_4309);
or U4957 (N_4957,N_4289,N_4322);
nand U4958 (N_4958,N_4119,N_4234);
xor U4959 (N_4959,N_4057,N_4328);
or U4960 (N_4960,N_4323,N_4414);
nand U4961 (N_4961,N_4036,N_4107);
or U4962 (N_4962,N_4228,N_4116);
nor U4963 (N_4963,N_4359,N_4443);
nand U4964 (N_4964,N_4226,N_4387);
and U4965 (N_4965,N_4486,N_4219);
xor U4966 (N_4966,N_4393,N_4215);
nand U4967 (N_4967,N_4411,N_4147);
nand U4968 (N_4968,N_4153,N_4332);
nor U4969 (N_4969,N_4341,N_4427);
or U4970 (N_4970,N_4355,N_4239);
or U4971 (N_4971,N_4211,N_4352);
xnor U4972 (N_4972,N_4298,N_4247);
or U4973 (N_4973,N_4137,N_4080);
xnor U4974 (N_4974,N_4265,N_4343);
xor U4975 (N_4975,N_4064,N_4324);
nand U4976 (N_4976,N_4319,N_4406);
xor U4977 (N_4977,N_4374,N_4486);
or U4978 (N_4978,N_4095,N_4232);
or U4979 (N_4979,N_4313,N_4330);
or U4980 (N_4980,N_4048,N_4072);
xnor U4981 (N_4981,N_4010,N_4369);
or U4982 (N_4982,N_4411,N_4211);
and U4983 (N_4983,N_4164,N_4152);
nor U4984 (N_4984,N_4487,N_4345);
nor U4985 (N_4985,N_4364,N_4147);
and U4986 (N_4986,N_4173,N_4251);
nor U4987 (N_4987,N_4236,N_4356);
nand U4988 (N_4988,N_4100,N_4207);
nand U4989 (N_4989,N_4230,N_4117);
or U4990 (N_4990,N_4302,N_4340);
nand U4991 (N_4991,N_4089,N_4389);
nand U4992 (N_4992,N_4063,N_4072);
nand U4993 (N_4993,N_4468,N_4379);
nor U4994 (N_4994,N_4460,N_4144);
xnor U4995 (N_4995,N_4234,N_4027);
nor U4996 (N_4996,N_4307,N_4297);
and U4997 (N_4997,N_4280,N_4405);
nand U4998 (N_4998,N_4188,N_4150);
nand U4999 (N_4999,N_4269,N_4163);
nor U5000 (N_5000,N_4626,N_4615);
nand U5001 (N_5001,N_4887,N_4653);
xnor U5002 (N_5002,N_4902,N_4972);
xnor U5003 (N_5003,N_4776,N_4666);
xnor U5004 (N_5004,N_4889,N_4517);
or U5005 (N_5005,N_4960,N_4511);
xor U5006 (N_5006,N_4981,N_4595);
and U5007 (N_5007,N_4967,N_4996);
and U5008 (N_5008,N_4513,N_4735);
xnor U5009 (N_5009,N_4877,N_4699);
nor U5010 (N_5010,N_4540,N_4624);
nor U5011 (N_5011,N_4806,N_4752);
or U5012 (N_5012,N_4682,N_4849);
or U5013 (N_5013,N_4733,N_4777);
nand U5014 (N_5014,N_4717,N_4828);
nand U5015 (N_5015,N_4893,N_4597);
nor U5016 (N_5016,N_4944,N_4696);
and U5017 (N_5017,N_4954,N_4724);
and U5018 (N_5018,N_4775,N_4676);
and U5019 (N_5019,N_4557,N_4690);
and U5020 (N_5020,N_4781,N_4876);
or U5021 (N_5021,N_4815,N_4727);
xnor U5022 (N_5022,N_4922,N_4942);
nand U5023 (N_5023,N_4501,N_4945);
or U5024 (N_5024,N_4659,N_4589);
xnor U5025 (N_5025,N_4612,N_4567);
and U5026 (N_5026,N_4951,N_4573);
or U5027 (N_5027,N_4519,N_4785);
and U5028 (N_5028,N_4587,N_4883);
nor U5029 (N_5029,N_4533,N_4535);
xnor U5030 (N_5030,N_4793,N_4962);
nor U5031 (N_5031,N_4641,N_4616);
or U5032 (N_5032,N_4753,N_4810);
xor U5033 (N_5033,N_4860,N_4576);
nand U5034 (N_5034,N_4681,N_4609);
nand U5035 (N_5035,N_4780,N_4614);
xnor U5036 (N_5036,N_4526,N_4644);
nand U5037 (N_5037,N_4739,N_4797);
and U5038 (N_5038,N_4854,N_4636);
nor U5039 (N_5039,N_4741,N_4697);
or U5040 (N_5040,N_4857,N_4961);
xor U5041 (N_5041,N_4886,N_4863);
nor U5042 (N_5042,N_4968,N_4610);
nand U5043 (N_5043,N_4756,N_4822);
or U5044 (N_5044,N_4904,N_4999);
xnor U5045 (N_5045,N_4670,N_4723);
nand U5046 (N_5046,N_4840,N_4901);
and U5047 (N_5047,N_4900,N_4584);
xnor U5048 (N_5048,N_4619,N_4873);
nand U5049 (N_5049,N_4834,N_4936);
nand U5050 (N_5050,N_4563,N_4649);
nor U5051 (N_5051,N_4665,N_4829);
xnor U5052 (N_5052,N_4928,N_4694);
and U5053 (N_5053,N_4508,N_4738);
nor U5054 (N_5054,N_4941,N_4695);
and U5055 (N_5055,N_4891,N_4599);
xor U5056 (N_5056,N_4805,N_4537);
or U5057 (N_5057,N_4570,N_4707);
xor U5058 (N_5058,N_4965,N_4506);
or U5059 (N_5059,N_4532,N_4946);
nor U5060 (N_5060,N_4939,N_4716);
and U5061 (N_5061,N_4835,N_4890);
and U5062 (N_5062,N_4958,N_4927);
and U5063 (N_5063,N_4850,N_4663);
or U5064 (N_5064,N_4705,N_4995);
and U5065 (N_5065,N_4825,N_4830);
nand U5066 (N_5066,N_4748,N_4955);
xnor U5067 (N_5067,N_4843,N_4948);
nor U5068 (N_5068,N_4507,N_4611);
xor U5069 (N_5069,N_4865,N_4648);
xnor U5070 (N_5070,N_4847,N_4868);
and U5071 (N_5071,N_4505,N_4711);
nand U5072 (N_5072,N_4767,N_4755);
nor U5073 (N_5073,N_4687,N_4879);
or U5074 (N_5074,N_4510,N_4866);
xor U5075 (N_5075,N_4754,N_4637);
nand U5076 (N_5076,N_4730,N_4527);
and U5077 (N_5077,N_4542,N_4977);
nand U5078 (N_5078,N_4565,N_4969);
nor U5079 (N_5079,N_4633,N_4926);
nand U5080 (N_5080,N_4924,N_4983);
nand U5081 (N_5081,N_4623,N_4971);
and U5082 (N_5082,N_4523,N_4861);
xnor U5083 (N_5083,N_4818,N_4832);
xor U5084 (N_5084,N_4745,N_4836);
nor U5085 (N_5085,N_4635,N_4545);
and U5086 (N_5086,N_4655,N_4602);
nand U5087 (N_5087,N_4638,N_4562);
nand U5088 (N_5088,N_4543,N_4575);
nand U5089 (N_5089,N_4817,N_4680);
nor U5090 (N_5090,N_4782,N_4598);
nand U5091 (N_5091,N_4524,N_4892);
and U5092 (N_5092,N_4862,N_4988);
and U5093 (N_5093,N_4980,N_4729);
nor U5094 (N_5094,N_4622,N_4952);
nor U5095 (N_5095,N_4558,N_4837);
and U5096 (N_5096,N_4959,N_4634);
nor U5097 (N_5097,N_4693,N_4908);
xnor U5098 (N_5098,N_4726,N_4544);
xor U5099 (N_5099,N_4888,N_4809);
nand U5100 (N_5100,N_4677,N_4600);
and U5101 (N_5101,N_4552,N_4645);
and U5102 (N_5102,N_4715,N_4783);
or U5103 (N_5103,N_4630,N_4798);
xnor U5104 (N_5104,N_4728,N_4931);
nor U5105 (N_5105,N_4606,N_4539);
xor U5106 (N_5106,N_4846,N_4502);
nand U5107 (N_5107,N_4974,N_4536);
nor U5108 (N_5108,N_4607,N_4702);
and U5109 (N_5109,N_4761,N_4827);
or U5110 (N_5110,N_4564,N_4521);
xor U5111 (N_5111,N_4773,N_4935);
or U5112 (N_5112,N_4559,N_4732);
and U5113 (N_5113,N_4566,N_4604);
nor U5114 (N_5114,N_4803,N_4885);
nand U5115 (N_5115,N_4763,N_4950);
nor U5116 (N_5116,N_4579,N_4642);
or U5117 (N_5117,N_4656,N_4672);
xnor U5118 (N_5118,N_4929,N_4758);
and U5119 (N_5119,N_4593,N_4821);
or U5120 (N_5120,N_4640,N_4875);
nand U5121 (N_5121,N_4590,N_4601);
xor U5122 (N_5122,N_4986,N_4736);
and U5123 (N_5123,N_4826,N_4578);
nor U5124 (N_5124,N_4743,N_4910);
xnor U5125 (N_5125,N_4720,N_4686);
or U5126 (N_5126,N_4842,N_4778);
and U5127 (N_5127,N_4975,N_4899);
and U5128 (N_5128,N_4966,N_4867);
or U5129 (N_5129,N_4963,N_4852);
nor U5130 (N_5130,N_4884,N_4794);
nand U5131 (N_5131,N_4799,N_4774);
xor U5132 (N_5132,N_4874,N_4800);
xor U5133 (N_5133,N_4770,N_4554);
nor U5134 (N_5134,N_4768,N_4631);
nor U5135 (N_5135,N_4594,N_4500);
or U5136 (N_5136,N_4920,N_4664);
nand U5137 (N_5137,N_4534,N_4700);
xor U5138 (N_5138,N_4779,N_4982);
or U5139 (N_5139,N_4549,N_4667);
and U5140 (N_5140,N_4679,N_4514);
nand U5141 (N_5141,N_4515,N_4701);
and U5142 (N_5142,N_4998,N_4762);
nor U5143 (N_5143,N_4674,N_4628);
xnor U5144 (N_5144,N_4940,N_4571);
or U5145 (N_5145,N_4586,N_4504);
nor U5146 (N_5146,N_4522,N_4790);
or U5147 (N_5147,N_4683,N_4871);
or U5148 (N_5148,N_4880,N_4831);
nand U5149 (N_5149,N_4646,N_4509);
or U5150 (N_5150,N_4786,N_4503);
xor U5151 (N_5151,N_4561,N_4529);
and U5152 (N_5152,N_4660,N_4851);
nand U5153 (N_5153,N_4807,N_4916);
or U5154 (N_5154,N_4569,N_4572);
or U5155 (N_5155,N_4629,N_4698);
xor U5156 (N_5156,N_4792,N_4719);
and U5157 (N_5157,N_4917,N_4930);
nand U5158 (N_5158,N_4546,N_4650);
or U5159 (N_5159,N_4744,N_4872);
nor U5160 (N_5160,N_4556,N_4788);
xor U5161 (N_5161,N_4978,N_4627);
or U5162 (N_5162,N_4751,N_4620);
and U5163 (N_5163,N_4956,N_4688);
nand U5164 (N_5164,N_4905,N_4613);
or U5165 (N_5165,N_4750,N_4734);
or U5166 (N_5166,N_4553,N_4881);
nand U5167 (N_5167,N_4765,N_4909);
and U5168 (N_5168,N_4772,N_4985);
and U5169 (N_5169,N_4903,N_4764);
nor U5170 (N_5170,N_4704,N_4555);
or U5171 (N_5171,N_4512,N_4516);
and U5172 (N_5172,N_4823,N_4560);
nand U5173 (N_5173,N_4551,N_4990);
nand U5174 (N_5174,N_4858,N_4964);
xnor U5175 (N_5175,N_4970,N_4538);
and U5176 (N_5176,N_4870,N_4824);
xnor U5177 (N_5177,N_4541,N_4808);
and U5178 (N_5178,N_4859,N_4918);
nor U5179 (N_5179,N_4662,N_4685);
nand U5180 (N_5180,N_4796,N_4617);
nand U5181 (N_5181,N_4991,N_4855);
nand U5182 (N_5182,N_4520,N_4819);
xnor U5183 (N_5183,N_4530,N_4947);
and U5184 (N_5184,N_4895,N_4742);
xor U5185 (N_5185,N_4864,N_4913);
or U5186 (N_5186,N_4596,N_4839);
nand U5187 (N_5187,N_4856,N_4771);
or U5188 (N_5188,N_4591,N_4784);
xor U5189 (N_5189,N_4993,N_4582);
nor U5190 (N_5190,N_4789,N_4923);
nor U5191 (N_5191,N_4643,N_4731);
xnor U5192 (N_5192,N_4992,N_4804);
xnor U5193 (N_5193,N_4976,N_4932);
nor U5194 (N_5194,N_4583,N_4907);
xor U5195 (N_5195,N_4746,N_4605);
or U5196 (N_5196,N_4713,N_4673);
or U5197 (N_5197,N_4737,N_4703);
or U5198 (N_5198,N_4618,N_4878);
and U5199 (N_5199,N_4925,N_4671);
nor U5200 (N_5200,N_4911,N_4897);
nand U5201 (N_5201,N_4749,N_4580);
xnor U5202 (N_5202,N_4957,N_4661);
or U5203 (N_5203,N_4984,N_4647);
nand U5204 (N_5204,N_4651,N_4848);
nand U5205 (N_5205,N_4548,N_4709);
nand U5206 (N_5206,N_4833,N_4791);
nor U5207 (N_5207,N_4938,N_4933);
xor U5208 (N_5208,N_4987,N_4937);
or U5209 (N_5209,N_4675,N_4853);
and U5210 (N_5210,N_4654,N_4816);
xor U5211 (N_5211,N_4531,N_4915);
and U5212 (N_5212,N_4801,N_4588);
and U5213 (N_5213,N_4625,N_4740);
and U5214 (N_5214,N_4639,N_4997);
and U5215 (N_5215,N_4657,N_4760);
xnor U5216 (N_5216,N_4652,N_4706);
xnor U5217 (N_5217,N_4994,N_4844);
and U5218 (N_5218,N_4919,N_4518);
or U5219 (N_5219,N_4898,N_4906);
nor U5220 (N_5220,N_4632,N_4795);
or U5221 (N_5221,N_4802,N_4550);
nor U5222 (N_5222,N_4766,N_4581);
nand U5223 (N_5223,N_4882,N_4691);
xor U5224 (N_5224,N_4525,N_4812);
or U5225 (N_5225,N_4896,N_4621);
or U5226 (N_5226,N_4714,N_4759);
nor U5227 (N_5227,N_4953,N_4841);
or U5228 (N_5228,N_4914,N_4814);
xor U5229 (N_5229,N_4547,N_4989);
xor U5230 (N_5230,N_4921,N_4592);
or U5231 (N_5231,N_4820,N_4668);
or U5232 (N_5232,N_4838,N_4722);
nand U5233 (N_5233,N_4568,N_4574);
xor U5234 (N_5234,N_4811,N_4712);
and U5235 (N_5235,N_4973,N_4585);
or U5236 (N_5236,N_4757,N_4658);
xor U5237 (N_5237,N_4678,N_4692);
or U5238 (N_5238,N_4725,N_4943);
nand U5239 (N_5239,N_4934,N_4710);
nor U5240 (N_5240,N_4528,N_4845);
nor U5241 (N_5241,N_4603,N_4669);
and U5242 (N_5242,N_4718,N_4747);
nand U5243 (N_5243,N_4813,N_4869);
and U5244 (N_5244,N_4721,N_4979);
and U5245 (N_5245,N_4577,N_4769);
nand U5246 (N_5246,N_4787,N_4689);
and U5247 (N_5247,N_4912,N_4894);
nor U5248 (N_5248,N_4949,N_4708);
nor U5249 (N_5249,N_4608,N_4684);
xor U5250 (N_5250,N_4948,N_4920);
or U5251 (N_5251,N_4857,N_4814);
and U5252 (N_5252,N_4716,N_4692);
xor U5253 (N_5253,N_4747,N_4734);
or U5254 (N_5254,N_4612,N_4695);
nor U5255 (N_5255,N_4964,N_4955);
nand U5256 (N_5256,N_4583,N_4589);
nor U5257 (N_5257,N_4609,N_4536);
nand U5258 (N_5258,N_4793,N_4891);
nor U5259 (N_5259,N_4579,N_4597);
nor U5260 (N_5260,N_4834,N_4880);
nand U5261 (N_5261,N_4540,N_4926);
and U5262 (N_5262,N_4935,N_4652);
nand U5263 (N_5263,N_4502,N_4925);
or U5264 (N_5264,N_4962,N_4661);
xnor U5265 (N_5265,N_4916,N_4978);
nor U5266 (N_5266,N_4598,N_4681);
and U5267 (N_5267,N_4978,N_4639);
and U5268 (N_5268,N_4804,N_4756);
and U5269 (N_5269,N_4710,N_4773);
nand U5270 (N_5270,N_4515,N_4541);
nand U5271 (N_5271,N_4800,N_4697);
xor U5272 (N_5272,N_4996,N_4810);
xor U5273 (N_5273,N_4635,N_4728);
xor U5274 (N_5274,N_4522,N_4563);
nor U5275 (N_5275,N_4523,N_4897);
nand U5276 (N_5276,N_4893,N_4768);
and U5277 (N_5277,N_4949,N_4678);
or U5278 (N_5278,N_4805,N_4891);
nand U5279 (N_5279,N_4571,N_4697);
xnor U5280 (N_5280,N_4685,N_4953);
nor U5281 (N_5281,N_4803,N_4516);
nor U5282 (N_5282,N_4851,N_4635);
and U5283 (N_5283,N_4562,N_4954);
xor U5284 (N_5284,N_4521,N_4892);
nand U5285 (N_5285,N_4874,N_4776);
or U5286 (N_5286,N_4954,N_4816);
nor U5287 (N_5287,N_4592,N_4804);
xor U5288 (N_5288,N_4607,N_4967);
nand U5289 (N_5289,N_4778,N_4599);
and U5290 (N_5290,N_4542,N_4823);
nor U5291 (N_5291,N_4574,N_4929);
and U5292 (N_5292,N_4578,N_4613);
or U5293 (N_5293,N_4541,N_4708);
and U5294 (N_5294,N_4819,N_4897);
and U5295 (N_5295,N_4977,N_4547);
nand U5296 (N_5296,N_4999,N_4692);
and U5297 (N_5297,N_4577,N_4567);
nand U5298 (N_5298,N_4540,N_4644);
nand U5299 (N_5299,N_4656,N_4963);
or U5300 (N_5300,N_4894,N_4932);
and U5301 (N_5301,N_4805,N_4540);
xor U5302 (N_5302,N_4708,N_4506);
and U5303 (N_5303,N_4610,N_4939);
nor U5304 (N_5304,N_4846,N_4528);
and U5305 (N_5305,N_4736,N_4649);
or U5306 (N_5306,N_4569,N_4927);
nand U5307 (N_5307,N_4673,N_4961);
nor U5308 (N_5308,N_4810,N_4627);
xnor U5309 (N_5309,N_4663,N_4692);
xor U5310 (N_5310,N_4685,N_4966);
nor U5311 (N_5311,N_4540,N_4734);
nand U5312 (N_5312,N_4990,N_4867);
nand U5313 (N_5313,N_4752,N_4812);
and U5314 (N_5314,N_4972,N_4833);
nand U5315 (N_5315,N_4972,N_4814);
and U5316 (N_5316,N_4727,N_4730);
or U5317 (N_5317,N_4940,N_4800);
nor U5318 (N_5318,N_4718,N_4982);
nor U5319 (N_5319,N_4823,N_4645);
nor U5320 (N_5320,N_4828,N_4562);
and U5321 (N_5321,N_4763,N_4773);
nand U5322 (N_5322,N_4831,N_4525);
and U5323 (N_5323,N_4712,N_4640);
nor U5324 (N_5324,N_4784,N_4799);
xnor U5325 (N_5325,N_4661,N_4734);
nor U5326 (N_5326,N_4600,N_4725);
or U5327 (N_5327,N_4921,N_4769);
xor U5328 (N_5328,N_4824,N_4861);
or U5329 (N_5329,N_4702,N_4517);
or U5330 (N_5330,N_4820,N_4794);
nor U5331 (N_5331,N_4541,N_4985);
or U5332 (N_5332,N_4751,N_4574);
nand U5333 (N_5333,N_4928,N_4626);
or U5334 (N_5334,N_4532,N_4828);
or U5335 (N_5335,N_4870,N_4923);
and U5336 (N_5336,N_4807,N_4500);
nor U5337 (N_5337,N_4826,N_4666);
nor U5338 (N_5338,N_4838,N_4996);
xor U5339 (N_5339,N_4950,N_4873);
xor U5340 (N_5340,N_4745,N_4681);
nor U5341 (N_5341,N_4873,N_4990);
nand U5342 (N_5342,N_4867,N_4515);
nand U5343 (N_5343,N_4575,N_4999);
and U5344 (N_5344,N_4771,N_4957);
nand U5345 (N_5345,N_4647,N_4981);
nor U5346 (N_5346,N_4573,N_4982);
and U5347 (N_5347,N_4680,N_4723);
and U5348 (N_5348,N_4861,N_4881);
xnor U5349 (N_5349,N_4549,N_4948);
or U5350 (N_5350,N_4869,N_4699);
and U5351 (N_5351,N_4793,N_4752);
and U5352 (N_5352,N_4623,N_4812);
and U5353 (N_5353,N_4888,N_4647);
xnor U5354 (N_5354,N_4619,N_4792);
or U5355 (N_5355,N_4836,N_4928);
and U5356 (N_5356,N_4829,N_4684);
nor U5357 (N_5357,N_4600,N_4506);
and U5358 (N_5358,N_4732,N_4793);
nand U5359 (N_5359,N_4578,N_4662);
nor U5360 (N_5360,N_4958,N_4643);
nand U5361 (N_5361,N_4870,N_4852);
nand U5362 (N_5362,N_4882,N_4816);
nand U5363 (N_5363,N_4734,N_4741);
nor U5364 (N_5364,N_4828,N_4610);
and U5365 (N_5365,N_4758,N_4747);
nor U5366 (N_5366,N_4682,N_4641);
nor U5367 (N_5367,N_4656,N_4698);
or U5368 (N_5368,N_4635,N_4526);
or U5369 (N_5369,N_4641,N_4649);
and U5370 (N_5370,N_4590,N_4840);
and U5371 (N_5371,N_4553,N_4724);
nand U5372 (N_5372,N_4753,N_4985);
or U5373 (N_5373,N_4574,N_4740);
nor U5374 (N_5374,N_4699,N_4584);
or U5375 (N_5375,N_4521,N_4970);
nand U5376 (N_5376,N_4717,N_4982);
nor U5377 (N_5377,N_4805,N_4530);
and U5378 (N_5378,N_4812,N_4643);
and U5379 (N_5379,N_4931,N_4774);
and U5380 (N_5380,N_4862,N_4585);
nor U5381 (N_5381,N_4739,N_4600);
nor U5382 (N_5382,N_4510,N_4685);
and U5383 (N_5383,N_4548,N_4808);
xor U5384 (N_5384,N_4836,N_4768);
and U5385 (N_5385,N_4581,N_4690);
and U5386 (N_5386,N_4664,N_4863);
nand U5387 (N_5387,N_4740,N_4524);
nand U5388 (N_5388,N_4625,N_4887);
xnor U5389 (N_5389,N_4601,N_4999);
and U5390 (N_5390,N_4646,N_4782);
xor U5391 (N_5391,N_4955,N_4822);
and U5392 (N_5392,N_4585,N_4991);
and U5393 (N_5393,N_4801,N_4863);
xnor U5394 (N_5394,N_4869,N_4508);
or U5395 (N_5395,N_4737,N_4835);
nor U5396 (N_5396,N_4708,N_4797);
or U5397 (N_5397,N_4811,N_4636);
or U5398 (N_5398,N_4514,N_4680);
nor U5399 (N_5399,N_4682,N_4645);
and U5400 (N_5400,N_4834,N_4815);
and U5401 (N_5401,N_4692,N_4960);
nand U5402 (N_5402,N_4813,N_4630);
or U5403 (N_5403,N_4602,N_4728);
xor U5404 (N_5404,N_4972,N_4811);
or U5405 (N_5405,N_4575,N_4898);
nand U5406 (N_5406,N_4804,N_4831);
nor U5407 (N_5407,N_4947,N_4674);
nor U5408 (N_5408,N_4511,N_4767);
and U5409 (N_5409,N_4924,N_4831);
xor U5410 (N_5410,N_4816,N_4697);
nor U5411 (N_5411,N_4805,N_4884);
nand U5412 (N_5412,N_4535,N_4796);
xnor U5413 (N_5413,N_4823,N_4818);
nand U5414 (N_5414,N_4929,N_4676);
nand U5415 (N_5415,N_4910,N_4986);
or U5416 (N_5416,N_4574,N_4987);
or U5417 (N_5417,N_4512,N_4902);
xnor U5418 (N_5418,N_4961,N_4893);
nand U5419 (N_5419,N_4755,N_4789);
and U5420 (N_5420,N_4579,N_4740);
or U5421 (N_5421,N_4837,N_4976);
nor U5422 (N_5422,N_4700,N_4968);
nor U5423 (N_5423,N_4515,N_4634);
or U5424 (N_5424,N_4944,N_4578);
xnor U5425 (N_5425,N_4984,N_4825);
or U5426 (N_5426,N_4814,N_4971);
and U5427 (N_5427,N_4547,N_4790);
xor U5428 (N_5428,N_4736,N_4662);
nor U5429 (N_5429,N_4784,N_4607);
nor U5430 (N_5430,N_4778,N_4621);
xnor U5431 (N_5431,N_4518,N_4572);
or U5432 (N_5432,N_4812,N_4924);
or U5433 (N_5433,N_4570,N_4801);
nor U5434 (N_5434,N_4541,N_4884);
or U5435 (N_5435,N_4835,N_4818);
or U5436 (N_5436,N_4687,N_4563);
and U5437 (N_5437,N_4511,N_4716);
xnor U5438 (N_5438,N_4910,N_4736);
and U5439 (N_5439,N_4785,N_4692);
or U5440 (N_5440,N_4942,N_4554);
or U5441 (N_5441,N_4785,N_4914);
xor U5442 (N_5442,N_4654,N_4906);
or U5443 (N_5443,N_4926,N_4584);
nand U5444 (N_5444,N_4655,N_4548);
xnor U5445 (N_5445,N_4685,N_4906);
or U5446 (N_5446,N_4553,N_4647);
nor U5447 (N_5447,N_4813,N_4931);
and U5448 (N_5448,N_4801,N_4950);
nor U5449 (N_5449,N_4670,N_4676);
and U5450 (N_5450,N_4895,N_4671);
nor U5451 (N_5451,N_4648,N_4730);
nor U5452 (N_5452,N_4710,N_4694);
and U5453 (N_5453,N_4587,N_4991);
or U5454 (N_5454,N_4570,N_4637);
or U5455 (N_5455,N_4728,N_4762);
nand U5456 (N_5456,N_4829,N_4934);
nor U5457 (N_5457,N_4667,N_4690);
nand U5458 (N_5458,N_4807,N_4545);
and U5459 (N_5459,N_4988,N_4775);
xor U5460 (N_5460,N_4757,N_4561);
nor U5461 (N_5461,N_4729,N_4748);
nor U5462 (N_5462,N_4612,N_4686);
and U5463 (N_5463,N_4974,N_4768);
and U5464 (N_5464,N_4729,N_4509);
nor U5465 (N_5465,N_4874,N_4617);
or U5466 (N_5466,N_4752,N_4662);
or U5467 (N_5467,N_4601,N_4663);
and U5468 (N_5468,N_4528,N_4869);
nand U5469 (N_5469,N_4556,N_4545);
xor U5470 (N_5470,N_4540,N_4942);
nor U5471 (N_5471,N_4975,N_4906);
nor U5472 (N_5472,N_4708,N_4777);
or U5473 (N_5473,N_4881,N_4790);
and U5474 (N_5474,N_4678,N_4793);
nor U5475 (N_5475,N_4792,N_4610);
nor U5476 (N_5476,N_4743,N_4586);
nand U5477 (N_5477,N_4535,N_4915);
or U5478 (N_5478,N_4880,N_4910);
xor U5479 (N_5479,N_4553,N_4947);
and U5480 (N_5480,N_4717,N_4963);
or U5481 (N_5481,N_4791,N_4618);
or U5482 (N_5482,N_4779,N_4576);
nand U5483 (N_5483,N_4682,N_4792);
or U5484 (N_5484,N_4574,N_4961);
and U5485 (N_5485,N_4884,N_4813);
or U5486 (N_5486,N_4895,N_4554);
nand U5487 (N_5487,N_4712,N_4652);
and U5488 (N_5488,N_4500,N_4714);
nor U5489 (N_5489,N_4853,N_4896);
or U5490 (N_5490,N_4778,N_4872);
and U5491 (N_5491,N_4664,N_4652);
and U5492 (N_5492,N_4579,N_4630);
nor U5493 (N_5493,N_4841,N_4739);
and U5494 (N_5494,N_4532,N_4658);
or U5495 (N_5495,N_4523,N_4888);
xor U5496 (N_5496,N_4747,N_4902);
or U5497 (N_5497,N_4772,N_4681);
nor U5498 (N_5498,N_4957,N_4558);
and U5499 (N_5499,N_4624,N_4834);
xnor U5500 (N_5500,N_5319,N_5046);
or U5501 (N_5501,N_5404,N_5010);
or U5502 (N_5502,N_5284,N_5176);
nor U5503 (N_5503,N_5166,N_5138);
or U5504 (N_5504,N_5260,N_5235);
or U5505 (N_5505,N_5106,N_5208);
xor U5506 (N_5506,N_5369,N_5354);
nor U5507 (N_5507,N_5253,N_5469);
and U5508 (N_5508,N_5024,N_5121);
xnor U5509 (N_5509,N_5108,N_5221);
nand U5510 (N_5510,N_5393,N_5009);
or U5511 (N_5511,N_5465,N_5174);
nand U5512 (N_5512,N_5231,N_5136);
or U5513 (N_5513,N_5325,N_5360);
and U5514 (N_5514,N_5190,N_5335);
nor U5515 (N_5515,N_5286,N_5130);
and U5516 (N_5516,N_5264,N_5448);
nor U5517 (N_5517,N_5498,N_5236);
nor U5518 (N_5518,N_5409,N_5116);
or U5519 (N_5519,N_5328,N_5275);
nand U5520 (N_5520,N_5165,N_5449);
nand U5521 (N_5521,N_5445,N_5374);
and U5522 (N_5522,N_5279,N_5234);
xor U5523 (N_5523,N_5471,N_5333);
nor U5524 (N_5524,N_5071,N_5431);
nand U5525 (N_5525,N_5497,N_5287);
or U5526 (N_5526,N_5371,N_5454);
and U5527 (N_5527,N_5285,N_5394);
and U5528 (N_5528,N_5062,N_5340);
and U5529 (N_5529,N_5467,N_5400);
or U5530 (N_5530,N_5204,N_5159);
nand U5531 (N_5531,N_5091,N_5178);
or U5532 (N_5532,N_5154,N_5455);
or U5533 (N_5533,N_5392,N_5044);
or U5534 (N_5534,N_5278,N_5385);
nand U5535 (N_5535,N_5429,N_5492);
nand U5536 (N_5536,N_5306,N_5050);
and U5537 (N_5537,N_5148,N_5119);
xnor U5538 (N_5538,N_5143,N_5086);
or U5539 (N_5539,N_5414,N_5035);
and U5540 (N_5540,N_5218,N_5053);
or U5541 (N_5541,N_5270,N_5037);
xnor U5542 (N_5542,N_5216,N_5293);
or U5543 (N_5543,N_5280,N_5334);
and U5544 (N_5544,N_5161,N_5141);
nand U5545 (N_5545,N_5361,N_5418);
xor U5546 (N_5546,N_5380,N_5348);
xor U5547 (N_5547,N_5080,N_5359);
xnor U5548 (N_5548,N_5459,N_5002);
nor U5549 (N_5549,N_5479,N_5470);
xnor U5550 (N_5550,N_5382,N_5100);
nand U5551 (N_5551,N_5255,N_5489);
nand U5552 (N_5552,N_5128,N_5312);
nand U5553 (N_5553,N_5281,N_5142);
and U5554 (N_5554,N_5115,N_5257);
nand U5555 (N_5555,N_5324,N_5378);
xor U5556 (N_5556,N_5242,N_5343);
or U5557 (N_5557,N_5314,N_5038);
xor U5558 (N_5558,N_5363,N_5329);
xnor U5559 (N_5559,N_5464,N_5357);
and U5560 (N_5560,N_5188,N_5277);
nand U5561 (N_5561,N_5177,N_5132);
xnor U5562 (N_5562,N_5366,N_5391);
and U5563 (N_5563,N_5456,N_5070);
and U5564 (N_5564,N_5321,N_5230);
nand U5565 (N_5565,N_5107,N_5039);
and U5566 (N_5566,N_5054,N_5346);
or U5567 (N_5567,N_5384,N_5043);
or U5568 (N_5568,N_5463,N_5135);
and U5569 (N_5569,N_5376,N_5105);
nor U5570 (N_5570,N_5494,N_5124);
or U5571 (N_5571,N_5152,N_5205);
nor U5572 (N_5572,N_5092,N_5004);
nand U5573 (N_5573,N_5118,N_5224);
or U5574 (N_5574,N_5447,N_5308);
nand U5575 (N_5575,N_5090,N_5273);
and U5576 (N_5576,N_5422,N_5491);
nand U5577 (N_5577,N_5434,N_5087);
or U5578 (N_5578,N_5327,N_5261);
or U5579 (N_5579,N_5020,N_5432);
nor U5580 (N_5580,N_5297,N_5419);
nor U5581 (N_5581,N_5453,N_5396);
or U5582 (N_5582,N_5149,N_5219);
and U5583 (N_5583,N_5248,N_5114);
xnor U5584 (N_5584,N_5078,N_5095);
or U5585 (N_5585,N_5215,N_5322);
and U5586 (N_5586,N_5067,N_5077);
xor U5587 (N_5587,N_5049,N_5424);
and U5588 (N_5588,N_5047,N_5075);
or U5589 (N_5589,N_5304,N_5232);
nor U5590 (N_5590,N_5294,N_5249);
nor U5591 (N_5591,N_5162,N_5401);
and U5592 (N_5592,N_5478,N_5330);
nor U5593 (N_5593,N_5341,N_5290);
nand U5594 (N_5594,N_5191,N_5407);
xor U5595 (N_5595,N_5229,N_5405);
xor U5596 (N_5596,N_5256,N_5225);
and U5597 (N_5597,N_5093,N_5320);
xor U5598 (N_5598,N_5250,N_5496);
nand U5599 (N_5599,N_5423,N_5227);
and U5600 (N_5600,N_5417,N_5182);
nor U5601 (N_5601,N_5365,N_5458);
xnor U5602 (N_5602,N_5164,N_5094);
or U5603 (N_5603,N_5019,N_5487);
or U5604 (N_5604,N_5157,N_5355);
or U5605 (N_5605,N_5347,N_5103);
xnor U5606 (N_5606,N_5018,N_5473);
nand U5607 (N_5607,N_5362,N_5084);
nand U5608 (N_5608,N_5042,N_5339);
and U5609 (N_5609,N_5207,N_5315);
and U5610 (N_5610,N_5307,N_5083);
xnor U5611 (N_5611,N_5033,N_5263);
nor U5612 (N_5612,N_5029,N_5451);
and U5613 (N_5613,N_5425,N_5126);
or U5614 (N_5614,N_5428,N_5476);
and U5615 (N_5615,N_5021,N_5433);
or U5616 (N_5616,N_5001,N_5301);
nand U5617 (N_5617,N_5298,N_5482);
xor U5618 (N_5618,N_5233,N_5475);
and U5619 (N_5619,N_5056,N_5140);
nor U5620 (N_5620,N_5079,N_5197);
nor U5621 (N_5621,N_5439,N_5151);
nor U5622 (N_5622,N_5317,N_5436);
nand U5623 (N_5623,N_5055,N_5254);
and U5624 (N_5624,N_5012,N_5258);
nand U5625 (N_5625,N_5032,N_5125);
nand U5626 (N_5626,N_5303,N_5222);
and U5627 (N_5627,N_5377,N_5201);
xor U5628 (N_5628,N_5367,N_5403);
nor U5629 (N_5629,N_5438,N_5446);
xnor U5630 (N_5630,N_5203,N_5379);
and U5631 (N_5631,N_5063,N_5052);
and U5632 (N_5632,N_5060,N_5192);
xor U5633 (N_5633,N_5402,N_5206);
nor U5634 (N_5634,N_5210,N_5059);
nor U5635 (N_5635,N_5170,N_5408);
nand U5636 (N_5636,N_5189,N_5241);
or U5637 (N_5637,N_5299,N_5318);
xor U5638 (N_5638,N_5295,N_5370);
and U5639 (N_5639,N_5416,N_5477);
xor U5640 (N_5640,N_5072,N_5238);
nor U5641 (N_5641,N_5336,N_5326);
nand U5642 (N_5642,N_5276,N_5274);
xor U5643 (N_5643,N_5111,N_5430);
or U5644 (N_5644,N_5167,N_5171);
nor U5645 (N_5645,N_5386,N_5183);
and U5646 (N_5646,N_5082,N_5110);
or U5647 (N_5647,N_5443,N_5244);
xnor U5648 (N_5648,N_5265,N_5389);
nand U5649 (N_5649,N_5472,N_5123);
nor U5650 (N_5650,N_5466,N_5160);
nand U5651 (N_5651,N_5495,N_5102);
nand U5652 (N_5652,N_5209,N_5017);
nor U5653 (N_5653,N_5368,N_5185);
and U5654 (N_5654,N_5351,N_5342);
or U5655 (N_5655,N_5006,N_5096);
nor U5656 (N_5656,N_5015,N_5169);
xnor U5657 (N_5657,N_5112,N_5145);
or U5658 (N_5658,N_5271,N_5283);
and U5659 (N_5659,N_5193,N_5031);
and U5660 (N_5660,N_5202,N_5133);
xor U5661 (N_5661,N_5442,N_5099);
xor U5662 (N_5662,N_5127,N_5023);
or U5663 (N_5663,N_5117,N_5129);
xnor U5664 (N_5664,N_5291,N_5440);
and U5665 (N_5665,N_5486,N_5139);
or U5666 (N_5666,N_5187,N_5410);
and U5667 (N_5667,N_5034,N_5251);
xor U5668 (N_5668,N_5228,N_5484);
and U5669 (N_5669,N_5337,N_5252);
nand U5670 (N_5670,N_5057,N_5302);
and U5671 (N_5671,N_5457,N_5296);
nor U5672 (N_5672,N_5247,N_5485);
or U5673 (N_5673,N_5122,N_5309);
or U5674 (N_5674,N_5134,N_5350);
nor U5675 (N_5675,N_5217,N_5068);
nand U5676 (N_5676,N_5113,N_5088);
and U5677 (N_5677,N_5172,N_5040);
xnor U5678 (N_5678,N_5499,N_5226);
nand U5679 (N_5679,N_5313,N_5069);
or U5680 (N_5680,N_5311,N_5437);
and U5681 (N_5681,N_5461,N_5013);
and U5682 (N_5682,N_5267,N_5364);
nand U5683 (N_5683,N_5268,N_5011);
or U5684 (N_5684,N_5194,N_5098);
nor U5685 (N_5685,N_5353,N_5289);
and U5686 (N_5686,N_5007,N_5196);
nand U5687 (N_5687,N_5156,N_5213);
xor U5688 (N_5688,N_5181,N_5008);
xnor U5689 (N_5689,N_5237,N_5460);
nand U5690 (N_5690,N_5358,N_5173);
xor U5691 (N_5691,N_5085,N_5051);
nor U5692 (N_5692,N_5005,N_5488);
nand U5693 (N_5693,N_5199,N_5421);
nand U5694 (N_5694,N_5345,N_5089);
nor U5695 (N_5695,N_5045,N_5109);
nor U5696 (N_5696,N_5387,N_5212);
or U5697 (N_5697,N_5323,N_5398);
nand U5698 (N_5698,N_5066,N_5305);
and U5699 (N_5699,N_5146,N_5468);
or U5700 (N_5700,N_5144,N_5406);
and U5701 (N_5701,N_5027,N_5356);
xor U5702 (N_5702,N_5158,N_5101);
nor U5703 (N_5703,N_5184,N_5214);
or U5704 (N_5704,N_5061,N_5344);
and U5705 (N_5705,N_5450,N_5331);
nor U5706 (N_5706,N_5220,N_5081);
or U5707 (N_5707,N_5474,N_5014);
and U5708 (N_5708,N_5316,N_5420);
nand U5709 (N_5709,N_5399,N_5168);
or U5710 (N_5710,N_5462,N_5211);
nor U5711 (N_5711,N_5065,N_5016);
or U5712 (N_5712,N_5383,N_5239);
nor U5713 (N_5713,N_5003,N_5452);
or U5714 (N_5714,N_5163,N_5246);
or U5715 (N_5715,N_5180,N_5435);
nor U5716 (N_5716,N_5076,N_5349);
nor U5717 (N_5717,N_5375,N_5153);
and U5718 (N_5718,N_5397,N_5155);
or U5719 (N_5719,N_5272,N_5381);
and U5720 (N_5720,N_5058,N_5022);
nand U5721 (N_5721,N_5372,N_5395);
and U5722 (N_5722,N_5310,N_5292);
xnor U5723 (N_5723,N_5444,N_5412);
or U5724 (N_5724,N_5259,N_5137);
nor U5725 (N_5725,N_5048,N_5390);
nor U5726 (N_5726,N_5000,N_5411);
xnor U5727 (N_5727,N_5373,N_5097);
nor U5728 (N_5728,N_5198,N_5240);
or U5729 (N_5729,N_5426,N_5104);
nand U5730 (N_5730,N_5441,N_5288);
nand U5731 (N_5731,N_5282,N_5036);
nand U5732 (N_5732,N_5415,N_5223);
nand U5733 (N_5733,N_5200,N_5064);
nand U5734 (N_5734,N_5266,N_5332);
nor U5735 (N_5735,N_5041,N_5427);
and U5736 (N_5736,N_5245,N_5269);
nor U5737 (N_5737,N_5480,N_5179);
xor U5738 (N_5738,N_5074,N_5150);
nand U5739 (N_5739,N_5025,N_5338);
nor U5740 (N_5740,N_5483,N_5388);
or U5741 (N_5741,N_5243,N_5147);
xor U5742 (N_5742,N_5175,N_5262);
nor U5743 (N_5743,N_5300,N_5352);
xor U5744 (N_5744,N_5120,N_5131);
xnor U5745 (N_5745,N_5493,N_5413);
nand U5746 (N_5746,N_5186,N_5026);
nor U5747 (N_5747,N_5030,N_5073);
xor U5748 (N_5748,N_5195,N_5490);
or U5749 (N_5749,N_5481,N_5028);
nor U5750 (N_5750,N_5453,N_5480);
nor U5751 (N_5751,N_5112,N_5101);
or U5752 (N_5752,N_5241,N_5201);
or U5753 (N_5753,N_5160,N_5401);
or U5754 (N_5754,N_5156,N_5270);
nand U5755 (N_5755,N_5171,N_5249);
nor U5756 (N_5756,N_5189,N_5329);
nor U5757 (N_5757,N_5035,N_5232);
nand U5758 (N_5758,N_5245,N_5338);
xnor U5759 (N_5759,N_5004,N_5389);
nand U5760 (N_5760,N_5146,N_5178);
or U5761 (N_5761,N_5276,N_5393);
nand U5762 (N_5762,N_5302,N_5426);
nand U5763 (N_5763,N_5148,N_5009);
or U5764 (N_5764,N_5346,N_5487);
nor U5765 (N_5765,N_5130,N_5309);
or U5766 (N_5766,N_5186,N_5132);
xor U5767 (N_5767,N_5233,N_5358);
nor U5768 (N_5768,N_5421,N_5184);
xnor U5769 (N_5769,N_5343,N_5488);
nor U5770 (N_5770,N_5209,N_5342);
nand U5771 (N_5771,N_5493,N_5136);
and U5772 (N_5772,N_5266,N_5313);
nor U5773 (N_5773,N_5283,N_5077);
nor U5774 (N_5774,N_5355,N_5280);
xor U5775 (N_5775,N_5122,N_5014);
xor U5776 (N_5776,N_5464,N_5117);
nor U5777 (N_5777,N_5023,N_5104);
xor U5778 (N_5778,N_5227,N_5452);
nor U5779 (N_5779,N_5369,N_5027);
nor U5780 (N_5780,N_5139,N_5167);
nor U5781 (N_5781,N_5103,N_5312);
or U5782 (N_5782,N_5344,N_5295);
nand U5783 (N_5783,N_5496,N_5069);
nand U5784 (N_5784,N_5295,N_5393);
nand U5785 (N_5785,N_5093,N_5035);
and U5786 (N_5786,N_5462,N_5156);
xnor U5787 (N_5787,N_5032,N_5191);
and U5788 (N_5788,N_5185,N_5240);
xnor U5789 (N_5789,N_5467,N_5364);
xnor U5790 (N_5790,N_5230,N_5311);
and U5791 (N_5791,N_5273,N_5012);
nand U5792 (N_5792,N_5397,N_5323);
nand U5793 (N_5793,N_5384,N_5434);
xor U5794 (N_5794,N_5169,N_5420);
xor U5795 (N_5795,N_5255,N_5083);
nand U5796 (N_5796,N_5458,N_5383);
and U5797 (N_5797,N_5395,N_5251);
xor U5798 (N_5798,N_5342,N_5334);
nand U5799 (N_5799,N_5121,N_5260);
and U5800 (N_5800,N_5498,N_5141);
nand U5801 (N_5801,N_5224,N_5317);
or U5802 (N_5802,N_5411,N_5385);
and U5803 (N_5803,N_5416,N_5376);
xnor U5804 (N_5804,N_5095,N_5009);
xnor U5805 (N_5805,N_5478,N_5137);
nand U5806 (N_5806,N_5314,N_5071);
xor U5807 (N_5807,N_5472,N_5092);
xor U5808 (N_5808,N_5317,N_5346);
and U5809 (N_5809,N_5054,N_5163);
or U5810 (N_5810,N_5177,N_5309);
nor U5811 (N_5811,N_5349,N_5348);
xor U5812 (N_5812,N_5092,N_5289);
xor U5813 (N_5813,N_5051,N_5271);
nand U5814 (N_5814,N_5098,N_5246);
nor U5815 (N_5815,N_5466,N_5265);
nand U5816 (N_5816,N_5463,N_5196);
xnor U5817 (N_5817,N_5306,N_5243);
or U5818 (N_5818,N_5400,N_5334);
nand U5819 (N_5819,N_5263,N_5378);
nor U5820 (N_5820,N_5497,N_5260);
and U5821 (N_5821,N_5035,N_5421);
and U5822 (N_5822,N_5134,N_5289);
or U5823 (N_5823,N_5409,N_5267);
nor U5824 (N_5824,N_5255,N_5021);
xnor U5825 (N_5825,N_5110,N_5322);
or U5826 (N_5826,N_5210,N_5170);
nand U5827 (N_5827,N_5342,N_5082);
and U5828 (N_5828,N_5220,N_5103);
or U5829 (N_5829,N_5031,N_5394);
or U5830 (N_5830,N_5023,N_5007);
or U5831 (N_5831,N_5367,N_5249);
or U5832 (N_5832,N_5499,N_5306);
nand U5833 (N_5833,N_5431,N_5018);
xnor U5834 (N_5834,N_5272,N_5348);
and U5835 (N_5835,N_5116,N_5130);
or U5836 (N_5836,N_5454,N_5118);
xor U5837 (N_5837,N_5239,N_5465);
and U5838 (N_5838,N_5350,N_5405);
nand U5839 (N_5839,N_5169,N_5129);
nor U5840 (N_5840,N_5349,N_5235);
nor U5841 (N_5841,N_5012,N_5172);
or U5842 (N_5842,N_5079,N_5242);
nor U5843 (N_5843,N_5066,N_5434);
nor U5844 (N_5844,N_5407,N_5468);
and U5845 (N_5845,N_5448,N_5330);
or U5846 (N_5846,N_5065,N_5055);
nand U5847 (N_5847,N_5455,N_5446);
nand U5848 (N_5848,N_5023,N_5486);
xnor U5849 (N_5849,N_5454,N_5165);
or U5850 (N_5850,N_5194,N_5053);
and U5851 (N_5851,N_5363,N_5060);
and U5852 (N_5852,N_5437,N_5332);
and U5853 (N_5853,N_5169,N_5334);
or U5854 (N_5854,N_5054,N_5295);
nand U5855 (N_5855,N_5209,N_5370);
nor U5856 (N_5856,N_5080,N_5420);
nand U5857 (N_5857,N_5273,N_5255);
nor U5858 (N_5858,N_5011,N_5333);
nor U5859 (N_5859,N_5255,N_5334);
or U5860 (N_5860,N_5212,N_5362);
or U5861 (N_5861,N_5122,N_5267);
and U5862 (N_5862,N_5415,N_5023);
or U5863 (N_5863,N_5344,N_5069);
nor U5864 (N_5864,N_5316,N_5010);
nor U5865 (N_5865,N_5013,N_5407);
and U5866 (N_5866,N_5017,N_5109);
and U5867 (N_5867,N_5102,N_5008);
nand U5868 (N_5868,N_5457,N_5066);
xor U5869 (N_5869,N_5450,N_5078);
or U5870 (N_5870,N_5189,N_5423);
xor U5871 (N_5871,N_5371,N_5168);
xor U5872 (N_5872,N_5248,N_5231);
nor U5873 (N_5873,N_5350,N_5351);
xor U5874 (N_5874,N_5288,N_5450);
and U5875 (N_5875,N_5440,N_5061);
nor U5876 (N_5876,N_5475,N_5419);
and U5877 (N_5877,N_5462,N_5319);
and U5878 (N_5878,N_5209,N_5182);
or U5879 (N_5879,N_5435,N_5385);
xor U5880 (N_5880,N_5328,N_5454);
nand U5881 (N_5881,N_5001,N_5104);
or U5882 (N_5882,N_5421,N_5033);
nand U5883 (N_5883,N_5351,N_5166);
nand U5884 (N_5884,N_5037,N_5040);
and U5885 (N_5885,N_5088,N_5335);
or U5886 (N_5886,N_5089,N_5432);
nand U5887 (N_5887,N_5340,N_5472);
xnor U5888 (N_5888,N_5386,N_5365);
and U5889 (N_5889,N_5159,N_5099);
nand U5890 (N_5890,N_5067,N_5054);
nand U5891 (N_5891,N_5180,N_5097);
xnor U5892 (N_5892,N_5249,N_5299);
and U5893 (N_5893,N_5133,N_5455);
nor U5894 (N_5894,N_5241,N_5228);
or U5895 (N_5895,N_5436,N_5416);
nand U5896 (N_5896,N_5484,N_5492);
and U5897 (N_5897,N_5462,N_5443);
or U5898 (N_5898,N_5051,N_5451);
xnor U5899 (N_5899,N_5413,N_5222);
and U5900 (N_5900,N_5146,N_5357);
or U5901 (N_5901,N_5432,N_5293);
xor U5902 (N_5902,N_5192,N_5049);
nor U5903 (N_5903,N_5204,N_5373);
nor U5904 (N_5904,N_5304,N_5262);
xor U5905 (N_5905,N_5101,N_5177);
and U5906 (N_5906,N_5426,N_5151);
and U5907 (N_5907,N_5237,N_5359);
and U5908 (N_5908,N_5495,N_5343);
nor U5909 (N_5909,N_5426,N_5381);
and U5910 (N_5910,N_5451,N_5353);
nand U5911 (N_5911,N_5141,N_5169);
nand U5912 (N_5912,N_5080,N_5121);
nand U5913 (N_5913,N_5256,N_5069);
xnor U5914 (N_5914,N_5200,N_5025);
xnor U5915 (N_5915,N_5187,N_5269);
and U5916 (N_5916,N_5223,N_5300);
and U5917 (N_5917,N_5212,N_5048);
nor U5918 (N_5918,N_5179,N_5241);
xnor U5919 (N_5919,N_5023,N_5424);
nand U5920 (N_5920,N_5318,N_5099);
or U5921 (N_5921,N_5112,N_5497);
and U5922 (N_5922,N_5190,N_5101);
xor U5923 (N_5923,N_5130,N_5170);
xnor U5924 (N_5924,N_5497,N_5454);
nor U5925 (N_5925,N_5039,N_5420);
and U5926 (N_5926,N_5054,N_5397);
or U5927 (N_5927,N_5303,N_5314);
nand U5928 (N_5928,N_5279,N_5347);
nand U5929 (N_5929,N_5333,N_5416);
nor U5930 (N_5930,N_5277,N_5143);
and U5931 (N_5931,N_5005,N_5214);
xnor U5932 (N_5932,N_5401,N_5332);
xnor U5933 (N_5933,N_5118,N_5230);
nand U5934 (N_5934,N_5130,N_5473);
nor U5935 (N_5935,N_5374,N_5289);
nand U5936 (N_5936,N_5076,N_5131);
and U5937 (N_5937,N_5215,N_5136);
xor U5938 (N_5938,N_5395,N_5183);
and U5939 (N_5939,N_5036,N_5290);
and U5940 (N_5940,N_5359,N_5171);
xnor U5941 (N_5941,N_5365,N_5215);
xor U5942 (N_5942,N_5111,N_5265);
and U5943 (N_5943,N_5004,N_5404);
nand U5944 (N_5944,N_5356,N_5470);
or U5945 (N_5945,N_5469,N_5216);
xor U5946 (N_5946,N_5201,N_5187);
and U5947 (N_5947,N_5126,N_5019);
xor U5948 (N_5948,N_5435,N_5263);
xor U5949 (N_5949,N_5048,N_5164);
or U5950 (N_5950,N_5256,N_5260);
nor U5951 (N_5951,N_5089,N_5389);
xor U5952 (N_5952,N_5393,N_5394);
nand U5953 (N_5953,N_5178,N_5493);
or U5954 (N_5954,N_5256,N_5359);
and U5955 (N_5955,N_5310,N_5420);
and U5956 (N_5956,N_5321,N_5411);
xor U5957 (N_5957,N_5229,N_5121);
or U5958 (N_5958,N_5350,N_5022);
and U5959 (N_5959,N_5359,N_5453);
nand U5960 (N_5960,N_5489,N_5267);
nor U5961 (N_5961,N_5422,N_5154);
nor U5962 (N_5962,N_5358,N_5287);
nor U5963 (N_5963,N_5137,N_5397);
or U5964 (N_5964,N_5437,N_5150);
and U5965 (N_5965,N_5108,N_5300);
nor U5966 (N_5966,N_5252,N_5162);
nand U5967 (N_5967,N_5034,N_5116);
xor U5968 (N_5968,N_5043,N_5492);
xor U5969 (N_5969,N_5038,N_5486);
and U5970 (N_5970,N_5086,N_5163);
nand U5971 (N_5971,N_5201,N_5145);
or U5972 (N_5972,N_5474,N_5104);
nand U5973 (N_5973,N_5301,N_5180);
nand U5974 (N_5974,N_5450,N_5113);
and U5975 (N_5975,N_5092,N_5175);
nor U5976 (N_5976,N_5136,N_5019);
or U5977 (N_5977,N_5082,N_5452);
nor U5978 (N_5978,N_5139,N_5160);
xor U5979 (N_5979,N_5000,N_5281);
or U5980 (N_5980,N_5370,N_5172);
nand U5981 (N_5981,N_5354,N_5304);
nand U5982 (N_5982,N_5041,N_5083);
and U5983 (N_5983,N_5107,N_5069);
and U5984 (N_5984,N_5428,N_5110);
and U5985 (N_5985,N_5109,N_5013);
xor U5986 (N_5986,N_5499,N_5445);
nor U5987 (N_5987,N_5128,N_5345);
xor U5988 (N_5988,N_5256,N_5192);
and U5989 (N_5989,N_5152,N_5130);
nand U5990 (N_5990,N_5253,N_5399);
nor U5991 (N_5991,N_5344,N_5390);
and U5992 (N_5992,N_5248,N_5039);
and U5993 (N_5993,N_5494,N_5256);
or U5994 (N_5994,N_5071,N_5038);
nand U5995 (N_5995,N_5288,N_5030);
or U5996 (N_5996,N_5386,N_5134);
and U5997 (N_5997,N_5296,N_5136);
and U5998 (N_5998,N_5304,N_5435);
or U5999 (N_5999,N_5014,N_5142);
or U6000 (N_6000,N_5833,N_5721);
xor U6001 (N_6001,N_5914,N_5691);
nor U6002 (N_6002,N_5918,N_5698);
nor U6003 (N_6003,N_5774,N_5553);
and U6004 (N_6004,N_5621,N_5814);
xnor U6005 (N_6005,N_5931,N_5762);
and U6006 (N_6006,N_5637,N_5883);
xnor U6007 (N_6007,N_5937,N_5759);
xnor U6008 (N_6008,N_5878,N_5566);
nand U6009 (N_6009,N_5732,N_5563);
xor U6010 (N_6010,N_5982,N_5990);
or U6011 (N_6011,N_5654,N_5502);
nand U6012 (N_6012,N_5555,N_5934);
nor U6013 (N_6013,N_5796,N_5890);
or U6014 (N_6014,N_5632,N_5564);
or U6015 (N_6015,N_5987,N_5584);
or U6016 (N_6016,N_5751,N_5784);
nand U6017 (N_6017,N_5678,N_5813);
nand U6018 (N_6018,N_5783,N_5744);
nand U6019 (N_6019,N_5792,N_5529);
and U6020 (N_6020,N_5627,N_5623);
nand U6021 (N_6021,N_5945,N_5899);
xor U6022 (N_6022,N_5800,N_5794);
or U6023 (N_6023,N_5970,N_5981);
or U6024 (N_6024,N_5745,N_5993);
and U6025 (N_6025,N_5786,N_5935);
xor U6026 (N_6026,N_5765,N_5595);
nand U6027 (N_6027,N_5709,N_5518);
and U6028 (N_6028,N_5609,N_5825);
xor U6029 (N_6029,N_5941,N_5689);
xor U6030 (N_6030,N_5870,N_5871);
nand U6031 (N_6031,N_5634,N_5548);
and U6032 (N_6032,N_5582,N_5509);
and U6033 (N_6033,N_5718,N_5618);
nand U6034 (N_6034,N_5706,N_5948);
xor U6035 (N_6035,N_5644,N_5638);
xnor U6036 (N_6036,N_5926,N_5873);
and U6037 (N_6037,N_5598,N_5722);
or U6038 (N_6038,N_5554,N_5608);
nand U6039 (N_6039,N_5600,N_5785);
nand U6040 (N_6040,N_5953,N_5967);
and U6041 (N_6041,N_5612,N_5647);
and U6042 (N_6042,N_5975,N_5979);
xnor U6043 (N_6043,N_5697,N_5592);
nand U6044 (N_6044,N_5674,N_5865);
xnor U6045 (N_6045,N_5779,N_5604);
xnor U6046 (N_6046,N_5500,N_5806);
nand U6047 (N_6047,N_5606,N_5530);
xor U6048 (N_6048,N_5940,N_5610);
and U6049 (N_6049,N_5725,N_5620);
and U6050 (N_6050,N_5716,N_5665);
xor U6051 (N_6051,N_5594,N_5547);
xnor U6052 (N_6052,N_5572,N_5950);
xnor U6053 (N_6053,N_5636,N_5943);
xor U6054 (N_6054,N_5843,N_5954);
xor U6055 (N_6055,N_5642,N_5903);
nand U6056 (N_6056,N_5649,N_5817);
nand U6057 (N_6057,N_5687,N_5590);
nand U6058 (N_6058,N_5570,N_5551);
nand U6059 (N_6059,N_5753,N_5655);
and U6060 (N_6060,N_5882,N_5850);
and U6061 (N_6061,N_5910,N_5846);
or U6062 (N_6062,N_5720,N_5963);
nand U6063 (N_6063,N_5780,N_5856);
and U6064 (N_6064,N_5781,N_5991);
nor U6065 (N_6065,N_5675,N_5503);
nor U6066 (N_6066,N_5640,N_5690);
xor U6067 (N_6067,N_5809,N_5888);
and U6068 (N_6068,N_5701,N_5578);
nand U6069 (N_6069,N_5648,N_5695);
xor U6070 (N_6070,N_5580,N_5605);
or U6071 (N_6071,N_5911,N_5629);
and U6072 (N_6072,N_5521,N_5558);
or U6073 (N_6073,N_5810,N_5556);
or U6074 (N_6074,N_5520,N_5879);
xnor U6075 (N_6075,N_5599,N_5836);
xor U6076 (N_6076,N_5686,N_5524);
xnor U6077 (N_6077,N_5681,N_5896);
and U6078 (N_6078,N_5908,N_5626);
xnor U6079 (N_6079,N_5992,N_5522);
or U6080 (N_6080,N_5557,N_5874);
nor U6081 (N_6081,N_5651,N_5912);
or U6082 (N_6082,N_5624,N_5545);
or U6083 (N_6083,N_5876,N_5951);
and U6084 (N_6084,N_5907,N_5985);
or U6085 (N_6085,N_5579,N_5597);
nand U6086 (N_6086,N_5776,N_5507);
nand U6087 (N_6087,N_5510,N_5740);
and U6088 (N_6088,N_5864,N_5639);
nand U6089 (N_6089,N_5615,N_5826);
or U6090 (N_6090,N_5897,N_5552);
xor U6091 (N_6091,N_5757,N_5965);
xnor U6092 (N_6092,N_5508,N_5657);
nor U6093 (N_6093,N_5544,N_5733);
xnor U6094 (N_6094,N_5787,N_5671);
nand U6095 (N_6095,N_5891,N_5688);
nor U6096 (N_6096,N_5962,N_5708);
nand U6097 (N_6097,N_5616,N_5887);
and U6098 (N_6098,N_5677,N_5822);
nor U6099 (N_6099,N_5568,N_5669);
xnor U6100 (N_6100,N_5512,N_5724);
or U6101 (N_6101,N_5501,N_5866);
or U6102 (N_6102,N_5834,N_5946);
or U6103 (N_6103,N_5760,N_5643);
and U6104 (N_6104,N_5575,N_5535);
or U6105 (N_6105,N_5995,N_5567);
nand U6106 (N_6106,N_5761,N_5904);
and U6107 (N_6107,N_5944,N_5603);
xnor U6108 (N_6108,N_5875,N_5956);
or U6109 (N_6109,N_5952,N_5569);
or U6110 (N_6110,N_5924,N_5628);
and U6111 (N_6111,N_5881,N_5829);
xnor U6112 (N_6112,N_5898,N_5742);
and U6113 (N_6113,N_5949,N_5998);
and U6114 (N_6114,N_5617,N_5583);
nand U6115 (N_6115,N_5892,N_5772);
and U6116 (N_6116,N_5619,N_5702);
nand U6117 (N_6117,N_5939,N_5607);
and U6118 (N_6118,N_5596,N_5523);
and U6119 (N_6119,N_5798,N_5775);
xnor U6120 (N_6120,N_5917,N_5923);
and U6121 (N_6121,N_5727,N_5506);
nor U6122 (N_6122,N_5820,N_5828);
xor U6123 (N_6123,N_5532,N_5816);
xor U6124 (N_6124,N_5700,N_5710);
xor U6125 (N_6125,N_5679,N_5539);
or U6126 (N_6126,N_5673,N_5812);
nor U6127 (N_6127,N_5738,N_5755);
nor U6128 (N_6128,N_5540,N_5515);
xor U6129 (N_6129,N_5747,N_5593);
and U6130 (N_6130,N_5758,N_5703);
and U6131 (N_6131,N_5505,N_5957);
nor U6132 (N_6132,N_5659,N_5611);
and U6133 (N_6133,N_5531,N_5750);
and U6134 (N_6134,N_5735,N_5748);
and U6135 (N_6135,N_5831,N_5805);
or U6136 (N_6136,N_5662,N_5823);
nor U6137 (N_6137,N_5516,N_5771);
nor U6138 (N_6138,N_5633,N_5630);
nand U6139 (N_6139,N_5656,N_5801);
and U6140 (N_6140,N_5857,N_5546);
or U6141 (N_6141,N_5631,N_5999);
and U6142 (N_6142,N_5601,N_5676);
or U6143 (N_6143,N_5901,N_5730);
nand U6144 (N_6144,N_5538,N_5811);
nand U6145 (N_6145,N_5562,N_5561);
and U6146 (N_6146,N_5707,N_5723);
or U6147 (N_6147,N_5932,N_5928);
or U6148 (N_6148,N_5622,N_5537);
or U6149 (N_6149,N_5880,N_5713);
and U6150 (N_6150,N_5541,N_5574);
xor U6151 (N_6151,N_5858,N_5737);
xnor U6152 (N_6152,N_5902,N_5915);
or U6153 (N_6153,N_5715,N_5922);
xnor U6154 (N_6154,N_5602,N_5684);
xor U6155 (N_6155,N_5646,N_5877);
or U6156 (N_6156,N_5872,N_5667);
nor U6157 (N_6157,N_5534,N_5849);
nor U6158 (N_6158,N_5799,N_5625);
nor U6159 (N_6159,N_5573,N_5756);
xnor U6160 (N_6160,N_5894,N_5986);
or U6161 (N_6161,N_5900,N_5519);
xnor U6162 (N_6162,N_5851,N_5696);
nand U6163 (N_6163,N_5788,N_5886);
nand U6164 (N_6164,N_5895,N_5841);
xnor U6165 (N_6165,N_5978,N_5885);
xor U6166 (N_6166,N_5514,N_5925);
and U6167 (N_6167,N_5893,N_5905);
nand U6168 (N_6168,N_5955,N_5581);
and U6169 (N_6169,N_5842,N_5848);
nor U6170 (N_6170,N_5921,N_5614);
xnor U6171 (N_6171,N_5980,N_5704);
and U6172 (N_6172,N_5752,N_5726);
and U6173 (N_6173,N_5773,N_5528);
nand U6174 (N_6174,N_5571,N_5728);
nor U6175 (N_6175,N_5741,N_5853);
nand U6176 (N_6176,N_5746,N_5861);
nand U6177 (N_6177,N_5793,N_5961);
nor U6178 (N_6178,N_5658,N_5652);
nand U6179 (N_6179,N_5835,N_5818);
xor U6180 (N_6180,N_5807,N_5795);
nor U6181 (N_6181,N_5588,N_5560);
and U6182 (N_6182,N_5804,N_5743);
xnor U6183 (N_6183,N_5971,N_5692);
nor U6184 (N_6184,N_5803,N_5739);
and U6185 (N_6185,N_5790,N_5916);
nand U6186 (N_6186,N_5536,N_5769);
or U6187 (N_6187,N_5821,N_5717);
and U6188 (N_6188,N_5832,N_5827);
nand U6189 (N_6189,N_5854,N_5670);
nand U6190 (N_6190,N_5712,N_5942);
xnor U6191 (N_6191,N_5525,N_5960);
or U6192 (N_6192,N_5973,N_5550);
and U6193 (N_6193,N_5984,N_5641);
nor U6194 (N_6194,N_5837,N_5542);
and U6195 (N_6195,N_5683,N_5653);
nor U6196 (N_6196,N_5966,N_5969);
and U6197 (N_6197,N_5768,N_5947);
xnor U6198 (N_6198,N_5889,N_5736);
and U6199 (N_6199,N_5577,N_5513);
nand U6200 (N_6200,N_5770,N_5936);
or U6201 (N_6201,N_5789,N_5693);
nor U6202 (N_6202,N_5974,N_5906);
nand U6203 (N_6203,N_5933,N_5958);
and U6204 (N_6204,N_5983,N_5996);
nor U6205 (N_6205,N_5972,N_5685);
xnor U6206 (N_6206,N_5526,N_5533);
and U6207 (N_6207,N_5797,N_5791);
and U6208 (N_6208,N_5543,N_5587);
nand U6209 (N_6209,N_5668,N_5977);
or U6210 (N_6210,N_5860,N_5719);
xor U6211 (N_6211,N_5591,N_5782);
nand U6212 (N_6212,N_5613,N_5929);
nand U6213 (N_6213,N_5680,N_5920);
nand U6214 (N_6214,N_5824,N_5855);
and U6215 (N_6215,N_5650,N_5714);
or U6216 (N_6216,N_5863,N_5549);
xor U6217 (N_6217,N_5839,N_5682);
nor U6218 (N_6218,N_5576,N_5734);
xor U6219 (N_6219,N_5959,N_5527);
or U6220 (N_6220,N_5927,N_5729);
and U6221 (N_6221,N_5847,N_5504);
and U6222 (N_6222,N_5666,N_5994);
xnor U6223 (N_6223,N_5808,N_5661);
and U6224 (N_6224,N_5845,N_5919);
nand U6225 (N_6225,N_5913,N_5589);
nor U6226 (N_6226,N_5645,N_5664);
nand U6227 (N_6227,N_5859,N_5672);
nor U6228 (N_6228,N_5711,N_5767);
or U6229 (N_6229,N_5517,N_5586);
xnor U6230 (N_6230,N_5862,N_5559);
or U6231 (N_6231,N_5699,N_5989);
nor U6232 (N_6232,N_5635,N_5868);
or U6233 (N_6233,N_5660,N_5511);
nor U6234 (N_6234,N_5778,N_5694);
and U6235 (N_6235,N_5815,N_5867);
nor U6236 (N_6236,N_5777,N_5964);
nor U6237 (N_6237,N_5968,N_5705);
or U6238 (N_6238,N_5997,N_5585);
xnor U6239 (N_6239,N_5754,N_5766);
xnor U6240 (N_6240,N_5764,N_5884);
nand U6241 (N_6241,N_5763,N_5930);
xnor U6242 (N_6242,N_5749,N_5830);
xor U6243 (N_6243,N_5852,N_5976);
xnor U6244 (N_6244,N_5869,N_5909);
nor U6245 (N_6245,N_5731,N_5838);
xnor U6246 (N_6246,N_5840,N_5938);
nor U6247 (N_6247,N_5844,N_5663);
and U6248 (N_6248,N_5802,N_5565);
and U6249 (N_6249,N_5819,N_5988);
nand U6250 (N_6250,N_5930,N_5990);
nand U6251 (N_6251,N_5639,N_5539);
and U6252 (N_6252,N_5842,N_5574);
nand U6253 (N_6253,N_5922,N_5671);
and U6254 (N_6254,N_5604,N_5581);
nand U6255 (N_6255,N_5938,N_5874);
nor U6256 (N_6256,N_5847,N_5887);
and U6257 (N_6257,N_5908,N_5895);
nand U6258 (N_6258,N_5589,N_5876);
nor U6259 (N_6259,N_5730,N_5915);
xnor U6260 (N_6260,N_5565,N_5567);
or U6261 (N_6261,N_5834,N_5708);
and U6262 (N_6262,N_5749,N_5996);
or U6263 (N_6263,N_5686,N_5715);
or U6264 (N_6264,N_5883,N_5938);
or U6265 (N_6265,N_5826,N_5825);
and U6266 (N_6266,N_5644,N_5796);
nor U6267 (N_6267,N_5546,N_5882);
and U6268 (N_6268,N_5607,N_5517);
nor U6269 (N_6269,N_5874,N_5695);
nand U6270 (N_6270,N_5667,N_5825);
nor U6271 (N_6271,N_5873,N_5507);
nand U6272 (N_6272,N_5964,N_5811);
xnor U6273 (N_6273,N_5738,N_5703);
nor U6274 (N_6274,N_5796,N_5781);
nand U6275 (N_6275,N_5989,N_5870);
and U6276 (N_6276,N_5864,N_5969);
or U6277 (N_6277,N_5902,N_5967);
and U6278 (N_6278,N_5808,N_5576);
or U6279 (N_6279,N_5535,N_5581);
xor U6280 (N_6280,N_5533,N_5692);
nor U6281 (N_6281,N_5842,N_5547);
nor U6282 (N_6282,N_5623,N_5704);
xor U6283 (N_6283,N_5638,N_5895);
xnor U6284 (N_6284,N_5953,N_5973);
xnor U6285 (N_6285,N_5878,N_5689);
xor U6286 (N_6286,N_5973,N_5874);
nand U6287 (N_6287,N_5737,N_5763);
nand U6288 (N_6288,N_5971,N_5749);
xor U6289 (N_6289,N_5602,N_5943);
or U6290 (N_6290,N_5592,N_5947);
xor U6291 (N_6291,N_5843,N_5728);
or U6292 (N_6292,N_5970,N_5772);
xnor U6293 (N_6293,N_5788,N_5836);
nand U6294 (N_6294,N_5775,N_5611);
or U6295 (N_6295,N_5968,N_5848);
xor U6296 (N_6296,N_5685,N_5862);
nand U6297 (N_6297,N_5838,N_5645);
or U6298 (N_6298,N_5539,N_5833);
nor U6299 (N_6299,N_5784,N_5706);
xor U6300 (N_6300,N_5990,N_5952);
or U6301 (N_6301,N_5760,N_5572);
nand U6302 (N_6302,N_5916,N_5918);
xnor U6303 (N_6303,N_5941,N_5678);
or U6304 (N_6304,N_5505,N_5983);
nor U6305 (N_6305,N_5693,N_5610);
and U6306 (N_6306,N_5758,N_5981);
or U6307 (N_6307,N_5914,N_5539);
and U6308 (N_6308,N_5922,N_5551);
nand U6309 (N_6309,N_5817,N_5805);
xor U6310 (N_6310,N_5542,N_5999);
nor U6311 (N_6311,N_5564,N_5710);
or U6312 (N_6312,N_5782,N_5659);
or U6313 (N_6313,N_5834,N_5607);
or U6314 (N_6314,N_5599,N_5895);
or U6315 (N_6315,N_5736,N_5651);
xor U6316 (N_6316,N_5726,N_5723);
xor U6317 (N_6317,N_5836,N_5964);
and U6318 (N_6318,N_5547,N_5670);
xnor U6319 (N_6319,N_5925,N_5886);
and U6320 (N_6320,N_5588,N_5585);
or U6321 (N_6321,N_5505,N_5930);
nor U6322 (N_6322,N_5690,N_5554);
or U6323 (N_6323,N_5904,N_5541);
xor U6324 (N_6324,N_5615,N_5857);
nor U6325 (N_6325,N_5903,N_5697);
nand U6326 (N_6326,N_5618,N_5972);
or U6327 (N_6327,N_5957,N_5711);
and U6328 (N_6328,N_5668,N_5681);
and U6329 (N_6329,N_5745,N_5672);
and U6330 (N_6330,N_5640,N_5968);
nor U6331 (N_6331,N_5645,N_5659);
xor U6332 (N_6332,N_5627,N_5720);
or U6333 (N_6333,N_5987,N_5960);
xnor U6334 (N_6334,N_5957,N_5941);
or U6335 (N_6335,N_5549,N_5713);
and U6336 (N_6336,N_5780,N_5692);
xnor U6337 (N_6337,N_5822,N_5552);
xor U6338 (N_6338,N_5784,N_5587);
and U6339 (N_6339,N_5797,N_5937);
nand U6340 (N_6340,N_5580,N_5999);
and U6341 (N_6341,N_5762,N_5896);
nand U6342 (N_6342,N_5895,N_5965);
or U6343 (N_6343,N_5873,N_5701);
and U6344 (N_6344,N_5635,N_5567);
or U6345 (N_6345,N_5888,N_5784);
nor U6346 (N_6346,N_5967,N_5543);
nor U6347 (N_6347,N_5500,N_5879);
and U6348 (N_6348,N_5535,N_5985);
or U6349 (N_6349,N_5764,N_5678);
and U6350 (N_6350,N_5948,N_5635);
xnor U6351 (N_6351,N_5738,N_5829);
and U6352 (N_6352,N_5642,N_5708);
or U6353 (N_6353,N_5627,N_5574);
and U6354 (N_6354,N_5517,N_5674);
or U6355 (N_6355,N_5917,N_5903);
xor U6356 (N_6356,N_5856,N_5980);
nor U6357 (N_6357,N_5611,N_5925);
or U6358 (N_6358,N_5688,N_5780);
xor U6359 (N_6359,N_5835,N_5644);
nand U6360 (N_6360,N_5758,N_5551);
and U6361 (N_6361,N_5934,N_5881);
xor U6362 (N_6362,N_5652,N_5569);
nor U6363 (N_6363,N_5807,N_5930);
or U6364 (N_6364,N_5508,N_5962);
or U6365 (N_6365,N_5567,N_5983);
or U6366 (N_6366,N_5618,N_5877);
nand U6367 (N_6367,N_5738,N_5677);
nand U6368 (N_6368,N_5933,N_5997);
nor U6369 (N_6369,N_5691,N_5886);
nor U6370 (N_6370,N_5581,N_5653);
nand U6371 (N_6371,N_5639,N_5595);
xnor U6372 (N_6372,N_5510,N_5848);
or U6373 (N_6373,N_5513,N_5602);
or U6374 (N_6374,N_5972,N_5559);
nand U6375 (N_6375,N_5901,N_5661);
xnor U6376 (N_6376,N_5782,N_5975);
and U6377 (N_6377,N_5637,N_5777);
nor U6378 (N_6378,N_5732,N_5986);
nor U6379 (N_6379,N_5750,N_5752);
nand U6380 (N_6380,N_5708,N_5795);
and U6381 (N_6381,N_5952,N_5615);
nand U6382 (N_6382,N_5808,N_5716);
and U6383 (N_6383,N_5508,N_5546);
and U6384 (N_6384,N_5712,N_5626);
and U6385 (N_6385,N_5836,N_5557);
xor U6386 (N_6386,N_5751,N_5573);
or U6387 (N_6387,N_5850,N_5849);
nor U6388 (N_6388,N_5765,N_5871);
and U6389 (N_6389,N_5556,N_5904);
nor U6390 (N_6390,N_5779,N_5805);
nor U6391 (N_6391,N_5779,N_5749);
nand U6392 (N_6392,N_5625,N_5994);
xnor U6393 (N_6393,N_5831,N_5665);
nor U6394 (N_6394,N_5778,N_5851);
nor U6395 (N_6395,N_5933,N_5914);
or U6396 (N_6396,N_5814,N_5856);
nand U6397 (N_6397,N_5615,N_5738);
xnor U6398 (N_6398,N_5684,N_5937);
nor U6399 (N_6399,N_5883,N_5655);
nand U6400 (N_6400,N_5909,N_5663);
nor U6401 (N_6401,N_5564,N_5761);
and U6402 (N_6402,N_5752,N_5540);
nand U6403 (N_6403,N_5701,N_5697);
or U6404 (N_6404,N_5684,N_5849);
nor U6405 (N_6405,N_5903,N_5529);
or U6406 (N_6406,N_5585,N_5798);
or U6407 (N_6407,N_5739,N_5572);
or U6408 (N_6408,N_5717,N_5782);
and U6409 (N_6409,N_5752,N_5890);
or U6410 (N_6410,N_5855,N_5809);
or U6411 (N_6411,N_5743,N_5599);
or U6412 (N_6412,N_5867,N_5671);
nand U6413 (N_6413,N_5978,N_5626);
nand U6414 (N_6414,N_5858,N_5682);
nand U6415 (N_6415,N_5969,N_5580);
and U6416 (N_6416,N_5799,N_5790);
and U6417 (N_6417,N_5739,N_5771);
nand U6418 (N_6418,N_5716,N_5846);
xnor U6419 (N_6419,N_5685,N_5818);
xnor U6420 (N_6420,N_5955,N_5861);
and U6421 (N_6421,N_5994,N_5748);
and U6422 (N_6422,N_5984,N_5964);
nor U6423 (N_6423,N_5776,N_5747);
xnor U6424 (N_6424,N_5804,N_5566);
nor U6425 (N_6425,N_5924,N_5527);
or U6426 (N_6426,N_5798,N_5826);
xnor U6427 (N_6427,N_5556,N_5560);
nand U6428 (N_6428,N_5734,N_5975);
and U6429 (N_6429,N_5667,N_5850);
or U6430 (N_6430,N_5885,N_5976);
nand U6431 (N_6431,N_5502,N_5687);
or U6432 (N_6432,N_5780,N_5744);
or U6433 (N_6433,N_5961,N_5981);
and U6434 (N_6434,N_5748,N_5639);
nand U6435 (N_6435,N_5703,N_5905);
or U6436 (N_6436,N_5887,N_5976);
and U6437 (N_6437,N_5647,N_5635);
xor U6438 (N_6438,N_5646,N_5547);
nor U6439 (N_6439,N_5820,N_5559);
or U6440 (N_6440,N_5606,N_5896);
nor U6441 (N_6441,N_5530,N_5670);
nor U6442 (N_6442,N_5548,N_5740);
nand U6443 (N_6443,N_5994,N_5832);
nor U6444 (N_6444,N_5584,N_5796);
nor U6445 (N_6445,N_5964,N_5669);
or U6446 (N_6446,N_5628,N_5580);
and U6447 (N_6447,N_5896,N_5974);
xnor U6448 (N_6448,N_5772,N_5775);
xor U6449 (N_6449,N_5770,N_5922);
or U6450 (N_6450,N_5973,N_5607);
or U6451 (N_6451,N_5795,N_5877);
nand U6452 (N_6452,N_5718,N_5658);
or U6453 (N_6453,N_5611,N_5774);
nor U6454 (N_6454,N_5551,N_5647);
nand U6455 (N_6455,N_5507,N_5519);
nor U6456 (N_6456,N_5784,N_5599);
and U6457 (N_6457,N_5945,N_5626);
nor U6458 (N_6458,N_5843,N_5523);
or U6459 (N_6459,N_5806,N_5736);
and U6460 (N_6460,N_5919,N_5896);
or U6461 (N_6461,N_5939,N_5876);
and U6462 (N_6462,N_5784,N_5896);
xor U6463 (N_6463,N_5928,N_5533);
and U6464 (N_6464,N_5924,N_5587);
nand U6465 (N_6465,N_5949,N_5907);
nor U6466 (N_6466,N_5600,N_5692);
nor U6467 (N_6467,N_5831,N_5978);
and U6468 (N_6468,N_5605,N_5876);
or U6469 (N_6469,N_5504,N_5598);
and U6470 (N_6470,N_5536,N_5991);
and U6471 (N_6471,N_5777,N_5560);
nor U6472 (N_6472,N_5736,N_5548);
nand U6473 (N_6473,N_5921,N_5728);
or U6474 (N_6474,N_5601,N_5577);
or U6475 (N_6475,N_5884,N_5733);
and U6476 (N_6476,N_5546,N_5784);
nor U6477 (N_6477,N_5681,N_5795);
xor U6478 (N_6478,N_5657,N_5707);
xnor U6479 (N_6479,N_5739,N_5928);
or U6480 (N_6480,N_5920,N_5526);
or U6481 (N_6481,N_5892,N_5519);
or U6482 (N_6482,N_5587,N_5898);
nor U6483 (N_6483,N_5652,N_5620);
xnor U6484 (N_6484,N_5514,N_5699);
nand U6485 (N_6485,N_5633,N_5652);
and U6486 (N_6486,N_5840,N_5614);
nor U6487 (N_6487,N_5872,N_5985);
nor U6488 (N_6488,N_5580,N_5825);
or U6489 (N_6489,N_5507,N_5854);
nor U6490 (N_6490,N_5849,N_5950);
xnor U6491 (N_6491,N_5883,N_5690);
and U6492 (N_6492,N_5723,N_5995);
and U6493 (N_6493,N_5883,N_5617);
and U6494 (N_6494,N_5715,N_5847);
and U6495 (N_6495,N_5534,N_5574);
nor U6496 (N_6496,N_5650,N_5537);
nand U6497 (N_6497,N_5616,N_5635);
nand U6498 (N_6498,N_5806,N_5888);
nor U6499 (N_6499,N_5806,N_5521);
nand U6500 (N_6500,N_6183,N_6044);
and U6501 (N_6501,N_6050,N_6496);
xnor U6502 (N_6502,N_6179,N_6222);
nand U6503 (N_6503,N_6214,N_6078);
and U6504 (N_6504,N_6051,N_6278);
nand U6505 (N_6505,N_6149,N_6389);
and U6506 (N_6506,N_6104,N_6087);
and U6507 (N_6507,N_6211,N_6369);
and U6508 (N_6508,N_6128,N_6441);
nand U6509 (N_6509,N_6386,N_6410);
xor U6510 (N_6510,N_6338,N_6210);
nand U6511 (N_6511,N_6471,N_6446);
xnor U6512 (N_6512,N_6006,N_6216);
nand U6513 (N_6513,N_6094,N_6141);
and U6514 (N_6514,N_6140,N_6480);
xnor U6515 (N_6515,N_6220,N_6405);
nor U6516 (N_6516,N_6106,N_6137);
xnor U6517 (N_6517,N_6492,N_6292);
nor U6518 (N_6518,N_6150,N_6105);
nand U6519 (N_6519,N_6375,N_6270);
and U6520 (N_6520,N_6299,N_6248);
nor U6521 (N_6521,N_6314,N_6444);
xnor U6522 (N_6522,N_6483,N_6181);
or U6523 (N_6523,N_6407,N_6343);
and U6524 (N_6524,N_6316,N_6059);
nor U6525 (N_6525,N_6239,N_6194);
or U6526 (N_6526,N_6182,N_6024);
xor U6527 (N_6527,N_6479,N_6086);
nand U6528 (N_6528,N_6171,N_6250);
xnor U6529 (N_6529,N_6322,N_6038);
or U6530 (N_6530,N_6377,N_6459);
or U6531 (N_6531,N_6302,N_6075);
nand U6532 (N_6532,N_6157,N_6116);
or U6533 (N_6533,N_6247,N_6174);
and U6534 (N_6534,N_6062,N_6258);
nor U6535 (N_6535,N_6445,N_6262);
nor U6536 (N_6536,N_6436,N_6234);
or U6537 (N_6537,N_6039,N_6199);
and U6538 (N_6538,N_6019,N_6259);
xor U6539 (N_6539,N_6148,N_6030);
nor U6540 (N_6540,N_6068,N_6219);
or U6541 (N_6541,N_6365,N_6451);
nand U6542 (N_6542,N_6497,N_6448);
nor U6543 (N_6543,N_6452,N_6387);
xnor U6544 (N_6544,N_6393,N_6423);
nor U6545 (N_6545,N_6133,N_6111);
xor U6546 (N_6546,N_6466,N_6282);
nor U6547 (N_6547,N_6224,N_6486);
and U6548 (N_6548,N_6409,N_6154);
nand U6549 (N_6549,N_6455,N_6072);
or U6550 (N_6550,N_6127,N_6303);
or U6551 (N_6551,N_6095,N_6485);
xnor U6552 (N_6552,N_6090,N_6306);
or U6553 (N_6553,N_6424,N_6240);
nand U6554 (N_6554,N_6065,N_6165);
nand U6555 (N_6555,N_6131,N_6110);
nor U6556 (N_6556,N_6256,N_6053);
and U6557 (N_6557,N_6443,N_6473);
nand U6558 (N_6558,N_6034,N_6162);
or U6559 (N_6559,N_6073,N_6435);
or U6560 (N_6560,N_6012,N_6226);
nor U6561 (N_6561,N_6016,N_6212);
and U6562 (N_6562,N_6061,N_6176);
or U6563 (N_6563,N_6231,N_6469);
nand U6564 (N_6564,N_6070,N_6488);
or U6565 (N_6565,N_6201,N_6396);
or U6566 (N_6566,N_6121,N_6359);
nor U6567 (N_6567,N_6376,N_6287);
nand U6568 (N_6568,N_6045,N_6402);
nand U6569 (N_6569,N_6472,N_6146);
xor U6570 (N_6570,N_6002,N_6232);
nor U6571 (N_6571,N_6193,N_6168);
nand U6572 (N_6572,N_6261,N_6196);
nand U6573 (N_6573,N_6271,N_6124);
and U6574 (N_6574,N_6321,N_6029);
nor U6575 (N_6575,N_6081,N_6041);
and U6576 (N_6576,N_6301,N_6099);
xnor U6577 (N_6577,N_6253,N_6429);
nor U6578 (N_6578,N_6427,N_6358);
or U6579 (N_6579,N_6384,N_6371);
or U6580 (N_6580,N_6163,N_6257);
and U6581 (N_6581,N_6112,N_6098);
nand U6582 (N_6582,N_6333,N_6060);
xor U6583 (N_6583,N_6113,N_6103);
nand U6584 (N_6584,N_6122,N_6372);
xnor U6585 (N_6585,N_6380,N_6033);
xnor U6586 (N_6586,N_6138,N_6277);
nor U6587 (N_6587,N_6330,N_6318);
and U6588 (N_6588,N_6374,N_6312);
nand U6589 (N_6589,N_6433,N_6323);
or U6590 (N_6590,N_6067,N_6191);
nor U6591 (N_6591,N_6209,N_6093);
xnor U6592 (N_6592,N_6144,N_6342);
xnor U6593 (N_6593,N_6079,N_6378);
or U6594 (N_6594,N_6197,N_6421);
nand U6595 (N_6595,N_6326,N_6390);
xor U6596 (N_6596,N_6289,N_6419);
or U6597 (N_6597,N_6047,N_6015);
or U6598 (N_6598,N_6428,N_6238);
nand U6599 (N_6599,N_6468,N_6017);
nor U6600 (N_6600,N_6458,N_6170);
nand U6601 (N_6601,N_6102,N_6158);
nor U6602 (N_6602,N_6223,N_6225);
nand U6603 (N_6603,N_6130,N_6349);
nor U6604 (N_6604,N_6005,N_6252);
nor U6605 (N_6605,N_6432,N_6217);
xor U6606 (N_6606,N_6273,N_6023);
nand U6607 (N_6607,N_6331,N_6119);
nor U6608 (N_6608,N_6063,N_6208);
and U6609 (N_6609,N_6412,N_6481);
nand U6610 (N_6610,N_6195,N_6007);
or U6611 (N_6611,N_6042,N_6276);
or U6612 (N_6612,N_6319,N_6032);
nor U6613 (N_6613,N_6244,N_6484);
or U6614 (N_6614,N_6324,N_6001);
nor U6615 (N_6615,N_6453,N_6340);
nand U6616 (N_6616,N_6354,N_6398);
and U6617 (N_6617,N_6494,N_6064);
nand U6618 (N_6618,N_6279,N_6037);
xor U6619 (N_6619,N_6177,N_6052);
or U6620 (N_6620,N_6311,N_6403);
nor U6621 (N_6621,N_6228,N_6281);
and U6622 (N_6622,N_6080,N_6255);
or U6623 (N_6623,N_6266,N_6101);
and U6624 (N_6624,N_6397,N_6304);
xnor U6625 (N_6625,N_6313,N_6077);
nor U6626 (N_6626,N_6031,N_6198);
nor U6627 (N_6627,N_6339,N_6348);
xnor U6628 (N_6628,N_6309,N_6392);
nor U6629 (N_6629,N_6178,N_6352);
and U6630 (N_6630,N_6013,N_6009);
and U6631 (N_6631,N_6260,N_6167);
nor U6632 (N_6632,N_6329,N_6213);
nor U6633 (N_6633,N_6000,N_6344);
xnor U6634 (N_6634,N_6418,N_6003);
or U6635 (N_6635,N_6251,N_6347);
nand U6636 (N_6636,N_6118,N_6020);
xor U6637 (N_6637,N_6120,N_6074);
nor U6638 (N_6638,N_6026,N_6477);
nor U6639 (N_6639,N_6430,N_6341);
nor U6640 (N_6640,N_6391,N_6125);
nor U6641 (N_6641,N_6159,N_6114);
nor U6642 (N_6642,N_6334,N_6490);
xnor U6643 (N_6643,N_6230,N_6058);
nand U6644 (N_6644,N_6487,N_6462);
or U6645 (N_6645,N_6464,N_6164);
and U6646 (N_6646,N_6385,N_6237);
and U6647 (N_6647,N_6294,N_6283);
nand U6648 (N_6648,N_6373,N_6189);
or U6649 (N_6649,N_6284,N_6350);
nor U6650 (N_6650,N_6335,N_6272);
xor U6651 (N_6651,N_6014,N_6117);
xnor U6652 (N_6652,N_6227,N_6035);
and U6653 (N_6653,N_6202,N_6285);
nand U6654 (N_6654,N_6361,N_6245);
nor U6655 (N_6655,N_6265,N_6450);
nand U6656 (N_6656,N_6221,N_6143);
or U6657 (N_6657,N_6246,N_6040);
nand U6658 (N_6658,N_6097,N_6442);
nand U6659 (N_6659,N_6091,N_6153);
nor U6660 (N_6660,N_6475,N_6243);
xnor U6661 (N_6661,N_6152,N_6394);
or U6662 (N_6662,N_6315,N_6470);
nand U6663 (N_6663,N_6379,N_6155);
nor U6664 (N_6664,N_6115,N_6425);
and U6665 (N_6665,N_6305,N_6493);
xnor U6666 (N_6666,N_6242,N_6132);
xnor U6667 (N_6667,N_6204,N_6401);
or U6668 (N_6668,N_6346,N_6463);
and U6669 (N_6669,N_6076,N_6188);
and U6670 (N_6670,N_6293,N_6416);
and U6671 (N_6671,N_6461,N_6046);
or U6672 (N_6672,N_6018,N_6085);
xnor U6673 (N_6673,N_6071,N_6139);
and U6674 (N_6674,N_6404,N_6364);
nand U6675 (N_6675,N_6160,N_6362);
nand U6676 (N_6676,N_6215,N_6190);
and U6677 (N_6677,N_6172,N_6439);
xnor U6678 (N_6678,N_6192,N_6021);
xor U6679 (N_6679,N_6382,N_6022);
and U6680 (N_6680,N_6482,N_6298);
xor U6681 (N_6681,N_6291,N_6355);
and U6682 (N_6682,N_6109,N_6100);
and U6683 (N_6683,N_6082,N_6426);
xnor U6684 (N_6684,N_6366,N_6142);
or U6685 (N_6685,N_6084,N_6413);
or U6686 (N_6686,N_6048,N_6328);
or U6687 (N_6687,N_6028,N_6356);
nand U6688 (N_6688,N_6325,N_6107);
or U6689 (N_6689,N_6476,N_6057);
and U6690 (N_6690,N_6205,N_6357);
nor U6691 (N_6691,N_6096,N_6367);
xnor U6692 (N_6692,N_6495,N_6145);
or U6693 (N_6693,N_6186,N_6417);
or U6694 (N_6694,N_6456,N_6310);
xnor U6695 (N_6695,N_6307,N_6011);
or U6696 (N_6696,N_6200,N_6414);
xnor U6697 (N_6697,N_6184,N_6054);
nand U6698 (N_6698,N_6489,N_6056);
or U6699 (N_6699,N_6411,N_6465);
or U6700 (N_6700,N_6088,N_6268);
nor U6701 (N_6701,N_6108,N_6351);
and U6702 (N_6702,N_6336,N_6235);
or U6703 (N_6703,N_6136,N_6254);
xor U6704 (N_6704,N_6241,N_6434);
nor U6705 (N_6705,N_6089,N_6449);
nor U6706 (N_6706,N_6457,N_6129);
nor U6707 (N_6707,N_6010,N_6236);
or U6708 (N_6708,N_6498,N_6092);
or U6709 (N_6709,N_6368,N_6437);
nor U6710 (N_6710,N_6274,N_6438);
or U6711 (N_6711,N_6297,N_6055);
nor U6712 (N_6712,N_6218,N_6267);
or U6713 (N_6713,N_6083,N_6151);
and U6714 (N_6714,N_6460,N_6169);
nor U6715 (N_6715,N_6135,N_6175);
and U6716 (N_6716,N_6156,N_6173);
and U6717 (N_6717,N_6406,N_6049);
nor U6718 (N_6718,N_6290,N_6286);
and U6719 (N_6719,N_6295,N_6499);
and U6720 (N_6720,N_6317,N_6415);
nand U6721 (N_6721,N_6491,N_6206);
nor U6722 (N_6722,N_6381,N_6370);
nor U6723 (N_6723,N_6025,N_6467);
nor U6724 (N_6724,N_6383,N_6280);
nor U6725 (N_6725,N_6440,N_6422);
nor U6726 (N_6726,N_6263,N_6275);
xnor U6727 (N_6727,N_6147,N_6043);
or U6728 (N_6728,N_6269,N_6069);
xnor U6729 (N_6729,N_6288,N_6388);
nor U6730 (N_6730,N_6134,N_6345);
nor U6731 (N_6731,N_6431,N_6264);
and U6732 (N_6732,N_6420,N_6180);
and U6733 (N_6733,N_6008,N_6185);
xor U6734 (N_6734,N_6123,N_6187);
or U6735 (N_6735,N_6400,N_6399);
and U6736 (N_6736,N_6004,N_6036);
xor U6737 (N_6737,N_6327,N_6332);
and U6738 (N_6738,N_6308,N_6360);
and U6739 (N_6739,N_6161,N_6027);
xor U6740 (N_6740,N_6203,N_6296);
or U6741 (N_6741,N_6300,N_6126);
or U6742 (N_6742,N_6395,N_6066);
or U6743 (N_6743,N_6363,N_6166);
nand U6744 (N_6744,N_6337,N_6454);
nor U6745 (N_6745,N_6478,N_6474);
nand U6746 (N_6746,N_6249,N_6233);
xor U6747 (N_6747,N_6447,N_6229);
or U6748 (N_6748,N_6320,N_6207);
nor U6749 (N_6749,N_6353,N_6408);
nand U6750 (N_6750,N_6391,N_6471);
and U6751 (N_6751,N_6051,N_6219);
or U6752 (N_6752,N_6259,N_6059);
and U6753 (N_6753,N_6481,N_6032);
xnor U6754 (N_6754,N_6316,N_6260);
and U6755 (N_6755,N_6151,N_6338);
nor U6756 (N_6756,N_6060,N_6033);
and U6757 (N_6757,N_6372,N_6272);
or U6758 (N_6758,N_6456,N_6010);
nor U6759 (N_6759,N_6367,N_6036);
nand U6760 (N_6760,N_6418,N_6360);
or U6761 (N_6761,N_6297,N_6044);
xnor U6762 (N_6762,N_6282,N_6420);
nor U6763 (N_6763,N_6009,N_6029);
and U6764 (N_6764,N_6332,N_6416);
or U6765 (N_6765,N_6268,N_6105);
nand U6766 (N_6766,N_6258,N_6429);
nor U6767 (N_6767,N_6301,N_6456);
nand U6768 (N_6768,N_6301,N_6298);
nand U6769 (N_6769,N_6048,N_6322);
xor U6770 (N_6770,N_6018,N_6154);
nand U6771 (N_6771,N_6026,N_6272);
or U6772 (N_6772,N_6486,N_6079);
nor U6773 (N_6773,N_6007,N_6314);
and U6774 (N_6774,N_6388,N_6344);
nand U6775 (N_6775,N_6276,N_6084);
nand U6776 (N_6776,N_6136,N_6429);
nand U6777 (N_6777,N_6485,N_6104);
and U6778 (N_6778,N_6346,N_6317);
or U6779 (N_6779,N_6378,N_6383);
xor U6780 (N_6780,N_6439,N_6093);
nand U6781 (N_6781,N_6383,N_6490);
and U6782 (N_6782,N_6298,N_6280);
nand U6783 (N_6783,N_6074,N_6189);
or U6784 (N_6784,N_6093,N_6420);
or U6785 (N_6785,N_6050,N_6387);
xnor U6786 (N_6786,N_6255,N_6485);
and U6787 (N_6787,N_6313,N_6070);
and U6788 (N_6788,N_6050,N_6427);
nand U6789 (N_6789,N_6028,N_6349);
xor U6790 (N_6790,N_6074,N_6222);
and U6791 (N_6791,N_6074,N_6028);
xor U6792 (N_6792,N_6302,N_6284);
and U6793 (N_6793,N_6386,N_6091);
and U6794 (N_6794,N_6377,N_6111);
and U6795 (N_6795,N_6261,N_6029);
nor U6796 (N_6796,N_6389,N_6025);
xnor U6797 (N_6797,N_6453,N_6401);
or U6798 (N_6798,N_6058,N_6379);
nand U6799 (N_6799,N_6410,N_6210);
and U6800 (N_6800,N_6319,N_6270);
and U6801 (N_6801,N_6219,N_6205);
or U6802 (N_6802,N_6049,N_6373);
and U6803 (N_6803,N_6162,N_6168);
nand U6804 (N_6804,N_6478,N_6117);
xnor U6805 (N_6805,N_6406,N_6465);
or U6806 (N_6806,N_6258,N_6106);
or U6807 (N_6807,N_6127,N_6273);
or U6808 (N_6808,N_6133,N_6448);
or U6809 (N_6809,N_6237,N_6280);
xnor U6810 (N_6810,N_6350,N_6052);
xnor U6811 (N_6811,N_6333,N_6444);
and U6812 (N_6812,N_6483,N_6137);
nand U6813 (N_6813,N_6465,N_6152);
and U6814 (N_6814,N_6030,N_6168);
nor U6815 (N_6815,N_6401,N_6254);
xnor U6816 (N_6816,N_6186,N_6129);
nor U6817 (N_6817,N_6112,N_6316);
nand U6818 (N_6818,N_6219,N_6163);
or U6819 (N_6819,N_6496,N_6484);
xnor U6820 (N_6820,N_6111,N_6436);
and U6821 (N_6821,N_6121,N_6497);
or U6822 (N_6822,N_6458,N_6311);
and U6823 (N_6823,N_6143,N_6385);
and U6824 (N_6824,N_6287,N_6464);
nand U6825 (N_6825,N_6352,N_6205);
nor U6826 (N_6826,N_6011,N_6368);
xor U6827 (N_6827,N_6437,N_6180);
and U6828 (N_6828,N_6470,N_6466);
nor U6829 (N_6829,N_6048,N_6470);
nor U6830 (N_6830,N_6474,N_6029);
and U6831 (N_6831,N_6207,N_6097);
or U6832 (N_6832,N_6018,N_6299);
or U6833 (N_6833,N_6088,N_6296);
and U6834 (N_6834,N_6462,N_6171);
nor U6835 (N_6835,N_6338,N_6426);
nor U6836 (N_6836,N_6299,N_6439);
and U6837 (N_6837,N_6208,N_6410);
nand U6838 (N_6838,N_6046,N_6105);
nor U6839 (N_6839,N_6409,N_6115);
nor U6840 (N_6840,N_6300,N_6384);
xnor U6841 (N_6841,N_6176,N_6022);
xnor U6842 (N_6842,N_6013,N_6361);
nand U6843 (N_6843,N_6309,N_6116);
or U6844 (N_6844,N_6063,N_6367);
xnor U6845 (N_6845,N_6165,N_6018);
xnor U6846 (N_6846,N_6108,N_6222);
xor U6847 (N_6847,N_6067,N_6110);
nand U6848 (N_6848,N_6470,N_6185);
nor U6849 (N_6849,N_6359,N_6279);
and U6850 (N_6850,N_6174,N_6335);
or U6851 (N_6851,N_6242,N_6335);
or U6852 (N_6852,N_6148,N_6380);
nand U6853 (N_6853,N_6289,N_6252);
nand U6854 (N_6854,N_6333,N_6222);
or U6855 (N_6855,N_6283,N_6177);
or U6856 (N_6856,N_6040,N_6043);
xor U6857 (N_6857,N_6227,N_6294);
nor U6858 (N_6858,N_6367,N_6346);
nand U6859 (N_6859,N_6191,N_6477);
nor U6860 (N_6860,N_6195,N_6362);
or U6861 (N_6861,N_6181,N_6137);
and U6862 (N_6862,N_6271,N_6483);
or U6863 (N_6863,N_6158,N_6355);
nor U6864 (N_6864,N_6029,N_6319);
nor U6865 (N_6865,N_6154,N_6462);
xor U6866 (N_6866,N_6144,N_6217);
nor U6867 (N_6867,N_6299,N_6285);
nand U6868 (N_6868,N_6268,N_6336);
nand U6869 (N_6869,N_6023,N_6220);
and U6870 (N_6870,N_6057,N_6403);
and U6871 (N_6871,N_6002,N_6399);
nand U6872 (N_6872,N_6029,N_6121);
or U6873 (N_6873,N_6291,N_6401);
xnor U6874 (N_6874,N_6190,N_6129);
nor U6875 (N_6875,N_6374,N_6079);
or U6876 (N_6876,N_6084,N_6201);
or U6877 (N_6877,N_6106,N_6490);
nor U6878 (N_6878,N_6195,N_6457);
and U6879 (N_6879,N_6351,N_6015);
xnor U6880 (N_6880,N_6457,N_6413);
nand U6881 (N_6881,N_6318,N_6354);
and U6882 (N_6882,N_6196,N_6185);
and U6883 (N_6883,N_6362,N_6458);
nor U6884 (N_6884,N_6250,N_6188);
nand U6885 (N_6885,N_6111,N_6052);
nor U6886 (N_6886,N_6065,N_6044);
and U6887 (N_6887,N_6376,N_6226);
or U6888 (N_6888,N_6346,N_6157);
nand U6889 (N_6889,N_6436,N_6488);
nand U6890 (N_6890,N_6347,N_6128);
nand U6891 (N_6891,N_6008,N_6454);
or U6892 (N_6892,N_6284,N_6062);
and U6893 (N_6893,N_6486,N_6356);
xnor U6894 (N_6894,N_6305,N_6490);
and U6895 (N_6895,N_6178,N_6133);
xor U6896 (N_6896,N_6392,N_6454);
nor U6897 (N_6897,N_6061,N_6358);
nand U6898 (N_6898,N_6327,N_6095);
nand U6899 (N_6899,N_6112,N_6296);
and U6900 (N_6900,N_6362,N_6034);
nand U6901 (N_6901,N_6007,N_6149);
and U6902 (N_6902,N_6134,N_6460);
and U6903 (N_6903,N_6149,N_6101);
xnor U6904 (N_6904,N_6336,N_6209);
nor U6905 (N_6905,N_6298,N_6074);
xor U6906 (N_6906,N_6363,N_6468);
nor U6907 (N_6907,N_6050,N_6280);
nand U6908 (N_6908,N_6175,N_6090);
nor U6909 (N_6909,N_6064,N_6047);
or U6910 (N_6910,N_6479,N_6048);
xor U6911 (N_6911,N_6396,N_6161);
or U6912 (N_6912,N_6050,N_6362);
nand U6913 (N_6913,N_6364,N_6245);
xor U6914 (N_6914,N_6050,N_6000);
nor U6915 (N_6915,N_6333,N_6495);
xnor U6916 (N_6916,N_6073,N_6385);
nand U6917 (N_6917,N_6210,N_6200);
or U6918 (N_6918,N_6405,N_6011);
and U6919 (N_6919,N_6012,N_6319);
xor U6920 (N_6920,N_6401,N_6473);
nand U6921 (N_6921,N_6064,N_6256);
or U6922 (N_6922,N_6012,N_6129);
nor U6923 (N_6923,N_6309,N_6161);
xor U6924 (N_6924,N_6227,N_6276);
and U6925 (N_6925,N_6026,N_6120);
xor U6926 (N_6926,N_6068,N_6242);
xor U6927 (N_6927,N_6041,N_6393);
xor U6928 (N_6928,N_6232,N_6287);
nor U6929 (N_6929,N_6310,N_6382);
nand U6930 (N_6930,N_6218,N_6237);
xnor U6931 (N_6931,N_6415,N_6245);
and U6932 (N_6932,N_6219,N_6157);
or U6933 (N_6933,N_6328,N_6049);
xor U6934 (N_6934,N_6249,N_6401);
xnor U6935 (N_6935,N_6084,N_6441);
xor U6936 (N_6936,N_6493,N_6078);
nand U6937 (N_6937,N_6386,N_6218);
and U6938 (N_6938,N_6428,N_6313);
or U6939 (N_6939,N_6469,N_6094);
nand U6940 (N_6940,N_6000,N_6428);
nand U6941 (N_6941,N_6348,N_6085);
xnor U6942 (N_6942,N_6372,N_6352);
nand U6943 (N_6943,N_6380,N_6093);
xnor U6944 (N_6944,N_6094,N_6190);
xnor U6945 (N_6945,N_6143,N_6210);
nor U6946 (N_6946,N_6417,N_6495);
xor U6947 (N_6947,N_6254,N_6413);
nor U6948 (N_6948,N_6427,N_6267);
and U6949 (N_6949,N_6207,N_6315);
nand U6950 (N_6950,N_6101,N_6333);
xnor U6951 (N_6951,N_6421,N_6160);
nand U6952 (N_6952,N_6437,N_6238);
or U6953 (N_6953,N_6215,N_6108);
or U6954 (N_6954,N_6145,N_6119);
and U6955 (N_6955,N_6174,N_6406);
nand U6956 (N_6956,N_6188,N_6105);
xor U6957 (N_6957,N_6296,N_6035);
nand U6958 (N_6958,N_6038,N_6053);
and U6959 (N_6959,N_6292,N_6284);
or U6960 (N_6960,N_6144,N_6275);
and U6961 (N_6961,N_6187,N_6403);
nor U6962 (N_6962,N_6243,N_6111);
nor U6963 (N_6963,N_6064,N_6382);
or U6964 (N_6964,N_6325,N_6401);
xnor U6965 (N_6965,N_6281,N_6285);
or U6966 (N_6966,N_6157,N_6024);
xor U6967 (N_6967,N_6166,N_6158);
nand U6968 (N_6968,N_6364,N_6447);
and U6969 (N_6969,N_6156,N_6263);
nand U6970 (N_6970,N_6317,N_6142);
or U6971 (N_6971,N_6106,N_6342);
xor U6972 (N_6972,N_6027,N_6321);
nor U6973 (N_6973,N_6209,N_6161);
and U6974 (N_6974,N_6262,N_6233);
and U6975 (N_6975,N_6270,N_6088);
nand U6976 (N_6976,N_6208,N_6486);
nor U6977 (N_6977,N_6446,N_6369);
nor U6978 (N_6978,N_6448,N_6477);
or U6979 (N_6979,N_6161,N_6162);
nor U6980 (N_6980,N_6289,N_6259);
or U6981 (N_6981,N_6328,N_6229);
nor U6982 (N_6982,N_6498,N_6257);
nor U6983 (N_6983,N_6043,N_6046);
nor U6984 (N_6984,N_6196,N_6153);
nor U6985 (N_6985,N_6333,N_6483);
nor U6986 (N_6986,N_6297,N_6131);
nor U6987 (N_6987,N_6358,N_6155);
or U6988 (N_6988,N_6347,N_6419);
or U6989 (N_6989,N_6015,N_6290);
nor U6990 (N_6990,N_6463,N_6397);
or U6991 (N_6991,N_6108,N_6179);
or U6992 (N_6992,N_6215,N_6076);
nand U6993 (N_6993,N_6298,N_6178);
xnor U6994 (N_6994,N_6213,N_6342);
xor U6995 (N_6995,N_6144,N_6263);
nand U6996 (N_6996,N_6079,N_6376);
and U6997 (N_6997,N_6160,N_6049);
nor U6998 (N_6998,N_6242,N_6014);
nand U6999 (N_6999,N_6492,N_6283);
or U7000 (N_7000,N_6609,N_6970);
nand U7001 (N_7001,N_6670,N_6753);
or U7002 (N_7002,N_6747,N_6566);
nand U7003 (N_7003,N_6636,N_6667);
or U7004 (N_7004,N_6589,N_6990);
nor U7005 (N_7005,N_6529,N_6762);
nand U7006 (N_7006,N_6552,N_6783);
or U7007 (N_7007,N_6554,N_6645);
xor U7008 (N_7008,N_6941,N_6958);
and U7009 (N_7009,N_6822,N_6683);
and U7010 (N_7010,N_6768,N_6874);
or U7011 (N_7011,N_6885,N_6847);
nand U7012 (N_7012,N_6731,N_6812);
and U7013 (N_7013,N_6980,N_6844);
nand U7014 (N_7014,N_6692,N_6916);
xnor U7015 (N_7015,N_6788,N_6843);
and U7016 (N_7016,N_6543,N_6930);
nor U7017 (N_7017,N_6948,N_6635);
and U7018 (N_7018,N_6903,N_6611);
and U7019 (N_7019,N_6946,N_6549);
xnor U7020 (N_7020,N_6957,N_6520);
nor U7021 (N_7021,N_6926,N_6833);
nor U7022 (N_7022,N_6621,N_6974);
or U7023 (N_7023,N_6514,N_6653);
nor U7024 (N_7024,N_6976,N_6921);
xor U7025 (N_7025,N_6913,N_6672);
or U7026 (N_7026,N_6890,N_6760);
nor U7027 (N_7027,N_6593,N_6709);
nor U7028 (N_7028,N_6513,N_6892);
xor U7029 (N_7029,N_6633,N_6869);
and U7030 (N_7030,N_6713,N_6715);
xor U7031 (N_7031,N_6956,N_6909);
or U7032 (N_7032,N_6527,N_6615);
nor U7033 (N_7033,N_6998,N_6853);
and U7034 (N_7034,N_6984,N_6969);
xor U7035 (N_7035,N_6684,N_6639);
nor U7036 (N_7036,N_6729,N_6938);
and U7037 (N_7037,N_6877,N_6779);
nor U7038 (N_7038,N_6894,N_6603);
or U7039 (N_7039,N_6682,N_6900);
nor U7040 (N_7040,N_6710,N_6735);
nor U7041 (N_7041,N_6761,N_6570);
or U7042 (N_7042,N_6977,N_6604);
or U7043 (N_7043,N_6986,N_6596);
and U7044 (N_7044,N_6581,N_6521);
or U7045 (N_7045,N_6632,N_6919);
or U7046 (N_7046,N_6789,N_6696);
and U7047 (N_7047,N_6988,N_6910);
nor U7048 (N_7048,N_6775,N_6584);
nand U7049 (N_7049,N_6944,N_6524);
and U7050 (N_7050,N_6823,N_6902);
or U7051 (N_7051,N_6719,N_6698);
and U7052 (N_7052,N_6975,N_6810);
or U7053 (N_7053,N_6734,N_6748);
nor U7054 (N_7054,N_6883,N_6935);
or U7055 (N_7055,N_6700,N_6891);
nor U7056 (N_7056,N_6914,N_6758);
nand U7057 (N_7057,N_6863,N_6732);
nor U7058 (N_7058,N_6950,N_6691);
nor U7059 (N_7059,N_6506,N_6716);
and U7060 (N_7060,N_6781,N_6537);
nand U7061 (N_7061,N_6848,N_6817);
nor U7062 (N_7062,N_6959,N_6583);
or U7063 (N_7063,N_6787,N_6996);
and U7064 (N_7064,N_6790,N_6804);
xnor U7065 (N_7065,N_6786,N_6896);
or U7066 (N_7066,N_6556,N_6824);
nand U7067 (N_7067,N_6539,N_6547);
xnor U7068 (N_7068,N_6749,N_6928);
and U7069 (N_7069,N_6982,N_6846);
nor U7070 (N_7070,N_6881,N_6931);
nand U7071 (N_7071,N_6802,N_6852);
nor U7072 (N_7072,N_6867,N_6771);
and U7073 (N_7073,N_6523,N_6736);
xnor U7074 (N_7074,N_6967,N_6569);
nand U7075 (N_7075,N_6945,N_6884);
or U7076 (N_7076,N_6654,N_6655);
nor U7077 (N_7077,N_6859,N_6536);
or U7078 (N_7078,N_6851,N_6507);
or U7079 (N_7079,N_6849,N_6580);
xor U7080 (N_7080,N_6857,N_6837);
or U7081 (N_7081,N_6707,N_6972);
nor U7082 (N_7082,N_6586,N_6668);
xor U7083 (N_7083,N_6567,N_6688);
xor U7084 (N_7084,N_6770,N_6600);
nand U7085 (N_7085,N_6991,N_6803);
nand U7086 (N_7086,N_6755,N_6727);
nor U7087 (N_7087,N_6625,N_6590);
nand U7088 (N_7088,N_6840,N_6829);
nor U7089 (N_7089,N_6582,N_6797);
and U7090 (N_7090,N_6693,N_6622);
and U7091 (N_7091,N_6659,N_6773);
nand U7092 (N_7092,N_6535,N_6985);
nand U7093 (N_7093,N_6557,N_6888);
or U7094 (N_7094,N_6687,N_6597);
nor U7095 (N_7095,N_6951,N_6871);
nor U7096 (N_7096,N_6978,N_6801);
and U7097 (N_7097,N_6784,N_6799);
and U7098 (N_7098,N_6598,N_6875);
or U7099 (N_7099,N_6664,N_6546);
or U7100 (N_7100,N_6726,N_6947);
xor U7101 (N_7101,N_6511,N_6897);
nor U7102 (N_7102,N_6893,N_6872);
nor U7103 (N_7103,N_6793,N_6968);
xor U7104 (N_7104,N_6887,N_6652);
or U7105 (N_7105,N_6518,N_6809);
or U7106 (N_7106,N_6765,N_6669);
or U7107 (N_7107,N_6943,N_6689);
xnor U7108 (N_7108,N_6724,N_6505);
nand U7109 (N_7109,N_6854,N_6515);
xnor U7110 (N_7110,N_6678,N_6530);
or U7111 (N_7111,N_6638,N_6563);
nor U7112 (N_7112,N_6798,N_6745);
xor U7113 (N_7113,N_6973,N_6791);
nor U7114 (N_7114,N_6658,N_6531);
xor U7115 (N_7115,N_6911,N_6647);
and U7116 (N_7116,N_6594,N_6895);
nand U7117 (N_7117,N_6725,N_6800);
nor U7118 (N_7118,N_6516,N_6585);
nand U7119 (N_7119,N_6508,N_6627);
nand U7120 (N_7120,N_6751,N_6929);
nor U7121 (N_7121,N_6856,N_6733);
nor U7122 (N_7122,N_6607,N_6963);
or U7123 (N_7123,N_6741,N_6677);
or U7124 (N_7124,N_6522,N_6836);
nand U7125 (N_7125,N_6721,N_6559);
or U7126 (N_7126,N_6954,N_6631);
nor U7127 (N_7127,N_6780,N_6744);
or U7128 (N_7128,N_6839,N_6966);
xnor U7129 (N_7129,N_6899,N_6663);
and U7130 (N_7130,N_6542,N_6572);
and U7131 (N_7131,N_6702,N_6595);
or U7132 (N_7132,N_6739,N_6772);
nor U7133 (N_7133,N_6993,N_6901);
and U7134 (N_7134,N_6608,N_6861);
xnor U7135 (N_7135,N_6953,N_6905);
or U7136 (N_7136,N_6813,N_6728);
or U7137 (N_7137,N_6917,N_6828);
xor U7138 (N_7138,N_6740,N_6746);
and U7139 (N_7139,N_6971,N_6553);
and U7140 (N_7140,N_6835,N_6961);
and U7141 (N_7141,N_6940,N_6525);
and U7142 (N_7142,N_6936,N_6876);
nor U7143 (N_7143,N_6866,N_6960);
or U7144 (N_7144,N_6679,N_6845);
xnor U7145 (N_7145,N_6767,N_6695);
nand U7146 (N_7146,N_6757,N_6564);
or U7147 (N_7147,N_6685,N_6722);
nor U7148 (N_7148,N_6738,N_6955);
nor U7149 (N_7149,N_6922,N_6540);
or U7150 (N_7150,N_6898,N_6612);
and U7151 (N_7151,N_6640,N_6614);
xnor U7152 (N_7152,N_6561,N_6532);
xor U7153 (N_7153,N_6742,N_6879);
or U7154 (N_7154,N_6643,N_6510);
nand U7155 (N_7155,N_6701,N_6509);
nor U7156 (N_7156,N_6634,N_6648);
nand U7157 (N_7157,N_6816,N_6754);
nor U7158 (N_7158,N_6550,N_6592);
nand U7159 (N_7159,N_6806,N_6785);
nand U7160 (N_7160,N_6656,N_6660);
nor U7161 (N_7161,N_6952,N_6576);
nor U7162 (N_7162,N_6651,N_6807);
or U7163 (N_7163,N_6626,N_6811);
xnor U7164 (N_7164,N_6720,N_6878);
or U7165 (N_7165,N_6964,N_6665);
and U7166 (N_7166,N_6575,N_6934);
and U7167 (N_7167,N_6618,N_6674);
nor U7168 (N_7168,N_6920,N_6662);
or U7169 (N_7169,N_6841,N_6826);
nor U7170 (N_7170,N_6610,N_6711);
and U7171 (N_7171,N_6686,N_6661);
or U7172 (N_7172,N_6602,N_6965);
or U7173 (N_7173,N_6743,N_6574);
or U7174 (N_7174,N_6657,N_6825);
xor U7175 (N_7175,N_6619,N_6578);
nor U7176 (N_7176,N_6766,N_6503);
and U7177 (N_7177,N_6927,N_6551);
xnor U7178 (N_7178,N_6855,N_6699);
and U7179 (N_7179,N_6915,N_6568);
nor U7180 (N_7180,N_6992,N_6796);
and U7181 (N_7181,N_6939,N_6752);
and U7182 (N_7182,N_6962,N_6886);
or U7183 (N_7183,N_6889,N_6868);
xnor U7184 (N_7184,N_6694,N_6932);
and U7185 (N_7185,N_6577,N_6650);
nor U7186 (N_7186,N_6666,N_6778);
and U7187 (N_7187,N_6500,N_6642);
nor U7188 (N_7188,N_6620,N_6723);
and U7189 (N_7189,N_6544,N_6565);
nor U7190 (N_7190,N_6805,N_6533);
nor U7191 (N_7191,N_6641,N_6850);
or U7192 (N_7192,N_6925,N_6912);
nor U7193 (N_7193,N_6907,N_6862);
xnor U7194 (N_7194,N_6571,N_6599);
and U7195 (N_7195,N_6528,N_6808);
nand U7196 (N_7196,N_6923,N_6649);
nor U7197 (N_7197,N_6512,N_6504);
and U7198 (N_7198,N_6794,N_6933);
and U7199 (N_7199,N_6776,N_6541);
and U7200 (N_7200,N_6646,N_6579);
or U7201 (N_7201,N_6750,N_6830);
xor U7202 (N_7202,N_6999,N_6774);
nand U7203 (N_7203,N_6601,N_6995);
nor U7204 (N_7204,N_6832,N_6681);
or U7205 (N_7205,N_6623,N_6777);
xor U7206 (N_7206,N_6827,N_6834);
xnor U7207 (N_7207,N_6587,N_6987);
and U7208 (N_7208,N_6819,N_6795);
xnor U7209 (N_7209,N_6924,N_6842);
or U7210 (N_7210,N_6558,N_6624);
or U7211 (N_7211,N_6949,N_6637);
nand U7212 (N_7212,N_6942,N_6981);
and U7213 (N_7213,N_6821,N_6997);
xnor U7214 (N_7214,N_6555,N_6979);
or U7215 (N_7215,N_6697,N_6573);
xnor U7216 (N_7216,N_6769,N_6838);
or U7217 (N_7217,N_6671,N_6673);
xnor U7218 (N_7218,N_6718,N_6545);
or U7219 (N_7219,N_6613,N_6763);
and U7220 (N_7220,N_6880,N_6534);
nand U7221 (N_7221,N_6918,N_6764);
xor U7222 (N_7222,N_6588,N_6994);
xor U7223 (N_7223,N_6538,N_6882);
and U7224 (N_7224,N_6680,N_6616);
nor U7225 (N_7225,N_6717,N_6782);
and U7226 (N_7226,N_6870,N_6906);
nand U7227 (N_7227,N_6708,N_6937);
xor U7228 (N_7228,N_6703,N_6873);
or U7229 (N_7229,N_6860,N_6864);
or U7230 (N_7230,N_6737,N_6858);
nand U7231 (N_7231,N_6526,N_6831);
and U7232 (N_7232,N_6519,N_6814);
nand U7233 (N_7233,N_6675,N_6548);
nand U7234 (N_7234,N_6676,N_6983);
nor U7235 (N_7235,N_6818,N_6617);
nor U7236 (N_7236,N_6606,N_6706);
or U7237 (N_7237,N_6792,N_6904);
and U7238 (N_7238,N_6501,N_6628);
nand U7239 (N_7239,N_6759,N_6502);
xnor U7240 (N_7240,N_6989,N_6690);
nand U7241 (N_7241,N_6820,N_6704);
xnor U7242 (N_7242,N_6630,N_6517);
and U7243 (N_7243,N_6591,N_6730);
or U7244 (N_7244,N_6644,N_6705);
xor U7245 (N_7245,N_6629,N_6714);
xnor U7246 (N_7246,N_6865,N_6562);
nand U7247 (N_7247,N_6815,N_6605);
nand U7248 (N_7248,N_6560,N_6756);
nor U7249 (N_7249,N_6712,N_6908);
xnor U7250 (N_7250,N_6740,N_6755);
or U7251 (N_7251,N_6683,N_6659);
and U7252 (N_7252,N_6863,N_6730);
or U7253 (N_7253,N_6804,N_6828);
xor U7254 (N_7254,N_6631,N_6550);
nand U7255 (N_7255,N_6688,N_6813);
xor U7256 (N_7256,N_6987,N_6787);
or U7257 (N_7257,N_6607,N_6624);
and U7258 (N_7258,N_6510,N_6640);
xor U7259 (N_7259,N_6940,N_6754);
nand U7260 (N_7260,N_6934,N_6849);
nand U7261 (N_7261,N_6931,N_6525);
nand U7262 (N_7262,N_6859,N_6966);
nor U7263 (N_7263,N_6520,N_6928);
and U7264 (N_7264,N_6510,N_6895);
xnor U7265 (N_7265,N_6662,N_6882);
and U7266 (N_7266,N_6873,N_6698);
and U7267 (N_7267,N_6987,N_6669);
and U7268 (N_7268,N_6733,N_6844);
nand U7269 (N_7269,N_6946,N_6517);
nor U7270 (N_7270,N_6745,N_6985);
nand U7271 (N_7271,N_6765,N_6925);
xor U7272 (N_7272,N_6864,N_6927);
xor U7273 (N_7273,N_6798,N_6512);
nand U7274 (N_7274,N_6945,N_6938);
and U7275 (N_7275,N_6565,N_6506);
nand U7276 (N_7276,N_6930,N_6941);
or U7277 (N_7277,N_6528,N_6500);
and U7278 (N_7278,N_6818,N_6700);
nor U7279 (N_7279,N_6967,N_6811);
nor U7280 (N_7280,N_6966,N_6718);
xor U7281 (N_7281,N_6706,N_6769);
and U7282 (N_7282,N_6864,N_6571);
and U7283 (N_7283,N_6831,N_6638);
or U7284 (N_7284,N_6992,N_6535);
xnor U7285 (N_7285,N_6629,N_6723);
nand U7286 (N_7286,N_6730,N_6712);
nor U7287 (N_7287,N_6886,N_6746);
nand U7288 (N_7288,N_6854,N_6570);
and U7289 (N_7289,N_6816,N_6982);
nor U7290 (N_7290,N_6708,N_6529);
or U7291 (N_7291,N_6936,N_6712);
and U7292 (N_7292,N_6614,N_6563);
nand U7293 (N_7293,N_6591,N_6802);
xor U7294 (N_7294,N_6908,N_6799);
or U7295 (N_7295,N_6535,N_6801);
nand U7296 (N_7296,N_6803,N_6809);
nor U7297 (N_7297,N_6796,N_6798);
nand U7298 (N_7298,N_6768,N_6937);
xor U7299 (N_7299,N_6828,N_6767);
nand U7300 (N_7300,N_6729,N_6863);
nor U7301 (N_7301,N_6913,N_6657);
or U7302 (N_7302,N_6602,N_6661);
or U7303 (N_7303,N_6868,N_6832);
nand U7304 (N_7304,N_6564,N_6531);
nand U7305 (N_7305,N_6822,N_6902);
and U7306 (N_7306,N_6897,N_6592);
nor U7307 (N_7307,N_6724,N_6841);
nand U7308 (N_7308,N_6603,N_6664);
xor U7309 (N_7309,N_6861,N_6739);
nand U7310 (N_7310,N_6955,N_6937);
or U7311 (N_7311,N_6700,N_6702);
xnor U7312 (N_7312,N_6509,N_6775);
xnor U7313 (N_7313,N_6744,N_6953);
and U7314 (N_7314,N_6765,N_6554);
xor U7315 (N_7315,N_6586,N_6581);
xor U7316 (N_7316,N_6574,N_6923);
nor U7317 (N_7317,N_6795,N_6959);
or U7318 (N_7318,N_6642,N_6727);
and U7319 (N_7319,N_6807,N_6869);
nand U7320 (N_7320,N_6745,N_6511);
and U7321 (N_7321,N_6689,N_6744);
nand U7322 (N_7322,N_6956,N_6736);
and U7323 (N_7323,N_6526,N_6953);
nor U7324 (N_7324,N_6717,N_6509);
nor U7325 (N_7325,N_6915,N_6877);
nand U7326 (N_7326,N_6807,N_6933);
nor U7327 (N_7327,N_6891,N_6581);
nor U7328 (N_7328,N_6780,N_6966);
nor U7329 (N_7329,N_6763,N_6975);
and U7330 (N_7330,N_6543,N_6530);
or U7331 (N_7331,N_6807,N_6747);
xnor U7332 (N_7332,N_6760,N_6909);
nand U7333 (N_7333,N_6780,N_6564);
nor U7334 (N_7334,N_6716,N_6919);
and U7335 (N_7335,N_6833,N_6618);
or U7336 (N_7336,N_6607,N_6603);
or U7337 (N_7337,N_6656,N_6614);
or U7338 (N_7338,N_6896,N_6818);
xor U7339 (N_7339,N_6791,N_6655);
nand U7340 (N_7340,N_6564,N_6714);
or U7341 (N_7341,N_6513,N_6937);
nor U7342 (N_7342,N_6822,N_6581);
nor U7343 (N_7343,N_6772,N_6549);
and U7344 (N_7344,N_6994,N_6896);
xor U7345 (N_7345,N_6932,N_6522);
and U7346 (N_7346,N_6833,N_6856);
xnor U7347 (N_7347,N_6501,N_6790);
nor U7348 (N_7348,N_6884,N_6798);
nand U7349 (N_7349,N_6622,N_6906);
nand U7350 (N_7350,N_6913,N_6626);
and U7351 (N_7351,N_6954,N_6515);
or U7352 (N_7352,N_6549,N_6782);
xnor U7353 (N_7353,N_6630,N_6651);
and U7354 (N_7354,N_6884,N_6700);
and U7355 (N_7355,N_6681,N_6842);
nand U7356 (N_7356,N_6501,N_6849);
and U7357 (N_7357,N_6573,N_6676);
and U7358 (N_7358,N_6763,N_6956);
nand U7359 (N_7359,N_6569,N_6829);
nand U7360 (N_7360,N_6807,N_6530);
nor U7361 (N_7361,N_6538,N_6844);
or U7362 (N_7362,N_6879,N_6918);
nand U7363 (N_7363,N_6679,N_6745);
nand U7364 (N_7364,N_6501,N_6649);
nand U7365 (N_7365,N_6693,N_6754);
nor U7366 (N_7366,N_6862,N_6963);
nand U7367 (N_7367,N_6737,N_6579);
xnor U7368 (N_7368,N_6670,N_6605);
or U7369 (N_7369,N_6565,N_6957);
xor U7370 (N_7370,N_6791,N_6803);
nor U7371 (N_7371,N_6867,N_6514);
nand U7372 (N_7372,N_6694,N_6523);
xnor U7373 (N_7373,N_6664,N_6666);
nor U7374 (N_7374,N_6932,N_6588);
nor U7375 (N_7375,N_6928,N_6500);
and U7376 (N_7376,N_6783,N_6949);
nand U7377 (N_7377,N_6701,N_6512);
xnor U7378 (N_7378,N_6705,N_6936);
nor U7379 (N_7379,N_6567,N_6861);
nand U7380 (N_7380,N_6815,N_6544);
or U7381 (N_7381,N_6633,N_6577);
nand U7382 (N_7382,N_6631,N_6763);
nor U7383 (N_7383,N_6909,N_6658);
or U7384 (N_7384,N_6976,N_6864);
or U7385 (N_7385,N_6688,N_6739);
nand U7386 (N_7386,N_6985,N_6962);
nor U7387 (N_7387,N_6980,N_6610);
or U7388 (N_7388,N_6988,N_6547);
or U7389 (N_7389,N_6754,N_6920);
nand U7390 (N_7390,N_6609,N_6558);
xor U7391 (N_7391,N_6946,N_6835);
and U7392 (N_7392,N_6527,N_6656);
and U7393 (N_7393,N_6554,N_6971);
or U7394 (N_7394,N_6625,N_6651);
xor U7395 (N_7395,N_6682,N_6867);
xor U7396 (N_7396,N_6527,N_6719);
nor U7397 (N_7397,N_6719,N_6656);
or U7398 (N_7398,N_6660,N_6686);
nor U7399 (N_7399,N_6603,N_6829);
xnor U7400 (N_7400,N_6974,N_6806);
and U7401 (N_7401,N_6768,N_6781);
and U7402 (N_7402,N_6655,N_6850);
nor U7403 (N_7403,N_6663,N_6505);
and U7404 (N_7404,N_6747,N_6750);
nand U7405 (N_7405,N_6590,N_6912);
xnor U7406 (N_7406,N_6989,N_6922);
nor U7407 (N_7407,N_6838,N_6812);
nand U7408 (N_7408,N_6726,N_6782);
nand U7409 (N_7409,N_6528,N_6854);
nor U7410 (N_7410,N_6563,N_6883);
nor U7411 (N_7411,N_6580,N_6569);
xnor U7412 (N_7412,N_6741,N_6597);
or U7413 (N_7413,N_6647,N_6798);
and U7414 (N_7414,N_6522,N_6627);
nand U7415 (N_7415,N_6605,N_6828);
nor U7416 (N_7416,N_6507,N_6668);
and U7417 (N_7417,N_6595,N_6563);
or U7418 (N_7418,N_6548,N_6682);
and U7419 (N_7419,N_6759,N_6522);
and U7420 (N_7420,N_6745,N_6906);
nor U7421 (N_7421,N_6992,N_6573);
and U7422 (N_7422,N_6599,N_6851);
nand U7423 (N_7423,N_6544,N_6752);
and U7424 (N_7424,N_6571,N_6685);
nand U7425 (N_7425,N_6902,N_6890);
nand U7426 (N_7426,N_6533,N_6665);
or U7427 (N_7427,N_6860,N_6836);
nand U7428 (N_7428,N_6820,N_6909);
nand U7429 (N_7429,N_6980,N_6627);
nand U7430 (N_7430,N_6802,N_6514);
or U7431 (N_7431,N_6913,N_6690);
nor U7432 (N_7432,N_6611,N_6530);
or U7433 (N_7433,N_6920,N_6937);
xnor U7434 (N_7434,N_6967,N_6995);
xnor U7435 (N_7435,N_6508,N_6583);
nand U7436 (N_7436,N_6738,N_6544);
and U7437 (N_7437,N_6505,N_6511);
and U7438 (N_7438,N_6588,N_6933);
nor U7439 (N_7439,N_6990,N_6971);
or U7440 (N_7440,N_6800,N_6959);
or U7441 (N_7441,N_6911,N_6683);
nor U7442 (N_7442,N_6647,N_6531);
nand U7443 (N_7443,N_6933,N_6558);
nand U7444 (N_7444,N_6699,N_6794);
nand U7445 (N_7445,N_6813,N_6504);
nand U7446 (N_7446,N_6732,N_6590);
nor U7447 (N_7447,N_6885,N_6991);
nor U7448 (N_7448,N_6931,N_6672);
xor U7449 (N_7449,N_6930,N_6555);
xor U7450 (N_7450,N_6513,N_6716);
or U7451 (N_7451,N_6670,N_6529);
and U7452 (N_7452,N_6582,N_6825);
and U7453 (N_7453,N_6655,N_6544);
and U7454 (N_7454,N_6901,N_6593);
xor U7455 (N_7455,N_6695,N_6586);
nor U7456 (N_7456,N_6711,N_6959);
xnor U7457 (N_7457,N_6834,N_6726);
xor U7458 (N_7458,N_6515,N_6878);
and U7459 (N_7459,N_6648,N_6718);
or U7460 (N_7460,N_6976,N_6552);
and U7461 (N_7461,N_6753,N_6626);
nand U7462 (N_7462,N_6514,N_6846);
and U7463 (N_7463,N_6923,N_6773);
or U7464 (N_7464,N_6505,N_6766);
and U7465 (N_7465,N_6861,N_6822);
and U7466 (N_7466,N_6577,N_6918);
nand U7467 (N_7467,N_6690,N_6544);
nand U7468 (N_7468,N_6605,N_6550);
nand U7469 (N_7469,N_6854,N_6700);
or U7470 (N_7470,N_6988,N_6652);
or U7471 (N_7471,N_6910,N_6679);
or U7472 (N_7472,N_6899,N_6972);
and U7473 (N_7473,N_6962,N_6652);
nor U7474 (N_7474,N_6958,N_6883);
xnor U7475 (N_7475,N_6807,N_6595);
xnor U7476 (N_7476,N_6680,N_6970);
nand U7477 (N_7477,N_6612,N_6880);
nand U7478 (N_7478,N_6766,N_6935);
nor U7479 (N_7479,N_6587,N_6920);
or U7480 (N_7480,N_6871,N_6874);
xnor U7481 (N_7481,N_6772,N_6533);
nor U7482 (N_7482,N_6995,N_6780);
nor U7483 (N_7483,N_6923,N_6799);
nor U7484 (N_7484,N_6588,N_6679);
and U7485 (N_7485,N_6874,N_6699);
nor U7486 (N_7486,N_6583,N_6913);
nor U7487 (N_7487,N_6696,N_6954);
or U7488 (N_7488,N_6825,N_6609);
or U7489 (N_7489,N_6524,N_6631);
or U7490 (N_7490,N_6964,N_6912);
and U7491 (N_7491,N_6780,N_6894);
xor U7492 (N_7492,N_6853,N_6602);
or U7493 (N_7493,N_6559,N_6568);
nor U7494 (N_7494,N_6668,N_6752);
nand U7495 (N_7495,N_6734,N_6573);
xnor U7496 (N_7496,N_6566,N_6960);
and U7497 (N_7497,N_6841,N_6682);
xnor U7498 (N_7498,N_6664,N_6602);
and U7499 (N_7499,N_6740,N_6744);
and U7500 (N_7500,N_7052,N_7216);
or U7501 (N_7501,N_7431,N_7400);
nand U7502 (N_7502,N_7307,N_7011);
nand U7503 (N_7503,N_7451,N_7221);
xor U7504 (N_7504,N_7212,N_7463);
xor U7505 (N_7505,N_7142,N_7094);
or U7506 (N_7506,N_7024,N_7432);
nand U7507 (N_7507,N_7344,N_7032);
nor U7508 (N_7508,N_7040,N_7046);
xor U7509 (N_7509,N_7272,N_7487);
nor U7510 (N_7510,N_7115,N_7398);
nand U7511 (N_7511,N_7045,N_7028);
or U7512 (N_7512,N_7181,N_7140);
and U7513 (N_7513,N_7076,N_7002);
or U7514 (N_7514,N_7320,N_7240);
xnor U7515 (N_7515,N_7061,N_7030);
nand U7516 (N_7516,N_7298,N_7244);
xnor U7517 (N_7517,N_7009,N_7437);
or U7518 (N_7518,N_7004,N_7389);
or U7519 (N_7519,N_7475,N_7311);
or U7520 (N_7520,N_7473,N_7452);
xnor U7521 (N_7521,N_7044,N_7427);
or U7522 (N_7522,N_7305,N_7302);
or U7523 (N_7523,N_7345,N_7268);
nor U7524 (N_7524,N_7332,N_7394);
and U7525 (N_7525,N_7019,N_7148);
or U7526 (N_7526,N_7039,N_7220);
or U7527 (N_7527,N_7472,N_7163);
nor U7528 (N_7528,N_7100,N_7343);
or U7529 (N_7529,N_7361,N_7410);
nand U7530 (N_7530,N_7481,N_7217);
nand U7531 (N_7531,N_7036,N_7084);
xnor U7532 (N_7532,N_7326,N_7342);
xor U7533 (N_7533,N_7278,N_7460);
nor U7534 (N_7534,N_7152,N_7459);
or U7535 (N_7535,N_7286,N_7055);
nand U7536 (N_7536,N_7064,N_7035);
and U7537 (N_7537,N_7359,N_7421);
and U7538 (N_7538,N_7494,N_7187);
or U7539 (N_7539,N_7129,N_7294);
xor U7540 (N_7540,N_7133,N_7368);
nand U7541 (N_7541,N_7488,N_7184);
xnor U7542 (N_7542,N_7419,N_7139);
nand U7543 (N_7543,N_7116,N_7000);
xnor U7544 (N_7544,N_7276,N_7218);
nor U7545 (N_7545,N_7103,N_7053);
or U7546 (N_7546,N_7396,N_7380);
and U7547 (N_7547,N_7141,N_7373);
nor U7548 (N_7548,N_7067,N_7464);
nor U7549 (N_7549,N_7243,N_7239);
xnor U7550 (N_7550,N_7153,N_7223);
xnor U7551 (N_7551,N_7209,N_7059);
xnor U7552 (N_7552,N_7438,N_7407);
and U7553 (N_7553,N_7378,N_7334);
nand U7554 (N_7554,N_7126,N_7377);
or U7555 (N_7555,N_7467,N_7238);
nor U7556 (N_7556,N_7333,N_7071);
and U7557 (N_7557,N_7079,N_7446);
and U7558 (N_7558,N_7424,N_7093);
nor U7559 (N_7559,N_7253,N_7308);
or U7560 (N_7560,N_7428,N_7470);
xor U7561 (N_7561,N_7247,N_7476);
xnor U7562 (N_7562,N_7062,N_7074);
and U7563 (N_7563,N_7168,N_7383);
nand U7564 (N_7564,N_7448,N_7083);
or U7565 (N_7565,N_7167,N_7189);
and U7566 (N_7566,N_7191,N_7007);
or U7567 (N_7567,N_7041,N_7297);
xnor U7568 (N_7568,N_7327,N_7402);
and U7569 (N_7569,N_7310,N_7204);
xor U7570 (N_7570,N_7114,N_7082);
and U7571 (N_7571,N_7117,N_7057);
nor U7572 (N_7572,N_7202,N_7252);
and U7573 (N_7573,N_7051,N_7095);
xnor U7574 (N_7574,N_7384,N_7158);
and U7575 (N_7575,N_7162,N_7441);
nand U7576 (N_7576,N_7119,N_7483);
or U7577 (N_7577,N_7374,N_7038);
or U7578 (N_7578,N_7034,N_7322);
nand U7579 (N_7579,N_7329,N_7492);
nand U7580 (N_7580,N_7183,N_7185);
nor U7581 (N_7581,N_7399,N_7224);
nand U7582 (N_7582,N_7275,N_7290);
nand U7583 (N_7583,N_7109,N_7208);
and U7584 (N_7584,N_7257,N_7449);
and U7585 (N_7585,N_7161,N_7490);
nor U7586 (N_7586,N_7242,N_7271);
xor U7587 (N_7587,N_7409,N_7496);
and U7588 (N_7588,N_7469,N_7425);
xnor U7589 (N_7589,N_7358,N_7482);
nor U7590 (N_7590,N_7430,N_7388);
xnor U7591 (N_7591,N_7113,N_7391);
xor U7592 (N_7592,N_7145,N_7304);
nor U7593 (N_7593,N_7027,N_7186);
nor U7594 (N_7594,N_7069,N_7371);
nor U7595 (N_7595,N_7146,N_7177);
nor U7596 (N_7596,N_7347,N_7321);
or U7597 (N_7597,N_7078,N_7331);
and U7598 (N_7598,N_7241,N_7269);
xnor U7599 (N_7599,N_7013,N_7154);
xnor U7600 (N_7600,N_7401,N_7107);
and U7601 (N_7601,N_7435,N_7357);
and U7602 (N_7602,N_7077,N_7075);
or U7603 (N_7603,N_7102,N_7376);
and U7604 (N_7604,N_7413,N_7325);
or U7605 (N_7605,N_7337,N_7447);
and U7606 (N_7606,N_7461,N_7457);
nand U7607 (N_7607,N_7355,N_7065);
nor U7608 (N_7608,N_7196,N_7287);
nand U7609 (N_7609,N_7335,N_7166);
nor U7610 (N_7610,N_7215,N_7106);
nor U7611 (N_7611,N_7160,N_7281);
nor U7612 (N_7612,N_7037,N_7291);
or U7613 (N_7613,N_7289,N_7439);
nor U7614 (N_7614,N_7063,N_7245);
nand U7615 (N_7615,N_7336,N_7198);
nand U7616 (N_7616,N_7403,N_7200);
and U7617 (N_7617,N_7135,N_7195);
or U7618 (N_7618,N_7203,N_7293);
xnor U7619 (N_7619,N_7128,N_7073);
or U7620 (N_7620,N_7138,N_7232);
nand U7621 (N_7621,N_7414,N_7277);
and U7622 (N_7622,N_7043,N_7426);
nand U7623 (N_7623,N_7453,N_7156);
xnor U7624 (N_7624,N_7248,N_7338);
and U7625 (N_7625,N_7340,N_7369);
and U7626 (N_7626,N_7025,N_7354);
or U7627 (N_7627,N_7348,N_7323);
nor U7628 (N_7628,N_7349,N_7397);
nand U7629 (N_7629,N_7315,N_7370);
nand U7630 (N_7630,N_7246,N_7033);
nand U7631 (N_7631,N_7176,N_7270);
and U7632 (N_7632,N_7143,N_7020);
or U7633 (N_7633,N_7211,N_7003);
and U7634 (N_7634,N_7405,N_7468);
or U7635 (N_7635,N_7412,N_7456);
xor U7636 (N_7636,N_7282,N_7018);
and U7637 (N_7637,N_7406,N_7295);
nor U7638 (N_7638,N_7173,N_7454);
nand U7639 (N_7639,N_7471,N_7313);
or U7640 (N_7640,N_7021,N_7360);
or U7641 (N_7641,N_7324,N_7207);
nand U7642 (N_7642,N_7047,N_7008);
nand U7643 (N_7643,N_7192,N_7292);
nor U7644 (N_7644,N_7480,N_7171);
nor U7645 (N_7645,N_7060,N_7352);
and U7646 (N_7646,N_7120,N_7404);
xnor U7647 (N_7647,N_7070,N_7267);
nand U7648 (N_7648,N_7134,N_7213);
or U7649 (N_7649,N_7089,N_7462);
and U7650 (N_7650,N_7111,N_7101);
xor U7651 (N_7651,N_7306,N_7085);
nor U7652 (N_7652,N_7440,N_7390);
or U7653 (N_7653,N_7118,N_7042);
xor U7654 (N_7654,N_7231,N_7386);
or U7655 (N_7655,N_7288,N_7251);
xnor U7656 (N_7656,N_7300,N_7010);
nand U7657 (N_7657,N_7097,N_7048);
xnor U7658 (N_7658,N_7182,N_7341);
nor U7659 (N_7659,N_7169,N_7236);
and U7660 (N_7660,N_7266,N_7445);
xnor U7661 (N_7661,N_7458,N_7455);
or U7662 (N_7662,N_7433,N_7144);
nor U7663 (N_7663,N_7350,N_7316);
nor U7664 (N_7664,N_7127,N_7026);
nor U7665 (N_7665,N_7318,N_7249);
xnor U7666 (N_7666,N_7356,N_7014);
nand U7667 (N_7667,N_7328,N_7330);
nand U7668 (N_7668,N_7372,N_7319);
and U7669 (N_7669,N_7180,N_7222);
or U7670 (N_7670,N_7050,N_7493);
xor U7671 (N_7671,N_7382,N_7484);
or U7672 (N_7672,N_7080,N_7339);
and U7673 (N_7673,N_7365,N_7489);
or U7674 (N_7674,N_7104,N_7068);
nor U7675 (N_7675,N_7017,N_7193);
and U7676 (N_7676,N_7006,N_7346);
and U7677 (N_7677,N_7015,N_7029);
nor U7678 (N_7678,N_7299,N_7314);
and U7679 (N_7679,N_7112,N_7258);
nor U7680 (N_7680,N_7124,N_7172);
nand U7681 (N_7681,N_7157,N_7479);
xnor U7682 (N_7682,N_7049,N_7132);
or U7683 (N_7683,N_7175,N_7385);
and U7684 (N_7684,N_7417,N_7150);
or U7685 (N_7685,N_7229,N_7283);
or U7686 (N_7686,N_7205,N_7081);
xnor U7687 (N_7687,N_7091,N_7194);
and U7688 (N_7688,N_7178,N_7174);
and U7689 (N_7689,N_7056,N_7442);
or U7690 (N_7690,N_7263,N_7273);
or U7691 (N_7691,N_7147,N_7265);
or U7692 (N_7692,N_7197,N_7415);
nor U7693 (N_7693,N_7498,N_7123);
or U7694 (N_7694,N_7199,N_7170);
nor U7695 (N_7695,N_7495,N_7429);
nand U7696 (N_7696,N_7230,N_7317);
nand U7697 (N_7697,N_7225,N_7309);
nor U7698 (N_7698,N_7096,N_7416);
nand U7699 (N_7699,N_7086,N_7279);
xor U7700 (N_7700,N_7436,N_7227);
nand U7701 (N_7701,N_7485,N_7151);
xor U7702 (N_7702,N_7408,N_7363);
nand U7703 (N_7703,N_7450,N_7131);
and U7704 (N_7704,N_7274,N_7098);
or U7705 (N_7705,N_7280,N_7353);
nor U7706 (N_7706,N_7214,N_7165);
or U7707 (N_7707,N_7159,N_7054);
or U7708 (N_7708,N_7110,N_7023);
nand U7709 (N_7709,N_7022,N_7201);
nor U7710 (N_7710,N_7137,N_7234);
xor U7711 (N_7711,N_7387,N_7179);
nor U7712 (N_7712,N_7235,N_7058);
and U7713 (N_7713,N_7233,N_7303);
xor U7714 (N_7714,N_7255,N_7420);
xnor U7715 (N_7715,N_7136,N_7190);
nor U7716 (N_7716,N_7066,N_7099);
xnor U7717 (N_7717,N_7226,N_7121);
nand U7718 (N_7718,N_7087,N_7262);
or U7719 (N_7719,N_7395,N_7250);
xnor U7720 (N_7720,N_7497,N_7005);
or U7721 (N_7721,N_7375,N_7351);
and U7722 (N_7722,N_7219,N_7422);
and U7723 (N_7723,N_7465,N_7379);
nand U7724 (N_7724,N_7108,N_7254);
or U7725 (N_7725,N_7256,N_7092);
or U7726 (N_7726,N_7155,N_7486);
xor U7727 (N_7727,N_7001,N_7474);
and U7728 (N_7728,N_7392,N_7364);
and U7729 (N_7729,N_7122,N_7149);
or U7730 (N_7730,N_7264,N_7125);
nor U7731 (N_7731,N_7411,N_7296);
nand U7732 (N_7732,N_7499,N_7393);
and U7733 (N_7733,N_7418,N_7228);
nor U7734 (N_7734,N_7362,N_7284);
nand U7735 (N_7735,N_7444,N_7012);
nand U7736 (N_7736,N_7105,N_7381);
nor U7737 (N_7737,N_7491,N_7466);
nor U7738 (N_7738,N_7072,N_7188);
and U7739 (N_7739,N_7301,N_7164);
xor U7740 (N_7740,N_7285,N_7434);
nand U7741 (N_7741,N_7477,N_7130);
or U7742 (N_7742,N_7260,N_7423);
nor U7743 (N_7743,N_7312,N_7237);
or U7744 (N_7744,N_7031,N_7016);
or U7745 (N_7745,N_7090,N_7443);
xor U7746 (N_7746,N_7478,N_7367);
nand U7747 (N_7747,N_7366,N_7206);
nand U7748 (N_7748,N_7259,N_7088);
xnor U7749 (N_7749,N_7210,N_7261);
or U7750 (N_7750,N_7242,N_7284);
xnor U7751 (N_7751,N_7161,N_7234);
nand U7752 (N_7752,N_7088,N_7101);
xor U7753 (N_7753,N_7313,N_7262);
nor U7754 (N_7754,N_7012,N_7141);
and U7755 (N_7755,N_7001,N_7494);
nand U7756 (N_7756,N_7456,N_7149);
or U7757 (N_7757,N_7056,N_7399);
or U7758 (N_7758,N_7184,N_7031);
nor U7759 (N_7759,N_7206,N_7169);
nand U7760 (N_7760,N_7262,N_7307);
nor U7761 (N_7761,N_7034,N_7368);
nor U7762 (N_7762,N_7098,N_7265);
xnor U7763 (N_7763,N_7117,N_7035);
or U7764 (N_7764,N_7462,N_7339);
and U7765 (N_7765,N_7300,N_7038);
or U7766 (N_7766,N_7088,N_7038);
or U7767 (N_7767,N_7235,N_7001);
and U7768 (N_7768,N_7412,N_7010);
nand U7769 (N_7769,N_7099,N_7499);
nor U7770 (N_7770,N_7440,N_7409);
xnor U7771 (N_7771,N_7405,N_7474);
or U7772 (N_7772,N_7025,N_7207);
nor U7773 (N_7773,N_7492,N_7079);
and U7774 (N_7774,N_7181,N_7051);
or U7775 (N_7775,N_7098,N_7003);
and U7776 (N_7776,N_7488,N_7125);
or U7777 (N_7777,N_7034,N_7291);
and U7778 (N_7778,N_7304,N_7323);
xnor U7779 (N_7779,N_7172,N_7241);
nor U7780 (N_7780,N_7334,N_7442);
xor U7781 (N_7781,N_7163,N_7415);
or U7782 (N_7782,N_7284,N_7387);
nor U7783 (N_7783,N_7265,N_7029);
and U7784 (N_7784,N_7448,N_7247);
xor U7785 (N_7785,N_7050,N_7256);
xor U7786 (N_7786,N_7241,N_7198);
nor U7787 (N_7787,N_7483,N_7152);
or U7788 (N_7788,N_7382,N_7415);
or U7789 (N_7789,N_7378,N_7027);
or U7790 (N_7790,N_7319,N_7450);
or U7791 (N_7791,N_7424,N_7018);
or U7792 (N_7792,N_7353,N_7144);
and U7793 (N_7793,N_7112,N_7177);
nand U7794 (N_7794,N_7490,N_7015);
nand U7795 (N_7795,N_7141,N_7130);
nand U7796 (N_7796,N_7329,N_7226);
or U7797 (N_7797,N_7488,N_7205);
xor U7798 (N_7798,N_7417,N_7234);
nor U7799 (N_7799,N_7279,N_7337);
nand U7800 (N_7800,N_7467,N_7064);
or U7801 (N_7801,N_7250,N_7144);
and U7802 (N_7802,N_7333,N_7260);
xnor U7803 (N_7803,N_7433,N_7003);
nor U7804 (N_7804,N_7127,N_7181);
nor U7805 (N_7805,N_7368,N_7328);
and U7806 (N_7806,N_7120,N_7452);
nor U7807 (N_7807,N_7250,N_7253);
xnor U7808 (N_7808,N_7434,N_7447);
xor U7809 (N_7809,N_7306,N_7309);
or U7810 (N_7810,N_7370,N_7111);
nand U7811 (N_7811,N_7121,N_7106);
xor U7812 (N_7812,N_7017,N_7464);
or U7813 (N_7813,N_7472,N_7074);
nor U7814 (N_7814,N_7492,N_7080);
nand U7815 (N_7815,N_7086,N_7462);
or U7816 (N_7816,N_7322,N_7429);
nor U7817 (N_7817,N_7358,N_7021);
or U7818 (N_7818,N_7450,N_7446);
nor U7819 (N_7819,N_7045,N_7201);
nand U7820 (N_7820,N_7287,N_7485);
xor U7821 (N_7821,N_7329,N_7349);
nand U7822 (N_7822,N_7493,N_7146);
xor U7823 (N_7823,N_7325,N_7490);
nor U7824 (N_7824,N_7027,N_7374);
or U7825 (N_7825,N_7059,N_7489);
or U7826 (N_7826,N_7269,N_7333);
nor U7827 (N_7827,N_7231,N_7149);
nand U7828 (N_7828,N_7167,N_7425);
or U7829 (N_7829,N_7005,N_7297);
and U7830 (N_7830,N_7393,N_7247);
or U7831 (N_7831,N_7020,N_7232);
and U7832 (N_7832,N_7259,N_7284);
or U7833 (N_7833,N_7001,N_7350);
nor U7834 (N_7834,N_7006,N_7110);
and U7835 (N_7835,N_7426,N_7244);
nand U7836 (N_7836,N_7313,N_7015);
and U7837 (N_7837,N_7470,N_7122);
or U7838 (N_7838,N_7200,N_7389);
nor U7839 (N_7839,N_7303,N_7011);
or U7840 (N_7840,N_7043,N_7384);
nand U7841 (N_7841,N_7463,N_7177);
and U7842 (N_7842,N_7481,N_7416);
xor U7843 (N_7843,N_7296,N_7133);
or U7844 (N_7844,N_7128,N_7133);
or U7845 (N_7845,N_7314,N_7322);
xor U7846 (N_7846,N_7227,N_7489);
nor U7847 (N_7847,N_7082,N_7021);
xnor U7848 (N_7848,N_7310,N_7262);
and U7849 (N_7849,N_7467,N_7435);
nand U7850 (N_7850,N_7263,N_7484);
xnor U7851 (N_7851,N_7471,N_7457);
and U7852 (N_7852,N_7332,N_7352);
and U7853 (N_7853,N_7039,N_7020);
xnor U7854 (N_7854,N_7202,N_7423);
nor U7855 (N_7855,N_7395,N_7376);
nor U7856 (N_7856,N_7464,N_7481);
or U7857 (N_7857,N_7327,N_7436);
and U7858 (N_7858,N_7070,N_7340);
nand U7859 (N_7859,N_7352,N_7337);
or U7860 (N_7860,N_7382,N_7219);
nand U7861 (N_7861,N_7138,N_7314);
or U7862 (N_7862,N_7305,N_7391);
xor U7863 (N_7863,N_7224,N_7086);
nor U7864 (N_7864,N_7341,N_7200);
nor U7865 (N_7865,N_7128,N_7025);
nand U7866 (N_7866,N_7017,N_7104);
nand U7867 (N_7867,N_7097,N_7358);
nand U7868 (N_7868,N_7135,N_7273);
nand U7869 (N_7869,N_7026,N_7477);
or U7870 (N_7870,N_7439,N_7126);
and U7871 (N_7871,N_7141,N_7411);
nand U7872 (N_7872,N_7024,N_7172);
and U7873 (N_7873,N_7052,N_7287);
xnor U7874 (N_7874,N_7060,N_7117);
and U7875 (N_7875,N_7489,N_7346);
nor U7876 (N_7876,N_7207,N_7425);
or U7877 (N_7877,N_7333,N_7351);
xor U7878 (N_7878,N_7171,N_7491);
nor U7879 (N_7879,N_7323,N_7145);
or U7880 (N_7880,N_7142,N_7091);
nor U7881 (N_7881,N_7028,N_7228);
nand U7882 (N_7882,N_7419,N_7063);
and U7883 (N_7883,N_7022,N_7228);
nor U7884 (N_7884,N_7449,N_7055);
nor U7885 (N_7885,N_7488,N_7476);
or U7886 (N_7886,N_7084,N_7231);
nor U7887 (N_7887,N_7268,N_7086);
and U7888 (N_7888,N_7175,N_7422);
or U7889 (N_7889,N_7270,N_7458);
xnor U7890 (N_7890,N_7253,N_7165);
nand U7891 (N_7891,N_7193,N_7317);
nand U7892 (N_7892,N_7067,N_7355);
nor U7893 (N_7893,N_7113,N_7445);
and U7894 (N_7894,N_7030,N_7246);
and U7895 (N_7895,N_7301,N_7109);
or U7896 (N_7896,N_7409,N_7248);
and U7897 (N_7897,N_7226,N_7235);
or U7898 (N_7898,N_7248,N_7493);
xnor U7899 (N_7899,N_7158,N_7109);
or U7900 (N_7900,N_7364,N_7139);
or U7901 (N_7901,N_7449,N_7311);
and U7902 (N_7902,N_7477,N_7268);
and U7903 (N_7903,N_7280,N_7119);
nor U7904 (N_7904,N_7481,N_7128);
and U7905 (N_7905,N_7066,N_7423);
xnor U7906 (N_7906,N_7433,N_7335);
nand U7907 (N_7907,N_7498,N_7336);
nor U7908 (N_7908,N_7327,N_7468);
nor U7909 (N_7909,N_7253,N_7340);
xnor U7910 (N_7910,N_7099,N_7285);
and U7911 (N_7911,N_7424,N_7054);
nand U7912 (N_7912,N_7485,N_7185);
nand U7913 (N_7913,N_7453,N_7456);
nand U7914 (N_7914,N_7452,N_7203);
nor U7915 (N_7915,N_7329,N_7365);
nand U7916 (N_7916,N_7386,N_7265);
nand U7917 (N_7917,N_7489,N_7169);
or U7918 (N_7918,N_7341,N_7299);
and U7919 (N_7919,N_7484,N_7201);
nor U7920 (N_7920,N_7404,N_7163);
or U7921 (N_7921,N_7137,N_7301);
and U7922 (N_7922,N_7040,N_7419);
nand U7923 (N_7923,N_7337,N_7050);
or U7924 (N_7924,N_7160,N_7317);
or U7925 (N_7925,N_7015,N_7323);
xnor U7926 (N_7926,N_7098,N_7473);
xor U7927 (N_7927,N_7413,N_7109);
or U7928 (N_7928,N_7498,N_7475);
xor U7929 (N_7929,N_7152,N_7155);
and U7930 (N_7930,N_7063,N_7458);
nand U7931 (N_7931,N_7034,N_7220);
nor U7932 (N_7932,N_7146,N_7316);
or U7933 (N_7933,N_7147,N_7056);
nor U7934 (N_7934,N_7443,N_7261);
nand U7935 (N_7935,N_7430,N_7163);
nand U7936 (N_7936,N_7105,N_7062);
xnor U7937 (N_7937,N_7098,N_7429);
nand U7938 (N_7938,N_7086,N_7490);
and U7939 (N_7939,N_7214,N_7223);
nor U7940 (N_7940,N_7398,N_7021);
xor U7941 (N_7941,N_7428,N_7224);
or U7942 (N_7942,N_7366,N_7186);
and U7943 (N_7943,N_7197,N_7322);
and U7944 (N_7944,N_7085,N_7308);
xnor U7945 (N_7945,N_7000,N_7427);
and U7946 (N_7946,N_7360,N_7069);
nand U7947 (N_7947,N_7154,N_7001);
or U7948 (N_7948,N_7059,N_7468);
nor U7949 (N_7949,N_7019,N_7128);
nand U7950 (N_7950,N_7033,N_7208);
nand U7951 (N_7951,N_7285,N_7237);
nand U7952 (N_7952,N_7137,N_7440);
nand U7953 (N_7953,N_7052,N_7088);
nor U7954 (N_7954,N_7351,N_7231);
nor U7955 (N_7955,N_7008,N_7494);
nand U7956 (N_7956,N_7025,N_7246);
or U7957 (N_7957,N_7073,N_7120);
and U7958 (N_7958,N_7097,N_7104);
xnor U7959 (N_7959,N_7290,N_7158);
nor U7960 (N_7960,N_7242,N_7101);
nor U7961 (N_7961,N_7202,N_7009);
nor U7962 (N_7962,N_7270,N_7193);
xnor U7963 (N_7963,N_7372,N_7011);
or U7964 (N_7964,N_7462,N_7082);
and U7965 (N_7965,N_7434,N_7382);
nand U7966 (N_7966,N_7077,N_7210);
or U7967 (N_7967,N_7098,N_7067);
or U7968 (N_7968,N_7355,N_7043);
and U7969 (N_7969,N_7277,N_7177);
nand U7970 (N_7970,N_7369,N_7421);
or U7971 (N_7971,N_7234,N_7217);
nand U7972 (N_7972,N_7100,N_7011);
or U7973 (N_7973,N_7342,N_7423);
nor U7974 (N_7974,N_7048,N_7456);
or U7975 (N_7975,N_7308,N_7286);
or U7976 (N_7976,N_7479,N_7026);
or U7977 (N_7977,N_7120,N_7330);
nand U7978 (N_7978,N_7263,N_7391);
or U7979 (N_7979,N_7412,N_7047);
and U7980 (N_7980,N_7050,N_7442);
nor U7981 (N_7981,N_7136,N_7077);
or U7982 (N_7982,N_7357,N_7045);
or U7983 (N_7983,N_7212,N_7100);
xnor U7984 (N_7984,N_7440,N_7064);
nor U7985 (N_7985,N_7288,N_7386);
and U7986 (N_7986,N_7497,N_7058);
nor U7987 (N_7987,N_7465,N_7385);
or U7988 (N_7988,N_7071,N_7028);
and U7989 (N_7989,N_7352,N_7241);
and U7990 (N_7990,N_7080,N_7118);
and U7991 (N_7991,N_7240,N_7188);
nand U7992 (N_7992,N_7183,N_7392);
nand U7993 (N_7993,N_7112,N_7293);
or U7994 (N_7994,N_7456,N_7422);
or U7995 (N_7995,N_7040,N_7028);
xor U7996 (N_7996,N_7271,N_7338);
nand U7997 (N_7997,N_7204,N_7209);
xnor U7998 (N_7998,N_7106,N_7322);
and U7999 (N_7999,N_7378,N_7331);
xnor U8000 (N_8000,N_7740,N_7999);
nand U8001 (N_8001,N_7530,N_7536);
nand U8002 (N_8002,N_7787,N_7823);
xnor U8003 (N_8003,N_7622,N_7901);
and U8004 (N_8004,N_7966,N_7567);
or U8005 (N_8005,N_7576,N_7902);
xnor U8006 (N_8006,N_7569,N_7839);
nor U8007 (N_8007,N_7580,N_7851);
or U8008 (N_8008,N_7503,N_7977);
nor U8009 (N_8009,N_7895,N_7518);
nand U8010 (N_8010,N_7770,N_7693);
and U8011 (N_8011,N_7786,N_7736);
nor U8012 (N_8012,N_7613,N_7689);
nand U8013 (N_8013,N_7719,N_7645);
xnor U8014 (N_8014,N_7991,N_7983);
or U8015 (N_8015,N_7961,N_7779);
and U8016 (N_8016,N_7629,N_7612);
nor U8017 (N_8017,N_7735,N_7637);
nand U8018 (N_8018,N_7797,N_7739);
nand U8019 (N_8019,N_7701,N_7582);
nand U8020 (N_8020,N_7638,N_7842);
nand U8021 (N_8021,N_7877,N_7956);
or U8022 (N_8022,N_7650,N_7552);
nor U8023 (N_8023,N_7863,N_7684);
and U8024 (N_8024,N_7834,N_7831);
nand U8025 (N_8025,N_7812,N_7568);
and U8026 (N_8026,N_7829,N_7540);
or U8027 (N_8027,N_7625,N_7950);
and U8028 (N_8028,N_7601,N_7589);
nor U8029 (N_8029,N_7727,N_7942);
nor U8030 (N_8030,N_7690,N_7686);
nand U8031 (N_8031,N_7941,N_7705);
or U8032 (N_8032,N_7820,N_7913);
xor U8033 (N_8033,N_7806,N_7971);
and U8034 (N_8034,N_7720,N_7677);
and U8035 (N_8035,N_7934,N_7867);
nand U8036 (N_8036,N_7709,N_7696);
and U8037 (N_8037,N_7874,N_7879);
and U8038 (N_8038,N_7657,N_7848);
or U8039 (N_8039,N_7938,N_7716);
nand U8040 (N_8040,N_7781,N_7918);
nand U8041 (N_8041,N_7746,N_7558);
or U8042 (N_8042,N_7575,N_7703);
or U8043 (N_8043,N_7973,N_7619);
and U8044 (N_8044,N_7549,N_7949);
nor U8045 (N_8045,N_7960,N_7868);
and U8046 (N_8046,N_7544,N_7803);
nor U8047 (N_8047,N_7923,N_7826);
nand U8048 (N_8048,N_7886,N_7987);
nand U8049 (N_8049,N_7509,N_7627);
or U8050 (N_8050,N_7832,N_7931);
or U8051 (N_8051,N_7870,N_7771);
and U8052 (N_8052,N_7587,N_7539);
or U8053 (N_8053,N_7741,N_7819);
nand U8054 (N_8054,N_7535,N_7533);
nand U8055 (N_8055,N_7715,N_7651);
and U8056 (N_8056,N_7501,N_7976);
or U8057 (N_8057,N_7659,N_7556);
xor U8058 (N_8058,N_7598,N_7850);
xor U8059 (N_8059,N_7652,N_7808);
nand U8060 (N_8060,N_7661,N_7989);
nand U8061 (N_8061,N_7745,N_7835);
nor U8062 (N_8062,N_7626,N_7892);
nand U8063 (N_8063,N_7752,N_7898);
xor U8064 (N_8064,N_7673,N_7981);
nor U8065 (N_8065,N_7641,N_7609);
and U8066 (N_8066,N_7856,N_7714);
or U8067 (N_8067,N_7665,N_7880);
nand U8068 (N_8068,N_7744,N_7894);
nor U8069 (N_8069,N_7859,N_7517);
and U8070 (N_8070,N_7882,N_7708);
nand U8071 (N_8071,N_7506,N_7970);
nand U8072 (N_8072,N_7957,N_7513);
and U8073 (N_8073,N_7699,N_7920);
and U8074 (N_8074,N_7852,N_7907);
nor U8075 (N_8075,N_7903,N_7774);
nand U8076 (N_8076,N_7900,N_7982);
xor U8077 (N_8077,N_7995,N_7769);
xor U8078 (N_8078,N_7633,N_7584);
nor U8079 (N_8079,N_7700,N_7878);
nor U8080 (N_8080,N_7897,N_7866);
xor U8081 (N_8081,N_7847,N_7909);
nand U8082 (N_8082,N_7554,N_7801);
xnor U8083 (N_8083,N_7908,N_7534);
or U8084 (N_8084,N_7743,N_7630);
or U8085 (N_8085,N_7671,N_7865);
nor U8086 (N_8086,N_7845,N_7573);
and U8087 (N_8087,N_7564,N_7804);
xor U8088 (N_8088,N_7784,N_7610);
or U8089 (N_8089,N_7818,N_7994);
xor U8090 (N_8090,N_7937,N_7927);
and U8091 (N_8091,N_7644,N_7559);
or U8092 (N_8092,N_7723,N_7667);
or U8093 (N_8093,N_7821,N_7572);
or U8094 (N_8094,N_7563,N_7911);
nor U8095 (N_8095,N_7551,N_7958);
nor U8096 (N_8096,N_7597,N_7824);
nand U8097 (N_8097,N_7545,N_7749);
xnor U8098 (N_8098,N_7682,N_7537);
nor U8099 (N_8099,N_7516,N_7574);
and U8100 (N_8100,N_7924,N_7791);
or U8101 (N_8101,N_7946,N_7777);
xnor U8102 (N_8102,N_7663,N_7889);
nor U8103 (N_8103,N_7766,N_7944);
xor U8104 (N_8104,N_7793,N_7706);
or U8105 (N_8105,N_7760,N_7730);
nor U8106 (N_8106,N_7802,N_7885);
or U8107 (N_8107,N_7822,N_7595);
nand U8108 (N_8108,N_7840,N_7914);
or U8109 (N_8109,N_7617,N_7658);
nand U8110 (N_8110,N_7899,N_7917);
and U8111 (N_8111,N_7594,N_7577);
xnor U8112 (N_8112,N_7881,N_7546);
and U8113 (N_8113,N_7768,N_7952);
and U8114 (N_8114,N_7562,N_7904);
and U8115 (N_8115,N_7861,N_7732);
nand U8116 (N_8116,N_7519,N_7916);
nand U8117 (N_8117,N_7986,N_7799);
and U8118 (N_8118,N_7890,N_7965);
nand U8119 (N_8119,N_7759,N_7765);
xor U8120 (N_8120,N_7853,N_7500);
nor U8121 (N_8121,N_7997,N_7883);
and U8122 (N_8122,N_7836,N_7733);
or U8123 (N_8123,N_7581,N_7600);
or U8124 (N_8124,N_7555,N_7921);
xnor U8125 (N_8125,N_7943,N_7541);
or U8126 (N_8126,N_7707,N_7547);
nor U8127 (N_8127,N_7816,N_7713);
nor U8128 (N_8128,N_7968,N_7782);
nor U8129 (N_8129,N_7578,N_7694);
xnor U8130 (N_8130,N_7754,N_7685);
or U8131 (N_8131,N_7928,N_7653);
nand U8132 (N_8132,N_7849,N_7620);
nor U8133 (N_8133,N_7514,N_7725);
nor U8134 (N_8134,N_7930,N_7654);
nor U8135 (N_8135,N_7543,N_7773);
or U8136 (N_8136,N_7825,N_7811);
nand U8137 (N_8137,N_7583,N_7596);
and U8138 (N_8138,N_7523,N_7862);
xor U8139 (N_8139,N_7756,N_7721);
or U8140 (N_8140,N_7758,N_7993);
nor U8141 (N_8141,N_7691,N_7780);
xnor U8142 (N_8142,N_7929,N_7967);
and U8143 (N_8143,N_7527,N_7557);
or U8144 (N_8144,N_7794,N_7912);
xnor U8145 (N_8145,N_7675,N_7750);
nand U8146 (N_8146,N_7717,N_7615);
and U8147 (N_8147,N_7896,N_7510);
nor U8148 (N_8148,N_7778,N_7800);
nand U8149 (N_8149,N_7979,N_7603);
or U8150 (N_8150,N_7962,N_7692);
nor U8151 (N_8151,N_7593,N_7783);
or U8152 (N_8152,N_7560,N_7605);
xnor U8153 (N_8153,N_7790,N_7525);
nor U8154 (N_8154,N_7586,N_7561);
and U8155 (N_8155,N_7712,N_7634);
or U8156 (N_8156,N_7992,N_7642);
nor U8157 (N_8157,N_7767,N_7975);
xor U8158 (N_8158,N_7954,N_7963);
nand U8159 (N_8159,N_7893,N_7502);
xnor U8160 (N_8160,N_7761,N_7742);
or U8161 (N_8161,N_7591,N_7857);
xnor U8162 (N_8162,N_7672,N_7662);
xor U8163 (N_8163,N_7623,N_7817);
nand U8164 (N_8164,N_7538,N_7932);
xnor U8165 (N_8165,N_7762,N_7726);
nand U8166 (N_8166,N_7796,N_7570);
nand U8167 (N_8167,N_7649,N_7854);
and U8168 (N_8168,N_7830,N_7520);
or U8169 (N_8169,N_7788,N_7905);
nand U8170 (N_8170,N_7515,N_7776);
and U8171 (N_8171,N_7674,N_7844);
xor U8172 (N_8172,N_7805,N_7599);
and U8173 (N_8173,N_7687,N_7953);
nand U8174 (N_8174,N_7608,N_7676);
and U8175 (N_8175,N_7571,N_7951);
or U8176 (N_8176,N_7925,N_7566);
nor U8177 (N_8177,N_7876,N_7646);
and U8178 (N_8178,N_7734,N_7656);
or U8179 (N_8179,N_7698,N_7526);
nor U8180 (N_8180,N_7606,N_7512);
or U8181 (N_8181,N_7948,N_7919);
nor U8182 (N_8182,N_7984,N_7604);
nand U8183 (N_8183,N_7548,N_7959);
and U8184 (N_8184,N_7611,N_7636);
or U8185 (N_8185,N_7872,N_7990);
and U8186 (N_8186,N_7910,N_7504);
or U8187 (N_8187,N_7521,N_7933);
nor U8188 (N_8188,N_7813,N_7647);
nor U8189 (N_8189,N_7710,N_7731);
and U8190 (N_8190,N_7585,N_7843);
and U8191 (N_8191,N_7751,N_7532);
and U8192 (N_8192,N_7639,N_7680);
nor U8193 (N_8193,N_7632,N_7669);
and U8194 (N_8194,N_7624,N_7827);
nand U8195 (N_8195,N_7565,N_7670);
and U8196 (N_8196,N_7855,N_7964);
nor U8197 (N_8197,N_7815,N_7947);
or U8198 (N_8198,N_7763,N_7755);
and U8199 (N_8199,N_7785,N_7722);
and U8200 (N_8200,N_7996,N_7508);
or U8201 (N_8201,N_7764,N_7858);
nand U8202 (N_8202,N_7798,N_7621);
or U8203 (N_8203,N_7860,N_7747);
or U8204 (N_8204,N_7795,N_7884);
and U8205 (N_8205,N_7915,N_7607);
xor U8206 (N_8206,N_7511,N_7814);
or U8207 (N_8207,N_7697,N_7792);
and U8208 (N_8208,N_7875,N_7678);
and U8209 (N_8209,N_7969,N_7688);
nand U8210 (N_8210,N_7702,N_7704);
and U8211 (N_8211,N_7728,N_7891);
xor U8212 (N_8212,N_7998,N_7550);
nand U8213 (N_8213,N_7757,N_7588);
nand U8214 (N_8214,N_7592,N_7939);
nor U8215 (N_8215,N_7887,N_7945);
xor U8216 (N_8216,N_7524,N_7666);
nor U8217 (N_8217,N_7590,N_7837);
or U8218 (N_8218,N_7789,N_7980);
and U8219 (N_8219,N_7628,N_7873);
nand U8220 (N_8220,N_7936,N_7972);
nand U8221 (N_8221,N_7664,N_7528);
or U8222 (N_8222,N_7955,N_7888);
or U8223 (N_8223,N_7974,N_7655);
nand U8224 (N_8224,N_7640,N_7711);
and U8225 (N_8225,N_7846,N_7507);
nand U8226 (N_8226,N_7505,N_7668);
and U8227 (N_8227,N_7579,N_7869);
nor U8228 (N_8228,N_7695,N_7738);
nor U8229 (N_8229,N_7737,N_7522);
nand U8230 (N_8230,N_7616,N_7833);
nor U8231 (N_8231,N_7871,N_7940);
xnor U8232 (N_8232,N_7828,N_7807);
nor U8233 (N_8233,N_7810,N_7926);
and U8234 (N_8234,N_7838,N_7841);
nor U8235 (N_8235,N_7643,N_7775);
xnor U8236 (N_8236,N_7922,N_7935);
nor U8237 (N_8237,N_7724,N_7602);
nor U8238 (N_8238,N_7531,N_7635);
xor U8239 (N_8239,N_7864,N_7988);
nor U8240 (N_8240,N_7542,N_7985);
or U8241 (N_8241,N_7648,N_7978);
nand U8242 (N_8242,N_7772,N_7660);
nand U8243 (N_8243,N_7753,N_7679);
or U8244 (N_8244,N_7631,N_7718);
nand U8245 (N_8245,N_7809,N_7529);
and U8246 (N_8246,N_7748,N_7614);
and U8247 (N_8247,N_7681,N_7729);
xnor U8248 (N_8248,N_7683,N_7553);
nor U8249 (N_8249,N_7906,N_7618);
or U8250 (N_8250,N_7851,N_7543);
nand U8251 (N_8251,N_7812,N_7730);
xor U8252 (N_8252,N_7568,N_7500);
nor U8253 (N_8253,N_7650,N_7820);
and U8254 (N_8254,N_7541,N_7519);
or U8255 (N_8255,N_7787,N_7613);
or U8256 (N_8256,N_7945,N_7682);
nor U8257 (N_8257,N_7613,N_7826);
or U8258 (N_8258,N_7955,N_7975);
nor U8259 (N_8259,N_7807,N_7832);
nor U8260 (N_8260,N_7717,N_7660);
and U8261 (N_8261,N_7929,N_7813);
nor U8262 (N_8262,N_7710,N_7848);
or U8263 (N_8263,N_7848,N_7641);
xor U8264 (N_8264,N_7666,N_7532);
or U8265 (N_8265,N_7522,N_7546);
or U8266 (N_8266,N_7732,N_7920);
or U8267 (N_8267,N_7846,N_7624);
xor U8268 (N_8268,N_7728,N_7851);
and U8269 (N_8269,N_7554,N_7572);
or U8270 (N_8270,N_7972,N_7664);
nand U8271 (N_8271,N_7593,N_7618);
or U8272 (N_8272,N_7534,N_7824);
xnor U8273 (N_8273,N_7798,N_7903);
xor U8274 (N_8274,N_7563,N_7599);
and U8275 (N_8275,N_7513,N_7984);
or U8276 (N_8276,N_7512,N_7789);
xor U8277 (N_8277,N_7537,N_7956);
nor U8278 (N_8278,N_7864,N_7654);
or U8279 (N_8279,N_7841,N_7797);
nor U8280 (N_8280,N_7863,N_7758);
or U8281 (N_8281,N_7577,N_7870);
and U8282 (N_8282,N_7674,N_7741);
xnor U8283 (N_8283,N_7765,N_7902);
or U8284 (N_8284,N_7536,N_7936);
xnor U8285 (N_8285,N_7551,N_7586);
nand U8286 (N_8286,N_7776,N_7635);
nor U8287 (N_8287,N_7649,N_7968);
nor U8288 (N_8288,N_7967,N_7732);
nand U8289 (N_8289,N_7524,N_7955);
nand U8290 (N_8290,N_7852,N_7762);
or U8291 (N_8291,N_7620,N_7942);
xnor U8292 (N_8292,N_7508,N_7772);
xnor U8293 (N_8293,N_7987,N_7878);
and U8294 (N_8294,N_7646,N_7932);
nand U8295 (N_8295,N_7680,N_7572);
nor U8296 (N_8296,N_7500,N_7995);
xor U8297 (N_8297,N_7864,N_7611);
and U8298 (N_8298,N_7739,N_7700);
xor U8299 (N_8299,N_7565,N_7533);
xor U8300 (N_8300,N_7854,N_7857);
xor U8301 (N_8301,N_7940,N_7501);
nor U8302 (N_8302,N_7932,N_7694);
nand U8303 (N_8303,N_7852,N_7862);
or U8304 (N_8304,N_7911,N_7741);
nand U8305 (N_8305,N_7748,N_7652);
xnor U8306 (N_8306,N_7874,N_7906);
and U8307 (N_8307,N_7964,N_7570);
nand U8308 (N_8308,N_7750,N_7500);
nand U8309 (N_8309,N_7931,N_7791);
or U8310 (N_8310,N_7934,N_7705);
nand U8311 (N_8311,N_7515,N_7997);
xor U8312 (N_8312,N_7858,N_7615);
nand U8313 (N_8313,N_7719,N_7595);
nand U8314 (N_8314,N_7701,N_7921);
or U8315 (N_8315,N_7564,N_7654);
or U8316 (N_8316,N_7620,N_7600);
nand U8317 (N_8317,N_7558,N_7859);
xor U8318 (N_8318,N_7798,N_7681);
nor U8319 (N_8319,N_7967,N_7623);
and U8320 (N_8320,N_7944,N_7646);
nor U8321 (N_8321,N_7761,N_7989);
or U8322 (N_8322,N_7680,N_7561);
nand U8323 (N_8323,N_7954,N_7609);
nor U8324 (N_8324,N_7965,N_7705);
nand U8325 (N_8325,N_7723,N_7588);
xor U8326 (N_8326,N_7533,N_7792);
nand U8327 (N_8327,N_7862,N_7628);
xor U8328 (N_8328,N_7965,N_7856);
or U8329 (N_8329,N_7798,N_7744);
nand U8330 (N_8330,N_7814,N_7633);
nor U8331 (N_8331,N_7666,N_7831);
nor U8332 (N_8332,N_7594,N_7838);
xnor U8333 (N_8333,N_7980,N_7687);
nand U8334 (N_8334,N_7502,N_7947);
nor U8335 (N_8335,N_7842,N_7900);
or U8336 (N_8336,N_7691,N_7991);
or U8337 (N_8337,N_7943,N_7736);
or U8338 (N_8338,N_7510,N_7982);
and U8339 (N_8339,N_7648,N_7847);
xnor U8340 (N_8340,N_7676,N_7585);
xor U8341 (N_8341,N_7652,N_7510);
nor U8342 (N_8342,N_7862,N_7696);
or U8343 (N_8343,N_7736,N_7679);
nor U8344 (N_8344,N_7763,N_7533);
or U8345 (N_8345,N_7616,N_7906);
nor U8346 (N_8346,N_7630,N_7553);
nand U8347 (N_8347,N_7747,N_7570);
and U8348 (N_8348,N_7925,N_7698);
xor U8349 (N_8349,N_7533,N_7680);
or U8350 (N_8350,N_7557,N_7637);
nor U8351 (N_8351,N_7661,N_7910);
or U8352 (N_8352,N_7889,N_7548);
nor U8353 (N_8353,N_7953,N_7832);
and U8354 (N_8354,N_7999,N_7904);
and U8355 (N_8355,N_7784,N_7517);
and U8356 (N_8356,N_7822,N_7828);
or U8357 (N_8357,N_7547,N_7619);
and U8358 (N_8358,N_7849,N_7811);
or U8359 (N_8359,N_7779,N_7883);
nor U8360 (N_8360,N_7964,N_7839);
and U8361 (N_8361,N_7890,N_7748);
nor U8362 (N_8362,N_7978,N_7916);
xor U8363 (N_8363,N_7944,N_7986);
and U8364 (N_8364,N_7506,N_7971);
nor U8365 (N_8365,N_7658,N_7806);
and U8366 (N_8366,N_7798,N_7630);
nand U8367 (N_8367,N_7917,N_7927);
and U8368 (N_8368,N_7622,N_7877);
and U8369 (N_8369,N_7890,N_7835);
nand U8370 (N_8370,N_7531,N_7817);
nand U8371 (N_8371,N_7690,N_7556);
nor U8372 (N_8372,N_7931,N_7628);
nor U8373 (N_8373,N_7907,N_7638);
and U8374 (N_8374,N_7510,N_7552);
nor U8375 (N_8375,N_7813,N_7915);
xor U8376 (N_8376,N_7791,N_7608);
and U8377 (N_8377,N_7868,N_7510);
nor U8378 (N_8378,N_7686,N_7720);
xnor U8379 (N_8379,N_7744,N_7863);
nor U8380 (N_8380,N_7500,N_7603);
or U8381 (N_8381,N_7951,N_7919);
xnor U8382 (N_8382,N_7963,N_7551);
and U8383 (N_8383,N_7961,N_7513);
nor U8384 (N_8384,N_7899,N_7556);
nand U8385 (N_8385,N_7996,N_7673);
nand U8386 (N_8386,N_7545,N_7986);
xor U8387 (N_8387,N_7666,N_7552);
nand U8388 (N_8388,N_7639,N_7760);
xnor U8389 (N_8389,N_7637,N_7992);
nand U8390 (N_8390,N_7697,N_7965);
or U8391 (N_8391,N_7800,N_7747);
xnor U8392 (N_8392,N_7885,N_7940);
xnor U8393 (N_8393,N_7871,N_7801);
nor U8394 (N_8394,N_7530,N_7935);
and U8395 (N_8395,N_7561,N_7621);
and U8396 (N_8396,N_7583,N_7575);
nor U8397 (N_8397,N_7946,N_7709);
and U8398 (N_8398,N_7944,N_7796);
or U8399 (N_8399,N_7678,N_7512);
nor U8400 (N_8400,N_7840,N_7941);
nand U8401 (N_8401,N_7530,N_7541);
nand U8402 (N_8402,N_7667,N_7974);
nand U8403 (N_8403,N_7849,N_7594);
and U8404 (N_8404,N_7977,N_7729);
nand U8405 (N_8405,N_7646,N_7612);
nor U8406 (N_8406,N_7909,N_7795);
xor U8407 (N_8407,N_7565,N_7923);
or U8408 (N_8408,N_7860,N_7855);
nor U8409 (N_8409,N_7789,N_7723);
and U8410 (N_8410,N_7777,N_7795);
or U8411 (N_8411,N_7938,N_7959);
or U8412 (N_8412,N_7722,N_7816);
nor U8413 (N_8413,N_7663,N_7996);
nand U8414 (N_8414,N_7596,N_7694);
nor U8415 (N_8415,N_7722,N_7556);
nor U8416 (N_8416,N_7705,N_7998);
nor U8417 (N_8417,N_7986,N_7947);
nand U8418 (N_8418,N_7626,N_7944);
and U8419 (N_8419,N_7683,N_7760);
and U8420 (N_8420,N_7649,N_7893);
nand U8421 (N_8421,N_7579,N_7981);
xor U8422 (N_8422,N_7816,N_7760);
or U8423 (N_8423,N_7517,N_7729);
xor U8424 (N_8424,N_7708,N_7876);
and U8425 (N_8425,N_7941,N_7758);
nand U8426 (N_8426,N_7543,N_7823);
and U8427 (N_8427,N_7819,N_7962);
nand U8428 (N_8428,N_7922,N_7698);
xnor U8429 (N_8429,N_7779,N_7694);
nand U8430 (N_8430,N_7604,N_7852);
nor U8431 (N_8431,N_7753,N_7887);
nand U8432 (N_8432,N_7774,N_7712);
nand U8433 (N_8433,N_7894,N_7767);
and U8434 (N_8434,N_7884,N_7506);
nand U8435 (N_8435,N_7733,N_7646);
xor U8436 (N_8436,N_7564,N_7649);
or U8437 (N_8437,N_7837,N_7996);
or U8438 (N_8438,N_7726,N_7903);
nor U8439 (N_8439,N_7524,N_7918);
xnor U8440 (N_8440,N_7761,N_7525);
and U8441 (N_8441,N_7799,N_7982);
or U8442 (N_8442,N_7622,N_7748);
or U8443 (N_8443,N_7664,N_7673);
or U8444 (N_8444,N_7812,N_7531);
nand U8445 (N_8445,N_7813,N_7695);
xor U8446 (N_8446,N_7784,N_7549);
nor U8447 (N_8447,N_7849,N_7961);
xor U8448 (N_8448,N_7763,N_7893);
xor U8449 (N_8449,N_7934,N_7564);
and U8450 (N_8450,N_7814,N_7759);
nand U8451 (N_8451,N_7867,N_7577);
and U8452 (N_8452,N_7976,N_7646);
and U8453 (N_8453,N_7752,N_7561);
nand U8454 (N_8454,N_7961,N_7895);
nor U8455 (N_8455,N_7678,N_7704);
and U8456 (N_8456,N_7573,N_7770);
nand U8457 (N_8457,N_7975,N_7740);
xor U8458 (N_8458,N_7806,N_7736);
or U8459 (N_8459,N_7883,N_7533);
or U8460 (N_8460,N_7673,N_7501);
and U8461 (N_8461,N_7774,N_7665);
or U8462 (N_8462,N_7762,N_7626);
and U8463 (N_8463,N_7765,N_7747);
xnor U8464 (N_8464,N_7954,N_7989);
nand U8465 (N_8465,N_7597,N_7854);
and U8466 (N_8466,N_7961,N_7928);
and U8467 (N_8467,N_7867,N_7630);
nand U8468 (N_8468,N_7827,N_7837);
or U8469 (N_8469,N_7843,N_7706);
xnor U8470 (N_8470,N_7693,N_7773);
or U8471 (N_8471,N_7777,N_7990);
or U8472 (N_8472,N_7630,N_7655);
xor U8473 (N_8473,N_7775,N_7858);
nor U8474 (N_8474,N_7844,N_7513);
nand U8475 (N_8475,N_7721,N_7747);
nand U8476 (N_8476,N_7783,N_7599);
and U8477 (N_8477,N_7772,N_7690);
nand U8478 (N_8478,N_7641,N_7608);
xnor U8479 (N_8479,N_7625,N_7764);
or U8480 (N_8480,N_7560,N_7545);
xnor U8481 (N_8481,N_7817,N_7899);
nor U8482 (N_8482,N_7656,N_7879);
nand U8483 (N_8483,N_7850,N_7748);
nor U8484 (N_8484,N_7779,N_7846);
or U8485 (N_8485,N_7781,N_7702);
xor U8486 (N_8486,N_7898,N_7926);
xnor U8487 (N_8487,N_7638,N_7823);
or U8488 (N_8488,N_7540,N_7909);
nor U8489 (N_8489,N_7743,N_7842);
xor U8490 (N_8490,N_7505,N_7710);
and U8491 (N_8491,N_7549,N_7590);
xnor U8492 (N_8492,N_7716,N_7520);
nand U8493 (N_8493,N_7548,N_7969);
and U8494 (N_8494,N_7683,N_7839);
xor U8495 (N_8495,N_7905,N_7761);
nand U8496 (N_8496,N_7509,N_7506);
nand U8497 (N_8497,N_7763,N_7577);
or U8498 (N_8498,N_7913,N_7614);
or U8499 (N_8499,N_7605,N_7823);
or U8500 (N_8500,N_8104,N_8237);
nand U8501 (N_8501,N_8098,N_8396);
and U8502 (N_8502,N_8190,N_8319);
and U8503 (N_8503,N_8035,N_8217);
xnor U8504 (N_8504,N_8475,N_8373);
and U8505 (N_8505,N_8064,N_8078);
nor U8506 (N_8506,N_8378,N_8377);
nor U8507 (N_8507,N_8218,N_8052);
nand U8508 (N_8508,N_8390,N_8456);
nor U8509 (N_8509,N_8366,N_8438);
nor U8510 (N_8510,N_8461,N_8256);
nor U8511 (N_8511,N_8106,N_8315);
and U8512 (N_8512,N_8087,N_8358);
nand U8513 (N_8513,N_8299,N_8292);
and U8514 (N_8514,N_8150,N_8123);
or U8515 (N_8515,N_8092,N_8443);
nand U8516 (N_8516,N_8304,N_8155);
or U8517 (N_8517,N_8004,N_8447);
nand U8518 (N_8518,N_8355,N_8048);
nand U8519 (N_8519,N_8433,N_8327);
nor U8520 (N_8520,N_8334,N_8049);
xnor U8521 (N_8521,N_8259,N_8057);
nor U8522 (N_8522,N_8027,N_8129);
and U8523 (N_8523,N_8130,N_8338);
nor U8524 (N_8524,N_8464,N_8419);
xor U8525 (N_8525,N_8127,N_8308);
nor U8526 (N_8526,N_8229,N_8216);
nor U8527 (N_8527,N_8252,N_8287);
nand U8528 (N_8528,N_8008,N_8241);
nor U8529 (N_8529,N_8249,N_8303);
nand U8530 (N_8530,N_8069,N_8286);
nand U8531 (N_8531,N_8149,N_8487);
or U8532 (N_8532,N_8036,N_8339);
xor U8533 (N_8533,N_8430,N_8258);
and U8534 (N_8534,N_8455,N_8290);
and U8535 (N_8535,N_8289,N_8172);
nand U8536 (N_8536,N_8121,N_8265);
or U8537 (N_8537,N_8103,N_8264);
or U8538 (N_8538,N_8293,N_8174);
and U8539 (N_8539,N_8335,N_8016);
nand U8540 (N_8540,N_8126,N_8143);
nand U8541 (N_8541,N_8105,N_8146);
and U8542 (N_8542,N_8062,N_8240);
nor U8543 (N_8543,N_8221,N_8294);
xor U8544 (N_8544,N_8242,N_8496);
and U8545 (N_8545,N_8158,N_8090);
nand U8546 (N_8546,N_8117,N_8428);
and U8547 (N_8547,N_8326,N_8457);
and U8548 (N_8548,N_8368,N_8344);
and U8549 (N_8549,N_8023,N_8115);
or U8550 (N_8550,N_8009,N_8370);
and U8551 (N_8551,N_8454,N_8312);
or U8552 (N_8552,N_8097,N_8040);
nand U8553 (N_8553,N_8215,N_8450);
or U8554 (N_8554,N_8184,N_8107);
xnor U8555 (N_8555,N_8300,N_8236);
nor U8556 (N_8556,N_8230,N_8422);
xor U8557 (N_8557,N_8210,N_8360);
nor U8558 (N_8558,N_8266,N_8177);
or U8559 (N_8559,N_8141,N_8403);
nor U8560 (N_8560,N_8047,N_8369);
nor U8561 (N_8561,N_8188,N_8185);
xnor U8562 (N_8562,N_8269,N_8387);
nor U8563 (N_8563,N_8473,N_8257);
nand U8564 (N_8564,N_8192,N_8212);
and U8565 (N_8565,N_8099,N_8267);
and U8566 (N_8566,N_8271,N_8182);
nand U8567 (N_8567,N_8323,N_8291);
and U8568 (N_8568,N_8477,N_8043);
nor U8569 (N_8569,N_8284,N_8091);
xnor U8570 (N_8570,N_8166,N_8305);
nor U8571 (N_8571,N_8181,N_8262);
or U8572 (N_8572,N_8139,N_8371);
nand U8573 (N_8573,N_8239,N_8316);
nor U8574 (N_8574,N_8214,N_8353);
and U8575 (N_8575,N_8119,N_8154);
nor U8576 (N_8576,N_8122,N_8364);
nand U8577 (N_8577,N_8484,N_8152);
nor U8578 (N_8578,N_8356,N_8399);
xor U8579 (N_8579,N_8169,N_8045);
nor U8580 (N_8580,N_8025,N_8082);
nor U8581 (N_8581,N_8354,N_8317);
nor U8582 (N_8582,N_8398,N_8075);
or U8583 (N_8583,N_8320,N_8379);
or U8584 (N_8584,N_8272,N_8228);
nor U8585 (N_8585,N_8467,N_8163);
nor U8586 (N_8586,N_8111,N_8478);
xnor U8587 (N_8587,N_8383,N_8493);
and U8588 (N_8588,N_8005,N_8440);
nor U8589 (N_8589,N_8222,N_8298);
xnor U8590 (N_8590,N_8275,N_8248);
and U8591 (N_8591,N_8223,N_8088);
and U8592 (N_8592,N_8160,N_8365);
nand U8593 (N_8593,N_8101,N_8426);
nand U8594 (N_8594,N_8448,N_8451);
and U8595 (N_8595,N_8498,N_8311);
xor U8596 (N_8596,N_8157,N_8238);
or U8597 (N_8597,N_8072,N_8077);
or U8598 (N_8598,N_8019,N_8283);
nor U8599 (N_8599,N_8193,N_8226);
nor U8600 (N_8600,N_8296,N_8156);
nor U8601 (N_8601,N_8109,N_8034);
and U8602 (N_8602,N_8254,N_8110);
and U8603 (N_8603,N_8061,N_8246);
nor U8604 (N_8604,N_8322,N_8056);
xor U8605 (N_8605,N_8164,N_8011);
nor U8606 (N_8606,N_8260,N_8488);
xnor U8607 (N_8607,N_8471,N_8423);
or U8608 (N_8608,N_8279,N_8026);
and U8609 (N_8609,N_8499,N_8065);
or U8610 (N_8610,N_8268,N_8132);
or U8611 (N_8611,N_8205,N_8341);
or U8612 (N_8612,N_8147,N_8250);
nor U8613 (N_8613,N_8017,N_8060);
or U8614 (N_8614,N_8466,N_8452);
xor U8615 (N_8615,N_8395,N_8435);
xor U8616 (N_8616,N_8337,N_8000);
xor U8617 (N_8617,N_8243,N_8424);
or U8618 (N_8618,N_8118,N_8108);
or U8619 (N_8619,N_8384,N_8407);
or U8620 (N_8620,N_8083,N_8148);
xnor U8621 (N_8621,N_8191,N_8231);
or U8622 (N_8622,N_8436,N_8161);
nor U8623 (N_8623,N_8372,N_8028);
nand U8624 (N_8624,N_8142,N_8325);
nor U8625 (N_8625,N_8495,N_8458);
nor U8626 (N_8626,N_8136,N_8282);
nand U8627 (N_8627,N_8054,N_8389);
xnor U8628 (N_8628,N_8417,N_8225);
and U8629 (N_8629,N_8100,N_8168);
or U8630 (N_8630,N_8213,N_8336);
nand U8631 (N_8631,N_8491,N_8469);
or U8632 (N_8632,N_8261,N_8459);
nand U8633 (N_8633,N_8093,N_8081);
nand U8634 (N_8634,N_8202,N_8444);
nor U8635 (N_8635,N_8067,N_8402);
xnor U8636 (N_8636,N_8324,N_8410);
nand U8637 (N_8637,N_8055,N_8328);
or U8638 (N_8638,N_8421,N_8412);
and U8639 (N_8639,N_8489,N_8362);
and U8640 (N_8640,N_8196,N_8232);
xor U8641 (N_8641,N_8073,N_8183);
and U8642 (N_8642,N_8037,N_8363);
xor U8643 (N_8643,N_8058,N_8297);
xnor U8644 (N_8644,N_8434,N_8138);
xor U8645 (N_8645,N_8442,N_8010);
xor U8646 (N_8646,N_8413,N_8041);
nor U8647 (N_8647,N_8432,N_8197);
nor U8648 (N_8648,N_8050,N_8276);
xor U8649 (N_8649,N_8140,N_8361);
nand U8650 (N_8650,N_8391,N_8474);
xnor U8651 (N_8651,N_8176,N_8167);
and U8652 (N_8652,N_8032,N_8318);
or U8653 (N_8653,N_8219,N_8144);
nand U8654 (N_8654,N_8253,N_8033);
nor U8655 (N_8655,N_8018,N_8255);
nor U8656 (N_8656,N_8281,N_8482);
nand U8657 (N_8657,N_8408,N_8472);
nor U8658 (N_8658,N_8002,N_8483);
xnor U8659 (N_8659,N_8173,N_8089);
xnor U8660 (N_8660,N_8420,N_8234);
or U8661 (N_8661,N_8114,N_8351);
and U8662 (N_8662,N_8494,N_8427);
or U8663 (N_8663,N_8020,N_8051);
nor U8664 (N_8664,N_8381,N_8063);
nand U8665 (N_8665,N_8347,N_8367);
xnor U8666 (N_8666,N_8079,N_8352);
nor U8667 (N_8667,N_8480,N_8330);
nand U8668 (N_8668,N_8128,N_8302);
and U8669 (N_8669,N_8321,N_8343);
nor U8670 (N_8670,N_8388,N_8416);
and U8671 (N_8671,N_8080,N_8340);
or U8672 (N_8672,N_8171,N_8460);
or U8673 (N_8673,N_8096,N_8277);
or U8674 (N_8674,N_8007,N_8084);
or U8675 (N_8675,N_8178,N_8059);
or U8676 (N_8676,N_8431,N_8309);
nor U8677 (N_8677,N_8074,N_8314);
xor U8678 (N_8678,N_8235,N_8039);
or U8679 (N_8679,N_8208,N_8453);
nor U8680 (N_8680,N_8003,N_8001);
nor U8681 (N_8681,N_8263,N_8134);
or U8682 (N_8682,N_8200,N_8310);
or U8683 (N_8683,N_8313,N_8331);
nor U8684 (N_8684,N_8006,N_8245);
or U8685 (N_8685,N_8382,N_8463);
nor U8686 (N_8686,N_8301,N_8195);
nand U8687 (N_8687,N_8186,N_8125);
xnor U8688 (N_8688,N_8346,N_8042);
and U8689 (N_8689,N_8076,N_8247);
and U8690 (N_8690,N_8224,N_8179);
or U8691 (N_8691,N_8014,N_8405);
xnor U8692 (N_8692,N_8386,N_8068);
or U8693 (N_8693,N_8170,N_8029);
or U8694 (N_8694,N_8203,N_8220);
and U8695 (N_8695,N_8085,N_8165);
xnor U8696 (N_8696,N_8332,N_8449);
nand U8697 (N_8697,N_8359,N_8116);
nor U8698 (N_8698,N_8429,N_8492);
and U8699 (N_8699,N_8415,N_8206);
nor U8700 (N_8700,N_8465,N_8151);
nor U8701 (N_8701,N_8329,N_8476);
and U8702 (N_8702,N_8046,N_8095);
and U8703 (N_8703,N_8374,N_8044);
or U8704 (N_8704,N_8446,N_8112);
or U8705 (N_8705,N_8445,N_8401);
xnor U8706 (N_8706,N_8189,N_8133);
or U8707 (N_8707,N_8497,N_8350);
and U8708 (N_8708,N_8113,N_8479);
nor U8709 (N_8709,N_8333,N_8102);
and U8710 (N_8710,N_8071,N_8175);
or U8711 (N_8711,N_8066,N_8306);
xor U8712 (N_8712,N_8295,N_8012);
nor U8713 (N_8713,N_8024,N_8437);
or U8714 (N_8714,N_8481,N_8031);
nor U8715 (N_8715,N_8207,N_8038);
and U8716 (N_8716,N_8439,N_8021);
xnor U8717 (N_8717,N_8404,N_8270);
nand U8718 (N_8718,N_8385,N_8380);
and U8719 (N_8719,N_8227,N_8411);
xnor U8720 (N_8720,N_8274,N_8209);
or U8721 (N_8721,N_8486,N_8485);
or U8722 (N_8722,N_8376,N_8397);
or U8723 (N_8723,N_8120,N_8400);
xnor U8724 (N_8724,N_8392,N_8131);
or U8725 (N_8725,N_8375,N_8288);
xnor U8726 (N_8726,N_8345,N_8462);
nand U8727 (N_8727,N_8357,N_8280);
xor U8728 (N_8728,N_8251,N_8053);
nand U8729 (N_8729,N_8194,N_8285);
and U8730 (N_8730,N_8470,N_8137);
or U8731 (N_8731,N_8418,N_8393);
xnor U8732 (N_8732,N_8342,N_8425);
xor U8733 (N_8733,N_8409,N_8414);
nor U8734 (N_8734,N_8441,N_8468);
xnor U8735 (N_8735,N_8013,N_8030);
nand U8736 (N_8736,N_8394,N_8348);
nor U8737 (N_8737,N_8406,N_8145);
xor U8738 (N_8738,N_8187,N_8233);
and U8739 (N_8739,N_8198,N_8273);
or U8740 (N_8740,N_8201,N_8159);
nand U8741 (N_8741,N_8135,N_8015);
nor U8742 (N_8742,N_8204,N_8086);
nor U8743 (N_8743,N_8349,N_8199);
or U8744 (N_8744,N_8180,N_8124);
xor U8745 (N_8745,N_8490,N_8094);
nor U8746 (N_8746,N_8162,N_8278);
nand U8747 (N_8747,N_8307,N_8244);
or U8748 (N_8748,N_8070,N_8022);
nor U8749 (N_8749,N_8153,N_8211);
xor U8750 (N_8750,N_8401,N_8324);
or U8751 (N_8751,N_8130,N_8452);
and U8752 (N_8752,N_8087,N_8075);
xor U8753 (N_8753,N_8431,N_8013);
xnor U8754 (N_8754,N_8141,N_8242);
nor U8755 (N_8755,N_8164,N_8321);
or U8756 (N_8756,N_8138,N_8393);
and U8757 (N_8757,N_8156,N_8108);
xnor U8758 (N_8758,N_8219,N_8074);
and U8759 (N_8759,N_8115,N_8439);
or U8760 (N_8760,N_8396,N_8485);
or U8761 (N_8761,N_8040,N_8248);
nand U8762 (N_8762,N_8286,N_8042);
nor U8763 (N_8763,N_8278,N_8011);
or U8764 (N_8764,N_8234,N_8071);
and U8765 (N_8765,N_8170,N_8346);
nor U8766 (N_8766,N_8236,N_8175);
or U8767 (N_8767,N_8413,N_8288);
or U8768 (N_8768,N_8364,N_8169);
nand U8769 (N_8769,N_8486,N_8137);
nor U8770 (N_8770,N_8199,N_8289);
nor U8771 (N_8771,N_8378,N_8371);
and U8772 (N_8772,N_8394,N_8441);
xor U8773 (N_8773,N_8033,N_8199);
nand U8774 (N_8774,N_8417,N_8384);
xor U8775 (N_8775,N_8292,N_8210);
xnor U8776 (N_8776,N_8411,N_8255);
xnor U8777 (N_8777,N_8479,N_8119);
xor U8778 (N_8778,N_8169,N_8043);
or U8779 (N_8779,N_8062,N_8087);
nor U8780 (N_8780,N_8485,N_8298);
or U8781 (N_8781,N_8020,N_8089);
nand U8782 (N_8782,N_8250,N_8412);
nand U8783 (N_8783,N_8130,N_8461);
nand U8784 (N_8784,N_8465,N_8051);
and U8785 (N_8785,N_8410,N_8128);
or U8786 (N_8786,N_8498,N_8128);
nand U8787 (N_8787,N_8144,N_8121);
or U8788 (N_8788,N_8395,N_8331);
xnor U8789 (N_8789,N_8485,N_8083);
and U8790 (N_8790,N_8136,N_8083);
or U8791 (N_8791,N_8304,N_8461);
or U8792 (N_8792,N_8139,N_8088);
and U8793 (N_8793,N_8065,N_8350);
nor U8794 (N_8794,N_8396,N_8455);
nor U8795 (N_8795,N_8409,N_8271);
or U8796 (N_8796,N_8143,N_8048);
nand U8797 (N_8797,N_8409,N_8295);
and U8798 (N_8798,N_8490,N_8062);
nand U8799 (N_8799,N_8070,N_8000);
nand U8800 (N_8800,N_8189,N_8482);
nand U8801 (N_8801,N_8058,N_8445);
xnor U8802 (N_8802,N_8064,N_8399);
nand U8803 (N_8803,N_8134,N_8078);
or U8804 (N_8804,N_8384,N_8252);
nand U8805 (N_8805,N_8076,N_8263);
and U8806 (N_8806,N_8381,N_8069);
or U8807 (N_8807,N_8143,N_8364);
nand U8808 (N_8808,N_8088,N_8195);
xnor U8809 (N_8809,N_8042,N_8071);
and U8810 (N_8810,N_8010,N_8229);
and U8811 (N_8811,N_8140,N_8004);
xor U8812 (N_8812,N_8335,N_8286);
and U8813 (N_8813,N_8331,N_8069);
xnor U8814 (N_8814,N_8377,N_8043);
and U8815 (N_8815,N_8459,N_8417);
or U8816 (N_8816,N_8084,N_8400);
and U8817 (N_8817,N_8047,N_8173);
or U8818 (N_8818,N_8351,N_8060);
or U8819 (N_8819,N_8345,N_8174);
or U8820 (N_8820,N_8054,N_8082);
and U8821 (N_8821,N_8156,N_8239);
or U8822 (N_8822,N_8009,N_8077);
nor U8823 (N_8823,N_8135,N_8487);
nor U8824 (N_8824,N_8209,N_8342);
nand U8825 (N_8825,N_8147,N_8299);
and U8826 (N_8826,N_8299,N_8273);
nand U8827 (N_8827,N_8052,N_8272);
and U8828 (N_8828,N_8220,N_8044);
or U8829 (N_8829,N_8478,N_8444);
and U8830 (N_8830,N_8452,N_8460);
and U8831 (N_8831,N_8453,N_8385);
nor U8832 (N_8832,N_8239,N_8383);
nor U8833 (N_8833,N_8023,N_8258);
nand U8834 (N_8834,N_8360,N_8135);
nand U8835 (N_8835,N_8458,N_8008);
nand U8836 (N_8836,N_8483,N_8348);
xnor U8837 (N_8837,N_8133,N_8173);
nand U8838 (N_8838,N_8274,N_8260);
nand U8839 (N_8839,N_8128,N_8049);
nand U8840 (N_8840,N_8296,N_8100);
and U8841 (N_8841,N_8263,N_8398);
nand U8842 (N_8842,N_8178,N_8305);
nand U8843 (N_8843,N_8116,N_8132);
or U8844 (N_8844,N_8247,N_8394);
and U8845 (N_8845,N_8477,N_8394);
or U8846 (N_8846,N_8402,N_8411);
and U8847 (N_8847,N_8304,N_8121);
xor U8848 (N_8848,N_8401,N_8307);
xor U8849 (N_8849,N_8162,N_8024);
nor U8850 (N_8850,N_8204,N_8368);
nand U8851 (N_8851,N_8012,N_8142);
or U8852 (N_8852,N_8170,N_8466);
xnor U8853 (N_8853,N_8433,N_8271);
nand U8854 (N_8854,N_8409,N_8258);
or U8855 (N_8855,N_8142,N_8191);
nand U8856 (N_8856,N_8265,N_8489);
xor U8857 (N_8857,N_8443,N_8221);
and U8858 (N_8858,N_8267,N_8178);
and U8859 (N_8859,N_8219,N_8067);
nand U8860 (N_8860,N_8136,N_8284);
nand U8861 (N_8861,N_8010,N_8041);
xnor U8862 (N_8862,N_8141,N_8248);
nor U8863 (N_8863,N_8048,N_8284);
xnor U8864 (N_8864,N_8044,N_8284);
or U8865 (N_8865,N_8180,N_8198);
or U8866 (N_8866,N_8157,N_8141);
xor U8867 (N_8867,N_8196,N_8433);
xnor U8868 (N_8868,N_8422,N_8410);
xnor U8869 (N_8869,N_8152,N_8446);
or U8870 (N_8870,N_8166,N_8369);
and U8871 (N_8871,N_8480,N_8173);
and U8872 (N_8872,N_8351,N_8184);
nand U8873 (N_8873,N_8143,N_8386);
and U8874 (N_8874,N_8200,N_8124);
nand U8875 (N_8875,N_8405,N_8001);
and U8876 (N_8876,N_8327,N_8089);
and U8877 (N_8877,N_8036,N_8319);
and U8878 (N_8878,N_8297,N_8152);
and U8879 (N_8879,N_8011,N_8230);
or U8880 (N_8880,N_8067,N_8024);
and U8881 (N_8881,N_8005,N_8091);
xnor U8882 (N_8882,N_8011,N_8163);
nand U8883 (N_8883,N_8019,N_8499);
xor U8884 (N_8884,N_8260,N_8400);
nand U8885 (N_8885,N_8366,N_8187);
xor U8886 (N_8886,N_8267,N_8137);
nor U8887 (N_8887,N_8491,N_8161);
xnor U8888 (N_8888,N_8488,N_8180);
xnor U8889 (N_8889,N_8216,N_8088);
nor U8890 (N_8890,N_8195,N_8314);
or U8891 (N_8891,N_8496,N_8051);
and U8892 (N_8892,N_8293,N_8357);
nand U8893 (N_8893,N_8424,N_8094);
or U8894 (N_8894,N_8201,N_8278);
nand U8895 (N_8895,N_8277,N_8016);
nor U8896 (N_8896,N_8014,N_8323);
or U8897 (N_8897,N_8384,N_8382);
or U8898 (N_8898,N_8098,N_8131);
nand U8899 (N_8899,N_8433,N_8376);
or U8900 (N_8900,N_8037,N_8256);
xnor U8901 (N_8901,N_8377,N_8097);
nor U8902 (N_8902,N_8273,N_8424);
or U8903 (N_8903,N_8097,N_8010);
nand U8904 (N_8904,N_8019,N_8062);
nand U8905 (N_8905,N_8356,N_8165);
nor U8906 (N_8906,N_8025,N_8193);
xor U8907 (N_8907,N_8339,N_8418);
and U8908 (N_8908,N_8022,N_8092);
nand U8909 (N_8909,N_8415,N_8161);
xnor U8910 (N_8910,N_8409,N_8084);
nor U8911 (N_8911,N_8323,N_8090);
xnor U8912 (N_8912,N_8419,N_8122);
nand U8913 (N_8913,N_8387,N_8161);
or U8914 (N_8914,N_8089,N_8085);
and U8915 (N_8915,N_8258,N_8135);
and U8916 (N_8916,N_8245,N_8269);
xnor U8917 (N_8917,N_8374,N_8187);
nor U8918 (N_8918,N_8325,N_8178);
xnor U8919 (N_8919,N_8248,N_8266);
or U8920 (N_8920,N_8091,N_8453);
nand U8921 (N_8921,N_8364,N_8145);
xor U8922 (N_8922,N_8027,N_8223);
and U8923 (N_8923,N_8233,N_8033);
xor U8924 (N_8924,N_8266,N_8016);
or U8925 (N_8925,N_8462,N_8246);
or U8926 (N_8926,N_8447,N_8255);
xnor U8927 (N_8927,N_8387,N_8147);
xor U8928 (N_8928,N_8404,N_8136);
nand U8929 (N_8929,N_8399,N_8324);
xnor U8930 (N_8930,N_8011,N_8369);
nor U8931 (N_8931,N_8476,N_8496);
or U8932 (N_8932,N_8062,N_8039);
and U8933 (N_8933,N_8204,N_8212);
nand U8934 (N_8934,N_8212,N_8074);
xor U8935 (N_8935,N_8305,N_8268);
xnor U8936 (N_8936,N_8182,N_8368);
nand U8937 (N_8937,N_8496,N_8224);
and U8938 (N_8938,N_8420,N_8149);
xnor U8939 (N_8939,N_8471,N_8079);
nand U8940 (N_8940,N_8118,N_8491);
nand U8941 (N_8941,N_8129,N_8174);
and U8942 (N_8942,N_8184,N_8181);
nand U8943 (N_8943,N_8347,N_8411);
or U8944 (N_8944,N_8473,N_8047);
nand U8945 (N_8945,N_8015,N_8445);
nand U8946 (N_8946,N_8000,N_8181);
nor U8947 (N_8947,N_8073,N_8482);
nor U8948 (N_8948,N_8027,N_8387);
xnor U8949 (N_8949,N_8235,N_8180);
nor U8950 (N_8950,N_8432,N_8226);
nor U8951 (N_8951,N_8018,N_8412);
xor U8952 (N_8952,N_8026,N_8289);
or U8953 (N_8953,N_8373,N_8200);
xor U8954 (N_8954,N_8205,N_8393);
and U8955 (N_8955,N_8233,N_8111);
xnor U8956 (N_8956,N_8198,N_8335);
or U8957 (N_8957,N_8457,N_8467);
xnor U8958 (N_8958,N_8260,N_8106);
xnor U8959 (N_8959,N_8186,N_8037);
xnor U8960 (N_8960,N_8378,N_8242);
or U8961 (N_8961,N_8474,N_8479);
nor U8962 (N_8962,N_8070,N_8191);
nand U8963 (N_8963,N_8006,N_8296);
or U8964 (N_8964,N_8438,N_8307);
nand U8965 (N_8965,N_8113,N_8494);
nand U8966 (N_8966,N_8147,N_8253);
nor U8967 (N_8967,N_8224,N_8280);
or U8968 (N_8968,N_8194,N_8036);
nand U8969 (N_8969,N_8049,N_8316);
nor U8970 (N_8970,N_8086,N_8092);
nor U8971 (N_8971,N_8139,N_8137);
or U8972 (N_8972,N_8330,N_8438);
xnor U8973 (N_8973,N_8140,N_8092);
or U8974 (N_8974,N_8159,N_8186);
nand U8975 (N_8975,N_8390,N_8426);
nor U8976 (N_8976,N_8037,N_8208);
nor U8977 (N_8977,N_8384,N_8243);
or U8978 (N_8978,N_8458,N_8071);
xor U8979 (N_8979,N_8206,N_8089);
or U8980 (N_8980,N_8007,N_8299);
nand U8981 (N_8981,N_8123,N_8327);
and U8982 (N_8982,N_8249,N_8243);
and U8983 (N_8983,N_8294,N_8058);
nor U8984 (N_8984,N_8012,N_8086);
and U8985 (N_8985,N_8014,N_8126);
xor U8986 (N_8986,N_8384,N_8242);
xnor U8987 (N_8987,N_8296,N_8354);
xnor U8988 (N_8988,N_8449,N_8499);
xnor U8989 (N_8989,N_8022,N_8491);
nor U8990 (N_8990,N_8298,N_8137);
xnor U8991 (N_8991,N_8458,N_8436);
nand U8992 (N_8992,N_8291,N_8069);
and U8993 (N_8993,N_8100,N_8379);
and U8994 (N_8994,N_8469,N_8166);
nand U8995 (N_8995,N_8192,N_8320);
and U8996 (N_8996,N_8175,N_8336);
nand U8997 (N_8997,N_8419,N_8305);
nor U8998 (N_8998,N_8251,N_8191);
and U8999 (N_8999,N_8067,N_8365);
nand U9000 (N_9000,N_8515,N_8717);
or U9001 (N_9001,N_8520,N_8591);
and U9002 (N_9002,N_8748,N_8756);
nand U9003 (N_9003,N_8995,N_8564);
xnor U9004 (N_9004,N_8736,N_8543);
xor U9005 (N_9005,N_8858,N_8853);
or U9006 (N_9006,N_8801,N_8529);
xnor U9007 (N_9007,N_8873,N_8811);
and U9008 (N_9008,N_8940,N_8552);
and U9009 (N_9009,N_8592,N_8677);
nand U9010 (N_9010,N_8810,N_8542);
or U9011 (N_9011,N_8854,N_8663);
nand U9012 (N_9012,N_8944,N_8720);
xor U9013 (N_9013,N_8544,N_8759);
nand U9014 (N_9014,N_8583,N_8766);
nor U9015 (N_9015,N_8604,N_8704);
nor U9016 (N_9016,N_8749,N_8540);
and U9017 (N_9017,N_8545,N_8934);
and U9018 (N_9018,N_8897,N_8670);
and U9019 (N_9019,N_8613,N_8723);
nor U9020 (N_9020,N_8728,N_8951);
xnor U9021 (N_9021,N_8846,N_8697);
xnor U9022 (N_9022,N_8595,N_8538);
nor U9023 (N_9023,N_8968,N_8903);
and U9024 (N_9024,N_8913,N_8554);
nor U9025 (N_9025,N_8840,N_8737);
nor U9026 (N_9026,N_8949,N_8767);
xnor U9027 (N_9027,N_8816,N_8547);
nand U9028 (N_9028,N_8505,N_8539);
nand U9029 (N_9029,N_8946,N_8974);
xnor U9030 (N_9030,N_8805,N_8863);
nand U9031 (N_9031,N_8660,N_8667);
xor U9032 (N_9032,N_8878,N_8651);
and U9033 (N_9033,N_8513,N_8841);
nand U9034 (N_9034,N_8718,N_8608);
or U9035 (N_9035,N_8981,N_8632);
nor U9036 (N_9036,N_8813,N_8674);
nand U9037 (N_9037,N_8626,N_8711);
and U9038 (N_9038,N_8818,N_8644);
or U9039 (N_9039,N_8987,N_8790);
or U9040 (N_9040,N_8933,N_8762);
xor U9041 (N_9041,N_8834,N_8923);
nand U9042 (N_9042,N_8849,N_8957);
xnor U9043 (N_9043,N_8652,N_8610);
or U9044 (N_9044,N_8500,N_8628);
nor U9045 (N_9045,N_8605,N_8734);
nand U9046 (N_9046,N_8796,N_8585);
nor U9047 (N_9047,N_8931,N_8916);
nand U9048 (N_9048,N_8708,N_8765);
nor U9049 (N_9049,N_8690,N_8795);
xnor U9050 (N_9050,N_8636,N_8941);
xnor U9051 (N_9051,N_8984,N_8550);
or U9052 (N_9052,N_8568,N_8825);
or U9053 (N_9053,N_8609,N_8694);
nand U9054 (N_9054,N_8990,N_8577);
xnor U9055 (N_9055,N_8800,N_8565);
nand U9056 (N_9056,N_8950,N_8623);
xnor U9057 (N_9057,N_8537,N_8803);
xnor U9058 (N_9058,N_8664,N_8955);
or U9059 (N_9059,N_8893,N_8735);
or U9060 (N_9060,N_8860,N_8647);
and U9061 (N_9061,N_8606,N_8689);
nand U9062 (N_9062,N_8861,N_8641);
or U9063 (N_9063,N_8837,N_8721);
xor U9064 (N_9064,N_8649,N_8738);
nand U9065 (N_9065,N_8832,N_8902);
nor U9066 (N_9066,N_8774,N_8502);
nor U9067 (N_9067,N_8822,N_8959);
xnor U9068 (N_9068,N_8899,N_8522);
or U9069 (N_9069,N_8914,N_8943);
or U9070 (N_9070,N_8619,N_8926);
or U9071 (N_9071,N_8730,N_8905);
nor U9072 (N_9072,N_8952,N_8947);
xor U9073 (N_9073,N_8971,N_8625);
xnor U9074 (N_9074,N_8722,N_8732);
and U9075 (N_9075,N_8920,N_8885);
or U9076 (N_9076,N_8586,N_8703);
xor U9077 (N_9077,N_8872,N_8999);
nor U9078 (N_9078,N_8699,N_8904);
nor U9079 (N_9079,N_8668,N_8692);
xor U9080 (N_9080,N_8615,N_8646);
or U9081 (N_9081,N_8534,N_8526);
nor U9082 (N_9082,N_8870,N_8880);
nand U9083 (N_9083,N_8714,N_8935);
nand U9084 (N_9084,N_8693,N_8638);
or U9085 (N_9085,N_8953,N_8620);
or U9086 (N_9086,N_8852,N_8763);
or U9087 (N_9087,N_8927,N_8700);
nor U9088 (N_9088,N_8936,N_8998);
nor U9089 (N_9089,N_8910,N_8921);
nor U9090 (N_9090,N_8603,N_8976);
xor U9091 (N_9091,N_8525,N_8826);
or U9092 (N_9092,N_8973,N_8675);
and U9093 (N_9093,N_8876,N_8574);
or U9094 (N_9094,N_8843,N_8584);
and U9095 (N_9095,N_8895,N_8977);
or U9096 (N_9096,N_8508,N_8573);
and U9097 (N_9097,N_8922,N_8869);
xnor U9098 (N_9098,N_8633,N_8889);
or U9099 (N_9099,N_8909,N_8798);
and U9100 (N_9100,N_8563,N_8655);
nand U9101 (N_9101,N_8958,N_8888);
xnor U9102 (N_9102,N_8978,N_8676);
nand U9103 (N_9103,N_8925,N_8965);
xnor U9104 (N_9104,N_8740,N_8776);
nand U9105 (N_9105,N_8601,N_8530);
nand U9106 (N_9106,N_8682,N_8580);
xor U9107 (N_9107,N_8960,N_8553);
xor U9108 (N_9108,N_8919,N_8746);
xor U9109 (N_9109,N_8777,N_8764);
xnor U9110 (N_9110,N_8627,N_8611);
nor U9111 (N_9111,N_8679,N_8572);
and U9112 (N_9112,N_8653,N_8862);
or U9113 (N_9113,N_8836,N_8607);
or U9114 (N_9114,N_8648,N_8982);
nor U9115 (N_9115,N_8928,N_8596);
xor U9116 (N_9116,N_8614,N_8719);
nor U9117 (N_9117,N_8794,N_8569);
and U9118 (N_9118,N_8503,N_8850);
or U9119 (N_9119,N_8900,N_8937);
xor U9120 (N_9120,N_8656,N_8890);
nor U9121 (N_9121,N_8879,N_8710);
nor U9122 (N_9122,N_8908,N_8932);
or U9123 (N_9123,N_8597,N_8793);
or U9124 (N_9124,N_8906,N_8709);
nand U9125 (N_9125,N_8696,N_8779);
and U9126 (N_9126,N_8823,N_8678);
nand U9127 (N_9127,N_8686,N_8961);
and U9128 (N_9128,N_8504,N_8851);
or U9129 (N_9129,N_8871,N_8802);
nand U9130 (N_9130,N_8594,N_8966);
xor U9131 (N_9131,N_8575,N_8929);
or U9132 (N_9132,N_8657,N_8831);
nor U9133 (N_9133,N_8681,N_8556);
and U9134 (N_9134,N_8833,N_8555);
xnor U9135 (N_9135,N_8877,N_8654);
and U9136 (N_9136,N_8570,N_8804);
or U9137 (N_9137,N_8988,N_8726);
and U9138 (N_9138,N_8839,N_8698);
nand U9139 (N_9139,N_8635,N_8578);
and U9140 (N_9140,N_8784,N_8775);
nand U9141 (N_9141,N_8848,N_8874);
nand U9142 (N_9142,N_8770,N_8857);
or U9143 (N_9143,N_8758,N_8993);
xnor U9144 (N_9144,N_8817,N_8750);
xnor U9145 (N_9145,N_8600,N_8673);
or U9146 (N_9146,N_8602,N_8662);
and U9147 (N_9147,N_8989,N_8742);
and U9148 (N_9148,N_8842,N_8576);
xor U9149 (N_9149,N_8789,N_8518);
nand U9150 (N_9150,N_8745,N_8512);
or U9151 (N_9151,N_8938,N_8821);
nand U9152 (N_9152,N_8808,N_8685);
and U9153 (N_9153,N_8669,N_8886);
xnor U9154 (N_9154,N_8561,N_8942);
and U9155 (N_9155,N_8992,N_8658);
or U9156 (N_9156,N_8672,N_8918);
or U9157 (N_9157,N_8524,N_8593);
nor U9158 (N_9158,N_8954,N_8680);
or U9159 (N_9159,N_8743,N_8713);
nor U9160 (N_9160,N_8812,N_8637);
and U9161 (N_9161,N_8797,N_8536);
xor U9162 (N_9162,N_8744,N_8773);
xnor U9163 (N_9163,N_8924,N_8639);
or U9164 (N_9164,N_8519,N_8769);
nor U9165 (N_9165,N_8754,N_8780);
nand U9166 (N_9166,N_8571,N_8621);
and U9167 (N_9167,N_8566,N_8969);
nor U9168 (N_9168,N_8671,N_8791);
or U9169 (N_9169,N_8716,N_8650);
or U9170 (N_9170,N_8781,N_8807);
nor U9171 (N_9171,N_8972,N_8645);
xnor U9172 (N_9172,N_8859,N_8772);
xor U9173 (N_9173,N_8891,N_8617);
nor U9174 (N_9174,N_8917,N_8514);
or U9175 (N_9175,N_8741,N_8975);
xnor U9176 (N_9176,N_8867,N_8847);
nand U9177 (N_9177,N_8962,N_8531);
and U9178 (N_9178,N_8588,N_8546);
nand U9179 (N_9179,N_8541,N_8579);
nor U9180 (N_9180,N_8630,N_8548);
nand U9181 (N_9181,N_8629,N_8752);
or U9182 (N_9182,N_8640,N_8901);
xnor U9183 (N_9183,N_8631,N_8830);
and U9184 (N_9184,N_8930,N_8915);
xor U9185 (N_9185,N_8517,N_8815);
nand U9186 (N_9186,N_8963,N_8567);
or U9187 (N_9187,N_8523,N_8875);
xor U9188 (N_9188,N_8991,N_8911);
or U9189 (N_9189,N_8727,N_8533);
and U9190 (N_9190,N_8970,N_8760);
and U9191 (N_9191,N_8562,N_8516);
nor U9192 (N_9192,N_8828,N_8997);
or U9193 (N_9193,N_8509,N_8856);
xor U9194 (N_9194,N_8755,N_8898);
nor U9195 (N_9195,N_8616,N_8896);
and U9196 (N_9196,N_8783,N_8642);
xor U9197 (N_9197,N_8824,N_8715);
xnor U9198 (N_9198,N_8835,N_8753);
nor U9199 (N_9199,N_8598,N_8590);
and U9200 (N_9200,N_8844,N_8587);
and U9201 (N_9201,N_8507,N_8884);
nor U9202 (N_9202,N_8612,N_8622);
nand U9203 (N_9203,N_8751,N_8739);
and U9204 (N_9204,N_8551,N_8712);
nand U9205 (N_9205,N_8820,N_8799);
or U9206 (N_9206,N_8864,N_8892);
nand U9207 (N_9207,N_8589,N_8964);
and U9208 (N_9208,N_8829,N_8643);
or U9209 (N_9209,N_8560,N_8691);
xor U9210 (N_9210,N_8986,N_8707);
nand U9211 (N_9211,N_8939,N_8967);
xnor U9212 (N_9212,N_8535,N_8788);
nor U9213 (N_9213,N_8532,N_8894);
xnor U9214 (N_9214,N_8666,N_8787);
xnor U9215 (N_9215,N_8865,N_8702);
and U9216 (N_9216,N_8948,N_8582);
nand U9217 (N_9217,N_8725,N_8527);
or U9218 (N_9218,N_8729,N_8511);
or U9219 (N_9219,N_8785,N_8747);
xor U9220 (N_9220,N_8809,N_8731);
or U9221 (N_9221,N_8855,N_8684);
and U9222 (N_9222,N_8687,N_8501);
nor U9223 (N_9223,N_8706,N_8701);
and U9224 (N_9224,N_8506,N_8806);
and U9225 (N_9225,N_8881,N_8665);
nor U9226 (N_9226,N_8979,N_8634);
xor U9227 (N_9227,N_8771,N_8945);
xor U9228 (N_9228,N_8549,N_8761);
or U9229 (N_9229,N_8778,N_8782);
nand U9230 (N_9230,N_8528,N_8883);
xor U9231 (N_9231,N_8827,N_8599);
xnor U9232 (N_9232,N_8866,N_8996);
or U9233 (N_9233,N_8956,N_8882);
and U9234 (N_9234,N_8819,N_8558);
nor U9235 (N_9235,N_8983,N_8994);
xor U9236 (N_9236,N_8559,N_8624);
nand U9237 (N_9237,N_8695,N_8768);
or U9238 (N_9238,N_8912,N_8618);
xor U9239 (N_9239,N_8814,N_8683);
nor U9240 (N_9240,N_8980,N_8659);
or U9241 (N_9241,N_8521,N_8845);
or U9242 (N_9242,N_8838,N_8705);
nor U9243 (N_9243,N_8557,N_8907);
and U9244 (N_9244,N_8724,N_8661);
and U9245 (N_9245,N_8887,N_8786);
nor U9246 (N_9246,N_8688,N_8985);
nor U9247 (N_9247,N_8510,N_8757);
or U9248 (N_9248,N_8733,N_8868);
and U9249 (N_9249,N_8792,N_8581);
or U9250 (N_9250,N_8773,N_8622);
and U9251 (N_9251,N_8690,N_8671);
nand U9252 (N_9252,N_8988,N_8930);
or U9253 (N_9253,N_8974,N_8894);
or U9254 (N_9254,N_8908,N_8737);
xor U9255 (N_9255,N_8795,N_8706);
and U9256 (N_9256,N_8804,N_8708);
or U9257 (N_9257,N_8847,N_8994);
nand U9258 (N_9258,N_8545,N_8685);
nor U9259 (N_9259,N_8821,N_8750);
and U9260 (N_9260,N_8994,N_8567);
nor U9261 (N_9261,N_8705,N_8750);
and U9262 (N_9262,N_8980,N_8933);
xnor U9263 (N_9263,N_8916,N_8602);
nor U9264 (N_9264,N_8664,N_8591);
nor U9265 (N_9265,N_8792,N_8935);
nor U9266 (N_9266,N_8997,N_8807);
nand U9267 (N_9267,N_8511,N_8864);
or U9268 (N_9268,N_8876,N_8726);
or U9269 (N_9269,N_8996,N_8652);
nor U9270 (N_9270,N_8780,N_8849);
xor U9271 (N_9271,N_8961,N_8551);
or U9272 (N_9272,N_8695,N_8621);
xor U9273 (N_9273,N_8747,N_8844);
nor U9274 (N_9274,N_8779,N_8590);
nand U9275 (N_9275,N_8933,N_8834);
and U9276 (N_9276,N_8841,N_8709);
xnor U9277 (N_9277,N_8522,N_8864);
and U9278 (N_9278,N_8918,N_8929);
nand U9279 (N_9279,N_8857,N_8758);
and U9280 (N_9280,N_8511,N_8589);
and U9281 (N_9281,N_8504,N_8956);
and U9282 (N_9282,N_8845,N_8981);
xnor U9283 (N_9283,N_8713,N_8817);
and U9284 (N_9284,N_8796,N_8739);
and U9285 (N_9285,N_8747,N_8880);
or U9286 (N_9286,N_8806,N_8790);
and U9287 (N_9287,N_8781,N_8557);
nand U9288 (N_9288,N_8541,N_8789);
nand U9289 (N_9289,N_8777,N_8851);
nor U9290 (N_9290,N_8713,N_8825);
or U9291 (N_9291,N_8566,N_8751);
xnor U9292 (N_9292,N_8785,N_8859);
or U9293 (N_9293,N_8634,N_8735);
or U9294 (N_9294,N_8728,N_8642);
and U9295 (N_9295,N_8502,N_8925);
xnor U9296 (N_9296,N_8574,N_8817);
nor U9297 (N_9297,N_8961,N_8944);
nand U9298 (N_9298,N_8702,N_8614);
or U9299 (N_9299,N_8593,N_8979);
and U9300 (N_9300,N_8575,N_8674);
nor U9301 (N_9301,N_8742,N_8563);
and U9302 (N_9302,N_8723,N_8841);
nand U9303 (N_9303,N_8704,N_8535);
nand U9304 (N_9304,N_8591,N_8547);
nand U9305 (N_9305,N_8912,N_8993);
nand U9306 (N_9306,N_8937,N_8707);
nor U9307 (N_9307,N_8718,N_8604);
xor U9308 (N_9308,N_8795,N_8972);
or U9309 (N_9309,N_8771,N_8943);
or U9310 (N_9310,N_8704,N_8758);
nand U9311 (N_9311,N_8923,N_8505);
nor U9312 (N_9312,N_8503,N_8654);
nor U9313 (N_9313,N_8947,N_8679);
or U9314 (N_9314,N_8630,N_8622);
nor U9315 (N_9315,N_8881,N_8875);
nor U9316 (N_9316,N_8882,N_8850);
nand U9317 (N_9317,N_8686,N_8996);
and U9318 (N_9318,N_8790,N_8971);
or U9319 (N_9319,N_8743,N_8615);
nand U9320 (N_9320,N_8587,N_8607);
or U9321 (N_9321,N_8868,N_8813);
xnor U9322 (N_9322,N_8651,N_8688);
or U9323 (N_9323,N_8737,N_8571);
or U9324 (N_9324,N_8536,N_8978);
xnor U9325 (N_9325,N_8748,N_8738);
xor U9326 (N_9326,N_8697,N_8555);
or U9327 (N_9327,N_8717,N_8639);
or U9328 (N_9328,N_8771,N_8608);
nor U9329 (N_9329,N_8964,N_8846);
and U9330 (N_9330,N_8925,N_8501);
nor U9331 (N_9331,N_8611,N_8634);
nor U9332 (N_9332,N_8543,N_8585);
nand U9333 (N_9333,N_8798,N_8971);
nor U9334 (N_9334,N_8958,N_8800);
and U9335 (N_9335,N_8896,N_8803);
and U9336 (N_9336,N_8559,N_8833);
xnor U9337 (N_9337,N_8902,N_8812);
and U9338 (N_9338,N_8617,N_8558);
and U9339 (N_9339,N_8659,N_8901);
or U9340 (N_9340,N_8878,N_8697);
nor U9341 (N_9341,N_8940,N_8559);
or U9342 (N_9342,N_8545,N_8906);
nand U9343 (N_9343,N_8982,N_8742);
and U9344 (N_9344,N_8521,N_8784);
nor U9345 (N_9345,N_8872,N_8767);
nor U9346 (N_9346,N_8767,N_8799);
or U9347 (N_9347,N_8677,N_8630);
or U9348 (N_9348,N_8751,N_8764);
or U9349 (N_9349,N_8811,N_8505);
or U9350 (N_9350,N_8928,N_8574);
or U9351 (N_9351,N_8507,N_8848);
xnor U9352 (N_9352,N_8934,N_8610);
nor U9353 (N_9353,N_8834,N_8694);
or U9354 (N_9354,N_8840,N_8559);
or U9355 (N_9355,N_8714,N_8713);
or U9356 (N_9356,N_8660,N_8558);
and U9357 (N_9357,N_8847,N_8840);
or U9358 (N_9358,N_8697,N_8888);
nor U9359 (N_9359,N_8724,N_8763);
or U9360 (N_9360,N_8659,N_8736);
and U9361 (N_9361,N_8565,N_8941);
nand U9362 (N_9362,N_8595,N_8562);
nand U9363 (N_9363,N_8685,N_8627);
xnor U9364 (N_9364,N_8688,N_8601);
or U9365 (N_9365,N_8743,N_8984);
nand U9366 (N_9366,N_8902,N_8778);
or U9367 (N_9367,N_8546,N_8656);
nand U9368 (N_9368,N_8537,N_8921);
or U9369 (N_9369,N_8768,N_8604);
xor U9370 (N_9370,N_8551,N_8838);
and U9371 (N_9371,N_8716,N_8527);
nand U9372 (N_9372,N_8892,N_8923);
nor U9373 (N_9373,N_8870,N_8863);
nand U9374 (N_9374,N_8708,N_8636);
nor U9375 (N_9375,N_8695,N_8651);
or U9376 (N_9376,N_8688,N_8597);
or U9377 (N_9377,N_8985,N_8716);
nor U9378 (N_9378,N_8503,N_8864);
and U9379 (N_9379,N_8800,N_8713);
xnor U9380 (N_9380,N_8851,N_8894);
xnor U9381 (N_9381,N_8541,N_8660);
xor U9382 (N_9382,N_8808,N_8791);
and U9383 (N_9383,N_8588,N_8574);
and U9384 (N_9384,N_8975,N_8577);
or U9385 (N_9385,N_8700,N_8634);
and U9386 (N_9386,N_8813,N_8714);
nand U9387 (N_9387,N_8525,N_8750);
nand U9388 (N_9388,N_8538,N_8509);
or U9389 (N_9389,N_8686,N_8554);
and U9390 (N_9390,N_8535,N_8859);
or U9391 (N_9391,N_8748,N_8938);
nor U9392 (N_9392,N_8672,N_8711);
or U9393 (N_9393,N_8556,N_8809);
nor U9394 (N_9394,N_8909,N_8615);
nor U9395 (N_9395,N_8541,N_8719);
and U9396 (N_9396,N_8807,N_8875);
and U9397 (N_9397,N_8924,N_8634);
or U9398 (N_9398,N_8568,N_8578);
or U9399 (N_9399,N_8760,N_8753);
or U9400 (N_9400,N_8894,N_8771);
nor U9401 (N_9401,N_8563,N_8678);
or U9402 (N_9402,N_8555,N_8564);
and U9403 (N_9403,N_8890,N_8800);
and U9404 (N_9404,N_8796,N_8807);
nand U9405 (N_9405,N_8508,N_8965);
and U9406 (N_9406,N_8835,N_8927);
and U9407 (N_9407,N_8862,N_8656);
xor U9408 (N_9408,N_8598,N_8564);
or U9409 (N_9409,N_8868,N_8748);
nand U9410 (N_9410,N_8617,N_8607);
and U9411 (N_9411,N_8687,N_8768);
nand U9412 (N_9412,N_8856,N_8602);
or U9413 (N_9413,N_8919,N_8811);
or U9414 (N_9414,N_8886,N_8894);
nor U9415 (N_9415,N_8598,N_8529);
nand U9416 (N_9416,N_8744,N_8679);
and U9417 (N_9417,N_8829,N_8726);
xor U9418 (N_9418,N_8634,N_8612);
xor U9419 (N_9419,N_8991,N_8987);
nand U9420 (N_9420,N_8775,N_8996);
nor U9421 (N_9421,N_8662,N_8754);
nor U9422 (N_9422,N_8892,N_8572);
and U9423 (N_9423,N_8703,N_8953);
xor U9424 (N_9424,N_8603,N_8748);
nor U9425 (N_9425,N_8749,N_8986);
or U9426 (N_9426,N_8518,N_8868);
or U9427 (N_9427,N_8696,N_8614);
or U9428 (N_9428,N_8576,N_8766);
or U9429 (N_9429,N_8978,N_8578);
or U9430 (N_9430,N_8942,N_8775);
and U9431 (N_9431,N_8873,N_8719);
and U9432 (N_9432,N_8924,N_8741);
and U9433 (N_9433,N_8814,N_8576);
nand U9434 (N_9434,N_8969,N_8821);
and U9435 (N_9435,N_8778,N_8769);
xor U9436 (N_9436,N_8669,N_8827);
xnor U9437 (N_9437,N_8876,N_8833);
nor U9438 (N_9438,N_8900,N_8809);
or U9439 (N_9439,N_8872,N_8517);
xor U9440 (N_9440,N_8798,N_8966);
nor U9441 (N_9441,N_8839,N_8792);
xnor U9442 (N_9442,N_8525,N_8659);
and U9443 (N_9443,N_8693,N_8765);
nor U9444 (N_9444,N_8621,N_8968);
nand U9445 (N_9445,N_8569,N_8567);
nor U9446 (N_9446,N_8845,N_8750);
nand U9447 (N_9447,N_8972,N_8572);
or U9448 (N_9448,N_8504,N_8575);
and U9449 (N_9449,N_8765,N_8934);
or U9450 (N_9450,N_8795,N_8618);
or U9451 (N_9451,N_8915,N_8709);
nor U9452 (N_9452,N_8652,N_8851);
nand U9453 (N_9453,N_8883,N_8746);
nor U9454 (N_9454,N_8952,N_8851);
xor U9455 (N_9455,N_8567,N_8749);
nor U9456 (N_9456,N_8500,N_8568);
or U9457 (N_9457,N_8884,N_8547);
xnor U9458 (N_9458,N_8817,N_8542);
nand U9459 (N_9459,N_8813,N_8961);
xor U9460 (N_9460,N_8921,N_8754);
and U9461 (N_9461,N_8992,N_8568);
xnor U9462 (N_9462,N_8697,N_8658);
nor U9463 (N_9463,N_8873,N_8971);
xnor U9464 (N_9464,N_8650,N_8811);
xnor U9465 (N_9465,N_8732,N_8757);
or U9466 (N_9466,N_8652,N_8585);
and U9467 (N_9467,N_8925,N_8530);
and U9468 (N_9468,N_8919,N_8874);
and U9469 (N_9469,N_8886,N_8517);
xor U9470 (N_9470,N_8658,N_8609);
xor U9471 (N_9471,N_8830,N_8691);
xnor U9472 (N_9472,N_8974,N_8576);
or U9473 (N_9473,N_8742,N_8589);
nand U9474 (N_9474,N_8504,N_8643);
xnor U9475 (N_9475,N_8992,N_8639);
nand U9476 (N_9476,N_8524,N_8580);
and U9477 (N_9477,N_8812,N_8956);
nand U9478 (N_9478,N_8525,N_8507);
and U9479 (N_9479,N_8672,N_8850);
nor U9480 (N_9480,N_8899,N_8690);
and U9481 (N_9481,N_8829,N_8819);
and U9482 (N_9482,N_8943,N_8924);
and U9483 (N_9483,N_8714,N_8539);
and U9484 (N_9484,N_8545,N_8507);
or U9485 (N_9485,N_8868,N_8931);
or U9486 (N_9486,N_8816,N_8699);
xnor U9487 (N_9487,N_8664,N_8727);
xnor U9488 (N_9488,N_8855,N_8579);
or U9489 (N_9489,N_8653,N_8784);
nor U9490 (N_9490,N_8858,N_8677);
nand U9491 (N_9491,N_8752,N_8852);
nand U9492 (N_9492,N_8511,N_8929);
nor U9493 (N_9493,N_8913,N_8805);
and U9494 (N_9494,N_8587,N_8708);
nor U9495 (N_9495,N_8842,N_8700);
or U9496 (N_9496,N_8653,N_8516);
or U9497 (N_9497,N_8695,N_8761);
nor U9498 (N_9498,N_8522,N_8615);
nand U9499 (N_9499,N_8822,N_8663);
nand U9500 (N_9500,N_9446,N_9271);
nor U9501 (N_9501,N_9292,N_9257);
or U9502 (N_9502,N_9469,N_9295);
or U9503 (N_9503,N_9357,N_9433);
xnor U9504 (N_9504,N_9392,N_9289);
and U9505 (N_9505,N_9494,N_9479);
or U9506 (N_9506,N_9437,N_9442);
or U9507 (N_9507,N_9455,N_9454);
nand U9508 (N_9508,N_9167,N_9421);
and U9509 (N_9509,N_9112,N_9407);
xor U9510 (N_9510,N_9283,N_9351);
nand U9511 (N_9511,N_9377,N_9113);
and U9512 (N_9512,N_9200,N_9320);
nor U9513 (N_9513,N_9001,N_9426);
nor U9514 (N_9514,N_9187,N_9337);
nor U9515 (N_9515,N_9157,N_9169);
nor U9516 (N_9516,N_9290,N_9011);
nand U9517 (N_9517,N_9405,N_9156);
and U9518 (N_9518,N_9419,N_9341);
nand U9519 (N_9519,N_9353,N_9339);
xnor U9520 (N_9520,N_9024,N_9010);
xnor U9521 (N_9521,N_9012,N_9141);
xnor U9522 (N_9522,N_9054,N_9122);
xnor U9523 (N_9523,N_9161,N_9155);
nand U9524 (N_9524,N_9043,N_9067);
xor U9525 (N_9525,N_9018,N_9131);
nor U9526 (N_9526,N_9160,N_9338);
xor U9527 (N_9527,N_9499,N_9017);
xnor U9528 (N_9528,N_9406,N_9014);
or U9529 (N_9529,N_9287,N_9291);
or U9530 (N_9530,N_9171,N_9129);
xor U9531 (N_9531,N_9366,N_9094);
nand U9532 (N_9532,N_9095,N_9227);
nand U9533 (N_9533,N_9253,N_9117);
nand U9534 (N_9534,N_9428,N_9116);
xnor U9535 (N_9535,N_9209,N_9079);
or U9536 (N_9536,N_9127,N_9281);
and U9537 (N_9537,N_9464,N_9324);
nor U9538 (N_9538,N_9432,N_9163);
nor U9539 (N_9539,N_9177,N_9027);
nor U9540 (N_9540,N_9175,N_9246);
and U9541 (N_9541,N_9435,N_9233);
and U9542 (N_9542,N_9026,N_9234);
nor U9543 (N_9543,N_9189,N_9279);
nor U9544 (N_9544,N_9180,N_9068);
and U9545 (N_9545,N_9195,N_9041);
nand U9546 (N_9546,N_9363,N_9472);
and U9547 (N_9547,N_9052,N_9359);
or U9548 (N_9548,N_9044,N_9051);
nand U9549 (N_9549,N_9184,N_9459);
nor U9550 (N_9550,N_9130,N_9329);
nand U9551 (N_9551,N_9013,N_9456);
nor U9552 (N_9552,N_9140,N_9276);
nand U9553 (N_9553,N_9417,N_9096);
or U9554 (N_9554,N_9458,N_9274);
and U9555 (N_9555,N_9321,N_9275);
and U9556 (N_9556,N_9286,N_9089);
and U9557 (N_9557,N_9237,N_9016);
and U9558 (N_9558,N_9115,N_9465);
and U9559 (N_9559,N_9362,N_9389);
or U9560 (N_9560,N_9133,N_9202);
nor U9561 (N_9561,N_9425,N_9106);
or U9562 (N_9562,N_9396,N_9258);
nand U9563 (N_9563,N_9100,N_9288);
or U9564 (N_9564,N_9046,N_9444);
xnor U9565 (N_9565,N_9420,N_9380);
or U9566 (N_9566,N_9092,N_9272);
xor U9567 (N_9567,N_9213,N_9222);
xor U9568 (N_9568,N_9042,N_9144);
nand U9569 (N_9569,N_9020,N_9206);
and U9570 (N_9570,N_9404,N_9193);
xnor U9571 (N_9571,N_9293,N_9102);
or U9572 (N_9572,N_9343,N_9109);
and U9573 (N_9573,N_9235,N_9008);
xnor U9574 (N_9574,N_9086,N_9039);
nor U9575 (N_9575,N_9267,N_9118);
nand U9576 (N_9576,N_9152,N_9153);
nand U9577 (N_9577,N_9378,N_9101);
nor U9578 (N_9578,N_9284,N_9422);
or U9579 (N_9579,N_9004,N_9361);
nand U9580 (N_9580,N_9477,N_9123);
or U9581 (N_9581,N_9326,N_9305);
xnor U9582 (N_9582,N_9059,N_9074);
or U9583 (N_9583,N_9229,N_9344);
nor U9584 (N_9584,N_9262,N_9453);
or U9585 (N_9585,N_9137,N_9081);
nor U9586 (N_9586,N_9483,N_9447);
nor U9587 (N_9587,N_9440,N_9073);
or U9588 (N_9588,N_9280,N_9098);
xor U9589 (N_9589,N_9040,N_9255);
and U9590 (N_9590,N_9121,N_9108);
or U9591 (N_9591,N_9402,N_9217);
xor U9592 (N_9592,N_9358,N_9119);
or U9593 (N_9593,N_9000,N_9260);
xnor U9594 (N_9594,N_9078,N_9037);
nor U9595 (N_9595,N_9087,N_9250);
or U9596 (N_9596,N_9110,N_9179);
or U9597 (N_9597,N_9069,N_9379);
nor U9598 (N_9598,N_9176,N_9308);
xnor U9599 (N_9599,N_9247,N_9307);
xor U9600 (N_9600,N_9450,N_9397);
xor U9601 (N_9601,N_9007,N_9231);
and U9602 (N_9602,N_9249,N_9104);
nand U9603 (N_9603,N_9266,N_9304);
or U9604 (N_9604,N_9080,N_9076);
xnor U9605 (N_9605,N_9224,N_9057);
nand U9606 (N_9606,N_9369,N_9452);
and U9607 (N_9607,N_9436,N_9107);
or U9608 (N_9608,N_9265,N_9294);
and U9609 (N_9609,N_9375,N_9314);
nor U9610 (N_9610,N_9482,N_9252);
xnor U9611 (N_9611,N_9411,N_9120);
or U9612 (N_9612,N_9461,N_9315);
and U9613 (N_9613,N_9484,N_9047);
nand U9614 (N_9614,N_9487,N_9225);
nor U9615 (N_9615,N_9423,N_9226);
nor U9616 (N_9616,N_9316,N_9241);
nor U9617 (N_9617,N_9395,N_9408);
and U9618 (N_9618,N_9198,N_9090);
or U9619 (N_9619,N_9055,N_9489);
xnor U9620 (N_9620,N_9356,N_9170);
nor U9621 (N_9621,N_9063,N_9413);
nand U9622 (N_9622,N_9478,N_9273);
xnor U9623 (N_9623,N_9188,N_9062);
and U9624 (N_9624,N_9302,N_9238);
xor U9625 (N_9625,N_9221,N_9345);
or U9626 (N_9626,N_9475,N_9135);
nand U9627 (N_9627,N_9367,N_9165);
and U9628 (N_9628,N_9263,N_9480);
or U9629 (N_9629,N_9330,N_9201);
nor U9630 (N_9630,N_9021,N_9053);
or U9631 (N_9631,N_9003,N_9497);
nand U9632 (N_9632,N_9332,N_9325);
or U9633 (N_9633,N_9498,N_9309);
xnor U9634 (N_9634,N_9083,N_9441);
xnor U9635 (N_9635,N_9173,N_9323);
nand U9636 (N_9636,N_9372,N_9145);
xnor U9637 (N_9637,N_9311,N_9183);
nor U9638 (N_9638,N_9493,N_9216);
nor U9639 (N_9639,N_9070,N_9409);
nand U9640 (N_9640,N_9399,N_9390);
or U9641 (N_9641,N_9207,N_9105);
and U9642 (N_9642,N_9354,N_9211);
xnor U9643 (N_9643,N_9139,N_9306);
xnor U9644 (N_9644,N_9296,N_9410);
xnor U9645 (N_9645,N_9005,N_9485);
or U9646 (N_9646,N_9150,N_9097);
nor U9647 (N_9647,N_9383,N_9085);
nand U9648 (N_9648,N_9429,N_9335);
xnor U9649 (N_9649,N_9300,N_9032);
and U9650 (N_9650,N_9182,N_9158);
and U9651 (N_9651,N_9319,N_9091);
nand U9652 (N_9652,N_9072,N_9387);
nand U9653 (N_9653,N_9278,N_9495);
nor U9654 (N_9654,N_9168,N_9365);
xnor U9655 (N_9655,N_9125,N_9342);
nand U9656 (N_9656,N_9268,N_9393);
and U9657 (N_9657,N_9214,N_9371);
nand U9658 (N_9658,N_9414,N_9232);
nor U9659 (N_9659,N_9394,N_9285);
nor U9660 (N_9660,N_9270,N_9208);
nor U9661 (N_9661,N_9025,N_9449);
nor U9662 (N_9662,N_9303,N_9259);
or U9663 (N_9663,N_9488,N_9033);
nor U9664 (N_9664,N_9126,N_9088);
and U9665 (N_9665,N_9071,N_9240);
nor U9666 (N_9666,N_9203,N_9355);
nor U9667 (N_9667,N_9061,N_9148);
and U9668 (N_9668,N_9467,N_9333);
and U9669 (N_9669,N_9142,N_9384);
or U9670 (N_9670,N_9373,N_9015);
nand U9671 (N_9671,N_9199,N_9212);
xnor U9672 (N_9672,N_9049,N_9388);
and U9673 (N_9673,N_9022,N_9256);
nand U9674 (N_9674,N_9299,N_9077);
nor U9675 (N_9675,N_9151,N_9205);
nor U9676 (N_9676,N_9269,N_9243);
or U9677 (N_9677,N_9374,N_9236);
xnor U9678 (N_9678,N_9242,N_9261);
nor U9679 (N_9679,N_9164,N_9154);
nand U9680 (N_9680,N_9382,N_9481);
xor U9681 (N_9681,N_9223,N_9192);
or U9682 (N_9682,N_9058,N_9368);
xnor U9683 (N_9683,N_9111,N_9196);
nand U9684 (N_9684,N_9386,N_9434);
and U9685 (N_9685,N_9491,N_9451);
or U9686 (N_9686,N_9317,N_9381);
nand U9687 (N_9687,N_9204,N_9313);
and U9688 (N_9688,N_9476,N_9401);
or U9689 (N_9689,N_9029,N_9282);
nand U9690 (N_9690,N_9416,N_9438);
nor U9691 (N_9691,N_9009,N_9376);
nor U9692 (N_9692,N_9471,N_9370);
or U9693 (N_9693,N_9352,N_9132);
or U9694 (N_9694,N_9385,N_9463);
or U9695 (N_9695,N_9347,N_9348);
nand U9696 (N_9696,N_9066,N_9473);
nor U9697 (N_9697,N_9228,N_9172);
and U9698 (N_9698,N_9492,N_9084);
and U9699 (N_9699,N_9099,N_9220);
nor U9700 (N_9700,N_9103,N_9138);
xor U9701 (N_9701,N_9346,N_9418);
nand U9702 (N_9702,N_9210,N_9350);
nor U9703 (N_9703,N_9298,N_9230);
nor U9704 (N_9704,N_9430,N_9400);
nand U9705 (N_9705,N_9297,N_9082);
nand U9706 (N_9706,N_9143,N_9219);
or U9707 (N_9707,N_9254,N_9178);
nor U9708 (N_9708,N_9439,N_9065);
xor U9709 (N_9709,N_9186,N_9159);
nor U9710 (N_9710,N_9050,N_9312);
nand U9711 (N_9711,N_9457,N_9136);
xnor U9712 (N_9712,N_9490,N_9443);
nor U9713 (N_9713,N_9060,N_9364);
xnor U9714 (N_9714,N_9190,N_9251);
xor U9715 (N_9715,N_9462,N_9336);
nand U9716 (N_9716,N_9093,N_9166);
or U9717 (N_9717,N_9124,N_9215);
nand U9718 (N_9718,N_9075,N_9028);
xnor U9719 (N_9719,N_9239,N_9470);
nor U9720 (N_9720,N_9244,N_9162);
and U9721 (N_9721,N_9328,N_9002);
nand U9722 (N_9722,N_9149,N_9030);
and U9723 (N_9723,N_9334,N_9398);
nor U9724 (N_9724,N_9128,N_9277);
nor U9725 (N_9725,N_9048,N_9448);
nor U9726 (N_9726,N_9006,N_9349);
and U9727 (N_9727,N_9019,N_9486);
xor U9728 (N_9728,N_9424,N_9264);
nand U9729 (N_9729,N_9340,N_9056);
nand U9730 (N_9730,N_9218,N_9301);
nand U9731 (N_9731,N_9248,N_9331);
or U9732 (N_9732,N_9460,N_9431);
or U9733 (N_9733,N_9391,N_9194);
nor U9734 (N_9734,N_9036,N_9310);
and U9735 (N_9735,N_9031,N_9191);
and U9736 (N_9736,N_9322,N_9147);
or U9737 (N_9737,N_9474,N_9427);
or U9738 (N_9738,N_9415,N_9064);
nor U9739 (N_9739,N_9403,N_9023);
nor U9740 (N_9740,N_9360,N_9038);
nor U9741 (N_9741,N_9445,N_9197);
or U9742 (N_9742,N_9327,N_9468);
xor U9743 (N_9743,N_9045,N_9466);
xor U9744 (N_9744,N_9174,N_9146);
nand U9745 (N_9745,N_9035,N_9412);
xor U9746 (N_9746,N_9496,N_9114);
nand U9747 (N_9747,N_9185,N_9034);
xnor U9748 (N_9748,N_9318,N_9134);
and U9749 (N_9749,N_9245,N_9181);
xnor U9750 (N_9750,N_9086,N_9487);
nor U9751 (N_9751,N_9442,N_9337);
nand U9752 (N_9752,N_9353,N_9367);
nor U9753 (N_9753,N_9304,N_9095);
xnor U9754 (N_9754,N_9092,N_9078);
nand U9755 (N_9755,N_9424,N_9092);
xor U9756 (N_9756,N_9221,N_9164);
xnor U9757 (N_9757,N_9201,N_9439);
or U9758 (N_9758,N_9276,N_9473);
nor U9759 (N_9759,N_9266,N_9442);
nand U9760 (N_9760,N_9138,N_9064);
or U9761 (N_9761,N_9294,N_9050);
nor U9762 (N_9762,N_9306,N_9068);
nand U9763 (N_9763,N_9424,N_9372);
xor U9764 (N_9764,N_9313,N_9081);
and U9765 (N_9765,N_9447,N_9379);
and U9766 (N_9766,N_9485,N_9151);
or U9767 (N_9767,N_9274,N_9026);
nand U9768 (N_9768,N_9159,N_9156);
or U9769 (N_9769,N_9416,N_9486);
or U9770 (N_9770,N_9076,N_9398);
nor U9771 (N_9771,N_9401,N_9137);
xnor U9772 (N_9772,N_9072,N_9448);
and U9773 (N_9773,N_9292,N_9428);
nand U9774 (N_9774,N_9301,N_9037);
nand U9775 (N_9775,N_9238,N_9325);
and U9776 (N_9776,N_9338,N_9318);
and U9777 (N_9777,N_9023,N_9469);
or U9778 (N_9778,N_9327,N_9187);
xor U9779 (N_9779,N_9082,N_9232);
nand U9780 (N_9780,N_9290,N_9199);
nand U9781 (N_9781,N_9352,N_9098);
xor U9782 (N_9782,N_9468,N_9122);
nor U9783 (N_9783,N_9492,N_9221);
nor U9784 (N_9784,N_9221,N_9199);
or U9785 (N_9785,N_9341,N_9349);
or U9786 (N_9786,N_9294,N_9442);
nand U9787 (N_9787,N_9349,N_9131);
nor U9788 (N_9788,N_9071,N_9445);
or U9789 (N_9789,N_9274,N_9364);
or U9790 (N_9790,N_9205,N_9493);
and U9791 (N_9791,N_9251,N_9404);
and U9792 (N_9792,N_9336,N_9315);
and U9793 (N_9793,N_9481,N_9124);
and U9794 (N_9794,N_9089,N_9315);
or U9795 (N_9795,N_9376,N_9162);
or U9796 (N_9796,N_9094,N_9476);
or U9797 (N_9797,N_9252,N_9474);
or U9798 (N_9798,N_9213,N_9015);
or U9799 (N_9799,N_9288,N_9253);
xnor U9800 (N_9800,N_9414,N_9393);
or U9801 (N_9801,N_9390,N_9494);
or U9802 (N_9802,N_9312,N_9070);
and U9803 (N_9803,N_9339,N_9101);
nand U9804 (N_9804,N_9216,N_9444);
nand U9805 (N_9805,N_9234,N_9113);
nor U9806 (N_9806,N_9349,N_9168);
xor U9807 (N_9807,N_9122,N_9490);
xor U9808 (N_9808,N_9471,N_9354);
nand U9809 (N_9809,N_9469,N_9350);
nand U9810 (N_9810,N_9491,N_9058);
or U9811 (N_9811,N_9150,N_9166);
nand U9812 (N_9812,N_9311,N_9462);
or U9813 (N_9813,N_9057,N_9252);
nand U9814 (N_9814,N_9261,N_9279);
xnor U9815 (N_9815,N_9489,N_9283);
nand U9816 (N_9816,N_9309,N_9189);
xnor U9817 (N_9817,N_9244,N_9492);
or U9818 (N_9818,N_9338,N_9186);
and U9819 (N_9819,N_9053,N_9471);
and U9820 (N_9820,N_9208,N_9085);
xnor U9821 (N_9821,N_9159,N_9210);
xnor U9822 (N_9822,N_9042,N_9211);
and U9823 (N_9823,N_9164,N_9210);
nand U9824 (N_9824,N_9076,N_9475);
nand U9825 (N_9825,N_9110,N_9490);
and U9826 (N_9826,N_9015,N_9135);
nand U9827 (N_9827,N_9435,N_9006);
xnor U9828 (N_9828,N_9108,N_9174);
nand U9829 (N_9829,N_9389,N_9080);
nor U9830 (N_9830,N_9112,N_9205);
or U9831 (N_9831,N_9111,N_9322);
nor U9832 (N_9832,N_9319,N_9374);
or U9833 (N_9833,N_9327,N_9167);
nand U9834 (N_9834,N_9060,N_9498);
nand U9835 (N_9835,N_9303,N_9460);
or U9836 (N_9836,N_9041,N_9304);
nand U9837 (N_9837,N_9123,N_9284);
xor U9838 (N_9838,N_9389,N_9240);
xor U9839 (N_9839,N_9164,N_9040);
xor U9840 (N_9840,N_9162,N_9368);
or U9841 (N_9841,N_9279,N_9463);
xor U9842 (N_9842,N_9373,N_9157);
xor U9843 (N_9843,N_9269,N_9113);
and U9844 (N_9844,N_9165,N_9334);
or U9845 (N_9845,N_9406,N_9254);
xor U9846 (N_9846,N_9135,N_9120);
or U9847 (N_9847,N_9247,N_9071);
xnor U9848 (N_9848,N_9217,N_9395);
xor U9849 (N_9849,N_9065,N_9300);
nor U9850 (N_9850,N_9311,N_9454);
or U9851 (N_9851,N_9169,N_9121);
or U9852 (N_9852,N_9036,N_9037);
nand U9853 (N_9853,N_9489,N_9429);
or U9854 (N_9854,N_9041,N_9408);
xnor U9855 (N_9855,N_9073,N_9385);
or U9856 (N_9856,N_9159,N_9070);
nor U9857 (N_9857,N_9290,N_9213);
or U9858 (N_9858,N_9153,N_9248);
and U9859 (N_9859,N_9046,N_9282);
nand U9860 (N_9860,N_9499,N_9361);
and U9861 (N_9861,N_9064,N_9123);
xnor U9862 (N_9862,N_9035,N_9467);
nand U9863 (N_9863,N_9150,N_9481);
or U9864 (N_9864,N_9027,N_9379);
nand U9865 (N_9865,N_9496,N_9388);
nor U9866 (N_9866,N_9417,N_9099);
or U9867 (N_9867,N_9342,N_9311);
or U9868 (N_9868,N_9067,N_9402);
and U9869 (N_9869,N_9332,N_9189);
or U9870 (N_9870,N_9324,N_9272);
and U9871 (N_9871,N_9248,N_9297);
nand U9872 (N_9872,N_9443,N_9068);
and U9873 (N_9873,N_9475,N_9426);
or U9874 (N_9874,N_9403,N_9183);
xnor U9875 (N_9875,N_9226,N_9064);
xnor U9876 (N_9876,N_9038,N_9146);
nor U9877 (N_9877,N_9012,N_9207);
and U9878 (N_9878,N_9123,N_9372);
nand U9879 (N_9879,N_9436,N_9072);
nor U9880 (N_9880,N_9222,N_9404);
xor U9881 (N_9881,N_9212,N_9093);
or U9882 (N_9882,N_9158,N_9446);
and U9883 (N_9883,N_9044,N_9083);
and U9884 (N_9884,N_9298,N_9461);
nor U9885 (N_9885,N_9131,N_9423);
nor U9886 (N_9886,N_9424,N_9014);
or U9887 (N_9887,N_9346,N_9116);
xor U9888 (N_9888,N_9412,N_9467);
nor U9889 (N_9889,N_9263,N_9352);
xnor U9890 (N_9890,N_9109,N_9435);
xnor U9891 (N_9891,N_9122,N_9167);
xnor U9892 (N_9892,N_9218,N_9238);
nand U9893 (N_9893,N_9267,N_9290);
and U9894 (N_9894,N_9178,N_9396);
and U9895 (N_9895,N_9380,N_9287);
or U9896 (N_9896,N_9276,N_9440);
nand U9897 (N_9897,N_9288,N_9237);
nand U9898 (N_9898,N_9083,N_9035);
nor U9899 (N_9899,N_9339,N_9069);
and U9900 (N_9900,N_9296,N_9193);
xor U9901 (N_9901,N_9006,N_9433);
and U9902 (N_9902,N_9207,N_9078);
nor U9903 (N_9903,N_9015,N_9004);
nand U9904 (N_9904,N_9426,N_9241);
or U9905 (N_9905,N_9108,N_9301);
xor U9906 (N_9906,N_9424,N_9438);
xor U9907 (N_9907,N_9239,N_9041);
nor U9908 (N_9908,N_9489,N_9087);
or U9909 (N_9909,N_9171,N_9461);
xnor U9910 (N_9910,N_9107,N_9085);
and U9911 (N_9911,N_9187,N_9194);
nor U9912 (N_9912,N_9129,N_9251);
xnor U9913 (N_9913,N_9082,N_9435);
or U9914 (N_9914,N_9181,N_9166);
nor U9915 (N_9915,N_9200,N_9022);
xor U9916 (N_9916,N_9474,N_9497);
or U9917 (N_9917,N_9401,N_9381);
or U9918 (N_9918,N_9039,N_9221);
nand U9919 (N_9919,N_9075,N_9398);
or U9920 (N_9920,N_9263,N_9079);
xnor U9921 (N_9921,N_9311,N_9011);
or U9922 (N_9922,N_9265,N_9440);
nand U9923 (N_9923,N_9340,N_9046);
and U9924 (N_9924,N_9423,N_9358);
or U9925 (N_9925,N_9235,N_9499);
and U9926 (N_9926,N_9163,N_9293);
xor U9927 (N_9927,N_9315,N_9081);
nand U9928 (N_9928,N_9116,N_9230);
nand U9929 (N_9929,N_9172,N_9108);
xor U9930 (N_9930,N_9438,N_9172);
xnor U9931 (N_9931,N_9342,N_9253);
and U9932 (N_9932,N_9059,N_9455);
nor U9933 (N_9933,N_9249,N_9377);
nand U9934 (N_9934,N_9325,N_9118);
nand U9935 (N_9935,N_9457,N_9028);
nor U9936 (N_9936,N_9251,N_9333);
xor U9937 (N_9937,N_9428,N_9071);
nand U9938 (N_9938,N_9305,N_9193);
nor U9939 (N_9939,N_9146,N_9200);
or U9940 (N_9940,N_9049,N_9144);
nand U9941 (N_9941,N_9124,N_9202);
and U9942 (N_9942,N_9039,N_9144);
or U9943 (N_9943,N_9282,N_9257);
nand U9944 (N_9944,N_9275,N_9044);
and U9945 (N_9945,N_9254,N_9488);
and U9946 (N_9946,N_9056,N_9368);
nand U9947 (N_9947,N_9404,N_9129);
and U9948 (N_9948,N_9352,N_9156);
nand U9949 (N_9949,N_9403,N_9484);
and U9950 (N_9950,N_9428,N_9472);
or U9951 (N_9951,N_9141,N_9037);
nor U9952 (N_9952,N_9044,N_9137);
xnor U9953 (N_9953,N_9325,N_9389);
nor U9954 (N_9954,N_9353,N_9444);
and U9955 (N_9955,N_9075,N_9222);
or U9956 (N_9956,N_9274,N_9262);
or U9957 (N_9957,N_9275,N_9499);
or U9958 (N_9958,N_9121,N_9350);
nor U9959 (N_9959,N_9193,N_9231);
or U9960 (N_9960,N_9409,N_9226);
and U9961 (N_9961,N_9246,N_9397);
nand U9962 (N_9962,N_9318,N_9012);
and U9963 (N_9963,N_9328,N_9498);
or U9964 (N_9964,N_9471,N_9361);
nand U9965 (N_9965,N_9296,N_9034);
or U9966 (N_9966,N_9304,N_9023);
and U9967 (N_9967,N_9228,N_9275);
nand U9968 (N_9968,N_9202,N_9225);
and U9969 (N_9969,N_9237,N_9231);
or U9970 (N_9970,N_9203,N_9307);
nand U9971 (N_9971,N_9337,N_9221);
nand U9972 (N_9972,N_9106,N_9384);
nand U9973 (N_9973,N_9157,N_9253);
xnor U9974 (N_9974,N_9013,N_9216);
nor U9975 (N_9975,N_9367,N_9358);
or U9976 (N_9976,N_9026,N_9006);
xor U9977 (N_9977,N_9197,N_9358);
nand U9978 (N_9978,N_9036,N_9024);
nor U9979 (N_9979,N_9283,N_9481);
nand U9980 (N_9980,N_9107,N_9135);
nor U9981 (N_9981,N_9414,N_9389);
and U9982 (N_9982,N_9153,N_9146);
or U9983 (N_9983,N_9264,N_9392);
or U9984 (N_9984,N_9436,N_9286);
or U9985 (N_9985,N_9014,N_9429);
xnor U9986 (N_9986,N_9202,N_9176);
or U9987 (N_9987,N_9352,N_9253);
nand U9988 (N_9988,N_9104,N_9251);
nand U9989 (N_9989,N_9431,N_9342);
and U9990 (N_9990,N_9375,N_9049);
xor U9991 (N_9991,N_9413,N_9363);
nand U9992 (N_9992,N_9444,N_9219);
nor U9993 (N_9993,N_9196,N_9499);
and U9994 (N_9994,N_9394,N_9457);
nand U9995 (N_9995,N_9064,N_9361);
nor U9996 (N_9996,N_9266,N_9392);
xor U9997 (N_9997,N_9367,N_9197);
nand U9998 (N_9998,N_9295,N_9407);
nor U9999 (N_9999,N_9073,N_9391);
xor U10000 (N_10000,N_9968,N_9746);
and U10001 (N_10001,N_9615,N_9669);
nand U10002 (N_10002,N_9963,N_9725);
nor U10003 (N_10003,N_9506,N_9837);
nand U10004 (N_10004,N_9905,N_9886);
or U10005 (N_10005,N_9976,N_9643);
and U10006 (N_10006,N_9564,N_9620);
nand U10007 (N_10007,N_9881,N_9740);
xor U10008 (N_10008,N_9890,N_9668);
and U10009 (N_10009,N_9546,N_9505);
or U10010 (N_10010,N_9532,N_9866);
nor U10011 (N_10011,N_9846,N_9551);
and U10012 (N_10012,N_9629,N_9747);
xor U10013 (N_10013,N_9941,N_9695);
nor U10014 (N_10014,N_9992,N_9859);
xor U10015 (N_10015,N_9541,N_9875);
or U10016 (N_10016,N_9873,N_9673);
xor U10017 (N_10017,N_9853,N_9674);
nor U10018 (N_10018,N_9844,N_9533);
nand U10019 (N_10019,N_9775,N_9809);
xnor U10020 (N_10020,N_9504,N_9694);
or U10021 (N_10021,N_9978,N_9940);
nor U10022 (N_10022,N_9582,N_9958);
or U10023 (N_10023,N_9681,N_9655);
nand U10024 (N_10024,N_9787,N_9573);
xor U10025 (N_10025,N_9901,N_9675);
xnor U10026 (N_10026,N_9916,N_9852);
nand U10027 (N_10027,N_9628,N_9501);
nor U10028 (N_10028,N_9788,N_9634);
nand U10029 (N_10029,N_9765,N_9715);
nand U10030 (N_10030,N_9748,N_9945);
xor U10031 (N_10031,N_9516,N_9662);
xor U10032 (N_10032,N_9847,N_9585);
or U10033 (N_10033,N_9816,N_9897);
xnor U10034 (N_10034,N_9648,N_9800);
and U10035 (N_10035,N_9979,N_9697);
nand U10036 (N_10036,N_9909,N_9636);
and U10037 (N_10037,N_9927,N_9877);
xor U10038 (N_10038,N_9796,N_9828);
xor U10039 (N_10039,N_9749,N_9601);
and U10040 (N_10040,N_9913,N_9754);
and U10041 (N_10041,N_9821,N_9861);
nand U10042 (N_10042,N_9633,N_9528);
nor U10043 (N_10043,N_9683,N_9760);
and U10044 (N_10044,N_9857,N_9918);
nand U10045 (N_10045,N_9574,N_9892);
or U10046 (N_10046,N_9584,N_9562);
nand U10047 (N_10047,N_9794,N_9649);
or U10048 (N_10048,N_9680,N_9708);
xnor U10049 (N_10049,N_9772,N_9540);
xor U10050 (N_10050,N_9935,N_9621);
xnor U10051 (N_10051,N_9825,N_9845);
nand U10052 (N_10052,N_9991,N_9730);
and U10053 (N_10053,N_9961,N_9572);
nand U10054 (N_10054,N_9952,N_9616);
and U10055 (N_10055,N_9637,N_9849);
and U10056 (N_10056,N_9666,N_9783);
nor U10057 (N_10057,N_9781,N_9842);
nand U10058 (N_10058,N_9644,N_9594);
xnor U10059 (N_10059,N_9670,N_9738);
nor U10060 (N_10060,N_9508,N_9936);
nand U10061 (N_10061,N_9630,N_9811);
xnor U10062 (N_10062,N_9595,N_9672);
nand U10063 (N_10063,N_9663,N_9912);
xor U10064 (N_10064,N_9704,N_9512);
nand U10065 (N_10065,N_9509,N_9706);
nand U10066 (N_10066,N_9997,N_9851);
or U10067 (N_10067,N_9947,N_9566);
nor U10068 (N_10068,N_9972,N_9946);
xnor U10069 (N_10069,N_9719,N_9870);
or U10070 (N_10070,N_9780,N_9915);
or U10071 (N_10071,N_9711,N_9826);
nor U10072 (N_10072,N_9969,N_9898);
and U10073 (N_10073,N_9654,N_9640);
xnor U10074 (N_10074,N_9676,N_9503);
nand U10075 (N_10075,N_9933,N_9613);
or U10076 (N_10076,N_9980,N_9717);
or U10077 (N_10077,N_9771,N_9661);
and U10078 (N_10078,N_9885,N_9657);
xor U10079 (N_10079,N_9538,N_9750);
nand U10080 (N_10080,N_9843,N_9510);
or U10081 (N_10081,N_9819,N_9549);
and U10082 (N_10082,N_9865,N_9959);
or U10083 (N_10083,N_9838,N_9756);
or U10084 (N_10084,N_9822,N_9544);
nor U10085 (N_10085,N_9815,N_9710);
nand U10086 (N_10086,N_9688,N_9735);
nand U10087 (N_10087,N_9949,N_9656);
or U10088 (N_10088,N_9817,N_9966);
xor U10089 (N_10089,N_9728,N_9632);
xor U10090 (N_10090,N_9893,N_9791);
xor U10091 (N_10091,N_9736,N_9593);
and U10092 (N_10092,N_9827,N_9526);
and U10093 (N_10093,N_9626,N_9934);
or U10094 (N_10094,N_9888,N_9718);
xnor U10095 (N_10095,N_9721,N_9555);
nand U10096 (N_10096,N_9962,N_9923);
or U10097 (N_10097,N_9587,N_9539);
nand U10098 (N_10098,N_9967,N_9970);
nand U10099 (N_10099,N_9753,N_9926);
and U10100 (N_10100,N_9906,N_9502);
nand U10101 (N_10101,N_9563,N_9999);
and U10102 (N_10102,N_9521,N_9820);
nand U10103 (N_10103,N_9611,N_9910);
and U10104 (N_10104,N_9589,N_9884);
and U10105 (N_10105,N_9872,N_9922);
nand U10106 (N_10106,N_9790,N_9543);
xor U10107 (N_10107,N_9763,N_9651);
xor U10108 (N_10108,N_9659,N_9698);
or U10109 (N_10109,N_9863,N_9841);
and U10110 (N_10110,N_9565,N_9530);
and U10111 (N_10111,N_9802,N_9829);
nand U10112 (N_10112,N_9642,N_9995);
or U10113 (N_10113,N_9631,N_9939);
nand U10114 (N_10114,N_9732,N_9557);
nor U10115 (N_10115,N_9840,N_9617);
nand U10116 (N_10116,N_9578,N_9804);
xnor U10117 (N_10117,N_9824,N_9702);
xor U10118 (N_10118,N_9950,N_9646);
nor U10119 (N_10119,N_9994,N_9786);
and U10120 (N_10120,N_9925,N_9887);
or U10121 (N_10121,N_9839,N_9696);
nand U10122 (N_10122,N_9973,N_9832);
or U10123 (N_10123,N_9591,N_9801);
or U10124 (N_10124,N_9712,N_9608);
or U10125 (N_10125,N_9560,N_9686);
xor U10126 (N_10126,N_9592,N_9511);
nor U10127 (N_10127,N_9977,N_9514);
and U10128 (N_10128,N_9720,N_9998);
nand U10129 (N_10129,N_9836,N_9685);
nand U10130 (N_10130,N_9938,N_9729);
nor U10131 (N_10131,N_9924,N_9814);
xnor U10132 (N_10132,N_9583,N_9773);
nor U10133 (N_10133,N_9792,N_9757);
nand U10134 (N_10134,N_9567,N_9919);
xor U10135 (N_10135,N_9951,N_9990);
nor U10136 (N_10136,N_9982,N_9606);
nor U10137 (N_10137,N_9871,N_9568);
or U10138 (N_10138,N_9907,N_9818);
and U10139 (N_10139,N_9603,N_9895);
xor U10140 (N_10140,N_9722,N_9577);
nor U10141 (N_10141,N_9614,N_9806);
and U10142 (N_10142,N_9525,N_9707);
or U10143 (N_10143,N_9709,N_9914);
xnor U10144 (N_10144,N_9580,N_9547);
and U10145 (N_10145,N_9625,N_9727);
xnor U10146 (N_10146,N_9904,N_9799);
xor U10147 (N_10147,N_9768,N_9988);
xnor U10148 (N_10148,N_9974,N_9553);
or U10149 (N_10149,N_9678,N_9784);
or U10150 (N_10150,N_9536,N_9855);
and U10151 (N_10151,N_9523,N_9703);
xor U10152 (N_10152,N_9743,N_9679);
xor U10153 (N_10153,N_9548,N_9745);
nand U10154 (N_10154,N_9894,N_9627);
and U10155 (N_10155,N_9689,N_9987);
or U10156 (N_10156,N_9879,N_9575);
nand U10157 (N_10157,N_9789,N_9986);
or U10158 (N_10158,N_9953,N_9714);
xnor U10159 (N_10159,N_9535,N_9891);
xor U10160 (N_10160,N_9902,N_9604);
xor U10161 (N_10161,N_9724,N_9831);
or U10162 (N_10162,N_9652,N_9639);
and U10163 (N_10163,N_9778,N_9571);
nand U10164 (N_10164,N_9527,N_9758);
and U10165 (N_10165,N_9954,N_9742);
nor U10166 (N_10166,N_9860,N_9880);
xnor U10167 (N_10167,N_9975,N_9684);
xnor U10168 (N_10168,N_9660,N_9576);
and U10169 (N_10169,N_9984,N_9600);
xor U10170 (N_10170,N_9705,N_9807);
or U10171 (N_10171,N_9653,N_9751);
nand U10172 (N_10172,N_9797,N_9713);
or U10173 (N_10173,N_9744,N_9638);
xnor U10174 (N_10174,N_9609,N_9700);
xnor U10175 (N_10175,N_9833,N_9687);
nand U10176 (N_10176,N_9948,N_9517);
nand U10177 (N_10177,N_9597,N_9518);
and U10178 (N_10178,N_9964,N_9943);
and U10179 (N_10179,N_9782,N_9917);
or U10180 (N_10180,N_9739,N_9699);
nand U10181 (N_10181,N_9607,N_9776);
nor U10182 (N_10182,N_9764,N_9647);
and U10183 (N_10183,N_9579,N_9513);
or U10184 (N_10184,N_9928,N_9691);
nand U10185 (N_10185,N_9610,N_9590);
and U10186 (N_10186,N_9779,N_9955);
nor U10187 (N_10187,N_9692,N_9622);
and U10188 (N_10188,N_9876,N_9701);
or U10189 (N_10189,N_9883,N_9542);
or U10190 (N_10190,N_9612,N_9965);
and U10191 (N_10191,N_9889,N_9682);
xor U10192 (N_10192,N_9723,N_9920);
and U10193 (N_10193,N_9500,N_9671);
xnor U10194 (N_10194,N_9645,N_9805);
xor U10195 (N_10195,N_9869,N_9769);
or U10196 (N_10196,N_9731,N_9856);
and U10197 (N_10197,N_9561,N_9664);
and U10198 (N_10198,N_9900,N_9677);
xnor U10199 (N_10199,N_9770,N_9996);
nor U10200 (N_10200,N_9619,N_9529);
nor U10201 (N_10201,N_9911,N_9774);
nor U10202 (N_10202,N_9605,N_9602);
or U10203 (N_10203,N_9850,N_9569);
or U10204 (N_10204,N_9868,N_9823);
nor U10205 (N_10205,N_9848,N_9534);
nand U10206 (N_10206,N_9766,N_9921);
xor U10207 (N_10207,N_9858,N_9785);
xor U10208 (N_10208,N_9864,N_9767);
xor U10209 (N_10209,N_9930,N_9777);
nor U10210 (N_10210,N_9741,N_9795);
nand U10211 (N_10211,N_9650,N_9588);
nand U10212 (N_10212,N_9618,N_9808);
and U10213 (N_10213,N_9899,N_9903);
xor U10214 (N_10214,N_9545,N_9641);
or U10215 (N_10215,N_9929,N_9862);
or U10216 (N_10216,N_9524,N_9874);
or U10217 (N_10217,N_9599,N_9623);
or U10218 (N_10218,N_9798,N_9882);
nand U10219 (N_10219,N_9944,N_9624);
or U10220 (N_10220,N_9693,N_9762);
nor U10221 (N_10221,N_9793,N_9830);
xnor U10222 (N_10222,N_9983,N_9810);
or U10223 (N_10223,N_9985,N_9667);
xor U10224 (N_10224,N_9598,N_9755);
xor U10225 (N_10225,N_9531,N_9556);
nor U10226 (N_10226,N_9665,N_9554);
nand U10227 (N_10227,N_9956,N_9957);
xnor U10228 (N_10228,N_9908,N_9522);
and U10229 (N_10229,N_9581,N_9981);
or U10230 (N_10230,N_9552,N_9507);
nand U10231 (N_10231,N_9570,N_9726);
and U10232 (N_10232,N_9759,N_9812);
and U10233 (N_10233,N_9537,N_9896);
nand U10234 (N_10234,N_9716,N_9586);
nor U10235 (N_10235,N_9559,N_9854);
or U10236 (N_10236,N_9519,N_9515);
nor U10237 (N_10237,N_9971,N_9867);
and U10238 (N_10238,N_9993,N_9937);
nor U10239 (N_10239,N_9989,N_9931);
and U10240 (N_10240,N_9878,N_9813);
nor U10241 (N_10241,N_9737,N_9734);
and U10242 (N_10242,N_9733,N_9752);
or U10243 (N_10243,N_9635,N_9761);
or U10244 (N_10244,N_9803,N_9658);
or U10245 (N_10245,N_9834,N_9835);
or U10246 (N_10246,N_9596,N_9942);
nor U10247 (N_10247,N_9550,N_9690);
and U10248 (N_10248,N_9932,N_9558);
and U10249 (N_10249,N_9520,N_9960);
nand U10250 (N_10250,N_9704,N_9962);
nor U10251 (N_10251,N_9871,N_9915);
nand U10252 (N_10252,N_9844,N_9942);
xor U10253 (N_10253,N_9846,N_9779);
xnor U10254 (N_10254,N_9956,N_9719);
or U10255 (N_10255,N_9738,N_9928);
xnor U10256 (N_10256,N_9988,N_9790);
nand U10257 (N_10257,N_9569,N_9693);
or U10258 (N_10258,N_9549,N_9672);
nand U10259 (N_10259,N_9824,N_9820);
nor U10260 (N_10260,N_9793,N_9643);
xnor U10261 (N_10261,N_9712,N_9716);
xor U10262 (N_10262,N_9914,N_9853);
and U10263 (N_10263,N_9881,N_9886);
nor U10264 (N_10264,N_9707,N_9817);
xor U10265 (N_10265,N_9868,N_9745);
and U10266 (N_10266,N_9522,N_9711);
nand U10267 (N_10267,N_9828,N_9780);
nor U10268 (N_10268,N_9547,N_9684);
or U10269 (N_10269,N_9954,N_9721);
xnor U10270 (N_10270,N_9793,N_9524);
nand U10271 (N_10271,N_9754,N_9670);
and U10272 (N_10272,N_9910,N_9908);
or U10273 (N_10273,N_9737,N_9840);
and U10274 (N_10274,N_9538,N_9881);
nor U10275 (N_10275,N_9919,N_9535);
or U10276 (N_10276,N_9534,N_9596);
nor U10277 (N_10277,N_9862,N_9688);
xor U10278 (N_10278,N_9879,N_9738);
and U10279 (N_10279,N_9650,N_9758);
or U10280 (N_10280,N_9513,N_9783);
or U10281 (N_10281,N_9868,N_9998);
and U10282 (N_10282,N_9864,N_9798);
and U10283 (N_10283,N_9550,N_9939);
or U10284 (N_10284,N_9979,N_9953);
and U10285 (N_10285,N_9937,N_9979);
nor U10286 (N_10286,N_9765,N_9817);
nor U10287 (N_10287,N_9854,N_9888);
nand U10288 (N_10288,N_9577,N_9930);
and U10289 (N_10289,N_9540,N_9882);
nand U10290 (N_10290,N_9526,N_9806);
nor U10291 (N_10291,N_9708,N_9582);
or U10292 (N_10292,N_9880,N_9925);
nand U10293 (N_10293,N_9690,N_9658);
nand U10294 (N_10294,N_9912,N_9803);
nand U10295 (N_10295,N_9530,N_9937);
or U10296 (N_10296,N_9866,N_9834);
xnor U10297 (N_10297,N_9941,N_9975);
nand U10298 (N_10298,N_9930,N_9552);
and U10299 (N_10299,N_9684,N_9611);
and U10300 (N_10300,N_9655,N_9996);
xnor U10301 (N_10301,N_9555,N_9706);
xor U10302 (N_10302,N_9615,N_9879);
xnor U10303 (N_10303,N_9576,N_9543);
and U10304 (N_10304,N_9645,N_9585);
nor U10305 (N_10305,N_9962,N_9859);
and U10306 (N_10306,N_9500,N_9944);
or U10307 (N_10307,N_9877,N_9514);
or U10308 (N_10308,N_9525,N_9604);
nor U10309 (N_10309,N_9662,N_9554);
and U10310 (N_10310,N_9611,N_9884);
nand U10311 (N_10311,N_9936,N_9536);
xnor U10312 (N_10312,N_9993,N_9841);
xnor U10313 (N_10313,N_9696,N_9716);
nor U10314 (N_10314,N_9884,N_9814);
or U10315 (N_10315,N_9668,N_9784);
nor U10316 (N_10316,N_9995,N_9526);
nor U10317 (N_10317,N_9892,N_9575);
and U10318 (N_10318,N_9781,N_9684);
or U10319 (N_10319,N_9915,N_9787);
nand U10320 (N_10320,N_9631,N_9994);
and U10321 (N_10321,N_9617,N_9641);
nor U10322 (N_10322,N_9588,N_9589);
and U10323 (N_10323,N_9980,N_9530);
nand U10324 (N_10324,N_9929,N_9948);
nand U10325 (N_10325,N_9918,N_9745);
and U10326 (N_10326,N_9945,N_9948);
and U10327 (N_10327,N_9741,N_9794);
xor U10328 (N_10328,N_9661,N_9576);
xor U10329 (N_10329,N_9669,N_9957);
or U10330 (N_10330,N_9533,N_9850);
or U10331 (N_10331,N_9824,N_9908);
nor U10332 (N_10332,N_9603,N_9628);
or U10333 (N_10333,N_9865,N_9890);
or U10334 (N_10334,N_9736,N_9755);
and U10335 (N_10335,N_9817,N_9835);
or U10336 (N_10336,N_9734,N_9559);
or U10337 (N_10337,N_9974,N_9765);
xnor U10338 (N_10338,N_9706,N_9648);
nand U10339 (N_10339,N_9950,N_9949);
nand U10340 (N_10340,N_9972,N_9548);
xor U10341 (N_10341,N_9642,N_9729);
or U10342 (N_10342,N_9985,N_9804);
or U10343 (N_10343,N_9655,N_9553);
and U10344 (N_10344,N_9803,N_9638);
and U10345 (N_10345,N_9858,N_9512);
and U10346 (N_10346,N_9554,N_9854);
xnor U10347 (N_10347,N_9858,N_9939);
nand U10348 (N_10348,N_9859,N_9843);
or U10349 (N_10349,N_9895,N_9992);
or U10350 (N_10350,N_9573,N_9823);
and U10351 (N_10351,N_9902,N_9851);
nor U10352 (N_10352,N_9973,N_9785);
nand U10353 (N_10353,N_9744,N_9972);
nor U10354 (N_10354,N_9630,N_9788);
xnor U10355 (N_10355,N_9583,N_9606);
and U10356 (N_10356,N_9587,N_9850);
nor U10357 (N_10357,N_9752,N_9563);
and U10358 (N_10358,N_9711,N_9512);
nand U10359 (N_10359,N_9819,N_9730);
and U10360 (N_10360,N_9714,N_9701);
and U10361 (N_10361,N_9739,N_9516);
or U10362 (N_10362,N_9760,N_9764);
or U10363 (N_10363,N_9586,N_9582);
and U10364 (N_10364,N_9856,N_9593);
or U10365 (N_10365,N_9566,N_9722);
nor U10366 (N_10366,N_9698,N_9526);
nand U10367 (N_10367,N_9933,N_9729);
and U10368 (N_10368,N_9949,N_9612);
or U10369 (N_10369,N_9601,N_9754);
xnor U10370 (N_10370,N_9943,N_9939);
and U10371 (N_10371,N_9646,N_9598);
xnor U10372 (N_10372,N_9803,N_9928);
and U10373 (N_10373,N_9591,N_9731);
or U10374 (N_10374,N_9720,N_9993);
nor U10375 (N_10375,N_9924,N_9722);
xnor U10376 (N_10376,N_9718,N_9530);
xor U10377 (N_10377,N_9810,N_9663);
and U10378 (N_10378,N_9501,N_9522);
nor U10379 (N_10379,N_9973,N_9661);
or U10380 (N_10380,N_9646,N_9865);
and U10381 (N_10381,N_9703,N_9970);
nand U10382 (N_10382,N_9964,N_9826);
and U10383 (N_10383,N_9920,N_9852);
or U10384 (N_10384,N_9977,N_9745);
and U10385 (N_10385,N_9582,N_9652);
xor U10386 (N_10386,N_9847,N_9605);
nand U10387 (N_10387,N_9661,N_9761);
and U10388 (N_10388,N_9767,N_9906);
or U10389 (N_10389,N_9688,N_9549);
and U10390 (N_10390,N_9967,N_9641);
or U10391 (N_10391,N_9734,N_9776);
or U10392 (N_10392,N_9829,N_9898);
or U10393 (N_10393,N_9841,N_9599);
nand U10394 (N_10394,N_9967,N_9651);
nor U10395 (N_10395,N_9960,N_9895);
or U10396 (N_10396,N_9964,N_9833);
and U10397 (N_10397,N_9828,N_9583);
nand U10398 (N_10398,N_9635,N_9774);
xor U10399 (N_10399,N_9768,N_9972);
nand U10400 (N_10400,N_9610,N_9719);
xor U10401 (N_10401,N_9773,N_9511);
and U10402 (N_10402,N_9965,N_9841);
xnor U10403 (N_10403,N_9834,N_9761);
or U10404 (N_10404,N_9581,N_9979);
nor U10405 (N_10405,N_9714,N_9660);
nand U10406 (N_10406,N_9885,N_9916);
and U10407 (N_10407,N_9991,N_9912);
xor U10408 (N_10408,N_9944,N_9926);
xor U10409 (N_10409,N_9900,N_9954);
xnor U10410 (N_10410,N_9676,N_9669);
xor U10411 (N_10411,N_9901,N_9740);
and U10412 (N_10412,N_9988,N_9820);
and U10413 (N_10413,N_9711,N_9527);
xor U10414 (N_10414,N_9919,N_9617);
and U10415 (N_10415,N_9711,N_9508);
or U10416 (N_10416,N_9781,N_9810);
nor U10417 (N_10417,N_9687,N_9919);
nand U10418 (N_10418,N_9973,N_9871);
nand U10419 (N_10419,N_9692,N_9671);
xor U10420 (N_10420,N_9696,N_9763);
nand U10421 (N_10421,N_9552,N_9889);
nor U10422 (N_10422,N_9610,N_9864);
or U10423 (N_10423,N_9527,N_9885);
or U10424 (N_10424,N_9974,N_9774);
nand U10425 (N_10425,N_9818,N_9564);
nand U10426 (N_10426,N_9585,N_9914);
or U10427 (N_10427,N_9848,N_9582);
nor U10428 (N_10428,N_9765,N_9902);
xor U10429 (N_10429,N_9982,N_9894);
xnor U10430 (N_10430,N_9695,N_9946);
nand U10431 (N_10431,N_9595,N_9899);
or U10432 (N_10432,N_9735,N_9760);
nand U10433 (N_10433,N_9609,N_9678);
or U10434 (N_10434,N_9891,N_9905);
and U10435 (N_10435,N_9836,N_9617);
xnor U10436 (N_10436,N_9686,N_9881);
or U10437 (N_10437,N_9971,N_9595);
and U10438 (N_10438,N_9754,N_9954);
or U10439 (N_10439,N_9909,N_9891);
or U10440 (N_10440,N_9966,N_9560);
or U10441 (N_10441,N_9776,N_9632);
and U10442 (N_10442,N_9875,N_9884);
nand U10443 (N_10443,N_9970,N_9609);
xor U10444 (N_10444,N_9730,N_9979);
or U10445 (N_10445,N_9701,N_9509);
nand U10446 (N_10446,N_9546,N_9836);
or U10447 (N_10447,N_9749,N_9779);
nand U10448 (N_10448,N_9528,N_9515);
or U10449 (N_10449,N_9809,N_9840);
nor U10450 (N_10450,N_9852,N_9577);
nand U10451 (N_10451,N_9651,N_9951);
nor U10452 (N_10452,N_9961,N_9585);
nand U10453 (N_10453,N_9618,N_9626);
nand U10454 (N_10454,N_9736,N_9792);
nor U10455 (N_10455,N_9829,N_9630);
xor U10456 (N_10456,N_9900,N_9690);
nor U10457 (N_10457,N_9644,N_9556);
nor U10458 (N_10458,N_9798,N_9892);
and U10459 (N_10459,N_9681,N_9722);
xor U10460 (N_10460,N_9748,N_9895);
xor U10461 (N_10461,N_9991,N_9583);
and U10462 (N_10462,N_9861,N_9537);
or U10463 (N_10463,N_9867,N_9728);
xnor U10464 (N_10464,N_9577,N_9902);
and U10465 (N_10465,N_9798,N_9607);
xnor U10466 (N_10466,N_9884,N_9908);
xnor U10467 (N_10467,N_9592,N_9898);
and U10468 (N_10468,N_9664,N_9674);
nor U10469 (N_10469,N_9878,N_9779);
and U10470 (N_10470,N_9800,N_9647);
nor U10471 (N_10471,N_9643,N_9885);
nand U10472 (N_10472,N_9662,N_9550);
and U10473 (N_10473,N_9604,N_9729);
nor U10474 (N_10474,N_9791,N_9932);
or U10475 (N_10475,N_9554,N_9604);
nor U10476 (N_10476,N_9528,N_9883);
xnor U10477 (N_10477,N_9714,N_9738);
xor U10478 (N_10478,N_9954,N_9882);
and U10479 (N_10479,N_9570,N_9772);
nand U10480 (N_10480,N_9686,N_9927);
nor U10481 (N_10481,N_9794,N_9833);
nand U10482 (N_10482,N_9724,N_9965);
and U10483 (N_10483,N_9965,N_9614);
nor U10484 (N_10484,N_9873,N_9573);
nand U10485 (N_10485,N_9795,N_9935);
nand U10486 (N_10486,N_9704,N_9676);
nor U10487 (N_10487,N_9546,N_9963);
and U10488 (N_10488,N_9938,N_9870);
and U10489 (N_10489,N_9782,N_9750);
nand U10490 (N_10490,N_9831,N_9646);
and U10491 (N_10491,N_9905,N_9873);
and U10492 (N_10492,N_9927,N_9837);
xor U10493 (N_10493,N_9950,N_9657);
nor U10494 (N_10494,N_9914,N_9801);
or U10495 (N_10495,N_9737,N_9826);
xnor U10496 (N_10496,N_9633,N_9761);
xnor U10497 (N_10497,N_9795,N_9532);
nand U10498 (N_10498,N_9896,N_9995);
nand U10499 (N_10499,N_9697,N_9994);
and U10500 (N_10500,N_10130,N_10403);
nor U10501 (N_10501,N_10010,N_10018);
nor U10502 (N_10502,N_10248,N_10094);
or U10503 (N_10503,N_10032,N_10286);
and U10504 (N_10504,N_10292,N_10146);
nor U10505 (N_10505,N_10391,N_10361);
and U10506 (N_10506,N_10468,N_10377);
nand U10507 (N_10507,N_10435,N_10327);
xnor U10508 (N_10508,N_10356,N_10069);
and U10509 (N_10509,N_10229,N_10158);
xor U10510 (N_10510,N_10288,N_10009);
nand U10511 (N_10511,N_10124,N_10054);
nand U10512 (N_10512,N_10352,N_10350);
nor U10513 (N_10513,N_10488,N_10285);
nand U10514 (N_10514,N_10460,N_10154);
or U10515 (N_10515,N_10145,N_10001);
xnor U10516 (N_10516,N_10030,N_10077);
nand U10517 (N_10517,N_10104,N_10021);
or U10518 (N_10518,N_10493,N_10078);
xor U10519 (N_10519,N_10193,N_10392);
and U10520 (N_10520,N_10024,N_10448);
nor U10521 (N_10521,N_10406,N_10422);
nand U10522 (N_10522,N_10036,N_10483);
xor U10523 (N_10523,N_10242,N_10423);
or U10524 (N_10524,N_10125,N_10174);
nand U10525 (N_10525,N_10137,N_10291);
or U10526 (N_10526,N_10050,N_10041);
or U10527 (N_10527,N_10359,N_10026);
and U10528 (N_10528,N_10425,N_10385);
and U10529 (N_10529,N_10357,N_10038);
nand U10530 (N_10530,N_10005,N_10378);
and U10531 (N_10531,N_10322,N_10070);
and U10532 (N_10532,N_10358,N_10340);
xor U10533 (N_10533,N_10366,N_10139);
xnor U10534 (N_10534,N_10035,N_10263);
nand U10535 (N_10535,N_10328,N_10397);
xnor U10536 (N_10536,N_10049,N_10197);
and U10537 (N_10537,N_10179,N_10445);
and U10538 (N_10538,N_10386,N_10341);
nor U10539 (N_10539,N_10266,N_10113);
and U10540 (N_10540,N_10134,N_10310);
xnor U10541 (N_10541,N_10043,N_10096);
nand U10542 (N_10542,N_10478,N_10467);
or U10543 (N_10543,N_10415,N_10167);
xnor U10544 (N_10544,N_10123,N_10066);
nor U10545 (N_10545,N_10244,N_10007);
nand U10546 (N_10546,N_10469,N_10063);
and U10547 (N_10547,N_10017,N_10439);
nand U10548 (N_10548,N_10101,N_10308);
nand U10549 (N_10549,N_10337,N_10162);
xnor U10550 (N_10550,N_10323,N_10354);
xor U10551 (N_10551,N_10087,N_10164);
nor U10552 (N_10552,N_10325,N_10486);
or U10553 (N_10553,N_10264,N_10304);
xnor U10554 (N_10554,N_10080,N_10060);
nand U10555 (N_10555,N_10287,N_10100);
nand U10556 (N_10556,N_10110,N_10349);
or U10557 (N_10557,N_10437,N_10471);
nor U10558 (N_10558,N_10008,N_10099);
nor U10559 (N_10559,N_10331,N_10499);
and U10560 (N_10560,N_10442,N_10417);
nand U10561 (N_10561,N_10213,N_10138);
xor U10562 (N_10562,N_10398,N_10204);
nand U10563 (N_10563,N_10491,N_10321);
nand U10564 (N_10564,N_10275,N_10208);
nand U10565 (N_10565,N_10192,N_10219);
nand U10566 (N_10566,N_10045,N_10128);
and U10567 (N_10567,N_10294,N_10269);
xor U10568 (N_10568,N_10476,N_10053);
xnor U10569 (N_10569,N_10402,N_10132);
nor U10570 (N_10570,N_10481,N_10084);
and U10571 (N_10571,N_10133,N_10334);
nor U10572 (N_10572,N_10474,N_10159);
or U10573 (N_10573,N_10303,N_10025);
nand U10574 (N_10574,N_10450,N_10117);
or U10575 (N_10575,N_10419,N_10072);
nor U10576 (N_10576,N_10245,N_10314);
nand U10577 (N_10577,N_10028,N_10335);
or U10578 (N_10578,N_10367,N_10426);
nand U10579 (N_10579,N_10014,N_10225);
nor U10580 (N_10580,N_10153,N_10176);
nand U10581 (N_10581,N_10458,N_10027);
xor U10582 (N_10582,N_10233,N_10401);
and U10583 (N_10583,N_10037,N_10180);
nand U10584 (N_10584,N_10140,N_10297);
nand U10585 (N_10585,N_10268,N_10424);
nand U10586 (N_10586,N_10163,N_10353);
xor U10587 (N_10587,N_10272,N_10102);
nor U10588 (N_10588,N_10383,N_10156);
nor U10589 (N_10589,N_10231,N_10372);
and U10590 (N_10590,N_10347,N_10108);
xnor U10591 (N_10591,N_10393,N_10190);
nor U10592 (N_10592,N_10195,N_10273);
nand U10593 (N_10593,N_10236,N_10224);
and U10594 (N_10594,N_10056,N_10409);
and U10595 (N_10595,N_10183,N_10047);
nor U10596 (N_10596,N_10355,N_10243);
xor U10597 (N_10597,N_10451,N_10390);
nor U10598 (N_10598,N_10251,N_10332);
or U10599 (N_10599,N_10440,N_10370);
and U10600 (N_10600,N_10112,N_10387);
nor U10601 (N_10601,N_10492,N_10170);
nor U10602 (N_10602,N_10345,N_10189);
and U10603 (N_10603,N_10414,N_10147);
xor U10604 (N_10604,N_10067,N_10057);
nor U10605 (N_10605,N_10295,N_10438);
or U10606 (N_10606,N_10201,N_10453);
or U10607 (N_10607,N_10166,N_10121);
nand U10608 (N_10608,N_10120,N_10033);
or U10609 (N_10609,N_10324,N_10346);
and U10610 (N_10610,N_10342,N_10211);
or U10611 (N_10611,N_10181,N_10305);
nor U10612 (N_10612,N_10062,N_10296);
xor U10613 (N_10613,N_10301,N_10312);
xor U10614 (N_10614,N_10384,N_10118);
or U10615 (N_10615,N_10022,N_10092);
nor U10616 (N_10616,N_10237,N_10215);
nor U10617 (N_10617,N_10119,N_10441);
or U10618 (N_10618,N_10234,N_10299);
and U10619 (N_10619,N_10200,N_10226);
nand U10620 (N_10620,N_10380,N_10116);
nand U10621 (N_10621,N_10326,N_10319);
and U10622 (N_10622,N_10052,N_10184);
nand U10623 (N_10623,N_10114,N_10498);
or U10624 (N_10624,N_10457,N_10316);
nand U10625 (N_10625,N_10465,N_10240);
or U10626 (N_10626,N_10186,N_10279);
xor U10627 (N_10627,N_10191,N_10065);
or U10628 (N_10628,N_10339,N_10443);
nand U10629 (N_10629,N_10489,N_10048);
and U10630 (N_10630,N_10004,N_10046);
and U10631 (N_10631,N_10088,N_10259);
nor U10632 (N_10632,N_10461,N_10472);
nor U10633 (N_10633,N_10430,N_10407);
xnor U10634 (N_10634,N_10280,N_10462);
nand U10635 (N_10635,N_10011,N_10320);
nand U10636 (N_10636,N_10330,N_10307);
nand U10637 (N_10637,N_10455,N_10157);
xor U10638 (N_10638,N_10408,N_10188);
or U10639 (N_10639,N_10029,N_10362);
xor U10640 (N_10640,N_10012,N_10459);
nor U10641 (N_10641,N_10228,N_10329);
xor U10642 (N_10642,N_10389,N_10013);
and U10643 (N_10643,N_10484,N_10253);
and U10644 (N_10644,N_10115,N_10371);
nor U10645 (N_10645,N_10106,N_10098);
or U10646 (N_10646,N_10250,N_10388);
xnor U10647 (N_10647,N_10238,N_10428);
nand U10648 (N_10648,N_10196,N_10381);
nor U10649 (N_10649,N_10351,N_10434);
and U10650 (N_10650,N_10107,N_10207);
nand U10651 (N_10651,N_10271,N_10141);
and U10652 (N_10652,N_10126,N_10258);
or U10653 (N_10653,N_10071,N_10464);
and U10654 (N_10654,N_10494,N_10475);
and U10655 (N_10655,N_10374,N_10270);
xnor U10656 (N_10656,N_10416,N_10187);
nor U10657 (N_10657,N_10223,N_10218);
and U10658 (N_10658,N_10427,N_10410);
or U10659 (N_10659,N_10477,N_10260);
nand U10660 (N_10660,N_10293,N_10436);
or U10661 (N_10661,N_10160,N_10040);
xnor U10662 (N_10662,N_10306,N_10411);
xnor U10663 (N_10663,N_10470,N_10143);
nand U10664 (N_10664,N_10122,N_10252);
and U10665 (N_10665,N_10148,N_10487);
nor U10666 (N_10666,N_10210,N_10479);
xor U10667 (N_10667,N_10379,N_10344);
and U10668 (N_10668,N_10485,N_10421);
nand U10669 (N_10669,N_10282,N_10198);
and U10670 (N_10670,N_10267,N_10221);
and U10671 (N_10671,N_10175,N_10151);
xnor U10672 (N_10672,N_10375,N_10463);
nand U10673 (N_10673,N_10220,N_10290);
nand U10674 (N_10674,N_10097,N_10480);
nand U10675 (N_10675,N_10418,N_10311);
or U10676 (N_10676,N_10222,N_10149);
or U10677 (N_10677,N_10278,N_10168);
and U10678 (N_10678,N_10254,N_10336);
nand U10679 (N_10679,N_10034,N_10194);
xnor U10680 (N_10680,N_10249,N_10111);
nand U10681 (N_10681,N_10216,N_10274);
and U10682 (N_10682,N_10109,N_10203);
nand U10683 (N_10683,N_10085,N_10083);
or U10684 (N_10684,N_10217,N_10169);
nor U10685 (N_10685,N_10042,N_10456);
xor U10686 (N_10686,N_10142,N_10413);
nor U10687 (N_10687,N_10338,N_10079);
xor U10688 (N_10688,N_10230,N_10348);
nand U10689 (N_10689,N_10241,N_10039);
xor U10690 (N_10690,N_10093,N_10343);
nand U10691 (N_10691,N_10182,N_10281);
and U10692 (N_10692,N_10400,N_10006);
nand U10693 (N_10693,N_10257,N_10232);
or U10694 (N_10694,N_10177,N_10202);
or U10695 (N_10695,N_10076,N_10432);
and U10696 (N_10696,N_10064,N_10394);
and U10697 (N_10697,N_10497,N_10382);
nand U10698 (N_10698,N_10444,N_10061);
and U10699 (N_10699,N_10089,N_10256);
and U10700 (N_10700,N_10373,N_10205);
nor U10701 (N_10701,N_10317,N_10129);
and U10702 (N_10702,N_10276,N_10090);
xnor U10703 (N_10703,N_10300,N_10496);
nand U10704 (N_10704,N_10412,N_10454);
nor U10705 (N_10705,N_10068,N_10212);
nand U10706 (N_10706,N_10262,N_10227);
nor U10707 (N_10707,N_10135,N_10150);
nor U10708 (N_10708,N_10309,N_10058);
xor U10709 (N_10709,N_10405,N_10003);
xnor U10710 (N_10710,N_10247,N_10433);
nand U10711 (N_10711,N_10482,N_10277);
nor U10712 (N_10712,N_10265,N_10395);
or U10713 (N_10713,N_10446,N_10452);
or U10714 (N_10714,N_10173,N_10165);
xnor U10715 (N_10715,N_10246,N_10074);
nor U10716 (N_10716,N_10131,N_10044);
nor U10717 (N_10717,N_10073,N_10155);
or U10718 (N_10718,N_10368,N_10209);
and U10719 (N_10719,N_10144,N_10081);
and U10720 (N_10720,N_10283,N_10313);
or U10721 (N_10721,N_10429,N_10161);
nor U10722 (N_10722,N_10095,N_10495);
and U10723 (N_10723,N_10086,N_10015);
nand U10724 (N_10724,N_10214,N_10399);
or U10725 (N_10725,N_10082,N_10051);
nand U10726 (N_10726,N_10261,N_10365);
or U10727 (N_10727,N_10055,N_10447);
and U10728 (N_10728,N_10364,N_10023);
nand U10729 (N_10729,N_10376,N_10420);
and U10730 (N_10730,N_10103,N_10431);
xor U10731 (N_10731,N_10473,N_10136);
nor U10732 (N_10732,N_10369,N_10333);
nand U10733 (N_10733,N_10178,N_10315);
nand U10734 (N_10734,N_10185,N_10127);
and U10735 (N_10735,N_10002,N_10031);
nor U10736 (N_10736,N_10000,N_10363);
xnor U10737 (N_10737,N_10152,N_10302);
nor U10738 (N_10738,N_10235,N_10020);
or U10739 (N_10739,N_10019,N_10075);
xor U10740 (N_10740,N_10091,N_10059);
nand U10741 (N_10741,N_10404,N_10105);
nor U10742 (N_10742,N_10490,N_10206);
or U10743 (N_10743,N_10289,N_10199);
and U10744 (N_10744,N_10171,N_10016);
and U10745 (N_10745,N_10172,N_10298);
or U10746 (N_10746,N_10255,N_10284);
or U10747 (N_10747,N_10239,N_10466);
or U10748 (N_10748,N_10449,N_10318);
and U10749 (N_10749,N_10396,N_10360);
nor U10750 (N_10750,N_10376,N_10138);
and U10751 (N_10751,N_10463,N_10498);
nand U10752 (N_10752,N_10015,N_10133);
nor U10753 (N_10753,N_10217,N_10478);
or U10754 (N_10754,N_10330,N_10147);
xor U10755 (N_10755,N_10265,N_10427);
nand U10756 (N_10756,N_10155,N_10257);
nor U10757 (N_10757,N_10476,N_10195);
nand U10758 (N_10758,N_10239,N_10218);
nor U10759 (N_10759,N_10462,N_10432);
or U10760 (N_10760,N_10324,N_10129);
nand U10761 (N_10761,N_10298,N_10023);
xnor U10762 (N_10762,N_10303,N_10343);
nor U10763 (N_10763,N_10366,N_10306);
or U10764 (N_10764,N_10157,N_10234);
and U10765 (N_10765,N_10418,N_10206);
nor U10766 (N_10766,N_10260,N_10367);
xor U10767 (N_10767,N_10055,N_10105);
and U10768 (N_10768,N_10105,N_10204);
nand U10769 (N_10769,N_10260,N_10248);
nor U10770 (N_10770,N_10066,N_10250);
and U10771 (N_10771,N_10047,N_10218);
nor U10772 (N_10772,N_10460,N_10434);
xor U10773 (N_10773,N_10402,N_10459);
nor U10774 (N_10774,N_10230,N_10461);
xnor U10775 (N_10775,N_10402,N_10012);
nor U10776 (N_10776,N_10483,N_10104);
or U10777 (N_10777,N_10364,N_10471);
nand U10778 (N_10778,N_10237,N_10179);
nor U10779 (N_10779,N_10327,N_10351);
nor U10780 (N_10780,N_10365,N_10173);
nor U10781 (N_10781,N_10374,N_10260);
and U10782 (N_10782,N_10398,N_10381);
nor U10783 (N_10783,N_10243,N_10453);
nand U10784 (N_10784,N_10366,N_10207);
and U10785 (N_10785,N_10458,N_10409);
or U10786 (N_10786,N_10142,N_10371);
xnor U10787 (N_10787,N_10463,N_10011);
nand U10788 (N_10788,N_10243,N_10315);
or U10789 (N_10789,N_10239,N_10047);
xnor U10790 (N_10790,N_10394,N_10018);
or U10791 (N_10791,N_10359,N_10463);
nor U10792 (N_10792,N_10439,N_10422);
or U10793 (N_10793,N_10399,N_10255);
or U10794 (N_10794,N_10414,N_10053);
nor U10795 (N_10795,N_10480,N_10439);
or U10796 (N_10796,N_10411,N_10010);
xor U10797 (N_10797,N_10068,N_10472);
xor U10798 (N_10798,N_10289,N_10304);
xnor U10799 (N_10799,N_10411,N_10260);
or U10800 (N_10800,N_10439,N_10483);
xor U10801 (N_10801,N_10474,N_10162);
xor U10802 (N_10802,N_10391,N_10316);
and U10803 (N_10803,N_10314,N_10187);
or U10804 (N_10804,N_10278,N_10406);
and U10805 (N_10805,N_10265,N_10309);
nor U10806 (N_10806,N_10455,N_10268);
nor U10807 (N_10807,N_10118,N_10387);
nor U10808 (N_10808,N_10287,N_10106);
or U10809 (N_10809,N_10290,N_10090);
and U10810 (N_10810,N_10492,N_10261);
nor U10811 (N_10811,N_10124,N_10203);
xor U10812 (N_10812,N_10361,N_10182);
or U10813 (N_10813,N_10382,N_10016);
or U10814 (N_10814,N_10414,N_10127);
nor U10815 (N_10815,N_10399,N_10175);
and U10816 (N_10816,N_10447,N_10451);
xnor U10817 (N_10817,N_10287,N_10007);
xnor U10818 (N_10818,N_10302,N_10037);
or U10819 (N_10819,N_10003,N_10051);
nor U10820 (N_10820,N_10022,N_10224);
or U10821 (N_10821,N_10258,N_10182);
xor U10822 (N_10822,N_10163,N_10304);
and U10823 (N_10823,N_10466,N_10245);
xor U10824 (N_10824,N_10288,N_10446);
and U10825 (N_10825,N_10387,N_10074);
nor U10826 (N_10826,N_10141,N_10063);
and U10827 (N_10827,N_10192,N_10100);
or U10828 (N_10828,N_10290,N_10408);
nor U10829 (N_10829,N_10004,N_10373);
xnor U10830 (N_10830,N_10405,N_10217);
and U10831 (N_10831,N_10198,N_10068);
and U10832 (N_10832,N_10336,N_10067);
nand U10833 (N_10833,N_10033,N_10337);
xnor U10834 (N_10834,N_10346,N_10278);
or U10835 (N_10835,N_10367,N_10148);
nand U10836 (N_10836,N_10486,N_10028);
nand U10837 (N_10837,N_10427,N_10376);
nor U10838 (N_10838,N_10181,N_10046);
nor U10839 (N_10839,N_10462,N_10416);
xnor U10840 (N_10840,N_10413,N_10268);
nand U10841 (N_10841,N_10074,N_10232);
nand U10842 (N_10842,N_10196,N_10262);
xor U10843 (N_10843,N_10237,N_10299);
or U10844 (N_10844,N_10125,N_10294);
or U10845 (N_10845,N_10064,N_10166);
and U10846 (N_10846,N_10118,N_10122);
xor U10847 (N_10847,N_10305,N_10000);
xor U10848 (N_10848,N_10240,N_10093);
nand U10849 (N_10849,N_10035,N_10290);
nand U10850 (N_10850,N_10376,N_10100);
nor U10851 (N_10851,N_10469,N_10306);
nor U10852 (N_10852,N_10094,N_10383);
xnor U10853 (N_10853,N_10372,N_10396);
and U10854 (N_10854,N_10162,N_10150);
and U10855 (N_10855,N_10317,N_10384);
xnor U10856 (N_10856,N_10416,N_10365);
nor U10857 (N_10857,N_10420,N_10388);
nand U10858 (N_10858,N_10067,N_10395);
nor U10859 (N_10859,N_10066,N_10343);
xor U10860 (N_10860,N_10338,N_10248);
or U10861 (N_10861,N_10146,N_10389);
or U10862 (N_10862,N_10447,N_10352);
nand U10863 (N_10863,N_10339,N_10277);
and U10864 (N_10864,N_10018,N_10159);
and U10865 (N_10865,N_10398,N_10308);
or U10866 (N_10866,N_10197,N_10126);
and U10867 (N_10867,N_10075,N_10174);
or U10868 (N_10868,N_10271,N_10105);
and U10869 (N_10869,N_10356,N_10491);
nor U10870 (N_10870,N_10096,N_10469);
xnor U10871 (N_10871,N_10007,N_10236);
and U10872 (N_10872,N_10078,N_10162);
and U10873 (N_10873,N_10082,N_10436);
nand U10874 (N_10874,N_10257,N_10136);
xnor U10875 (N_10875,N_10405,N_10013);
nor U10876 (N_10876,N_10082,N_10143);
nor U10877 (N_10877,N_10108,N_10155);
nor U10878 (N_10878,N_10145,N_10417);
and U10879 (N_10879,N_10438,N_10431);
xnor U10880 (N_10880,N_10016,N_10114);
and U10881 (N_10881,N_10267,N_10270);
xnor U10882 (N_10882,N_10217,N_10399);
or U10883 (N_10883,N_10011,N_10493);
or U10884 (N_10884,N_10214,N_10029);
nor U10885 (N_10885,N_10437,N_10320);
xor U10886 (N_10886,N_10459,N_10359);
nand U10887 (N_10887,N_10245,N_10216);
xnor U10888 (N_10888,N_10110,N_10249);
nand U10889 (N_10889,N_10360,N_10113);
or U10890 (N_10890,N_10302,N_10139);
nor U10891 (N_10891,N_10415,N_10346);
nand U10892 (N_10892,N_10080,N_10082);
or U10893 (N_10893,N_10252,N_10400);
xor U10894 (N_10894,N_10186,N_10188);
or U10895 (N_10895,N_10448,N_10228);
xnor U10896 (N_10896,N_10342,N_10222);
or U10897 (N_10897,N_10166,N_10323);
and U10898 (N_10898,N_10370,N_10377);
or U10899 (N_10899,N_10093,N_10018);
and U10900 (N_10900,N_10217,N_10302);
or U10901 (N_10901,N_10380,N_10062);
nor U10902 (N_10902,N_10162,N_10347);
nand U10903 (N_10903,N_10203,N_10316);
xor U10904 (N_10904,N_10302,N_10170);
nand U10905 (N_10905,N_10187,N_10165);
xnor U10906 (N_10906,N_10073,N_10283);
nor U10907 (N_10907,N_10260,N_10099);
and U10908 (N_10908,N_10100,N_10498);
and U10909 (N_10909,N_10063,N_10087);
xor U10910 (N_10910,N_10489,N_10078);
and U10911 (N_10911,N_10280,N_10176);
and U10912 (N_10912,N_10212,N_10485);
or U10913 (N_10913,N_10360,N_10333);
nand U10914 (N_10914,N_10083,N_10229);
and U10915 (N_10915,N_10417,N_10453);
xnor U10916 (N_10916,N_10288,N_10390);
and U10917 (N_10917,N_10037,N_10301);
and U10918 (N_10918,N_10393,N_10497);
or U10919 (N_10919,N_10280,N_10097);
nor U10920 (N_10920,N_10338,N_10349);
or U10921 (N_10921,N_10210,N_10417);
and U10922 (N_10922,N_10419,N_10409);
or U10923 (N_10923,N_10462,N_10463);
nand U10924 (N_10924,N_10365,N_10357);
or U10925 (N_10925,N_10424,N_10022);
xnor U10926 (N_10926,N_10224,N_10181);
nor U10927 (N_10927,N_10210,N_10444);
nand U10928 (N_10928,N_10141,N_10090);
xor U10929 (N_10929,N_10302,N_10241);
and U10930 (N_10930,N_10184,N_10243);
or U10931 (N_10931,N_10270,N_10430);
nor U10932 (N_10932,N_10045,N_10375);
and U10933 (N_10933,N_10147,N_10304);
and U10934 (N_10934,N_10001,N_10058);
and U10935 (N_10935,N_10341,N_10243);
nor U10936 (N_10936,N_10357,N_10077);
and U10937 (N_10937,N_10324,N_10472);
nand U10938 (N_10938,N_10149,N_10331);
nand U10939 (N_10939,N_10160,N_10058);
nor U10940 (N_10940,N_10038,N_10456);
xor U10941 (N_10941,N_10009,N_10282);
xor U10942 (N_10942,N_10180,N_10322);
or U10943 (N_10943,N_10350,N_10269);
nand U10944 (N_10944,N_10304,N_10478);
nor U10945 (N_10945,N_10304,N_10459);
xor U10946 (N_10946,N_10080,N_10028);
or U10947 (N_10947,N_10381,N_10414);
xnor U10948 (N_10948,N_10147,N_10044);
and U10949 (N_10949,N_10488,N_10240);
nand U10950 (N_10950,N_10308,N_10471);
and U10951 (N_10951,N_10371,N_10311);
or U10952 (N_10952,N_10319,N_10004);
or U10953 (N_10953,N_10282,N_10096);
nor U10954 (N_10954,N_10214,N_10174);
or U10955 (N_10955,N_10223,N_10422);
or U10956 (N_10956,N_10425,N_10138);
and U10957 (N_10957,N_10020,N_10301);
nand U10958 (N_10958,N_10364,N_10104);
nand U10959 (N_10959,N_10118,N_10038);
xnor U10960 (N_10960,N_10066,N_10197);
xor U10961 (N_10961,N_10488,N_10341);
or U10962 (N_10962,N_10179,N_10146);
xnor U10963 (N_10963,N_10101,N_10003);
or U10964 (N_10964,N_10336,N_10043);
or U10965 (N_10965,N_10420,N_10097);
xnor U10966 (N_10966,N_10080,N_10374);
and U10967 (N_10967,N_10295,N_10431);
or U10968 (N_10968,N_10433,N_10248);
nand U10969 (N_10969,N_10346,N_10420);
and U10970 (N_10970,N_10122,N_10093);
xor U10971 (N_10971,N_10326,N_10059);
nand U10972 (N_10972,N_10090,N_10374);
and U10973 (N_10973,N_10330,N_10440);
nor U10974 (N_10974,N_10344,N_10390);
or U10975 (N_10975,N_10297,N_10132);
and U10976 (N_10976,N_10079,N_10398);
nand U10977 (N_10977,N_10014,N_10392);
nand U10978 (N_10978,N_10372,N_10206);
and U10979 (N_10979,N_10052,N_10337);
xnor U10980 (N_10980,N_10126,N_10388);
nor U10981 (N_10981,N_10076,N_10158);
or U10982 (N_10982,N_10029,N_10197);
and U10983 (N_10983,N_10050,N_10344);
xor U10984 (N_10984,N_10453,N_10266);
and U10985 (N_10985,N_10283,N_10124);
and U10986 (N_10986,N_10459,N_10286);
nand U10987 (N_10987,N_10253,N_10383);
and U10988 (N_10988,N_10232,N_10197);
xor U10989 (N_10989,N_10118,N_10258);
and U10990 (N_10990,N_10089,N_10230);
or U10991 (N_10991,N_10283,N_10293);
nand U10992 (N_10992,N_10176,N_10317);
xor U10993 (N_10993,N_10433,N_10246);
and U10994 (N_10994,N_10124,N_10207);
nand U10995 (N_10995,N_10065,N_10120);
nor U10996 (N_10996,N_10137,N_10005);
nand U10997 (N_10997,N_10484,N_10130);
nor U10998 (N_10998,N_10495,N_10145);
nand U10999 (N_10999,N_10251,N_10392);
nor U11000 (N_11000,N_10887,N_10915);
xor U11001 (N_11001,N_10654,N_10787);
nand U11002 (N_11002,N_10619,N_10753);
nand U11003 (N_11003,N_10940,N_10867);
nor U11004 (N_11004,N_10873,N_10883);
or U11005 (N_11005,N_10569,N_10895);
and U11006 (N_11006,N_10502,N_10960);
nor U11007 (N_11007,N_10522,N_10967);
and U11008 (N_11008,N_10637,N_10585);
nor U11009 (N_11009,N_10956,N_10570);
nor U11010 (N_11010,N_10648,N_10812);
and U11011 (N_11011,N_10652,N_10731);
nand U11012 (N_11012,N_10545,N_10728);
or U11013 (N_11013,N_10732,N_10508);
and U11014 (N_11014,N_10893,N_10532);
nand U11015 (N_11015,N_10699,N_10751);
nor U11016 (N_11016,N_10938,N_10797);
xor U11017 (N_11017,N_10922,N_10771);
xnor U11018 (N_11018,N_10607,N_10580);
or U11019 (N_11019,N_10818,N_10576);
nor U11020 (N_11020,N_10624,N_10941);
nor U11021 (N_11021,N_10840,N_10602);
nor U11022 (N_11022,N_10593,N_10944);
and U11023 (N_11023,N_10558,N_10513);
and U11024 (N_11024,N_10655,N_10662);
xor U11025 (N_11025,N_10843,N_10889);
and U11026 (N_11026,N_10746,N_10794);
and U11027 (N_11027,N_10671,N_10703);
nor U11028 (N_11028,N_10519,N_10788);
or U11029 (N_11029,N_10864,N_10804);
nor U11030 (N_11030,N_10733,N_10988);
xor U11031 (N_11031,N_10600,N_10912);
and U11032 (N_11032,N_10505,N_10695);
nor U11033 (N_11033,N_10852,N_10793);
xnor U11034 (N_11034,N_10808,N_10782);
xor U11035 (N_11035,N_10752,N_10589);
xor U11036 (N_11036,N_10716,N_10924);
or U11037 (N_11037,N_10996,N_10884);
or U11038 (N_11038,N_10875,N_10528);
nor U11039 (N_11039,N_10544,N_10838);
xnor U11040 (N_11040,N_10575,N_10772);
and U11041 (N_11041,N_10696,N_10994);
nor U11042 (N_11042,N_10972,N_10830);
nand U11043 (N_11043,N_10786,N_10650);
and U11044 (N_11044,N_10835,N_10869);
and U11045 (N_11045,N_10621,N_10574);
and U11046 (N_11046,N_10891,N_10809);
xnor U11047 (N_11047,N_10937,N_10507);
nand U11048 (N_11048,N_10791,N_10849);
nand U11049 (N_11049,N_10511,N_10689);
or U11050 (N_11050,N_10634,N_10641);
nor U11051 (N_11051,N_10820,N_10706);
xnor U11052 (N_11052,N_10881,N_10712);
xor U11053 (N_11053,N_10659,N_10720);
nand U11054 (N_11054,N_10799,N_10853);
xnor U11055 (N_11055,N_10845,N_10743);
nor U11056 (N_11056,N_10635,N_10737);
nand U11057 (N_11057,N_10890,N_10504);
nor U11058 (N_11058,N_10563,N_10954);
and U11059 (N_11059,N_10568,N_10773);
xnor U11060 (N_11060,N_10640,N_10935);
nor U11061 (N_11061,N_10665,N_10928);
nand U11062 (N_11062,N_10714,N_10827);
nor U11063 (N_11063,N_10630,N_10780);
nor U11064 (N_11064,N_10829,N_10584);
xor U11065 (N_11065,N_10821,N_10581);
or U11066 (N_11066,N_10586,N_10817);
nor U11067 (N_11067,N_10863,N_10579);
and U11068 (N_11068,N_10969,N_10717);
and U11069 (N_11069,N_10801,N_10764);
and U11070 (N_11070,N_10792,N_10595);
or U11071 (N_11071,N_10567,N_10930);
nor U11072 (N_11072,N_10936,N_10984);
nor U11073 (N_11073,N_10625,N_10949);
or U11074 (N_11074,N_10931,N_10880);
or U11075 (N_11075,N_10847,N_10987);
xor U11076 (N_11076,N_10705,N_10813);
nand U11077 (N_11077,N_10697,N_10747);
nand U11078 (N_11078,N_10521,N_10533);
and U11079 (N_11079,N_10514,N_10601);
nand U11080 (N_11080,N_10701,N_10748);
xnor U11081 (N_11081,N_10779,N_10740);
xnor U11082 (N_11082,N_10605,N_10768);
or U11083 (N_11083,N_10530,N_10707);
nand U11084 (N_11084,N_10932,N_10815);
nor U11085 (N_11085,N_10834,N_10738);
nand U11086 (N_11086,N_10807,N_10571);
nand U11087 (N_11087,N_10842,N_10620);
nor U11088 (N_11088,N_10672,N_10859);
xnor U11089 (N_11089,N_10814,N_10865);
and U11090 (N_11090,N_10874,N_10680);
xnor U11091 (N_11091,N_10550,N_10661);
nand U11092 (N_11092,N_10850,N_10905);
nor U11093 (N_11093,N_10965,N_10831);
and U11094 (N_11094,N_10908,N_10796);
or U11095 (N_11095,N_10693,N_10757);
nor U11096 (N_11096,N_10934,N_10633);
nand U11097 (N_11097,N_10876,N_10599);
and U11098 (N_11098,N_10755,N_10683);
or U11099 (N_11099,N_10682,N_10603);
nor U11100 (N_11100,N_10559,N_10989);
xor U11101 (N_11101,N_10911,N_10719);
or U11102 (N_11102,N_10708,N_10674);
xnor U11103 (N_11103,N_10704,N_10962);
and U11104 (N_11104,N_10841,N_10750);
nand U11105 (N_11105,N_10577,N_10933);
nor U11106 (N_11106,N_10778,N_10617);
nor U11107 (N_11107,N_10877,N_10993);
xnor U11108 (N_11108,N_10698,N_10610);
or U11109 (N_11109,N_10596,N_10973);
or U11110 (N_11110,N_10822,N_10556);
nand U11111 (N_11111,N_10702,N_10598);
or U11112 (N_11112,N_10977,N_10686);
or U11113 (N_11113,N_10961,N_10552);
or U11114 (N_11114,N_10770,N_10744);
nand U11115 (N_11115,N_10756,N_10979);
and U11116 (N_11116,N_10819,N_10958);
and U11117 (N_11117,N_10673,N_10690);
xnor U11118 (N_11118,N_10647,N_10613);
xnor U11119 (N_11119,N_10515,N_10542);
nand U11120 (N_11120,N_10668,N_10562);
or U11121 (N_11121,N_10612,N_10846);
nand U11122 (N_11122,N_10871,N_10675);
nor U11123 (N_11123,N_10543,N_10774);
xnor U11124 (N_11124,N_10734,N_10509);
or U11125 (N_11125,N_10629,N_10651);
nor U11126 (N_11126,N_10526,N_10622);
and U11127 (N_11127,N_10836,N_10573);
and U11128 (N_11128,N_10833,N_10541);
and U11129 (N_11129,N_10649,N_10646);
or U11130 (N_11130,N_10857,N_10946);
nor U11131 (N_11131,N_10520,N_10991);
or U11132 (N_11132,N_10534,N_10798);
nand U11133 (N_11133,N_10644,N_10909);
xnor U11134 (N_11134,N_10529,N_10806);
nor U11135 (N_11135,N_10614,N_10828);
nor U11136 (N_11136,N_10826,N_10844);
nand U11137 (N_11137,N_10759,N_10945);
and U11138 (N_11138,N_10546,N_10766);
and U11139 (N_11139,N_10561,N_10862);
or U11140 (N_11140,N_10523,N_10992);
or U11141 (N_11141,N_10892,N_10726);
or U11142 (N_11142,N_10762,N_10555);
nor U11143 (N_11143,N_10872,N_10676);
nand U11144 (N_11144,N_10926,N_10564);
nor U11145 (N_11145,N_10653,N_10710);
and U11146 (N_11146,N_10525,N_10692);
nor U11147 (N_11147,N_10899,N_10777);
nor U11148 (N_11148,N_10642,N_10512);
nor U11149 (N_11149,N_10506,N_10951);
or U11150 (N_11150,N_10975,N_10535);
nor U11151 (N_11151,N_10837,N_10623);
and U11152 (N_11152,N_10725,N_10832);
xor U11153 (N_11153,N_10735,N_10709);
or U11154 (N_11154,N_10615,N_10700);
nor U11155 (N_11155,N_10897,N_10914);
or U11156 (N_11156,N_10611,N_10670);
nand U11157 (N_11157,N_10885,N_10667);
xnor U11158 (N_11158,N_10549,N_10959);
or U11159 (N_11159,N_10723,N_10587);
xor U11160 (N_11160,N_10636,N_10910);
nor U11161 (N_11161,N_10594,N_10628);
nand U11162 (N_11162,N_10810,N_10886);
xor U11163 (N_11163,N_10982,N_10694);
and U11164 (N_11164,N_10904,N_10921);
xor U11165 (N_11165,N_10537,N_10663);
or U11166 (N_11166,N_10964,N_10816);
nand U11167 (N_11167,N_10868,N_10824);
nand U11168 (N_11168,N_10953,N_10627);
or U11169 (N_11169,N_10551,N_10785);
or U11170 (N_11170,N_10981,N_10531);
nor U11171 (N_11171,N_10974,N_10896);
nor U11172 (N_11172,N_10554,N_10998);
nand U11173 (N_11173,N_10729,N_10741);
nand U11174 (N_11174,N_10583,N_10966);
xnor U11175 (N_11175,N_10643,N_10848);
nand U11176 (N_11176,N_10855,N_10894);
nand U11177 (N_11177,N_10727,N_10803);
nor U11178 (N_11178,N_10986,N_10898);
and U11179 (N_11179,N_10811,N_10538);
xor U11180 (N_11180,N_10769,N_10524);
xor U11181 (N_11181,N_10913,N_10645);
xnor U11182 (N_11182,N_10767,N_10968);
nor U11183 (N_11183,N_10547,N_10781);
or U11184 (N_11184,N_10681,N_10618);
nor U11185 (N_11185,N_10919,N_10878);
nor U11186 (N_11186,N_10608,N_10970);
nand U11187 (N_11187,N_10632,N_10943);
and U11188 (N_11188,N_10666,N_10678);
or U11189 (N_11189,N_10906,N_10939);
nand U11190 (N_11190,N_10501,N_10963);
nand U11191 (N_11191,N_10656,N_10660);
nor U11192 (N_11192,N_10825,N_10997);
and U11193 (N_11193,N_10858,N_10900);
nand U11194 (N_11194,N_10925,N_10687);
and U11195 (N_11195,N_10664,N_10510);
or U11196 (N_11196,N_10592,N_10578);
nor U11197 (N_11197,N_10917,N_10783);
xnor U11198 (N_11198,N_10518,N_10861);
xor U11199 (N_11199,N_10823,N_10918);
xor U11200 (N_11200,N_10980,N_10742);
or U11201 (N_11201,N_10999,N_10761);
nor U11202 (N_11202,N_10718,N_10609);
nor U11203 (N_11203,N_10950,N_10947);
and U11204 (N_11204,N_10749,N_10800);
and U11205 (N_11205,N_10923,N_10606);
nor U11206 (N_11206,N_10669,N_10775);
nand U11207 (N_11207,N_10776,N_10948);
or U11208 (N_11208,N_10907,N_10685);
nor U11209 (N_11209,N_10548,N_10839);
xnor U11210 (N_11210,N_10553,N_10860);
nand U11211 (N_11211,N_10715,N_10721);
or U11212 (N_11212,N_10978,N_10745);
xnor U11213 (N_11213,N_10888,N_10902);
nor U11214 (N_11214,N_10955,N_10527);
xnor U11215 (N_11215,N_10597,N_10503);
and U11216 (N_11216,N_10572,N_10638);
xor U11217 (N_11217,N_10679,N_10856);
nor U11218 (N_11218,N_10730,N_10851);
or U11219 (N_11219,N_10976,N_10626);
and U11220 (N_11220,N_10582,N_10657);
xor U11221 (N_11221,N_10983,N_10631);
nor U11222 (N_11222,N_10539,N_10942);
xnor U11223 (N_11223,N_10879,N_10739);
and U11224 (N_11224,N_10736,N_10557);
or U11225 (N_11225,N_10517,N_10802);
and U11226 (N_11226,N_10684,N_10540);
and U11227 (N_11227,N_10560,N_10927);
nand U11228 (N_11228,N_10536,N_10870);
xnor U11229 (N_11229,N_10591,N_10903);
xnor U11230 (N_11230,N_10795,N_10758);
or U11231 (N_11231,N_10985,N_10588);
and U11232 (N_11232,N_10995,N_10854);
and U11233 (N_11233,N_10957,N_10500);
and U11234 (N_11234,N_10590,N_10566);
nor U11235 (N_11235,N_10866,N_10916);
nand U11236 (N_11236,N_10565,N_10990);
nor U11237 (N_11237,N_10604,N_10790);
nand U11238 (N_11238,N_10929,N_10971);
and U11239 (N_11239,N_10754,N_10516);
nand U11240 (N_11240,N_10920,N_10805);
nand U11241 (N_11241,N_10713,N_10691);
xor U11242 (N_11242,N_10677,N_10722);
nand U11243 (N_11243,N_10784,N_10901);
xor U11244 (N_11244,N_10789,N_10763);
nor U11245 (N_11245,N_10724,N_10765);
and U11246 (N_11246,N_10711,N_10760);
nor U11247 (N_11247,N_10688,N_10658);
nor U11248 (N_11248,N_10882,N_10952);
or U11249 (N_11249,N_10639,N_10616);
nand U11250 (N_11250,N_10871,N_10961);
nand U11251 (N_11251,N_10605,N_10977);
and U11252 (N_11252,N_10831,N_10526);
nor U11253 (N_11253,N_10541,N_10826);
and U11254 (N_11254,N_10699,N_10816);
xor U11255 (N_11255,N_10802,N_10928);
and U11256 (N_11256,N_10769,N_10613);
and U11257 (N_11257,N_10580,N_10836);
nor U11258 (N_11258,N_10593,N_10760);
or U11259 (N_11259,N_10863,N_10587);
and U11260 (N_11260,N_10597,N_10909);
nand U11261 (N_11261,N_10628,N_10959);
or U11262 (N_11262,N_10809,N_10652);
nor U11263 (N_11263,N_10524,N_10652);
or U11264 (N_11264,N_10909,N_10984);
and U11265 (N_11265,N_10875,N_10816);
nand U11266 (N_11266,N_10661,N_10949);
nor U11267 (N_11267,N_10910,N_10799);
and U11268 (N_11268,N_10506,N_10829);
or U11269 (N_11269,N_10664,N_10993);
or U11270 (N_11270,N_10652,N_10862);
xnor U11271 (N_11271,N_10847,N_10672);
and U11272 (N_11272,N_10960,N_10677);
nand U11273 (N_11273,N_10785,N_10848);
and U11274 (N_11274,N_10942,N_10637);
xor U11275 (N_11275,N_10872,N_10730);
and U11276 (N_11276,N_10933,N_10946);
or U11277 (N_11277,N_10536,N_10902);
xor U11278 (N_11278,N_10994,N_10568);
xnor U11279 (N_11279,N_10884,N_10866);
xor U11280 (N_11280,N_10742,N_10921);
nand U11281 (N_11281,N_10642,N_10877);
and U11282 (N_11282,N_10983,N_10699);
xor U11283 (N_11283,N_10723,N_10958);
nand U11284 (N_11284,N_10639,N_10604);
nand U11285 (N_11285,N_10502,N_10970);
nor U11286 (N_11286,N_10591,N_10824);
or U11287 (N_11287,N_10802,N_10519);
xnor U11288 (N_11288,N_10805,N_10997);
nand U11289 (N_11289,N_10682,N_10848);
nand U11290 (N_11290,N_10717,N_10762);
nand U11291 (N_11291,N_10850,N_10658);
and U11292 (N_11292,N_10848,N_10567);
xor U11293 (N_11293,N_10837,N_10678);
and U11294 (N_11294,N_10555,N_10557);
or U11295 (N_11295,N_10551,N_10898);
xor U11296 (N_11296,N_10927,N_10501);
and U11297 (N_11297,N_10860,N_10844);
nor U11298 (N_11298,N_10530,N_10787);
or U11299 (N_11299,N_10694,N_10510);
nor U11300 (N_11300,N_10525,N_10900);
xor U11301 (N_11301,N_10723,N_10818);
xnor U11302 (N_11302,N_10904,N_10579);
xnor U11303 (N_11303,N_10693,N_10636);
xnor U11304 (N_11304,N_10710,N_10959);
and U11305 (N_11305,N_10822,N_10903);
or U11306 (N_11306,N_10734,N_10982);
nand U11307 (N_11307,N_10908,N_10827);
nand U11308 (N_11308,N_10862,N_10739);
and U11309 (N_11309,N_10981,N_10510);
nor U11310 (N_11310,N_10798,N_10616);
xor U11311 (N_11311,N_10927,N_10662);
nand U11312 (N_11312,N_10994,N_10876);
nand U11313 (N_11313,N_10552,N_10538);
or U11314 (N_11314,N_10910,N_10651);
nor U11315 (N_11315,N_10814,N_10710);
or U11316 (N_11316,N_10997,N_10692);
nor U11317 (N_11317,N_10991,N_10680);
nand U11318 (N_11318,N_10591,N_10792);
or U11319 (N_11319,N_10664,N_10603);
nand U11320 (N_11320,N_10576,N_10628);
nor U11321 (N_11321,N_10728,N_10645);
xor U11322 (N_11322,N_10534,N_10986);
or U11323 (N_11323,N_10926,N_10858);
or U11324 (N_11324,N_10688,N_10794);
or U11325 (N_11325,N_10980,N_10824);
nand U11326 (N_11326,N_10792,N_10936);
nor U11327 (N_11327,N_10734,N_10777);
and U11328 (N_11328,N_10601,N_10837);
and U11329 (N_11329,N_10847,N_10977);
nor U11330 (N_11330,N_10747,N_10770);
nand U11331 (N_11331,N_10591,N_10680);
nand U11332 (N_11332,N_10973,N_10801);
and U11333 (N_11333,N_10795,N_10522);
xor U11334 (N_11334,N_10762,N_10617);
xnor U11335 (N_11335,N_10574,N_10650);
nand U11336 (N_11336,N_10653,N_10830);
and U11337 (N_11337,N_10976,N_10915);
and U11338 (N_11338,N_10997,N_10808);
nor U11339 (N_11339,N_10883,N_10524);
or U11340 (N_11340,N_10574,N_10578);
nor U11341 (N_11341,N_10704,N_10695);
nor U11342 (N_11342,N_10557,N_10672);
nor U11343 (N_11343,N_10551,N_10659);
nand U11344 (N_11344,N_10768,N_10577);
or U11345 (N_11345,N_10832,N_10768);
nor U11346 (N_11346,N_10631,N_10889);
xor U11347 (N_11347,N_10703,N_10827);
xnor U11348 (N_11348,N_10981,N_10566);
nand U11349 (N_11349,N_10962,N_10859);
nor U11350 (N_11350,N_10693,N_10755);
and U11351 (N_11351,N_10725,N_10575);
and U11352 (N_11352,N_10562,N_10783);
and U11353 (N_11353,N_10837,N_10878);
and U11354 (N_11354,N_10653,N_10769);
xnor U11355 (N_11355,N_10989,N_10783);
nand U11356 (N_11356,N_10520,N_10500);
or U11357 (N_11357,N_10951,N_10733);
xnor U11358 (N_11358,N_10804,N_10641);
and U11359 (N_11359,N_10621,N_10976);
xor U11360 (N_11360,N_10760,N_10563);
or U11361 (N_11361,N_10575,N_10603);
and U11362 (N_11362,N_10597,N_10686);
nor U11363 (N_11363,N_10852,N_10679);
and U11364 (N_11364,N_10886,N_10921);
xnor U11365 (N_11365,N_10662,N_10645);
nand U11366 (N_11366,N_10626,N_10556);
or U11367 (N_11367,N_10991,N_10546);
or U11368 (N_11368,N_10772,N_10955);
nand U11369 (N_11369,N_10723,N_10815);
xnor U11370 (N_11370,N_10867,N_10638);
and U11371 (N_11371,N_10964,N_10614);
nor U11372 (N_11372,N_10950,N_10815);
nand U11373 (N_11373,N_10792,N_10788);
and U11374 (N_11374,N_10735,N_10580);
xnor U11375 (N_11375,N_10854,N_10682);
xor U11376 (N_11376,N_10615,N_10881);
xor U11377 (N_11377,N_10716,N_10547);
nand U11378 (N_11378,N_10860,N_10936);
nor U11379 (N_11379,N_10930,N_10992);
or U11380 (N_11380,N_10889,N_10594);
xnor U11381 (N_11381,N_10676,N_10605);
xor U11382 (N_11382,N_10623,N_10749);
or U11383 (N_11383,N_10982,N_10903);
or U11384 (N_11384,N_10676,N_10538);
nand U11385 (N_11385,N_10928,N_10911);
xnor U11386 (N_11386,N_10754,N_10569);
and U11387 (N_11387,N_10872,N_10621);
and U11388 (N_11388,N_10732,N_10841);
or U11389 (N_11389,N_10993,N_10927);
or U11390 (N_11390,N_10602,N_10615);
nand U11391 (N_11391,N_10652,N_10821);
nor U11392 (N_11392,N_10647,N_10650);
and U11393 (N_11393,N_10694,N_10655);
nor U11394 (N_11394,N_10646,N_10787);
or U11395 (N_11395,N_10561,N_10932);
or U11396 (N_11396,N_10702,N_10711);
nand U11397 (N_11397,N_10823,N_10800);
nand U11398 (N_11398,N_10787,N_10920);
and U11399 (N_11399,N_10780,N_10529);
xnor U11400 (N_11400,N_10846,N_10749);
nand U11401 (N_11401,N_10998,N_10783);
xor U11402 (N_11402,N_10940,N_10744);
and U11403 (N_11403,N_10764,N_10608);
or U11404 (N_11404,N_10703,N_10745);
and U11405 (N_11405,N_10615,N_10807);
or U11406 (N_11406,N_10543,N_10601);
or U11407 (N_11407,N_10897,N_10847);
nor U11408 (N_11408,N_10547,N_10734);
or U11409 (N_11409,N_10560,N_10589);
nand U11410 (N_11410,N_10509,N_10859);
nor U11411 (N_11411,N_10565,N_10513);
and U11412 (N_11412,N_10628,N_10508);
nand U11413 (N_11413,N_10542,N_10748);
nor U11414 (N_11414,N_10705,N_10866);
nand U11415 (N_11415,N_10940,N_10844);
and U11416 (N_11416,N_10660,N_10535);
nand U11417 (N_11417,N_10825,N_10991);
xor U11418 (N_11418,N_10826,N_10603);
or U11419 (N_11419,N_10804,N_10780);
nand U11420 (N_11420,N_10715,N_10969);
xor U11421 (N_11421,N_10663,N_10812);
and U11422 (N_11422,N_10913,N_10655);
nand U11423 (N_11423,N_10671,N_10904);
nand U11424 (N_11424,N_10997,N_10856);
xnor U11425 (N_11425,N_10622,N_10903);
nand U11426 (N_11426,N_10577,N_10687);
or U11427 (N_11427,N_10925,N_10663);
nor U11428 (N_11428,N_10505,N_10515);
or U11429 (N_11429,N_10570,N_10868);
xnor U11430 (N_11430,N_10915,N_10912);
nor U11431 (N_11431,N_10666,N_10585);
nor U11432 (N_11432,N_10555,N_10621);
or U11433 (N_11433,N_10529,N_10695);
xor U11434 (N_11434,N_10871,N_10926);
and U11435 (N_11435,N_10519,N_10940);
and U11436 (N_11436,N_10909,N_10707);
and U11437 (N_11437,N_10743,N_10916);
and U11438 (N_11438,N_10977,N_10938);
xnor U11439 (N_11439,N_10788,N_10646);
nand U11440 (N_11440,N_10872,N_10572);
or U11441 (N_11441,N_10732,N_10541);
nand U11442 (N_11442,N_10827,N_10984);
xnor U11443 (N_11443,N_10758,N_10951);
xnor U11444 (N_11444,N_10865,N_10873);
nor U11445 (N_11445,N_10882,N_10910);
xnor U11446 (N_11446,N_10513,N_10651);
and U11447 (N_11447,N_10967,N_10959);
and U11448 (N_11448,N_10756,N_10543);
xor U11449 (N_11449,N_10952,N_10722);
xor U11450 (N_11450,N_10868,N_10791);
nor U11451 (N_11451,N_10871,N_10822);
or U11452 (N_11452,N_10656,N_10796);
or U11453 (N_11453,N_10541,N_10879);
nand U11454 (N_11454,N_10944,N_10551);
or U11455 (N_11455,N_10942,N_10640);
and U11456 (N_11456,N_10960,N_10915);
or U11457 (N_11457,N_10526,N_10967);
xnor U11458 (N_11458,N_10863,N_10944);
xnor U11459 (N_11459,N_10987,N_10960);
nor U11460 (N_11460,N_10991,N_10671);
and U11461 (N_11461,N_10787,N_10714);
nor U11462 (N_11462,N_10692,N_10585);
xor U11463 (N_11463,N_10938,N_10888);
xnor U11464 (N_11464,N_10582,N_10507);
nand U11465 (N_11465,N_10668,N_10986);
xor U11466 (N_11466,N_10795,N_10603);
and U11467 (N_11467,N_10673,N_10628);
and U11468 (N_11468,N_10557,N_10751);
and U11469 (N_11469,N_10934,N_10521);
nor U11470 (N_11470,N_10984,N_10893);
or U11471 (N_11471,N_10984,N_10675);
nand U11472 (N_11472,N_10683,N_10656);
nand U11473 (N_11473,N_10543,N_10915);
xnor U11474 (N_11474,N_10662,N_10667);
xor U11475 (N_11475,N_10939,N_10600);
xnor U11476 (N_11476,N_10884,N_10928);
nand U11477 (N_11477,N_10589,N_10568);
xor U11478 (N_11478,N_10904,N_10701);
or U11479 (N_11479,N_10995,N_10549);
and U11480 (N_11480,N_10904,N_10979);
nand U11481 (N_11481,N_10922,N_10952);
xor U11482 (N_11482,N_10774,N_10526);
nand U11483 (N_11483,N_10950,N_10504);
xnor U11484 (N_11484,N_10773,N_10688);
and U11485 (N_11485,N_10930,N_10935);
and U11486 (N_11486,N_10964,N_10590);
nor U11487 (N_11487,N_10697,N_10661);
or U11488 (N_11488,N_10550,N_10592);
or U11489 (N_11489,N_10546,N_10872);
and U11490 (N_11490,N_10836,N_10600);
and U11491 (N_11491,N_10623,N_10937);
or U11492 (N_11492,N_10592,N_10647);
xnor U11493 (N_11493,N_10967,N_10924);
xor U11494 (N_11494,N_10748,N_10924);
nor U11495 (N_11495,N_10548,N_10948);
nor U11496 (N_11496,N_10992,N_10923);
nor U11497 (N_11497,N_10586,N_10789);
xnor U11498 (N_11498,N_10949,N_10711);
nand U11499 (N_11499,N_10859,N_10784);
xnor U11500 (N_11500,N_11342,N_11238);
nand U11501 (N_11501,N_11141,N_11318);
or U11502 (N_11502,N_11057,N_11220);
nand U11503 (N_11503,N_11052,N_11275);
or U11504 (N_11504,N_11295,N_11451);
nand U11505 (N_11505,N_11330,N_11251);
or U11506 (N_11506,N_11065,N_11440);
or U11507 (N_11507,N_11142,N_11150);
or U11508 (N_11508,N_11023,N_11077);
nand U11509 (N_11509,N_11037,N_11305);
nand U11510 (N_11510,N_11045,N_11331);
nor U11511 (N_11511,N_11063,N_11343);
nor U11512 (N_11512,N_11496,N_11125);
xor U11513 (N_11513,N_11061,N_11226);
nor U11514 (N_11514,N_11394,N_11247);
and U11515 (N_11515,N_11152,N_11472);
or U11516 (N_11516,N_11400,N_11326);
or U11517 (N_11517,N_11283,N_11172);
xor U11518 (N_11518,N_11461,N_11200);
xor U11519 (N_11519,N_11216,N_11107);
or U11520 (N_11520,N_11431,N_11372);
and U11521 (N_11521,N_11104,N_11294);
or U11522 (N_11522,N_11351,N_11462);
xor U11523 (N_11523,N_11457,N_11064);
nor U11524 (N_11524,N_11194,N_11098);
nor U11525 (N_11525,N_11156,N_11430);
xnor U11526 (N_11526,N_11232,N_11270);
or U11527 (N_11527,N_11006,N_11427);
xor U11528 (N_11528,N_11178,N_11022);
or U11529 (N_11529,N_11079,N_11284);
or U11530 (N_11530,N_11231,N_11035);
nand U11531 (N_11531,N_11480,N_11073);
and U11532 (N_11532,N_11004,N_11467);
and U11533 (N_11533,N_11367,N_11137);
xnor U11534 (N_11534,N_11187,N_11448);
or U11535 (N_11535,N_11222,N_11008);
or U11536 (N_11536,N_11016,N_11429);
and U11537 (N_11537,N_11191,N_11197);
nand U11538 (N_11538,N_11375,N_11076);
or U11539 (N_11539,N_11258,N_11227);
nand U11540 (N_11540,N_11031,N_11425);
nor U11541 (N_11541,N_11285,N_11129);
nor U11542 (N_11542,N_11420,N_11252);
nor U11543 (N_11543,N_11248,N_11074);
or U11544 (N_11544,N_11368,N_11167);
and U11545 (N_11545,N_11289,N_11051);
and U11546 (N_11546,N_11335,N_11328);
xor U11547 (N_11547,N_11358,N_11366);
nand U11548 (N_11548,N_11382,N_11039);
and U11549 (N_11549,N_11403,N_11376);
nor U11550 (N_11550,N_11101,N_11445);
and U11551 (N_11551,N_11314,N_11133);
nor U11552 (N_11552,N_11166,N_11319);
or U11553 (N_11553,N_11207,N_11396);
or U11554 (N_11554,N_11334,N_11301);
xnor U11555 (N_11555,N_11032,N_11347);
or U11556 (N_11556,N_11114,N_11482);
xnor U11557 (N_11557,N_11264,N_11340);
or U11558 (N_11558,N_11219,N_11488);
nand U11559 (N_11559,N_11249,N_11266);
nor U11560 (N_11560,N_11139,N_11424);
xor U11561 (N_11561,N_11091,N_11069);
xnor U11562 (N_11562,N_11337,N_11447);
or U11563 (N_11563,N_11071,N_11164);
and U11564 (N_11564,N_11109,N_11265);
xnor U11565 (N_11565,N_11182,N_11174);
nand U11566 (N_11566,N_11170,N_11214);
or U11567 (N_11567,N_11315,N_11393);
nand U11568 (N_11568,N_11213,N_11279);
nor U11569 (N_11569,N_11009,N_11134);
or U11570 (N_11570,N_11345,N_11409);
nand U11571 (N_11571,N_11365,N_11381);
nor U11572 (N_11572,N_11446,N_11012);
xor U11573 (N_11573,N_11014,N_11128);
nor U11574 (N_11574,N_11397,N_11422);
or U11575 (N_11575,N_11269,N_11388);
nand U11576 (N_11576,N_11370,N_11309);
and U11577 (N_11577,N_11276,N_11286);
xnor U11578 (N_11578,N_11384,N_11307);
nand U11579 (N_11579,N_11383,N_11498);
or U11580 (N_11580,N_11288,N_11239);
nand U11581 (N_11581,N_11161,N_11005);
xnor U11582 (N_11582,N_11413,N_11070);
and U11583 (N_11583,N_11020,N_11291);
nand U11584 (N_11584,N_11481,N_11210);
or U11585 (N_11585,N_11120,N_11089);
nand U11586 (N_11586,N_11123,N_11416);
xor U11587 (N_11587,N_11303,N_11323);
and U11588 (N_11588,N_11463,N_11362);
or U11589 (N_11589,N_11281,N_11024);
nor U11590 (N_11590,N_11329,N_11453);
nor U11591 (N_11591,N_11296,N_11179);
or U11592 (N_11592,N_11349,N_11059);
nand U11593 (N_11593,N_11243,N_11072);
or U11594 (N_11594,N_11293,N_11302);
or U11595 (N_11595,N_11456,N_11162);
nor U11596 (N_11596,N_11483,N_11352);
nor U11597 (N_11597,N_11298,N_11404);
nor U11598 (N_11598,N_11183,N_11184);
nand U11599 (N_11599,N_11452,N_11121);
xnor U11600 (N_11600,N_11157,N_11459);
and U11601 (N_11601,N_11475,N_11245);
or U11602 (N_11602,N_11021,N_11414);
xnor U11603 (N_11603,N_11113,N_11019);
nand U11604 (N_11604,N_11111,N_11398);
nor U11605 (N_11605,N_11437,N_11188);
and U11606 (N_11606,N_11173,N_11148);
or U11607 (N_11607,N_11122,N_11435);
or U11608 (N_11608,N_11218,N_11344);
and U11609 (N_11609,N_11190,N_11259);
nor U11610 (N_11610,N_11067,N_11225);
xor U11611 (N_11611,N_11242,N_11158);
nand U11612 (N_11612,N_11084,N_11105);
or U11613 (N_11613,N_11208,N_11441);
or U11614 (N_11614,N_11412,N_11272);
nand U11615 (N_11615,N_11085,N_11401);
xor U11616 (N_11616,N_11353,N_11055);
and U11617 (N_11617,N_11075,N_11405);
and U11618 (N_11618,N_11479,N_11257);
and U11619 (N_11619,N_11277,N_11086);
xnor U11620 (N_11620,N_11081,N_11465);
nand U11621 (N_11621,N_11038,N_11095);
nor U11622 (N_11622,N_11028,N_11237);
nand U11623 (N_11623,N_11324,N_11262);
xnor U11624 (N_11624,N_11357,N_11003);
and U11625 (N_11625,N_11325,N_11018);
nor U11626 (N_11626,N_11127,N_11499);
or U11627 (N_11627,N_11118,N_11491);
xor U11628 (N_11628,N_11332,N_11348);
nand U11629 (N_11629,N_11449,N_11477);
xnor U11630 (N_11630,N_11374,N_11322);
nor U11631 (N_11631,N_11092,N_11093);
xnor U11632 (N_11632,N_11115,N_11406);
and U11633 (N_11633,N_11470,N_11147);
nor U11634 (N_11634,N_11389,N_11175);
xor U11635 (N_11635,N_11390,N_11436);
xnor U11636 (N_11636,N_11155,N_11246);
xnor U11637 (N_11637,N_11131,N_11198);
nand U11638 (N_11638,N_11407,N_11354);
or U11639 (N_11639,N_11025,N_11181);
xor U11640 (N_11640,N_11117,N_11078);
nor U11641 (N_11641,N_11240,N_11203);
nor U11642 (N_11642,N_11364,N_11485);
nor U11643 (N_11643,N_11042,N_11165);
nand U11644 (N_11644,N_11391,N_11495);
nand U11645 (N_11645,N_11377,N_11244);
nand U11646 (N_11646,N_11316,N_11317);
nand U11647 (N_11647,N_11228,N_11419);
nand U11648 (N_11648,N_11177,N_11168);
nand U11649 (N_11649,N_11490,N_11468);
nor U11650 (N_11650,N_11224,N_11153);
nor U11651 (N_11651,N_11029,N_11356);
nor U11652 (N_11652,N_11080,N_11094);
nand U11653 (N_11653,N_11410,N_11255);
xor U11654 (N_11654,N_11209,N_11484);
nor U11655 (N_11655,N_11333,N_11434);
xnor U11656 (N_11656,N_11492,N_11408);
xor U11657 (N_11657,N_11169,N_11135);
or U11658 (N_11658,N_11221,N_11215);
nand U11659 (N_11659,N_11015,N_11359);
xor U11660 (N_11660,N_11493,N_11017);
and U11661 (N_11661,N_11455,N_11106);
xor U11662 (N_11662,N_11320,N_11268);
and U11663 (N_11663,N_11146,N_11471);
nor U11664 (N_11664,N_11185,N_11066);
xor U11665 (N_11665,N_11379,N_11083);
nor U11666 (N_11666,N_11151,N_11474);
or U11667 (N_11667,N_11062,N_11116);
nor U11668 (N_11668,N_11274,N_11000);
nand U11669 (N_11669,N_11371,N_11196);
and U11670 (N_11670,N_11442,N_11068);
nor U11671 (N_11671,N_11217,N_11176);
and U11672 (N_11672,N_11261,N_11439);
nor U11673 (N_11673,N_11464,N_11205);
or U11674 (N_11674,N_11103,N_11466);
xnor U11675 (N_11675,N_11204,N_11234);
nand U11676 (N_11676,N_11049,N_11233);
or U11677 (N_11677,N_11201,N_11088);
or U11678 (N_11678,N_11102,N_11327);
or U11679 (N_11679,N_11361,N_11050);
nor U11680 (N_11680,N_11056,N_11013);
or U11681 (N_11681,N_11282,N_11236);
nand U11682 (N_11682,N_11206,N_11159);
and U11683 (N_11683,N_11273,N_11469);
or U11684 (N_11684,N_11360,N_11443);
xor U11685 (N_11685,N_11087,N_11421);
xnor U11686 (N_11686,N_11260,N_11423);
or U11687 (N_11687,N_11369,N_11189);
nand U11688 (N_11688,N_11418,N_11223);
nor U11689 (N_11689,N_11486,N_11041);
and U11690 (N_11690,N_11180,N_11034);
nor U11691 (N_11691,N_11411,N_11494);
and U11692 (N_11692,N_11138,N_11432);
and U11693 (N_11693,N_11202,N_11476);
or U11694 (N_11694,N_11163,N_11195);
xnor U11695 (N_11695,N_11011,N_11054);
and U11696 (N_11696,N_11082,N_11438);
nand U11697 (N_11697,N_11036,N_11254);
nor U11698 (N_11698,N_11132,N_11280);
xnor U11699 (N_11699,N_11338,N_11256);
and U11700 (N_11700,N_11110,N_11497);
or U11701 (N_11701,N_11350,N_11415);
xor U11702 (N_11702,N_11136,N_11212);
xor U11703 (N_11703,N_11140,N_11230);
and U11704 (N_11704,N_11100,N_11058);
nor U11705 (N_11705,N_11399,N_11473);
nand U11706 (N_11706,N_11363,N_11428);
nand U11707 (N_11707,N_11312,N_11160);
nand U11708 (N_11708,N_11060,N_11460);
and U11709 (N_11709,N_11043,N_11311);
nand U11710 (N_11710,N_11308,N_11186);
nand U11711 (N_11711,N_11002,N_11253);
or U11712 (N_11712,N_11395,N_11297);
and U11713 (N_11713,N_11053,N_11454);
nor U11714 (N_11714,N_11292,N_11355);
xor U11715 (N_11715,N_11033,N_11433);
nor U11716 (N_11716,N_11001,N_11306);
and U11717 (N_11717,N_11386,N_11199);
xnor U11718 (N_11718,N_11030,N_11380);
xnor U11719 (N_11719,N_11321,N_11241);
or U11720 (N_11720,N_11192,N_11046);
or U11721 (N_11721,N_11007,N_11097);
nand U11722 (N_11722,N_11047,N_11385);
nor U11723 (N_11723,N_11278,N_11149);
xor U11724 (N_11724,N_11341,N_11267);
nand U11725 (N_11725,N_11271,N_11108);
or U11726 (N_11726,N_11339,N_11044);
xnor U11727 (N_11727,N_11229,N_11171);
or U11728 (N_11728,N_11426,N_11145);
nor U11729 (N_11729,N_11250,N_11450);
xor U11730 (N_11730,N_11387,N_11124);
nand U11731 (N_11731,N_11287,N_11126);
or U11732 (N_11732,N_11112,N_11026);
nand U11733 (N_11733,N_11402,N_11300);
or U11734 (N_11734,N_11304,N_11487);
xor U11735 (N_11735,N_11027,N_11010);
and U11736 (N_11736,N_11290,N_11099);
and U11737 (N_11737,N_11313,N_11048);
nor U11738 (N_11738,N_11392,N_11478);
nor U11739 (N_11739,N_11489,N_11336);
nor U11740 (N_11740,N_11040,N_11154);
nor U11741 (N_11741,N_11444,N_11144);
nand U11742 (N_11742,N_11090,N_11458);
xor U11743 (N_11743,N_11373,N_11130);
and U11744 (N_11744,N_11310,N_11193);
and U11745 (N_11745,N_11096,N_11235);
nand U11746 (N_11746,N_11346,N_11143);
or U11747 (N_11747,N_11211,N_11299);
xnor U11748 (N_11748,N_11119,N_11378);
and U11749 (N_11749,N_11417,N_11263);
nor U11750 (N_11750,N_11000,N_11224);
or U11751 (N_11751,N_11281,N_11258);
or U11752 (N_11752,N_11452,N_11435);
nor U11753 (N_11753,N_11399,N_11283);
nand U11754 (N_11754,N_11072,N_11347);
nand U11755 (N_11755,N_11469,N_11373);
xor U11756 (N_11756,N_11386,N_11169);
nand U11757 (N_11757,N_11407,N_11194);
or U11758 (N_11758,N_11320,N_11319);
xor U11759 (N_11759,N_11414,N_11137);
nand U11760 (N_11760,N_11177,N_11378);
or U11761 (N_11761,N_11216,N_11003);
nor U11762 (N_11762,N_11304,N_11139);
and U11763 (N_11763,N_11365,N_11147);
nor U11764 (N_11764,N_11324,N_11396);
nor U11765 (N_11765,N_11089,N_11344);
and U11766 (N_11766,N_11358,N_11064);
xor U11767 (N_11767,N_11489,N_11421);
and U11768 (N_11768,N_11282,N_11407);
nor U11769 (N_11769,N_11101,N_11035);
and U11770 (N_11770,N_11122,N_11320);
or U11771 (N_11771,N_11293,N_11307);
nor U11772 (N_11772,N_11061,N_11281);
and U11773 (N_11773,N_11149,N_11425);
nand U11774 (N_11774,N_11148,N_11454);
xnor U11775 (N_11775,N_11337,N_11378);
nor U11776 (N_11776,N_11205,N_11414);
nor U11777 (N_11777,N_11447,N_11437);
and U11778 (N_11778,N_11149,N_11460);
and U11779 (N_11779,N_11197,N_11176);
and U11780 (N_11780,N_11114,N_11059);
xnor U11781 (N_11781,N_11056,N_11330);
nor U11782 (N_11782,N_11147,N_11091);
or U11783 (N_11783,N_11484,N_11433);
xor U11784 (N_11784,N_11490,N_11013);
nor U11785 (N_11785,N_11377,N_11167);
or U11786 (N_11786,N_11274,N_11040);
xor U11787 (N_11787,N_11312,N_11290);
and U11788 (N_11788,N_11063,N_11053);
or U11789 (N_11789,N_11247,N_11401);
and U11790 (N_11790,N_11252,N_11363);
nor U11791 (N_11791,N_11077,N_11394);
or U11792 (N_11792,N_11246,N_11054);
and U11793 (N_11793,N_11215,N_11328);
or U11794 (N_11794,N_11030,N_11196);
nand U11795 (N_11795,N_11437,N_11302);
xor U11796 (N_11796,N_11472,N_11104);
and U11797 (N_11797,N_11289,N_11424);
or U11798 (N_11798,N_11483,N_11190);
xor U11799 (N_11799,N_11227,N_11368);
or U11800 (N_11800,N_11006,N_11123);
nand U11801 (N_11801,N_11437,N_11309);
xor U11802 (N_11802,N_11443,N_11135);
nor U11803 (N_11803,N_11039,N_11084);
nor U11804 (N_11804,N_11281,N_11304);
nor U11805 (N_11805,N_11265,N_11239);
xnor U11806 (N_11806,N_11236,N_11013);
xor U11807 (N_11807,N_11324,N_11491);
and U11808 (N_11808,N_11347,N_11069);
nand U11809 (N_11809,N_11199,N_11205);
or U11810 (N_11810,N_11383,N_11016);
and U11811 (N_11811,N_11302,N_11016);
nor U11812 (N_11812,N_11004,N_11486);
nor U11813 (N_11813,N_11247,N_11495);
and U11814 (N_11814,N_11151,N_11032);
nand U11815 (N_11815,N_11110,N_11429);
nand U11816 (N_11816,N_11466,N_11008);
nand U11817 (N_11817,N_11342,N_11471);
nor U11818 (N_11818,N_11484,N_11321);
nor U11819 (N_11819,N_11018,N_11394);
and U11820 (N_11820,N_11495,N_11286);
xnor U11821 (N_11821,N_11164,N_11338);
nand U11822 (N_11822,N_11072,N_11138);
and U11823 (N_11823,N_11043,N_11188);
or U11824 (N_11824,N_11333,N_11423);
nand U11825 (N_11825,N_11317,N_11217);
nand U11826 (N_11826,N_11224,N_11333);
and U11827 (N_11827,N_11351,N_11159);
and U11828 (N_11828,N_11082,N_11129);
nor U11829 (N_11829,N_11308,N_11322);
and U11830 (N_11830,N_11334,N_11220);
or U11831 (N_11831,N_11036,N_11163);
or U11832 (N_11832,N_11354,N_11153);
or U11833 (N_11833,N_11049,N_11347);
or U11834 (N_11834,N_11035,N_11450);
nand U11835 (N_11835,N_11038,N_11140);
nand U11836 (N_11836,N_11449,N_11181);
nor U11837 (N_11837,N_11225,N_11291);
and U11838 (N_11838,N_11387,N_11251);
xor U11839 (N_11839,N_11373,N_11200);
nor U11840 (N_11840,N_11000,N_11346);
or U11841 (N_11841,N_11310,N_11062);
and U11842 (N_11842,N_11497,N_11289);
or U11843 (N_11843,N_11055,N_11490);
nor U11844 (N_11844,N_11253,N_11136);
nor U11845 (N_11845,N_11049,N_11044);
or U11846 (N_11846,N_11499,N_11075);
nand U11847 (N_11847,N_11030,N_11327);
or U11848 (N_11848,N_11200,N_11014);
xor U11849 (N_11849,N_11286,N_11378);
xor U11850 (N_11850,N_11000,N_11297);
and U11851 (N_11851,N_11416,N_11117);
xor U11852 (N_11852,N_11261,N_11289);
nand U11853 (N_11853,N_11321,N_11018);
nand U11854 (N_11854,N_11038,N_11428);
nor U11855 (N_11855,N_11220,N_11222);
and U11856 (N_11856,N_11207,N_11397);
nor U11857 (N_11857,N_11446,N_11300);
and U11858 (N_11858,N_11499,N_11198);
xor U11859 (N_11859,N_11094,N_11058);
or U11860 (N_11860,N_11078,N_11294);
xnor U11861 (N_11861,N_11105,N_11044);
or U11862 (N_11862,N_11306,N_11318);
nand U11863 (N_11863,N_11423,N_11495);
nor U11864 (N_11864,N_11354,N_11119);
nor U11865 (N_11865,N_11378,N_11406);
and U11866 (N_11866,N_11178,N_11450);
xor U11867 (N_11867,N_11205,N_11164);
or U11868 (N_11868,N_11254,N_11302);
or U11869 (N_11869,N_11290,N_11018);
nor U11870 (N_11870,N_11178,N_11090);
and U11871 (N_11871,N_11285,N_11263);
nor U11872 (N_11872,N_11488,N_11367);
or U11873 (N_11873,N_11450,N_11036);
nor U11874 (N_11874,N_11199,N_11051);
nor U11875 (N_11875,N_11195,N_11123);
nand U11876 (N_11876,N_11412,N_11241);
nor U11877 (N_11877,N_11243,N_11166);
nand U11878 (N_11878,N_11425,N_11115);
nand U11879 (N_11879,N_11009,N_11088);
nor U11880 (N_11880,N_11025,N_11048);
nand U11881 (N_11881,N_11042,N_11136);
and U11882 (N_11882,N_11009,N_11499);
xnor U11883 (N_11883,N_11019,N_11264);
or U11884 (N_11884,N_11132,N_11006);
and U11885 (N_11885,N_11017,N_11172);
and U11886 (N_11886,N_11247,N_11369);
xor U11887 (N_11887,N_11410,N_11236);
or U11888 (N_11888,N_11422,N_11368);
or U11889 (N_11889,N_11229,N_11041);
xor U11890 (N_11890,N_11071,N_11246);
and U11891 (N_11891,N_11284,N_11050);
nor U11892 (N_11892,N_11362,N_11457);
and U11893 (N_11893,N_11100,N_11384);
nor U11894 (N_11894,N_11493,N_11499);
nand U11895 (N_11895,N_11023,N_11301);
xor U11896 (N_11896,N_11292,N_11331);
or U11897 (N_11897,N_11373,N_11384);
xor U11898 (N_11898,N_11219,N_11458);
or U11899 (N_11899,N_11166,N_11007);
xnor U11900 (N_11900,N_11053,N_11433);
nor U11901 (N_11901,N_11149,N_11496);
nand U11902 (N_11902,N_11108,N_11467);
nor U11903 (N_11903,N_11222,N_11434);
nand U11904 (N_11904,N_11490,N_11036);
nand U11905 (N_11905,N_11054,N_11111);
nor U11906 (N_11906,N_11317,N_11332);
xnor U11907 (N_11907,N_11441,N_11265);
and U11908 (N_11908,N_11057,N_11162);
xnor U11909 (N_11909,N_11404,N_11449);
xnor U11910 (N_11910,N_11347,N_11352);
xnor U11911 (N_11911,N_11325,N_11141);
nand U11912 (N_11912,N_11186,N_11245);
xnor U11913 (N_11913,N_11080,N_11310);
nand U11914 (N_11914,N_11355,N_11377);
xnor U11915 (N_11915,N_11190,N_11045);
nand U11916 (N_11916,N_11059,N_11181);
xnor U11917 (N_11917,N_11433,N_11015);
xnor U11918 (N_11918,N_11431,N_11429);
xnor U11919 (N_11919,N_11357,N_11459);
nor U11920 (N_11920,N_11202,N_11017);
xor U11921 (N_11921,N_11313,N_11488);
and U11922 (N_11922,N_11129,N_11049);
and U11923 (N_11923,N_11086,N_11381);
nor U11924 (N_11924,N_11442,N_11327);
nand U11925 (N_11925,N_11295,N_11255);
or U11926 (N_11926,N_11400,N_11419);
and U11927 (N_11927,N_11302,N_11193);
nor U11928 (N_11928,N_11001,N_11092);
nand U11929 (N_11929,N_11244,N_11345);
xnor U11930 (N_11930,N_11031,N_11372);
xnor U11931 (N_11931,N_11275,N_11082);
or U11932 (N_11932,N_11168,N_11171);
nand U11933 (N_11933,N_11245,N_11131);
nand U11934 (N_11934,N_11121,N_11224);
nand U11935 (N_11935,N_11411,N_11470);
or U11936 (N_11936,N_11385,N_11068);
xor U11937 (N_11937,N_11369,N_11100);
xnor U11938 (N_11938,N_11452,N_11142);
or U11939 (N_11939,N_11409,N_11054);
nor U11940 (N_11940,N_11340,N_11285);
and U11941 (N_11941,N_11226,N_11234);
xnor U11942 (N_11942,N_11310,N_11318);
nor U11943 (N_11943,N_11118,N_11282);
xnor U11944 (N_11944,N_11068,N_11105);
nor U11945 (N_11945,N_11349,N_11019);
xor U11946 (N_11946,N_11245,N_11003);
nand U11947 (N_11947,N_11483,N_11453);
xor U11948 (N_11948,N_11345,N_11233);
nor U11949 (N_11949,N_11275,N_11319);
and U11950 (N_11950,N_11222,N_11440);
xnor U11951 (N_11951,N_11157,N_11036);
or U11952 (N_11952,N_11481,N_11224);
nand U11953 (N_11953,N_11056,N_11099);
and U11954 (N_11954,N_11030,N_11419);
xor U11955 (N_11955,N_11404,N_11492);
nand U11956 (N_11956,N_11464,N_11091);
nor U11957 (N_11957,N_11242,N_11169);
nand U11958 (N_11958,N_11343,N_11162);
or U11959 (N_11959,N_11350,N_11435);
and U11960 (N_11960,N_11087,N_11201);
nand U11961 (N_11961,N_11228,N_11352);
and U11962 (N_11962,N_11301,N_11046);
or U11963 (N_11963,N_11323,N_11204);
nand U11964 (N_11964,N_11265,N_11131);
nor U11965 (N_11965,N_11170,N_11139);
xnor U11966 (N_11966,N_11374,N_11093);
xnor U11967 (N_11967,N_11333,N_11022);
nand U11968 (N_11968,N_11224,N_11222);
nand U11969 (N_11969,N_11080,N_11478);
xnor U11970 (N_11970,N_11248,N_11336);
and U11971 (N_11971,N_11408,N_11451);
nor U11972 (N_11972,N_11231,N_11122);
and U11973 (N_11973,N_11390,N_11448);
nand U11974 (N_11974,N_11177,N_11364);
xor U11975 (N_11975,N_11099,N_11247);
and U11976 (N_11976,N_11405,N_11096);
nand U11977 (N_11977,N_11307,N_11417);
nand U11978 (N_11978,N_11462,N_11245);
and U11979 (N_11979,N_11368,N_11409);
xnor U11980 (N_11980,N_11257,N_11338);
and U11981 (N_11981,N_11023,N_11123);
nand U11982 (N_11982,N_11212,N_11461);
nand U11983 (N_11983,N_11436,N_11186);
xor U11984 (N_11984,N_11254,N_11199);
nor U11985 (N_11985,N_11009,N_11276);
or U11986 (N_11986,N_11004,N_11140);
nor U11987 (N_11987,N_11254,N_11401);
or U11988 (N_11988,N_11072,N_11338);
nor U11989 (N_11989,N_11368,N_11128);
or U11990 (N_11990,N_11017,N_11097);
nor U11991 (N_11991,N_11288,N_11245);
nand U11992 (N_11992,N_11390,N_11120);
nor U11993 (N_11993,N_11000,N_11318);
xnor U11994 (N_11994,N_11210,N_11106);
and U11995 (N_11995,N_11040,N_11360);
and U11996 (N_11996,N_11340,N_11470);
or U11997 (N_11997,N_11486,N_11472);
or U11998 (N_11998,N_11439,N_11122);
xnor U11999 (N_11999,N_11133,N_11303);
and U12000 (N_12000,N_11832,N_11805);
xnor U12001 (N_12001,N_11607,N_11559);
nand U12002 (N_12002,N_11591,N_11955);
xor U12003 (N_12003,N_11595,N_11814);
nand U12004 (N_12004,N_11572,N_11554);
xor U12005 (N_12005,N_11630,N_11867);
xor U12006 (N_12006,N_11958,N_11889);
or U12007 (N_12007,N_11503,N_11584);
xnor U12008 (N_12008,N_11544,N_11558);
xnor U12009 (N_12009,N_11516,N_11648);
nor U12010 (N_12010,N_11605,N_11632);
and U12011 (N_12011,N_11946,N_11986);
xnor U12012 (N_12012,N_11667,N_11862);
nor U12013 (N_12013,N_11570,N_11762);
and U12014 (N_12014,N_11902,N_11615);
and U12015 (N_12015,N_11880,N_11787);
and U12016 (N_12016,N_11643,N_11614);
nand U12017 (N_12017,N_11977,N_11852);
xor U12018 (N_12018,N_11789,N_11758);
nor U12019 (N_12019,N_11903,N_11702);
nor U12020 (N_12020,N_11690,N_11984);
or U12021 (N_12021,N_11836,N_11779);
nand U12022 (N_12022,N_11709,N_11991);
and U12023 (N_12023,N_11749,N_11565);
or U12024 (N_12024,N_11786,N_11775);
nor U12025 (N_12025,N_11788,N_11937);
nor U12026 (N_12026,N_11526,N_11750);
nand U12027 (N_12027,N_11560,N_11695);
or U12028 (N_12028,N_11699,N_11849);
and U12029 (N_12029,N_11881,N_11670);
nor U12030 (N_12030,N_11914,N_11548);
and U12031 (N_12031,N_11776,N_11864);
nand U12032 (N_12032,N_11590,N_11797);
or U12033 (N_12033,N_11523,N_11649);
xnor U12034 (N_12034,N_11997,N_11541);
nand U12035 (N_12035,N_11638,N_11803);
and U12036 (N_12036,N_11957,N_11688);
or U12037 (N_12037,N_11891,N_11571);
nand U12038 (N_12038,N_11680,N_11748);
nor U12039 (N_12039,N_11785,N_11936);
xor U12040 (N_12040,N_11794,N_11520);
nand U12041 (N_12041,N_11925,N_11932);
or U12042 (N_12042,N_11698,N_11765);
nand U12043 (N_12043,N_11641,N_11989);
or U12044 (N_12044,N_11979,N_11964);
nor U12045 (N_12045,N_11700,N_11943);
nand U12046 (N_12046,N_11692,N_11965);
nor U12047 (N_12047,N_11568,N_11747);
xnor U12048 (N_12048,N_11713,N_11701);
or U12049 (N_12049,N_11752,N_11655);
xnor U12050 (N_12050,N_11961,N_11743);
and U12051 (N_12051,N_11625,N_11509);
nand U12052 (N_12052,N_11987,N_11974);
nor U12053 (N_12053,N_11766,N_11998);
xnor U12054 (N_12054,N_11740,N_11642);
nor U12055 (N_12055,N_11848,N_11825);
or U12056 (N_12056,N_11622,N_11751);
or U12057 (N_12057,N_11816,N_11873);
nor U12058 (N_12058,N_11679,N_11736);
nand U12059 (N_12059,N_11725,N_11610);
xor U12060 (N_12060,N_11950,N_11659);
nor U12061 (N_12061,N_11988,N_11899);
nand U12062 (N_12062,N_11773,N_11598);
xnor U12063 (N_12063,N_11589,N_11744);
and U12064 (N_12064,N_11715,N_11636);
nand U12065 (N_12065,N_11954,N_11968);
and U12066 (N_12066,N_11710,N_11745);
nor U12067 (N_12067,N_11846,N_11871);
and U12068 (N_12068,N_11795,N_11578);
or U12069 (N_12069,N_11634,N_11663);
nand U12070 (N_12070,N_11983,N_11831);
xor U12071 (N_12071,N_11627,N_11637);
or U12072 (N_12072,N_11962,N_11582);
nand U12073 (N_12073,N_11791,N_11518);
or U12074 (N_12074,N_11819,N_11556);
nor U12075 (N_12075,N_11818,N_11777);
nor U12076 (N_12076,N_11539,N_11618);
xor U12077 (N_12077,N_11916,N_11729);
xor U12078 (N_12078,N_11919,N_11868);
and U12079 (N_12079,N_11508,N_11728);
nand U12080 (N_12080,N_11529,N_11697);
xnor U12081 (N_12081,N_11500,N_11804);
nor U12082 (N_12082,N_11938,N_11769);
nand U12083 (N_12083,N_11992,N_11647);
nor U12084 (N_12084,N_11908,N_11826);
nand U12085 (N_12085,N_11893,N_11858);
and U12086 (N_12086,N_11672,N_11857);
or U12087 (N_12087,N_11907,N_11808);
and U12088 (N_12088,N_11685,N_11521);
nor U12089 (N_12089,N_11756,N_11874);
nor U12090 (N_12090,N_11575,N_11809);
nand U12091 (N_12091,N_11802,N_11976);
xor U12092 (N_12092,N_11592,N_11682);
nor U12093 (N_12093,N_11928,N_11723);
nor U12094 (N_12094,N_11985,N_11612);
or U12095 (N_12095,N_11904,N_11927);
or U12096 (N_12096,N_11501,N_11734);
xor U12097 (N_12097,N_11597,N_11629);
nand U12098 (N_12098,N_11675,N_11882);
nor U12099 (N_12099,N_11604,N_11973);
or U12100 (N_12100,N_11945,N_11707);
xnor U12101 (N_12101,N_11566,N_11872);
nand U12102 (N_12102,N_11757,N_11549);
xnor U12103 (N_12103,N_11912,N_11942);
nor U12104 (N_12104,N_11854,N_11801);
or U12105 (N_12105,N_11845,N_11909);
xor U12106 (N_12106,N_11761,N_11822);
or U12107 (N_12107,N_11514,N_11877);
xnor U12108 (N_12108,N_11948,N_11719);
and U12109 (N_12109,N_11658,N_11533);
and U12110 (N_12110,N_11623,N_11724);
nor U12111 (N_12111,N_11673,N_11579);
nand U12112 (N_12112,N_11800,N_11553);
and U12113 (N_12113,N_11731,N_11755);
and U12114 (N_12114,N_11890,N_11653);
xnor U12115 (N_12115,N_11897,N_11654);
xor U12116 (N_12116,N_11617,N_11609);
and U12117 (N_12117,N_11567,N_11995);
nor U12118 (N_12118,N_11841,N_11537);
or U12119 (N_12119,N_11703,N_11650);
xnor U12120 (N_12120,N_11684,N_11967);
nor U12121 (N_12121,N_11810,N_11674);
or U12122 (N_12122,N_11771,N_11917);
or U12123 (N_12123,N_11662,N_11522);
and U12124 (N_12124,N_11531,N_11865);
xor U12125 (N_12125,N_11821,N_11830);
or U12126 (N_12126,N_11887,N_11746);
xnor U12127 (N_12127,N_11990,N_11913);
and U12128 (N_12128,N_11677,N_11633);
nor U12129 (N_12129,N_11660,N_11823);
nor U12130 (N_12130,N_11534,N_11820);
or U12131 (N_12131,N_11645,N_11827);
or U12132 (N_12132,N_11896,N_11982);
or U12133 (N_12133,N_11910,N_11861);
nor U12134 (N_12134,N_11644,N_11513);
nand U12135 (N_12135,N_11798,N_11770);
nor U12136 (N_12136,N_11711,N_11969);
xor U12137 (N_12137,N_11953,N_11866);
nand U12138 (N_12138,N_11878,N_11714);
xor U12139 (N_12139,N_11915,N_11599);
xnor U12140 (N_12140,N_11905,N_11602);
or U12141 (N_12141,N_11753,N_11506);
and U12142 (N_12142,N_11737,N_11894);
xnor U12143 (N_12143,N_11895,N_11828);
and U12144 (N_12144,N_11524,N_11975);
and U12145 (N_12145,N_11883,N_11726);
nor U12146 (N_12146,N_11721,N_11657);
xor U12147 (N_12147,N_11806,N_11519);
or U12148 (N_12148,N_11718,N_11666);
xor U12149 (N_12149,N_11603,N_11535);
nand U12150 (N_12150,N_11708,N_11628);
nor U12151 (N_12151,N_11515,N_11525);
and U12152 (N_12152,N_11594,N_11840);
xnor U12153 (N_12153,N_11952,N_11671);
nor U12154 (N_12154,N_11817,N_11920);
or U12155 (N_12155,N_11507,N_11542);
nand U12156 (N_12156,N_11853,N_11767);
xnor U12157 (N_12157,N_11783,N_11661);
nor U12158 (N_12158,N_11547,N_11716);
xnor U12159 (N_12159,N_11621,N_11624);
nand U12160 (N_12160,N_11935,N_11576);
nand U12161 (N_12161,N_11730,N_11669);
nor U12162 (N_12162,N_11530,N_11781);
xnor U12163 (N_12163,N_11586,N_11562);
nand U12164 (N_12164,N_11620,N_11839);
nor U12165 (N_12165,N_11900,N_11855);
nor U12166 (N_12166,N_11834,N_11956);
nor U12167 (N_12167,N_11687,N_11563);
nand U12168 (N_12168,N_11712,N_11838);
xor U12169 (N_12169,N_11664,N_11886);
and U12170 (N_12170,N_11504,N_11811);
and U12171 (N_12171,N_11600,N_11898);
or U12172 (N_12172,N_11583,N_11735);
and U12173 (N_12173,N_11933,N_11835);
or U12174 (N_12174,N_11668,N_11999);
xnor U12175 (N_12175,N_11588,N_11875);
and U12176 (N_12176,N_11739,N_11829);
or U12177 (N_12177,N_11843,N_11860);
nand U12178 (N_12178,N_11812,N_11683);
and U12179 (N_12179,N_11646,N_11678);
nand U12180 (N_12180,N_11601,N_11574);
nor U12181 (N_12181,N_11815,N_11686);
or U12182 (N_12182,N_11869,N_11764);
and U12183 (N_12183,N_11742,N_11759);
nor U12184 (N_12184,N_11930,N_11652);
xnor U12185 (N_12185,N_11512,N_11606);
xnor U12186 (N_12186,N_11774,N_11727);
or U12187 (N_12187,N_11705,N_11924);
and U12188 (N_12188,N_11611,N_11613);
or U12189 (N_12189,N_11884,N_11931);
or U12190 (N_12190,N_11545,N_11717);
xnor U12191 (N_12191,N_11778,N_11859);
or U12192 (N_12192,N_11694,N_11780);
or U12193 (N_12193,N_11921,N_11901);
nor U12194 (N_12194,N_11844,N_11966);
nor U12195 (N_12195,N_11577,N_11824);
nor U12196 (N_12196,N_11656,N_11741);
and U12197 (N_12197,N_11510,N_11635);
xnor U12198 (N_12198,N_11517,N_11947);
nor U12199 (N_12199,N_11546,N_11596);
nor U12200 (N_12200,N_11790,N_11842);
xnor U12201 (N_12201,N_11934,N_11555);
nand U12202 (N_12202,N_11782,N_11911);
nor U12203 (N_12203,N_11813,N_11906);
nand U12204 (N_12204,N_11505,N_11940);
and U12205 (N_12205,N_11949,N_11651);
xor U12206 (N_12206,N_11550,N_11768);
nor U12207 (N_12207,N_11996,N_11527);
xnor U12208 (N_12208,N_11951,N_11793);
and U12209 (N_12209,N_11754,N_11978);
or U12210 (N_12210,N_11941,N_11631);
nand U12211 (N_12211,N_11885,N_11959);
xnor U12212 (N_12212,N_11619,N_11561);
nand U12213 (N_12213,N_11792,N_11939);
nand U12214 (N_12214,N_11720,N_11640);
and U12215 (N_12215,N_11929,N_11693);
nand U12216 (N_12216,N_11837,N_11851);
xnor U12217 (N_12217,N_11502,N_11540);
nor U12218 (N_12218,N_11923,N_11552);
and U12219 (N_12219,N_11980,N_11944);
nor U12220 (N_12220,N_11888,N_11922);
nor U12221 (N_12221,N_11608,N_11532);
and U12222 (N_12222,N_11665,N_11689);
xnor U12223 (N_12223,N_11760,N_11963);
or U12224 (N_12224,N_11536,N_11993);
xnor U12225 (N_12225,N_11863,N_11681);
or U12226 (N_12226,N_11918,N_11580);
and U12227 (N_12227,N_11732,N_11528);
or U12228 (N_12228,N_11970,N_11799);
and U12229 (N_12229,N_11543,N_11994);
or U12230 (N_12230,N_11733,N_11639);
nand U12231 (N_12231,N_11972,N_11850);
nand U12232 (N_12232,N_11879,N_11870);
and U12233 (N_12233,N_11847,N_11772);
or U12234 (N_12234,N_11691,N_11971);
nand U12235 (N_12235,N_11511,N_11616);
or U12236 (N_12236,N_11981,N_11876);
nand U12237 (N_12237,N_11807,N_11704);
xor U12238 (N_12238,N_11581,N_11796);
and U12239 (N_12239,N_11593,N_11587);
and U12240 (N_12240,N_11676,N_11960);
or U12241 (N_12241,N_11706,N_11763);
nand U12242 (N_12242,N_11569,N_11557);
xor U12243 (N_12243,N_11585,N_11892);
and U12244 (N_12244,N_11626,N_11564);
and U12245 (N_12245,N_11738,N_11784);
or U12246 (N_12246,N_11926,N_11538);
xnor U12247 (N_12247,N_11833,N_11856);
xnor U12248 (N_12248,N_11696,N_11551);
nand U12249 (N_12249,N_11722,N_11573);
nor U12250 (N_12250,N_11753,N_11978);
and U12251 (N_12251,N_11993,N_11550);
nor U12252 (N_12252,N_11555,N_11945);
and U12253 (N_12253,N_11780,N_11639);
or U12254 (N_12254,N_11841,N_11741);
or U12255 (N_12255,N_11783,N_11713);
nand U12256 (N_12256,N_11635,N_11525);
and U12257 (N_12257,N_11640,N_11858);
nor U12258 (N_12258,N_11663,N_11896);
nand U12259 (N_12259,N_11645,N_11777);
xnor U12260 (N_12260,N_11799,N_11858);
or U12261 (N_12261,N_11534,N_11635);
nand U12262 (N_12262,N_11889,N_11699);
nand U12263 (N_12263,N_11889,N_11665);
and U12264 (N_12264,N_11652,N_11882);
or U12265 (N_12265,N_11505,N_11565);
nor U12266 (N_12266,N_11613,N_11824);
or U12267 (N_12267,N_11994,N_11584);
or U12268 (N_12268,N_11730,N_11658);
nor U12269 (N_12269,N_11821,N_11693);
nand U12270 (N_12270,N_11960,N_11952);
and U12271 (N_12271,N_11927,N_11530);
nand U12272 (N_12272,N_11847,N_11986);
xnor U12273 (N_12273,N_11852,N_11891);
nand U12274 (N_12274,N_11578,N_11930);
nand U12275 (N_12275,N_11749,N_11960);
xor U12276 (N_12276,N_11811,N_11747);
or U12277 (N_12277,N_11505,N_11719);
nand U12278 (N_12278,N_11652,N_11978);
nor U12279 (N_12279,N_11797,N_11618);
nor U12280 (N_12280,N_11536,N_11547);
xor U12281 (N_12281,N_11964,N_11764);
xnor U12282 (N_12282,N_11513,N_11637);
nand U12283 (N_12283,N_11845,N_11643);
nor U12284 (N_12284,N_11844,N_11750);
and U12285 (N_12285,N_11787,N_11799);
and U12286 (N_12286,N_11528,N_11814);
xnor U12287 (N_12287,N_11904,N_11905);
or U12288 (N_12288,N_11878,N_11511);
and U12289 (N_12289,N_11628,N_11786);
or U12290 (N_12290,N_11555,N_11900);
or U12291 (N_12291,N_11718,N_11536);
or U12292 (N_12292,N_11845,N_11816);
and U12293 (N_12293,N_11761,N_11811);
nor U12294 (N_12294,N_11854,N_11812);
nor U12295 (N_12295,N_11980,N_11733);
and U12296 (N_12296,N_11526,N_11800);
and U12297 (N_12297,N_11698,N_11838);
nand U12298 (N_12298,N_11764,N_11936);
xor U12299 (N_12299,N_11640,N_11738);
nand U12300 (N_12300,N_11692,N_11962);
or U12301 (N_12301,N_11623,N_11659);
nand U12302 (N_12302,N_11634,N_11869);
nand U12303 (N_12303,N_11903,N_11740);
and U12304 (N_12304,N_11985,N_11545);
xor U12305 (N_12305,N_11994,N_11761);
and U12306 (N_12306,N_11646,N_11633);
and U12307 (N_12307,N_11880,N_11543);
and U12308 (N_12308,N_11779,N_11596);
or U12309 (N_12309,N_11560,N_11898);
and U12310 (N_12310,N_11592,N_11796);
or U12311 (N_12311,N_11817,N_11925);
nor U12312 (N_12312,N_11934,N_11745);
nor U12313 (N_12313,N_11849,N_11562);
nand U12314 (N_12314,N_11924,N_11594);
xor U12315 (N_12315,N_11528,N_11839);
xnor U12316 (N_12316,N_11860,N_11633);
and U12317 (N_12317,N_11656,N_11611);
nand U12318 (N_12318,N_11721,N_11647);
nor U12319 (N_12319,N_11931,N_11999);
nand U12320 (N_12320,N_11526,N_11662);
nor U12321 (N_12321,N_11634,N_11803);
and U12322 (N_12322,N_11837,N_11769);
or U12323 (N_12323,N_11814,N_11997);
xnor U12324 (N_12324,N_11720,N_11737);
and U12325 (N_12325,N_11566,N_11555);
or U12326 (N_12326,N_11971,N_11582);
xnor U12327 (N_12327,N_11700,N_11900);
and U12328 (N_12328,N_11568,N_11848);
or U12329 (N_12329,N_11784,N_11987);
nand U12330 (N_12330,N_11656,N_11551);
nor U12331 (N_12331,N_11992,N_11558);
or U12332 (N_12332,N_11898,N_11977);
and U12333 (N_12333,N_11882,N_11991);
or U12334 (N_12334,N_11707,N_11782);
and U12335 (N_12335,N_11624,N_11797);
or U12336 (N_12336,N_11516,N_11745);
and U12337 (N_12337,N_11583,N_11882);
nand U12338 (N_12338,N_11545,N_11890);
nor U12339 (N_12339,N_11785,N_11592);
and U12340 (N_12340,N_11953,N_11629);
or U12341 (N_12341,N_11854,N_11667);
nand U12342 (N_12342,N_11767,N_11827);
or U12343 (N_12343,N_11561,N_11742);
or U12344 (N_12344,N_11881,N_11916);
nand U12345 (N_12345,N_11574,N_11845);
and U12346 (N_12346,N_11574,N_11752);
or U12347 (N_12347,N_11774,N_11710);
nor U12348 (N_12348,N_11541,N_11533);
or U12349 (N_12349,N_11709,N_11877);
nand U12350 (N_12350,N_11934,N_11847);
nor U12351 (N_12351,N_11648,N_11724);
xor U12352 (N_12352,N_11543,N_11785);
nand U12353 (N_12353,N_11545,N_11962);
and U12354 (N_12354,N_11799,N_11643);
or U12355 (N_12355,N_11686,N_11693);
xnor U12356 (N_12356,N_11898,N_11787);
nor U12357 (N_12357,N_11962,N_11677);
nand U12358 (N_12358,N_11816,N_11893);
or U12359 (N_12359,N_11961,N_11888);
nand U12360 (N_12360,N_11738,N_11654);
and U12361 (N_12361,N_11618,N_11736);
nand U12362 (N_12362,N_11557,N_11528);
and U12363 (N_12363,N_11817,N_11585);
xnor U12364 (N_12364,N_11567,N_11550);
xnor U12365 (N_12365,N_11970,N_11899);
nand U12366 (N_12366,N_11823,N_11657);
or U12367 (N_12367,N_11528,N_11565);
or U12368 (N_12368,N_11741,N_11529);
nand U12369 (N_12369,N_11700,N_11665);
nand U12370 (N_12370,N_11884,N_11715);
nand U12371 (N_12371,N_11830,N_11634);
and U12372 (N_12372,N_11780,N_11949);
nor U12373 (N_12373,N_11837,N_11790);
or U12374 (N_12374,N_11801,N_11905);
or U12375 (N_12375,N_11770,N_11577);
and U12376 (N_12376,N_11740,N_11896);
nor U12377 (N_12377,N_11733,N_11751);
or U12378 (N_12378,N_11810,N_11653);
and U12379 (N_12379,N_11651,N_11897);
nand U12380 (N_12380,N_11830,N_11683);
xnor U12381 (N_12381,N_11655,N_11836);
xnor U12382 (N_12382,N_11602,N_11700);
nor U12383 (N_12383,N_11728,N_11725);
nor U12384 (N_12384,N_11775,N_11544);
or U12385 (N_12385,N_11697,N_11970);
or U12386 (N_12386,N_11505,N_11957);
and U12387 (N_12387,N_11610,N_11790);
or U12388 (N_12388,N_11781,N_11830);
nand U12389 (N_12389,N_11709,N_11678);
or U12390 (N_12390,N_11655,N_11932);
and U12391 (N_12391,N_11547,N_11971);
or U12392 (N_12392,N_11866,N_11614);
nand U12393 (N_12393,N_11863,N_11689);
xor U12394 (N_12394,N_11823,N_11912);
nor U12395 (N_12395,N_11834,N_11917);
nor U12396 (N_12396,N_11966,N_11621);
and U12397 (N_12397,N_11677,N_11569);
and U12398 (N_12398,N_11752,N_11849);
nand U12399 (N_12399,N_11566,N_11543);
nor U12400 (N_12400,N_11653,N_11535);
or U12401 (N_12401,N_11684,N_11600);
or U12402 (N_12402,N_11536,N_11518);
or U12403 (N_12403,N_11905,N_11505);
nor U12404 (N_12404,N_11810,N_11713);
xor U12405 (N_12405,N_11924,N_11853);
or U12406 (N_12406,N_11967,N_11894);
or U12407 (N_12407,N_11804,N_11722);
nand U12408 (N_12408,N_11601,N_11951);
nor U12409 (N_12409,N_11912,N_11970);
or U12410 (N_12410,N_11557,N_11821);
nor U12411 (N_12411,N_11808,N_11931);
nor U12412 (N_12412,N_11842,N_11731);
nand U12413 (N_12413,N_11515,N_11718);
and U12414 (N_12414,N_11597,N_11772);
or U12415 (N_12415,N_11728,N_11775);
xnor U12416 (N_12416,N_11814,N_11850);
xnor U12417 (N_12417,N_11953,N_11942);
and U12418 (N_12418,N_11722,N_11539);
and U12419 (N_12419,N_11611,N_11727);
nand U12420 (N_12420,N_11882,N_11811);
xnor U12421 (N_12421,N_11865,N_11550);
xnor U12422 (N_12422,N_11905,N_11618);
nand U12423 (N_12423,N_11662,N_11915);
nor U12424 (N_12424,N_11624,N_11931);
nand U12425 (N_12425,N_11915,N_11513);
and U12426 (N_12426,N_11796,N_11621);
xnor U12427 (N_12427,N_11836,N_11964);
nand U12428 (N_12428,N_11733,N_11802);
nor U12429 (N_12429,N_11592,N_11750);
or U12430 (N_12430,N_11898,N_11973);
xnor U12431 (N_12431,N_11608,N_11653);
or U12432 (N_12432,N_11621,N_11817);
nor U12433 (N_12433,N_11881,N_11850);
and U12434 (N_12434,N_11798,N_11515);
nand U12435 (N_12435,N_11587,N_11601);
xnor U12436 (N_12436,N_11903,N_11514);
xor U12437 (N_12437,N_11531,N_11884);
and U12438 (N_12438,N_11660,N_11856);
xor U12439 (N_12439,N_11583,N_11963);
nand U12440 (N_12440,N_11968,N_11859);
nand U12441 (N_12441,N_11824,N_11562);
nand U12442 (N_12442,N_11898,N_11954);
xor U12443 (N_12443,N_11910,N_11836);
and U12444 (N_12444,N_11937,N_11838);
nand U12445 (N_12445,N_11880,N_11590);
nor U12446 (N_12446,N_11773,N_11767);
xnor U12447 (N_12447,N_11870,N_11669);
or U12448 (N_12448,N_11627,N_11884);
and U12449 (N_12449,N_11942,N_11908);
nor U12450 (N_12450,N_11619,N_11533);
xnor U12451 (N_12451,N_11635,N_11984);
nand U12452 (N_12452,N_11835,N_11849);
xnor U12453 (N_12453,N_11590,N_11935);
nor U12454 (N_12454,N_11738,N_11756);
nand U12455 (N_12455,N_11990,N_11904);
xor U12456 (N_12456,N_11529,N_11613);
and U12457 (N_12457,N_11759,N_11506);
xor U12458 (N_12458,N_11883,N_11711);
nand U12459 (N_12459,N_11500,N_11548);
or U12460 (N_12460,N_11954,N_11616);
nand U12461 (N_12461,N_11756,N_11821);
or U12462 (N_12462,N_11783,N_11503);
nor U12463 (N_12463,N_11860,N_11753);
nand U12464 (N_12464,N_11705,N_11935);
and U12465 (N_12465,N_11652,N_11953);
nand U12466 (N_12466,N_11539,N_11532);
or U12467 (N_12467,N_11896,N_11685);
xnor U12468 (N_12468,N_11568,N_11959);
nor U12469 (N_12469,N_11760,N_11730);
nor U12470 (N_12470,N_11878,N_11735);
and U12471 (N_12471,N_11759,N_11548);
and U12472 (N_12472,N_11604,N_11784);
xor U12473 (N_12473,N_11565,N_11964);
and U12474 (N_12474,N_11527,N_11702);
nand U12475 (N_12475,N_11936,N_11845);
or U12476 (N_12476,N_11906,N_11992);
xor U12477 (N_12477,N_11759,N_11724);
or U12478 (N_12478,N_11513,N_11615);
and U12479 (N_12479,N_11678,N_11799);
and U12480 (N_12480,N_11756,N_11808);
nand U12481 (N_12481,N_11869,N_11981);
xor U12482 (N_12482,N_11654,N_11512);
xor U12483 (N_12483,N_11993,N_11950);
or U12484 (N_12484,N_11688,N_11684);
nor U12485 (N_12485,N_11970,N_11991);
nand U12486 (N_12486,N_11923,N_11564);
xnor U12487 (N_12487,N_11659,N_11752);
or U12488 (N_12488,N_11782,N_11561);
or U12489 (N_12489,N_11538,N_11860);
and U12490 (N_12490,N_11838,N_11550);
nor U12491 (N_12491,N_11972,N_11812);
nor U12492 (N_12492,N_11754,N_11751);
nand U12493 (N_12493,N_11503,N_11524);
xor U12494 (N_12494,N_11745,N_11631);
nand U12495 (N_12495,N_11820,N_11961);
and U12496 (N_12496,N_11756,N_11982);
nand U12497 (N_12497,N_11983,N_11762);
and U12498 (N_12498,N_11664,N_11834);
nor U12499 (N_12499,N_11974,N_11678);
or U12500 (N_12500,N_12340,N_12427);
xnor U12501 (N_12501,N_12419,N_12399);
and U12502 (N_12502,N_12064,N_12172);
nor U12503 (N_12503,N_12263,N_12103);
or U12504 (N_12504,N_12290,N_12133);
or U12505 (N_12505,N_12489,N_12412);
and U12506 (N_12506,N_12137,N_12358);
nand U12507 (N_12507,N_12291,N_12052);
or U12508 (N_12508,N_12210,N_12081);
nor U12509 (N_12509,N_12475,N_12136);
nor U12510 (N_12510,N_12249,N_12048);
and U12511 (N_12511,N_12491,N_12192);
and U12512 (N_12512,N_12084,N_12104);
or U12513 (N_12513,N_12023,N_12378);
and U12514 (N_12514,N_12314,N_12303);
xor U12515 (N_12515,N_12339,N_12001);
nand U12516 (N_12516,N_12117,N_12486);
nor U12517 (N_12517,N_12197,N_12383);
and U12518 (N_12518,N_12119,N_12158);
xor U12519 (N_12519,N_12363,N_12444);
nor U12520 (N_12520,N_12224,N_12376);
or U12521 (N_12521,N_12413,N_12390);
xor U12522 (N_12522,N_12037,N_12415);
and U12523 (N_12523,N_12016,N_12080);
or U12524 (N_12524,N_12306,N_12464);
or U12525 (N_12525,N_12150,N_12068);
nand U12526 (N_12526,N_12253,N_12195);
nand U12527 (N_12527,N_12267,N_12047);
and U12528 (N_12528,N_12129,N_12442);
nand U12529 (N_12529,N_12176,N_12184);
or U12530 (N_12530,N_12327,N_12416);
or U12531 (N_12531,N_12452,N_12186);
nand U12532 (N_12532,N_12086,N_12035);
or U12533 (N_12533,N_12331,N_12190);
xor U12534 (N_12534,N_12252,N_12438);
nand U12535 (N_12535,N_12468,N_12005);
nor U12536 (N_12536,N_12402,N_12270);
and U12537 (N_12537,N_12496,N_12209);
xor U12538 (N_12538,N_12387,N_12418);
and U12539 (N_12539,N_12020,N_12228);
and U12540 (N_12540,N_12424,N_12189);
nor U12541 (N_12541,N_12124,N_12012);
xnor U12542 (N_12542,N_12349,N_12221);
or U12543 (N_12543,N_12346,N_12410);
xor U12544 (N_12544,N_12149,N_12227);
nor U12545 (N_12545,N_12330,N_12066);
nor U12546 (N_12546,N_12436,N_12059);
and U12547 (N_12547,N_12159,N_12146);
or U12548 (N_12548,N_12070,N_12040);
and U12549 (N_12549,N_12374,N_12166);
nor U12550 (N_12550,N_12431,N_12089);
or U12551 (N_12551,N_12026,N_12043);
or U12552 (N_12552,N_12126,N_12131);
nor U12553 (N_12553,N_12213,N_12193);
nor U12554 (N_12554,N_12113,N_12147);
nand U12555 (N_12555,N_12140,N_12063);
and U12556 (N_12556,N_12203,N_12044);
or U12557 (N_12557,N_12440,N_12022);
or U12558 (N_12558,N_12432,N_12214);
or U12559 (N_12559,N_12353,N_12328);
or U12560 (N_12560,N_12277,N_12407);
or U12561 (N_12561,N_12251,N_12036);
nand U12562 (N_12562,N_12487,N_12187);
nand U12563 (N_12563,N_12217,N_12139);
or U12564 (N_12564,N_12498,N_12460);
nor U12565 (N_12565,N_12456,N_12259);
and U12566 (N_12566,N_12458,N_12342);
or U12567 (N_12567,N_12401,N_12337);
xor U12568 (N_12568,N_12058,N_12151);
xor U12569 (N_12569,N_12205,N_12334);
or U12570 (N_12570,N_12076,N_12007);
or U12571 (N_12571,N_12038,N_12138);
or U12572 (N_12572,N_12361,N_12125);
or U12573 (N_12573,N_12162,N_12073);
nor U12574 (N_12574,N_12074,N_12031);
nor U12575 (N_12575,N_12307,N_12426);
xnor U12576 (N_12576,N_12042,N_12481);
and U12577 (N_12577,N_12274,N_12313);
nand U12578 (N_12578,N_12451,N_12144);
or U12579 (N_12579,N_12114,N_12380);
and U12580 (N_12580,N_12127,N_12148);
nor U12581 (N_12581,N_12317,N_12386);
and U12582 (N_12582,N_12208,N_12061);
and U12583 (N_12583,N_12196,N_12371);
and U12584 (N_12584,N_12108,N_12397);
nand U12585 (N_12585,N_12493,N_12072);
or U12586 (N_12586,N_12478,N_12260);
nand U12587 (N_12587,N_12429,N_12006);
or U12588 (N_12588,N_12321,N_12312);
or U12589 (N_12589,N_12485,N_12299);
and U12590 (N_12590,N_12320,N_12135);
nor U12591 (N_12591,N_12100,N_12335);
or U12592 (N_12592,N_12441,N_12134);
nand U12593 (N_12593,N_12204,N_12128);
nand U12594 (N_12594,N_12461,N_12098);
nand U12595 (N_12595,N_12230,N_12246);
or U12596 (N_12596,N_12102,N_12421);
xnor U12597 (N_12597,N_12293,N_12300);
and U12598 (N_12598,N_12264,N_12094);
nand U12599 (N_12599,N_12060,N_12428);
and U12600 (N_12600,N_12041,N_12409);
or U12601 (N_12601,N_12477,N_12046);
nand U12602 (N_12602,N_12240,N_12369);
and U12603 (N_12603,N_12014,N_12411);
and U12604 (N_12604,N_12261,N_12474);
nand U12605 (N_12605,N_12356,N_12381);
and U12606 (N_12606,N_12338,N_12430);
xor U12607 (N_12607,N_12311,N_12237);
xnor U12608 (N_12608,N_12165,N_12179);
xor U12609 (N_12609,N_12341,N_12155);
or U12610 (N_12610,N_12142,N_12010);
xnor U12611 (N_12611,N_12333,N_12123);
or U12612 (N_12612,N_12229,N_12202);
nand U12613 (N_12613,N_12292,N_12265);
xor U12614 (N_12614,N_12211,N_12198);
or U12615 (N_12615,N_12395,N_12071);
or U12616 (N_12616,N_12112,N_12082);
and U12617 (N_12617,N_12285,N_12011);
and U12618 (N_12618,N_12301,N_12078);
or U12619 (N_12619,N_12017,N_12178);
and U12620 (N_12620,N_12247,N_12174);
nor U12621 (N_12621,N_12352,N_12188);
nand U12622 (N_12622,N_12473,N_12169);
xnor U12623 (N_12623,N_12212,N_12105);
nor U12624 (N_12624,N_12236,N_12233);
nand U12625 (N_12625,N_12302,N_12281);
xnor U12626 (N_12626,N_12465,N_12258);
nor U12627 (N_12627,N_12053,N_12450);
or U12628 (N_12628,N_12110,N_12215);
and U12629 (N_12629,N_12479,N_12091);
xor U12630 (N_12630,N_12075,N_12490);
nor U12631 (N_12631,N_12122,N_12287);
nand U12632 (N_12632,N_12408,N_12153);
xor U12633 (N_12633,N_12488,N_12218);
and U12634 (N_12634,N_12201,N_12015);
xnor U12635 (N_12635,N_12294,N_12360);
nor U12636 (N_12636,N_12289,N_12455);
and U12637 (N_12637,N_12282,N_12154);
xor U12638 (N_12638,N_12457,N_12373);
xnor U12639 (N_12639,N_12482,N_12167);
and U12640 (N_12640,N_12183,N_12002);
and U12641 (N_12641,N_12389,N_12404);
xor U12642 (N_12642,N_12405,N_12400);
xor U12643 (N_12643,N_12045,N_12120);
nor U12644 (N_12644,N_12365,N_12003);
nor U12645 (N_12645,N_12284,N_12454);
nor U12646 (N_12646,N_12050,N_12069);
or U12647 (N_12647,N_12238,N_12362);
nand U12648 (N_12648,N_12051,N_12396);
nand U12649 (N_12649,N_12370,N_12034);
nand U12650 (N_12650,N_12472,N_12226);
nand U12651 (N_12651,N_12445,N_12152);
and U12652 (N_12652,N_12161,N_12173);
xor U12653 (N_12653,N_12029,N_12325);
nor U12654 (N_12654,N_12276,N_12297);
nor U12655 (N_12655,N_12250,N_12350);
xor U12656 (N_12656,N_12296,N_12298);
and U12657 (N_12657,N_12033,N_12262);
nor U12658 (N_12658,N_12171,N_12255);
or U12659 (N_12659,N_12241,N_12185);
nand U12660 (N_12660,N_12199,N_12336);
or U12661 (N_12661,N_12109,N_12470);
or U12662 (N_12662,N_12182,N_12326);
xor U12663 (N_12663,N_12057,N_12004);
xnor U12664 (N_12664,N_12375,N_12106);
xor U12665 (N_12665,N_12160,N_12025);
or U12666 (N_12666,N_12272,N_12434);
and U12667 (N_12667,N_12476,N_12433);
and U12668 (N_12668,N_12083,N_12239);
and U12669 (N_12669,N_12000,N_12480);
nand U12670 (N_12670,N_12175,N_12315);
nor U12671 (N_12671,N_12008,N_12095);
xor U12672 (N_12672,N_12207,N_12484);
or U12673 (N_12673,N_12268,N_12448);
or U12674 (N_12674,N_12027,N_12379);
nand U12675 (N_12675,N_12459,N_12039);
or U12676 (N_12676,N_12355,N_12273);
nor U12677 (N_12677,N_12013,N_12271);
xnor U12678 (N_12678,N_12345,N_12388);
xnor U12679 (N_12679,N_12425,N_12223);
xor U12680 (N_12680,N_12087,N_12449);
nand U12681 (N_12681,N_12168,N_12093);
nand U12682 (N_12682,N_12055,N_12366);
xor U12683 (N_12683,N_12435,N_12032);
xnor U12684 (N_12684,N_12367,N_12414);
nand U12685 (N_12685,N_12235,N_12107);
or U12686 (N_12686,N_12248,N_12288);
nand U12687 (N_12687,N_12024,N_12329);
and U12688 (N_12688,N_12181,N_12280);
nand U12689 (N_12689,N_12446,N_12420);
or U12690 (N_12690,N_12206,N_12332);
nor U12691 (N_12691,N_12049,N_12225);
and U12692 (N_12692,N_12382,N_12077);
xor U12693 (N_12693,N_12157,N_12219);
and U12694 (N_12694,N_12088,N_12111);
nand U12695 (N_12695,N_12132,N_12417);
xor U12696 (N_12696,N_12090,N_12121);
and U12697 (N_12697,N_12368,N_12234);
xnor U12698 (N_12698,N_12056,N_12391);
xor U12699 (N_12699,N_12466,N_12347);
xor U12700 (N_12700,N_12101,N_12164);
nor U12701 (N_12701,N_12453,N_12232);
and U12702 (N_12702,N_12309,N_12304);
xor U12703 (N_12703,N_12257,N_12143);
xnor U12704 (N_12704,N_12286,N_12021);
nand U12705 (N_12705,N_12319,N_12085);
and U12706 (N_12706,N_12385,N_12141);
xor U12707 (N_12707,N_12495,N_12494);
nand U12708 (N_12708,N_12191,N_12009);
xor U12709 (N_12709,N_12357,N_12254);
or U12710 (N_12710,N_12471,N_12359);
nor U12711 (N_12711,N_12463,N_12092);
nor U12712 (N_12712,N_12200,N_12406);
nand U12713 (N_12713,N_12403,N_12062);
nor U12714 (N_12714,N_12243,N_12364);
and U12715 (N_12715,N_12115,N_12310);
or U12716 (N_12716,N_12469,N_12447);
or U12717 (N_12717,N_12256,N_12439);
nand U12718 (N_12718,N_12028,N_12318);
and U12719 (N_12719,N_12295,N_12492);
nand U12720 (N_12720,N_12499,N_12096);
and U12721 (N_12721,N_12323,N_12018);
and U12722 (N_12722,N_12269,N_12392);
and U12723 (N_12723,N_12170,N_12266);
and U12724 (N_12724,N_12030,N_12220);
nor U12725 (N_12725,N_12384,N_12423);
nor U12726 (N_12726,N_12462,N_12279);
nand U12727 (N_12727,N_12079,N_12422);
xnor U12728 (N_12728,N_12097,N_12324);
nand U12729 (N_12729,N_12322,N_12305);
nor U12730 (N_12730,N_12443,N_12354);
and U12731 (N_12731,N_12242,N_12437);
or U12732 (N_12732,N_12194,N_12372);
nor U12733 (N_12733,N_12216,N_12483);
xor U12734 (N_12734,N_12308,N_12467);
xor U12735 (N_12735,N_12065,N_12231);
and U12736 (N_12736,N_12278,N_12118);
or U12737 (N_12737,N_12067,N_12497);
xnor U12738 (N_12738,N_12222,N_12145);
or U12739 (N_12739,N_12393,N_12343);
xor U12740 (N_12740,N_12344,N_12394);
and U12741 (N_12741,N_12116,N_12398);
nand U12742 (N_12742,N_12244,N_12099);
or U12743 (N_12743,N_12156,N_12348);
nor U12744 (N_12744,N_12130,N_12377);
xnor U12745 (N_12745,N_12180,N_12275);
nor U12746 (N_12746,N_12316,N_12163);
nand U12747 (N_12747,N_12351,N_12019);
nor U12748 (N_12748,N_12283,N_12054);
nor U12749 (N_12749,N_12245,N_12177);
and U12750 (N_12750,N_12310,N_12377);
nand U12751 (N_12751,N_12330,N_12311);
and U12752 (N_12752,N_12010,N_12086);
and U12753 (N_12753,N_12441,N_12299);
xor U12754 (N_12754,N_12298,N_12490);
xor U12755 (N_12755,N_12389,N_12062);
nand U12756 (N_12756,N_12110,N_12227);
or U12757 (N_12757,N_12314,N_12079);
nor U12758 (N_12758,N_12085,N_12174);
nand U12759 (N_12759,N_12220,N_12393);
xnor U12760 (N_12760,N_12294,N_12498);
and U12761 (N_12761,N_12205,N_12287);
and U12762 (N_12762,N_12096,N_12339);
xor U12763 (N_12763,N_12356,N_12067);
nor U12764 (N_12764,N_12196,N_12231);
nor U12765 (N_12765,N_12187,N_12196);
or U12766 (N_12766,N_12068,N_12200);
nand U12767 (N_12767,N_12482,N_12428);
xor U12768 (N_12768,N_12349,N_12387);
or U12769 (N_12769,N_12031,N_12446);
xor U12770 (N_12770,N_12428,N_12194);
nor U12771 (N_12771,N_12016,N_12492);
xnor U12772 (N_12772,N_12397,N_12186);
xnor U12773 (N_12773,N_12123,N_12083);
xnor U12774 (N_12774,N_12005,N_12419);
xnor U12775 (N_12775,N_12296,N_12345);
and U12776 (N_12776,N_12365,N_12335);
nor U12777 (N_12777,N_12375,N_12272);
xnor U12778 (N_12778,N_12120,N_12180);
nand U12779 (N_12779,N_12308,N_12330);
and U12780 (N_12780,N_12186,N_12399);
nand U12781 (N_12781,N_12059,N_12416);
and U12782 (N_12782,N_12299,N_12465);
nor U12783 (N_12783,N_12479,N_12201);
nor U12784 (N_12784,N_12270,N_12150);
or U12785 (N_12785,N_12314,N_12299);
or U12786 (N_12786,N_12385,N_12257);
nand U12787 (N_12787,N_12270,N_12458);
and U12788 (N_12788,N_12302,N_12038);
xnor U12789 (N_12789,N_12117,N_12418);
xor U12790 (N_12790,N_12232,N_12212);
nand U12791 (N_12791,N_12414,N_12450);
nor U12792 (N_12792,N_12228,N_12469);
or U12793 (N_12793,N_12091,N_12174);
or U12794 (N_12794,N_12492,N_12122);
nor U12795 (N_12795,N_12034,N_12221);
nand U12796 (N_12796,N_12211,N_12276);
or U12797 (N_12797,N_12478,N_12170);
xnor U12798 (N_12798,N_12068,N_12450);
nand U12799 (N_12799,N_12331,N_12483);
xnor U12800 (N_12800,N_12262,N_12378);
nand U12801 (N_12801,N_12179,N_12106);
and U12802 (N_12802,N_12138,N_12021);
nor U12803 (N_12803,N_12418,N_12043);
or U12804 (N_12804,N_12328,N_12329);
or U12805 (N_12805,N_12497,N_12206);
xor U12806 (N_12806,N_12247,N_12403);
and U12807 (N_12807,N_12445,N_12027);
and U12808 (N_12808,N_12399,N_12086);
xor U12809 (N_12809,N_12488,N_12327);
nor U12810 (N_12810,N_12481,N_12380);
nor U12811 (N_12811,N_12089,N_12324);
nor U12812 (N_12812,N_12245,N_12466);
xnor U12813 (N_12813,N_12271,N_12162);
or U12814 (N_12814,N_12368,N_12385);
nor U12815 (N_12815,N_12360,N_12122);
nand U12816 (N_12816,N_12306,N_12282);
nor U12817 (N_12817,N_12167,N_12076);
or U12818 (N_12818,N_12118,N_12043);
nand U12819 (N_12819,N_12469,N_12102);
xnor U12820 (N_12820,N_12220,N_12091);
nand U12821 (N_12821,N_12089,N_12053);
and U12822 (N_12822,N_12246,N_12200);
xor U12823 (N_12823,N_12292,N_12127);
nand U12824 (N_12824,N_12214,N_12238);
or U12825 (N_12825,N_12467,N_12007);
nor U12826 (N_12826,N_12499,N_12188);
and U12827 (N_12827,N_12289,N_12041);
xnor U12828 (N_12828,N_12401,N_12308);
and U12829 (N_12829,N_12192,N_12459);
nand U12830 (N_12830,N_12216,N_12259);
nand U12831 (N_12831,N_12307,N_12446);
or U12832 (N_12832,N_12022,N_12268);
nand U12833 (N_12833,N_12459,N_12261);
xnor U12834 (N_12834,N_12129,N_12174);
and U12835 (N_12835,N_12293,N_12364);
xor U12836 (N_12836,N_12143,N_12079);
and U12837 (N_12837,N_12128,N_12066);
nor U12838 (N_12838,N_12404,N_12377);
and U12839 (N_12839,N_12073,N_12053);
and U12840 (N_12840,N_12078,N_12198);
nor U12841 (N_12841,N_12275,N_12044);
or U12842 (N_12842,N_12391,N_12251);
xnor U12843 (N_12843,N_12060,N_12167);
and U12844 (N_12844,N_12435,N_12368);
nand U12845 (N_12845,N_12013,N_12169);
or U12846 (N_12846,N_12316,N_12136);
or U12847 (N_12847,N_12000,N_12383);
xor U12848 (N_12848,N_12443,N_12382);
or U12849 (N_12849,N_12451,N_12231);
and U12850 (N_12850,N_12246,N_12030);
nor U12851 (N_12851,N_12376,N_12040);
nand U12852 (N_12852,N_12113,N_12355);
xnor U12853 (N_12853,N_12266,N_12323);
nand U12854 (N_12854,N_12351,N_12084);
nor U12855 (N_12855,N_12435,N_12494);
nor U12856 (N_12856,N_12277,N_12440);
nor U12857 (N_12857,N_12473,N_12308);
or U12858 (N_12858,N_12187,N_12399);
and U12859 (N_12859,N_12231,N_12121);
xor U12860 (N_12860,N_12149,N_12191);
and U12861 (N_12861,N_12350,N_12266);
or U12862 (N_12862,N_12290,N_12296);
or U12863 (N_12863,N_12095,N_12260);
or U12864 (N_12864,N_12434,N_12188);
or U12865 (N_12865,N_12361,N_12035);
xor U12866 (N_12866,N_12039,N_12082);
nand U12867 (N_12867,N_12475,N_12456);
and U12868 (N_12868,N_12413,N_12472);
xnor U12869 (N_12869,N_12489,N_12407);
nand U12870 (N_12870,N_12172,N_12112);
xnor U12871 (N_12871,N_12362,N_12451);
nand U12872 (N_12872,N_12030,N_12237);
or U12873 (N_12873,N_12174,N_12405);
nand U12874 (N_12874,N_12099,N_12142);
nand U12875 (N_12875,N_12075,N_12015);
nand U12876 (N_12876,N_12293,N_12113);
xor U12877 (N_12877,N_12164,N_12200);
nand U12878 (N_12878,N_12452,N_12283);
nor U12879 (N_12879,N_12407,N_12405);
nor U12880 (N_12880,N_12347,N_12165);
nand U12881 (N_12881,N_12231,N_12158);
xor U12882 (N_12882,N_12182,N_12321);
nand U12883 (N_12883,N_12262,N_12365);
or U12884 (N_12884,N_12362,N_12007);
nand U12885 (N_12885,N_12238,N_12156);
nand U12886 (N_12886,N_12069,N_12060);
xor U12887 (N_12887,N_12127,N_12144);
nor U12888 (N_12888,N_12260,N_12304);
xor U12889 (N_12889,N_12104,N_12182);
nand U12890 (N_12890,N_12054,N_12115);
xnor U12891 (N_12891,N_12380,N_12033);
nand U12892 (N_12892,N_12372,N_12253);
xor U12893 (N_12893,N_12381,N_12105);
and U12894 (N_12894,N_12250,N_12343);
xnor U12895 (N_12895,N_12323,N_12041);
or U12896 (N_12896,N_12056,N_12184);
xnor U12897 (N_12897,N_12315,N_12136);
xnor U12898 (N_12898,N_12479,N_12308);
nand U12899 (N_12899,N_12151,N_12449);
and U12900 (N_12900,N_12220,N_12157);
nand U12901 (N_12901,N_12409,N_12053);
xnor U12902 (N_12902,N_12372,N_12396);
or U12903 (N_12903,N_12114,N_12384);
nor U12904 (N_12904,N_12169,N_12442);
xor U12905 (N_12905,N_12448,N_12288);
and U12906 (N_12906,N_12279,N_12346);
nand U12907 (N_12907,N_12108,N_12126);
nor U12908 (N_12908,N_12215,N_12124);
nor U12909 (N_12909,N_12267,N_12229);
xor U12910 (N_12910,N_12445,N_12279);
xor U12911 (N_12911,N_12331,N_12130);
nor U12912 (N_12912,N_12090,N_12067);
and U12913 (N_12913,N_12431,N_12399);
nor U12914 (N_12914,N_12214,N_12270);
xnor U12915 (N_12915,N_12475,N_12304);
nand U12916 (N_12916,N_12484,N_12139);
or U12917 (N_12917,N_12405,N_12137);
and U12918 (N_12918,N_12311,N_12294);
and U12919 (N_12919,N_12175,N_12193);
nand U12920 (N_12920,N_12383,N_12038);
or U12921 (N_12921,N_12259,N_12071);
nor U12922 (N_12922,N_12414,N_12412);
and U12923 (N_12923,N_12278,N_12029);
nand U12924 (N_12924,N_12268,N_12384);
xor U12925 (N_12925,N_12048,N_12155);
or U12926 (N_12926,N_12342,N_12147);
nor U12927 (N_12927,N_12433,N_12150);
or U12928 (N_12928,N_12209,N_12420);
nand U12929 (N_12929,N_12491,N_12277);
nor U12930 (N_12930,N_12225,N_12457);
nand U12931 (N_12931,N_12179,N_12448);
or U12932 (N_12932,N_12375,N_12072);
nand U12933 (N_12933,N_12234,N_12249);
or U12934 (N_12934,N_12397,N_12030);
and U12935 (N_12935,N_12215,N_12115);
or U12936 (N_12936,N_12386,N_12484);
nor U12937 (N_12937,N_12369,N_12247);
nand U12938 (N_12938,N_12310,N_12328);
nand U12939 (N_12939,N_12147,N_12225);
nor U12940 (N_12940,N_12063,N_12393);
xor U12941 (N_12941,N_12289,N_12038);
nand U12942 (N_12942,N_12494,N_12459);
nand U12943 (N_12943,N_12429,N_12062);
nor U12944 (N_12944,N_12232,N_12458);
nand U12945 (N_12945,N_12372,N_12425);
or U12946 (N_12946,N_12254,N_12437);
nand U12947 (N_12947,N_12025,N_12268);
nor U12948 (N_12948,N_12117,N_12052);
xor U12949 (N_12949,N_12083,N_12074);
nand U12950 (N_12950,N_12015,N_12056);
nand U12951 (N_12951,N_12159,N_12240);
xnor U12952 (N_12952,N_12114,N_12341);
or U12953 (N_12953,N_12315,N_12405);
nand U12954 (N_12954,N_12272,N_12489);
and U12955 (N_12955,N_12133,N_12452);
nor U12956 (N_12956,N_12441,N_12488);
xor U12957 (N_12957,N_12293,N_12430);
xor U12958 (N_12958,N_12401,N_12346);
or U12959 (N_12959,N_12026,N_12085);
xor U12960 (N_12960,N_12090,N_12259);
nor U12961 (N_12961,N_12328,N_12262);
nor U12962 (N_12962,N_12438,N_12379);
nor U12963 (N_12963,N_12028,N_12099);
xor U12964 (N_12964,N_12353,N_12116);
xnor U12965 (N_12965,N_12144,N_12431);
xnor U12966 (N_12966,N_12117,N_12219);
or U12967 (N_12967,N_12383,N_12267);
xor U12968 (N_12968,N_12200,N_12077);
xor U12969 (N_12969,N_12028,N_12097);
and U12970 (N_12970,N_12099,N_12419);
nand U12971 (N_12971,N_12402,N_12264);
xnor U12972 (N_12972,N_12305,N_12400);
xnor U12973 (N_12973,N_12342,N_12201);
nand U12974 (N_12974,N_12492,N_12253);
and U12975 (N_12975,N_12450,N_12124);
xnor U12976 (N_12976,N_12254,N_12158);
or U12977 (N_12977,N_12050,N_12415);
or U12978 (N_12978,N_12456,N_12200);
nor U12979 (N_12979,N_12014,N_12259);
nor U12980 (N_12980,N_12168,N_12275);
nor U12981 (N_12981,N_12161,N_12307);
or U12982 (N_12982,N_12225,N_12484);
nand U12983 (N_12983,N_12326,N_12095);
nand U12984 (N_12984,N_12409,N_12304);
xor U12985 (N_12985,N_12072,N_12196);
or U12986 (N_12986,N_12097,N_12376);
xnor U12987 (N_12987,N_12084,N_12183);
xnor U12988 (N_12988,N_12282,N_12247);
or U12989 (N_12989,N_12434,N_12005);
xor U12990 (N_12990,N_12434,N_12159);
nor U12991 (N_12991,N_12463,N_12458);
and U12992 (N_12992,N_12466,N_12417);
and U12993 (N_12993,N_12079,N_12341);
or U12994 (N_12994,N_12315,N_12458);
or U12995 (N_12995,N_12413,N_12133);
nand U12996 (N_12996,N_12115,N_12105);
and U12997 (N_12997,N_12370,N_12192);
xnor U12998 (N_12998,N_12091,N_12316);
and U12999 (N_12999,N_12057,N_12254);
or U13000 (N_13000,N_12995,N_12635);
nand U13001 (N_13001,N_12863,N_12557);
nor U13002 (N_13002,N_12563,N_12924);
nor U13003 (N_13003,N_12744,N_12939);
nor U13004 (N_13004,N_12595,N_12884);
and U13005 (N_13005,N_12773,N_12653);
or U13006 (N_13006,N_12975,N_12720);
or U13007 (N_13007,N_12928,N_12614);
and U13008 (N_13008,N_12938,N_12901);
and U13009 (N_13009,N_12840,N_12687);
or U13010 (N_13010,N_12780,N_12997);
and U13011 (N_13011,N_12526,N_12979);
and U13012 (N_13012,N_12971,N_12804);
or U13013 (N_13013,N_12588,N_12564);
or U13014 (N_13014,N_12590,N_12655);
nand U13015 (N_13015,N_12981,N_12959);
or U13016 (N_13016,N_12611,N_12560);
nand U13017 (N_13017,N_12820,N_12775);
or U13018 (N_13018,N_12838,N_12945);
and U13019 (N_13019,N_12671,N_12865);
nor U13020 (N_13020,N_12950,N_12629);
nand U13021 (N_13021,N_12509,N_12737);
and U13022 (N_13022,N_12692,N_12507);
nor U13023 (N_13023,N_12679,N_12736);
or U13024 (N_13024,N_12685,N_12941);
nand U13025 (N_13025,N_12639,N_12801);
nand U13026 (N_13026,N_12962,N_12841);
nand U13027 (N_13027,N_12721,N_12643);
xnor U13028 (N_13028,N_12880,N_12922);
nand U13029 (N_13029,N_12872,N_12828);
xor U13030 (N_13030,N_12681,N_12920);
or U13031 (N_13031,N_12553,N_12642);
nor U13032 (N_13032,N_12836,N_12790);
and U13033 (N_13033,N_12559,N_12600);
xnor U13034 (N_13034,N_12711,N_12667);
xor U13035 (N_13035,N_12532,N_12960);
and U13036 (N_13036,N_12758,N_12571);
nand U13037 (N_13037,N_12527,N_12967);
nand U13038 (N_13038,N_12934,N_12662);
xor U13039 (N_13039,N_12911,N_12965);
nand U13040 (N_13040,N_12796,N_12558);
and U13041 (N_13041,N_12786,N_12550);
and U13042 (N_13042,N_12803,N_12594);
nor U13043 (N_13043,N_12705,N_12634);
xnor U13044 (N_13044,N_12624,N_12751);
nand U13045 (N_13045,N_12940,N_12556);
nor U13046 (N_13046,N_12930,N_12536);
nand U13047 (N_13047,N_12622,N_12544);
xnor U13048 (N_13048,N_12718,N_12715);
and U13049 (N_13049,N_12889,N_12937);
nand U13050 (N_13050,N_12907,N_12980);
nor U13051 (N_13051,N_12579,N_12759);
nor U13052 (N_13052,N_12998,N_12730);
or U13053 (N_13053,N_12762,N_12593);
nor U13054 (N_13054,N_12787,N_12973);
nor U13055 (N_13055,N_12910,N_12645);
nor U13056 (N_13056,N_12764,N_12996);
nand U13057 (N_13057,N_12626,N_12505);
nand U13058 (N_13058,N_12688,N_12742);
and U13059 (N_13059,N_12848,N_12649);
or U13060 (N_13060,N_12956,N_12784);
xnor U13061 (N_13061,N_12504,N_12983);
or U13062 (N_13062,N_12750,N_12729);
xnor U13063 (N_13063,N_12931,N_12621);
nand U13064 (N_13064,N_12680,N_12670);
xor U13065 (N_13065,N_12761,N_12968);
nand U13066 (N_13066,N_12943,N_12904);
xor U13067 (N_13067,N_12716,N_12808);
or U13068 (N_13068,N_12854,N_12619);
and U13069 (N_13069,N_12748,N_12990);
xor U13070 (N_13070,N_12502,N_12807);
nand U13071 (N_13071,N_12881,N_12800);
nor U13072 (N_13072,N_12599,N_12949);
xnor U13073 (N_13073,N_12731,N_12749);
and U13074 (N_13074,N_12852,N_12704);
xor U13075 (N_13075,N_12540,N_12942);
or U13076 (N_13076,N_12678,N_12978);
nand U13077 (N_13077,N_12992,N_12798);
xnor U13078 (N_13078,N_12900,N_12699);
xnor U13079 (N_13079,N_12517,N_12914);
and U13080 (N_13080,N_12974,N_12581);
and U13081 (N_13081,N_12876,N_12972);
nand U13082 (N_13082,N_12646,N_12933);
nor U13083 (N_13083,N_12651,N_12893);
or U13084 (N_13084,N_12617,N_12637);
nand U13085 (N_13085,N_12862,N_12586);
xor U13086 (N_13086,N_12991,N_12948);
or U13087 (N_13087,N_12506,N_12817);
nor U13088 (N_13088,N_12732,N_12908);
or U13089 (N_13089,N_12955,N_12897);
nor U13090 (N_13090,N_12896,N_12735);
or U13091 (N_13091,N_12603,N_12669);
xnor U13092 (N_13092,N_12944,N_12714);
or U13093 (N_13093,N_12562,N_12812);
or U13094 (N_13094,N_12584,N_12832);
xnor U13095 (N_13095,N_12551,N_12977);
xor U13096 (N_13096,N_12608,N_12964);
nand U13097 (N_13097,N_12636,N_12576);
and U13098 (N_13098,N_12604,N_12906);
nand U13099 (N_13099,N_12878,N_12976);
xor U13100 (N_13100,N_12641,N_12805);
or U13101 (N_13101,N_12706,N_12696);
and U13102 (N_13102,N_12849,N_12923);
nand U13103 (N_13103,N_12886,N_12674);
nor U13104 (N_13104,N_12697,N_12548);
xor U13105 (N_13105,N_12754,N_12885);
and U13106 (N_13106,N_12850,N_12902);
xor U13107 (N_13107,N_12961,N_12656);
xnor U13108 (N_13108,N_12779,N_12592);
xor U13109 (N_13109,N_12567,N_12665);
or U13110 (N_13110,N_12632,N_12745);
and U13111 (N_13111,N_12830,N_12606);
xnor U13112 (N_13112,N_12768,N_12726);
nand U13113 (N_13113,N_12905,N_12628);
or U13114 (N_13114,N_12657,N_12609);
xor U13115 (N_13115,N_12503,N_12508);
or U13116 (N_13116,N_12575,N_12763);
nand U13117 (N_13117,N_12733,N_12501);
xor U13118 (N_13118,N_12554,N_12539);
xor U13119 (N_13119,N_12756,N_12822);
or U13120 (N_13120,N_12932,N_12515);
nor U13121 (N_13121,N_12587,N_12627);
nand U13122 (N_13122,N_12895,N_12658);
nand U13123 (N_13123,N_12882,N_12666);
nor U13124 (N_13124,N_12698,N_12694);
nor U13125 (N_13125,N_12861,N_12710);
xor U13126 (N_13126,N_12552,N_12788);
xnor U13127 (N_13127,N_12925,N_12695);
nor U13128 (N_13128,N_12534,N_12597);
nor U13129 (N_13129,N_12859,N_12953);
or U13130 (N_13130,N_12811,N_12612);
xnor U13131 (N_13131,N_12774,N_12545);
or U13132 (N_13132,N_12985,N_12668);
nor U13133 (N_13133,N_12578,N_12982);
nor U13134 (N_13134,N_12712,N_12633);
or U13135 (N_13135,N_12677,N_12568);
xnor U13136 (N_13136,N_12989,N_12707);
nand U13137 (N_13137,N_12821,N_12566);
nand U13138 (N_13138,N_12647,N_12858);
xnor U13139 (N_13139,N_12638,N_12512);
xnor U13140 (N_13140,N_12855,N_12814);
xnor U13141 (N_13141,N_12969,N_12722);
nand U13142 (N_13142,N_12792,N_12795);
or U13143 (N_13143,N_12834,N_12672);
or U13144 (N_13144,N_12570,N_12625);
or U13145 (N_13145,N_12868,N_12951);
nand U13146 (N_13146,N_12823,N_12760);
and U13147 (N_13147,N_12912,N_12815);
nand U13148 (N_13148,N_12739,N_12782);
nand U13149 (N_13149,N_12755,N_12853);
or U13150 (N_13150,N_12987,N_12644);
and U13151 (N_13151,N_12778,N_12824);
or U13152 (N_13152,N_12802,N_12675);
xnor U13153 (N_13153,N_12913,N_12500);
or U13154 (N_13154,N_12719,N_12767);
nand U13155 (N_13155,N_12877,N_12766);
nand U13156 (N_13156,N_12577,N_12874);
and U13157 (N_13157,N_12518,N_12869);
nand U13158 (N_13158,N_12631,N_12839);
and U13159 (N_13159,N_12591,N_12819);
nand U13160 (N_13160,N_12918,N_12607);
or U13161 (N_13161,N_12569,N_12806);
and U13162 (N_13162,N_12986,N_12957);
or U13163 (N_13163,N_12522,N_12521);
nor U13164 (N_13164,N_12988,N_12542);
xor U13165 (N_13165,N_12583,N_12528);
nand U13166 (N_13166,N_12511,N_12873);
nor U13167 (N_13167,N_12724,N_12531);
nor U13168 (N_13168,N_12999,N_12818);
nand U13169 (N_13169,N_12602,N_12516);
nor U13170 (N_13170,N_12827,N_12851);
xnor U13171 (N_13171,N_12682,N_12741);
and U13172 (N_13172,N_12894,N_12615);
or U13173 (N_13173,N_12809,N_12776);
xor U13174 (N_13174,N_12860,N_12689);
and U13175 (N_13175,N_12966,N_12867);
nor U13176 (N_13176,N_12752,N_12845);
xor U13177 (N_13177,N_12525,N_12630);
nor U13178 (N_13178,N_12623,N_12921);
nand U13179 (N_13179,N_12984,N_12535);
xnor U13180 (N_13180,N_12856,N_12746);
or U13181 (N_13181,N_12797,N_12582);
xor U13182 (N_13182,N_12572,N_12700);
and U13183 (N_13183,N_12772,N_12728);
and U13184 (N_13184,N_12793,N_12529);
nand U13185 (N_13185,N_12654,N_12813);
xor U13186 (N_13186,N_12747,N_12866);
or U13187 (N_13187,N_12713,N_12601);
and U13188 (N_13188,N_12777,N_12618);
xnor U13189 (N_13189,N_12909,N_12791);
xor U13190 (N_13190,N_12514,N_12616);
and U13191 (N_13191,N_12783,N_12829);
xor U13192 (N_13192,N_12701,N_12541);
nor U13193 (N_13193,N_12650,N_12844);
and U13194 (N_13194,N_12826,N_12640);
xor U13195 (N_13195,N_12598,N_12993);
and U13196 (N_13196,N_12958,N_12947);
or U13197 (N_13197,N_12919,N_12898);
nand U13198 (N_13198,N_12530,N_12843);
and U13199 (N_13199,N_12652,N_12709);
nor U13200 (N_13200,N_12875,N_12927);
nand U13201 (N_13201,N_12952,N_12660);
and U13202 (N_13202,N_12613,N_12676);
and U13203 (N_13203,N_12847,N_12725);
nor U13204 (N_13204,N_12580,N_12963);
nor U13205 (N_13205,N_12693,N_12871);
nor U13206 (N_13206,N_12543,N_12717);
nor U13207 (N_13207,N_12753,N_12864);
or U13208 (N_13208,N_12870,N_12520);
nor U13209 (N_13209,N_12887,N_12661);
nor U13210 (N_13210,N_12994,N_12890);
nand U13211 (N_13211,N_12831,N_12757);
nand U13212 (N_13212,N_12589,N_12596);
or U13213 (N_13213,N_12835,N_12523);
and U13214 (N_13214,N_12903,N_12538);
or U13215 (N_13215,N_12664,N_12799);
or U13216 (N_13216,N_12703,N_12574);
and U13217 (N_13217,N_12702,N_12892);
and U13218 (N_13218,N_12565,N_12781);
and U13219 (N_13219,N_12683,N_12555);
nand U13220 (N_13220,N_12561,N_12769);
and U13221 (N_13221,N_12765,N_12946);
nand U13222 (N_13222,N_12620,N_12743);
nor U13223 (N_13223,N_12794,N_12857);
nor U13224 (N_13224,N_12659,N_12610);
and U13225 (N_13225,N_12684,N_12842);
nand U13226 (N_13226,N_12810,N_12690);
and U13227 (N_13227,N_12936,N_12708);
xnor U13228 (N_13228,N_12929,N_12519);
or U13229 (N_13229,N_12916,N_12883);
and U13230 (N_13230,N_12510,N_12816);
or U13231 (N_13231,N_12585,N_12546);
or U13232 (N_13232,N_12513,N_12663);
and U13233 (N_13233,N_12573,N_12771);
and U13234 (N_13234,N_12734,N_12537);
nand U13235 (N_13235,N_12846,N_12648);
and U13236 (N_13236,N_12888,N_12549);
nor U13237 (N_13237,N_12673,N_12891);
or U13238 (N_13238,N_12970,N_12789);
and U13239 (N_13239,N_12605,N_12740);
nor U13240 (N_13240,N_12935,N_12533);
and U13241 (N_13241,N_12825,N_12954);
and U13242 (N_13242,N_12547,N_12686);
nor U13243 (N_13243,N_12785,N_12524);
nor U13244 (N_13244,N_12915,N_12926);
and U13245 (N_13245,N_12723,N_12899);
and U13246 (N_13246,N_12691,N_12917);
xnor U13247 (N_13247,N_12738,N_12770);
nand U13248 (N_13248,N_12727,N_12833);
xnor U13249 (N_13249,N_12837,N_12879);
nor U13250 (N_13250,N_12757,N_12991);
and U13251 (N_13251,N_12643,N_12574);
xor U13252 (N_13252,N_12792,N_12884);
xnor U13253 (N_13253,N_12675,N_12556);
and U13254 (N_13254,N_12585,N_12788);
xor U13255 (N_13255,N_12623,N_12526);
nand U13256 (N_13256,N_12592,N_12812);
nand U13257 (N_13257,N_12517,N_12838);
xnor U13258 (N_13258,N_12739,N_12691);
and U13259 (N_13259,N_12600,N_12942);
or U13260 (N_13260,N_12809,N_12681);
and U13261 (N_13261,N_12545,N_12710);
nand U13262 (N_13262,N_12840,N_12596);
xor U13263 (N_13263,N_12764,N_12963);
nor U13264 (N_13264,N_12882,N_12704);
xnor U13265 (N_13265,N_12577,N_12527);
xnor U13266 (N_13266,N_12958,N_12502);
or U13267 (N_13267,N_12948,N_12753);
and U13268 (N_13268,N_12883,N_12851);
nand U13269 (N_13269,N_12982,N_12693);
or U13270 (N_13270,N_12733,N_12522);
nor U13271 (N_13271,N_12964,N_12603);
xor U13272 (N_13272,N_12530,N_12798);
nand U13273 (N_13273,N_12965,N_12879);
or U13274 (N_13274,N_12628,N_12646);
nand U13275 (N_13275,N_12923,N_12698);
nand U13276 (N_13276,N_12589,N_12627);
nor U13277 (N_13277,N_12803,N_12959);
and U13278 (N_13278,N_12808,N_12962);
and U13279 (N_13279,N_12514,N_12620);
or U13280 (N_13280,N_12825,N_12829);
nor U13281 (N_13281,N_12966,N_12604);
or U13282 (N_13282,N_12798,N_12809);
xnor U13283 (N_13283,N_12820,N_12556);
nand U13284 (N_13284,N_12516,N_12776);
or U13285 (N_13285,N_12661,N_12918);
xor U13286 (N_13286,N_12921,N_12747);
xor U13287 (N_13287,N_12723,N_12554);
or U13288 (N_13288,N_12636,N_12620);
nand U13289 (N_13289,N_12613,N_12538);
or U13290 (N_13290,N_12953,N_12950);
or U13291 (N_13291,N_12628,N_12620);
nand U13292 (N_13292,N_12854,N_12747);
nor U13293 (N_13293,N_12692,N_12591);
and U13294 (N_13294,N_12588,N_12749);
nand U13295 (N_13295,N_12915,N_12987);
and U13296 (N_13296,N_12738,N_12979);
and U13297 (N_13297,N_12967,N_12955);
and U13298 (N_13298,N_12863,N_12567);
nor U13299 (N_13299,N_12685,N_12960);
and U13300 (N_13300,N_12511,N_12671);
nor U13301 (N_13301,N_12662,N_12865);
nor U13302 (N_13302,N_12727,N_12731);
nand U13303 (N_13303,N_12877,N_12931);
xor U13304 (N_13304,N_12704,N_12858);
or U13305 (N_13305,N_12657,N_12592);
xnor U13306 (N_13306,N_12856,N_12940);
and U13307 (N_13307,N_12726,N_12663);
or U13308 (N_13308,N_12739,N_12753);
xor U13309 (N_13309,N_12800,N_12858);
or U13310 (N_13310,N_12915,N_12956);
nand U13311 (N_13311,N_12886,N_12947);
or U13312 (N_13312,N_12873,N_12520);
or U13313 (N_13313,N_12729,N_12942);
and U13314 (N_13314,N_12738,N_12736);
nand U13315 (N_13315,N_12925,N_12941);
nand U13316 (N_13316,N_12719,N_12940);
xor U13317 (N_13317,N_12640,N_12750);
xnor U13318 (N_13318,N_12590,N_12532);
and U13319 (N_13319,N_12694,N_12812);
or U13320 (N_13320,N_12793,N_12579);
xnor U13321 (N_13321,N_12588,N_12700);
nand U13322 (N_13322,N_12714,N_12893);
nor U13323 (N_13323,N_12637,N_12894);
nand U13324 (N_13324,N_12974,N_12890);
nor U13325 (N_13325,N_12770,N_12922);
nor U13326 (N_13326,N_12772,N_12976);
and U13327 (N_13327,N_12752,N_12508);
nor U13328 (N_13328,N_12538,N_12611);
or U13329 (N_13329,N_12827,N_12504);
nor U13330 (N_13330,N_12630,N_12959);
nand U13331 (N_13331,N_12819,N_12820);
nor U13332 (N_13332,N_12615,N_12607);
or U13333 (N_13333,N_12965,N_12874);
xor U13334 (N_13334,N_12792,N_12507);
or U13335 (N_13335,N_12953,N_12947);
or U13336 (N_13336,N_12972,N_12624);
and U13337 (N_13337,N_12695,N_12515);
xnor U13338 (N_13338,N_12638,N_12912);
and U13339 (N_13339,N_12618,N_12617);
nand U13340 (N_13340,N_12572,N_12774);
nand U13341 (N_13341,N_12516,N_12829);
nor U13342 (N_13342,N_12642,N_12882);
or U13343 (N_13343,N_12683,N_12900);
xnor U13344 (N_13344,N_12857,N_12694);
xor U13345 (N_13345,N_12519,N_12737);
or U13346 (N_13346,N_12565,N_12544);
nor U13347 (N_13347,N_12504,N_12760);
nand U13348 (N_13348,N_12620,N_12776);
nor U13349 (N_13349,N_12555,N_12800);
nor U13350 (N_13350,N_12835,N_12842);
nand U13351 (N_13351,N_12509,N_12570);
nand U13352 (N_13352,N_12523,N_12799);
xnor U13353 (N_13353,N_12540,N_12965);
nor U13354 (N_13354,N_12774,N_12603);
or U13355 (N_13355,N_12540,N_12782);
or U13356 (N_13356,N_12639,N_12557);
xnor U13357 (N_13357,N_12797,N_12847);
and U13358 (N_13358,N_12502,N_12903);
and U13359 (N_13359,N_12790,N_12534);
nand U13360 (N_13360,N_12673,N_12515);
or U13361 (N_13361,N_12787,N_12771);
nand U13362 (N_13362,N_12577,N_12722);
xnor U13363 (N_13363,N_12643,N_12903);
xnor U13364 (N_13364,N_12636,N_12767);
xnor U13365 (N_13365,N_12730,N_12797);
xor U13366 (N_13366,N_12921,N_12666);
nor U13367 (N_13367,N_12532,N_12950);
xnor U13368 (N_13368,N_12866,N_12833);
nand U13369 (N_13369,N_12748,N_12940);
xor U13370 (N_13370,N_12643,N_12797);
nor U13371 (N_13371,N_12836,N_12638);
nand U13372 (N_13372,N_12817,N_12965);
nand U13373 (N_13373,N_12647,N_12967);
nor U13374 (N_13374,N_12746,N_12581);
xor U13375 (N_13375,N_12670,N_12903);
nand U13376 (N_13376,N_12516,N_12523);
xor U13377 (N_13377,N_12614,N_12602);
nand U13378 (N_13378,N_12787,N_12583);
nand U13379 (N_13379,N_12558,N_12618);
xnor U13380 (N_13380,N_12752,N_12667);
and U13381 (N_13381,N_12766,N_12642);
xor U13382 (N_13382,N_12576,N_12868);
and U13383 (N_13383,N_12985,N_12926);
or U13384 (N_13384,N_12721,N_12607);
nand U13385 (N_13385,N_12552,N_12532);
or U13386 (N_13386,N_12505,N_12805);
nand U13387 (N_13387,N_12637,N_12641);
nor U13388 (N_13388,N_12586,N_12563);
nand U13389 (N_13389,N_12760,N_12578);
xor U13390 (N_13390,N_12770,N_12521);
xnor U13391 (N_13391,N_12758,N_12874);
and U13392 (N_13392,N_12591,N_12945);
and U13393 (N_13393,N_12636,N_12523);
nor U13394 (N_13394,N_12950,N_12534);
nor U13395 (N_13395,N_12812,N_12977);
xnor U13396 (N_13396,N_12501,N_12902);
nor U13397 (N_13397,N_12563,N_12589);
nand U13398 (N_13398,N_12510,N_12532);
nand U13399 (N_13399,N_12653,N_12601);
nor U13400 (N_13400,N_12741,N_12779);
nor U13401 (N_13401,N_12658,N_12500);
xnor U13402 (N_13402,N_12642,N_12720);
nor U13403 (N_13403,N_12610,N_12648);
and U13404 (N_13404,N_12777,N_12901);
xnor U13405 (N_13405,N_12877,N_12743);
nand U13406 (N_13406,N_12695,N_12674);
and U13407 (N_13407,N_12940,N_12904);
xor U13408 (N_13408,N_12978,N_12927);
and U13409 (N_13409,N_12820,N_12648);
nor U13410 (N_13410,N_12714,N_12799);
and U13411 (N_13411,N_12664,N_12606);
or U13412 (N_13412,N_12944,N_12872);
nand U13413 (N_13413,N_12679,N_12904);
nand U13414 (N_13414,N_12791,N_12517);
or U13415 (N_13415,N_12796,N_12617);
nand U13416 (N_13416,N_12805,N_12960);
nand U13417 (N_13417,N_12819,N_12922);
or U13418 (N_13418,N_12904,N_12715);
nand U13419 (N_13419,N_12606,N_12642);
nand U13420 (N_13420,N_12991,N_12916);
and U13421 (N_13421,N_12584,N_12572);
and U13422 (N_13422,N_12767,N_12510);
nor U13423 (N_13423,N_12520,N_12806);
and U13424 (N_13424,N_12833,N_12606);
nand U13425 (N_13425,N_12571,N_12646);
or U13426 (N_13426,N_12846,N_12620);
or U13427 (N_13427,N_12707,N_12548);
nand U13428 (N_13428,N_12628,N_12788);
nand U13429 (N_13429,N_12746,N_12571);
and U13430 (N_13430,N_12623,N_12741);
or U13431 (N_13431,N_12806,N_12970);
xnor U13432 (N_13432,N_12582,N_12638);
nand U13433 (N_13433,N_12800,N_12854);
nand U13434 (N_13434,N_12671,N_12683);
nand U13435 (N_13435,N_12706,N_12702);
nor U13436 (N_13436,N_12891,N_12529);
or U13437 (N_13437,N_12908,N_12694);
nand U13438 (N_13438,N_12843,N_12697);
xor U13439 (N_13439,N_12764,N_12818);
and U13440 (N_13440,N_12956,N_12855);
nand U13441 (N_13441,N_12828,N_12681);
and U13442 (N_13442,N_12898,N_12589);
nand U13443 (N_13443,N_12533,N_12632);
xnor U13444 (N_13444,N_12564,N_12956);
nand U13445 (N_13445,N_12953,N_12790);
nor U13446 (N_13446,N_12722,N_12971);
and U13447 (N_13447,N_12804,N_12909);
and U13448 (N_13448,N_12629,N_12580);
nor U13449 (N_13449,N_12669,N_12799);
nand U13450 (N_13450,N_12802,N_12649);
nand U13451 (N_13451,N_12823,N_12660);
or U13452 (N_13452,N_12755,N_12945);
nor U13453 (N_13453,N_12658,N_12939);
or U13454 (N_13454,N_12871,N_12787);
and U13455 (N_13455,N_12961,N_12511);
and U13456 (N_13456,N_12728,N_12586);
or U13457 (N_13457,N_12544,N_12633);
nand U13458 (N_13458,N_12950,N_12979);
xnor U13459 (N_13459,N_12536,N_12524);
xor U13460 (N_13460,N_12875,N_12919);
and U13461 (N_13461,N_12545,N_12819);
xor U13462 (N_13462,N_12983,N_12828);
nor U13463 (N_13463,N_12635,N_12664);
nand U13464 (N_13464,N_12751,N_12747);
and U13465 (N_13465,N_12766,N_12885);
and U13466 (N_13466,N_12801,N_12643);
nand U13467 (N_13467,N_12900,N_12867);
or U13468 (N_13468,N_12900,N_12696);
nand U13469 (N_13469,N_12518,N_12998);
or U13470 (N_13470,N_12920,N_12899);
nand U13471 (N_13471,N_12813,N_12820);
xnor U13472 (N_13472,N_12591,N_12779);
xor U13473 (N_13473,N_12902,N_12543);
nor U13474 (N_13474,N_12904,N_12581);
xnor U13475 (N_13475,N_12899,N_12708);
nand U13476 (N_13476,N_12726,N_12538);
nor U13477 (N_13477,N_12554,N_12760);
nor U13478 (N_13478,N_12749,N_12805);
nor U13479 (N_13479,N_12941,N_12596);
nand U13480 (N_13480,N_12948,N_12523);
and U13481 (N_13481,N_12511,N_12613);
or U13482 (N_13482,N_12941,N_12541);
or U13483 (N_13483,N_12615,N_12999);
nand U13484 (N_13484,N_12789,N_12786);
nand U13485 (N_13485,N_12858,N_12797);
or U13486 (N_13486,N_12601,N_12616);
and U13487 (N_13487,N_12940,N_12660);
and U13488 (N_13488,N_12957,N_12626);
nand U13489 (N_13489,N_12918,N_12612);
xor U13490 (N_13490,N_12626,N_12801);
and U13491 (N_13491,N_12556,N_12515);
nor U13492 (N_13492,N_12693,N_12712);
nor U13493 (N_13493,N_12851,N_12602);
and U13494 (N_13494,N_12933,N_12898);
nor U13495 (N_13495,N_12765,N_12809);
or U13496 (N_13496,N_12867,N_12958);
nor U13497 (N_13497,N_12993,N_12549);
and U13498 (N_13498,N_12564,N_12943);
or U13499 (N_13499,N_12823,N_12969);
nand U13500 (N_13500,N_13273,N_13081);
nor U13501 (N_13501,N_13169,N_13205);
or U13502 (N_13502,N_13385,N_13298);
xnor U13503 (N_13503,N_13319,N_13292);
xor U13504 (N_13504,N_13410,N_13179);
or U13505 (N_13505,N_13208,N_13226);
nand U13506 (N_13506,N_13204,N_13196);
nor U13507 (N_13507,N_13177,N_13009);
xnor U13508 (N_13508,N_13444,N_13098);
xor U13509 (N_13509,N_13291,N_13035);
nor U13510 (N_13510,N_13055,N_13408);
and U13511 (N_13511,N_13371,N_13173);
and U13512 (N_13512,N_13224,N_13010);
and U13513 (N_13513,N_13090,N_13360);
or U13514 (N_13514,N_13482,N_13181);
and U13515 (N_13515,N_13490,N_13282);
nor U13516 (N_13516,N_13242,N_13419);
nor U13517 (N_13517,N_13341,N_13174);
nor U13518 (N_13518,N_13237,N_13138);
or U13519 (N_13519,N_13150,N_13072);
nor U13520 (N_13520,N_13347,N_13143);
nand U13521 (N_13521,N_13076,N_13175);
nand U13522 (N_13522,N_13266,N_13418);
or U13523 (N_13523,N_13421,N_13002);
xnor U13524 (N_13524,N_13469,N_13137);
nand U13525 (N_13525,N_13272,N_13032);
nor U13526 (N_13526,N_13440,N_13331);
nor U13527 (N_13527,N_13160,N_13313);
xnor U13528 (N_13528,N_13463,N_13489);
xnor U13529 (N_13529,N_13267,N_13301);
and U13530 (N_13530,N_13077,N_13379);
and U13531 (N_13531,N_13353,N_13052);
nor U13532 (N_13532,N_13369,N_13387);
nor U13533 (N_13533,N_13258,N_13212);
nor U13534 (N_13534,N_13484,N_13193);
nor U13535 (N_13535,N_13308,N_13039);
nor U13536 (N_13536,N_13265,N_13280);
or U13537 (N_13537,N_13164,N_13498);
xor U13538 (N_13538,N_13136,N_13453);
nand U13539 (N_13539,N_13108,N_13378);
nor U13540 (N_13540,N_13465,N_13185);
nor U13541 (N_13541,N_13405,N_13257);
nand U13542 (N_13542,N_13167,N_13183);
and U13543 (N_13543,N_13247,N_13470);
xor U13544 (N_13544,N_13261,N_13097);
xor U13545 (N_13545,N_13485,N_13404);
and U13546 (N_13546,N_13399,N_13071);
xor U13547 (N_13547,N_13094,N_13320);
xnor U13548 (N_13548,N_13087,N_13023);
or U13549 (N_13549,N_13244,N_13445);
nand U13550 (N_13550,N_13386,N_13065);
xnor U13551 (N_13551,N_13284,N_13295);
nor U13552 (N_13552,N_13105,N_13102);
or U13553 (N_13553,N_13434,N_13158);
nor U13554 (N_13554,N_13134,N_13152);
nor U13555 (N_13555,N_13423,N_13277);
xor U13556 (N_13556,N_13232,N_13088);
xnor U13557 (N_13557,N_13154,N_13384);
nand U13558 (N_13558,N_13229,N_13262);
and U13559 (N_13559,N_13159,N_13231);
and U13560 (N_13560,N_13031,N_13011);
nor U13561 (N_13561,N_13316,N_13122);
or U13562 (N_13562,N_13448,N_13178);
nor U13563 (N_13563,N_13468,N_13307);
nor U13564 (N_13564,N_13142,N_13441);
nor U13565 (N_13565,N_13157,N_13328);
and U13566 (N_13566,N_13424,N_13220);
xnor U13567 (N_13567,N_13491,N_13367);
xnor U13568 (N_13568,N_13104,N_13171);
xor U13569 (N_13569,N_13117,N_13151);
and U13570 (N_13570,N_13051,N_13390);
and U13571 (N_13571,N_13056,N_13343);
xor U13572 (N_13572,N_13166,N_13275);
xor U13573 (N_13573,N_13001,N_13141);
and U13574 (N_13574,N_13462,N_13380);
or U13575 (N_13575,N_13078,N_13344);
xor U13576 (N_13576,N_13372,N_13354);
nand U13577 (N_13577,N_13330,N_13206);
xnor U13578 (N_13578,N_13398,N_13082);
xor U13579 (N_13579,N_13403,N_13063);
nor U13580 (N_13580,N_13127,N_13113);
or U13581 (N_13581,N_13207,N_13172);
and U13582 (N_13582,N_13073,N_13057);
or U13583 (N_13583,N_13163,N_13228);
nor U13584 (N_13584,N_13333,N_13309);
xor U13585 (N_13585,N_13483,N_13436);
and U13586 (N_13586,N_13210,N_13191);
nor U13587 (N_13587,N_13439,N_13288);
xor U13588 (N_13588,N_13299,N_13070);
or U13589 (N_13589,N_13040,N_13402);
and U13590 (N_13590,N_13480,N_13250);
nor U13591 (N_13591,N_13176,N_13279);
nand U13592 (N_13592,N_13192,N_13416);
xor U13593 (N_13593,N_13050,N_13361);
and U13594 (N_13594,N_13359,N_13047);
xnor U13595 (N_13595,N_13114,N_13452);
xor U13596 (N_13596,N_13148,N_13116);
or U13597 (N_13597,N_13446,N_13096);
nor U13598 (N_13598,N_13281,N_13129);
xnor U13599 (N_13599,N_13198,N_13409);
nor U13600 (N_13600,N_13199,N_13217);
nand U13601 (N_13601,N_13488,N_13411);
xnor U13602 (N_13602,N_13425,N_13429);
or U13603 (N_13603,N_13135,N_13287);
xor U13604 (N_13604,N_13451,N_13252);
nor U13605 (N_13605,N_13365,N_13486);
xnor U13606 (N_13606,N_13044,N_13240);
xor U13607 (N_13607,N_13132,N_13092);
nor U13608 (N_13608,N_13374,N_13155);
and U13609 (N_13609,N_13251,N_13373);
or U13610 (N_13610,N_13459,N_13025);
xnor U13611 (N_13611,N_13464,N_13222);
nor U13612 (N_13612,N_13302,N_13115);
nand U13613 (N_13613,N_13391,N_13059);
and U13614 (N_13614,N_13190,N_13254);
xor U13615 (N_13615,N_13165,N_13133);
and U13616 (N_13616,N_13417,N_13476);
nor U13617 (N_13617,N_13106,N_13213);
or U13618 (N_13618,N_13068,N_13013);
xor U13619 (N_13619,N_13188,N_13315);
nand U13620 (N_13620,N_13455,N_13269);
xnor U13621 (N_13621,N_13322,N_13321);
and U13622 (N_13622,N_13401,N_13350);
or U13623 (N_13623,N_13318,N_13022);
or U13624 (N_13624,N_13066,N_13332);
and U13625 (N_13625,N_13327,N_13437);
and U13626 (N_13626,N_13062,N_13238);
xor U13627 (N_13627,N_13060,N_13084);
or U13628 (N_13628,N_13110,N_13038);
or U13629 (N_13629,N_13368,N_13194);
nand U13630 (N_13630,N_13450,N_13026);
or U13631 (N_13631,N_13447,N_13495);
and U13632 (N_13632,N_13015,N_13381);
nand U13633 (N_13633,N_13442,N_13219);
or U13634 (N_13634,N_13477,N_13197);
xor U13635 (N_13635,N_13454,N_13089);
nand U13636 (N_13636,N_13189,N_13426);
and U13637 (N_13637,N_13339,N_13473);
and U13638 (N_13638,N_13306,N_13033);
nand U13639 (N_13639,N_13467,N_13103);
nor U13640 (N_13640,N_13085,N_13474);
and U13641 (N_13641,N_13305,N_13045);
nor U13642 (N_13642,N_13428,N_13407);
xor U13643 (N_13643,N_13336,N_13487);
nor U13644 (N_13644,N_13311,N_13000);
xnor U13645 (N_13645,N_13168,N_13120);
nor U13646 (N_13646,N_13256,N_13264);
and U13647 (N_13647,N_13364,N_13058);
nor U13648 (N_13648,N_13118,N_13420);
and U13649 (N_13649,N_13278,N_13180);
nand U13650 (N_13650,N_13221,N_13161);
nand U13651 (N_13651,N_13048,N_13121);
nor U13652 (N_13652,N_13170,N_13095);
and U13653 (N_13653,N_13294,N_13093);
nand U13654 (N_13654,N_13146,N_13021);
nor U13655 (N_13655,N_13124,N_13253);
nand U13656 (N_13656,N_13471,N_13494);
or U13657 (N_13657,N_13375,N_13144);
xnor U13658 (N_13658,N_13216,N_13140);
nor U13659 (N_13659,N_13415,N_13147);
or U13660 (N_13660,N_13126,N_13080);
nand U13661 (N_13661,N_13329,N_13314);
and U13662 (N_13662,N_13139,N_13304);
xor U13663 (N_13663,N_13388,N_13366);
xnor U13664 (N_13664,N_13182,N_13234);
nand U13665 (N_13665,N_13461,N_13432);
xnor U13666 (N_13666,N_13303,N_13458);
xnor U13667 (N_13667,N_13443,N_13069);
xnor U13668 (N_13668,N_13111,N_13112);
xnor U13669 (N_13669,N_13201,N_13492);
nor U13670 (N_13670,N_13227,N_13064);
or U13671 (N_13671,N_13355,N_13352);
nor U13672 (N_13672,N_13438,N_13422);
and U13673 (N_13673,N_13435,N_13406);
xor U13674 (N_13674,N_13061,N_13017);
xor U13675 (N_13675,N_13006,N_13335);
or U13676 (N_13676,N_13326,N_13259);
or U13677 (N_13677,N_13289,N_13260);
xor U13678 (N_13678,N_13083,N_13145);
nor U13679 (N_13679,N_13310,N_13184);
nand U13680 (N_13680,N_13382,N_13075);
nor U13681 (N_13681,N_13024,N_13430);
nand U13682 (N_13682,N_13358,N_13123);
and U13683 (N_13683,N_13338,N_13346);
or U13684 (N_13684,N_13394,N_13396);
xor U13685 (N_13685,N_13389,N_13186);
or U13686 (N_13686,N_13007,N_13345);
nand U13687 (N_13687,N_13107,N_13481);
nor U13688 (N_13688,N_13449,N_13153);
xnor U13689 (N_13689,N_13325,N_13392);
xor U13690 (N_13690,N_13255,N_13283);
nand U13691 (N_13691,N_13209,N_13297);
and U13692 (N_13692,N_13109,N_13427);
or U13693 (N_13693,N_13342,N_13285);
or U13694 (N_13694,N_13215,N_13431);
nor U13695 (N_13695,N_13334,N_13351);
nor U13696 (N_13696,N_13414,N_13067);
or U13697 (N_13697,N_13091,N_13036);
or U13698 (N_13698,N_13317,N_13018);
xnor U13699 (N_13699,N_13003,N_13475);
and U13700 (N_13700,N_13413,N_13323);
xnor U13701 (N_13701,N_13377,N_13005);
xor U13702 (N_13702,N_13041,N_13131);
and U13703 (N_13703,N_13263,N_13243);
or U13704 (N_13704,N_13400,N_13324);
xnor U13705 (N_13705,N_13187,N_13456);
xor U13706 (N_13706,N_13125,N_13357);
and U13707 (N_13707,N_13393,N_13499);
nand U13708 (N_13708,N_13312,N_13497);
xor U13709 (N_13709,N_13233,N_13012);
nand U13710 (N_13710,N_13466,N_13496);
nor U13711 (N_13711,N_13246,N_13472);
xor U13712 (N_13712,N_13079,N_13100);
and U13713 (N_13713,N_13099,N_13042);
or U13714 (N_13714,N_13030,N_13225);
or U13715 (N_13715,N_13296,N_13370);
and U13716 (N_13716,N_13202,N_13348);
nand U13717 (N_13717,N_13101,N_13074);
nand U13718 (N_13718,N_13004,N_13223);
nand U13719 (N_13719,N_13049,N_13239);
nand U13720 (N_13720,N_13363,N_13027);
xor U13721 (N_13721,N_13460,N_13214);
nor U13722 (N_13722,N_13195,N_13218);
or U13723 (N_13723,N_13046,N_13362);
nor U13724 (N_13724,N_13249,N_13293);
and U13725 (N_13725,N_13276,N_13300);
or U13726 (N_13726,N_13286,N_13119);
xor U13727 (N_13727,N_13156,N_13130);
or U13728 (N_13728,N_13034,N_13395);
nand U13729 (N_13729,N_13086,N_13037);
nor U13730 (N_13730,N_13433,N_13337);
xor U13731 (N_13731,N_13235,N_13271);
nand U13732 (N_13732,N_13478,N_13019);
nand U13733 (N_13733,N_13236,N_13457);
nor U13734 (N_13734,N_13054,N_13383);
nand U13735 (N_13735,N_13211,N_13270);
nor U13736 (N_13736,N_13028,N_13340);
nor U13737 (N_13737,N_13149,N_13162);
xnor U13738 (N_13738,N_13128,N_13016);
nor U13739 (N_13739,N_13020,N_13349);
and U13740 (N_13740,N_13043,N_13014);
or U13741 (N_13741,N_13290,N_13479);
or U13742 (N_13742,N_13241,N_13230);
and U13743 (N_13743,N_13268,N_13053);
nor U13744 (N_13744,N_13200,N_13356);
nand U13745 (N_13745,N_13376,N_13412);
and U13746 (N_13746,N_13008,N_13397);
xnor U13747 (N_13747,N_13245,N_13029);
nor U13748 (N_13748,N_13248,N_13203);
or U13749 (N_13749,N_13274,N_13493);
nand U13750 (N_13750,N_13451,N_13392);
nor U13751 (N_13751,N_13268,N_13486);
and U13752 (N_13752,N_13434,N_13231);
xnor U13753 (N_13753,N_13033,N_13261);
and U13754 (N_13754,N_13164,N_13007);
nand U13755 (N_13755,N_13391,N_13226);
nand U13756 (N_13756,N_13267,N_13217);
nor U13757 (N_13757,N_13317,N_13132);
nor U13758 (N_13758,N_13166,N_13029);
xnor U13759 (N_13759,N_13054,N_13109);
or U13760 (N_13760,N_13197,N_13003);
or U13761 (N_13761,N_13272,N_13422);
nor U13762 (N_13762,N_13388,N_13275);
nor U13763 (N_13763,N_13357,N_13304);
nor U13764 (N_13764,N_13365,N_13334);
nand U13765 (N_13765,N_13418,N_13446);
nor U13766 (N_13766,N_13134,N_13205);
nor U13767 (N_13767,N_13016,N_13415);
or U13768 (N_13768,N_13171,N_13422);
nand U13769 (N_13769,N_13059,N_13214);
or U13770 (N_13770,N_13021,N_13462);
or U13771 (N_13771,N_13423,N_13325);
xor U13772 (N_13772,N_13434,N_13378);
and U13773 (N_13773,N_13180,N_13376);
nand U13774 (N_13774,N_13254,N_13238);
nor U13775 (N_13775,N_13261,N_13377);
or U13776 (N_13776,N_13077,N_13439);
nand U13777 (N_13777,N_13247,N_13348);
nand U13778 (N_13778,N_13328,N_13447);
or U13779 (N_13779,N_13438,N_13321);
nand U13780 (N_13780,N_13443,N_13093);
and U13781 (N_13781,N_13139,N_13391);
and U13782 (N_13782,N_13426,N_13028);
and U13783 (N_13783,N_13331,N_13493);
xor U13784 (N_13784,N_13379,N_13439);
nand U13785 (N_13785,N_13322,N_13105);
or U13786 (N_13786,N_13089,N_13130);
or U13787 (N_13787,N_13434,N_13355);
xor U13788 (N_13788,N_13025,N_13036);
and U13789 (N_13789,N_13012,N_13413);
or U13790 (N_13790,N_13374,N_13087);
nand U13791 (N_13791,N_13475,N_13196);
nor U13792 (N_13792,N_13434,N_13069);
and U13793 (N_13793,N_13489,N_13438);
and U13794 (N_13794,N_13361,N_13290);
or U13795 (N_13795,N_13049,N_13399);
or U13796 (N_13796,N_13042,N_13058);
or U13797 (N_13797,N_13106,N_13055);
xor U13798 (N_13798,N_13042,N_13426);
and U13799 (N_13799,N_13042,N_13087);
nor U13800 (N_13800,N_13486,N_13140);
and U13801 (N_13801,N_13006,N_13005);
or U13802 (N_13802,N_13288,N_13066);
xnor U13803 (N_13803,N_13258,N_13340);
xnor U13804 (N_13804,N_13137,N_13315);
xnor U13805 (N_13805,N_13091,N_13155);
nor U13806 (N_13806,N_13142,N_13237);
nor U13807 (N_13807,N_13352,N_13264);
and U13808 (N_13808,N_13354,N_13311);
or U13809 (N_13809,N_13209,N_13138);
and U13810 (N_13810,N_13088,N_13121);
and U13811 (N_13811,N_13190,N_13066);
or U13812 (N_13812,N_13107,N_13405);
nand U13813 (N_13813,N_13281,N_13437);
xor U13814 (N_13814,N_13031,N_13390);
xnor U13815 (N_13815,N_13283,N_13371);
xor U13816 (N_13816,N_13308,N_13408);
or U13817 (N_13817,N_13142,N_13020);
nand U13818 (N_13818,N_13324,N_13062);
nor U13819 (N_13819,N_13347,N_13453);
xnor U13820 (N_13820,N_13289,N_13241);
nor U13821 (N_13821,N_13000,N_13413);
nor U13822 (N_13822,N_13417,N_13006);
nor U13823 (N_13823,N_13134,N_13190);
or U13824 (N_13824,N_13218,N_13169);
and U13825 (N_13825,N_13116,N_13440);
nand U13826 (N_13826,N_13191,N_13456);
nand U13827 (N_13827,N_13061,N_13320);
nor U13828 (N_13828,N_13322,N_13316);
or U13829 (N_13829,N_13393,N_13249);
nor U13830 (N_13830,N_13060,N_13438);
nor U13831 (N_13831,N_13113,N_13214);
nand U13832 (N_13832,N_13228,N_13447);
xnor U13833 (N_13833,N_13043,N_13030);
and U13834 (N_13834,N_13465,N_13289);
nor U13835 (N_13835,N_13296,N_13405);
nand U13836 (N_13836,N_13495,N_13443);
or U13837 (N_13837,N_13027,N_13245);
nand U13838 (N_13838,N_13337,N_13274);
nand U13839 (N_13839,N_13229,N_13111);
xor U13840 (N_13840,N_13246,N_13135);
or U13841 (N_13841,N_13309,N_13118);
xnor U13842 (N_13842,N_13346,N_13175);
and U13843 (N_13843,N_13397,N_13175);
xor U13844 (N_13844,N_13129,N_13371);
nand U13845 (N_13845,N_13241,N_13324);
and U13846 (N_13846,N_13354,N_13015);
nor U13847 (N_13847,N_13014,N_13311);
xnor U13848 (N_13848,N_13204,N_13209);
xnor U13849 (N_13849,N_13263,N_13269);
or U13850 (N_13850,N_13397,N_13326);
or U13851 (N_13851,N_13176,N_13207);
nand U13852 (N_13852,N_13266,N_13059);
or U13853 (N_13853,N_13223,N_13039);
or U13854 (N_13854,N_13287,N_13022);
and U13855 (N_13855,N_13472,N_13273);
or U13856 (N_13856,N_13296,N_13008);
nand U13857 (N_13857,N_13390,N_13407);
or U13858 (N_13858,N_13221,N_13217);
xnor U13859 (N_13859,N_13232,N_13108);
nand U13860 (N_13860,N_13323,N_13370);
xnor U13861 (N_13861,N_13193,N_13139);
nand U13862 (N_13862,N_13464,N_13382);
or U13863 (N_13863,N_13316,N_13352);
xnor U13864 (N_13864,N_13028,N_13146);
nand U13865 (N_13865,N_13306,N_13400);
nand U13866 (N_13866,N_13412,N_13453);
and U13867 (N_13867,N_13363,N_13107);
xnor U13868 (N_13868,N_13290,N_13187);
or U13869 (N_13869,N_13358,N_13201);
and U13870 (N_13870,N_13229,N_13171);
nand U13871 (N_13871,N_13326,N_13291);
xor U13872 (N_13872,N_13427,N_13432);
xor U13873 (N_13873,N_13416,N_13311);
and U13874 (N_13874,N_13403,N_13473);
xor U13875 (N_13875,N_13466,N_13040);
nand U13876 (N_13876,N_13285,N_13132);
xor U13877 (N_13877,N_13097,N_13167);
xnor U13878 (N_13878,N_13217,N_13315);
nand U13879 (N_13879,N_13209,N_13152);
and U13880 (N_13880,N_13317,N_13111);
nand U13881 (N_13881,N_13031,N_13350);
and U13882 (N_13882,N_13212,N_13319);
nor U13883 (N_13883,N_13420,N_13194);
xnor U13884 (N_13884,N_13040,N_13059);
xor U13885 (N_13885,N_13353,N_13478);
nor U13886 (N_13886,N_13185,N_13250);
nand U13887 (N_13887,N_13044,N_13239);
or U13888 (N_13888,N_13440,N_13251);
xor U13889 (N_13889,N_13317,N_13057);
xnor U13890 (N_13890,N_13198,N_13310);
and U13891 (N_13891,N_13437,N_13042);
xor U13892 (N_13892,N_13385,N_13238);
nand U13893 (N_13893,N_13144,N_13322);
xor U13894 (N_13894,N_13313,N_13427);
or U13895 (N_13895,N_13301,N_13039);
or U13896 (N_13896,N_13074,N_13332);
xor U13897 (N_13897,N_13245,N_13271);
nand U13898 (N_13898,N_13163,N_13277);
and U13899 (N_13899,N_13445,N_13127);
nor U13900 (N_13900,N_13040,N_13251);
xnor U13901 (N_13901,N_13412,N_13248);
nand U13902 (N_13902,N_13181,N_13038);
and U13903 (N_13903,N_13286,N_13239);
and U13904 (N_13904,N_13077,N_13464);
xnor U13905 (N_13905,N_13117,N_13193);
xnor U13906 (N_13906,N_13235,N_13068);
or U13907 (N_13907,N_13176,N_13400);
nor U13908 (N_13908,N_13186,N_13423);
nor U13909 (N_13909,N_13134,N_13457);
xor U13910 (N_13910,N_13013,N_13402);
or U13911 (N_13911,N_13472,N_13216);
nand U13912 (N_13912,N_13113,N_13242);
and U13913 (N_13913,N_13436,N_13454);
or U13914 (N_13914,N_13469,N_13481);
nor U13915 (N_13915,N_13051,N_13042);
nor U13916 (N_13916,N_13227,N_13099);
nand U13917 (N_13917,N_13264,N_13268);
or U13918 (N_13918,N_13354,N_13392);
nor U13919 (N_13919,N_13248,N_13311);
xnor U13920 (N_13920,N_13458,N_13052);
xor U13921 (N_13921,N_13430,N_13303);
xor U13922 (N_13922,N_13470,N_13314);
or U13923 (N_13923,N_13102,N_13465);
or U13924 (N_13924,N_13233,N_13045);
and U13925 (N_13925,N_13305,N_13231);
or U13926 (N_13926,N_13470,N_13051);
or U13927 (N_13927,N_13296,N_13423);
nand U13928 (N_13928,N_13067,N_13250);
and U13929 (N_13929,N_13134,N_13172);
and U13930 (N_13930,N_13148,N_13139);
nand U13931 (N_13931,N_13030,N_13211);
nor U13932 (N_13932,N_13452,N_13424);
and U13933 (N_13933,N_13281,N_13091);
nand U13934 (N_13934,N_13032,N_13025);
xnor U13935 (N_13935,N_13141,N_13142);
and U13936 (N_13936,N_13057,N_13123);
nor U13937 (N_13937,N_13396,N_13162);
or U13938 (N_13938,N_13405,N_13352);
nor U13939 (N_13939,N_13460,N_13189);
nand U13940 (N_13940,N_13121,N_13166);
xnor U13941 (N_13941,N_13110,N_13490);
or U13942 (N_13942,N_13213,N_13130);
nor U13943 (N_13943,N_13089,N_13084);
or U13944 (N_13944,N_13360,N_13269);
nand U13945 (N_13945,N_13335,N_13220);
xnor U13946 (N_13946,N_13211,N_13480);
nor U13947 (N_13947,N_13074,N_13182);
xnor U13948 (N_13948,N_13317,N_13212);
or U13949 (N_13949,N_13242,N_13277);
nor U13950 (N_13950,N_13410,N_13161);
nand U13951 (N_13951,N_13127,N_13079);
nand U13952 (N_13952,N_13371,N_13018);
or U13953 (N_13953,N_13082,N_13349);
nand U13954 (N_13954,N_13270,N_13412);
nor U13955 (N_13955,N_13241,N_13134);
and U13956 (N_13956,N_13392,N_13334);
nor U13957 (N_13957,N_13115,N_13243);
nand U13958 (N_13958,N_13150,N_13220);
or U13959 (N_13959,N_13223,N_13204);
and U13960 (N_13960,N_13192,N_13267);
or U13961 (N_13961,N_13285,N_13176);
or U13962 (N_13962,N_13353,N_13407);
nand U13963 (N_13963,N_13206,N_13085);
xnor U13964 (N_13964,N_13087,N_13181);
nor U13965 (N_13965,N_13081,N_13175);
or U13966 (N_13966,N_13300,N_13234);
nor U13967 (N_13967,N_13456,N_13467);
nor U13968 (N_13968,N_13248,N_13340);
nor U13969 (N_13969,N_13171,N_13313);
or U13970 (N_13970,N_13006,N_13032);
nor U13971 (N_13971,N_13286,N_13406);
xor U13972 (N_13972,N_13435,N_13110);
nand U13973 (N_13973,N_13258,N_13480);
or U13974 (N_13974,N_13245,N_13329);
nor U13975 (N_13975,N_13008,N_13321);
or U13976 (N_13976,N_13004,N_13447);
and U13977 (N_13977,N_13260,N_13084);
xnor U13978 (N_13978,N_13257,N_13014);
or U13979 (N_13979,N_13120,N_13286);
or U13980 (N_13980,N_13315,N_13293);
nand U13981 (N_13981,N_13340,N_13042);
xor U13982 (N_13982,N_13167,N_13054);
or U13983 (N_13983,N_13120,N_13250);
xor U13984 (N_13984,N_13291,N_13154);
nor U13985 (N_13985,N_13127,N_13095);
and U13986 (N_13986,N_13370,N_13343);
nand U13987 (N_13987,N_13169,N_13241);
nor U13988 (N_13988,N_13420,N_13048);
nor U13989 (N_13989,N_13306,N_13117);
xor U13990 (N_13990,N_13068,N_13114);
nor U13991 (N_13991,N_13113,N_13401);
nand U13992 (N_13992,N_13084,N_13360);
nor U13993 (N_13993,N_13132,N_13416);
xor U13994 (N_13994,N_13424,N_13112);
nor U13995 (N_13995,N_13379,N_13266);
xor U13996 (N_13996,N_13326,N_13447);
nor U13997 (N_13997,N_13419,N_13250);
xor U13998 (N_13998,N_13493,N_13097);
nand U13999 (N_13999,N_13473,N_13471);
xnor U14000 (N_14000,N_13917,N_13519);
xnor U14001 (N_14001,N_13801,N_13603);
and U14002 (N_14002,N_13778,N_13672);
nor U14003 (N_14003,N_13517,N_13851);
nand U14004 (N_14004,N_13654,N_13975);
xor U14005 (N_14005,N_13502,N_13749);
nor U14006 (N_14006,N_13667,N_13582);
nor U14007 (N_14007,N_13592,N_13837);
and U14008 (N_14008,N_13982,N_13561);
nand U14009 (N_14009,N_13538,N_13656);
and U14010 (N_14010,N_13703,N_13790);
nand U14011 (N_14011,N_13725,N_13512);
xnor U14012 (N_14012,N_13732,N_13552);
nor U14013 (N_14013,N_13729,N_13984);
and U14014 (N_14014,N_13613,N_13739);
nand U14015 (N_14015,N_13659,N_13840);
and U14016 (N_14016,N_13650,N_13946);
nor U14017 (N_14017,N_13506,N_13830);
nor U14018 (N_14018,N_13571,N_13641);
xor U14019 (N_14019,N_13677,N_13660);
xor U14020 (N_14020,N_13836,N_13541);
xnor U14021 (N_14021,N_13652,N_13748);
nand U14022 (N_14022,N_13935,N_13762);
nor U14023 (N_14023,N_13589,N_13817);
and U14024 (N_14024,N_13691,N_13776);
nand U14025 (N_14025,N_13990,N_13981);
xnor U14026 (N_14026,N_13915,N_13905);
or U14027 (N_14027,N_13598,N_13833);
nor U14028 (N_14028,N_13764,N_13713);
or U14029 (N_14029,N_13875,N_13528);
and U14030 (N_14030,N_13688,N_13838);
and U14031 (N_14031,N_13818,N_13923);
nand U14032 (N_14032,N_13756,N_13735);
nand U14033 (N_14033,N_13874,N_13721);
and U14034 (N_14034,N_13550,N_13900);
xor U14035 (N_14035,N_13763,N_13809);
nand U14036 (N_14036,N_13610,N_13546);
or U14037 (N_14037,N_13842,N_13861);
or U14038 (N_14038,N_13712,N_13924);
xor U14039 (N_14039,N_13886,N_13526);
nor U14040 (N_14040,N_13942,N_13616);
nand U14041 (N_14041,N_13683,N_13815);
nor U14042 (N_14042,N_13687,N_13821);
xnor U14043 (N_14043,N_13751,N_13773);
or U14044 (N_14044,N_13952,N_13642);
and U14045 (N_14045,N_13509,N_13588);
or U14046 (N_14046,N_13894,N_13774);
and U14047 (N_14047,N_13702,N_13564);
and U14048 (N_14048,N_13810,N_13898);
or U14049 (N_14049,N_13947,N_13661);
and U14050 (N_14050,N_13908,N_13991);
xnor U14051 (N_14051,N_13829,N_13822);
and U14052 (N_14052,N_13633,N_13951);
nand U14053 (N_14053,N_13843,N_13505);
or U14054 (N_14054,N_13602,N_13782);
nor U14055 (N_14055,N_13681,N_13578);
or U14056 (N_14056,N_13727,N_13568);
xnor U14057 (N_14057,N_13772,N_13783);
or U14058 (N_14058,N_13530,N_13812);
or U14059 (N_14059,N_13724,N_13954);
or U14060 (N_14060,N_13686,N_13963);
xor U14061 (N_14061,N_13577,N_13554);
nor U14062 (N_14062,N_13537,N_13918);
and U14063 (N_14063,N_13536,N_13959);
xor U14064 (N_14064,N_13555,N_13593);
nor U14065 (N_14065,N_13948,N_13586);
xor U14066 (N_14066,N_13730,N_13710);
xor U14067 (N_14067,N_13708,N_13580);
or U14068 (N_14068,N_13978,N_13707);
or U14069 (N_14069,N_13929,N_13912);
nand U14070 (N_14070,N_13844,N_13955);
nor U14071 (N_14071,N_13883,N_13698);
nor U14072 (N_14072,N_13863,N_13508);
or U14073 (N_14073,N_13716,N_13734);
and U14074 (N_14074,N_13547,N_13655);
nand U14075 (N_14075,N_13811,N_13871);
or U14076 (N_14076,N_13781,N_13969);
nand U14077 (N_14077,N_13722,N_13998);
xnor U14078 (N_14078,N_13945,N_13824);
and U14079 (N_14079,N_13662,N_13880);
nor U14080 (N_14080,N_13997,N_13666);
nand U14081 (N_14081,N_13866,N_13758);
or U14082 (N_14082,N_13849,N_13922);
nand U14083 (N_14083,N_13852,N_13609);
xnor U14084 (N_14084,N_13726,N_13839);
nor U14085 (N_14085,N_13545,N_13941);
or U14086 (N_14086,N_13621,N_13630);
or U14087 (N_14087,N_13738,N_13570);
nand U14088 (N_14088,N_13897,N_13983);
nor U14089 (N_14089,N_13544,N_13966);
xnor U14090 (N_14090,N_13827,N_13747);
nor U14091 (N_14091,N_13927,N_13717);
nand U14092 (N_14092,N_13961,N_13607);
and U14093 (N_14093,N_13744,N_13513);
nand U14094 (N_14094,N_13585,N_13524);
nor U14095 (N_14095,N_13514,N_13556);
nor U14096 (N_14096,N_13615,N_13757);
or U14097 (N_14097,N_13620,N_13792);
or U14098 (N_14098,N_13535,N_13803);
nand U14099 (N_14099,N_13916,N_13742);
nand U14100 (N_14100,N_13532,N_13933);
and U14101 (N_14101,N_13770,N_13551);
and U14102 (N_14102,N_13953,N_13521);
and U14103 (N_14103,N_13648,N_13807);
nor U14104 (N_14104,N_13902,N_13813);
or U14105 (N_14105,N_13657,N_13899);
and U14106 (N_14106,N_13701,N_13956);
and U14107 (N_14107,N_13507,N_13599);
xor U14108 (N_14108,N_13643,N_13796);
xor U14109 (N_14109,N_13765,N_13558);
xnor U14110 (N_14110,N_13925,N_13693);
or U14111 (N_14111,N_13706,N_13516);
nand U14112 (N_14112,N_13814,N_13549);
nand U14113 (N_14113,N_13854,N_13733);
and U14114 (N_14114,N_13569,N_13960);
and U14115 (N_14115,N_13575,N_13576);
nor U14116 (N_14116,N_13768,N_13943);
and U14117 (N_14117,N_13583,N_13913);
xnor U14118 (N_14118,N_13523,N_13649);
xnor U14119 (N_14119,N_13696,N_13623);
xnor U14120 (N_14120,N_13614,N_13759);
xnor U14121 (N_14121,N_13591,N_13850);
or U14122 (N_14122,N_13872,N_13936);
nand U14123 (N_14123,N_13937,N_13760);
nand U14124 (N_14124,N_13560,N_13685);
and U14125 (N_14125,N_13627,N_13789);
and U14126 (N_14126,N_13754,N_13786);
and U14127 (N_14127,N_13709,N_13835);
and U14128 (N_14128,N_13619,N_13563);
or U14129 (N_14129,N_13976,N_13846);
or U14130 (N_14130,N_13604,N_13767);
or U14131 (N_14131,N_13791,N_13825);
nand U14132 (N_14132,N_13992,N_13995);
nand U14133 (N_14133,N_13797,N_13629);
nand U14134 (N_14134,N_13664,N_13562);
or U14135 (N_14135,N_13973,N_13675);
nor U14136 (N_14136,N_13540,N_13679);
and U14137 (N_14137,N_13775,N_13845);
nand U14138 (N_14138,N_13719,N_13950);
or U14139 (N_14139,N_13893,N_13625);
nand U14140 (N_14140,N_13788,N_13670);
and U14141 (N_14141,N_13510,N_13635);
or U14142 (N_14142,N_13622,N_13868);
nand U14143 (N_14143,N_13731,N_13938);
and U14144 (N_14144,N_13596,N_13986);
and U14145 (N_14145,N_13503,N_13944);
xor U14146 (N_14146,N_13853,N_13873);
and U14147 (N_14147,N_13920,N_13699);
nor U14148 (N_14148,N_13634,N_13834);
and U14149 (N_14149,N_13971,N_13798);
nor U14150 (N_14150,N_13640,N_13799);
xnor U14151 (N_14151,N_13939,N_13780);
nor U14152 (N_14152,N_13674,N_13618);
or U14153 (N_14153,N_13889,N_13888);
or U14154 (N_14154,N_13881,N_13628);
xor U14155 (N_14155,N_13841,N_13645);
or U14156 (N_14156,N_13884,N_13753);
and U14157 (N_14157,N_13958,N_13794);
nand U14158 (N_14158,N_13785,N_13755);
nor U14159 (N_14159,N_13745,N_13793);
or U14160 (N_14160,N_13860,N_13877);
nor U14161 (N_14161,N_13636,N_13606);
nor U14162 (N_14162,N_13970,N_13581);
or U14163 (N_14163,N_13736,N_13631);
nand U14164 (N_14164,N_13740,N_13808);
nor U14165 (N_14165,N_13692,N_13921);
or U14166 (N_14166,N_13584,N_13644);
nand U14167 (N_14167,N_13892,N_13638);
nand U14168 (N_14168,N_13895,N_13587);
or U14169 (N_14169,N_13548,N_13689);
or U14170 (N_14170,N_13542,N_13879);
and U14171 (N_14171,N_13590,N_13704);
nor U14172 (N_14172,N_13940,N_13934);
and U14173 (N_14173,N_13847,N_13856);
or U14174 (N_14174,N_13676,N_13962);
nor U14175 (N_14175,N_13859,N_13910);
xnor U14176 (N_14176,N_13671,N_13529);
xor U14177 (N_14177,N_13926,N_13919);
and U14178 (N_14178,N_13994,N_13974);
xor U14179 (N_14179,N_13891,N_13769);
nor U14180 (N_14180,N_13565,N_13700);
and U14181 (N_14181,N_13601,N_13646);
nand U14182 (N_14182,N_13996,N_13826);
nor U14183 (N_14183,N_13848,N_13771);
or U14184 (N_14184,N_13515,N_13567);
or U14185 (N_14185,N_13608,N_13870);
nand U14186 (N_14186,N_13857,N_13624);
nor U14187 (N_14187,N_13539,N_13617);
or U14188 (N_14188,N_13658,N_13557);
and U14189 (N_14189,N_13743,N_13989);
or U14190 (N_14190,N_13795,N_13680);
and U14191 (N_14191,N_13858,N_13805);
nand U14192 (N_14192,N_13504,N_13965);
nor U14193 (N_14193,N_13885,N_13890);
nor U14194 (N_14194,N_13665,N_13720);
and U14195 (N_14195,N_13766,N_13876);
nor U14196 (N_14196,N_13887,N_13597);
and U14197 (N_14197,N_13728,N_13931);
nor U14198 (N_14198,N_13867,N_13914);
nor U14199 (N_14199,N_13626,N_13862);
or U14200 (N_14200,N_13779,N_13684);
or U14201 (N_14201,N_13579,N_13566);
nand U14202 (N_14202,N_13695,N_13559);
or U14203 (N_14203,N_13896,N_13500);
and U14204 (N_14204,N_13543,N_13741);
nand U14205 (N_14205,N_13800,N_13977);
xnor U14206 (N_14206,N_13611,N_13957);
xor U14207 (N_14207,N_13784,N_13705);
nor U14208 (N_14208,N_13632,N_13999);
xor U14209 (N_14209,N_13669,N_13663);
and U14210 (N_14210,N_13928,N_13682);
nor U14211 (N_14211,N_13527,N_13828);
or U14212 (N_14212,N_13715,N_13967);
xor U14213 (N_14213,N_13816,N_13534);
or U14214 (N_14214,N_13968,N_13746);
and U14215 (N_14215,N_13819,N_13711);
nand U14216 (N_14216,N_13651,N_13980);
xor U14217 (N_14217,N_13600,N_13949);
and U14218 (N_14218,N_13737,N_13653);
or U14219 (N_14219,N_13882,N_13972);
nand U14220 (N_14220,N_13911,N_13697);
nor U14221 (N_14221,N_13869,N_13639);
or U14222 (N_14222,N_13574,N_13752);
xnor U14223 (N_14223,N_13804,N_13907);
nand U14224 (N_14224,N_13694,N_13932);
nand U14225 (N_14225,N_13522,N_13802);
and U14226 (N_14226,N_13668,N_13906);
or U14227 (N_14227,N_13823,N_13964);
and U14228 (N_14228,N_13714,N_13988);
nand U14229 (N_14229,N_13903,N_13864);
or U14230 (N_14230,N_13637,N_13806);
or U14231 (N_14231,N_13750,N_13525);
nand U14232 (N_14232,N_13832,N_13531);
or U14233 (N_14233,N_13511,N_13985);
or U14234 (N_14234,N_13930,N_13612);
and U14235 (N_14235,N_13993,N_13787);
and U14236 (N_14236,N_13987,N_13777);
or U14237 (N_14237,N_13855,N_13979);
nor U14238 (N_14238,N_13572,N_13878);
and U14239 (N_14239,N_13723,N_13909);
and U14240 (N_14240,N_13718,N_13901);
nor U14241 (N_14241,N_13533,N_13553);
nand U14242 (N_14242,N_13820,N_13673);
nor U14243 (N_14243,N_13520,N_13690);
nand U14244 (N_14244,N_13594,N_13865);
or U14245 (N_14245,N_13573,N_13605);
or U14246 (N_14246,N_13761,N_13595);
xnor U14247 (N_14247,N_13678,N_13831);
xnor U14248 (N_14248,N_13647,N_13904);
xor U14249 (N_14249,N_13518,N_13501);
nand U14250 (N_14250,N_13615,N_13567);
nor U14251 (N_14251,N_13751,N_13768);
xnor U14252 (N_14252,N_13833,N_13712);
nand U14253 (N_14253,N_13635,N_13879);
or U14254 (N_14254,N_13515,N_13676);
and U14255 (N_14255,N_13752,N_13850);
nand U14256 (N_14256,N_13534,N_13854);
nor U14257 (N_14257,N_13933,N_13617);
nor U14258 (N_14258,N_13616,N_13813);
xor U14259 (N_14259,N_13930,N_13771);
and U14260 (N_14260,N_13724,N_13512);
nand U14261 (N_14261,N_13535,N_13545);
or U14262 (N_14262,N_13562,N_13741);
nand U14263 (N_14263,N_13748,N_13591);
nand U14264 (N_14264,N_13538,N_13757);
or U14265 (N_14265,N_13876,N_13930);
or U14266 (N_14266,N_13521,N_13861);
and U14267 (N_14267,N_13714,N_13890);
xor U14268 (N_14268,N_13751,N_13966);
xor U14269 (N_14269,N_13941,N_13762);
or U14270 (N_14270,N_13739,N_13720);
and U14271 (N_14271,N_13813,N_13793);
nand U14272 (N_14272,N_13913,N_13644);
or U14273 (N_14273,N_13648,N_13736);
nand U14274 (N_14274,N_13617,N_13681);
nand U14275 (N_14275,N_13752,N_13947);
nor U14276 (N_14276,N_13585,N_13851);
or U14277 (N_14277,N_13763,N_13560);
nand U14278 (N_14278,N_13551,N_13686);
nand U14279 (N_14279,N_13779,N_13832);
nor U14280 (N_14280,N_13722,N_13857);
or U14281 (N_14281,N_13991,N_13517);
nand U14282 (N_14282,N_13513,N_13882);
or U14283 (N_14283,N_13649,N_13947);
or U14284 (N_14284,N_13987,N_13945);
xnor U14285 (N_14285,N_13655,N_13608);
nand U14286 (N_14286,N_13951,N_13611);
and U14287 (N_14287,N_13966,N_13836);
nor U14288 (N_14288,N_13919,N_13869);
or U14289 (N_14289,N_13998,N_13822);
nor U14290 (N_14290,N_13598,N_13884);
nand U14291 (N_14291,N_13904,N_13643);
nand U14292 (N_14292,N_13905,N_13587);
nand U14293 (N_14293,N_13842,N_13512);
nor U14294 (N_14294,N_13640,N_13669);
xor U14295 (N_14295,N_13747,N_13751);
nor U14296 (N_14296,N_13820,N_13816);
xor U14297 (N_14297,N_13544,N_13560);
nand U14298 (N_14298,N_13922,N_13968);
nor U14299 (N_14299,N_13765,N_13502);
and U14300 (N_14300,N_13964,N_13798);
and U14301 (N_14301,N_13808,N_13794);
xnor U14302 (N_14302,N_13672,N_13925);
nand U14303 (N_14303,N_13536,N_13629);
and U14304 (N_14304,N_13815,N_13505);
xnor U14305 (N_14305,N_13881,N_13675);
xnor U14306 (N_14306,N_13822,N_13893);
xnor U14307 (N_14307,N_13786,N_13829);
or U14308 (N_14308,N_13956,N_13549);
nor U14309 (N_14309,N_13721,N_13924);
nand U14310 (N_14310,N_13602,N_13677);
xnor U14311 (N_14311,N_13714,N_13987);
xor U14312 (N_14312,N_13631,N_13660);
or U14313 (N_14313,N_13817,N_13572);
or U14314 (N_14314,N_13757,N_13713);
xnor U14315 (N_14315,N_13615,N_13910);
nor U14316 (N_14316,N_13782,N_13690);
nor U14317 (N_14317,N_13691,N_13914);
and U14318 (N_14318,N_13658,N_13609);
xnor U14319 (N_14319,N_13844,N_13924);
and U14320 (N_14320,N_13956,N_13877);
and U14321 (N_14321,N_13665,N_13507);
nor U14322 (N_14322,N_13917,N_13935);
or U14323 (N_14323,N_13715,N_13869);
xor U14324 (N_14324,N_13945,N_13600);
or U14325 (N_14325,N_13518,N_13725);
nor U14326 (N_14326,N_13821,N_13901);
or U14327 (N_14327,N_13520,N_13667);
nand U14328 (N_14328,N_13908,N_13756);
nand U14329 (N_14329,N_13637,N_13841);
xor U14330 (N_14330,N_13991,N_13728);
nor U14331 (N_14331,N_13670,N_13615);
and U14332 (N_14332,N_13728,N_13663);
xnor U14333 (N_14333,N_13561,N_13609);
xor U14334 (N_14334,N_13722,N_13505);
or U14335 (N_14335,N_13684,N_13920);
and U14336 (N_14336,N_13880,N_13532);
nor U14337 (N_14337,N_13541,N_13546);
nand U14338 (N_14338,N_13707,N_13873);
nand U14339 (N_14339,N_13500,N_13876);
nor U14340 (N_14340,N_13666,N_13714);
and U14341 (N_14341,N_13698,N_13869);
nor U14342 (N_14342,N_13837,N_13856);
and U14343 (N_14343,N_13634,N_13703);
xnor U14344 (N_14344,N_13996,N_13619);
or U14345 (N_14345,N_13634,N_13610);
nand U14346 (N_14346,N_13635,N_13728);
and U14347 (N_14347,N_13708,N_13755);
nor U14348 (N_14348,N_13840,N_13747);
and U14349 (N_14349,N_13681,N_13814);
or U14350 (N_14350,N_13610,N_13760);
nor U14351 (N_14351,N_13733,N_13661);
and U14352 (N_14352,N_13669,N_13765);
nand U14353 (N_14353,N_13704,N_13901);
nor U14354 (N_14354,N_13646,N_13875);
or U14355 (N_14355,N_13942,N_13742);
and U14356 (N_14356,N_13980,N_13711);
and U14357 (N_14357,N_13701,N_13909);
nor U14358 (N_14358,N_13810,N_13550);
nand U14359 (N_14359,N_13969,N_13853);
nand U14360 (N_14360,N_13904,N_13857);
and U14361 (N_14361,N_13917,N_13905);
nand U14362 (N_14362,N_13600,N_13613);
nand U14363 (N_14363,N_13849,N_13696);
nor U14364 (N_14364,N_13810,N_13764);
and U14365 (N_14365,N_13756,N_13512);
nor U14366 (N_14366,N_13620,N_13681);
or U14367 (N_14367,N_13864,N_13542);
and U14368 (N_14368,N_13993,N_13894);
or U14369 (N_14369,N_13574,N_13786);
or U14370 (N_14370,N_13822,N_13512);
and U14371 (N_14371,N_13581,N_13953);
and U14372 (N_14372,N_13765,N_13605);
and U14373 (N_14373,N_13679,N_13779);
nor U14374 (N_14374,N_13898,N_13971);
and U14375 (N_14375,N_13739,N_13856);
xnor U14376 (N_14376,N_13502,N_13705);
and U14377 (N_14377,N_13811,N_13693);
nand U14378 (N_14378,N_13705,N_13657);
xnor U14379 (N_14379,N_13823,N_13572);
and U14380 (N_14380,N_13856,N_13636);
nor U14381 (N_14381,N_13730,N_13501);
or U14382 (N_14382,N_13996,N_13675);
nand U14383 (N_14383,N_13712,N_13837);
xnor U14384 (N_14384,N_13905,N_13652);
or U14385 (N_14385,N_13743,N_13617);
nand U14386 (N_14386,N_13527,N_13603);
nor U14387 (N_14387,N_13903,N_13933);
nand U14388 (N_14388,N_13958,N_13527);
nor U14389 (N_14389,N_13886,N_13586);
xnor U14390 (N_14390,N_13848,N_13551);
nor U14391 (N_14391,N_13912,N_13892);
or U14392 (N_14392,N_13710,N_13800);
nand U14393 (N_14393,N_13527,N_13763);
nor U14394 (N_14394,N_13704,N_13681);
nand U14395 (N_14395,N_13907,N_13969);
nand U14396 (N_14396,N_13809,N_13891);
or U14397 (N_14397,N_13927,N_13544);
nor U14398 (N_14398,N_13631,N_13536);
or U14399 (N_14399,N_13948,N_13501);
and U14400 (N_14400,N_13577,N_13842);
and U14401 (N_14401,N_13588,N_13679);
and U14402 (N_14402,N_13838,N_13858);
or U14403 (N_14403,N_13930,N_13759);
nor U14404 (N_14404,N_13821,N_13684);
and U14405 (N_14405,N_13646,N_13673);
xnor U14406 (N_14406,N_13864,N_13872);
or U14407 (N_14407,N_13999,N_13906);
and U14408 (N_14408,N_13520,N_13894);
or U14409 (N_14409,N_13570,N_13889);
or U14410 (N_14410,N_13832,N_13830);
nor U14411 (N_14411,N_13505,N_13750);
or U14412 (N_14412,N_13821,N_13903);
nand U14413 (N_14413,N_13554,N_13536);
nand U14414 (N_14414,N_13820,N_13857);
xor U14415 (N_14415,N_13875,N_13799);
nand U14416 (N_14416,N_13531,N_13876);
or U14417 (N_14417,N_13654,N_13789);
nor U14418 (N_14418,N_13909,N_13570);
nor U14419 (N_14419,N_13609,N_13902);
xor U14420 (N_14420,N_13670,N_13834);
nand U14421 (N_14421,N_13600,N_13751);
and U14422 (N_14422,N_13661,N_13970);
and U14423 (N_14423,N_13615,N_13516);
and U14424 (N_14424,N_13943,N_13715);
nor U14425 (N_14425,N_13759,N_13630);
nand U14426 (N_14426,N_13662,N_13633);
nor U14427 (N_14427,N_13899,N_13826);
xnor U14428 (N_14428,N_13807,N_13511);
nand U14429 (N_14429,N_13610,N_13680);
nor U14430 (N_14430,N_13820,N_13516);
xor U14431 (N_14431,N_13972,N_13716);
and U14432 (N_14432,N_13677,N_13859);
xor U14433 (N_14433,N_13737,N_13738);
nor U14434 (N_14434,N_13679,N_13947);
nand U14435 (N_14435,N_13550,N_13892);
nand U14436 (N_14436,N_13836,N_13814);
nor U14437 (N_14437,N_13616,N_13937);
nor U14438 (N_14438,N_13619,N_13690);
xor U14439 (N_14439,N_13907,N_13537);
xor U14440 (N_14440,N_13800,N_13534);
and U14441 (N_14441,N_13965,N_13744);
nor U14442 (N_14442,N_13728,N_13639);
xnor U14443 (N_14443,N_13851,N_13790);
nand U14444 (N_14444,N_13820,N_13950);
xnor U14445 (N_14445,N_13531,N_13899);
xnor U14446 (N_14446,N_13843,N_13652);
nor U14447 (N_14447,N_13919,N_13837);
and U14448 (N_14448,N_13918,N_13804);
or U14449 (N_14449,N_13974,N_13798);
xnor U14450 (N_14450,N_13720,N_13540);
and U14451 (N_14451,N_13908,N_13948);
nor U14452 (N_14452,N_13558,N_13582);
nand U14453 (N_14453,N_13610,N_13624);
and U14454 (N_14454,N_13586,N_13854);
xor U14455 (N_14455,N_13659,N_13928);
and U14456 (N_14456,N_13550,N_13672);
xor U14457 (N_14457,N_13762,N_13610);
nor U14458 (N_14458,N_13585,N_13691);
nand U14459 (N_14459,N_13608,N_13725);
xnor U14460 (N_14460,N_13799,N_13874);
xnor U14461 (N_14461,N_13869,N_13816);
and U14462 (N_14462,N_13574,N_13922);
nand U14463 (N_14463,N_13523,N_13610);
nand U14464 (N_14464,N_13825,N_13770);
and U14465 (N_14465,N_13955,N_13869);
nor U14466 (N_14466,N_13967,N_13677);
nand U14467 (N_14467,N_13796,N_13585);
nand U14468 (N_14468,N_13940,N_13747);
or U14469 (N_14469,N_13772,N_13538);
nor U14470 (N_14470,N_13947,N_13627);
xnor U14471 (N_14471,N_13563,N_13831);
nand U14472 (N_14472,N_13920,N_13845);
xor U14473 (N_14473,N_13571,N_13920);
nor U14474 (N_14474,N_13730,N_13665);
or U14475 (N_14475,N_13594,N_13673);
nand U14476 (N_14476,N_13709,N_13702);
nand U14477 (N_14477,N_13822,N_13556);
and U14478 (N_14478,N_13984,N_13946);
or U14479 (N_14479,N_13636,N_13989);
nand U14480 (N_14480,N_13503,N_13695);
nor U14481 (N_14481,N_13641,N_13627);
nor U14482 (N_14482,N_13710,N_13793);
xnor U14483 (N_14483,N_13642,N_13651);
nor U14484 (N_14484,N_13572,N_13687);
or U14485 (N_14485,N_13820,N_13880);
nor U14486 (N_14486,N_13628,N_13625);
or U14487 (N_14487,N_13575,N_13867);
nand U14488 (N_14488,N_13659,N_13614);
and U14489 (N_14489,N_13912,N_13516);
nor U14490 (N_14490,N_13616,N_13739);
and U14491 (N_14491,N_13767,N_13948);
and U14492 (N_14492,N_13558,N_13560);
nand U14493 (N_14493,N_13528,N_13971);
nand U14494 (N_14494,N_13962,N_13853);
nand U14495 (N_14495,N_13564,N_13897);
xnor U14496 (N_14496,N_13926,N_13970);
nand U14497 (N_14497,N_13862,N_13541);
or U14498 (N_14498,N_13693,N_13876);
or U14499 (N_14499,N_13646,N_13869);
xnor U14500 (N_14500,N_14093,N_14181);
or U14501 (N_14501,N_14041,N_14052);
and U14502 (N_14502,N_14103,N_14154);
or U14503 (N_14503,N_14334,N_14010);
nor U14504 (N_14504,N_14194,N_14184);
and U14505 (N_14505,N_14222,N_14060);
and U14506 (N_14506,N_14243,N_14421);
and U14507 (N_14507,N_14162,N_14392);
xnor U14508 (N_14508,N_14206,N_14038);
or U14509 (N_14509,N_14488,N_14188);
nand U14510 (N_14510,N_14440,N_14067);
xnor U14511 (N_14511,N_14442,N_14346);
nand U14512 (N_14512,N_14470,N_14394);
nand U14513 (N_14513,N_14236,N_14028);
xnor U14514 (N_14514,N_14017,N_14201);
nor U14515 (N_14515,N_14172,N_14451);
nor U14516 (N_14516,N_14220,N_14102);
nor U14517 (N_14517,N_14111,N_14251);
xor U14518 (N_14518,N_14468,N_14433);
or U14519 (N_14519,N_14375,N_14146);
and U14520 (N_14520,N_14416,N_14225);
xnor U14521 (N_14521,N_14163,N_14305);
nor U14522 (N_14522,N_14139,N_14256);
nand U14523 (N_14523,N_14372,N_14486);
nand U14524 (N_14524,N_14192,N_14036);
nand U14525 (N_14525,N_14040,N_14325);
or U14526 (N_14526,N_14149,N_14310);
nand U14527 (N_14527,N_14293,N_14495);
and U14528 (N_14528,N_14483,N_14447);
nor U14529 (N_14529,N_14315,N_14368);
xnor U14530 (N_14530,N_14189,N_14354);
xor U14531 (N_14531,N_14330,N_14059);
nand U14532 (N_14532,N_14498,N_14101);
nor U14533 (N_14533,N_14492,N_14107);
and U14534 (N_14534,N_14185,N_14013);
and U14535 (N_14535,N_14113,N_14079);
nor U14536 (N_14536,N_14232,N_14365);
nor U14537 (N_14537,N_14098,N_14007);
xnor U14538 (N_14538,N_14340,N_14289);
and U14539 (N_14539,N_14396,N_14058);
nor U14540 (N_14540,N_14438,N_14360);
nand U14541 (N_14541,N_14001,N_14241);
nand U14542 (N_14542,N_14386,N_14155);
nor U14543 (N_14543,N_14444,N_14000);
and U14544 (N_14544,N_14202,N_14210);
xnor U14545 (N_14545,N_14323,N_14005);
and U14546 (N_14546,N_14458,N_14314);
and U14547 (N_14547,N_14078,N_14418);
nor U14548 (N_14548,N_14211,N_14459);
nor U14549 (N_14549,N_14395,N_14228);
nor U14550 (N_14550,N_14213,N_14247);
or U14551 (N_14551,N_14379,N_14095);
or U14552 (N_14552,N_14348,N_14429);
nand U14553 (N_14553,N_14385,N_14465);
nand U14554 (N_14554,N_14006,N_14384);
or U14555 (N_14555,N_14363,N_14134);
nor U14556 (N_14556,N_14439,N_14449);
and U14557 (N_14557,N_14034,N_14353);
nor U14558 (N_14558,N_14274,N_14303);
xor U14559 (N_14559,N_14481,N_14428);
and U14560 (N_14560,N_14357,N_14366);
nor U14561 (N_14561,N_14016,N_14089);
nand U14562 (N_14562,N_14435,N_14367);
or U14563 (N_14563,N_14491,N_14291);
or U14564 (N_14564,N_14473,N_14307);
xnor U14565 (N_14565,N_14086,N_14199);
and U14566 (N_14566,N_14132,N_14252);
nor U14567 (N_14567,N_14300,N_14180);
nor U14568 (N_14568,N_14341,N_14233);
nand U14569 (N_14569,N_14042,N_14264);
nand U14570 (N_14570,N_14441,N_14338);
nand U14571 (N_14571,N_14390,N_14302);
and U14572 (N_14572,N_14320,N_14182);
nor U14573 (N_14573,N_14335,N_14159);
xor U14574 (N_14574,N_14279,N_14499);
and U14575 (N_14575,N_14144,N_14455);
xnor U14576 (N_14576,N_14142,N_14286);
nand U14577 (N_14577,N_14343,N_14391);
or U14578 (N_14578,N_14110,N_14477);
xor U14579 (N_14579,N_14388,N_14200);
xor U14580 (N_14580,N_14258,N_14265);
xnor U14581 (N_14581,N_14061,N_14255);
xnor U14582 (N_14582,N_14167,N_14425);
and U14583 (N_14583,N_14071,N_14467);
and U14584 (N_14584,N_14209,N_14133);
xnor U14585 (N_14585,N_14328,N_14485);
xor U14586 (N_14586,N_14275,N_14246);
nor U14587 (N_14587,N_14108,N_14128);
and U14588 (N_14588,N_14178,N_14109);
nor U14589 (N_14589,N_14382,N_14044);
nor U14590 (N_14590,N_14074,N_14064);
xnor U14591 (N_14591,N_14053,N_14277);
or U14592 (N_14592,N_14020,N_14397);
nand U14593 (N_14593,N_14351,N_14411);
or U14594 (N_14594,N_14454,N_14126);
xor U14595 (N_14595,N_14179,N_14414);
nand U14596 (N_14596,N_14120,N_14245);
or U14597 (N_14597,N_14077,N_14267);
nand U14598 (N_14598,N_14280,N_14051);
or U14599 (N_14599,N_14035,N_14422);
xor U14600 (N_14600,N_14299,N_14032);
and U14601 (N_14601,N_14476,N_14461);
nand U14602 (N_14602,N_14378,N_14475);
and U14603 (N_14603,N_14065,N_14226);
or U14604 (N_14604,N_14099,N_14043);
and U14605 (N_14605,N_14446,N_14268);
nor U14606 (N_14606,N_14322,N_14118);
xnor U14607 (N_14607,N_14244,N_14436);
and U14608 (N_14608,N_14248,N_14023);
xor U14609 (N_14609,N_14494,N_14493);
nor U14610 (N_14610,N_14276,N_14057);
nand U14611 (N_14611,N_14153,N_14271);
nand U14612 (N_14612,N_14161,N_14229);
or U14613 (N_14613,N_14216,N_14009);
nor U14614 (N_14614,N_14138,N_14410);
xnor U14615 (N_14615,N_14249,N_14427);
nand U14616 (N_14616,N_14105,N_14272);
nand U14617 (N_14617,N_14084,N_14158);
nor U14618 (N_14618,N_14464,N_14266);
nor U14619 (N_14619,N_14301,N_14175);
xor U14620 (N_14620,N_14287,N_14297);
xnor U14621 (N_14621,N_14171,N_14219);
and U14622 (N_14622,N_14380,N_14104);
or U14623 (N_14623,N_14027,N_14457);
or U14624 (N_14624,N_14195,N_14047);
xor U14625 (N_14625,N_14092,N_14393);
or U14626 (N_14626,N_14137,N_14273);
xnor U14627 (N_14627,N_14448,N_14319);
or U14628 (N_14628,N_14140,N_14482);
nand U14629 (N_14629,N_14022,N_14069);
and U14630 (N_14630,N_14125,N_14176);
or U14631 (N_14631,N_14014,N_14193);
xnor U14632 (N_14632,N_14045,N_14318);
xnor U14633 (N_14633,N_14082,N_14203);
nand U14634 (N_14634,N_14381,N_14187);
or U14635 (N_14635,N_14344,N_14055);
nor U14636 (N_14636,N_14026,N_14260);
and U14637 (N_14637,N_14326,N_14288);
nand U14638 (N_14638,N_14298,N_14370);
nor U14639 (N_14639,N_14290,N_14037);
nand U14640 (N_14640,N_14173,N_14224);
xnor U14641 (N_14641,N_14062,N_14401);
or U14642 (N_14642,N_14164,N_14480);
nor U14643 (N_14643,N_14148,N_14090);
nand U14644 (N_14644,N_14431,N_14054);
nand U14645 (N_14645,N_14127,N_14313);
and U14646 (N_14646,N_14294,N_14150);
or U14647 (N_14647,N_14308,N_14129);
nor U14648 (N_14648,N_14371,N_14145);
nor U14649 (N_14649,N_14409,N_14204);
or U14650 (N_14650,N_14496,N_14445);
nand U14651 (N_14651,N_14143,N_14426);
xnor U14652 (N_14652,N_14408,N_14478);
or U14653 (N_14653,N_14490,N_14424);
and U14654 (N_14654,N_14282,N_14316);
xor U14655 (N_14655,N_14336,N_14355);
nor U14656 (N_14656,N_14072,N_14312);
or U14657 (N_14657,N_14234,N_14056);
xnor U14658 (N_14658,N_14434,N_14121);
xor U14659 (N_14659,N_14484,N_14135);
xor U14660 (N_14660,N_14170,N_14177);
xnor U14661 (N_14661,N_14471,N_14342);
nand U14662 (N_14662,N_14466,N_14106);
and U14663 (N_14663,N_14452,N_14327);
nor U14664 (N_14664,N_14430,N_14196);
and U14665 (N_14665,N_14221,N_14039);
nor U14666 (N_14666,N_14208,N_14281);
and U14667 (N_14667,N_14389,N_14004);
and U14668 (N_14668,N_14160,N_14031);
nor U14669 (N_14669,N_14050,N_14453);
nand U14670 (N_14670,N_14317,N_14021);
xnor U14671 (N_14671,N_14259,N_14304);
and U14672 (N_14672,N_14049,N_14024);
xnor U14673 (N_14673,N_14333,N_14091);
and U14674 (N_14674,N_14332,N_14151);
and U14675 (N_14675,N_14437,N_14112);
xnor U14676 (N_14676,N_14214,N_14474);
xor U14677 (N_14677,N_14420,N_14349);
xor U14678 (N_14678,N_14472,N_14130);
nand U14679 (N_14679,N_14169,N_14230);
nor U14680 (N_14680,N_14405,N_14076);
and U14681 (N_14681,N_14218,N_14331);
or U14682 (N_14682,N_14489,N_14403);
xor U14683 (N_14683,N_14124,N_14456);
nor U14684 (N_14684,N_14070,N_14399);
or U14685 (N_14685,N_14088,N_14460);
or U14686 (N_14686,N_14003,N_14407);
nor U14687 (N_14687,N_14269,N_14231);
xor U14688 (N_14688,N_14254,N_14237);
or U14689 (N_14689,N_14033,N_14345);
nand U14690 (N_14690,N_14008,N_14075);
and U14691 (N_14691,N_14183,N_14100);
and U14692 (N_14692,N_14207,N_14270);
nand U14693 (N_14693,N_14417,N_14463);
or U14694 (N_14694,N_14094,N_14066);
xnor U14695 (N_14695,N_14358,N_14415);
and U14696 (N_14696,N_14347,N_14283);
or U14697 (N_14697,N_14119,N_14398);
nand U14698 (N_14698,N_14097,N_14085);
xnor U14699 (N_14699,N_14165,N_14285);
or U14700 (N_14700,N_14292,N_14122);
or U14701 (N_14701,N_14350,N_14406);
nand U14702 (N_14702,N_14123,N_14262);
nand U14703 (N_14703,N_14174,N_14235);
xnor U14704 (N_14704,N_14046,N_14309);
xnor U14705 (N_14705,N_14450,N_14278);
nand U14706 (N_14706,N_14432,N_14156);
or U14707 (N_14707,N_14212,N_14030);
xor U14708 (N_14708,N_14402,N_14011);
or U14709 (N_14709,N_14240,N_14012);
or U14710 (N_14710,N_14131,N_14404);
xnor U14711 (N_14711,N_14073,N_14284);
nand U14712 (N_14712,N_14025,N_14157);
nand U14713 (N_14713,N_14369,N_14296);
xor U14714 (N_14714,N_14198,N_14015);
and U14715 (N_14715,N_14364,N_14413);
xor U14716 (N_14716,N_14115,N_14080);
xnor U14717 (N_14717,N_14215,N_14261);
or U14718 (N_14718,N_14400,N_14197);
and U14719 (N_14719,N_14019,N_14361);
nand U14720 (N_14720,N_14083,N_14242);
xor U14721 (N_14721,N_14339,N_14462);
xor U14722 (N_14722,N_14443,N_14311);
or U14723 (N_14723,N_14116,N_14306);
nor U14724 (N_14724,N_14227,N_14412);
nor U14725 (N_14725,N_14166,N_14352);
nor U14726 (N_14726,N_14356,N_14253);
nor U14727 (N_14727,N_14295,N_14487);
nand U14728 (N_14728,N_14029,N_14087);
nor U14729 (N_14729,N_14376,N_14324);
or U14730 (N_14730,N_14141,N_14190);
xnor U14731 (N_14731,N_14383,N_14250);
nand U14732 (N_14732,N_14423,N_14497);
nor U14733 (N_14733,N_14048,N_14321);
nand U14734 (N_14734,N_14373,N_14239);
xnor U14735 (N_14735,N_14096,N_14114);
nor U14736 (N_14736,N_14147,N_14117);
or U14737 (N_14737,N_14063,N_14018);
nand U14738 (N_14738,N_14068,N_14136);
or U14739 (N_14739,N_14359,N_14168);
nor U14740 (N_14740,N_14374,N_14257);
or U14741 (N_14741,N_14002,N_14081);
nor U14742 (N_14742,N_14362,N_14152);
or U14743 (N_14743,N_14223,N_14337);
xor U14744 (N_14744,N_14469,N_14191);
or U14745 (N_14745,N_14186,N_14479);
and U14746 (N_14746,N_14377,N_14263);
and U14747 (N_14747,N_14419,N_14205);
xor U14748 (N_14748,N_14329,N_14217);
or U14749 (N_14749,N_14238,N_14387);
and U14750 (N_14750,N_14134,N_14329);
and U14751 (N_14751,N_14163,N_14042);
or U14752 (N_14752,N_14109,N_14288);
and U14753 (N_14753,N_14276,N_14101);
and U14754 (N_14754,N_14416,N_14243);
xnor U14755 (N_14755,N_14444,N_14132);
and U14756 (N_14756,N_14012,N_14113);
and U14757 (N_14757,N_14298,N_14178);
nand U14758 (N_14758,N_14361,N_14327);
nand U14759 (N_14759,N_14118,N_14339);
and U14760 (N_14760,N_14050,N_14304);
nand U14761 (N_14761,N_14167,N_14211);
xor U14762 (N_14762,N_14351,N_14499);
and U14763 (N_14763,N_14137,N_14134);
nor U14764 (N_14764,N_14241,N_14273);
or U14765 (N_14765,N_14471,N_14319);
nand U14766 (N_14766,N_14050,N_14432);
nor U14767 (N_14767,N_14451,N_14345);
and U14768 (N_14768,N_14344,N_14241);
xor U14769 (N_14769,N_14101,N_14049);
or U14770 (N_14770,N_14061,N_14499);
nor U14771 (N_14771,N_14345,N_14167);
nand U14772 (N_14772,N_14296,N_14172);
or U14773 (N_14773,N_14483,N_14133);
xor U14774 (N_14774,N_14405,N_14416);
or U14775 (N_14775,N_14399,N_14260);
xnor U14776 (N_14776,N_14294,N_14149);
nand U14777 (N_14777,N_14425,N_14430);
nor U14778 (N_14778,N_14277,N_14069);
nor U14779 (N_14779,N_14384,N_14043);
nor U14780 (N_14780,N_14025,N_14463);
xor U14781 (N_14781,N_14394,N_14129);
nand U14782 (N_14782,N_14363,N_14227);
xor U14783 (N_14783,N_14022,N_14087);
nand U14784 (N_14784,N_14059,N_14443);
xnor U14785 (N_14785,N_14205,N_14483);
and U14786 (N_14786,N_14298,N_14465);
or U14787 (N_14787,N_14250,N_14271);
and U14788 (N_14788,N_14317,N_14453);
xnor U14789 (N_14789,N_14358,N_14429);
and U14790 (N_14790,N_14133,N_14452);
nor U14791 (N_14791,N_14228,N_14420);
nand U14792 (N_14792,N_14315,N_14265);
nor U14793 (N_14793,N_14009,N_14457);
and U14794 (N_14794,N_14384,N_14077);
or U14795 (N_14795,N_14464,N_14364);
nor U14796 (N_14796,N_14332,N_14470);
nor U14797 (N_14797,N_14469,N_14362);
nor U14798 (N_14798,N_14396,N_14317);
and U14799 (N_14799,N_14396,N_14212);
xnor U14800 (N_14800,N_14253,N_14446);
nand U14801 (N_14801,N_14391,N_14330);
nand U14802 (N_14802,N_14335,N_14147);
or U14803 (N_14803,N_14256,N_14325);
nand U14804 (N_14804,N_14052,N_14365);
and U14805 (N_14805,N_14079,N_14157);
and U14806 (N_14806,N_14476,N_14496);
xnor U14807 (N_14807,N_14289,N_14133);
and U14808 (N_14808,N_14294,N_14093);
nand U14809 (N_14809,N_14456,N_14397);
xnor U14810 (N_14810,N_14322,N_14359);
nand U14811 (N_14811,N_14102,N_14449);
nor U14812 (N_14812,N_14291,N_14273);
or U14813 (N_14813,N_14344,N_14326);
and U14814 (N_14814,N_14468,N_14144);
or U14815 (N_14815,N_14240,N_14105);
xor U14816 (N_14816,N_14485,N_14001);
or U14817 (N_14817,N_14229,N_14090);
or U14818 (N_14818,N_14370,N_14143);
nand U14819 (N_14819,N_14330,N_14006);
and U14820 (N_14820,N_14291,N_14308);
or U14821 (N_14821,N_14163,N_14409);
nand U14822 (N_14822,N_14390,N_14026);
and U14823 (N_14823,N_14078,N_14456);
or U14824 (N_14824,N_14082,N_14353);
and U14825 (N_14825,N_14243,N_14135);
or U14826 (N_14826,N_14481,N_14235);
xnor U14827 (N_14827,N_14322,N_14199);
xor U14828 (N_14828,N_14248,N_14192);
nand U14829 (N_14829,N_14174,N_14341);
nor U14830 (N_14830,N_14077,N_14246);
and U14831 (N_14831,N_14025,N_14389);
and U14832 (N_14832,N_14050,N_14061);
or U14833 (N_14833,N_14246,N_14440);
and U14834 (N_14834,N_14265,N_14395);
and U14835 (N_14835,N_14448,N_14331);
or U14836 (N_14836,N_14003,N_14424);
and U14837 (N_14837,N_14402,N_14375);
and U14838 (N_14838,N_14458,N_14442);
nand U14839 (N_14839,N_14061,N_14077);
nor U14840 (N_14840,N_14325,N_14271);
nand U14841 (N_14841,N_14352,N_14239);
and U14842 (N_14842,N_14201,N_14098);
nand U14843 (N_14843,N_14126,N_14343);
nand U14844 (N_14844,N_14194,N_14451);
nand U14845 (N_14845,N_14442,N_14062);
and U14846 (N_14846,N_14300,N_14351);
or U14847 (N_14847,N_14147,N_14438);
nor U14848 (N_14848,N_14413,N_14363);
xor U14849 (N_14849,N_14247,N_14167);
and U14850 (N_14850,N_14461,N_14279);
or U14851 (N_14851,N_14282,N_14310);
nand U14852 (N_14852,N_14221,N_14423);
nand U14853 (N_14853,N_14326,N_14246);
and U14854 (N_14854,N_14348,N_14499);
nand U14855 (N_14855,N_14473,N_14054);
and U14856 (N_14856,N_14052,N_14009);
or U14857 (N_14857,N_14228,N_14279);
nand U14858 (N_14858,N_14443,N_14404);
nor U14859 (N_14859,N_14426,N_14226);
xnor U14860 (N_14860,N_14041,N_14151);
xnor U14861 (N_14861,N_14329,N_14397);
and U14862 (N_14862,N_14313,N_14135);
nor U14863 (N_14863,N_14438,N_14093);
and U14864 (N_14864,N_14189,N_14359);
nand U14865 (N_14865,N_14466,N_14114);
and U14866 (N_14866,N_14135,N_14389);
xor U14867 (N_14867,N_14101,N_14271);
or U14868 (N_14868,N_14298,N_14378);
and U14869 (N_14869,N_14300,N_14089);
or U14870 (N_14870,N_14226,N_14085);
or U14871 (N_14871,N_14493,N_14393);
and U14872 (N_14872,N_14424,N_14227);
or U14873 (N_14873,N_14408,N_14410);
or U14874 (N_14874,N_14286,N_14038);
or U14875 (N_14875,N_14186,N_14099);
or U14876 (N_14876,N_14386,N_14422);
or U14877 (N_14877,N_14030,N_14055);
xor U14878 (N_14878,N_14089,N_14315);
xor U14879 (N_14879,N_14381,N_14274);
and U14880 (N_14880,N_14258,N_14494);
or U14881 (N_14881,N_14336,N_14325);
nand U14882 (N_14882,N_14322,N_14281);
or U14883 (N_14883,N_14195,N_14378);
nor U14884 (N_14884,N_14134,N_14451);
nor U14885 (N_14885,N_14242,N_14140);
nor U14886 (N_14886,N_14177,N_14153);
xnor U14887 (N_14887,N_14226,N_14353);
nand U14888 (N_14888,N_14260,N_14417);
xnor U14889 (N_14889,N_14103,N_14084);
or U14890 (N_14890,N_14105,N_14238);
and U14891 (N_14891,N_14281,N_14051);
nand U14892 (N_14892,N_14192,N_14060);
nor U14893 (N_14893,N_14069,N_14317);
and U14894 (N_14894,N_14270,N_14151);
xor U14895 (N_14895,N_14410,N_14496);
nor U14896 (N_14896,N_14111,N_14407);
nor U14897 (N_14897,N_14456,N_14424);
xor U14898 (N_14898,N_14359,N_14096);
and U14899 (N_14899,N_14227,N_14198);
xor U14900 (N_14900,N_14273,N_14470);
and U14901 (N_14901,N_14151,N_14108);
nand U14902 (N_14902,N_14233,N_14187);
and U14903 (N_14903,N_14066,N_14293);
nor U14904 (N_14904,N_14290,N_14331);
nor U14905 (N_14905,N_14358,N_14108);
nor U14906 (N_14906,N_14333,N_14482);
or U14907 (N_14907,N_14142,N_14073);
nand U14908 (N_14908,N_14465,N_14403);
nand U14909 (N_14909,N_14190,N_14205);
nor U14910 (N_14910,N_14158,N_14288);
nor U14911 (N_14911,N_14029,N_14377);
or U14912 (N_14912,N_14305,N_14129);
or U14913 (N_14913,N_14377,N_14097);
and U14914 (N_14914,N_14179,N_14354);
nand U14915 (N_14915,N_14458,N_14118);
and U14916 (N_14916,N_14206,N_14448);
and U14917 (N_14917,N_14006,N_14276);
xor U14918 (N_14918,N_14381,N_14382);
xnor U14919 (N_14919,N_14498,N_14337);
xnor U14920 (N_14920,N_14301,N_14072);
or U14921 (N_14921,N_14422,N_14235);
or U14922 (N_14922,N_14065,N_14123);
nor U14923 (N_14923,N_14105,N_14329);
or U14924 (N_14924,N_14321,N_14111);
nand U14925 (N_14925,N_14197,N_14029);
nor U14926 (N_14926,N_14388,N_14341);
nor U14927 (N_14927,N_14209,N_14446);
nor U14928 (N_14928,N_14472,N_14326);
nand U14929 (N_14929,N_14231,N_14342);
nand U14930 (N_14930,N_14227,N_14449);
nand U14931 (N_14931,N_14445,N_14247);
or U14932 (N_14932,N_14491,N_14420);
nand U14933 (N_14933,N_14312,N_14275);
nor U14934 (N_14934,N_14275,N_14130);
xor U14935 (N_14935,N_14177,N_14420);
and U14936 (N_14936,N_14051,N_14009);
nand U14937 (N_14937,N_14152,N_14143);
and U14938 (N_14938,N_14414,N_14220);
nor U14939 (N_14939,N_14330,N_14147);
nor U14940 (N_14940,N_14344,N_14202);
or U14941 (N_14941,N_14418,N_14236);
and U14942 (N_14942,N_14282,N_14307);
xor U14943 (N_14943,N_14413,N_14236);
and U14944 (N_14944,N_14286,N_14383);
nand U14945 (N_14945,N_14013,N_14301);
nor U14946 (N_14946,N_14281,N_14238);
nand U14947 (N_14947,N_14287,N_14352);
nand U14948 (N_14948,N_14298,N_14372);
nor U14949 (N_14949,N_14148,N_14061);
xnor U14950 (N_14950,N_14165,N_14104);
and U14951 (N_14951,N_14247,N_14376);
and U14952 (N_14952,N_14188,N_14484);
nand U14953 (N_14953,N_14232,N_14278);
nor U14954 (N_14954,N_14093,N_14470);
and U14955 (N_14955,N_14370,N_14092);
or U14956 (N_14956,N_14145,N_14386);
nand U14957 (N_14957,N_14173,N_14047);
nor U14958 (N_14958,N_14180,N_14408);
or U14959 (N_14959,N_14497,N_14406);
nand U14960 (N_14960,N_14061,N_14115);
or U14961 (N_14961,N_14471,N_14217);
or U14962 (N_14962,N_14470,N_14034);
or U14963 (N_14963,N_14095,N_14359);
xor U14964 (N_14964,N_14193,N_14226);
nor U14965 (N_14965,N_14422,N_14241);
nor U14966 (N_14966,N_14095,N_14443);
nand U14967 (N_14967,N_14090,N_14248);
and U14968 (N_14968,N_14421,N_14401);
xnor U14969 (N_14969,N_14026,N_14268);
and U14970 (N_14970,N_14041,N_14103);
nand U14971 (N_14971,N_14492,N_14347);
xor U14972 (N_14972,N_14117,N_14214);
nor U14973 (N_14973,N_14393,N_14229);
and U14974 (N_14974,N_14388,N_14437);
nor U14975 (N_14975,N_14191,N_14383);
xnor U14976 (N_14976,N_14325,N_14465);
xor U14977 (N_14977,N_14248,N_14393);
xnor U14978 (N_14978,N_14391,N_14357);
xor U14979 (N_14979,N_14051,N_14224);
nor U14980 (N_14980,N_14206,N_14099);
nor U14981 (N_14981,N_14291,N_14476);
nor U14982 (N_14982,N_14454,N_14094);
and U14983 (N_14983,N_14211,N_14033);
or U14984 (N_14984,N_14267,N_14430);
or U14985 (N_14985,N_14487,N_14337);
or U14986 (N_14986,N_14350,N_14460);
xor U14987 (N_14987,N_14428,N_14138);
nand U14988 (N_14988,N_14026,N_14455);
or U14989 (N_14989,N_14194,N_14140);
xnor U14990 (N_14990,N_14318,N_14382);
nor U14991 (N_14991,N_14131,N_14244);
or U14992 (N_14992,N_14429,N_14295);
nor U14993 (N_14993,N_14300,N_14413);
nand U14994 (N_14994,N_14469,N_14451);
nor U14995 (N_14995,N_14188,N_14398);
and U14996 (N_14996,N_14009,N_14169);
or U14997 (N_14997,N_14124,N_14310);
nor U14998 (N_14998,N_14340,N_14251);
and U14999 (N_14999,N_14050,N_14193);
and U15000 (N_15000,N_14895,N_14819);
nor U15001 (N_15001,N_14823,N_14655);
or U15002 (N_15002,N_14536,N_14618);
xnor U15003 (N_15003,N_14999,N_14758);
xnor U15004 (N_15004,N_14740,N_14575);
nor U15005 (N_15005,N_14573,N_14725);
xor U15006 (N_15006,N_14570,N_14809);
and U15007 (N_15007,N_14843,N_14961);
xor U15008 (N_15008,N_14764,N_14612);
nand U15009 (N_15009,N_14556,N_14718);
nand U15010 (N_15010,N_14840,N_14951);
xor U15011 (N_15011,N_14811,N_14514);
xor U15012 (N_15012,N_14945,N_14771);
or U15013 (N_15013,N_14683,N_14689);
or U15014 (N_15014,N_14878,N_14603);
and U15015 (N_15015,N_14883,N_14673);
or U15016 (N_15016,N_14555,N_14580);
nor U15017 (N_15017,N_14589,N_14972);
or U15018 (N_15018,N_14572,N_14942);
xnor U15019 (N_15019,N_14520,N_14682);
and U15020 (N_15020,N_14909,N_14834);
and U15021 (N_15021,N_14502,N_14808);
nor U15022 (N_15022,N_14513,N_14537);
xnor U15023 (N_15023,N_14962,N_14671);
xor U15024 (N_15024,N_14845,N_14893);
xnor U15025 (N_15025,N_14696,N_14896);
or U15026 (N_15026,N_14914,N_14892);
or U15027 (N_15027,N_14727,N_14676);
nand U15028 (N_15028,N_14897,N_14850);
xnor U15029 (N_15029,N_14783,N_14762);
xor U15030 (N_15030,N_14684,N_14623);
and U15031 (N_15031,N_14967,N_14544);
nand U15032 (N_15032,N_14692,N_14973);
and U15033 (N_15033,N_14855,N_14937);
nor U15034 (N_15034,N_14785,N_14821);
and U15035 (N_15035,N_14919,N_14759);
nand U15036 (N_15036,N_14630,N_14917);
xnor U15037 (N_15037,N_14867,N_14699);
or U15038 (N_15038,N_14741,N_14711);
xor U15039 (N_15039,N_14936,N_14516);
and U15040 (N_15040,N_14722,N_14985);
or U15041 (N_15041,N_14697,N_14698);
xnor U15042 (N_15042,N_14694,N_14990);
and U15043 (N_15043,N_14506,N_14702);
nor U15044 (N_15044,N_14902,N_14661);
nand U15045 (N_15045,N_14614,N_14719);
and U15046 (N_15046,N_14974,N_14866);
nor U15047 (N_15047,N_14779,N_14794);
nand U15048 (N_15048,N_14593,N_14549);
nor U15049 (N_15049,N_14775,N_14943);
and U15050 (N_15050,N_14731,N_14645);
and U15051 (N_15051,N_14828,N_14955);
nand U15052 (N_15052,N_14761,N_14713);
and U15053 (N_15053,N_14818,N_14568);
nor U15054 (N_15054,N_14726,N_14585);
xor U15055 (N_15055,N_14865,N_14879);
xor U15056 (N_15056,N_14611,N_14958);
xnor U15057 (N_15057,N_14838,N_14742);
nor U15058 (N_15058,N_14610,N_14939);
nand U15059 (N_15059,N_14515,N_14875);
and U15060 (N_15060,N_14748,N_14858);
and U15061 (N_15061,N_14518,N_14813);
nor U15062 (N_15062,N_14523,N_14924);
nor U15063 (N_15063,N_14640,N_14647);
and U15064 (N_15064,N_14721,N_14983);
nor U15065 (N_15065,N_14601,N_14591);
xor U15066 (N_15066,N_14929,N_14842);
and U15067 (N_15067,N_14859,N_14900);
xnor U15068 (N_15068,N_14534,N_14669);
nor U15069 (N_15069,N_14885,N_14869);
nor U15070 (N_15070,N_14784,N_14714);
nor U15071 (N_15071,N_14586,N_14795);
xor U15072 (N_15072,N_14712,N_14576);
and U15073 (N_15073,N_14932,N_14868);
nand U15074 (N_15074,N_14604,N_14801);
nor U15075 (N_15075,N_14639,N_14977);
xnor U15076 (N_15076,N_14982,N_14565);
nor U15077 (N_15077,N_14938,N_14826);
nor U15078 (N_15078,N_14531,N_14815);
nor U15079 (N_15079,N_14541,N_14677);
or U15080 (N_15080,N_14554,N_14501);
xor U15081 (N_15081,N_14707,N_14540);
or U15082 (N_15082,N_14927,N_14915);
xnor U15083 (N_15083,N_14642,N_14691);
or U15084 (N_15084,N_14563,N_14978);
nand U15085 (N_15085,N_14605,N_14754);
nand U15086 (N_15086,N_14786,N_14873);
nor U15087 (N_15087,N_14600,N_14538);
and U15088 (N_15088,N_14552,N_14728);
nor U15089 (N_15089,N_14646,N_14749);
or U15090 (N_15090,N_14899,N_14609);
or U15091 (N_15091,N_14856,N_14949);
nand U15092 (N_15092,N_14824,N_14629);
xor U15093 (N_15093,N_14874,N_14995);
nor U15094 (N_15094,N_14652,N_14948);
or U15095 (N_15095,N_14579,N_14720);
nand U15096 (N_15096,N_14527,N_14814);
xor U15097 (N_15097,N_14510,N_14577);
or U15098 (N_15098,N_14686,N_14539);
or U15099 (N_15099,N_14680,N_14916);
nand U15100 (N_15100,N_14690,N_14863);
nor U15101 (N_15101,N_14578,N_14964);
xnor U15102 (N_15102,N_14913,N_14559);
and U15103 (N_15103,N_14822,N_14947);
xor U15104 (N_15104,N_14550,N_14921);
nor U15105 (N_15105,N_14888,N_14566);
and U15106 (N_15106,N_14970,N_14653);
and U15107 (N_15107,N_14997,N_14649);
nor U15108 (N_15108,N_14812,N_14656);
xor U15109 (N_15109,N_14998,N_14674);
nor U15110 (N_15110,N_14700,N_14789);
or U15111 (N_15111,N_14980,N_14723);
nand U15112 (N_15112,N_14882,N_14852);
nand U15113 (N_15113,N_14993,N_14592);
nor U15114 (N_15114,N_14954,N_14542);
and U15115 (N_15115,N_14984,N_14525);
or U15116 (N_15116,N_14716,N_14912);
and U15117 (N_15117,N_14830,N_14880);
nand U15118 (N_15118,N_14839,N_14637);
nand U15119 (N_15119,N_14901,N_14767);
nand U15120 (N_15120,N_14654,N_14930);
or U15121 (N_15121,N_14791,N_14772);
xnor U15122 (N_15122,N_14807,N_14898);
and U15123 (N_15123,N_14597,N_14774);
nor U15124 (N_15124,N_14724,N_14551);
nor U15125 (N_15125,N_14991,N_14746);
and U15126 (N_15126,N_14768,N_14918);
and U15127 (N_15127,N_14827,N_14558);
or U15128 (N_15128,N_14756,N_14946);
and U15129 (N_15129,N_14848,N_14633);
nor U15130 (N_15130,N_14781,N_14735);
xor U15131 (N_15131,N_14667,N_14799);
nand U15132 (N_15132,N_14891,N_14574);
or U15133 (N_15133,N_14904,N_14619);
nor U15134 (N_15134,N_14910,N_14889);
xor U15135 (N_15135,N_14769,N_14533);
xnor U15136 (N_15136,N_14590,N_14928);
nor U15137 (N_15137,N_14715,N_14626);
or U15138 (N_15138,N_14975,N_14841);
xnor U15139 (N_15139,N_14968,N_14766);
or U15140 (N_15140,N_14695,N_14584);
nor U15141 (N_15141,N_14582,N_14734);
nand U15142 (N_15142,N_14624,N_14636);
nand U15143 (N_15143,N_14557,N_14934);
nand U15144 (N_15144,N_14641,N_14860);
nand U15145 (N_15145,N_14805,N_14744);
nand U15146 (N_15146,N_14569,N_14545);
nand U15147 (N_15147,N_14787,N_14836);
nand U15148 (N_15148,N_14599,N_14730);
nor U15149 (N_15149,N_14511,N_14509);
nand U15150 (N_15150,N_14562,N_14737);
nor U15151 (N_15151,N_14581,N_14923);
nand U15152 (N_15152,N_14595,N_14687);
xor U15153 (N_15153,N_14648,N_14663);
xor U15154 (N_15154,N_14672,N_14708);
nand U15155 (N_15155,N_14733,N_14810);
nand U15156 (N_15156,N_14616,N_14703);
xor U15157 (N_15157,N_14753,N_14598);
or U15158 (N_15158,N_14905,N_14522);
or U15159 (N_15159,N_14628,N_14956);
nand U15160 (N_15160,N_14802,N_14876);
or U15161 (N_15161,N_14662,N_14907);
xnor U15162 (N_15162,N_14906,N_14884);
xnor U15163 (N_15163,N_14681,N_14627);
nand U15164 (N_15164,N_14517,N_14894);
or U15165 (N_15165,N_14665,N_14931);
nand U15166 (N_15166,N_14659,N_14903);
and U15167 (N_15167,N_14857,N_14701);
nor U15168 (N_15168,N_14886,N_14816);
xnor U15169 (N_15169,N_14763,N_14751);
nor U15170 (N_15170,N_14911,N_14944);
or U15171 (N_15171,N_14844,N_14757);
or U15172 (N_15172,N_14793,N_14650);
and U15173 (N_15173,N_14871,N_14745);
or U15174 (N_15174,N_14685,N_14588);
nand U15175 (N_15175,N_14760,N_14941);
nand U15176 (N_15176,N_14804,N_14981);
xnor U15177 (N_15177,N_14853,N_14979);
and U15178 (N_15178,N_14803,N_14500);
or U15179 (N_15179,N_14738,N_14658);
and U15180 (N_15180,N_14782,N_14847);
xor U15181 (N_15181,N_14529,N_14553);
and U15182 (N_15182,N_14837,N_14908);
nor U15183 (N_15183,N_14966,N_14561);
xnor U15184 (N_15184,N_14583,N_14709);
and U15185 (N_15185,N_14688,N_14851);
nand U15186 (N_15186,N_14790,N_14528);
or U15187 (N_15187,N_14644,N_14953);
nand U15188 (N_15188,N_14959,N_14957);
and U15189 (N_15189,N_14776,N_14526);
xor U15190 (N_15190,N_14752,N_14988);
xor U15191 (N_15191,N_14987,N_14732);
and U15192 (N_15192,N_14971,N_14922);
or U15193 (N_15193,N_14770,N_14620);
or U15194 (N_15194,N_14831,N_14989);
and U15195 (N_15195,N_14530,N_14532);
or U15196 (N_15196,N_14773,N_14524);
and U15197 (N_15197,N_14567,N_14736);
nor U15198 (N_15198,N_14613,N_14710);
xor U15199 (N_15199,N_14704,N_14833);
nand U15200 (N_15200,N_14963,N_14854);
or U15201 (N_15201,N_14625,N_14777);
nand U15202 (N_15202,N_14564,N_14890);
and U15203 (N_15203,N_14606,N_14617);
nand U15204 (N_15204,N_14920,N_14615);
nor U15205 (N_15205,N_14634,N_14935);
nand U15206 (N_15206,N_14986,N_14643);
xnor U15207 (N_15207,N_14996,N_14675);
nor U15208 (N_15208,N_14832,N_14512);
xor U15209 (N_15209,N_14587,N_14792);
xnor U15210 (N_15210,N_14602,N_14846);
and U15211 (N_15211,N_14797,N_14668);
and U15212 (N_15212,N_14825,N_14705);
or U15213 (N_15213,N_14750,N_14806);
xor U15214 (N_15214,N_14950,N_14965);
nand U15215 (N_15215,N_14861,N_14817);
nor U15216 (N_15216,N_14664,N_14622);
xnor U15217 (N_15217,N_14925,N_14596);
xor U15218 (N_15218,N_14835,N_14706);
nand U15219 (N_15219,N_14849,N_14547);
and U15220 (N_15220,N_14829,N_14546);
or U15221 (N_15221,N_14505,N_14543);
xnor U15222 (N_15222,N_14679,N_14952);
or U15223 (N_15223,N_14635,N_14994);
or U15224 (N_15224,N_14631,N_14969);
or U15225 (N_15225,N_14670,N_14503);
and U15226 (N_15226,N_14594,N_14508);
nor U15227 (N_15227,N_14608,N_14666);
nor U15228 (N_15228,N_14881,N_14521);
nor U15229 (N_15229,N_14743,N_14877);
nand U15230 (N_15230,N_14507,N_14657);
nand U15231 (N_15231,N_14548,N_14870);
xnor U15232 (N_15232,N_14638,N_14504);
nand U15233 (N_15233,N_14739,N_14820);
xnor U15234 (N_15234,N_14519,N_14621);
nor U15235 (N_15235,N_14788,N_14571);
nand U15236 (N_15236,N_14780,N_14926);
nor U15237 (N_15237,N_14864,N_14862);
nor U15238 (N_15238,N_14607,N_14560);
nand U15239 (N_15239,N_14678,N_14632);
or U15240 (N_15240,N_14660,N_14798);
and U15241 (N_15241,N_14778,N_14535);
nor U15242 (N_15242,N_14933,N_14800);
nor U15243 (N_15243,N_14796,N_14717);
nand U15244 (N_15244,N_14693,N_14960);
nor U15245 (N_15245,N_14747,N_14651);
nor U15246 (N_15246,N_14887,N_14755);
nor U15247 (N_15247,N_14992,N_14765);
and U15248 (N_15248,N_14729,N_14872);
and U15249 (N_15249,N_14940,N_14976);
xor U15250 (N_15250,N_14712,N_14862);
nor U15251 (N_15251,N_14656,N_14713);
or U15252 (N_15252,N_14638,N_14737);
and U15253 (N_15253,N_14634,N_14604);
and U15254 (N_15254,N_14716,N_14666);
xnor U15255 (N_15255,N_14698,N_14846);
nor U15256 (N_15256,N_14744,N_14782);
and U15257 (N_15257,N_14686,N_14703);
or U15258 (N_15258,N_14788,N_14599);
or U15259 (N_15259,N_14722,N_14874);
nor U15260 (N_15260,N_14992,N_14877);
xor U15261 (N_15261,N_14900,N_14929);
nand U15262 (N_15262,N_14828,N_14529);
nor U15263 (N_15263,N_14593,N_14906);
or U15264 (N_15264,N_14912,N_14640);
xor U15265 (N_15265,N_14652,N_14786);
or U15266 (N_15266,N_14838,N_14713);
nor U15267 (N_15267,N_14548,N_14623);
or U15268 (N_15268,N_14800,N_14627);
nand U15269 (N_15269,N_14509,N_14968);
and U15270 (N_15270,N_14790,N_14957);
xnor U15271 (N_15271,N_14921,N_14710);
and U15272 (N_15272,N_14809,N_14981);
nand U15273 (N_15273,N_14772,N_14624);
xnor U15274 (N_15274,N_14787,N_14825);
or U15275 (N_15275,N_14667,N_14997);
nand U15276 (N_15276,N_14928,N_14580);
nand U15277 (N_15277,N_14904,N_14726);
or U15278 (N_15278,N_14615,N_14590);
nand U15279 (N_15279,N_14781,N_14536);
and U15280 (N_15280,N_14519,N_14598);
nand U15281 (N_15281,N_14684,N_14707);
nand U15282 (N_15282,N_14753,N_14965);
nand U15283 (N_15283,N_14926,N_14955);
or U15284 (N_15284,N_14528,N_14621);
nor U15285 (N_15285,N_14517,N_14811);
xor U15286 (N_15286,N_14566,N_14787);
or U15287 (N_15287,N_14995,N_14621);
xor U15288 (N_15288,N_14616,N_14599);
or U15289 (N_15289,N_14857,N_14585);
nor U15290 (N_15290,N_14539,N_14607);
nand U15291 (N_15291,N_14502,N_14723);
xor U15292 (N_15292,N_14562,N_14799);
or U15293 (N_15293,N_14974,N_14631);
and U15294 (N_15294,N_14512,N_14997);
and U15295 (N_15295,N_14779,N_14572);
nor U15296 (N_15296,N_14647,N_14741);
xor U15297 (N_15297,N_14734,N_14790);
xnor U15298 (N_15298,N_14771,N_14892);
nor U15299 (N_15299,N_14942,N_14805);
or U15300 (N_15300,N_14962,N_14971);
nor U15301 (N_15301,N_14996,N_14841);
nand U15302 (N_15302,N_14718,N_14899);
xor U15303 (N_15303,N_14717,N_14919);
or U15304 (N_15304,N_14849,N_14847);
and U15305 (N_15305,N_14802,N_14761);
nor U15306 (N_15306,N_14536,N_14631);
nand U15307 (N_15307,N_14974,N_14943);
and U15308 (N_15308,N_14828,N_14590);
nand U15309 (N_15309,N_14505,N_14646);
or U15310 (N_15310,N_14755,N_14813);
and U15311 (N_15311,N_14916,N_14824);
nand U15312 (N_15312,N_14572,N_14667);
nor U15313 (N_15313,N_14964,N_14698);
xor U15314 (N_15314,N_14779,N_14760);
nor U15315 (N_15315,N_14949,N_14757);
and U15316 (N_15316,N_14940,N_14519);
nand U15317 (N_15317,N_14992,N_14824);
and U15318 (N_15318,N_14986,N_14543);
nor U15319 (N_15319,N_14531,N_14821);
and U15320 (N_15320,N_14753,N_14974);
nor U15321 (N_15321,N_14896,N_14600);
and U15322 (N_15322,N_14585,N_14946);
and U15323 (N_15323,N_14937,N_14959);
or U15324 (N_15324,N_14883,N_14669);
nand U15325 (N_15325,N_14978,N_14998);
nand U15326 (N_15326,N_14671,N_14829);
nor U15327 (N_15327,N_14823,N_14989);
nand U15328 (N_15328,N_14602,N_14780);
and U15329 (N_15329,N_14713,N_14625);
nand U15330 (N_15330,N_14772,N_14634);
or U15331 (N_15331,N_14903,N_14600);
nor U15332 (N_15332,N_14938,N_14539);
nand U15333 (N_15333,N_14970,N_14837);
or U15334 (N_15334,N_14934,N_14602);
xor U15335 (N_15335,N_14782,N_14932);
and U15336 (N_15336,N_14942,N_14525);
nand U15337 (N_15337,N_14929,N_14702);
nor U15338 (N_15338,N_14697,N_14729);
nand U15339 (N_15339,N_14749,N_14503);
xnor U15340 (N_15340,N_14643,N_14735);
and U15341 (N_15341,N_14658,N_14919);
nand U15342 (N_15342,N_14700,N_14626);
and U15343 (N_15343,N_14539,N_14799);
nand U15344 (N_15344,N_14958,N_14894);
nor U15345 (N_15345,N_14998,N_14881);
nor U15346 (N_15346,N_14645,N_14696);
nand U15347 (N_15347,N_14848,N_14551);
nand U15348 (N_15348,N_14983,N_14549);
nor U15349 (N_15349,N_14636,N_14686);
or U15350 (N_15350,N_14769,N_14846);
and U15351 (N_15351,N_14742,N_14824);
or U15352 (N_15352,N_14785,N_14736);
nand U15353 (N_15353,N_14506,N_14630);
nor U15354 (N_15354,N_14537,N_14762);
nand U15355 (N_15355,N_14658,N_14982);
nor U15356 (N_15356,N_14513,N_14900);
or U15357 (N_15357,N_14834,N_14663);
nor U15358 (N_15358,N_14748,N_14854);
xor U15359 (N_15359,N_14765,N_14984);
or U15360 (N_15360,N_14507,N_14969);
nand U15361 (N_15361,N_14550,N_14905);
nand U15362 (N_15362,N_14748,N_14712);
nor U15363 (N_15363,N_14796,N_14803);
nor U15364 (N_15364,N_14756,N_14930);
and U15365 (N_15365,N_14510,N_14643);
xor U15366 (N_15366,N_14929,N_14616);
xor U15367 (N_15367,N_14832,N_14718);
nand U15368 (N_15368,N_14544,N_14928);
nand U15369 (N_15369,N_14598,N_14572);
xor U15370 (N_15370,N_14728,N_14947);
or U15371 (N_15371,N_14517,N_14738);
xnor U15372 (N_15372,N_14943,N_14736);
nor U15373 (N_15373,N_14573,N_14636);
xor U15374 (N_15374,N_14999,N_14976);
xnor U15375 (N_15375,N_14969,N_14749);
and U15376 (N_15376,N_14937,N_14973);
and U15377 (N_15377,N_14840,N_14916);
nand U15378 (N_15378,N_14735,N_14829);
nand U15379 (N_15379,N_14577,N_14956);
xor U15380 (N_15380,N_14787,N_14677);
xor U15381 (N_15381,N_14894,N_14812);
and U15382 (N_15382,N_14698,N_14710);
and U15383 (N_15383,N_14526,N_14742);
xnor U15384 (N_15384,N_14667,N_14605);
or U15385 (N_15385,N_14917,N_14874);
nor U15386 (N_15386,N_14776,N_14549);
nor U15387 (N_15387,N_14641,N_14622);
or U15388 (N_15388,N_14957,N_14838);
or U15389 (N_15389,N_14983,N_14803);
nor U15390 (N_15390,N_14807,N_14961);
or U15391 (N_15391,N_14963,N_14622);
or U15392 (N_15392,N_14780,N_14658);
nand U15393 (N_15393,N_14880,N_14647);
or U15394 (N_15394,N_14603,N_14618);
and U15395 (N_15395,N_14651,N_14700);
nor U15396 (N_15396,N_14579,N_14994);
xor U15397 (N_15397,N_14844,N_14645);
xor U15398 (N_15398,N_14822,N_14608);
xor U15399 (N_15399,N_14577,N_14751);
nor U15400 (N_15400,N_14880,N_14906);
xnor U15401 (N_15401,N_14928,N_14899);
or U15402 (N_15402,N_14700,N_14872);
and U15403 (N_15403,N_14597,N_14864);
and U15404 (N_15404,N_14922,N_14520);
nand U15405 (N_15405,N_14518,N_14753);
xnor U15406 (N_15406,N_14644,N_14756);
nor U15407 (N_15407,N_14676,N_14997);
or U15408 (N_15408,N_14503,N_14969);
nor U15409 (N_15409,N_14806,N_14616);
nand U15410 (N_15410,N_14593,N_14808);
nand U15411 (N_15411,N_14915,N_14666);
xor U15412 (N_15412,N_14908,N_14887);
xnor U15413 (N_15413,N_14980,N_14512);
nand U15414 (N_15414,N_14519,N_14733);
nor U15415 (N_15415,N_14691,N_14720);
and U15416 (N_15416,N_14608,N_14549);
or U15417 (N_15417,N_14582,N_14941);
nor U15418 (N_15418,N_14754,N_14995);
nand U15419 (N_15419,N_14909,N_14667);
nor U15420 (N_15420,N_14584,N_14668);
nor U15421 (N_15421,N_14749,N_14522);
nand U15422 (N_15422,N_14737,N_14618);
xnor U15423 (N_15423,N_14796,N_14830);
xor U15424 (N_15424,N_14658,N_14886);
nand U15425 (N_15425,N_14903,N_14999);
and U15426 (N_15426,N_14892,N_14750);
xor U15427 (N_15427,N_14628,N_14969);
nor U15428 (N_15428,N_14737,N_14686);
xor U15429 (N_15429,N_14531,N_14535);
and U15430 (N_15430,N_14991,N_14525);
nand U15431 (N_15431,N_14883,N_14719);
xnor U15432 (N_15432,N_14644,N_14505);
and U15433 (N_15433,N_14937,N_14604);
xor U15434 (N_15434,N_14653,N_14936);
or U15435 (N_15435,N_14597,N_14748);
xnor U15436 (N_15436,N_14573,N_14586);
nand U15437 (N_15437,N_14574,N_14736);
and U15438 (N_15438,N_14924,N_14859);
xor U15439 (N_15439,N_14621,N_14789);
nor U15440 (N_15440,N_14537,N_14823);
nor U15441 (N_15441,N_14909,N_14506);
nand U15442 (N_15442,N_14674,N_14839);
xnor U15443 (N_15443,N_14886,N_14652);
nor U15444 (N_15444,N_14575,N_14633);
xor U15445 (N_15445,N_14653,N_14881);
and U15446 (N_15446,N_14571,N_14607);
or U15447 (N_15447,N_14516,N_14688);
nand U15448 (N_15448,N_14567,N_14500);
nand U15449 (N_15449,N_14566,N_14889);
nor U15450 (N_15450,N_14897,N_14508);
or U15451 (N_15451,N_14987,N_14971);
xnor U15452 (N_15452,N_14527,N_14622);
and U15453 (N_15453,N_14559,N_14532);
and U15454 (N_15454,N_14916,N_14644);
or U15455 (N_15455,N_14940,N_14863);
and U15456 (N_15456,N_14880,N_14678);
xnor U15457 (N_15457,N_14680,N_14822);
xnor U15458 (N_15458,N_14866,N_14679);
or U15459 (N_15459,N_14507,N_14863);
or U15460 (N_15460,N_14996,N_14812);
xnor U15461 (N_15461,N_14892,N_14513);
nand U15462 (N_15462,N_14699,N_14720);
or U15463 (N_15463,N_14655,N_14777);
nand U15464 (N_15464,N_14665,N_14747);
and U15465 (N_15465,N_14570,N_14914);
and U15466 (N_15466,N_14882,N_14758);
and U15467 (N_15467,N_14882,N_14735);
xor U15468 (N_15468,N_14829,N_14995);
xor U15469 (N_15469,N_14588,N_14696);
nand U15470 (N_15470,N_14604,N_14792);
and U15471 (N_15471,N_14747,N_14813);
nor U15472 (N_15472,N_14581,N_14928);
nor U15473 (N_15473,N_14665,N_14830);
nor U15474 (N_15474,N_14941,N_14658);
and U15475 (N_15475,N_14651,N_14858);
or U15476 (N_15476,N_14796,N_14963);
xor U15477 (N_15477,N_14554,N_14758);
xor U15478 (N_15478,N_14786,N_14995);
or U15479 (N_15479,N_14690,N_14599);
or U15480 (N_15480,N_14521,N_14594);
nor U15481 (N_15481,N_14950,N_14734);
nor U15482 (N_15482,N_14786,N_14657);
nand U15483 (N_15483,N_14950,N_14581);
nor U15484 (N_15484,N_14883,N_14761);
nor U15485 (N_15485,N_14674,N_14950);
nand U15486 (N_15486,N_14878,N_14646);
and U15487 (N_15487,N_14626,N_14974);
and U15488 (N_15488,N_14555,N_14840);
or U15489 (N_15489,N_14774,N_14731);
and U15490 (N_15490,N_14797,N_14862);
nand U15491 (N_15491,N_14833,N_14553);
nand U15492 (N_15492,N_14831,N_14634);
nand U15493 (N_15493,N_14520,N_14582);
and U15494 (N_15494,N_14829,N_14850);
or U15495 (N_15495,N_14634,N_14811);
or U15496 (N_15496,N_14621,N_14837);
and U15497 (N_15497,N_14758,N_14822);
nand U15498 (N_15498,N_14827,N_14916);
nand U15499 (N_15499,N_14690,N_14692);
and U15500 (N_15500,N_15296,N_15210);
xor U15501 (N_15501,N_15272,N_15417);
nand U15502 (N_15502,N_15455,N_15448);
xnor U15503 (N_15503,N_15392,N_15173);
or U15504 (N_15504,N_15247,N_15015);
nor U15505 (N_15505,N_15342,N_15474);
nor U15506 (N_15506,N_15163,N_15424);
xnor U15507 (N_15507,N_15433,N_15345);
or U15508 (N_15508,N_15029,N_15236);
xor U15509 (N_15509,N_15361,N_15416);
and U15510 (N_15510,N_15081,N_15221);
nor U15511 (N_15511,N_15404,N_15134);
nor U15512 (N_15512,N_15079,N_15051);
and U15513 (N_15513,N_15386,N_15050);
or U15514 (N_15514,N_15205,N_15069);
nor U15515 (N_15515,N_15133,N_15352);
nand U15516 (N_15516,N_15160,N_15248);
and U15517 (N_15517,N_15409,N_15010);
nand U15518 (N_15518,N_15290,N_15240);
nor U15519 (N_15519,N_15207,N_15444);
or U15520 (N_15520,N_15231,N_15040);
or U15521 (N_15521,N_15182,N_15371);
nor U15522 (N_15522,N_15237,N_15279);
and U15523 (N_15523,N_15206,N_15262);
nand U15524 (N_15524,N_15251,N_15265);
nor U15525 (N_15525,N_15143,N_15036);
nor U15526 (N_15526,N_15198,N_15349);
or U15527 (N_15527,N_15309,N_15126);
xor U15528 (N_15528,N_15085,N_15074);
nor U15529 (N_15529,N_15067,N_15288);
xnor U15530 (N_15530,N_15273,N_15360);
nor U15531 (N_15531,N_15225,N_15099);
nor U15532 (N_15532,N_15289,N_15381);
nor U15533 (N_15533,N_15127,N_15440);
or U15534 (N_15534,N_15435,N_15249);
nor U15535 (N_15535,N_15108,N_15261);
and U15536 (N_15536,N_15496,N_15090);
xnor U15537 (N_15537,N_15239,N_15107);
nand U15538 (N_15538,N_15080,N_15009);
nand U15539 (N_15539,N_15006,N_15499);
or U15540 (N_15540,N_15203,N_15354);
nor U15541 (N_15541,N_15431,N_15411);
or U15542 (N_15542,N_15419,N_15170);
and U15543 (N_15543,N_15374,N_15162);
and U15544 (N_15544,N_15252,N_15280);
and U15545 (N_15545,N_15214,N_15175);
nor U15546 (N_15546,N_15087,N_15218);
or U15547 (N_15547,N_15318,N_15246);
nand U15548 (N_15548,N_15344,N_15234);
nor U15549 (N_15549,N_15057,N_15121);
xnor U15550 (N_15550,N_15233,N_15299);
nor U15551 (N_15551,N_15295,N_15105);
nand U15552 (N_15552,N_15412,N_15373);
nand U15553 (N_15553,N_15186,N_15358);
xnor U15554 (N_15554,N_15275,N_15042);
or U15555 (N_15555,N_15021,N_15140);
xnor U15556 (N_15556,N_15364,N_15190);
nor U15557 (N_15557,N_15285,N_15359);
and U15558 (N_15558,N_15227,N_15196);
nor U15559 (N_15559,N_15070,N_15307);
nor U15560 (N_15560,N_15314,N_15202);
nand U15561 (N_15561,N_15426,N_15348);
and U15562 (N_15562,N_15380,N_15365);
nor U15563 (N_15563,N_15018,N_15194);
or U15564 (N_15564,N_15473,N_15319);
nand U15565 (N_15565,N_15430,N_15291);
or U15566 (N_15566,N_15469,N_15331);
and U15567 (N_15567,N_15191,N_15128);
nor U15568 (N_15568,N_15475,N_15058);
or U15569 (N_15569,N_15024,N_15382);
nor U15570 (N_15570,N_15243,N_15420);
nor U15571 (N_15571,N_15068,N_15370);
nand U15572 (N_15572,N_15376,N_15283);
or U15573 (N_15573,N_15076,N_15379);
nand U15574 (N_15574,N_15428,N_15400);
nand U15575 (N_15575,N_15072,N_15315);
xor U15576 (N_15576,N_15393,N_15013);
or U15577 (N_15577,N_15366,N_15346);
xor U15578 (N_15578,N_15122,N_15429);
nor U15579 (N_15579,N_15446,N_15157);
nand U15580 (N_15580,N_15464,N_15481);
nand U15581 (N_15581,N_15350,N_15310);
nor U15582 (N_15582,N_15096,N_15181);
or U15583 (N_15583,N_15383,N_15049);
nor U15584 (N_15584,N_15384,N_15437);
nor U15585 (N_15585,N_15276,N_15211);
nand U15586 (N_15586,N_15438,N_15413);
or U15587 (N_15587,N_15063,N_15490);
nand U15588 (N_15588,N_15297,N_15269);
xor U15589 (N_15589,N_15031,N_15092);
nor U15590 (N_15590,N_15192,N_15375);
or U15591 (N_15591,N_15284,N_15415);
nand U15592 (N_15592,N_15369,N_15495);
nand U15593 (N_15593,N_15399,N_15098);
and U15594 (N_15594,N_15195,N_15264);
or U15595 (N_15595,N_15235,N_15391);
nor U15596 (N_15596,N_15476,N_15007);
xor U15597 (N_15597,N_15467,N_15322);
or U15598 (N_15598,N_15046,N_15165);
or U15599 (N_15599,N_15119,N_15439);
and U15600 (N_15600,N_15078,N_15317);
xnor U15601 (N_15601,N_15266,N_15082);
xnor U15602 (N_15602,N_15089,N_15213);
or U15603 (N_15603,N_15158,N_15253);
xor U15604 (N_15604,N_15362,N_15120);
nor U15605 (N_15605,N_15139,N_15418);
xnor U15606 (N_15606,N_15091,N_15093);
nand U15607 (N_15607,N_15044,N_15056);
nor U15608 (N_15608,N_15001,N_15212);
or U15609 (N_15609,N_15176,N_15189);
nor U15610 (N_15610,N_15335,N_15306);
and U15611 (N_15611,N_15197,N_15101);
or U15612 (N_15612,N_15377,N_15118);
or U15613 (N_15613,N_15449,N_15483);
or U15614 (N_15614,N_15151,N_15489);
xor U15615 (N_15615,N_15298,N_15124);
xor U15616 (N_15616,N_15268,N_15302);
or U15617 (N_15617,N_15325,N_15486);
nand U15618 (N_15618,N_15209,N_15232);
nand U15619 (N_15619,N_15421,N_15408);
nor U15620 (N_15620,N_15405,N_15330);
xnor U15621 (N_15621,N_15385,N_15311);
nor U15622 (N_15622,N_15432,N_15224);
and U15623 (N_15623,N_15368,N_15242);
and U15624 (N_15624,N_15323,N_15442);
xnor U15625 (N_15625,N_15294,N_15077);
and U15626 (N_15626,N_15111,N_15407);
and U15627 (N_15627,N_15187,N_15301);
nor U15628 (N_15628,N_15167,N_15447);
or U15629 (N_15629,N_15328,N_15088);
and U15630 (N_15630,N_15324,N_15329);
and U15631 (N_15631,N_15327,N_15491);
nand U15632 (N_15632,N_15129,N_15071);
nor U15633 (N_15633,N_15456,N_15398);
or U15634 (N_15634,N_15445,N_15263);
nand U15635 (N_15635,N_15028,N_15138);
nand U15636 (N_15636,N_15146,N_15113);
and U15637 (N_15637,N_15131,N_15177);
and U15638 (N_15638,N_15343,N_15367);
nand U15639 (N_15639,N_15389,N_15145);
and U15640 (N_15640,N_15450,N_15274);
nor U15641 (N_15641,N_15460,N_15498);
xor U15642 (N_15642,N_15406,N_15055);
and U15643 (N_15643,N_15023,N_15002);
and U15644 (N_15644,N_15132,N_15075);
or U15645 (N_15645,N_15008,N_15427);
and U15646 (N_15646,N_15403,N_15004);
and U15647 (N_15647,N_15463,N_15178);
or U15648 (N_15648,N_15270,N_15258);
nand U15649 (N_15649,N_15114,N_15397);
xor U15650 (N_15650,N_15104,N_15112);
and U15651 (N_15651,N_15462,N_15492);
and U15652 (N_15652,N_15100,N_15083);
and U15653 (N_15653,N_15395,N_15286);
xor U15654 (N_15654,N_15244,N_15410);
and U15655 (N_15655,N_15052,N_15137);
xnor U15656 (N_15656,N_15012,N_15060);
and U15657 (N_15657,N_15334,N_15135);
nand U15658 (N_15658,N_15480,N_15388);
or U15659 (N_15659,N_15153,N_15461);
or U15660 (N_15660,N_15171,N_15378);
nor U15661 (N_15661,N_15073,N_15230);
or U15662 (N_15662,N_15016,N_15441);
nor U15663 (N_15663,N_15027,N_15312);
xnor U15664 (N_15664,N_15017,N_15065);
nand U15665 (N_15665,N_15179,N_15148);
nor U15666 (N_15666,N_15292,N_15454);
xnor U15667 (N_15667,N_15493,N_15477);
and U15668 (N_15668,N_15147,N_15117);
nand U15669 (N_15669,N_15226,N_15372);
nand U15670 (N_15670,N_15106,N_15141);
and U15671 (N_15671,N_15000,N_15039);
or U15672 (N_15672,N_15183,N_15047);
and U15673 (N_15673,N_15037,N_15387);
nand U15674 (N_15674,N_15156,N_15256);
nor U15675 (N_15675,N_15351,N_15396);
nand U15676 (N_15676,N_15401,N_15340);
nand U15677 (N_15677,N_15423,N_15161);
xor U15678 (N_15678,N_15125,N_15453);
or U15679 (N_15679,N_15038,N_15390);
or U15680 (N_15680,N_15485,N_15219);
xnor U15681 (N_15681,N_15204,N_15086);
and U15682 (N_15682,N_15482,N_15245);
xnor U15683 (N_15683,N_15103,N_15308);
nor U15684 (N_15684,N_15061,N_15497);
nand U15685 (N_15685,N_15144,N_15479);
xnor U15686 (N_15686,N_15287,N_15193);
and U15687 (N_15687,N_15347,N_15130);
or U15688 (N_15688,N_15250,N_15005);
and U15689 (N_15689,N_15355,N_15281);
or U15690 (N_15690,N_15422,N_15303);
xnor U15691 (N_15691,N_15425,N_15316);
or U15692 (N_15692,N_15159,N_15468);
xor U15693 (N_15693,N_15466,N_15166);
and U15694 (N_15694,N_15172,N_15326);
xor U15695 (N_15695,N_15116,N_15267);
and U15696 (N_15696,N_15054,N_15115);
or U15697 (N_15697,N_15053,N_15164);
or U15698 (N_15698,N_15201,N_15142);
nand U15699 (N_15699,N_15020,N_15443);
nor U15700 (N_15700,N_15169,N_15110);
xnor U15701 (N_15701,N_15048,N_15084);
nand U15702 (N_15702,N_15019,N_15045);
nor U15703 (N_15703,N_15095,N_15259);
and U15704 (N_15704,N_15332,N_15282);
or U15705 (N_15705,N_15357,N_15488);
nor U15706 (N_15706,N_15168,N_15152);
xnor U15707 (N_15707,N_15033,N_15305);
nand U15708 (N_15708,N_15338,N_15472);
nand U15709 (N_15709,N_15136,N_15184);
and U15710 (N_15710,N_15313,N_15457);
nand U15711 (N_15711,N_15260,N_15026);
or U15712 (N_15712,N_15223,N_15032);
or U15713 (N_15713,N_15458,N_15321);
nand U15714 (N_15714,N_15222,N_15180);
nor U15715 (N_15715,N_15434,N_15339);
nand U15716 (N_15716,N_15320,N_15255);
and U15717 (N_15717,N_15241,N_15217);
or U15718 (N_15718,N_15011,N_15064);
nand U15719 (N_15719,N_15304,N_15238);
xor U15720 (N_15720,N_15254,N_15097);
or U15721 (N_15721,N_15353,N_15200);
nand U15722 (N_15722,N_15484,N_15478);
and U15723 (N_15723,N_15229,N_15034);
nor U15724 (N_15724,N_15300,N_15333);
nand U15725 (N_15725,N_15356,N_15271);
xor U15726 (N_15726,N_15436,N_15220);
nand U15727 (N_15727,N_15094,N_15337);
xor U15728 (N_15728,N_15394,N_15102);
xor U15729 (N_15729,N_15041,N_15470);
nand U15730 (N_15730,N_15025,N_15059);
and U15731 (N_15731,N_15471,N_15459);
or U15732 (N_15732,N_15452,N_15278);
and U15733 (N_15733,N_15465,N_15257);
or U15734 (N_15734,N_15208,N_15003);
xor U15735 (N_15735,N_15277,N_15066);
or U15736 (N_15736,N_15228,N_15109);
nand U15737 (N_15737,N_15451,N_15494);
xnor U15738 (N_15738,N_15043,N_15174);
nand U15739 (N_15739,N_15022,N_15030);
or U15740 (N_15740,N_15154,N_15199);
and U15741 (N_15741,N_15155,N_15216);
nor U15742 (N_15742,N_15402,N_15150);
nand U15743 (N_15743,N_15293,N_15149);
nand U15744 (N_15744,N_15215,N_15062);
nand U15745 (N_15745,N_15341,N_15336);
nor U15746 (N_15746,N_15123,N_15185);
nor U15747 (N_15747,N_15035,N_15188);
nand U15748 (N_15748,N_15014,N_15487);
or U15749 (N_15749,N_15363,N_15414);
xor U15750 (N_15750,N_15421,N_15447);
or U15751 (N_15751,N_15320,N_15022);
nand U15752 (N_15752,N_15142,N_15442);
and U15753 (N_15753,N_15341,N_15009);
nand U15754 (N_15754,N_15340,N_15252);
and U15755 (N_15755,N_15169,N_15423);
and U15756 (N_15756,N_15141,N_15153);
xor U15757 (N_15757,N_15236,N_15421);
xnor U15758 (N_15758,N_15258,N_15462);
or U15759 (N_15759,N_15264,N_15421);
and U15760 (N_15760,N_15341,N_15029);
nand U15761 (N_15761,N_15136,N_15412);
and U15762 (N_15762,N_15248,N_15349);
or U15763 (N_15763,N_15333,N_15471);
nand U15764 (N_15764,N_15445,N_15115);
nand U15765 (N_15765,N_15456,N_15393);
xnor U15766 (N_15766,N_15016,N_15434);
nor U15767 (N_15767,N_15450,N_15360);
and U15768 (N_15768,N_15039,N_15244);
xnor U15769 (N_15769,N_15005,N_15428);
and U15770 (N_15770,N_15471,N_15479);
nand U15771 (N_15771,N_15453,N_15329);
xor U15772 (N_15772,N_15423,N_15005);
or U15773 (N_15773,N_15276,N_15088);
xnor U15774 (N_15774,N_15040,N_15178);
or U15775 (N_15775,N_15213,N_15242);
nand U15776 (N_15776,N_15072,N_15238);
nand U15777 (N_15777,N_15315,N_15375);
and U15778 (N_15778,N_15117,N_15103);
xor U15779 (N_15779,N_15007,N_15337);
xor U15780 (N_15780,N_15444,N_15299);
nor U15781 (N_15781,N_15435,N_15280);
nand U15782 (N_15782,N_15126,N_15469);
and U15783 (N_15783,N_15181,N_15393);
nand U15784 (N_15784,N_15464,N_15235);
nor U15785 (N_15785,N_15189,N_15487);
or U15786 (N_15786,N_15148,N_15168);
nand U15787 (N_15787,N_15463,N_15128);
xor U15788 (N_15788,N_15318,N_15101);
xnor U15789 (N_15789,N_15342,N_15218);
xnor U15790 (N_15790,N_15401,N_15253);
nor U15791 (N_15791,N_15156,N_15121);
or U15792 (N_15792,N_15370,N_15013);
nand U15793 (N_15793,N_15345,N_15264);
xnor U15794 (N_15794,N_15297,N_15254);
xor U15795 (N_15795,N_15272,N_15339);
and U15796 (N_15796,N_15004,N_15162);
nand U15797 (N_15797,N_15467,N_15192);
xnor U15798 (N_15798,N_15251,N_15387);
or U15799 (N_15799,N_15489,N_15264);
xnor U15800 (N_15800,N_15223,N_15416);
nor U15801 (N_15801,N_15085,N_15098);
nand U15802 (N_15802,N_15251,N_15270);
or U15803 (N_15803,N_15315,N_15154);
nand U15804 (N_15804,N_15016,N_15012);
xnor U15805 (N_15805,N_15414,N_15320);
nor U15806 (N_15806,N_15181,N_15319);
or U15807 (N_15807,N_15193,N_15052);
nor U15808 (N_15808,N_15377,N_15239);
nor U15809 (N_15809,N_15015,N_15397);
and U15810 (N_15810,N_15493,N_15299);
nor U15811 (N_15811,N_15191,N_15295);
and U15812 (N_15812,N_15236,N_15313);
and U15813 (N_15813,N_15016,N_15020);
and U15814 (N_15814,N_15499,N_15227);
nor U15815 (N_15815,N_15493,N_15250);
xnor U15816 (N_15816,N_15400,N_15490);
nor U15817 (N_15817,N_15053,N_15165);
nor U15818 (N_15818,N_15040,N_15043);
and U15819 (N_15819,N_15034,N_15172);
xnor U15820 (N_15820,N_15336,N_15368);
nand U15821 (N_15821,N_15007,N_15289);
xor U15822 (N_15822,N_15194,N_15040);
and U15823 (N_15823,N_15117,N_15351);
or U15824 (N_15824,N_15170,N_15076);
or U15825 (N_15825,N_15198,N_15075);
and U15826 (N_15826,N_15347,N_15104);
xor U15827 (N_15827,N_15042,N_15388);
xor U15828 (N_15828,N_15320,N_15336);
xnor U15829 (N_15829,N_15170,N_15186);
or U15830 (N_15830,N_15419,N_15276);
nand U15831 (N_15831,N_15191,N_15351);
nand U15832 (N_15832,N_15275,N_15230);
xnor U15833 (N_15833,N_15007,N_15306);
xor U15834 (N_15834,N_15352,N_15321);
nand U15835 (N_15835,N_15212,N_15238);
nand U15836 (N_15836,N_15001,N_15049);
and U15837 (N_15837,N_15142,N_15035);
and U15838 (N_15838,N_15123,N_15361);
and U15839 (N_15839,N_15167,N_15182);
or U15840 (N_15840,N_15012,N_15179);
nor U15841 (N_15841,N_15281,N_15017);
nor U15842 (N_15842,N_15215,N_15425);
xnor U15843 (N_15843,N_15302,N_15036);
xor U15844 (N_15844,N_15152,N_15233);
nor U15845 (N_15845,N_15364,N_15237);
nand U15846 (N_15846,N_15087,N_15145);
nor U15847 (N_15847,N_15027,N_15049);
or U15848 (N_15848,N_15006,N_15000);
and U15849 (N_15849,N_15330,N_15223);
xnor U15850 (N_15850,N_15372,N_15486);
xor U15851 (N_15851,N_15047,N_15281);
nand U15852 (N_15852,N_15080,N_15302);
and U15853 (N_15853,N_15342,N_15097);
or U15854 (N_15854,N_15154,N_15172);
nor U15855 (N_15855,N_15273,N_15400);
nor U15856 (N_15856,N_15239,N_15180);
and U15857 (N_15857,N_15074,N_15411);
or U15858 (N_15858,N_15163,N_15357);
xor U15859 (N_15859,N_15096,N_15175);
and U15860 (N_15860,N_15048,N_15485);
nor U15861 (N_15861,N_15450,N_15302);
nand U15862 (N_15862,N_15086,N_15369);
or U15863 (N_15863,N_15024,N_15456);
xor U15864 (N_15864,N_15174,N_15413);
or U15865 (N_15865,N_15155,N_15400);
nand U15866 (N_15866,N_15199,N_15261);
and U15867 (N_15867,N_15352,N_15380);
or U15868 (N_15868,N_15275,N_15174);
and U15869 (N_15869,N_15208,N_15155);
nand U15870 (N_15870,N_15111,N_15161);
nor U15871 (N_15871,N_15130,N_15042);
or U15872 (N_15872,N_15478,N_15260);
nand U15873 (N_15873,N_15189,N_15007);
xor U15874 (N_15874,N_15100,N_15051);
and U15875 (N_15875,N_15225,N_15353);
nand U15876 (N_15876,N_15258,N_15115);
nand U15877 (N_15877,N_15131,N_15453);
and U15878 (N_15878,N_15200,N_15053);
xnor U15879 (N_15879,N_15243,N_15280);
nor U15880 (N_15880,N_15364,N_15158);
and U15881 (N_15881,N_15086,N_15003);
nor U15882 (N_15882,N_15424,N_15293);
or U15883 (N_15883,N_15334,N_15207);
nor U15884 (N_15884,N_15190,N_15102);
or U15885 (N_15885,N_15060,N_15050);
nor U15886 (N_15886,N_15247,N_15434);
or U15887 (N_15887,N_15265,N_15119);
xor U15888 (N_15888,N_15072,N_15457);
nand U15889 (N_15889,N_15333,N_15092);
nor U15890 (N_15890,N_15017,N_15447);
xnor U15891 (N_15891,N_15174,N_15015);
xor U15892 (N_15892,N_15314,N_15171);
or U15893 (N_15893,N_15113,N_15138);
or U15894 (N_15894,N_15070,N_15316);
and U15895 (N_15895,N_15089,N_15027);
xnor U15896 (N_15896,N_15023,N_15169);
nand U15897 (N_15897,N_15487,N_15171);
nor U15898 (N_15898,N_15369,N_15139);
xor U15899 (N_15899,N_15368,N_15494);
and U15900 (N_15900,N_15445,N_15371);
xnor U15901 (N_15901,N_15449,N_15319);
or U15902 (N_15902,N_15185,N_15352);
nand U15903 (N_15903,N_15220,N_15379);
or U15904 (N_15904,N_15350,N_15413);
nor U15905 (N_15905,N_15069,N_15023);
or U15906 (N_15906,N_15394,N_15042);
or U15907 (N_15907,N_15167,N_15352);
and U15908 (N_15908,N_15078,N_15022);
or U15909 (N_15909,N_15458,N_15245);
xor U15910 (N_15910,N_15140,N_15190);
nand U15911 (N_15911,N_15054,N_15171);
nor U15912 (N_15912,N_15420,N_15460);
xnor U15913 (N_15913,N_15248,N_15126);
or U15914 (N_15914,N_15015,N_15374);
xnor U15915 (N_15915,N_15413,N_15100);
nand U15916 (N_15916,N_15415,N_15444);
and U15917 (N_15917,N_15480,N_15496);
nor U15918 (N_15918,N_15022,N_15249);
nor U15919 (N_15919,N_15077,N_15375);
and U15920 (N_15920,N_15139,N_15215);
or U15921 (N_15921,N_15328,N_15360);
xor U15922 (N_15922,N_15359,N_15360);
and U15923 (N_15923,N_15097,N_15061);
nand U15924 (N_15924,N_15251,N_15451);
xnor U15925 (N_15925,N_15007,N_15039);
nand U15926 (N_15926,N_15049,N_15495);
nand U15927 (N_15927,N_15189,N_15451);
and U15928 (N_15928,N_15418,N_15297);
nor U15929 (N_15929,N_15190,N_15297);
or U15930 (N_15930,N_15377,N_15102);
xor U15931 (N_15931,N_15129,N_15346);
or U15932 (N_15932,N_15091,N_15212);
nor U15933 (N_15933,N_15137,N_15280);
nor U15934 (N_15934,N_15350,N_15003);
and U15935 (N_15935,N_15494,N_15114);
nor U15936 (N_15936,N_15005,N_15438);
xnor U15937 (N_15937,N_15127,N_15425);
nand U15938 (N_15938,N_15370,N_15427);
xnor U15939 (N_15939,N_15166,N_15332);
and U15940 (N_15940,N_15174,N_15262);
nor U15941 (N_15941,N_15078,N_15297);
nand U15942 (N_15942,N_15306,N_15295);
nor U15943 (N_15943,N_15397,N_15324);
or U15944 (N_15944,N_15393,N_15380);
nand U15945 (N_15945,N_15201,N_15455);
and U15946 (N_15946,N_15498,N_15180);
xnor U15947 (N_15947,N_15270,N_15007);
or U15948 (N_15948,N_15304,N_15234);
xor U15949 (N_15949,N_15042,N_15389);
xor U15950 (N_15950,N_15131,N_15208);
nor U15951 (N_15951,N_15142,N_15204);
or U15952 (N_15952,N_15190,N_15432);
xnor U15953 (N_15953,N_15373,N_15470);
xnor U15954 (N_15954,N_15275,N_15329);
and U15955 (N_15955,N_15389,N_15452);
or U15956 (N_15956,N_15366,N_15192);
or U15957 (N_15957,N_15483,N_15469);
nand U15958 (N_15958,N_15238,N_15101);
nand U15959 (N_15959,N_15034,N_15079);
nor U15960 (N_15960,N_15057,N_15309);
nor U15961 (N_15961,N_15055,N_15284);
xor U15962 (N_15962,N_15095,N_15484);
and U15963 (N_15963,N_15196,N_15454);
xor U15964 (N_15964,N_15130,N_15372);
and U15965 (N_15965,N_15067,N_15478);
nand U15966 (N_15966,N_15388,N_15111);
xor U15967 (N_15967,N_15205,N_15150);
and U15968 (N_15968,N_15061,N_15227);
and U15969 (N_15969,N_15476,N_15330);
or U15970 (N_15970,N_15073,N_15289);
xnor U15971 (N_15971,N_15433,N_15375);
and U15972 (N_15972,N_15036,N_15492);
or U15973 (N_15973,N_15428,N_15346);
xnor U15974 (N_15974,N_15220,N_15021);
or U15975 (N_15975,N_15335,N_15487);
nand U15976 (N_15976,N_15213,N_15048);
and U15977 (N_15977,N_15099,N_15156);
nand U15978 (N_15978,N_15286,N_15274);
nand U15979 (N_15979,N_15272,N_15302);
nand U15980 (N_15980,N_15375,N_15200);
or U15981 (N_15981,N_15102,N_15410);
nand U15982 (N_15982,N_15001,N_15054);
nand U15983 (N_15983,N_15395,N_15002);
or U15984 (N_15984,N_15207,N_15381);
and U15985 (N_15985,N_15210,N_15359);
and U15986 (N_15986,N_15167,N_15027);
and U15987 (N_15987,N_15465,N_15309);
or U15988 (N_15988,N_15088,N_15188);
nand U15989 (N_15989,N_15317,N_15266);
nand U15990 (N_15990,N_15025,N_15176);
xnor U15991 (N_15991,N_15095,N_15180);
nand U15992 (N_15992,N_15318,N_15085);
xnor U15993 (N_15993,N_15157,N_15009);
or U15994 (N_15994,N_15389,N_15118);
nand U15995 (N_15995,N_15301,N_15476);
nand U15996 (N_15996,N_15339,N_15145);
nand U15997 (N_15997,N_15203,N_15353);
or U15998 (N_15998,N_15048,N_15407);
xor U15999 (N_15999,N_15154,N_15439);
xor U16000 (N_16000,N_15609,N_15633);
and U16001 (N_16001,N_15900,N_15839);
xnor U16002 (N_16002,N_15576,N_15654);
nand U16003 (N_16003,N_15554,N_15750);
nand U16004 (N_16004,N_15563,N_15786);
nand U16005 (N_16005,N_15629,N_15909);
or U16006 (N_16006,N_15984,N_15624);
nand U16007 (N_16007,N_15587,N_15907);
nand U16008 (N_16008,N_15876,N_15809);
and U16009 (N_16009,N_15953,N_15598);
nor U16010 (N_16010,N_15664,N_15880);
and U16011 (N_16011,N_15978,N_15770);
nor U16012 (N_16012,N_15502,N_15673);
or U16013 (N_16013,N_15627,N_15704);
nand U16014 (N_16014,N_15542,N_15949);
and U16015 (N_16015,N_15814,N_15510);
xor U16016 (N_16016,N_15591,N_15776);
nor U16017 (N_16017,N_15637,N_15751);
or U16018 (N_16018,N_15929,N_15675);
nand U16019 (N_16019,N_15611,N_15742);
xnor U16020 (N_16020,N_15891,N_15877);
xor U16021 (N_16021,N_15834,N_15976);
or U16022 (N_16022,N_15560,N_15529);
or U16023 (N_16023,N_15740,N_15996);
xor U16024 (N_16024,N_15808,N_15728);
nor U16025 (N_16025,N_15551,N_15940);
and U16026 (N_16026,N_15754,N_15552);
or U16027 (N_16027,N_15562,N_15706);
nor U16028 (N_16028,N_15515,N_15570);
or U16029 (N_16029,N_15896,N_15720);
nor U16030 (N_16030,N_15730,N_15693);
nand U16031 (N_16031,N_15854,N_15852);
and U16032 (N_16032,N_15581,N_15614);
and U16033 (N_16033,N_15545,N_15979);
nand U16034 (N_16034,N_15606,N_15749);
nand U16035 (N_16035,N_15688,N_15862);
xor U16036 (N_16036,N_15710,N_15884);
and U16037 (N_16037,N_15847,N_15927);
or U16038 (N_16038,N_15861,N_15864);
nand U16039 (N_16039,N_15696,N_15731);
and U16040 (N_16040,N_15930,N_15500);
nor U16041 (N_16041,N_15863,N_15796);
or U16042 (N_16042,N_15868,N_15523);
nor U16043 (N_16043,N_15649,N_15842);
nand U16044 (N_16044,N_15859,N_15989);
xnor U16045 (N_16045,N_15805,N_15885);
nor U16046 (N_16046,N_15753,N_15518);
and U16047 (N_16047,N_15821,N_15780);
nor U16048 (N_16048,N_15958,N_15871);
and U16049 (N_16049,N_15916,N_15765);
xor U16050 (N_16050,N_15830,N_15875);
or U16051 (N_16051,N_15747,N_15759);
nor U16052 (N_16052,N_15746,N_15707);
and U16053 (N_16053,N_15959,N_15748);
or U16054 (N_16054,N_15509,N_15961);
or U16055 (N_16055,N_15666,N_15715);
or U16056 (N_16056,N_15535,N_15716);
nand U16057 (N_16057,N_15695,N_15744);
and U16058 (N_16058,N_15677,N_15787);
nor U16059 (N_16059,N_15691,N_15617);
xnor U16060 (N_16060,N_15967,N_15956);
nand U16061 (N_16061,N_15711,N_15572);
or U16062 (N_16062,N_15922,N_15840);
nor U16063 (N_16063,N_15950,N_15889);
or U16064 (N_16064,N_15827,N_15911);
and U16065 (N_16065,N_15969,N_15680);
and U16066 (N_16066,N_15504,N_15792);
nand U16067 (N_16067,N_15588,N_15766);
xnor U16068 (N_16068,N_15768,N_15771);
nand U16069 (N_16069,N_15812,N_15632);
nor U16070 (N_16070,N_15816,N_15619);
nand U16071 (N_16071,N_15557,N_15925);
or U16072 (N_16072,N_15685,N_15732);
nor U16073 (N_16073,N_15987,N_15917);
or U16074 (N_16074,N_15872,N_15756);
nor U16075 (N_16075,N_15952,N_15575);
and U16076 (N_16076,N_15908,N_15698);
nand U16077 (N_16077,N_15526,N_15752);
nand U16078 (N_16078,N_15628,N_15760);
xnor U16079 (N_16079,N_15806,N_15733);
nand U16080 (N_16080,N_15586,N_15717);
or U16081 (N_16081,N_15519,N_15874);
xnor U16082 (N_16082,N_15610,N_15517);
nor U16083 (N_16083,N_15574,N_15714);
and U16084 (N_16084,N_15726,N_15601);
or U16085 (N_16085,N_15946,N_15555);
or U16086 (N_16086,N_15886,N_15667);
nor U16087 (N_16087,N_15638,N_15836);
nor U16088 (N_16088,N_15799,N_15789);
nand U16089 (N_16089,N_15650,N_15681);
nor U16090 (N_16090,N_15924,N_15603);
nor U16091 (N_16091,N_15923,N_15790);
or U16092 (N_16092,N_15826,N_15920);
nand U16093 (N_16093,N_15735,N_15797);
xor U16094 (N_16094,N_15605,N_15738);
xor U16095 (N_16095,N_15699,N_15968);
and U16096 (N_16096,N_15912,N_15538);
nor U16097 (N_16097,N_15589,N_15620);
and U16098 (N_16098,N_15561,N_15604);
xor U16099 (N_16099,N_15837,N_15951);
nor U16100 (N_16100,N_15697,N_15965);
and U16101 (N_16101,N_15536,N_15833);
and U16102 (N_16102,N_15692,N_15762);
xor U16103 (N_16103,N_15646,N_15533);
and U16104 (N_16104,N_15943,N_15807);
or U16105 (N_16105,N_15682,N_15995);
or U16106 (N_16106,N_15516,N_15931);
nor U16107 (N_16107,N_15781,N_15981);
nor U16108 (N_16108,N_15919,N_15729);
nor U16109 (N_16109,N_15564,N_15937);
nand U16110 (N_16110,N_15530,N_15763);
nand U16111 (N_16111,N_15988,N_15823);
xnor U16112 (N_16112,N_15577,N_15566);
and U16113 (N_16113,N_15703,N_15773);
or U16114 (N_16114,N_15879,N_15855);
and U16115 (N_16115,N_15725,N_15843);
xor U16116 (N_16116,N_15565,N_15736);
xor U16117 (N_16117,N_15737,N_15921);
nor U16118 (N_16118,N_15901,N_15926);
and U16119 (N_16119,N_15625,N_15985);
and U16120 (N_16120,N_15878,N_15835);
xnor U16121 (N_16121,N_15801,N_15507);
nor U16122 (N_16122,N_15804,N_15665);
nor U16123 (N_16123,N_15743,N_15914);
nand U16124 (N_16124,N_15913,N_15870);
nor U16125 (N_16125,N_15903,N_15819);
or U16126 (N_16126,N_15669,N_15980);
and U16127 (N_16127,N_15838,N_15592);
nor U16128 (N_16128,N_15970,N_15676);
xor U16129 (N_16129,N_15569,N_15644);
xor U16130 (N_16130,N_15774,N_15986);
xor U16131 (N_16131,N_15656,N_15895);
nand U16132 (N_16132,N_15971,N_15820);
xor U16133 (N_16133,N_15899,N_15775);
and U16134 (N_16134,N_15558,N_15534);
nor U16135 (N_16135,N_15932,N_15898);
nand U16136 (N_16136,N_15573,N_15613);
and U16137 (N_16137,N_15977,N_15708);
nor U16138 (N_16138,N_15593,N_15630);
xor U16139 (N_16139,N_15544,N_15945);
nand U16140 (N_16140,N_15894,N_15689);
nand U16141 (N_16141,N_15778,N_15522);
nor U16142 (N_16142,N_15849,N_15687);
nor U16143 (N_16143,N_15853,N_15992);
or U16144 (N_16144,N_15905,N_15800);
nor U16145 (N_16145,N_15585,N_15767);
or U16146 (N_16146,N_15674,N_15739);
nor U16147 (N_16147,N_15506,N_15777);
nand U16148 (N_16148,N_15802,N_15648);
nor U16149 (N_16149,N_15531,N_15998);
nor U16150 (N_16150,N_15700,N_15634);
or U16151 (N_16151,N_15793,N_15663);
or U16152 (N_16152,N_15712,N_15865);
xor U16153 (N_16153,N_15636,N_15549);
nor U16154 (N_16154,N_15954,N_15660);
xnor U16155 (N_16155,N_15722,N_15906);
xor U16156 (N_16156,N_15813,N_15596);
and U16157 (N_16157,N_15694,N_15653);
nand U16158 (N_16158,N_15873,N_15524);
and U16159 (N_16159,N_15626,N_15607);
and U16160 (N_16160,N_15990,N_15643);
or U16161 (N_16161,N_15684,N_15546);
or U16162 (N_16162,N_15761,N_15672);
nand U16163 (N_16163,N_15599,N_15622);
nor U16164 (N_16164,N_15658,N_15709);
nor U16165 (N_16165,N_15825,N_15915);
nand U16166 (N_16166,N_15782,N_15616);
and U16167 (N_16167,N_15845,N_15982);
nor U16168 (N_16168,N_15822,N_15817);
xnor U16169 (N_16169,N_15942,N_15783);
nand U16170 (N_16170,N_15857,N_15850);
and U16171 (N_16171,N_15661,N_15897);
nand U16172 (N_16172,N_15727,N_15721);
and U16173 (N_16173,N_15974,N_15947);
nor U16174 (N_16174,N_15851,N_15784);
nand U16175 (N_16175,N_15972,N_15584);
nor U16176 (N_16176,N_15595,N_15505);
nand U16177 (N_16177,N_15764,N_15964);
nand U16178 (N_16178,N_15795,N_15983);
xnor U16179 (N_16179,N_15662,N_15893);
nand U16180 (N_16180,N_15939,N_15824);
or U16181 (N_16181,N_15679,N_15831);
xnor U16182 (N_16182,N_15844,N_15848);
and U16183 (N_16183,N_15973,N_15975);
xor U16184 (N_16184,N_15892,N_15828);
xor U16185 (N_16185,N_15623,N_15705);
xnor U16186 (N_16186,N_15723,N_15955);
nand U16187 (N_16187,N_15568,N_15772);
nand U16188 (N_16188,N_15579,N_15553);
nand U16189 (N_16189,N_15655,N_15541);
xnor U16190 (N_16190,N_15818,N_15659);
and U16191 (N_16191,N_15532,N_15769);
and U16192 (N_16192,N_15639,N_15527);
and U16193 (N_16193,N_15928,N_15741);
and U16194 (N_16194,N_15513,N_15548);
and U16195 (N_16195,N_15933,N_15668);
nor U16196 (N_16196,N_15944,N_15935);
nor U16197 (N_16197,N_15938,N_15652);
and U16198 (N_16198,N_15794,N_15583);
nor U16199 (N_16199,N_15631,N_15520);
nand U16200 (N_16200,N_15960,N_15671);
or U16201 (N_16201,N_15883,N_15811);
nand U16202 (N_16202,N_15580,N_15860);
xnor U16203 (N_16203,N_15963,N_15934);
nor U16204 (N_16204,N_15621,N_15597);
nand U16205 (N_16205,N_15642,N_15866);
xnor U16206 (N_16206,N_15719,N_15521);
nor U16207 (N_16207,N_15918,N_15525);
and U16208 (N_16208,N_15966,N_15724);
xor U16209 (N_16209,N_15501,N_15645);
or U16210 (N_16210,N_15999,N_15713);
xnor U16211 (N_16211,N_15991,N_15635);
or U16212 (N_16212,N_15612,N_15734);
nor U16213 (N_16213,N_15702,N_15791);
and U16214 (N_16214,N_15858,N_15647);
or U16215 (N_16215,N_15758,N_15641);
or U16216 (N_16216,N_15571,N_15832);
and U16217 (N_16217,N_15785,N_15602);
and U16218 (N_16218,N_15514,N_15547);
and U16219 (N_16219,N_15757,N_15718);
nand U16220 (N_16220,N_15888,N_15550);
xnor U16221 (N_16221,N_15678,N_15882);
nor U16222 (N_16222,N_15618,N_15528);
and U16223 (N_16223,N_15511,N_15829);
nor U16224 (N_16224,N_15537,N_15902);
or U16225 (N_16225,N_15890,N_15512);
nand U16226 (N_16226,N_15600,N_15904);
and U16227 (N_16227,N_15701,N_15810);
nand U16228 (N_16228,N_15543,N_15657);
and U16229 (N_16229,N_15841,N_15887);
nand U16230 (N_16230,N_15941,N_15683);
xor U16231 (N_16231,N_15539,N_15867);
xor U16232 (N_16232,N_15578,N_15615);
nand U16233 (N_16233,N_15856,N_15590);
nand U16234 (N_16234,N_15567,N_15846);
nand U16235 (N_16235,N_15910,N_15582);
nand U16236 (N_16236,N_15608,N_15503);
nor U16237 (N_16237,N_15957,N_15815);
and U16238 (N_16238,N_15640,N_15803);
xnor U16239 (N_16239,N_15779,N_15540);
xnor U16240 (N_16240,N_15869,N_15994);
xnor U16241 (N_16241,N_15690,N_15508);
xor U16242 (N_16242,N_15948,N_15788);
xor U16243 (N_16243,N_15556,N_15936);
xor U16244 (N_16244,N_15755,N_15997);
nand U16245 (N_16245,N_15798,N_15559);
xnor U16246 (N_16246,N_15881,N_15962);
or U16247 (N_16247,N_15594,N_15686);
and U16248 (N_16248,N_15651,N_15745);
or U16249 (N_16249,N_15670,N_15993);
nand U16250 (N_16250,N_15903,N_15536);
or U16251 (N_16251,N_15609,N_15931);
nand U16252 (N_16252,N_15631,N_15873);
nor U16253 (N_16253,N_15874,N_15668);
and U16254 (N_16254,N_15582,N_15756);
and U16255 (N_16255,N_15737,N_15734);
xor U16256 (N_16256,N_15724,N_15530);
and U16257 (N_16257,N_15693,N_15624);
nor U16258 (N_16258,N_15598,N_15775);
nor U16259 (N_16259,N_15727,N_15557);
or U16260 (N_16260,N_15594,N_15892);
nand U16261 (N_16261,N_15781,N_15567);
xor U16262 (N_16262,N_15816,N_15678);
xnor U16263 (N_16263,N_15712,N_15632);
xor U16264 (N_16264,N_15844,N_15701);
nor U16265 (N_16265,N_15702,N_15947);
or U16266 (N_16266,N_15754,N_15663);
nor U16267 (N_16267,N_15509,N_15891);
xor U16268 (N_16268,N_15538,N_15913);
nand U16269 (N_16269,N_15547,N_15623);
nand U16270 (N_16270,N_15848,N_15863);
nand U16271 (N_16271,N_15622,N_15886);
or U16272 (N_16272,N_15734,N_15765);
and U16273 (N_16273,N_15628,N_15972);
nand U16274 (N_16274,N_15951,N_15553);
and U16275 (N_16275,N_15814,N_15756);
nor U16276 (N_16276,N_15962,N_15678);
and U16277 (N_16277,N_15576,N_15823);
or U16278 (N_16278,N_15641,N_15769);
or U16279 (N_16279,N_15572,N_15504);
nor U16280 (N_16280,N_15865,N_15663);
nand U16281 (N_16281,N_15579,N_15842);
xnor U16282 (N_16282,N_15589,N_15712);
nand U16283 (N_16283,N_15503,N_15734);
nor U16284 (N_16284,N_15783,N_15633);
xor U16285 (N_16285,N_15664,N_15908);
nor U16286 (N_16286,N_15772,N_15901);
xnor U16287 (N_16287,N_15827,N_15599);
or U16288 (N_16288,N_15537,N_15680);
xor U16289 (N_16289,N_15633,N_15917);
xor U16290 (N_16290,N_15784,N_15823);
nor U16291 (N_16291,N_15652,N_15961);
xnor U16292 (N_16292,N_15936,N_15609);
and U16293 (N_16293,N_15660,N_15900);
nor U16294 (N_16294,N_15820,N_15604);
or U16295 (N_16295,N_15556,N_15875);
or U16296 (N_16296,N_15921,N_15500);
and U16297 (N_16297,N_15772,N_15954);
xor U16298 (N_16298,N_15802,N_15743);
and U16299 (N_16299,N_15584,N_15632);
xor U16300 (N_16300,N_15581,N_15560);
or U16301 (N_16301,N_15992,N_15867);
nor U16302 (N_16302,N_15970,N_15973);
or U16303 (N_16303,N_15655,N_15727);
xor U16304 (N_16304,N_15859,N_15548);
nor U16305 (N_16305,N_15540,N_15602);
xnor U16306 (N_16306,N_15632,N_15656);
or U16307 (N_16307,N_15863,N_15820);
xnor U16308 (N_16308,N_15787,N_15937);
and U16309 (N_16309,N_15947,N_15859);
or U16310 (N_16310,N_15943,N_15815);
nand U16311 (N_16311,N_15906,N_15894);
and U16312 (N_16312,N_15631,N_15990);
and U16313 (N_16313,N_15619,N_15525);
nor U16314 (N_16314,N_15645,N_15602);
or U16315 (N_16315,N_15590,N_15571);
nor U16316 (N_16316,N_15760,N_15797);
and U16317 (N_16317,N_15637,N_15636);
or U16318 (N_16318,N_15585,N_15729);
or U16319 (N_16319,N_15937,N_15516);
nand U16320 (N_16320,N_15961,N_15828);
nand U16321 (N_16321,N_15889,N_15998);
nor U16322 (N_16322,N_15872,N_15997);
xor U16323 (N_16323,N_15566,N_15922);
and U16324 (N_16324,N_15906,N_15794);
or U16325 (N_16325,N_15681,N_15680);
nor U16326 (N_16326,N_15847,N_15797);
xor U16327 (N_16327,N_15647,N_15729);
xnor U16328 (N_16328,N_15702,N_15768);
or U16329 (N_16329,N_15859,N_15880);
xor U16330 (N_16330,N_15501,N_15955);
nor U16331 (N_16331,N_15672,N_15920);
nor U16332 (N_16332,N_15860,N_15933);
nor U16333 (N_16333,N_15855,N_15637);
nand U16334 (N_16334,N_15880,N_15963);
nor U16335 (N_16335,N_15703,N_15976);
nor U16336 (N_16336,N_15881,N_15597);
xor U16337 (N_16337,N_15980,N_15982);
nand U16338 (N_16338,N_15641,N_15617);
nor U16339 (N_16339,N_15630,N_15950);
nor U16340 (N_16340,N_15662,N_15871);
nand U16341 (N_16341,N_15873,N_15531);
and U16342 (N_16342,N_15620,N_15676);
or U16343 (N_16343,N_15874,N_15878);
nor U16344 (N_16344,N_15736,N_15940);
nor U16345 (N_16345,N_15629,N_15795);
and U16346 (N_16346,N_15942,N_15872);
and U16347 (N_16347,N_15582,N_15639);
or U16348 (N_16348,N_15532,N_15759);
nand U16349 (N_16349,N_15749,N_15804);
nand U16350 (N_16350,N_15757,N_15579);
nand U16351 (N_16351,N_15742,N_15573);
xnor U16352 (N_16352,N_15718,N_15526);
nor U16353 (N_16353,N_15826,N_15541);
or U16354 (N_16354,N_15802,N_15967);
xnor U16355 (N_16355,N_15573,N_15529);
nand U16356 (N_16356,N_15542,N_15738);
xor U16357 (N_16357,N_15654,N_15735);
xnor U16358 (N_16358,N_15919,N_15591);
nor U16359 (N_16359,N_15636,N_15970);
and U16360 (N_16360,N_15627,N_15914);
xor U16361 (N_16361,N_15611,N_15691);
or U16362 (N_16362,N_15683,N_15538);
or U16363 (N_16363,N_15729,N_15931);
nor U16364 (N_16364,N_15790,N_15700);
nor U16365 (N_16365,N_15553,N_15530);
nor U16366 (N_16366,N_15876,N_15728);
xnor U16367 (N_16367,N_15693,N_15738);
nand U16368 (N_16368,N_15600,N_15728);
nand U16369 (N_16369,N_15553,N_15835);
xor U16370 (N_16370,N_15941,N_15598);
nor U16371 (N_16371,N_15751,N_15847);
nand U16372 (N_16372,N_15715,N_15904);
or U16373 (N_16373,N_15802,N_15663);
or U16374 (N_16374,N_15779,N_15642);
xor U16375 (N_16375,N_15909,N_15875);
and U16376 (N_16376,N_15510,N_15535);
or U16377 (N_16377,N_15731,N_15609);
nor U16378 (N_16378,N_15558,N_15514);
nor U16379 (N_16379,N_15505,N_15619);
nor U16380 (N_16380,N_15560,N_15930);
nor U16381 (N_16381,N_15724,N_15821);
xor U16382 (N_16382,N_15967,N_15594);
or U16383 (N_16383,N_15853,N_15815);
and U16384 (N_16384,N_15750,N_15767);
or U16385 (N_16385,N_15959,N_15905);
nand U16386 (N_16386,N_15611,N_15816);
xor U16387 (N_16387,N_15980,N_15515);
and U16388 (N_16388,N_15976,N_15766);
nand U16389 (N_16389,N_15890,N_15630);
nand U16390 (N_16390,N_15768,N_15753);
nor U16391 (N_16391,N_15955,N_15865);
nor U16392 (N_16392,N_15524,N_15705);
nor U16393 (N_16393,N_15996,N_15984);
or U16394 (N_16394,N_15892,N_15597);
nand U16395 (N_16395,N_15861,N_15693);
nor U16396 (N_16396,N_15888,N_15584);
nand U16397 (N_16397,N_15535,N_15655);
or U16398 (N_16398,N_15629,N_15761);
or U16399 (N_16399,N_15706,N_15969);
and U16400 (N_16400,N_15804,N_15510);
nand U16401 (N_16401,N_15968,N_15938);
or U16402 (N_16402,N_15907,N_15992);
and U16403 (N_16403,N_15950,N_15677);
nor U16404 (N_16404,N_15847,N_15627);
nand U16405 (N_16405,N_15710,N_15866);
nand U16406 (N_16406,N_15727,N_15862);
xnor U16407 (N_16407,N_15746,N_15699);
nor U16408 (N_16408,N_15799,N_15533);
xnor U16409 (N_16409,N_15827,N_15549);
and U16410 (N_16410,N_15763,N_15873);
and U16411 (N_16411,N_15602,N_15663);
and U16412 (N_16412,N_15698,N_15599);
nor U16413 (N_16413,N_15987,N_15760);
nor U16414 (N_16414,N_15913,N_15975);
and U16415 (N_16415,N_15889,N_15944);
nor U16416 (N_16416,N_15871,N_15818);
or U16417 (N_16417,N_15583,N_15983);
nor U16418 (N_16418,N_15722,N_15647);
or U16419 (N_16419,N_15503,N_15670);
and U16420 (N_16420,N_15553,N_15899);
nand U16421 (N_16421,N_15850,N_15997);
or U16422 (N_16422,N_15852,N_15950);
nand U16423 (N_16423,N_15826,N_15825);
or U16424 (N_16424,N_15845,N_15587);
xnor U16425 (N_16425,N_15726,N_15747);
nand U16426 (N_16426,N_15618,N_15578);
nor U16427 (N_16427,N_15628,N_15700);
xnor U16428 (N_16428,N_15886,N_15745);
nor U16429 (N_16429,N_15682,N_15603);
or U16430 (N_16430,N_15998,N_15548);
and U16431 (N_16431,N_15674,N_15910);
and U16432 (N_16432,N_15835,N_15780);
nand U16433 (N_16433,N_15674,N_15908);
nand U16434 (N_16434,N_15779,N_15880);
xor U16435 (N_16435,N_15801,N_15623);
xor U16436 (N_16436,N_15898,N_15974);
and U16437 (N_16437,N_15620,N_15771);
nand U16438 (N_16438,N_15993,N_15690);
or U16439 (N_16439,N_15843,N_15835);
and U16440 (N_16440,N_15770,N_15550);
and U16441 (N_16441,N_15640,N_15968);
nand U16442 (N_16442,N_15622,N_15905);
nand U16443 (N_16443,N_15704,N_15755);
nor U16444 (N_16444,N_15711,N_15896);
nand U16445 (N_16445,N_15932,N_15894);
xor U16446 (N_16446,N_15957,N_15990);
xor U16447 (N_16447,N_15666,N_15706);
nand U16448 (N_16448,N_15765,N_15775);
and U16449 (N_16449,N_15903,N_15845);
or U16450 (N_16450,N_15956,N_15772);
and U16451 (N_16451,N_15889,N_15783);
xnor U16452 (N_16452,N_15955,N_15545);
xnor U16453 (N_16453,N_15887,N_15700);
nor U16454 (N_16454,N_15925,N_15552);
and U16455 (N_16455,N_15571,N_15967);
nor U16456 (N_16456,N_15741,N_15935);
or U16457 (N_16457,N_15545,N_15735);
nand U16458 (N_16458,N_15823,N_15796);
nand U16459 (N_16459,N_15876,N_15597);
nor U16460 (N_16460,N_15888,N_15904);
or U16461 (N_16461,N_15902,N_15607);
nand U16462 (N_16462,N_15584,N_15758);
nor U16463 (N_16463,N_15857,N_15731);
or U16464 (N_16464,N_15601,N_15591);
nand U16465 (N_16465,N_15595,N_15585);
or U16466 (N_16466,N_15775,N_15865);
nor U16467 (N_16467,N_15544,N_15518);
nand U16468 (N_16468,N_15845,N_15960);
and U16469 (N_16469,N_15522,N_15752);
xor U16470 (N_16470,N_15847,N_15835);
nor U16471 (N_16471,N_15658,N_15712);
and U16472 (N_16472,N_15937,N_15975);
xnor U16473 (N_16473,N_15686,N_15777);
nor U16474 (N_16474,N_15606,N_15561);
nor U16475 (N_16475,N_15709,N_15639);
nor U16476 (N_16476,N_15630,N_15941);
and U16477 (N_16477,N_15868,N_15781);
xnor U16478 (N_16478,N_15872,N_15757);
or U16479 (N_16479,N_15549,N_15784);
xor U16480 (N_16480,N_15830,N_15682);
nand U16481 (N_16481,N_15589,N_15937);
and U16482 (N_16482,N_15628,N_15818);
or U16483 (N_16483,N_15810,N_15639);
nor U16484 (N_16484,N_15862,N_15595);
nor U16485 (N_16485,N_15811,N_15697);
xnor U16486 (N_16486,N_15560,N_15660);
xor U16487 (N_16487,N_15518,N_15832);
or U16488 (N_16488,N_15732,N_15844);
xor U16489 (N_16489,N_15754,N_15599);
and U16490 (N_16490,N_15616,N_15868);
xnor U16491 (N_16491,N_15778,N_15695);
nor U16492 (N_16492,N_15652,N_15808);
or U16493 (N_16493,N_15878,N_15574);
nor U16494 (N_16494,N_15826,N_15909);
nand U16495 (N_16495,N_15611,N_15799);
nand U16496 (N_16496,N_15549,N_15548);
nand U16497 (N_16497,N_15814,N_15530);
nor U16498 (N_16498,N_15909,N_15703);
and U16499 (N_16499,N_15717,N_15850);
xnor U16500 (N_16500,N_16477,N_16143);
nor U16501 (N_16501,N_16000,N_16237);
xnor U16502 (N_16502,N_16362,N_16469);
or U16503 (N_16503,N_16276,N_16031);
xor U16504 (N_16504,N_16486,N_16281);
and U16505 (N_16505,N_16400,N_16206);
xnor U16506 (N_16506,N_16351,N_16267);
nand U16507 (N_16507,N_16340,N_16204);
nor U16508 (N_16508,N_16091,N_16301);
and U16509 (N_16509,N_16138,N_16214);
or U16510 (N_16510,N_16103,N_16483);
nand U16511 (N_16511,N_16134,N_16336);
and U16512 (N_16512,N_16449,N_16024);
and U16513 (N_16513,N_16332,N_16217);
nor U16514 (N_16514,N_16361,N_16186);
and U16515 (N_16515,N_16093,N_16314);
and U16516 (N_16516,N_16233,N_16155);
or U16517 (N_16517,N_16323,N_16209);
or U16518 (N_16518,N_16460,N_16485);
xor U16519 (N_16519,N_16264,N_16028);
nor U16520 (N_16520,N_16411,N_16159);
xor U16521 (N_16521,N_16380,N_16303);
xor U16522 (N_16522,N_16350,N_16006);
and U16523 (N_16523,N_16354,N_16016);
xnor U16524 (N_16524,N_16240,N_16200);
nand U16525 (N_16525,N_16042,N_16359);
or U16526 (N_16526,N_16439,N_16215);
xnor U16527 (N_16527,N_16117,N_16320);
or U16528 (N_16528,N_16476,N_16481);
nor U16529 (N_16529,N_16269,N_16472);
or U16530 (N_16530,N_16297,N_16199);
and U16531 (N_16531,N_16089,N_16106);
nand U16532 (N_16532,N_16262,N_16223);
and U16533 (N_16533,N_16168,N_16410);
or U16534 (N_16534,N_16198,N_16007);
nand U16535 (N_16535,N_16309,N_16422);
nor U16536 (N_16536,N_16333,N_16498);
xor U16537 (N_16537,N_16337,N_16271);
nand U16538 (N_16538,N_16195,N_16428);
and U16539 (N_16539,N_16254,N_16107);
nand U16540 (N_16540,N_16265,N_16034);
or U16541 (N_16541,N_16352,N_16394);
nand U16542 (N_16542,N_16412,N_16471);
xor U16543 (N_16543,N_16136,N_16375);
nor U16544 (N_16544,N_16225,N_16196);
nor U16545 (N_16545,N_16389,N_16242);
nor U16546 (N_16546,N_16444,N_16310);
nor U16547 (N_16547,N_16404,N_16261);
or U16548 (N_16548,N_16355,N_16408);
or U16549 (N_16549,N_16423,N_16045);
nor U16550 (N_16550,N_16123,N_16192);
nand U16551 (N_16551,N_16231,N_16153);
and U16552 (N_16552,N_16181,N_16416);
nand U16553 (N_16553,N_16298,N_16221);
xnor U16554 (N_16554,N_16087,N_16292);
nand U16555 (N_16555,N_16270,N_16075);
and U16556 (N_16556,N_16245,N_16324);
and U16557 (N_16557,N_16207,N_16441);
or U16558 (N_16558,N_16210,N_16035);
xor U16559 (N_16559,N_16194,N_16437);
and U16560 (N_16560,N_16249,N_16274);
nand U16561 (N_16561,N_16147,N_16178);
xnor U16562 (N_16562,N_16029,N_16447);
xor U16563 (N_16563,N_16179,N_16120);
xor U16564 (N_16564,N_16014,N_16401);
nand U16565 (N_16565,N_16163,N_16373);
or U16566 (N_16566,N_16176,N_16406);
nor U16567 (N_16567,N_16005,N_16440);
nor U16568 (N_16568,N_16384,N_16219);
and U16569 (N_16569,N_16452,N_16046);
or U16570 (N_16570,N_16032,N_16479);
nand U16571 (N_16571,N_16497,N_16330);
or U16572 (N_16572,N_16213,N_16338);
nand U16573 (N_16573,N_16105,N_16258);
xnor U16574 (N_16574,N_16275,N_16125);
and U16575 (N_16575,N_16012,N_16429);
and U16576 (N_16576,N_16090,N_16312);
xnor U16577 (N_16577,N_16466,N_16057);
or U16578 (N_16578,N_16445,N_16432);
nor U16579 (N_16579,N_16252,N_16069);
nor U16580 (N_16580,N_16169,N_16442);
nor U16581 (N_16581,N_16288,N_16203);
xor U16582 (N_16582,N_16419,N_16054);
or U16583 (N_16583,N_16250,N_16454);
or U16584 (N_16584,N_16489,N_16174);
xnor U16585 (N_16585,N_16300,N_16119);
xnor U16586 (N_16586,N_16480,N_16130);
and U16587 (N_16587,N_16023,N_16084);
xnor U16588 (N_16588,N_16077,N_16074);
or U16589 (N_16589,N_16058,N_16049);
xnor U16590 (N_16590,N_16395,N_16073);
nor U16591 (N_16591,N_16173,N_16086);
and U16592 (N_16592,N_16451,N_16286);
or U16593 (N_16593,N_16154,N_16313);
xnor U16594 (N_16594,N_16279,N_16415);
and U16595 (N_16595,N_16094,N_16111);
xnor U16596 (N_16596,N_16450,N_16468);
nor U16597 (N_16597,N_16040,N_16290);
or U16598 (N_16598,N_16234,N_16294);
xor U16599 (N_16599,N_16396,N_16392);
or U16600 (N_16600,N_16438,N_16063);
nand U16601 (N_16601,N_16182,N_16374);
nand U16602 (N_16602,N_16293,N_16459);
nor U16603 (N_16603,N_16435,N_16295);
nor U16604 (N_16604,N_16030,N_16413);
or U16605 (N_16605,N_16342,N_16222);
or U16606 (N_16606,N_16331,N_16278);
nand U16607 (N_16607,N_16193,N_16305);
nor U16608 (N_16608,N_16358,N_16189);
or U16609 (N_16609,N_16284,N_16076);
nand U16610 (N_16610,N_16376,N_16236);
xor U16611 (N_16611,N_16443,N_16083);
or U16612 (N_16612,N_16257,N_16124);
xnor U16613 (N_16613,N_16280,N_16322);
nand U16614 (N_16614,N_16344,N_16088);
xnor U16615 (N_16615,N_16216,N_16446);
and U16616 (N_16616,N_16385,N_16047);
xnor U16617 (N_16617,N_16001,N_16140);
nand U16618 (N_16618,N_16414,N_16494);
nand U16619 (N_16619,N_16115,N_16455);
or U16620 (N_16620,N_16051,N_16363);
and U16621 (N_16621,N_16218,N_16127);
nor U16622 (N_16622,N_16418,N_16349);
xnor U16623 (N_16623,N_16048,N_16175);
or U16624 (N_16624,N_16244,N_16260);
and U16625 (N_16625,N_16318,N_16085);
nand U16626 (N_16626,N_16078,N_16139);
xor U16627 (N_16627,N_16038,N_16467);
nand U16628 (N_16628,N_16335,N_16167);
nor U16629 (N_16629,N_16329,N_16493);
xor U16630 (N_16630,N_16425,N_16378);
or U16631 (N_16631,N_16453,N_16360);
nand U16632 (N_16632,N_16059,N_16166);
nand U16633 (N_16633,N_16499,N_16171);
nor U16634 (N_16634,N_16431,N_16475);
or U16635 (N_16635,N_16304,N_16492);
and U16636 (N_16636,N_16356,N_16021);
xnor U16637 (N_16637,N_16017,N_16474);
nor U16638 (N_16638,N_16131,N_16496);
and U16639 (N_16639,N_16212,N_16104);
or U16640 (N_16640,N_16050,N_16190);
and U16641 (N_16641,N_16490,N_16132);
xor U16642 (N_16642,N_16272,N_16326);
or U16643 (N_16643,N_16135,N_16156);
nand U16644 (N_16644,N_16152,N_16162);
nand U16645 (N_16645,N_16239,N_16255);
and U16646 (N_16646,N_16161,N_16072);
nor U16647 (N_16647,N_16391,N_16388);
nand U16648 (N_16648,N_16037,N_16055);
and U16649 (N_16649,N_16064,N_16108);
or U16650 (N_16650,N_16427,N_16299);
nor U16651 (N_16651,N_16044,N_16387);
and U16652 (N_16652,N_16146,N_16113);
and U16653 (N_16653,N_16224,N_16319);
nor U16654 (N_16654,N_16381,N_16348);
or U16655 (N_16655,N_16092,N_16150);
or U16656 (N_16656,N_16316,N_16291);
nor U16657 (N_16657,N_16109,N_16398);
xor U16658 (N_16658,N_16263,N_16491);
and U16659 (N_16659,N_16371,N_16033);
xor U16660 (N_16660,N_16417,N_16142);
and U16661 (N_16661,N_16383,N_16367);
nand U16662 (N_16662,N_16235,N_16183);
nor U16663 (N_16663,N_16081,N_16112);
xnor U16664 (N_16664,N_16259,N_16025);
or U16665 (N_16665,N_16080,N_16266);
nand U16666 (N_16666,N_16019,N_16397);
and U16667 (N_16667,N_16434,N_16188);
and U16668 (N_16668,N_16296,N_16144);
nand U16669 (N_16669,N_16285,N_16053);
nand U16670 (N_16670,N_16379,N_16066);
nand U16671 (N_16671,N_16079,N_16495);
xor U16672 (N_16672,N_16121,N_16061);
nor U16673 (N_16673,N_16068,N_16015);
or U16674 (N_16674,N_16118,N_16470);
and U16675 (N_16675,N_16102,N_16230);
nor U16676 (N_16676,N_16339,N_16372);
or U16677 (N_16677,N_16448,N_16243);
xor U16678 (N_16678,N_16327,N_16287);
nand U16679 (N_16679,N_16165,N_16420);
and U16680 (N_16680,N_16343,N_16315);
xor U16681 (N_16681,N_16197,N_16185);
or U16682 (N_16682,N_16289,N_16036);
and U16683 (N_16683,N_16226,N_16082);
or U16684 (N_16684,N_16353,N_16070);
xor U16685 (N_16685,N_16211,N_16062);
xor U16686 (N_16686,N_16110,N_16020);
xor U16687 (N_16687,N_16457,N_16405);
nor U16688 (N_16688,N_16341,N_16399);
nand U16689 (N_16689,N_16201,N_16370);
nor U16690 (N_16690,N_16465,N_16191);
and U16691 (N_16691,N_16482,N_16402);
and U16692 (N_16692,N_16177,N_16462);
or U16693 (N_16693,N_16325,N_16277);
nand U16694 (N_16694,N_16357,N_16099);
xor U16695 (N_16695,N_16101,N_16056);
nand U16696 (N_16696,N_16334,N_16180);
and U16697 (N_16697,N_16008,N_16114);
xnor U16698 (N_16698,N_16365,N_16158);
and U16699 (N_16699,N_16386,N_16151);
and U16700 (N_16700,N_16238,N_16366);
nor U16701 (N_16701,N_16347,N_16393);
nand U16702 (N_16702,N_16227,N_16464);
or U16703 (N_16703,N_16463,N_16041);
nor U16704 (N_16704,N_16129,N_16039);
and U16705 (N_16705,N_16141,N_16052);
xnor U16706 (N_16706,N_16229,N_16247);
nand U16707 (N_16707,N_16018,N_16128);
xor U16708 (N_16708,N_16246,N_16009);
or U16709 (N_16709,N_16403,N_16208);
nor U16710 (N_16710,N_16251,N_16241);
and U16711 (N_16711,N_16306,N_16137);
nand U16712 (N_16712,N_16409,N_16478);
or U16713 (N_16713,N_16157,N_16202);
nand U16714 (N_16714,N_16433,N_16097);
xnor U16715 (N_16715,N_16407,N_16369);
nand U16716 (N_16716,N_16003,N_16382);
and U16717 (N_16717,N_16308,N_16095);
and U16718 (N_16718,N_16133,N_16011);
nor U16719 (N_16719,N_16328,N_16043);
nor U16720 (N_16720,N_16060,N_16172);
or U16721 (N_16721,N_16013,N_16065);
and U16722 (N_16722,N_16364,N_16377);
nor U16723 (N_16723,N_16148,N_16205);
nor U16724 (N_16724,N_16430,N_16248);
xor U16725 (N_16725,N_16002,N_16160);
or U16726 (N_16726,N_16164,N_16149);
or U16727 (N_16727,N_16100,N_16027);
xor U16728 (N_16728,N_16488,N_16346);
nand U16729 (N_16729,N_16187,N_16126);
nor U16730 (N_16730,N_16228,N_16022);
and U16731 (N_16731,N_16307,N_16426);
nand U16732 (N_16732,N_16484,N_16368);
or U16733 (N_16733,N_16004,N_16473);
nand U16734 (N_16734,N_16220,N_16282);
and U16735 (N_16735,N_16302,N_16421);
xor U16736 (N_16736,N_16145,N_16390);
or U16737 (N_16737,N_16317,N_16273);
and U16738 (N_16738,N_16461,N_16026);
nand U16739 (N_16739,N_16067,N_16096);
nand U16740 (N_16740,N_16311,N_16184);
nand U16741 (N_16741,N_16424,N_16345);
or U16742 (N_16742,N_16256,N_16071);
or U16743 (N_16743,N_16122,N_16268);
nand U16744 (N_16744,N_16010,N_16283);
or U16745 (N_16745,N_16458,N_16116);
or U16746 (N_16746,N_16232,N_16456);
nor U16747 (N_16747,N_16170,N_16436);
nand U16748 (N_16748,N_16253,N_16487);
xnor U16749 (N_16749,N_16321,N_16098);
and U16750 (N_16750,N_16492,N_16370);
or U16751 (N_16751,N_16410,N_16240);
and U16752 (N_16752,N_16036,N_16432);
and U16753 (N_16753,N_16267,N_16358);
and U16754 (N_16754,N_16055,N_16290);
and U16755 (N_16755,N_16238,N_16491);
nor U16756 (N_16756,N_16086,N_16332);
nor U16757 (N_16757,N_16376,N_16049);
xnor U16758 (N_16758,N_16247,N_16489);
xor U16759 (N_16759,N_16184,N_16488);
nand U16760 (N_16760,N_16255,N_16163);
xor U16761 (N_16761,N_16359,N_16173);
xnor U16762 (N_16762,N_16175,N_16297);
and U16763 (N_16763,N_16205,N_16249);
xnor U16764 (N_16764,N_16427,N_16297);
and U16765 (N_16765,N_16409,N_16093);
nand U16766 (N_16766,N_16387,N_16397);
xnor U16767 (N_16767,N_16125,N_16183);
nor U16768 (N_16768,N_16315,N_16101);
nand U16769 (N_16769,N_16188,N_16077);
and U16770 (N_16770,N_16122,N_16272);
nor U16771 (N_16771,N_16021,N_16311);
xnor U16772 (N_16772,N_16103,N_16011);
xnor U16773 (N_16773,N_16011,N_16090);
xor U16774 (N_16774,N_16036,N_16211);
nor U16775 (N_16775,N_16389,N_16178);
nor U16776 (N_16776,N_16218,N_16222);
or U16777 (N_16777,N_16395,N_16139);
nor U16778 (N_16778,N_16043,N_16481);
nor U16779 (N_16779,N_16202,N_16323);
xor U16780 (N_16780,N_16057,N_16043);
nor U16781 (N_16781,N_16309,N_16123);
nor U16782 (N_16782,N_16173,N_16300);
or U16783 (N_16783,N_16300,N_16212);
nand U16784 (N_16784,N_16204,N_16337);
or U16785 (N_16785,N_16403,N_16188);
xnor U16786 (N_16786,N_16111,N_16041);
nand U16787 (N_16787,N_16291,N_16343);
xor U16788 (N_16788,N_16338,N_16026);
or U16789 (N_16789,N_16247,N_16106);
nor U16790 (N_16790,N_16258,N_16413);
or U16791 (N_16791,N_16454,N_16238);
nand U16792 (N_16792,N_16431,N_16390);
and U16793 (N_16793,N_16370,N_16095);
nand U16794 (N_16794,N_16285,N_16206);
xnor U16795 (N_16795,N_16133,N_16233);
nor U16796 (N_16796,N_16405,N_16131);
xor U16797 (N_16797,N_16020,N_16306);
and U16798 (N_16798,N_16322,N_16146);
nor U16799 (N_16799,N_16261,N_16236);
nand U16800 (N_16800,N_16019,N_16407);
and U16801 (N_16801,N_16083,N_16063);
nand U16802 (N_16802,N_16263,N_16170);
nor U16803 (N_16803,N_16131,N_16445);
xnor U16804 (N_16804,N_16448,N_16423);
xnor U16805 (N_16805,N_16461,N_16242);
xnor U16806 (N_16806,N_16193,N_16131);
nor U16807 (N_16807,N_16205,N_16063);
or U16808 (N_16808,N_16014,N_16055);
or U16809 (N_16809,N_16108,N_16083);
xnor U16810 (N_16810,N_16133,N_16184);
or U16811 (N_16811,N_16466,N_16069);
nor U16812 (N_16812,N_16400,N_16010);
xnor U16813 (N_16813,N_16281,N_16187);
or U16814 (N_16814,N_16009,N_16161);
nand U16815 (N_16815,N_16205,N_16072);
nand U16816 (N_16816,N_16002,N_16327);
nand U16817 (N_16817,N_16139,N_16203);
and U16818 (N_16818,N_16476,N_16105);
xnor U16819 (N_16819,N_16105,N_16329);
or U16820 (N_16820,N_16208,N_16274);
and U16821 (N_16821,N_16305,N_16045);
xnor U16822 (N_16822,N_16346,N_16300);
xor U16823 (N_16823,N_16189,N_16240);
nor U16824 (N_16824,N_16028,N_16405);
nand U16825 (N_16825,N_16412,N_16074);
or U16826 (N_16826,N_16273,N_16103);
nand U16827 (N_16827,N_16053,N_16262);
nor U16828 (N_16828,N_16112,N_16220);
nand U16829 (N_16829,N_16280,N_16039);
nor U16830 (N_16830,N_16122,N_16106);
xnor U16831 (N_16831,N_16084,N_16027);
xnor U16832 (N_16832,N_16184,N_16418);
xnor U16833 (N_16833,N_16093,N_16070);
and U16834 (N_16834,N_16131,N_16400);
and U16835 (N_16835,N_16479,N_16376);
nand U16836 (N_16836,N_16065,N_16192);
nand U16837 (N_16837,N_16343,N_16483);
nor U16838 (N_16838,N_16462,N_16165);
nand U16839 (N_16839,N_16269,N_16009);
xor U16840 (N_16840,N_16492,N_16011);
xor U16841 (N_16841,N_16123,N_16086);
and U16842 (N_16842,N_16281,N_16006);
xor U16843 (N_16843,N_16048,N_16146);
or U16844 (N_16844,N_16285,N_16488);
nor U16845 (N_16845,N_16054,N_16263);
xnor U16846 (N_16846,N_16257,N_16239);
nand U16847 (N_16847,N_16044,N_16447);
nor U16848 (N_16848,N_16354,N_16186);
nand U16849 (N_16849,N_16085,N_16033);
nand U16850 (N_16850,N_16414,N_16283);
or U16851 (N_16851,N_16256,N_16101);
or U16852 (N_16852,N_16338,N_16188);
xnor U16853 (N_16853,N_16074,N_16141);
and U16854 (N_16854,N_16430,N_16363);
and U16855 (N_16855,N_16056,N_16480);
or U16856 (N_16856,N_16143,N_16285);
xor U16857 (N_16857,N_16340,N_16306);
or U16858 (N_16858,N_16161,N_16348);
xnor U16859 (N_16859,N_16189,N_16313);
and U16860 (N_16860,N_16272,N_16446);
nor U16861 (N_16861,N_16394,N_16342);
and U16862 (N_16862,N_16395,N_16089);
nand U16863 (N_16863,N_16232,N_16392);
xnor U16864 (N_16864,N_16458,N_16257);
or U16865 (N_16865,N_16006,N_16200);
xnor U16866 (N_16866,N_16211,N_16273);
and U16867 (N_16867,N_16258,N_16004);
nor U16868 (N_16868,N_16119,N_16058);
and U16869 (N_16869,N_16361,N_16483);
and U16870 (N_16870,N_16379,N_16308);
xnor U16871 (N_16871,N_16498,N_16056);
nand U16872 (N_16872,N_16027,N_16008);
or U16873 (N_16873,N_16258,N_16240);
and U16874 (N_16874,N_16370,N_16464);
xnor U16875 (N_16875,N_16122,N_16172);
and U16876 (N_16876,N_16296,N_16292);
or U16877 (N_16877,N_16057,N_16048);
xnor U16878 (N_16878,N_16295,N_16423);
or U16879 (N_16879,N_16151,N_16108);
and U16880 (N_16880,N_16171,N_16208);
xor U16881 (N_16881,N_16194,N_16249);
nor U16882 (N_16882,N_16172,N_16181);
nand U16883 (N_16883,N_16469,N_16015);
nand U16884 (N_16884,N_16315,N_16287);
nand U16885 (N_16885,N_16125,N_16496);
and U16886 (N_16886,N_16244,N_16331);
nand U16887 (N_16887,N_16480,N_16469);
or U16888 (N_16888,N_16399,N_16397);
xnor U16889 (N_16889,N_16439,N_16482);
xor U16890 (N_16890,N_16132,N_16289);
or U16891 (N_16891,N_16108,N_16245);
nor U16892 (N_16892,N_16313,N_16499);
and U16893 (N_16893,N_16415,N_16150);
nand U16894 (N_16894,N_16421,N_16301);
nor U16895 (N_16895,N_16429,N_16308);
nand U16896 (N_16896,N_16439,N_16278);
xnor U16897 (N_16897,N_16226,N_16253);
nand U16898 (N_16898,N_16121,N_16106);
nand U16899 (N_16899,N_16277,N_16192);
xor U16900 (N_16900,N_16028,N_16046);
nand U16901 (N_16901,N_16427,N_16160);
xnor U16902 (N_16902,N_16108,N_16435);
nor U16903 (N_16903,N_16489,N_16069);
and U16904 (N_16904,N_16092,N_16094);
or U16905 (N_16905,N_16236,N_16375);
nor U16906 (N_16906,N_16418,N_16062);
and U16907 (N_16907,N_16288,N_16457);
xnor U16908 (N_16908,N_16303,N_16130);
xnor U16909 (N_16909,N_16156,N_16188);
nand U16910 (N_16910,N_16466,N_16351);
nand U16911 (N_16911,N_16230,N_16136);
nor U16912 (N_16912,N_16310,N_16198);
or U16913 (N_16913,N_16258,N_16111);
nor U16914 (N_16914,N_16032,N_16417);
and U16915 (N_16915,N_16387,N_16075);
xnor U16916 (N_16916,N_16375,N_16175);
xor U16917 (N_16917,N_16079,N_16271);
nand U16918 (N_16918,N_16269,N_16197);
and U16919 (N_16919,N_16414,N_16261);
xnor U16920 (N_16920,N_16319,N_16315);
and U16921 (N_16921,N_16173,N_16054);
or U16922 (N_16922,N_16400,N_16394);
nor U16923 (N_16923,N_16447,N_16453);
nand U16924 (N_16924,N_16060,N_16123);
and U16925 (N_16925,N_16202,N_16263);
or U16926 (N_16926,N_16406,N_16035);
nand U16927 (N_16927,N_16029,N_16069);
or U16928 (N_16928,N_16036,N_16112);
or U16929 (N_16929,N_16387,N_16461);
nor U16930 (N_16930,N_16186,N_16445);
and U16931 (N_16931,N_16331,N_16077);
or U16932 (N_16932,N_16469,N_16282);
nor U16933 (N_16933,N_16025,N_16020);
xor U16934 (N_16934,N_16172,N_16068);
or U16935 (N_16935,N_16358,N_16036);
and U16936 (N_16936,N_16343,N_16481);
nand U16937 (N_16937,N_16221,N_16143);
and U16938 (N_16938,N_16113,N_16256);
or U16939 (N_16939,N_16497,N_16438);
nand U16940 (N_16940,N_16370,N_16153);
and U16941 (N_16941,N_16164,N_16303);
nand U16942 (N_16942,N_16172,N_16201);
and U16943 (N_16943,N_16407,N_16005);
or U16944 (N_16944,N_16076,N_16271);
nand U16945 (N_16945,N_16139,N_16169);
and U16946 (N_16946,N_16143,N_16457);
nor U16947 (N_16947,N_16032,N_16224);
xor U16948 (N_16948,N_16207,N_16133);
and U16949 (N_16949,N_16235,N_16402);
nand U16950 (N_16950,N_16448,N_16011);
nand U16951 (N_16951,N_16473,N_16092);
and U16952 (N_16952,N_16076,N_16340);
or U16953 (N_16953,N_16390,N_16113);
nand U16954 (N_16954,N_16477,N_16365);
nand U16955 (N_16955,N_16302,N_16174);
nand U16956 (N_16956,N_16185,N_16026);
or U16957 (N_16957,N_16016,N_16318);
or U16958 (N_16958,N_16246,N_16292);
nor U16959 (N_16959,N_16444,N_16258);
nand U16960 (N_16960,N_16144,N_16397);
or U16961 (N_16961,N_16433,N_16135);
or U16962 (N_16962,N_16035,N_16467);
nand U16963 (N_16963,N_16183,N_16032);
and U16964 (N_16964,N_16320,N_16015);
nor U16965 (N_16965,N_16093,N_16281);
nor U16966 (N_16966,N_16088,N_16485);
and U16967 (N_16967,N_16491,N_16432);
and U16968 (N_16968,N_16415,N_16333);
nand U16969 (N_16969,N_16089,N_16199);
nor U16970 (N_16970,N_16418,N_16483);
nand U16971 (N_16971,N_16160,N_16109);
or U16972 (N_16972,N_16156,N_16130);
nor U16973 (N_16973,N_16233,N_16009);
nand U16974 (N_16974,N_16032,N_16189);
and U16975 (N_16975,N_16147,N_16273);
xnor U16976 (N_16976,N_16062,N_16246);
xor U16977 (N_16977,N_16131,N_16111);
or U16978 (N_16978,N_16007,N_16297);
nor U16979 (N_16979,N_16157,N_16226);
or U16980 (N_16980,N_16231,N_16072);
xor U16981 (N_16981,N_16275,N_16317);
or U16982 (N_16982,N_16409,N_16191);
nand U16983 (N_16983,N_16234,N_16158);
and U16984 (N_16984,N_16472,N_16331);
or U16985 (N_16985,N_16445,N_16440);
and U16986 (N_16986,N_16030,N_16277);
nor U16987 (N_16987,N_16073,N_16339);
or U16988 (N_16988,N_16130,N_16277);
xnor U16989 (N_16989,N_16056,N_16007);
nand U16990 (N_16990,N_16387,N_16054);
or U16991 (N_16991,N_16409,N_16452);
nor U16992 (N_16992,N_16334,N_16023);
nand U16993 (N_16993,N_16490,N_16087);
and U16994 (N_16994,N_16481,N_16312);
nand U16995 (N_16995,N_16100,N_16035);
nor U16996 (N_16996,N_16276,N_16390);
and U16997 (N_16997,N_16145,N_16364);
or U16998 (N_16998,N_16490,N_16434);
and U16999 (N_16999,N_16105,N_16419);
or U17000 (N_17000,N_16650,N_16891);
and U17001 (N_17001,N_16642,N_16850);
nor U17002 (N_17002,N_16603,N_16592);
or U17003 (N_17003,N_16911,N_16829);
or U17004 (N_17004,N_16975,N_16768);
nand U17005 (N_17005,N_16969,N_16841);
or U17006 (N_17006,N_16851,N_16576);
or U17007 (N_17007,N_16888,N_16641);
xor U17008 (N_17008,N_16523,N_16818);
nor U17009 (N_17009,N_16549,N_16948);
nor U17010 (N_17010,N_16836,N_16540);
or U17011 (N_17011,N_16716,N_16725);
nor U17012 (N_17012,N_16628,N_16820);
or U17013 (N_17013,N_16580,N_16504);
xnor U17014 (N_17014,N_16532,N_16506);
xnor U17015 (N_17015,N_16552,N_16620);
and U17016 (N_17016,N_16800,N_16864);
and U17017 (N_17017,N_16584,N_16600);
xor U17018 (N_17018,N_16702,N_16508);
xnor U17019 (N_17019,N_16722,N_16717);
nor U17020 (N_17020,N_16846,N_16700);
xor U17021 (N_17021,N_16994,N_16827);
nor U17022 (N_17022,N_16723,N_16572);
or U17023 (N_17023,N_16941,N_16536);
or U17024 (N_17024,N_16714,N_16676);
nand U17025 (N_17025,N_16682,N_16883);
nand U17026 (N_17026,N_16654,N_16644);
and U17027 (N_17027,N_16880,N_16602);
nor U17028 (N_17028,N_16967,N_16885);
or U17029 (N_17029,N_16869,N_16957);
nand U17030 (N_17030,N_16806,N_16944);
nor U17031 (N_17031,N_16770,N_16742);
or U17032 (N_17032,N_16787,N_16597);
nor U17033 (N_17033,N_16908,N_16530);
nor U17034 (N_17034,N_16962,N_16838);
xor U17035 (N_17035,N_16522,N_16560);
xor U17036 (N_17036,N_16949,N_16807);
xnor U17037 (N_17037,N_16951,N_16637);
xor U17038 (N_17038,N_16832,N_16712);
nand U17039 (N_17039,N_16929,N_16866);
xor U17040 (N_17040,N_16614,N_16629);
nor U17041 (N_17041,N_16884,N_16808);
or U17042 (N_17042,N_16659,N_16855);
or U17043 (N_17043,N_16663,N_16879);
xor U17044 (N_17044,N_16652,N_16976);
and U17045 (N_17045,N_16763,N_16538);
and U17046 (N_17046,N_16664,N_16781);
nand U17047 (N_17047,N_16568,N_16814);
or U17048 (N_17048,N_16694,N_16871);
xor U17049 (N_17049,N_16837,N_16783);
xor U17050 (N_17050,N_16862,N_16860);
or U17051 (N_17051,N_16945,N_16968);
nor U17052 (N_17052,N_16713,N_16805);
and U17053 (N_17053,N_16925,N_16978);
nand U17054 (N_17054,N_16982,N_16639);
nand U17055 (N_17055,N_16749,N_16582);
or U17056 (N_17056,N_16902,N_16852);
nor U17057 (N_17057,N_16704,N_16821);
and U17058 (N_17058,N_16943,N_16526);
nor U17059 (N_17059,N_16502,N_16766);
and U17060 (N_17060,N_16686,N_16583);
xor U17061 (N_17061,N_16934,N_16971);
xnor U17062 (N_17062,N_16634,N_16559);
and U17063 (N_17063,N_16990,N_16824);
nor U17064 (N_17064,N_16692,N_16845);
nor U17065 (N_17065,N_16760,N_16701);
xnor U17066 (N_17066,N_16876,N_16550);
or U17067 (N_17067,N_16610,N_16563);
nor U17068 (N_17068,N_16615,N_16698);
and U17069 (N_17069,N_16589,N_16541);
or U17070 (N_17070,N_16985,N_16533);
nor U17071 (N_17071,N_16786,N_16525);
or U17072 (N_17072,N_16794,N_16791);
xnor U17073 (N_17073,N_16660,N_16816);
and U17074 (N_17074,N_16619,N_16956);
and U17075 (N_17075,N_16570,N_16581);
or U17076 (N_17076,N_16632,N_16859);
or U17077 (N_17077,N_16979,N_16656);
or U17078 (N_17078,N_16905,N_16718);
and U17079 (N_17079,N_16796,N_16733);
nand U17080 (N_17080,N_16882,N_16697);
xor U17081 (N_17081,N_16510,N_16801);
nand U17082 (N_17082,N_16752,N_16890);
nor U17083 (N_17083,N_16939,N_16542);
nor U17084 (N_17084,N_16761,N_16972);
nor U17085 (N_17085,N_16548,N_16566);
or U17086 (N_17086,N_16847,N_16710);
or U17087 (N_17087,N_16679,N_16907);
nor U17088 (N_17088,N_16622,N_16605);
or U17089 (N_17089,N_16735,N_16739);
or U17090 (N_17090,N_16731,N_16553);
or U17091 (N_17091,N_16751,N_16935);
xnor U17092 (N_17092,N_16771,N_16661);
or U17093 (N_17093,N_16591,N_16831);
xnor U17094 (N_17094,N_16812,N_16684);
nand U17095 (N_17095,N_16928,N_16789);
nor U17096 (N_17096,N_16782,N_16916);
and U17097 (N_17097,N_16788,N_16810);
or U17098 (N_17098,N_16987,N_16743);
or U17099 (N_17099,N_16547,N_16678);
and U17100 (N_17100,N_16887,N_16623);
xnor U17101 (N_17101,N_16625,N_16844);
nand U17102 (N_17102,N_16912,N_16728);
nor U17103 (N_17103,N_16598,N_16993);
nand U17104 (N_17104,N_16817,N_16609);
nand U17105 (N_17105,N_16587,N_16578);
xnor U17106 (N_17106,N_16618,N_16734);
and U17107 (N_17107,N_16670,N_16727);
nand U17108 (N_17108,N_16989,N_16558);
nand U17109 (N_17109,N_16653,N_16863);
nor U17110 (N_17110,N_16730,N_16937);
xnor U17111 (N_17111,N_16695,N_16872);
nand U17112 (N_17112,N_16640,N_16537);
nand U17113 (N_17113,N_16501,N_16953);
and U17114 (N_17114,N_16744,N_16999);
nor U17115 (N_17115,N_16569,N_16784);
nor U17116 (N_17116,N_16564,N_16726);
or U17117 (N_17117,N_16780,N_16599);
xnor U17118 (N_17118,N_16874,N_16843);
and U17119 (N_17119,N_16643,N_16966);
nor U17120 (N_17120,N_16936,N_16848);
xor U17121 (N_17121,N_16958,N_16938);
nand U17122 (N_17122,N_16724,N_16776);
nand U17123 (N_17123,N_16636,N_16970);
nor U17124 (N_17124,N_16804,N_16778);
nor U17125 (N_17125,N_16998,N_16894);
xor U17126 (N_17126,N_16895,N_16655);
nand U17127 (N_17127,N_16973,N_16903);
nor U17128 (N_17128,N_16875,N_16981);
and U17129 (N_17129,N_16608,N_16690);
nor U17130 (N_17130,N_16878,N_16516);
xor U17131 (N_17131,N_16899,N_16909);
nor U17132 (N_17132,N_16521,N_16915);
nor U17133 (N_17133,N_16834,N_16543);
or U17134 (N_17134,N_16961,N_16594);
nor U17135 (N_17135,N_16573,N_16896);
xor U17136 (N_17136,N_16685,N_16823);
xnor U17137 (N_17137,N_16666,N_16611);
or U17138 (N_17138,N_16940,N_16746);
or U17139 (N_17139,N_16926,N_16797);
and U17140 (N_17140,N_16767,N_16988);
nand U17141 (N_17141,N_16811,N_16507);
xor U17142 (N_17142,N_16631,N_16500);
or U17143 (N_17143,N_16930,N_16505);
or U17144 (N_17144,N_16921,N_16777);
and U17145 (N_17145,N_16539,N_16665);
xor U17146 (N_17146,N_16633,N_16853);
or U17147 (N_17147,N_16657,N_16849);
nor U17148 (N_17148,N_16842,N_16822);
and U17149 (N_17149,N_16952,N_16759);
nor U17150 (N_17150,N_16747,N_16520);
or U17151 (N_17151,N_16680,N_16933);
xnor U17152 (N_17152,N_16964,N_16986);
nand U17153 (N_17153,N_16877,N_16529);
nor U17154 (N_17154,N_16512,N_16906);
nand U17155 (N_17155,N_16828,N_16977);
nand U17156 (N_17156,N_16518,N_16901);
or U17157 (N_17157,N_16946,N_16544);
or U17158 (N_17158,N_16696,N_16980);
nor U17159 (N_17159,N_16960,N_16571);
nand U17160 (N_17160,N_16721,N_16719);
nor U17161 (N_17161,N_16865,N_16715);
xnor U17162 (N_17162,N_16813,N_16647);
or U17163 (N_17163,N_16511,N_16586);
and U17164 (N_17164,N_16554,N_16590);
xor U17165 (N_17165,N_16748,N_16606);
or U17166 (N_17166,N_16919,N_16681);
or U17167 (N_17167,N_16893,N_16914);
or U17168 (N_17168,N_16997,N_16509);
or U17169 (N_17169,N_16992,N_16840);
and U17170 (N_17170,N_16672,N_16658);
nor U17171 (N_17171,N_16924,N_16612);
nor U17172 (N_17172,N_16923,N_16826);
and U17173 (N_17173,N_16984,N_16892);
or U17174 (N_17174,N_16861,N_16668);
xnor U17175 (N_17175,N_16732,N_16708);
and U17176 (N_17176,N_16709,N_16870);
and U17177 (N_17177,N_16856,N_16996);
or U17178 (N_17178,N_16886,N_16833);
or U17179 (N_17179,N_16524,N_16562);
and U17180 (N_17180,N_16857,N_16764);
and U17181 (N_17181,N_16545,N_16556);
xor U17182 (N_17182,N_16792,N_16737);
nor U17183 (N_17183,N_16707,N_16942);
and U17184 (N_17184,N_16705,N_16900);
or U17185 (N_17185,N_16551,N_16630);
xnor U17186 (N_17186,N_16687,N_16624);
or U17187 (N_17187,N_16913,N_16617);
nand U17188 (N_17188,N_16585,N_16607);
nand U17189 (N_17189,N_16588,N_16677);
or U17190 (N_17190,N_16904,N_16755);
nand U17191 (N_17191,N_16762,N_16830);
xor U17192 (N_17192,N_16579,N_16503);
nand U17193 (N_17193,N_16881,N_16785);
or U17194 (N_17194,N_16897,N_16688);
nand U17195 (N_17195,N_16753,N_16621);
nor U17196 (N_17196,N_16574,N_16673);
or U17197 (N_17197,N_16867,N_16616);
nor U17198 (N_17198,N_16983,N_16635);
and U17199 (N_17199,N_16671,N_16674);
nor U17200 (N_17200,N_16745,N_16898);
xnor U17201 (N_17201,N_16662,N_16595);
xnor U17202 (N_17202,N_16645,N_16703);
nand U17203 (N_17203,N_16963,N_16527);
or U17204 (N_17204,N_16577,N_16575);
nand U17205 (N_17205,N_16738,N_16513);
nand U17206 (N_17206,N_16691,N_16922);
nor U17207 (N_17207,N_16803,N_16683);
xor U17208 (N_17208,N_16517,N_16754);
xnor U17209 (N_17209,N_16534,N_16531);
nor U17210 (N_17210,N_16868,N_16825);
and U17211 (N_17211,N_16561,N_16736);
nor U17212 (N_17212,N_16613,N_16995);
or U17213 (N_17213,N_16839,N_16918);
or U17214 (N_17214,N_16959,N_16950);
nor U17215 (N_17215,N_16910,N_16693);
and U17216 (N_17216,N_16515,N_16699);
or U17217 (N_17217,N_16798,N_16669);
or U17218 (N_17218,N_16858,N_16626);
xor U17219 (N_17219,N_16793,N_16648);
nand U17220 (N_17220,N_16773,N_16769);
xor U17221 (N_17221,N_16593,N_16774);
or U17222 (N_17222,N_16795,N_16651);
and U17223 (N_17223,N_16646,N_16689);
or U17224 (N_17224,N_16535,N_16756);
or U17225 (N_17225,N_16799,N_16889);
nor U17226 (N_17226,N_16775,N_16649);
or U17227 (N_17227,N_16557,N_16757);
nand U17228 (N_17228,N_16955,N_16974);
xnor U17229 (N_17229,N_16932,N_16604);
nor U17230 (N_17230,N_16931,N_16729);
nor U17231 (N_17231,N_16720,N_16706);
nor U17232 (N_17232,N_16991,N_16565);
or U17233 (N_17233,N_16740,N_16638);
and U17234 (N_17234,N_16667,N_16519);
nor U17235 (N_17235,N_16809,N_16920);
or U17236 (N_17236,N_16514,N_16835);
xor U17237 (N_17237,N_16675,N_16758);
or U17238 (N_17238,N_16815,N_16954);
xnor U17239 (N_17239,N_16627,N_16711);
and U17240 (N_17240,N_16567,N_16947);
nor U17241 (N_17241,N_16917,N_16765);
or U17242 (N_17242,N_16965,N_16596);
or U17243 (N_17243,N_16528,N_16741);
nand U17244 (N_17244,N_16854,N_16819);
and U17245 (N_17245,N_16873,N_16927);
nor U17246 (N_17246,N_16555,N_16802);
xnor U17247 (N_17247,N_16772,N_16546);
nor U17248 (N_17248,N_16779,N_16750);
and U17249 (N_17249,N_16601,N_16790);
nand U17250 (N_17250,N_16506,N_16706);
and U17251 (N_17251,N_16748,N_16874);
xor U17252 (N_17252,N_16902,N_16703);
xor U17253 (N_17253,N_16835,N_16786);
and U17254 (N_17254,N_16729,N_16990);
xnor U17255 (N_17255,N_16918,N_16545);
and U17256 (N_17256,N_16597,N_16876);
nor U17257 (N_17257,N_16699,N_16975);
nor U17258 (N_17258,N_16660,N_16843);
nor U17259 (N_17259,N_16749,N_16661);
nor U17260 (N_17260,N_16600,N_16738);
or U17261 (N_17261,N_16737,N_16584);
nor U17262 (N_17262,N_16619,N_16706);
or U17263 (N_17263,N_16695,N_16528);
nand U17264 (N_17264,N_16558,N_16718);
nand U17265 (N_17265,N_16924,N_16766);
or U17266 (N_17266,N_16521,N_16948);
nor U17267 (N_17267,N_16746,N_16511);
nand U17268 (N_17268,N_16589,N_16899);
xnor U17269 (N_17269,N_16897,N_16638);
nand U17270 (N_17270,N_16614,N_16745);
nand U17271 (N_17271,N_16668,N_16736);
nand U17272 (N_17272,N_16733,N_16663);
xnor U17273 (N_17273,N_16947,N_16897);
nor U17274 (N_17274,N_16637,N_16514);
and U17275 (N_17275,N_16830,N_16944);
xnor U17276 (N_17276,N_16616,N_16771);
nand U17277 (N_17277,N_16503,N_16600);
nor U17278 (N_17278,N_16842,N_16738);
nor U17279 (N_17279,N_16524,N_16505);
xor U17280 (N_17280,N_16875,N_16769);
nand U17281 (N_17281,N_16730,N_16656);
xnor U17282 (N_17282,N_16762,N_16911);
xor U17283 (N_17283,N_16509,N_16939);
xor U17284 (N_17284,N_16706,N_16569);
nand U17285 (N_17285,N_16920,N_16761);
nor U17286 (N_17286,N_16985,N_16755);
xor U17287 (N_17287,N_16738,N_16832);
nand U17288 (N_17288,N_16585,N_16781);
or U17289 (N_17289,N_16667,N_16679);
and U17290 (N_17290,N_16850,N_16727);
nand U17291 (N_17291,N_16640,N_16547);
nor U17292 (N_17292,N_16619,N_16726);
nor U17293 (N_17293,N_16842,N_16544);
or U17294 (N_17294,N_16767,N_16939);
or U17295 (N_17295,N_16734,N_16716);
and U17296 (N_17296,N_16904,N_16893);
nor U17297 (N_17297,N_16680,N_16738);
and U17298 (N_17298,N_16502,N_16585);
xor U17299 (N_17299,N_16587,N_16724);
nor U17300 (N_17300,N_16743,N_16884);
nor U17301 (N_17301,N_16547,N_16861);
and U17302 (N_17302,N_16798,N_16908);
or U17303 (N_17303,N_16661,N_16800);
nor U17304 (N_17304,N_16684,N_16920);
nor U17305 (N_17305,N_16917,N_16726);
or U17306 (N_17306,N_16598,N_16998);
nand U17307 (N_17307,N_16868,N_16762);
xor U17308 (N_17308,N_16649,N_16873);
xor U17309 (N_17309,N_16962,N_16815);
or U17310 (N_17310,N_16791,N_16989);
xor U17311 (N_17311,N_16672,N_16754);
nor U17312 (N_17312,N_16597,N_16830);
nor U17313 (N_17313,N_16824,N_16578);
or U17314 (N_17314,N_16799,N_16714);
nand U17315 (N_17315,N_16631,N_16993);
and U17316 (N_17316,N_16790,N_16746);
or U17317 (N_17317,N_16535,N_16544);
and U17318 (N_17318,N_16511,N_16540);
nor U17319 (N_17319,N_16605,N_16743);
xnor U17320 (N_17320,N_16973,N_16649);
xor U17321 (N_17321,N_16596,N_16744);
nand U17322 (N_17322,N_16620,N_16737);
and U17323 (N_17323,N_16632,N_16590);
and U17324 (N_17324,N_16848,N_16556);
or U17325 (N_17325,N_16797,N_16947);
xnor U17326 (N_17326,N_16931,N_16868);
and U17327 (N_17327,N_16697,N_16880);
nand U17328 (N_17328,N_16676,N_16897);
and U17329 (N_17329,N_16836,N_16589);
xnor U17330 (N_17330,N_16592,N_16913);
xor U17331 (N_17331,N_16703,N_16841);
nor U17332 (N_17332,N_16501,N_16579);
and U17333 (N_17333,N_16596,N_16865);
nand U17334 (N_17334,N_16931,N_16898);
nand U17335 (N_17335,N_16875,N_16912);
nand U17336 (N_17336,N_16524,N_16519);
nand U17337 (N_17337,N_16768,N_16867);
xor U17338 (N_17338,N_16779,N_16900);
or U17339 (N_17339,N_16811,N_16864);
nor U17340 (N_17340,N_16756,N_16732);
nand U17341 (N_17341,N_16569,N_16652);
nand U17342 (N_17342,N_16960,N_16658);
or U17343 (N_17343,N_16901,N_16995);
nand U17344 (N_17344,N_16686,N_16838);
and U17345 (N_17345,N_16609,N_16896);
or U17346 (N_17346,N_16773,N_16714);
xor U17347 (N_17347,N_16937,N_16873);
nor U17348 (N_17348,N_16640,N_16940);
nand U17349 (N_17349,N_16999,N_16692);
and U17350 (N_17350,N_16869,N_16523);
and U17351 (N_17351,N_16500,N_16913);
and U17352 (N_17352,N_16847,N_16556);
or U17353 (N_17353,N_16574,N_16645);
nor U17354 (N_17354,N_16949,N_16725);
or U17355 (N_17355,N_16931,N_16626);
nand U17356 (N_17356,N_16567,N_16912);
xnor U17357 (N_17357,N_16512,N_16870);
and U17358 (N_17358,N_16868,N_16808);
nand U17359 (N_17359,N_16666,N_16987);
or U17360 (N_17360,N_16737,N_16651);
or U17361 (N_17361,N_16549,N_16698);
nand U17362 (N_17362,N_16647,N_16797);
xor U17363 (N_17363,N_16586,N_16592);
xor U17364 (N_17364,N_16712,N_16861);
or U17365 (N_17365,N_16652,N_16534);
nand U17366 (N_17366,N_16935,N_16942);
nand U17367 (N_17367,N_16580,N_16914);
or U17368 (N_17368,N_16682,N_16622);
or U17369 (N_17369,N_16630,N_16729);
or U17370 (N_17370,N_16913,N_16902);
xor U17371 (N_17371,N_16845,N_16537);
or U17372 (N_17372,N_16967,N_16668);
nand U17373 (N_17373,N_16960,N_16634);
xnor U17374 (N_17374,N_16685,N_16510);
nand U17375 (N_17375,N_16793,N_16967);
xnor U17376 (N_17376,N_16808,N_16510);
and U17377 (N_17377,N_16945,N_16533);
nor U17378 (N_17378,N_16788,N_16897);
nor U17379 (N_17379,N_16759,N_16609);
or U17380 (N_17380,N_16570,N_16548);
and U17381 (N_17381,N_16908,N_16622);
or U17382 (N_17382,N_16598,N_16696);
nand U17383 (N_17383,N_16674,N_16519);
or U17384 (N_17384,N_16542,N_16897);
xor U17385 (N_17385,N_16887,N_16601);
nor U17386 (N_17386,N_16685,N_16972);
nor U17387 (N_17387,N_16881,N_16585);
or U17388 (N_17388,N_16583,N_16791);
nor U17389 (N_17389,N_16849,N_16925);
and U17390 (N_17390,N_16685,N_16847);
nor U17391 (N_17391,N_16913,N_16570);
and U17392 (N_17392,N_16504,N_16905);
and U17393 (N_17393,N_16580,N_16757);
nand U17394 (N_17394,N_16706,N_16559);
and U17395 (N_17395,N_16909,N_16949);
nand U17396 (N_17396,N_16911,N_16651);
nor U17397 (N_17397,N_16710,N_16889);
or U17398 (N_17398,N_16883,N_16839);
and U17399 (N_17399,N_16946,N_16859);
nor U17400 (N_17400,N_16578,N_16988);
nand U17401 (N_17401,N_16768,N_16589);
xor U17402 (N_17402,N_16689,N_16615);
nand U17403 (N_17403,N_16971,N_16729);
nor U17404 (N_17404,N_16583,N_16552);
xor U17405 (N_17405,N_16915,N_16702);
and U17406 (N_17406,N_16940,N_16828);
and U17407 (N_17407,N_16573,N_16612);
or U17408 (N_17408,N_16951,N_16862);
nand U17409 (N_17409,N_16521,N_16821);
nand U17410 (N_17410,N_16987,N_16684);
nor U17411 (N_17411,N_16565,N_16580);
xnor U17412 (N_17412,N_16578,N_16676);
nor U17413 (N_17413,N_16917,N_16715);
nor U17414 (N_17414,N_16789,N_16938);
and U17415 (N_17415,N_16552,N_16649);
nand U17416 (N_17416,N_16668,N_16516);
xnor U17417 (N_17417,N_16975,N_16966);
or U17418 (N_17418,N_16999,N_16828);
or U17419 (N_17419,N_16680,N_16562);
or U17420 (N_17420,N_16614,N_16937);
or U17421 (N_17421,N_16707,N_16857);
and U17422 (N_17422,N_16683,N_16677);
xor U17423 (N_17423,N_16879,N_16921);
or U17424 (N_17424,N_16641,N_16583);
nand U17425 (N_17425,N_16849,N_16616);
nor U17426 (N_17426,N_16780,N_16784);
xor U17427 (N_17427,N_16875,N_16639);
or U17428 (N_17428,N_16750,N_16741);
and U17429 (N_17429,N_16643,N_16866);
xnor U17430 (N_17430,N_16986,N_16719);
and U17431 (N_17431,N_16962,N_16857);
and U17432 (N_17432,N_16734,N_16635);
nor U17433 (N_17433,N_16816,N_16725);
xor U17434 (N_17434,N_16720,N_16820);
or U17435 (N_17435,N_16988,N_16616);
xor U17436 (N_17436,N_16613,N_16896);
xnor U17437 (N_17437,N_16710,N_16850);
xor U17438 (N_17438,N_16937,N_16900);
or U17439 (N_17439,N_16856,N_16518);
nand U17440 (N_17440,N_16925,N_16588);
xor U17441 (N_17441,N_16996,N_16789);
and U17442 (N_17442,N_16794,N_16784);
xor U17443 (N_17443,N_16961,N_16942);
xor U17444 (N_17444,N_16653,N_16804);
and U17445 (N_17445,N_16877,N_16931);
nor U17446 (N_17446,N_16849,N_16917);
and U17447 (N_17447,N_16803,N_16583);
nor U17448 (N_17448,N_16519,N_16988);
nand U17449 (N_17449,N_16618,N_16699);
nand U17450 (N_17450,N_16862,N_16850);
or U17451 (N_17451,N_16907,N_16824);
or U17452 (N_17452,N_16985,N_16541);
and U17453 (N_17453,N_16811,N_16675);
and U17454 (N_17454,N_16579,N_16748);
nor U17455 (N_17455,N_16515,N_16644);
nor U17456 (N_17456,N_16755,N_16544);
and U17457 (N_17457,N_16619,N_16836);
nand U17458 (N_17458,N_16767,N_16961);
nor U17459 (N_17459,N_16580,N_16836);
nor U17460 (N_17460,N_16898,N_16834);
and U17461 (N_17461,N_16818,N_16652);
or U17462 (N_17462,N_16699,N_16907);
and U17463 (N_17463,N_16983,N_16812);
nor U17464 (N_17464,N_16767,N_16569);
xnor U17465 (N_17465,N_16879,N_16651);
xor U17466 (N_17466,N_16744,N_16597);
and U17467 (N_17467,N_16582,N_16840);
or U17468 (N_17468,N_16511,N_16567);
nor U17469 (N_17469,N_16858,N_16806);
xnor U17470 (N_17470,N_16666,N_16668);
nor U17471 (N_17471,N_16994,N_16545);
nand U17472 (N_17472,N_16822,N_16612);
or U17473 (N_17473,N_16999,N_16869);
nand U17474 (N_17474,N_16836,N_16727);
or U17475 (N_17475,N_16918,N_16644);
or U17476 (N_17476,N_16858,N_16711);
or U17477 (N_17477,N_16532,N_16748);
nand U17478 (N_17478,N_16945,N_16658);
or U17479 (N_17479,N_16753,N_16790);
and U17480 (N_17480,N_16510,N_16979);
nor U17481 (N_17481,N_16807,N_16634);
nor U17482 (N_17482,N_16822,N_16883);
nand U17483 (N_17483,N_16596,N_16861);
and U17484 (N_17484,N_16987,N_16557);
xor U17485 (N_17485,N_16794,N_16988);
nand U17486 (N_17486,N_16918,N_16827);
nor U17487 (N_17487,N_16912,N_16984);
xnor U17488 (N_17488,N_16891,N_16657);
xor U17489 (N_17489,N_16504,N_16967);
nand U17490 (N_17490,N_16648,N_16540);
xnor U17491 (N_17491,N_16796,N_16805);
xor U17492 (N_17492,N_16729,N_16534);
xnor U17493 (N_17493,N_16573,N_16621);
or U17494 (N_17494,N_16704,N_16692);
and U17495 (N_17495,N_16925,N_16525);
xnor U17496 (N_17496,N_16587,N_16529);
nand U17497 (N_17497,N_16705,N_16785);
xor U17498 (N_17498,N_16670,N_16541);
and U17499 (N_17499,N_16874,N_16973);
nor U17500 (N_17500,N_17235,N_17357);
and U17501 (N_17501,N_17059,N_17405);
nand U17502 (N_17502,N_17363,N_17180);
and U17503 (N_17503,N_17300,N_17067);
xnor U17504 (N_17504,N_17491,N_17439);
nand U17505 (N_17505,N_17414,N_17062);
nor U17506 (N_17506,N_17438,N_17234);
nand U17507 (N_17507,N_17191,N_17375);
or U17508 (N_17508,N_17141,N_17273);
or U17509 (N_17509,N_17428,N_17205);
xnor U17510 (N_17510,N_17158,N_17098);
xnor U17511 (N_17511,N_17018,N_17167);
xnor U17512 (N_17512,N_17390,N_17053);
nor U17513 (N_17513,N_17242,N_17464);
xnor U17514 (N_17514,N_17123,N_17486);
or U17515 (N_17515,N_17055,N_17119);
or U17516 (N_17516,N_17407,N_17228);
nand U17517 (N_17517,N_17383,N_17259);
or U17518 (N_17518,N_17331,N_17134);
xor U17519 (N_17519,N_17083,N_17032);
nor U17520 (N_17520,N_17342,N_17297);
xnor U17521 (N_17521,N_17294,N_17366);
xnor U17522 (N_17522,N_17064,N_17304);
xnor U17523 (N_17523,N_17354,N_17254);
nand U17524 (N_17524,N_17328,N_17261);
nor U17525 (N_17525,N_17050,N_17310);
xor U17526 (N_17526,N_17468,N_17221);
and U17527 (N_17527,N_17105,N_17166);
and U17528 (N_17528,N_17135,N_17133);
and U17529 (N_17529,N_17301,N_17278);
or U17530 (N_17530,N_17217,N_17295);
nor U17531 (N_17531,N_17136,N_17401);
xnor U17532 (N_17532,N_17132,N_17449);
nor U17533 (N_17533,N_17475,N_17459);
nor U17534 (N_17534,N_17341,N_17125);
xor U17535 (N_17535,N_17356,N_17107);
nand U17536 (N_17536,N_17058,N_17084);
xor U17537 (N_17537,N_17418,N_17146);
or U17538 (N_17538,N_17149,N_17231);
and U17539 (N_17539,N_17121,N_17047);
xor U17540 (N_17540,N_17307,N_17264);
nor U17541 (N_17541,N_17026,N_17197);
nor U17542 (N_17542,N_17046,N_17040);
xor U17543 (N_17543,N_17049,N_17409);
xor U17544 (N_17544,N_17373,N_17408);
and U17545 (N_17545,N_17239,N_17493);
nand U17546 (N_17546,N_17069,N_17161);
xor U17547 (N_17547,N_17430,N_17332);
xor U17548 (N_17548,N_17226,N_17113);
or U17549 (N_17549,N_17483,N_17068);
xor U17550 (N_17550,N_17225,N_17413);
nand U17551 (N_17551,N_17453,N_17097);
or U17552 (N_17552,N_17402,N_17391);
and U17553 (N_17553,N_17024,N_17199);
nor U17554 (N_17554,N_17150,N_17292);
xnor U17555 (N_17555,N_17041,N_17089);
nand U17556 (N_17556,N_17033,N_17013);
nor U17557 (N_17557,N_17266,N_17017);
nor U17558 (N_17558,N_17496,N_17458);
nor U17559 (N_17559,N_17203,N_17284);
xnor U17560 (N_17560,N_17263,N_17081);
nand U17561 (N_17561,N_17382,N_17484);
nor U17562 (N_17562,N_17012,N_17425);
nand U17563 (N_17563,N_17060,N_17157);
nor U17564 (N_17564,N_17394,N_17378);
and U17565 (N_17565,N_17250,N_17204);
nand U17566 (N_17566,N_17175,N_17074);
nand U17567 (N_17567,N_17014,N_17201);
xnor U17568 (N_17568,N_17256,N_17063);
and U17569 (N_17569,N_17258,N_17351);
nand U17570 (N_17570,N_17127,N_17392);
or U17571 (N_17571,N_17082,N_17470);
nor U17572 (N_17572,N_17224,N_17202);
nor U17573 (N_17573,N_17303,N_17473);
nor U17574 (N_17574,N_17232,N_17372);
or U17575 (N_17575,N_17251,N_17183);
or U17576 (N_17576,N_17079,N_17309);
and U17577 (N_17577,N_17291,N_17109);
or U17578 (N_17578,N_17393,N_17164);
xnor U17579 (N_17579,N_17102,N_17466);
and U17580 (N_17580,N_17078,N_17478);
nor U17581 (N_17581,N_17450,N_17215);
nand U17582 (N_17582,N_17262,N_17115);
nor U17583 (N_17583,N_17156,N_17005);
or U17584 (N_17584,N_17282,N_17452);
xor U17585 (N_17585,N_17054,N_17056);
and U17586 (N_17586,N_17290,N_17344);
or U17587 (N_17587,N_17260,N_17369);
or U17588 (N_17588,N_17209,N_17417);
and U17589 (N_17589,N_17171,N_17360);
and U17590 (N_17590,N_17326,N_17008);
and U17591 (N_17591,N_17038,N_17039);
nor U17592 (N_17592,N_17349,N_17480);
nor U17593 (N_17593,N_17442,N_17311);
nand U17594 (N_17594,N_17306,N_17196);
xnor U17595 (N_17595,N_17463,N_17287);
nand U17596 (N_17596,N_17230,N_17359);
xor U17597 (N_17597,N_17370,N_17499);
and U17598 (N_17598,N_17118,N_17159);
xnor U17599 (N_17599,N_17437,N_17172);
nor U17600 (N_17600,N_17211,N_17030);
nor U17601 (N_17601,N_17147,N_17364);
nand U17602 (N_17602,N_17451,N_17052);
xor U17603 (N_17603,N_17412,N_17028);
nor U17604 (N_17604,N_17322,N_17044);
nor U17605 (N_17605,N_17387,N_17186);
or U17606 (N_17606,N_17333,N_17461);
and U17607 (N_17607,N_17286,N_17214);
nor U17608 (N_17608,N_17396,N_17419);
nand U17609 (N_17609,N_17381,N_17248);
or U17610 (N_17610,N_17080,N_17353);
nor U17611 (N_17611,N_17241,N_17155);
nand U17612 (N_17612,N_17208,N_17388);
and U17613 (N_17613,N_17189,N_17144);
nor U17614 (N_17614,N_17361,N_17010);
nor U17615 (N_17615,N_17091,N_17151);
and U17616 (N_17616,N_17482,N_17034);
and U17617 (N_17617,N_17243,N_17210);
nor U17618 (N_17618,N_17002,N_17374);
xor U17619 (N_17619,N_17007,N_17276);
and U17620 (N_17620,N_17448,N_17165);
nor U17621 (N_17621,N_17272,N_17368);
nand U17622 (N_17622,N_17179,N_17293);
or U17623 (N_17623,N_17497,N_17488);
nand U17624 (N_17624,N_17045,N_17317);
nand U17625 (N_17625,N_17339,N_17298);
nor U17626 (N_17626,N_17173,N_17296);
or U17627 (N_17627,N_17384,N_17397);
nor U17628 (N_17628,N_17350,N_17376);
and U17629 (N_17629,N_17399,N_17279);
xor U17630 (N_17630,N_17435,N_17267);
xor U17631 (N_17631,N_17443,N_17077);
nand U17632 (N_17632,N_17108,N_17335);
or U17633 (N_17633,N_17070,N_17492);
and U17634 (N_17634,N_17457,N_17330);
xor U17635 (N_17635,N_17145,N_17275);
nand U17636 (N_17636,N_17240,N_17462);
nand U17637 (N_17637,N_17410,N_17043);
nand U17638 (N_17638,N_17416,N_17093);
or U17639 (N_17639,N_17073,N_17142);
or U17640 (N_17640,N_17465,N_17244);
nor U17641 (N_17641,N_17117,N_17479);
or U17642 (N_17642,N_17444,N_17122);
xor U17643 (N_17643,N_17020,N_17222);
xnor U17644 (N_17644,N_17101,N_17498);
nor U17645 (N_17645,N_17269,N_17036);
and U17646 (N_17646,N_17429,N_17015);
and U17647 (N_17647,N_17371,N_17238);
xnor U17648 (N_17648,N_17398,N_17340);
nor U17649 (N_17649,N_17162,N_17087);
nor U17650 (N_17650,N_17207,N_17178);
nand U17651 (N_17651,N_17253,N_17403);
and U17652 (N_17652,N_17433,N_17111);
and U17653 (N_17653,N_17299,N_17312);
and U17654 (N_17654,N_17440,N_17346);
nor U17655 (N_17655,N_17386,N_17174);
xnor U17656 (N_17656,N_17138,N_17106);
nand U17657 (N_17657,N_17255,N_17424);
and U17658 (N_17658,N_17481,N_17185);
nand U17659 (N_17659,N_17427,N_17379);
nand U17660 (N_17660,N_17487,N_17358);
xnor U17661 (N_17661,N_17124,N_17200);
and U17662 (N_17662,N_17380,N_17277);
nand U17663 (N_17663,N_17229,N_17198);
xnor U17664 (N_17664,N_17065,N_17324);
nand U17665 (N_17665,N_17104,N_17152);
or U17666 (N_17666,N_17003,N_17153);
or U17667 (N_17667,N_17094,N_17103);
nand U17668 (N_17668,N_17423,N_17343);
and U17669 (N_17669,N_17137,N_17469);
nor U17670 (N_17670,N_17365,N_17216);
xor U17671 (N_17671,N_17170,N_17411);
xor U17672 (N_17672,N_17128,N_17195);
nand U17673 (N_17673,N_17004,N_17406);
nand U17674 (N_17674,N_17072,N_17130);
nand U17675 (N_17675,N_17252,N_17337);
nand U17676 (N_17676,N_17192,N_17131);
nor U17677 (N_17677,N_17057,N_17320);
and U17678 (N_17678,N_17329,N_17160);
nor U17679 (N_17679,N_17446,N_17110);
or U17680 (N_17680,N_17218,N_17494);
and U17681 (N_17681,N_17347,N_17400);
xor U17682 (N_17682,N_17169,N_17460);
xor U17683 (N_17683,N_17422,N_17318);
nand U17684 (N_17684,N_17177,N_17389);
nor U17685 (N_17685,N_17489,N_17431);
nand U17686 (N_17686,N_17313,N_17281);
or U17687 (N_17687,N_17323,N_17315);
and U17688 (N_17688,N_17247,N_17184);
xor U17689 (N_17689,N_17009,N_17420);
and U17690 (N_17690,N_17219,N_17114);
xor U17691 (N_17691,N_17445,N_17362);
nor U17692 (N_17692,N_17270,N_17176);
nor U17693 (N_17693,N_17436,N_17338);
or U17694 (N_17694,N_17071,N_17143);
nand U17695 (N_17695,N_17187,N_17120);
nor U17696 (N_17696,N_17265,N_17126);
nor U17697 (N_17697,N_17268,N_17285);
xnor U17698 (N_17698,N_17029,N_17289);
or U17699 (N_17699,N_17495,N_17139);
nor U17700 (N_17700,N_17181,N_17099);
xnor U17701 (N_17701,N_17352,N_17001);
xor U17702 (N_17702,N_17246,N_17377);
and U17703 (N_17703,N_17163,N_17140);
nand U17704 (N_17704,N_17095,N_17415);
nand U17705 (N_17705,N_17212,N_17245);
nor U17706 (N_17706,N_17336,N_17011);
nor U17707 (N_17707,N_17348,N_17100);
and U17708 (N_17708,N_17485,N_17085);
or U17709 (N_17709,N_17035,N_17021);
and U17710 (N_17710,N_17027,N_17325);
xnor U17711 (N_17711,N_17404,N_17148);
nor U17712 (N_17712,N_17314,N_17474);
xnor U17713 (N_17713,N_17447,N_17271);
nand U17714 (N_17714,N_17316,N_17233);
nand U17715 (N_17715,N_17037,N_17249);
or U17716 (N_17716,N_17455,N_17426);
xor U17717 (N_17717,N_17075,N_17319);
xor U17718 (N_17718,N_17395,N_17283);
nand U17719 (N_17719,N_17490,N_17237);
nor U17720 (N_17720,N_17334,N_17280);
xor U17721 (N_17721,N_17025,N_17385);
or U17722 (N_17722,N_17051,N_17193);
nor U17723 (N_17723,N_17477,N_17257);
or U17724 (N_17724,N_17454,N_17182);
xor U17725 (N_17725,N_17355,N_17112);
and U17726 (N_17726,N_17305,N_17194);
xnor U17727 (N_17727,N_17308,N_17129);
nand U17728 (N_17728,N_17288,N_17223);
or U17729 (N_17729,N_17220,N_17471);
and U17730 (N_17730,N_17154,N_17000);
or U17731 (N_17731,N_17345,N_17476);
or U17732 (N_17732,N_17092,N_17188);
or U17733 (N_17733,N_17088,N_17441);
and U17734 (N_17734,N_17274,N_17206);
nor U17735 (N_17735,N_17006,N_17090);
or U17736 (N_17736,N_17076,N_17472);
xnor U17737 (N_17737,N_17048,N_17213);
xor U17738 (N_17738,N_17302,N_17116);
or U17739 (N_17739,N_17227,N_17434);
xor U17740 (N_17740,N_17066,N_17421);
or U17741 (N_17741,N_17467,N_17168);
or U17742 (N_17742,N_17022,N_17456);
nand U17743 (N_17743,N_17031,N_17016);
and U17744 (N_17744,N_17327,N_17096);
xnor U17745 (N_17745,N_17019,N_17190);
nor U17746 (N_17746,N_17236,N_17432);
and U17747 (N_17747,N_17023,N_17086);
or U17748 (N_17748,N_17321,N_17367);
nand U17749 (N_17749,N_17042,N_17061);
xor U17750 (N_17750,N_17169,N_17323);
xnor U17751 (N_17751,N_17401,N_17285);
or U17752 (N_17752,N_17342,N_17253);
and U17753 (N_17753,N_17311,N_17017);
and U17754 (N_17754,N_17019,N_17040);
xnor U17755 (N_17755,N_17465,N_17488);
nor U17756 (N_17756,N_17240,N_17490);
xor U17757 (N_17757,N_17402,N_17489);
and U17758 (N_17758,N_17137,N_17441);
xnor U17759 (N_17759,N_17098,N_17291);
or U17760 (N_17760,N_17003,N_17420);
nor U17761 (N_17761,N_17085,N_17035);
nand U17762 (N_17762,N_17094,N_17338);
nand U17763 (N_17763,N_17034,N_17267);
xnor U17764 (N_17764,N_17292,N_17015);
or U17765 (N_17765,N_17275,N_17118);
or U17766 (N_17766,N_17468,N_17125);
and U17767 (N_17767,N_17019,N_17001);
and U17768 (N_17768,N_17324,N_17248);
or U17769 (N_17769,N_17320,N_17285);
and U17770 (N_17770,N_17021,N_17301);
or U17771 (N_17771,N_17441,N_17121);
nand U17772 (N_17772,N_17209,N_17242);
xor U17773 (N_17773,N_17481,N_17346);
and U17774 (N_17774,N_17238,N_17484);
and U17775 (N_17775,N_17325,N_17269);
nand U17776 (N_17776,N_17392,N_17228);
nand U17777 (N_17777,N_17444,N_17425);
nand U17778 (N_17778,N_17326,N_17484);
and U17779 (N_17779,N_17100,N_17093);
nand U17780 (N_17780,N_17335,N_17196);
nand U17781 (N_17781,N_17239,N_17468);
and U17782 (N_17782,N_17464,N_17314);
nor U17783 (N_17783,N_17496,N_17460);
or U17784 (N_17784,N_17215,N_17264);
and U17785 (N_17785,N_17270,N_17019);
or U17786 (N_17786,N_17001,N_17392);
and U17787 (N_17787,N_17159,N_17296);
xnor U17788 (N_17788,N_17234,N_17493);
or U17789 (N_17789,N_17302,N_17409);
xor U17790 (N_17790,N_17477,N_17299);
and U17791 (N_17791,N_17011,N_17099);
xnor U17792 (N_17792,N_17474,N_17198);
nor U17793 (N_17793,N_17330,N_17227);
nand U17794 (N_17794,N_17276,N_17329);
nor U17795 (N_17795,N_17494,N_17333);
xor U17796 (N_17796,N_17495,N_17131);
nor U17797 (N_17797,N_17354,N_17119);
nor U17798 (N_17798,N_17200,N_17184);
nand U17799 (N_17799,N_17472,N_17315);
xnor U17800 (N_17800,N_17030,N_17084);
or U17801 (N_17801,N_17118,N_17238);
xor U17802 (N_17802,N_17360,N_17274);
nor U17803 (N_17803,N_17365,N_17353);
nand U17804 (N_17804,N_17078,N_17062);
and U17805 (N_17805,N_17423,N_17107);
or U17806 (N_17806,N_17124,N_17305);
xor U17807 (N_17807,N_17369,N_17192);
nand U17808 (N_17808,N_17408,N_17466);
nand U17809 (N_17809,N_17346,N_17412);
nand U17810 (N_17810,N_17022,N_17416);
xnor U17811 (N_17811,N_17399,N_17443);
and U17812 (N_17812,N_17074,N_17073);
nand U17813 (N_17813,N_17223,N_17111);
and U17814 (N_17814,N_17094,N_17269);
nor U17815 (N_17815,N_17209,N_17004);
nand U17816 (N_17816,N_17294,N_17171);
nand U17817 (N_17817,N_17152,N_17384);
or U17818 (N_17818,N_17100,N_17249);
nand U17819 (N_17819,N_17233,N_17153);
or U17820 (N_17820,N_17148,N_17495);
and U17821 (N_17821,N_17053,N_17271);
or U17822 (N_17822,N_17175,N_17251);
nand U17823 (N_17823,N_17480,N_17352);
or U17824 (N_17824,N_17128,N_17306);
nand U17825 (N_17825,N_17035,N_17289);
nand U17826 (N_17826,N_17275,N_17074);
or U17827 (N_17827,N_17149,N_17362);
or U17828 (N_17828,N_17059,N_17142);
nand U17829 (N_17829,N_17138,N_17029);
nand U17830 (N_17830,N_17331,N_17018);
nor U17831 (N_17831,N_17247,N_17221);
or U17832 (N_17832,N_17319,N_17471);
nor U17833 (N_17833,N_17403,N_17339);
nor U17834 (N_17834,N_17081,N_17434);
nor U17835 (N_17835,N_17251,N_17433);
nand U17836 (N_17836,N_17112,N_17156);
xnor U17837 (N_17837,N_17187,N_17424);
and U17838 (N_17838,N_17360,N_17165);
nand U17839 (N_17839,N_17495,N_17493);
nand U17840 (N_17840,N_17180,N_17185);
nand U17841 (N_17841,N_17065,N_17298);
nand U17842 (N_17842,N_17257,N_17159);
xor U17843 (N_17843,N_17321,N_17238);
xnor U17844 (N_17844,N_17337,N_17154);
nor U17845 (N_17845,N_17118,N_17191);
nor U17846 (N_17846,N_17438,N_17293);
xnor U17847 (N_17847,N_17420,N_17263);
xor U17848 (N_17848,N_17320,N_17209);
nor U17849 (N_17849,N_17033,N_17163);
xor U17850 (N_17850,N_17106,N_17000);
and U17851 (N_17851,N_17303,N_17352);
or U17852 (N_17852,N_17449,N_17172);
xor U17853 (N_17853,N_17395,N_17488);
or U17854 (N_17854,N_17198,N_17157);
xnor U17855 (N_17855,N_17168,N_17386);
xor U17856 (N_17856,N_17403,N_17318);
or U17857 (N_17857,N_17452,N_17212);
and U17858 (N_17858,N_17105,N_17110);
nor U17859 (N_17859,N_17414,N_17119);
nor U17860 (N_17860,N_17316,N_17246);
and U17861 (N_17861,N_17310,N_17114);
or U17862 (N_17862,N_17463,N_17340);
nor U17863 (N_17863,N_17438,N_17246);
and U17864 (N_17864,N_17151,N_17156);
or U17865 (N_17865,N_17173,N_17394);
nand U17866 (N_17866,N_17148,N_17035);
or U17867 (N_17867,N_17475,N_17421);
xor U17868 (N_17868,N_17151,N_17043);
nand U17869 (N_17869,N_17076,N_17042);
and U17870 (N_17870,N_17416,N_17291);
nor U17871 (N_17871,N_17434,N_17041);
or U17872 (N_17872,N_17259,N_17004);
nand U17873 (N_17873,N_17157,N_17414);
nor U17874 (N_17874,N_17478,N_17020);
xor U17875 (N_17875,N_17195,N_17460);
or U17876 (N_17876,N_17372,N_17074);
and U17877 (N_17877,N_17203,N_17197);
xor U17878 (N_17878,N_17196,N_17125);
xor U17879 (N_17879,N_17052,N_17284);
xnor U17880 (N_17880,N_17332,N_17223);
or U17881 (N_17881,N_17200,N_17479);
or U17882 (N_17882,N_17383,N_17267);
nand U17883 (N_17883,N_17240,N_17202);
nand U17884 (N_17884,N_17224,N_17271);
or U17885 (N_17885,N_17331,N_17097);
nor U17886 (N_17886,N_17231,N_17498);
and U17887 (N_17887,N_17083,N_17048);
nor U17888 (N_17888,N_17430,N_17380);
nor U17889 (N_17889,N_17291,N_17128);
or U17890 (N_17890,N_17063,N_17327);
nand U17891 (N_17891,N_17078,N_17356);
nand U17892 (N_17892,N_17220,N_17139);
and U17893 (N_17893,N_17337,N_17300);
nand U17894 (N_17894,N_17178,N_17140);
or U17895 (N_17895,N_17080,N_17088);
or U17896 (N_17896,N_17384,N_17324);
xnor U17897 (N_17897,N_17475,N_17330);
or U17898 (N_17898,N_17017,N_17354);
xor U17899 (N_17899,N_17279,N_17045);
or U17900 (N_17900,N_17252,N_17343);
or U17901 (N_17901,N_17237,N_17102);
or U17902 (N_17902,N_17436,N_17127);
or U17903 (N_17903,N_17389,N_17354);
or U17904 (N_17904,N_17492,N_17005);
nand U17905 (N_17905,N_17330,N_17043);
nor U17906 (N_17906,N_17199,N_17174);
and U17907 (N_17907,N_17352,N_17126);
and U17908 (N_17908,N_17008,N_17113);
nand U17909 (N_17909,N_17257,N_17369);
nand U17910 (N_17910,N_17492,N_17249);
nand U17911 (N_17911,N_17106,N_17351);
xor U17912 (N_17912,N_17027,N_17074);
xnor U17913 (N_17913,N_17189,N_17335);
and U17914 (N_17914,N_17021,N_17074);
and U17915 (N_17915,N_17090,N_17353);
or U17916 (N_17916,N_17002,N_17115);
or U17917 (N_17917,N_17309,N_17185);
and U17918 (N_17918,N_17206,N_17306);
xor U17919 (N_17919,N_17499,N_17195);
or U17920 (N_17920,N_17072,N_17435);
and U17921 (N_17921,N_17161,N_17206);
nand U17922 (N_17922,N_17357,N_17177);
nor U17923 (N_17923,N_17135,N_17452);
nor U17924 (N_17924,N_17237,N_17247);
or U17925 (N_17925,N_17284,N_17021);
xor U17926 (N_17926,N_17094,N_17198);
and U17927 (N_17927,N_17313,N_17209);
xnor U17928 (N_17928,N_17400,N_17353);
nand U17929 (N_17929,N_17048,N_17165);
or U17930 (N_17930,N_17060,N_17201);
nand U17931 (N_17931,N_17312,N_17158);
nor U17932 (N_17932,N_17345,N_17195);
xnor U17933 (N_17933,N_17159,N_17189);
nor U17934 (N_17934,N_17288,N_17313);
nor U17935 (N_17935,N_17084,N_17266);
or U17936 (N_17936,N_17223,N_17485);
nor U17937 (N_17937,N_17312,N_17255);
nor U17938 (N_17938,N_17159,N_17039);
nor U17939 (N_17939,N_17091,N_17121);
and U17940 (N_17940,N_17221,N_17409);
and U17941 (N_17941,N_17148,N_17458);
and U17942 (N_17942,N_17359,N_17379);
or U17943 (N_17943,N_17027,N_17012);
or U17944 (N_17944,N_17469,N_17090);
nor U17945 (N_17945,N_17151,N_17315);
or U17946 (N_17946,N_17074,N_17208);
nand U17947 (N_17947,N_17432,N_17279);
or U17948 (N_17948,N_17091,N_17208);
xor U17949 (N_17949,N_17228,N_17010);
xor U17950 (N_17950,N_17375,N_17359);
or U17951 (N_17951,N_17172,N_17499);
or U17952 (N_17952,N_17282,N_17007);
nor U17953 (N_17953,N_17412,N_17139);
nor U17954 (N_17954,N_17013,N_17426);
nand U17955 (N_17955,N_17436,N_17213);
or U17956 (N_17956,N_17012,N_17173);
or U17957 (N_17957,N_17428,N_17058);
or U17958 (N_17958,N_17018,N_17240);
nor U17959 (N_17959,N_17045,N_17167);
or U17960 (N_17960,N_17006,N_17484);
nand U17961 (N_17961,N_17048,N_17449);
nand U17962 (N_17962,N_17435,N_17131);
nor U17963 (N_17963,N_17110,N_17219);
nor U17964 (N_17964,N_17365,N_17062);
xnor U17965 (N_17965,N_17211,N_17190);
or U17966 (N_17966,N_17015,N_17211);
nand U17967 (N_17967,N_17049,N_17082);
xor U17968 (N_17968,N_17148,N_17193);
and U17969 (N_17969,N_17032,N_17105);
nand U17970 (N_17970,N_17013,N_17103);
and U17971 (N_17971,N_17159,N_17273);
nand U17972 (N_17972,N_17088,N_17206);
or U17973 (N_17973,N_17430,N_17297);
xnor U17974 (N_17974,N_17433,N_17297);
xnor U17975 (N_17975,N_17300,N_17363);
nand U17976 (N_17976,N_17387,N_17209);
nand U17977 (N_17977,N_17257,N_17313);
nor U17978 (N_17978,N_17477,N_17286);
xnor U17979 (N_17979,N_17352,N_17362);
nor U17980 (N_17980,N_17203,N_17154);
or U17981 (N_17981,N_17160,N_17323);
and U17982 (N_17982,N_17068,N_17160);
nand U17983 (N_17983,N_17440,N_17100);
nor U17984 (N_17984,N_17104,N_17263);
nor U17985 (N_17985,N_17485,N_17341);
and U17986 (N_17986,N_17024,N_17221);
or U17987 (N_17987,N_17300,N_17144);
nand U17988 (N_17988,N_17062,N_17082);
xnor U17989 (N_17989,N_17083,N_17068);
nand U17990 (N_17990,N_17464,N_17395);
xor U17991 (N_17991,N_17382,N_17370);
xor U17992 (N_17992,N_17258,N_17417);
and U17993 (N_17993,N_17092,N_17255);
nand U17994 (N_17994,N_17106,N_17453);
and U17995 (N_17995,N_17041,N_17025);
nor U17996 (N_17996,N_17278,N_17302);
or U17997 (N_17997,N_17169,N_17069);
xor U17998 (N_17998,N_17252,N_17193);
or U17999 (N_17999,N_17475,N_17199);
or U18000 (N_18000,N_17769,N_17954);
or U18001 (N_18001,N_17902,N_17931);
xor U18002 (N_18002,N_17590,N_17539);
nor U18003 (N_18003,N_17973,N_17523);
xnor U18004 (N_18004,N_17659,N_17983);
or U18005 (N_18005,N_17682,N_17649);
nor U18006 (N_18006,N_17504,N_17640);
xor U18007 (N_18007,N_17577,N_17570);
nand U18008 (N_18008,N_17971,N_17788);
and U18009 (N_18009,N_17636,N_17595);
and U18010 (N_18010,N_17987,N_17917);
xor U18011 (N_18011,N_17869,N_17687);
nor U18012 (N_18012,N_17882,N_17540);
or U18013 (N_18013,N_17667,N_17646);
nand U18014 (N_18014,N_17740,N_17952);
nor U18015 (N_18015,N_17618,N_17516);
nand U18016 (N_18016,N_17819,N_17778);
xor U18017 (N_18017,N_17849,N_17858);
nor U18018 (N_18018,N_17548,N_17889);
nand U18019 (N_18019,N_17665,N_17745);
nand U18020 (N_18020,N_17519,N_17761);
and U18021 (N_18021,N_17837,N_17921);
or U18022 (N_18022,N_17907,N_17890);
nor U18023 (N_18023,N_17505,N_17965);
or U18024 (N_18024,N_17828,N_17552);
nand U18025 (N_18025,N_17768,N_17589);
or U18026 (N_18026,N_17868,N_17502);
nand U18027 (N_18027,N_17574,N_17556);
and U18028 (N_18028,N_17978,N_17863);
xor U18029 (N_18029,N_17753,N_17597);
nand U18030 (N_18030,N_17672,N_17859);
or U18031 (N_18031,N_17822,N_17609);
xor U18032 (N_18032,N_17695,N_17919);
xor U18033 (N_18033,N_17836,N_17898);
and U18034 (N_18034,N_17573,N_17885);
or U18035 (N_18035,N_17628,N_17817);
or U18036 (N_18036,N_17500,N_17830);
nor U18037 (N_18037,N_17801,N_17766);
nor U18038 (N_18038,N_17566,N_17881);
nand U18039 (N_18039,N_17661,N_17959);
nand U18040 (N_18040,N_17976,N_17823);
nor U18041 (N_18041,N_17873,N_17941);
nand U18042 (N_18042,N_17606,N_17707);
or U18043 (N_18043,N_17642,N_17758);
xnor U18044 (N_18044,N_17880,N_17664);
nor U18045 (N_18045,N_17694,N_17564);
nand U18046 (N_18046,N_17692,N_17608);
or U18047 (N_18047,N_17936,N_17816);
nand U18048 (N_18048,N_17621,N_17841);
xor U18049 (N_18049,N_17551,N_17612);
nand U18050 (N_18050,N_17793,N_17782);
nand U18051 (N_18051,N_17910,N_17512);
or U18052 (N_18052,N_17584,N_17704);
nor U18053 (N_18053,N_17940,N_17576);
nor U18054 (N_18054,N_17526,N_17767);
or U18055 (N_18055,N_17772,N_17805);
nor U18056 (N_18056,N_17698,N_17908);
nand U18057 (N_18057,N_17585,N_17645);
or U18058 (N_18058,N_17939,N_17755);
nor U18059 (N_18059,N_17815,N_17770);
or U18060 (N_18060,N_17938,N_17538);
nor U18061 (N_18061,N_17722,N_17529);
and U18062 (N_18062,N_17729,N_17688);
and U18063 (N_18063,N_17583,N_17776);
xnor U18064 (N_18064,N_17581,N_17660);
nand U18065 (N_18065,N_17797,N_17998);
nor U18066 (N_18066,N_17958,N_17943);
or U18067 (N_18067,N_17619,N_17629);
xnor U18068 (N_18068,N_17951,N_17721);
and U18069 (N_18069,N_17671,N_17835);
or U18070 (N_18070,N_17746,N_17634);
xnor U18071 (N_18071,N_17598,N_17826);
and U18072 (N_18072,N_17553,N_17541);
nor U18073 (N_18073,N_17732,N_17742);
nand U18074 (N_18074,N_17731,N_17897);
xor U18075 (N_18075,N_17783,N_17710);
and U18076 (N_18076,N_17592,N_17759);
and U18077 (N_18077,N_17903,N_17717);
or U18078 (N_18078,N_17864,N_17860);
xor U18079 (N_18079,N_17567,N_17674);
or U18080 (N_18080,N_17680,N_17794);
or U18081 (N_18081,N_17852,N_17879);
or U18082 (N_18082,N_17534,N_17525);
or U18083 (N_18083,N_17508,N_17914);
and U18084 (N_18084,N_17531,N_17637);
and U18085 (N_18085,N_17840,N_17888);
nor U18086 (N_18086,N_17850,N_17571);
nand U18087 (N_18087,N_17586,N_17594);
and U18088 (N_18088,N_17743,N_17773);
or U18089 (N_18089,N_17587,N_17896);
and U18090 (N_18090,N_17599,N_17503);
nor U18091 (N_18091,N_17994,N_17763);
or U18092 (N_18092,N_17984,N_17506);
xnor U18093 (N_18093,N_17517,N_17803);
and U18094 (N_18094,N_17878,N_17616);
or U18095 (N_18095,N_17832,N_17611);
nor U18096 (N_18096,N_17558,N_17877);
xnor U18097 (N_18097,N_17666,N_17510);
nand U18098 (N_18098,N_17668,N_17865);
nand U18099 (N_18099,N_17930,N_17949);
xnor U18100 (N_18100,N_17774,N_17686);
or U18101 (N_18101,N_17867,N_17604);
and U18102 (N_18102,N_17806,N_17675);
nand U18103 (N_18103,N_17990,N_17588);
or U18104 (N_18104,N_17739,N_17607);
nand U18105 (N_18105,N_17663,N_17824);
nand U18106 (N_18106,N_17677,N_17968);
nand U18107 (N_18107,N_17992,N_17886);
or U18108 (N_18108,N_17617,N_17762);
or U18109 (N_18109,N_17927,N_17545);
nand U18110 (N_18110,N_17969,N_17623);
nand U18111 (N_18111,N_17689,N_17981);
nand U18112 (N_18112,N_17842,N_17827);
and U18113 (N_18113,N_17808,N_17834);
and U18114 (N_18114,N_17575,N_17513);
or U18115 (N_18115,N_17653,N_17676);
and U18116 (N_18116,N_17765,N_17596);
or U18117 (N_18117,N_17874,N_17546);
and U18118 (N_18118,N_17855,N_17866);
and U18119 (N_18119,N_17802,N_17833);
nand U18120 (N_18120,N_17565,N_17955);
nor U18121 (N_18121,N_17848,N_17635);
nor U18122 (N_18122,N_17844,N_17651);
and U18123 (N_18123,N_17542,N_17647);
nand U18124 (N_18124,N_17738,N_17932);
and U18125 (N_18125,N_17970,N_17964);
and U18126 (N_18126,N_17948,N_17935);
or U18127 (N_18127,N_17925,N_17920);
nand U18128 (N_18128,N_17718,N_17963);
nor U18129 (N_18129,N_17654,N_17726);
and U18130 (N_18130,N_17875,N_17754);
nand U18131 (N_18131,N_17899,N_17533);
or U18132 (N_18132,N_17799,N_17893);
or U18133 (N_18133,N_17701,N_17625);
nor U18134 (N_18134,N_17792,N_17554);
or U18135 (N_18135,N_17632,N_17967);
xor U18136 (N_18136,N_17652,N_17580);
nor U18137 (N_18137,N_17934,N_17989);
and U18138 (N_18138,N_17961,N_17872);
nor U18139 (N_18139,N_17901,N_17702);
or U18140 (N_18140,N_17904,N_17536);
nand U18141 (N_18141,N_17501,N_17887);
and U18142 (N_18142,N_17800,N_17795);
nor U18143 (N_18143,N_17957,N_17557);
nand U18144 (N_18144,N_17915,N_17735);
xnor U18145 (N_18145,N_17627,N_17781);
nand U18146 (N_18146,N_17749,N_17857);
or U18147 (N_18147,N_17995,N_17514);
nand U18148 (N_18148,N_17991,N_17693);
xor U18149 (N_18149,N_17549,N_17518);
and U18150 (N_18150,N_17861,N_17714);
nor U18151 (N_18151,N_17535,N_17928);
or U18152 (N_18152,N_17979,N_17856);
nor U18153 (N_18153,N_17561,N_17560);
xor U18154 (N_18154,N_17945,N_17829);
nand U18155 (N_18155,N_17633,N_17751);
nand U18156 (N_18156,N_17960,N_17725);
nor U18157 (N_18157,N_17650,N_17747);
and U18158 (N_18158,N_17527,N_17602);
xor U18159 (N_18159,N_17734,N_17839);
nor U18160 (N_18160,N_17854,N_17699);
and U18161 (N_18161,N_17736,N_17831);
or U18162 (N_18162,N_17658,N_17923);
xor U18163 (N_18163,N_17522,N_17911);
and U18164 (N_18164,N_17891,N_17764);
and U18165 (N_18165,N_17809,N_17787);
and U18166 (N_18166,N_17511,N_17657);
or U18167 (N_18167,N_17845,N_17741);
nand U18168 (N_18168,N_17985,N_17784);
xnor U18169 (N_18169,N_17723,N_17638);
and U18170 (N_18170,N_17709,N_17543);
xor U18171 (N_18171,N_17988,N_17733);
nor U18172 (N_18172,N_17644,N_17563);
nand U18173 (N_18173,N_17670,N_17982);
xnor U18174 (N_18174,N_17613,N_17777);
and U18175 (N_18175,N_17748,N_17798);
or U18176 (N_18176,N_17821,N_17922);
nor U18177 (N_18177,N_17853,N_17700);
or U18178 (N_18178,N_17813,N_17509);
xor U18179 (N_18179,N_17532,N_17683);
nand U18180 (N_18180,N_17946,N_17847);
nor U18181 (N_18181,N_17883,N_17520);
nor U18182 (N_18182,N_17814,N_17953);
and U18183 (N_18183,N_17744,N_17622);
or U18184 (N_18184,N_17942,N_17944);
nor U18185 (N_18185,N_17624,N_17906);
xnor U18186 (N_18186,N_17547,N_17825);
or U18187 (N_18187,N_17591,N_17912);
nand U18188 (N_18188,N_17789,N_17843);
or U18189 (N_18189,N_17870,N_17615);
nand U18190 (N_18190,N_17977,N_17791);
xnor U18191 (N_18191,N_17641,N_17630);
or U18192 (N_18192,N_17892,N_17876);
and U18193 (N_18193,N_17924,N_17804);
xor U18194 (N_18194,N_17913,N_17697);
xor U18195 (N_18195,N_17610,N_17708);
or U18196 (N_18196,N_17956,N_17926);
xnor U18197 (N_18197,N_17673,N_17719);
or U18198 (N_18198,N_17796,N_17706);
and U18199 (N_18199,N_17681,N_17655);
xor U18200 (N_18200,N_17895,N_17662);
and U18201 (N_18201,N_17605,N_17997);
or U18202 (N_18202,N_17996,N_17716);
xor U18203 (N_18203,N_17684,N_17713);
or U18204 (N_18204,N_17947,N_17620);
nor U18205 (N_18205,N_17785,N_17728);
or U18206 (N_18206,N_17593,N_17559);
or U18207 (N_18207,N_17550,N_17750);
nor U18208 (N_18208,N_17614,N_17568);
or U18209 (N_18209,N_17918,N_17810);
nand U18210 (N_18210,N_17555,N_17929);
nand U18211 (N_18211,N_17937,N_17752);
nand U18212 (N_18212,N_17528,N_17669);
or U18213 (N_18213,N_17578,N_17537);
or U18214 (N_18214,N_17838,N_17724);
and U18215 (N_18215,N_17656,N_17603);
or U18216 (N_18216,N_17712,N_17962);
nand U18217 (N_18217,N_17703,N_17639);
nor U18218 (N_18218,N_17779,N_17786);
and U18219 (N_18219,N_17900,N_17507);
xnor U18220 (N_18220,N_17685,N_17648);
or U18221 (N_18221,N_17980,N_17679);
or U18222 (N_18222,N_17999,N_17757);
or U18223 (N_18223,N_17975,N_17760);
xnor U18224 (N_18224,N_17909,N_17544);
nand U18225 (N_18225,N_17771,N_17790);
and U18226 (N_18226,N_17530,N_17524);
xor U18227 (N_18227,N_17933,N_17811);
xor U18228 (N_18228,N_17950,N_17905);
nor U18229 (N_18229,N_17569,N_17851);
xor U18230 (N_18230,N_17572,N_17894);
nand U18231 (N_18231,N_17986,N_17626);
nand U18232 (N_18232,N_17862,N_17972);
nand U18233 (N_18233,N_17720,N_17582);
xor U18234 (N_18234,N_17756,N_17705);
xor U18235 (N_18235,N_17807,N_17727);
and U18236 (N_18236,N_17521,N_17715);
nor U18237 (N_18237,N_17515,N_17600);
nand U18238 (N_18238,N_17711,N_17775);
xor U18239 (N_18239,N_17974,N_17884);
xnor U18240 (N_18240,N_17820,N_17818);
or U18241 (N_18241,N_17871,N_17643);
or U18242 (N_18242,N_17631,N_17562);
and U18243 (N_18243,N_17737,N_17696);
nand U18244 (N_18244,N_17846,N_17601);
nand U18245 (N_18245,N_17966,N_17691);
xnor U18246 (N_18246,N_17690,N_17812);
nand U18247 (N_18247,N_17730,N_17993);
nor U18248 (N_18248,N_17780,N_17916);
nor U18249 (N_18249,N_17678,N_17579);
nor U18250 (N_18250,N_17518,N_17947);
nand U18251 (N_18251,N_17567,N_17652);
xnor U18252 (N_18252,N_17543,N_17587);
and U18253 (N_18253,N_17629,N_17564);
nor U18254 (N_18254,N_17764,N_17883);
nand U18255 (N_18255,N_17920,N_17684);
and U18256 (N_18256,N_17974,N_17759);
or U18257 (N_18257,N_17589,N_17968);
nand U18258 (N_18258,N_17707,N_17988);
nand U18259 (N_18259,N_17679,N_17785);
and U18260 (N_18260,N_17570,N_17860);
nor U18261 (N_18261,N_17607,N_17539);
or U18262 (N_18262,N_17854,N_17690);
and U18263 (N_18263,N_17795,N_17569);
xnor U18264 (N_18264,N_17557,N_17554);
and U18265 (N_18265,N_17887,N_17965);
nand U18266 (N_18266,N_17645,N_17532);
and U18267 (N_18267,N_17536,N_17751);
xnor U18268 (N_18268,N_17518,N_17599);
nand U18269 (N_18269,N_17680,N_17561);
or U18270 (N_18270,N_17925,N_17689);
nor U18271 (N_18271,N_17914,N_17722);
nor U18272 (N_18272,N_17566,N_17797);
xor U18273 (N_18273,N_17508,N_17741);
nor U18274 (N_18274,N_17877,N_17907);
and U18275 (N_18275,N_17841,N_17724);
xor U18276 (N_18276,N_17557,N_17696);
and U18277 (N_18277,N_17712,N_17934);
xnor U18278 (N_18278,N_17772,N_17521);
and U18279 (N_18279,N_17607,N_17813);
and U18280 (N_18280,N_17975,N_17921);
nor U18281 (N_18281,N_17942,N_17855);
and U18282 (N_18282,N_17944,N_17546);
nor U18283 (N_18283,N_17886,N_17572);
and U18284 (N_18284,N_17848,N_17720);
nand U18285 (N_18285,N_17681,N_17923);
and U18286 (N_18286,N_17616,N_17767);
nor U18287 (N_18287,N_17737,N_17560);
xor U18288 (N_18288,N_17844,N_17946);
or U18289 (N_18289,N_17987,N_17698);
nor U18290 (N_18290,N_17984,N_17629);
and U18291 (N_18291,N_17638,N_17759);
nor U18292 (N_18292,N_17816,N_17572);
nand U18293 (N_18293,N_17596,N_17544);
and U18294 (N_18294,N_17999,N_17578);
nor U18295 (N_18295,N_17824,N_17612);
xnor U18296 (N_18296,N_17654,N_17834);
nand U18297 (N_18297,N_17809,N_17909);
xnor U18298 (N_18298,N_17711,N_17687);
or U18299 (N_18299,N_17777,N_17881);
nand U18300 (N_18300,N_17573,N_17794);
nor U18301 (N_18301,N_17562,N_17651);
nand U18302 (N_18302,N_17850,N_17747);
or U18303 (N_18303,N_17934,N_17839);
xor U18304 (N_18304,N_17542,N_17727);
and U18305 (N_18305,N_17816,N_17834);
nand U18306 (N_18306,N_17990,N_17985);
xnor U18307 (N_18307,N_17697,N_17857);
nand U18308 (N_18308,N_17621,N_17954);
and U18309 (N_18309,N_17538,N_17790);
nand U18310 (N_18310,N_17986,N_17937);
nand U18311 (N_18311,N_17824,N_17771);
and U18312 (N_18312,N_17737,N_17672);
nor U18313 (N_18313,N_17722,N_17692);
and U18314 (N_18314,N_17703,N_17986);
or U18315 (N_18315,N_17745,N_17738);
nor U18316 (N_18316,N_17816,N_17900);
or U18317 (N_18317,N_17787,N_17646);
or U18318 (N_18318,N_17670,N_17809);
or U18319 (N_18319,N_17852,N_17660);
or U18320 (N_18320,N_17718,N_17653);
or U18321 (N_18321,N_17688,N_17799);
xnor U18322 (N_18322,N_17520,N_17617);
nand U18323 (N_18323,N_17623,N_17958);
nor U18324 (N_18324,N_17522,N_17711);
nor U18325 (N_18325,N_17748,N_17902);
nand U18326 (N_18326,N_17902,N_17566);
nand U18327 (N_18327,N_17839,N_17535);
nand U18328 (N_18328,N_17812,N_17781);
and U18329 (N_18329,N_17598,N_17861);
or U18330 (N_18330,N_17616,N_17796);
xor U18331 (N_18331,N_17852,N_17850);
or U18332 (N_18332,N_17792,N_17848);
xor U18333 (N_18333,N_17858,N_17640);
and U18334 (N_18334,N_17996,N_17566);
nor U18335 (N_18335,N_17883,N_17509);
xnor U18336 (N_18336,N_17965,N_17500);
and U18337 (N_18337,N_17993,N_17970);
nand U18338 (N_18338,N_17781,N_17679);
nor U18339 (N_18339,N_17907,N_17586);
nor U18340 (N_18340,N_17721,N_17713);
xnor U18341 (N_18341,N_17741,N_17656);
nor U18342 (N_18342,N_17909,N_17619);
nor U18343 (N_18343,N_17698,N_17950);
nand U18344 (N_18344,N_17697,N_17868);
and U18345 (N_18345,N_17671,N_17928);
nor U18346 (N_18346,N_17895,N_17943);
xnor U18347 (N_18347,N_17949,N_17942);
nand U18348 (N_18348,N_17774,N_17685);
and U18349 (N_18349,N_17796,N_17640);
or U18350 (N_18350,N_17856,N_17578);
and U18351 (N_18351,N_17601,N_17692);
nand U18352 (N_18352,N_17856,N_17558);
or U18353 (N_18353,N_17773,N_17507);
nand U18354 (N_18354,N_17661,N_17926);
nor U18355 (N_18355,N_17873,N_17915);
and U18356 (N_18356,N_17828,N_17946);
xor U18357 (N_18357,N_17694,N_17870);
nor U18358 (N_18358,N_17866,N_17512);
and U18359 (N_18359,N_17530,N_17790);
or U18360 (N_18360,N_17839,N_17656);
or U18361 (N_18361,N_17857,N_17910);
nor U18362 (N_18362,N_17905,N_17887);
nor U18363 (N_18363,N_17768,N_17711);
nand U18364 (N_18364,N_17662,N_17897);
nand U18365 (N_18365,N_17767,N_17989);
or U18366 (N_18366,N_17777,N_17601);
or U18367 (N_18367,N_17865,N_17535);
xor U18368 (N_18368,N_17955,N_17814);
or U18369 (N_18369,N_17645,N_17842);
or U18370 (N_18370,N_17503,N_17954);
nor U18371 (N_18371,N_17713,N_17503);
xnor U18372 (N_18372,N_17744,N_17734);
and U18373 (N_18373,N_17856,N_17905);
and U18374 (N_18374,N_17626,N_17677);
and U18375 (N_18375,N_17844,N_17629);
and U18376 (N_18376,N_17850,N_17920);
or U18377 (N_18377,N_17687,N_17617);
nor U18378 (N_18378,N_17535,N_17644);
nor U18379 (N_18379,N_17545,N_17887);
or U18380 (N_18380,N_17671,N_17709);
nor U18381 (N_18381,N_17549,N_17761);
nor U18382 (N_18382,N_17572,N_17752);
or U18383 (N_18383,N_17854,N_17868);
and U18384 (N_18384,N_17666,N_17776);
and U18385 (N_18385,N_17604,N_17853);
and U18386 (N_18386,N_17583,N_17719);
xnor U18387 (N_18387,N_17508,N_17519);
xnor U18388 (N_18388,N_17721,N_17764);
and U18389 (N_18389,N_17558,N_17591);
and U18390 (N_18390,N_17906,N_17815);
or U18391 (N_18391,N_17564,N_17728);
and U18392 (N_18392,N_17523,N_17974);
nand U18393 (N_18393,N_17849,N_17732);
or U18394 (N_18394,N_17965,N_17524);
or U18395 (N_18395,N_17653,N_17668);
nor U18396 (N_18396,N_17560,N_17538);
or U18397 (N_18397,N_17822,N_17687);
nand U18398 (N_18398,N_17572,N_17581);
or U18399 (N_18399,N_17721,N_17820);
and U18400 (N_18400,N_17910,N_17786);
and U18401 (N_18401,N_17751,N_17824);
nand U18402 (N_18402,N_17947,N_17905);
nand U18403 (N_18403,N_17586,N_17542);
nand U18404 (N_18404,N_17696,N_17781);
nand U18405 (N_18405,N_17888,N_17959);
and U18406 (N_18406,N_17997,N_17527);
and U18407 (N_18407,N_17815,N_17709);
xor U18408 (N_18408,N_17862,N_17579);
nor U18409 (N_18409,N_17733,N_17625);
nand U18410 (N_18410,N_17566,N_17863);
nor U18411 (N_18411,N_17976,N_17877);
or U18412 (N_18412,N_17952,N_17943);
nand U18413 (N_18413,N_17763,N_17536);
or U18414 (N_18414,N_17951,N_17641);
xnor U18415 (N_18415,N_17552,N_17762);
nor U18416 (N_18416,N_17729,N_17875);
nand U18417 (N_18417,N_17974,N_17644);
and U18418 (N_18418,N_17866,N_17632);
nand U18419 (N_18419,N_17942,N_17794);
xor U18420 (N_18420,N_17934,N_17674);
nor U18421 (N_18421,N_17954,N_17915);
xor U18422 (N_18422,N_17921,N_17656);
and U18423 (N_18423,N_17702,N_17771);
and U18424 (N_18424,N_17717,N_17632);
xnor U18425 (N_18425,N_17557,N_17669);
nor U18426 (N_18426,N_17624,N_17604);
or U18427 (N_18427,N_17856,N_17830);
xnor U18428 (N_18428,N_17620,N_17763);
xor U18429 (N_18429,N_17527,N_17575);
or U18430 (N_18430,N_17736,N_17961);
nor U18431 (N_18431,N_17878,N_17786);
xor U18432 (N_18432,N_17693,N_17778);
xnor U18433 (N_18433,N_17607,N_17515);
and U18434 (N_18434,N_17759,N_17743);
or U18435 (N_18435,N_17585,N_17822);
and U18436 (N_18436,N_17803,N_17846);
or U18437 (N_18437,N_17741,N_17919);
nand U18438 (N_18438,N_17614,N_17583);
or U18439 (N_18439,N_17623,N_17927);
nand U18440 (N_18440,N_17861,N_17715);
nand U18441 (N_18441,N_17797,N_17530);
xor U18442 (N_18442,N_17523,N_17610);
xor U18443 (N_18443,N_17906,N_17943);
nor U18444 (N_18444,N_17629,N_17676);
and U18445 (N_18445,N_17886,N_17756);
nor U18446 (N_18446,N_17890,N_17709);
or U18447 (N_18447,N_17635,N_17788);
nand U18448 (N_18448,N_17588,N_17855);
or U18449 (N_18449,N_17802,N_17765);
nor U18450 (N_18450,N_17769,N_17966);
xor U18451 (N_18451,N_17891,N_17763);
and U18452 (N_18452,N_17545,N_17845);
and U18453 (N_18453,N_17902,N_17550);
xnor U18454 (N_18454,N_17949,N_17843);
or U18455 (N_18455,N_17781,N_17928);
nor U18456 (N_18456,N_17752,N_17948);
nor U18457 (N_18457,N_17948,N_17642);
xor U18458 (N_18458,N_17555,N_17656);
nor U18459 (N_18459,N_17547,N_17716);
xnor U18460 (N_18460,N_17558,N_17765);
nor U18461 (N_18461,N_17696,N_17753);
nand U18462 (N_18462,N_17955,N_17612);
or U18463 (N_18463,N_17541,N_17641);
xor U18464 (N_18464,N_17631,N_17828);
nor U18465 (N_18465,N_17673,N_17831);
nand U18466 (N_18466,N_17848,N_17721);
and U18467 (N_18467,N_17654,N_17680);
nand U18468 (N_18468,N_17973,N_17601);
or U18469 (N_18469,N_17715,N_17695);
nand U18470 (N_18470,N_17843,N_17751);
or U18471 (N_18471,N_17966,N_17858);
xor U18472 (N_18472,N_17699,N_17667);
nand U18473 (N_18473,N_17534,N_17828);
xor U18474 (N_18474,N_17704,N_17750);
or U18475 (N_18475,N_17959,N_17641);
xnor U18476 (N_18476,N_17512,N_17875);
or U18477 (N_18477,N_17509,N_17954);
nor U18478 (N_18478,N_17675,N_17785);
nand U18479 (N_18479,N_17682,N_17908);
and U18480 (N_18480,N_17806,N_17835);
nor U18481 (N_18481,N_17780,N_17784);
nand U18482 (N_18482,N_17845,N_17929);
or U18483 (N_18483,N_17528,N_17612);
xnor U18484 (N_18484,N_17602,N_17655);
nor U18485 (N_18485,N_17842,N_17933);
xor U18486 (N_18486,N_17815,N_17910);
nor U18487 (N_18487,N_17808,N_17661);
xnor U18488 (N_18488,N_17524,N_17628);
or U18489 (N_18489,N_17812,N_17543);
and U18490 (N_18490,N_17676,N_17504);
or U18491 (N_18491,N_17888,N_17519);
or U18492 (N_18492,N_17943,N_17768);
nand U18493 (N_18493,N_17857,N_17792);
nand U18494 (N_18494,N_17909,N_17620);
nand U18495 (N_18495,N_17605,N_17510);
xor U18496 (N_18496,N_17910,N_17776);
nand U18497 (N_18497,N_17976,N_17960);
nor U18498 (N_18498,N_17734,N_17658);
nor U18499 (N_18499,N_17569,N_17612);
or U18500 (N_18500,N_18219,N_18101);
or U18501 (N_18501,N_18440,N_18343);
or U18502 (N_18502,N_18346,N_18194);
nand U18503 (N_18503,N_18102,N_18381);
and U18504 (N_18504,N_18248,N_18311);
nor U18505 (N_18505,N_18286,N_18023);
nand U18506 (N_18506,N_18062,N_18133);
and U18507 (N_18507,N_18277,N_18378);
xor U18508 (N_18508,N_18146,N_18353);
xnor U18509 (N_18509,N_18114,N_18349);
nand U18510 (N_18510,N_18425,N_18005);
and U18511 (N_18511,N_18070,N_18384);
and U18512 (N_18512,N_18010,N_18270);
nor U18513 (N_18513,N_18234,N_18181);
xor U18514 (N_18514,N_18161,N_18116);
xor U18515 (N_18515,N_18095,N_18345);
or U18516 (N_18516,N_18153,N_18058);
nand U18517 (N_18517,N_18092,N_18294);
nand U18518 (N_18518,N_18409,N_18035);
xor U18519 (N_18519,N_18064,N_18249);
and U18520 (N_18520,N_18229,N_18469);
or U18521 (N_18521,N_18218,N_18278);
nor U18522 (N_18522,N_18269,N_18486);
nor U18523 (N_18523,N_18372,N_18403);
or U18524 (N_18524,N_18006,N_18251);
nand U18525 (N_18525,N_18257,N_18460);
nor U18526 (N_18526,N_18106,N_18208);
nor U18527 (N_18527,N_18496,N_18475);
nor U18528 (N_18528,N_18029,N_18088);
xor U18529 (N_18529,N_18198,N_18163);
nand U18530 (N_18530,N_18437,N_18491);
or U18531 (N_18531,N_18043,N_18336);
and U18532 (N_18532,N_18463,N_18109);
nand U18533 (N_18533,N_18412,N_18283);
or U18534 (N_18534,N_18148,N_18124);
xnor U18535 (N_18535,N_18018,N_18150);
and U18536 (N_18536,N_18295,N_18305);
nand U18537 (N_18537,N_18388,N_18472);
and U18538 (N_18538,N_18480,N_18279);
xnor U18539 (N_18539,N_18433,N_18104);
nand U18540 (N_18540,N_18099,N_18021);
nand U18541 (N_18541,N_18326,N_18155);
xnor U18542 (N_18542,N_18327,N_18159);
nor U18543 (N_18543,N_18237,N_18459);
nor U18544 (N_18544,N_18306,N_18105);
or U18545 (N_18545,N_18351,N_18436);
xor U18546 (N_18546,N_18090,N_18377);
and U18547 (N_18547,N_18032,N_18273);
or U18548 (N_18548,N_18337,N_18189);
or U18549 (N_18549,N_18037,N_18074);
nand U18550 (N_18550,N_18495,N_18031);
nor U18551 (N_18551,N_18199,N_18158);
and U18552 (N_18552,N_18320,N_18473);
nand U18553 (N_18553,N_18331,N_18493);
and U18554 (N_18554,N_18003,N_18113);
nand U18555 (N_18555,N_18185,N_18197);
xnor U18556 (N_18556,N_18182,N_18147);
nor U18557 (N_18557,N_18135,N_18250);
nand U18558 (N_18558,N_18445,N_18324);
and U18559 (N_18559,N_18256,N_18371);
or U18560 (N_18560,N_18126,N_18276);
or U18561 (N_18561,N_18120,N_18167);
xnor U18562 (N_18562,N_18028,N_18030);
and U18563 (N_18563,N_18223,N_18117);
xor U18564 (N_18564,N_18338,N_18494);
nand U18565 (N_18565,N_18414,N_18369);
or U18566 (N_18566,N_18464,N_18390);
and U18567 (N_18567,N_18143,N_18456);
or U18568 (N_18568,N_18477,N_18179);
nand U18569 (N_18569,N_18356,N_18471);
and U18570 (N_18570,N_18368,N_18288);
xor U18571 (N_18571,N_18332,N_18044);
xor U18572 (N_18572,N_18290,N_18373);
or U18573 (N_18573,N_18103,N_18141);
and U18574 (N_18574,N_18068,N_18292);
nand U18575 (N_18575,N_18211,N_18057);
xnor U18576 (N_18576,N_18266,N_18089);
nand U18577 (N_18577,N_18022,N_18200);
nand U18578 (N_18578,N_18246,N_18393);
xnor U18579 (N_18579,N_18174,N_18192);
and U18580 (N_18580,N_18342,N_18479);
or U18581 (N_18581,N_18206,N_18461);
and U18582 (N_18582,N_18404,N_18056);
xnor U18583 (N_18583,N_18221,N_18415);
nand U18584 (N_18584,N_18462,N_18448);
nand U18585 (N_18585,N_18275,N_18304);
nor U18586 (N_18586,N_18291,N_18334);
nor U18587 (N_18587,N_18217,N_18301);
nor U18588 (N_18588,N_18222,N_18243);
nand U18589 (N_18589,N_18281,N_18367);
or U18590 (N_18590,N_18307,N_18115);
nand U18591 (N_18591,N_18019,N_18067);
nand U18592 (N_18592,N_18341,N_18376);
nor U18593 (N_18593,N_18072,N_18036);
and U18594 (N_18594,N_18386,N_18262);
and U18595 (N_18595,N_18157,N_18204);
or U18596 (N_18596,N_18165,N_18175);
nor U18597 (N_18597,N_18026,N_18258);
nand U18598 (N_18598,N_18357,N_18027);
nor U18599 (N_18599,N_18216,N_18065);
or U18600 (N_18600,N_18407,N_18212);
nor U18601 (N_18601,N_18140,N_18458);
xor U18602 (N_18602,N_18060,N_18100);
nand U18603 (N_18603,N_18033,N_18050);
and U18604 (N_18604,N_18419,N_18400);
or U18605 (N_18605,N_18255,N_18202);
and U18606 (N_18606,N_18394,N_18323);
nor U18607 (N_18607,N_18426,N_18122);
or U18608 (N_18608,N_18176,N_18144);
and U18609 (N_18609,N_18498,N_18130);
xor U18610 (N_18610,N_18254,N_18359);
nor U18611 (N_18611,N_18428,N_18466);
or U18612 (N_18612,N_18422,N_18151);
or U18613 (N_18613,N_18398,N_18309);
and U18614 (N_18614,N_18375,N_18240);
nor U18615 (N_18615,N_18438,N_18303);
or U18616 (N_18616,N_18449,N_18055);
or U18617 (N_18617,N_18042,N_18091);
and U18618 (N_18618,N_18228,N_18131);
and U18619 (N_18619,N_18423,N_18118);
or U18620 (N_18620,N_18329,N_18452);
and U18621 (N_18621,N_18396,N_18450);
nor U18622 (N_18622,N_18484,N_18340);
xnor U18623 (N_18623,N_18078,N_18352);
or U18624 (N_18624,N_18354,N_18287);
nand U18625 (N_18625,N_18085,N_18196);
xor U18626 (N_18626,N_18298,N_18024);
and U18627 (N_18627,N_18319,N_18280);
and U18628 (N_18628,N_18271,N_18052);
or U18629 (N_18629,N_18002,N_18007);
nor U18630 (N_18630,N_18402,N_18358);
nand U18631 (N_18631,N_18265,N_18107);
nand U18632 (N_18632,N_18132,N_18061);
nor U18633 (N_18633,N_18008,N_18125);
nand U18634 (N_18634,N_18312,N_18177);
and U18635 (N_18635,N_18186,N_18418);
xor U18636 (N_18636,N_18310,N_18264);
and U18637 (N_18637,N_18049,N_18427);
nand U18638 (N_18638,N_18205,N_18397);
nand U18639 (N_18639,N_18066,N_18039);
and U18640 (N_18640,N_18195,N_18015);
or U18641 (N_18641,N_18284,N_18213);
or U18642 (N_18642,N_18308,N_18134);
nand U18643 (N_18643,N_18227,N_18405);
nor U18644 (N_18644,N_18413,N_18365);
and U18645 (N_18645,N_18098,N_18421);
or U18646 (N_18646,N_18230,N_18434);
nor U18647 (N_18647,N_18017,N_18441);
nor U18648 (N_18648,N_18285,N_18226);
xor U18649 (N_18649,N_18382,N_18207);
or U18650 (N_18650,N_18457,N_18162);
or U18651 (N_18651,N_18333,N_18013);
and U18652 (N_18652,N_18478,N_18063);
xor U18653 (N_18653,N_18239,N_18451);
nand U18654 (N_18654,N_18267,N_18184);
or U18655 (N_18655,N_18083,N_18487);
or U18656 (N_18656,N_18489,N_18499);
nor U18657 (N_18657,N_18000,N_18417);
and U18658 (N_18658,N_18429,N_18096);
nor U18659 (N_18659,N_18314,N_18241);
and U18660 (N_18660,N_18317,N_18380);
nor U18661 (N_18661,N_18071,N_18047);
xor U18662 (N_18662,N_18087,N_18350);
nor U18663 (N_18663,N_18299,N_18045);
xnor U18664 (N_18664,N_18170,N_18112);
and U18665 (N_18665,N_18242,N_18411);
or U18666 (N_18666,N_18454,N_18416);
nand U18667 (N_18667,N_18391,N_18001);
nand U18668 (N_18668,N_18366,N_18059);
nand U18669 (N_18669,N_18447,N_18051);
nor U18670 (N_18670,N_18046,N_18318);
nor U18671 (N_18671,N_18300,N_18431);
xnor U18672 (N_18672,N_18020,N_18137);
and U18673 (N_18673,N_18444,N_18127);
and U18674 (N_18674,N_18172,N_18224);
nand U18675 (N_18675,N_18203,N_18016);
nor U18676 (N_18676,N_18041,N_18395);
nor U18677 (N_18677,N_18455,N_18481);
xnor U18678 (N_18678,N_18321,N_18316);
nand U18679 (N_18679,N_18123,N_18232);
and U18680 (N_18680,N_18210,N_18344);
nand U18681 (N_18681,N_18453,N_18108);
nor U18682 (N_18682,N_18183,N_18076);
or U18683 (N_18683,N_18328,N_18468);
nor U18684 (N_18684,N_18119,N_18214);
or U18685 (N_18685,N_18335,N_18121);
xnor U18686 (N_18686,N_18011,N_18110);
nand U18687 (N_18687,N_18111,N_18169);
xnor U18688 (N_18688,N_18439,N_18160);
nand U18689 (N_18689,N_18401,N_18152);
or U18690 (N_18690,N_18075,N_18399);
and U18691 (N_18691,N_18164,N_18430);
nor U18692 (N_18692,N_18077,N_18138);
and U18693 (N_18693,N_18355,N_18274);
nor U18694 (N_18694,N_18154,N_18231);
and U18695 (N_18695,N_18236,N_18081);
or U18696 (N_18696,N_18362,N_18410);
nand U18697 (N_18697,N_18424,N_18247);
nand U18698 (N_18698,N_18038,N_18190);
or U18699 (N_18699,N_18053,N_18315);
xor U18700 (N_18700,N_18379,N_18443);
xor U18701 (N_18701,N_18233,N_18173);
nor U18702 (N_18702,N_18476,N_18361);
or U18703 (N_18703,N_18220,N_18296);
nor U18704 (N_18704,N_18289,N_18432);
xor U18705 (N_18705,N_18235,N_18244);
nand U18706 (N_18706,N_18009,N_18313);
nor U18707 (N_18707,N_18209,N_18086);
nand U18708 (N_18708,N_18385,N_18128);
nand U18709 (N_18709,N_18339,N_18259);
and U18710 (N_18710,N_18492,N_18178);
nand U18711 (N_18711,N_18094,N_18082);
or U18712 (N_18712,N_18446,N_18282);
or U18713 (N_18713,N_18187,N_18191);
nor U18714 (N_18714,N_18048,N_18442);
nor U18715 (N_18715,N_18322,N_18215);
and U18716 (N_18716,N_18392,N_18483);
nor U18717 (N_18717,N_18406,N_18168);
and U18718 (N_18718,N_18485,N_18490);
nor U18719 (N_18719,N_18370,N_18383);
nand U18720 (N_18720,N_18347,N_18302);
nor U18721 (N_18721,N_18488,N_18420);
nor U18722 (N_18722,N_18166,N_18004);
and U18723 (N_18723,N_18482,N_18268);
nand U18724 (N_18724,N_18364,N_18054);
and U18725 (N_18725,N_18073,N_18293);
and U18726 (N_18726,N_18079,N_18080);
and U18727 (N_18727,N_18180,N_18139);
or U18728 (N_18728,N_18272,N_18156);
and U18729 (N_18729,N_18389,N_18193);
nand U18730 (N_18730,N_18408,N_18238);
nor U18731 (N_18731,N_18387,N_18136);
nand U18732 (N_18732,N_18012,N_18467);
nor U18733 (N_18733,N_18497,N_18474);
nand U18734 (N_18734,N_18245,N_18097);
nor U18735 (N_18735,N_18069,N_18260);
nor U18736 (N_18736,N_18325,N_18171);
xnor U18737 (N_18737,N_18201,N_18093);
or U18738 (N_18738,N_18145,N_18188);
xor U18739 (N_18739,N_18435,N_18297);
nor U18740 (N_18740,N_18025,N_18149);
nor U18741 (N_18741,N_18142,N_18129);
and U18742 (N_18742,N_18263,N_18363);
nor U18743 (N_18743,N_18225,N_18261);
xor U18744 (N_18744,N_18014,N_18470);
nand U18745 (N_18745,N_18374,N_18330);
nor U18746 (N_18746,N_18252,N_18040);
and U18747 (N_18747,N_18348,N_18465);
nor U18748 (N_18748,N_18084,N_18034);
xor U18749 (N_18749,N_18253,N_18360);
or U18750 (N_18750,N_18031,N_18090);
or U18751 (N_18751,N_18331,N_18244);
xor U18752 (N_18752,N_18427,N_18376);
and U18753 (N_18753,N_18283,N_18112);
and U18754 (N_18754,N_18134,N_18427);
or U18755 (N_18755,N_18317,N_18159);
and U18756 (N_18756,N_18384,N_18079);
nor U18757 (N_18757,N_18242,N_18211);
or U18758 (N_18758,N_18257,N_18148);
and U18759 (N_18759,N_18434,N_18365);
nand U18760 (N_18760,N_18379,N_18175);
nand U18761 (N_18761,N_18466,N_18348);
nand U18762 (N_18762,N_18228,N_18060);
nor U18763 (N_18763,N_18179,N_18488);
xor U18764 (N_18764,N_18364,N_18129);
nor U18765 (N_18765,N_18002,N_18453);
nor U18766 (N_18766,N_18039,N_18246);
xor U18767 (N_18767,N_18038,N_18336);
xor U18768 (N_18768,N_18270,N_18150);
xnor U18769 (N_18769,N_18300,N_18031);
or U18770 (N_18770,N_18310,N_18115);
nor U18771 (N_18771,N_18303,N_18007);
xor U18772 (N_18772,N_18485,N_18018);
or U18773 (N_18773,N_18484,N_18298);
nand U18774 (N_18774,N_18496,N_18398);
xnor U18775 (N_18775,N_18303,N_18262);
or U18776 (N_18776,N_18270,N_18120);
xor U18777 (N_18777,N_18106,N_18447);
or U18778 (N_18778,N_18218,N_18475);
and U18779 (N_18779,N_18340,N_18260);
and U18780 (N_18780,N_18374,N_18444);
nand U18781 (N_18781,N_18171,N_18380);
nand U18782 (N_18782,N_18428,N_18175);
nor U18783 (N_18783,N_18151,N_18499);
xnor U18784 (N_18784,N_18414,N_18205);
nand U18785 (N_18785,N_18447,N_18291);
nand U18786 (N_18786,N_18226,N_18389);
or U18787 (N_18787,N_18444,N_18440);
nor U18788 (N_18788,N_18290,N_18133);
nor U18789 (N_18789,N_18066,N_18160);
or U18790 (N_18790,N_18475,N_18391);
or U18791 (N_18791,N_18439,N_18397);
nand U18792 (N_18792,N_18265,N_18239);
nor U18793 (N_18793,N_18261,N_18324);
and U18794 (N_18794,N_18497,N_18424);
and U18795 (N_18795,N_18006,N_18198);
nor U18796 (N_18796,N_18193,N_18315);
nand U18797 (N_18797,N_18289,N_18268);
xor U18798 (N_18798,N_18009,N_18127);
xor U18799 (N_18799,N_18046,N_18392);
or U18800 (N_18800,N_18424,N_18174);
nor U18801 (N_18801,N_18227,N_18162);
or U18802 (N_18802,N_18131,N_18152);
nand U18803 (N_18803,N_18446,N_18494);
or U18804 (N_18804,N_18479,N_18387);
nand U18805 (N_18805,N_18369,N_18419);
and U18806 (N_18806,N_18450,N_18258);
or U18807 (N_18807,N_18012,N_18498);
nor U18808 (N_18808,N_18011,N_18460);
or U18809 (N_18809,N_18093,N_18367);
nor U18810 (N_18810,N_18028,N_18182);
nand U18811 (N_18811,N_18212,N_18071);
nand U18812 (N_18812,N_18023,N_18331);
or U18813 (N_18813,N_18364,N_18148);
nand U18814 (N_18814,N_18005,N_18251);
or U18815 (N_18815,N_18161,N_18476);
and U18816 (N_18816,N_18087,N_18286);
or U18817 (N_18817,N_18048,N_18086);
nand U18818 (N_18818,N_18017,N_18164);
xor U18819 (N_18819,N_18001,N_18189);
nand U18820 (N_18820,N_18150,N_18417);
or U18821 (N_18821,N_18430,N_18236);
and U18822 (N_18822,N_18047,N_18478);
or U18823 (N_18823,N_18215,N_18083);
nand U18824 (N_18824,N_18237,N_18244);
nand U18825 (N_18825,N_18051,N_18491);
and U18826 (N_18826,N_18145,N_18205);
and U18827 (N_18827,N_18139,N_18193);
nor U18828 (N_18828,N_18495,N_18261);
nor U18829 (N_18829,N_18351,N_18143);
and U18830 (N_18830,N_18330,N_18013);
or U18831 (N_18831,N_18417,N_18457);
nor U18832 (N_18832,N_18180,N_18248);
and U18833 (N_18833,N_18253,N_18015);
and U18834 (N_18834,N_18468,N_18223);
nand U18835 (N_18835,N_18391,N_18083);
and U18836 (N_18836,N_18346,N_18020);
or U18837 (N_18837,N_18226,N_18324);
or U18838 (N_18838,N_18497,N_18423);
nand U18839 (N_18839,N_18467,N_18314);
and U18840 (N_18840,N_18278,N_18248);
and U18841 (N_18841,N_18449,N_18003);
or U18842 (N_18842,N_18466,N_18471);
or U18843 (N_18843,N_18008,N_18175);
and U18844 (N_18844,N_18469,N_18442);
or U18845 (N_18845,N_18219,N_18081);
or U18846 (N_18846,N_18340,N_18068);
xor U18847 (N_18847,N_18033,N_18025);
and U18848 (N_18848,N_18370,N_18448);
nand U18849 (N_18849,N_18261,N_18088);
or U18850 (N_18850,N_18420,N_18453);
xor U18851 (N_18851,N_18309,N_18091);
nor U18852 (N_18852,N_18124,N_18447);
or U18853 (N_18853,N_18295,N_18194);
xor U18854 (N_18854,N_18239,N_18246);
and U18855 (N_18855,N_18372,N_18004);
nand U18856 (N_18856,N_18386,N_18301);
nor U18857 (N_18857,N_18128,N_18450);
nor U18858 (N_18858,N_18069,N_18273);
nor U18859 (N_18859,N_18014,N_18029);
and U18860 (N_18860,N_18215,N_18025);
and U18861 (N_18861,N_18408,N_18319);
and U18862 (N_18862,N_18413,N_18191);
nand U18863 (N_18863,N_18452,N_18435);
xor U18864 (N_18864,N_18366,N_18321);
or U18865 (N_18865,N_18031,N_18210);
xnor U18866 (N_18866,N_18114,N_18080);
nand U18867 (N_18867,N_18263,N_18106);
nor U18868 (N_18868,N_18321,N_18199);
nand U18869 (N_18869,N_18311,N_18230);
nor U18870 (N_18870,N_18246,N_18056);
nand U18871 (N_18871,N_18417,N_18178);
nand U18872 (N_18872,N_18204,N_18225);
xnor U18873 (N_18873,N_18325,N_18228);
nand U18874 (N_18874,N_18057,N_18400);
nand U18875 (N_18875,N_18044,N_18371);
or U18876 (N_18876,N_18425,N_18059);
or U18877 (N_18877,N_18012,N_18488);
and U18878 (N_18878,N_18111,N_18280);
and U18879 (N_18879,N_18148,N_18043);
nand U18880 (N_18880,N_18395,N_18088);
nor U18881 (N_18881,N_18370,N_18026);
nand U18882 (N_18882,N_18064,N_18118);
nand U18883 (N_18883,N_18250,N_18084);
nand U18884 (N_18884,N_18175,N_18197);
nor U18885 (N_18885,N_18261,N_18075);
nor U18886 (N_18886,N_18029,N_18333);
and U18887 (N_18887,N_18043,N_18455);
or U18888 (N_18888,N_18263,N_18059);
nand U18889 (N_18889,N_18074,N_18458);
and U18890 (N_18890,N_18285,N_18246);
xnor U18891 (N_18891,N_18362,N_18125);
nor U18892 (N_18892,N_18280,N_18333);
nor U18893 (N_18893,N_18332,N_18046);
and U18894 (N_18894,N_18430,N_18357);
xor U18895 (N_18895,N_18458,N_18016);
xnor U18896 (N_18896,N_18429,N_18409);
nor U18897 (N_18897,N_18307,N_18346);
nand U18898 (N_18898,N_18218,N_18150);
nand U18899 (N_18899,N_18446,N_18169);
and U18900 (N_18900,N_18408,N_18061);
xor U18901 (N_18901,N_18378,N_18374);
nor U18902 (N_18902,N_18196,N_18017);
nand U18903 (N_18903,N_18285,N_18456);
nor U18904 (N_18904,N_18405,N_18042);
nand U18905 (N_18905,N_18116,N_18465);
xnor U18906 (N_18906,N_18060,N_18138);
xor U18907 (N_18907,N_18285,N_18238);
xor U18908 (N_18908,N_18134,N_18383);
and U18909 (N_18909,N_18235,N_18383);
nand U18910 (N_18910,N_18358,N_18021);
or U18911 (N_18911,N_18468,N_18184);
nor U18912 (N_18912,N_18353,N_18019);
nor U18913 (N_18913,N_18461,N_18495);
nand U18914 (N_18914,N_18212,N_18351);
or U18915 (N_18915,N_18157,N_18192);
or U18916 (N_18916,N_18164,N_18439);
and U18917 (N_18917,N_18294,N_18024);
nor U18918 (N_18918,N_18160,N_18259);
or U18919 (N_18919,N_18039,N_18311);
nand U18920 (N_18920,N_18420,N_18431);
nand U18921 (N_18921,N_18076,N_18153);
or U18922 (N_18922,N_18180,N_18003);
or U18923 (N_18923,N_18229,N_18482);
and U18924 (N_18924,N_18388,N_18019);
nand U18925 (N_18925,N_18020,N_18301);
nand U18926 (N_18926,N_18209,N_18432);
and U18927 (N_18927,N_18065,N_18225);
nor U18928 (N_18928,N_18225,N_18030);
nand U18929 (N_18929,N_18368,N_18460);
nand U18930 (N_18930,N_18488,N_18389);
nor U18931 (N_18931,N_18200,N_18144);
and U18932 (N_18932,N_18342,N_18115);
and U18933 (N_18933,N_18437,N_18100);
or U18934 (N_18934,N_18044,N_18041);
or U18935 (N_18935,N_18151,N_18408);
nand U18936 (N_18936,N_18428,N_18066);
and U18937 (N_18937,N_18120,N_18422);
and U18938 (N_18938,N_18190,N_18136);
nor U18939 (N_18939,N_18293,N_18178);
nor U18940 (N_18940,N_18341,N_18084);
or U18941 (N_18941,N_18034,N_18465);
and U18942 (N_18942,N_18114,N_18118);
nor U18943 (N_18943,N_18098,N_18493);
xnor U18944 (N_18944,N_18214,N_18284);
or U18945 (N_18945,N_18472,N_18211);
xor U18946 (N_18946,N_18253,N_18214);
or U18947 (N_18947,N_18249,N_18409);
xor U18948 (N_18948,N_18242,N_18264);
nand U18949 (N_18949,N_18216,N_18496);
nor U18950 (N_18950,N_18452,N_18086);
or U18951 (N_18951,N_18365,N_18296);
xor U18952 (N_18952,N_18014,N_18119);
xnor U18953 (N_18953,N_18224,N_18290);
and U18954 (N_18954,N_18128,N_18252);
xor U18955 (N_18955,N_18321,N_18037);
xor U18956 (N_18956,N_18231,N_18143);
nand U18957 (N_18957,N_18121,N_18349);
and U18958 (N_18958,N_18030,N_18061);
nor U18959 (N_18959,N_18224,N_18146);
nand U18960 (N_18960,N_18030,N_18180);
and U18961 (N_18961,N_18423,N_18138);
and U18962 (N_18962,N_18187,N_18362);
nand U18963 (N_18963,N_18367,N_18328);
and U18964 (N_18964,N_18210,N_18149);
and U18965 (N_18965,N_18041,N_18055);
and U18966 (N_18966,N_18327,N_18241);
nand U18967 (N_18967,N_18081,N_18351);
or U18968 (N_18968,N_18089,N_18328);
xor U18969 (N_18969,N_18371,N_18413);
xor U18970 (N_18970,N_18078,N_18334);
or U18971 (N_18971,N_18407,N_18096);
nor U18972 (N_18972,N_18146,N_18291);
or U18973 (N_18973,N_18011,N_18078);
or U18974 (N_18974,N_18373,N_18053);
nor U18975 (N_18975,N_18156,N_18169);
nand U18976 (N_18976,N_18323,N_18441);
nor U18977 (N_18977,N_18482,N_18256);
nand U18978 (N_18978,N_18004,N_18299);
nand U18979 (N_18979,N_18483,N_18079);
or U18980 (N_18980,N_18157,N_18478);
and U18981 (N_18981,N_18290,N_18286);
nor U18982 (N_18982,N_18130,N_18384);
nor U18983 (N_18983,N_18120,N_18386);
and U18984 (N_18984,N_18480,N_18003);
or U18985 (N_18985,N_18042,N_18284);
nor U18986 (N_18986,N_18234,N_18306);
xor U18987 (N_18987,N_18131,N_18480);
or U18988 (N_18988,N_18415,N_18243);
or U18989 (N_18989,N_18238,N_18023);
or U18990 (N_18990,N_18372,N_18493);
xnor U18991 (N_18991,N_18208,N_18073);
xnor U18992 (N_18992,N_18225,N_18052);
nand U18993 (N_18993,N_18491,N_18027);
nand U18994 (N_18994,N_18190,N_18161);
and U18995 (N_18995,N_18447,N_18428);
nand U18996 (N_18996,N_18472,N_18054);
nand U18997 (N_18997,N_18302,N_18306);
xnor U18998 (N_18998,N_18030,N_18137);
xnor U18999 (N_18999,N_18277,N_18263);
or U19000 (N_19000,N_18554,N_18619);
and U19001 (N_19001,N_18520,N_18553);
xnor U19002 (N_19002,N_18519,N_18922);
and U19003 (N_19003,N_18610,N_18606);
or U19004 (N_19004,N_18693,N_18970);
xnor U19005 (N_19005,N_18683,N_18721);
nor U19006 (N_19006,N_18604,N_18704);
xnor U19007 (N_19007,N_18694,N_18812);
nand U19008 (N_19008,N_18873,N_18742);
and U19009 (N_19009,N_18673,N_18962);
or U19010 (N_19010,N_18695,N_18846);
nor U19011 (N_19011,N_18587,N_18515);
or U19012 (N_19012,N_18931,N_18884);
or U19013 (N_19013,N_18888,N_18923);
and U19014 (N_19014,N_18821,N_18995);
xnor U19015 (N_19015,N_18591,N_18682);
or U19016 (N_19016,N_18664,N_18790);
xor U19017 (N_19017,N_18893,N_18951);
nand U19018 (N_19018,N_18781,N_18711);
or U19019 (N_19019,N_18674,N_18533);
nand U19020 (N_19020,N_18942,N_18521);
or U19021 (N_19021,N_18615,N_18621);
nand U19022 (N_19022,N_18601,N_18551);
nand U19023 (N_19023,N_18799,N_18612);
and U19024 (N_19024,N_18902,N_18872);
nand U19025 (N_19025,N_18598,N_18581);
and U19026 (N_19026,N_18798,N_18728);
xor U19027 (N_19027,N_18500,N_18522);
nor U19028 (N_19028,N_18810,N_18958);
and U19029 (N_19029,N_18941,N_18676);
or U19030 (N_19030,N_18734,N_18933);
nor U19031 (N_19031,N_18572,N_18513);
nand U19032 (N_19032,N_18719,N_18785);
nand U19033 (N_19033,N_18649,N_18749);
nor U19034 (N_19034,N_18824,N_18978);
nor U19035 (N_19035,N_18705,N_18968);
nor U19036 (N_19036,N_18724,N_18715);
and U19037 (N_19037,N_18972,N_18917);
and U19038 (N_19038,N_18731,N_18563);
nor U19039 (N_19039,N_18633,N_18766);
xnor U19040 (N_19040,N_18752,N_18898);
xnor U19041 (N_19041,N_18539,N_18776);
nor U19042 (N_19042,N_18988,N_18758);
and U19043 (N_19043,N_18547,N_18773);
nand U19044 (N_19044,N_18618,N_18686);
and U19045 (N_19045,N_18955,N_18645);
xnor U19046 (N_19046,N_18573,N_18709);
xor U19047 (N_19047,N_18768,N_18748);
xor U19048 (N_19048,N_18518,N_18911);
nand U19049 (N_19049,N_18862,N_18813);
or U19050 (N_19050,N_18915,N_18526);
nor U19051 (N_19051,N_18895,N_18739);
xor U19052 (N_19052,N_18880,N_18580);
nand U19053 (N_19053,N_18878,N_18608);
nor U19054 (N_19054,N_18793,N_18842);
nand U19055 (N_19055,N_18900,N_18712);
nand U19056 (N_19056,N_18635,N_18623);
and U19057 (N_19057,N_18548,N_18871);
and U19058 (N_19058,N_18849,N_18613);
xor U19059 (N_19059,N_18909,N_18720);
and U19060 (N_19060,N_18885,N_18698);
nand U19061 (N_19061,N_18901,N_18946);
or U19062 (N_19062,N_18956,N_18675);
xor U19063 (N_19063,N_18718,N_18648);
or U19064 (N_19064,N_18779,N_18960);
nor U19065 (N_19065,N_18899,N_18541);
nor U19066 (N_19066,N_18945,N_18511);
xnor U19067 (N_19067,N_18882,N_18961);
xor U19068 (N_19068,N_18971,N_18701);
or U19069 (N_19069,N_18883,N_18908);
xor U19070 (N_19070,N_18887,N_18928);
nor U19071 (N_19071,N_18865,N_18544);
nand U19072 (N_19072,N_18636,N_18640);
nand U19073 (N_19073,N_18687,N_18528);
xor U19074 (N_19074,N_18751,N_18671);
xor U19075 (N_19075,N_18843,N_18796);
or U19076 (N_19076,N_18780,N_18927);
xnor U19077 (N_19077,N_18545,N_18523);
nand U19078 (N_19078,N_18628,N_18754);
xnor U19079 (N_19079,N_18969,N_18991);
nor U19080 (N_19080,N_18627,N_18723);
or U19081 (N_19081,N_18590,N_18658);
or U19082 (N_19082,N_18653,N_18987);
nor U19083 (N_19083,N_18557,N_18529);
xor U19084 (N_19084,N_18827,N_18730);
and U19085 (N_19085,N_18797,N_18907);
xnor U19086 (N_19086,N_18630,N_18947);
xor U19087 (N_19087,N_18722,N_18517);
nand U19088 (N_19088,N_18708,N_18857);
and U19089 (N_19089,N_18665,N_18912);
nor U19090 (N_19090,N_18875,N_18753);
or U19091 (N_19091,N_18575,N_18828);
or U19092 (N_19092,N_18836,N_18910);
nor U19093 (N_19093,N_18853,N_18784);
and U19094 (N_19094,N_18540,N_18592);
nor U19095 (N_19095,N_18772,N_18605);
nor U19096 (N_19096,N_18620,N_18765);
xnor U19097 (N_19097,N_18918,N_18763);
xnor U19098 (N_19098,N_18603,N_18770);
nor U19099 (N_19099,N_18670,N_18807);
nor U19100 (N_19100,N_18546,N_18789);
or U19101 (N_19101,N_18920,N_18644);
nand U19102 (N_19102,N_18850,N_18841);
and U19103 (N_19103,N_18959,N_18943);
or U19104 (N_19104,N_18626,N_18903);
nor U19105 (N_19105,N_18840,N_18607);
nor U19106 (N_19106,N_18527,N_18556);
xnor U19107 (N_19107,N_18937,N_18896);
nor U19108 (N_19108,N_18762,N_18576);
xnor U19109 (N_19109,N_18891,N_18974);
nor U19110 (N_19110,N_18510,N_18847);
nor U19111 (N_19111,N_18663,N_18584);
or U19112 (N_19112,N_18565,N_18655);
or U19113 (N_19113,N_18854,N_18594);
xor U19114 (N_19114,N_18999,N_18501);
or U19115 (N_19115,N_18889,N_18688);
or U19116 (N_19116,N_18870,N_18549);
and U19117 (N_19117,N_18732,N_18589);
nand U19118 (N_19118,N_18555,N_18746);
or U19119 (N_19119,N_18791,N_18713);
xnor U19120 (N_19120,N_18532,N_18769);
and U19121 (N_19121,N_18552,N_18823);
xnor U19122 (N_19122,N_18833,N_18818);
and U19123 (N_19123,N_18595,N_18690);
or U19124 (N_19124,N_18803,N_18678);
xnor U19125 (N_19125,N_18881,N_18795);
nor U19126 (N_19126,N_18760,N_18926);
or U19127 (N_19127,N_18866,N_18743);
or U19128 (N_19128,N_18778,N_18886);
and U19129 (N_19129,N_18935,N_18844);
nand U19130 (N_19130,N_18921,N_18602);
or U19131 (N_19131,N_18816,N_18736);
nor U19132 (N_19132,N_18574,N_18617);
xnor U19133 (N_19133,N_18984,N_18745);
or U19134 (N_19134,N_18906,N_18508);
nor U19135 (N_19135,N_18822,N_18535);
nand U19136 (N_19136,N_18782,N_18830);
nand U19137 (N_19137,N_18643,N_18578);
xor U19138 (N_19138,N_18503,N_18934);
or U19139 (N_19139,N_18764,N_18660);
nand U19140 (N_19140,N_18560,N_18794);
nor U19141 (N_19141,N_18979,N_18938);
xor U19142 (N_19142,N_18876,N_18516);
nand U19143 (N_19143,N_18838,N_18514);
xnor U19144 (N_19144,N_18976,N_18867);
nor U19145 (N_19145,N_18577,N_18505);
nand U19146 (N_19146,N_18642,N_18856);
and U19147 (N_19147,N_18756,N_18767);
nor U19148 (N_19148,N_18811,N_18894);
xnor U19149 (N_19149,N_18638,N_18629);
nand U19150 (N_19150,N_18659,N_18855);
and U19151 (N_19151,N_18940,N_18637);
nand U19152 (N_19152,N_18994,N_18869);
nor U19153 (N_19153,N_18692,N_18725);
nand U19154 (N_19154,N_18646,N_18877);
nand U19155 (N_19155,N_18634,N_18948);
nor U19156 (N_19156,N_18661,N_18861);
xnor U19157 (N_19157,N_18829,N_18509);
and U19158 (N_19158,N_18800,N_18845);
or U19159 (N_19159,N_18531,N_18863);
nor U19160 (N_19160,N_18801,N_18837);
nand U19161 (N_19161,N_18919,N_18975);
xnor U19162 (N_19162,N_18757,N_18691);
and U19163 (N_19163,N_18733,N_18814);
nor U19164 (N_19164,N_18859,N_18585);
xnor U19165 (N_19165,N_18562,N_18700);
nor U19166 (N_19166,N_18741,N_18936);
nand U19167 (N_19167,N_18890,N_18534);
nor U19168 (N_19168,N_18611,N_18667);
xor U19169 (N_19169,N_18666,N_18672);
nor U19170 (N_19170,N_18689,N_18860);
or U19171 (N_19171,N_18726,N_18831);
xor U19172 (N_19172,N_18788,N_18826);
nor U19173 (N_19173,N_18740,N_18706);
nor U19174 (N_19174,N_18771,N_18967);
xor U19175 (N_19175,N_18982,N_18750);
nor U19176 (N_19176,N_18806,N_18852);
nor U19177 (N_19177,N_18668,N_18593);
or U19178 (N_19178,N_18543,N_18817);
and U19179 (N_19179,N_18932,N_18697);
nand U19180 (N_19180,N_18680,N_18579);
or U19181 (N_19181,N_18625,N_18566);
nand U19182 (N_19182,N_18569,N_18977);
nor U19183 (N_19183,N_18662,N_18805);
nor U19184 (N_19184,N_18558,N_18568);
xnor U19185 (N_19185,N_18652,N_18567);
xor U19186 (N_19186,N_18996,N_18993);
or U19187 (N_19187,N_18989,N_18596);
nand U19188 (N_19188,N_18647,N_18622);
or U19189 (N_19189,N_18950,N_18819);
and U19190 (N_19190,N_18702,N_18949);
nor U19191 (N_19191,N_18542,N_18651);
or U19192 (N_19192,N_18583,N_18524);
and U19193 (N_19193,N_18707,N_18815);
xor U19194 (N_19194,N_18848,N_18744);
or U19195 (N_19195,N_18537,N_18858);
xor U19196 (N_19196,N_18997,N_18561);
nand U19197 (N_19197,N_18507,N_18808);
nor U19198 (N_19198,N_18998,N_18614);
and U19199 (N_19199,N_18973,N_18913);
xnor U19200 (N_19200,N_18820,N_18624);
and U19201 (N_19201,N_18964,N_18684);
and U19202 (N_19202,N_18747,N_18729);
or U19203 (N_19203,N_18939,N_18914);
nor U19204 (N_19204,N_18761,N_18929);
and U19205 (N_19205,N_18677,N_18657);
nor U19206 (N_19206,N_18953,N_18980);
or U19207 (N_19207,N_18930,N_18530);
xor U19208 (N_19208,N_18559,N_18506);
xnor U19209 (N_19209,N_18786,N_18755);
nor U19210 (N_19210,N_18650,N_18792);
or U19211 (N_19211,N_18609,N_18512);
and U19212 (N_19212,N_18835,N_18502);
and U19213 (N_19213,N_18990,N_18639);
or U19214 (N_19214,N_18868,N_18656);
nand U19215 (N_19215,N_18832,N_18892);
and U19216 (N_19216,N_18600,N_18654);
nand U19217 (N_19217,N_18703,N_18825);
and U19218 (N_19218,N_18957,N_18679);
or U19219 (N_19219,N_18632,N_18571);
xnor U19220 (N_19220,N_18802,N_18669);
nor U19221 (N_19221,N_18564,N_18925);
or U19222 (N_19222,N_18641,N_18735);
nand U19223 (N_19223,N_18570,N_18685);
xor U19224 (N_19224,N_18716,N_18965);
nor U19225 (N_19225,N_18874,N_18681);
or U19226 (N_19226,N_18981,N_18737);
nand U19227 (N_19227,N_18710,N_18834);
xnor U19228 (N_19228,N_18774,N_18983);
or U19229 (N_19229,N_18616,N_18954);
and U19230 (N_19230,N_18538,N_18963);
nand U19231 (N_19231,N_18588,N_18525);
nand U19232 (N_19232,N_18783,N_18727);
nor U19233 (N_19233,N_18864,N_18879);
nand U19234 (N_19234,N_18804,N_18985);
nand U19235 (N_19235,N_18986,N_18944);
or U19236 (N_19236,N_18597,N_18504);
nor U19237 (N_19237,N_18738,N_18759);
nand U19238 (N_19238,N_18897,N_18631);
xnor U19239 (N_19239,N_18952,N_18582);
nor U19240 (N_19240,N_18717,N_18966);
nand U19241 (N_19241,N_18851,N_18550);
or U19242 (N_19242,N_18775,N_18699);
or U19243 (N_19243,N_18787,N_18992);
and U19244 (N_19244,N_18696,N_18777);
and U19245 (N_19245,N_18599,N_18809);
xor U19246 (N_19246,N_18536,N_18916);
nand U19247 (N_19247,N_18839,N_18924);
xor U19248 (N_19248,N_18586,N_18904);
xnor U19249 (N_19249,N_18905,N_18714);
and U19250 (N_19250,N_18979,N_18645);
xor U19251 (N_19251,N_18675,N_18941);
or U19252 (N_19252,N_18800,N_18647);
xor U19253 (N_19253,N_18987,N_18651);
or U19254 (N_19254,N_18578,N_18626);
and U19255 (N_19255,N_18797,N_18914);
nand U19256 (N_19256,N_18658,N_18879);
or U19257 (N_19257,N_18685,N_18548);
nor U19258 (N_19258,N_18929,N_18678);
xor U19259 (N_19259,N_18876,N_18896);
or U19260 (N_19260,N_18502,N_18942);
or U19261 (N_19261,N_18795,N_18784);
nor U19262 (N_19262,N_18942,N_18608);
nor U19263 (N_19263,N_18907,N_18623);
or U19264 (N_19264,N_18558,N_18573);
xnor U19265 (N_19265,N_18902,N_18898);
xor U19266 (N_19266,N_18672,N_18559);
nand U19267 (N_19267,N_18678,N_18516);
or U19268 (N_19268,N_18574,N_18833);
nor U19269 (N_19269,N_18711,N_18605);
xnor U19270 (N_19270,N_18884,N_18940);
xnor U19271 (N_19271,N_18744,N_18696);
nand U19272 (N_19272,N_18897,N_18633);
or U19273 (N_19273,N_18711,N_18568);
or U19274 (N_19274,N_18956,N_18586);
and U19275 (N_19275,N_18526,N_18696);
or U19276 (N_19276,N_18620,N_18811);
or U19277 (N_19277,N_18655,N_18649);
and U19278 (N_19278,N_18804,N_18710);
and U19279 (N_19279,N_18979,N_18644);
and U19280 (N_19280,N_18928,N_18721);
or U19281 (N_19281,N_18829,N_18653);
and U19282 (N_19282,N_18742,N_18712);
nand U19283 (N_19283,N_18588,N_18575);
and U19284 (N_19284,N_18751,N_18756);
nor U19285 (N_19285,N_18745,N_18764);
or U19286 (N_19286,N_18926,N_18909);
nor U19287 (N_19287,N_18734,N_18947);
and U19288 (N_19288,N_18610,N_18670);
or U19289 (N_19289,N_18680,N_18534);
or U19290 (N_19290,N_18814,N_18769);
or U19291 (N_19291,N_18816,N_18947);
xor U19292 (N_19292,N_18915,N_18926);
and U19293 (N_19293,N_18770,N_18747);
nor U19294 (N_19294,N_18752,N_18937);
xor U19295 (N_19295,N_18787,N_18883);
or U19296 (N_19296,N_18518,N_18749);
xor U19297 (N_19297,N_18597,N_18544);
nand U19298 (N_19298,N_18636,N_18858);
and U19299 (N_19299,N_18819,N_18612);
and U19300 (N_19300,N_18668,N_18823);
xnor U19301 (N_19301,N_18548,N_18525);
and U19302 (N_19302,N_18929,N_18968);
or U19303 (N_19303,N_18811,N_18898);
nand U19304 (N_19304,N_18795,N_18605);
nand U19305 (N_19305,N_18912,N_18817);
nand U19306 (N_19306,N_18885,N_18967);
nand U19307 (N_19307,N_18654,N_18653);
and U19308 (N_19308,N_18670,N_18721);
xor U19309 (N_19309,N_18945,N_18804);
xnor U19310 (N_19310,N_18893,N_18988);
xnor U19311 (N_19311,N_18583,N_18610);
and U19312 (N_19312,N_18929,N_18559);
nand U19313 (N_19313,N_18699,N_18521);
xnor U19314 (N_19314,N_18816,N_18708);
nand U19315 (N_19315,N_18554,N_18515);
xor U19316 (N_19316,N_18780,N_18640);
xor U19317 (N_19317,N_18550,N_18677);
nor U19318 (N_19318,N_18722,N_18755);
and U19319 (N_19319,N_18712,N_18639);
nand U19320 (N_19320,N_18623,N_18689);
nor U19321 (N_19321,N_18790,N_18517);
and U19322 (N_19322,N_18676,N_18593);
xnor U19323 (N_19323,N_18889,N_18516);
xnor U19324 (N_19324,N_18746,N_18757);
nor U19325 (N_19325,N_18833,N_18535);
or U19326 (N_19326,N_18951,N_18860);
and U19327 (N_19327,N_18676,N_18818);
or U19328 (N_19328,N_18523,N_18571);
or U19329 (N_19329,N_18585,N_18655);
or U19330 (N_19330,N_18996,N_18650);
nand U19331 (N_19331,N_18821,N_18655);
nand U19332 (N_19332,N_18615,N_18875);
xnor U19333 (N_19333,N_18985,N_18658);
xnor U19334 (N_19334,N_18782,N_18822);
nor U19335 (N_19335,N_18707,N_18906);
nor U19336 (N_19336,N_18751,N_18771);
or U19337 (N_19337,N_18610,N_18809);
nor U19338 (N_19338,N_18586,N_18632);
nor U19339 (N_19339,N_18571,N_18700);
and U19340 (N_19340,N_18877,N_18582);
xnor U19341 (N_19341,N_18804,N_18586);
xnor U19342 (N_19342,N_18833,N_18721);
and U19343 (N_19343,N_18917,N_18645);
nand U19344 (N_19344,N_18930,N_18986);
xor U19345 (N_19345,N_18964,N_18957);
xor U19346 (N_19346,N_18572,N_18975);
and U19347 (N_19347,N_18943,N_18510);
and U19348 (N_19348,N_18653,N_18774);
and U19349 (N_19349,N_18599,N_18911);
xnor U19350 (N_19350,N_18713,N_18608);
xnor U19351 (N_19351,N_18566,N_18540);
nand U19352 (N_19352,N_18668,N_18538);
and U19353 (N_19353,N_18538,N_18757);
or U19354 (N_19354,N_18561,N_18698);
xnor U19355 (N_19355,N_18706,N_18823);
nor U19356 (N_19356,N_18978,N_18989);
nand U19357 (N_19357,N_18878,N_18877);
or U19358 (N_19358,N_18966,N_18871);
and U19359 (N_19359,N_18903,N_18828);
nor U19360 (N_19360,N_18569,N_18820);
nand U19361 (N_19361,N_18757,N_18668);
nor U19362 (N_19362,N_18532,N_18642);
and U19363 (N_19363,N_18529,N_18921);
nand U19364 (N_19364,N_18539,N_18876);
or U19365 (N_19365,N_18509,N_18526);
xor U19366 (N_19366,N_18607,N_18715);
and U19367 (N_19367,N_18833,N_18737);
xnor U19368 (N_19368,N_18828,N_18833);
nor U19369 (N_19369,N_18512,N_18840);
nor U19370 (N_19370,N_18951,N_18969);
and U19371 (N_19371,N_18721,N_18682);
and U19372 (N_19372,N_18634,N_18998);
and U19373 (N_19373,N_18772,N_18996);
xor U19374 (N_19374,N_18971,N_18746);
and U19375 (N_19375,N_18846,N_18904);
or U19376 (N_19376,N_18650,N_18604);
xor U19377 (N_19377,N_18907,N_18555);
and U19378 (N_19378,N_18993,N_18711);
xnor U19379 (N_19379,N_18568,N_18830);
and U19380 (N_19380,N_18721,N_18736);
nand U19381 (N_19381,N_18636,N_18501);
xnor U19382 (N_19382,N_18845,N_18527);
nor U19383 (N_19383,N_18762,N_18777);
and U19384 (N_19384,N_18640,N_18955);
xnor U19385 (N_19385,N_18598,N_18794);
xor U19386 (N_19386,N_18666,N_18765);
or U19387 (N_19387,N_18732,N_18564);
and U19388 (N_19388,N_18863,N_18793);
xor U19389 (N_19389,N_18939,N_18736);
xor U19390 (N_19390,N_18592,N_18963);
xnor U19391 (N_19391,N_18951,N_18844);
or U19392 (N_19392,N_18652,N_18792);
xnor U19393 (N_19393,N_18525,N_18669);
and U19394 (N_19394,N_18988,N_18932);
or U19395 (N_19395,N_18962,N_18798);
or U19396 (N_19396,N_18615,N_18766);
nand U19397 (N_19397,N_18666,N_18893);
nand U19398 (N_19398,N_18831,N_18789);
nor U19399 (N_19399,N_18961,N_18980);
nor U19400 (N_19400,N_18804,N_18566);
or U19401 (N_19401,N_18836,N_18644);
or U19402 (N_19402,N_18663,N_18855);
xnor U19403 (N_19403,N_18896,N_18881);
and U19404 (N_19404,N_18672,N_18791);
nand U19405 (N_19405,N_18787,N_18838);
and U19406 (N_19406,N_18897,N_18595);
nand U19407 (N_19407,N_18541,N_18829);
nor U19408 (N_19408,N_18513,N_18908);
nand U19409 (N_19409,N_18800,N_18509);
nand U19410 (N_19410,N_18873,N_18831);
nand U19411 (N_19411,N_18653,N_18806);
or U19412 (N_19412,N_18762,N_18678);
or U19413 (N_19413,N_18914,N_18973);
nor U19414 (N_19414,N_18939,N_18980);
nand U19415 (N_19415,N_18551,N_18887);
xnor U19416 (N_19416,N_18879,N_18921);
nand U19417 (N_19417,N_18786,N_18856);
and U19418 (N_19418,N_18709,N_18806);
or U19419 (N_19419,N_18533,N_18943);
and U19420 (N_19420,N_18981,N_18886);
nor U19421 (N_19421,N_18920,N_18685);
nand U19422 (N_19422,N_18833,N_18963);
and U19423 (N_19423,N_18916,N_18816);
nand U19424 (N_19424,N_18879,N_18916);
and U19425 (N_19425,N_18637,N_18515);
nand U19426 (N_19426,N_18646,N_18905);
xor U19427 (N_19427,N_18569,N_18918);
and U19428 (N_19428,N_18839,N_18637);
nand U19429 (N_19429,N_18650,N_18683);
or U19430 (N_19430,N_18779,N_18711);
nand U19431 (N_19431,N_18831,N_18601);
or U19432 (N_19432,N_18891,N_18869);
or U19433 (N_19433,N_18647,N_18957);
and U19434 (N_19434,N_18687,N_18864);
xnor U19435 (N_19435,N_18941,N_18920);
nand U19436 (N_19436,N_18747,N_18637);
xnor U19437 (N_19437,N_18609,N_18630);
xor U19438 (N_19438,N_18874,N_18897);
and U19439 (N_19439,N_18573,N_18857);
or U19440 (N_19440,N_18510,N_18699);
and U19441 (N_19441,N_18849,N_18503);
xnor U19442 (N_19442,N_18829,N_18809);
nand U19443 (N_19443,N_18816,N_18866);
nand U19444 (N_19444,N_18520,N_18802);
or U19445 (N_19445,N_18913,N_18546);
xor U19446 (N_19446,N_18859,N_18624);
and U19447 (N_19447,N_18634,N_18941);
or U19448 (N_19448,N_18617,N_18925);
nand U19449 (N_19449,N_18876,N_18972);
and U19450 (N_19450,N_18769,N_18590);
nand U19451 (N_19451,N_18643,N_18662);
nand U19452 (N_19452,N_18871,N_18701);
nand U19453 (N_19453,N_18886,N_18973);
xnor U19454 (N_19454,N_18847,N_18818);
and U19455 (N_19455,N_18768,N_18898);
or U19456 (N_19456,N_18873,N_18833);
nand U19457 (N_19457,N_18851,N_18578);
and U19458 (N_19458,N_18967,N_18983);
nand U19459 (N_19459,N_18679,N_18751);
nor U19460 (N_19460,N_18877,N_18707);
or U19461 (N_19461,N_18533,N_18634);
and U19462 (N_19462,N_18896,N_18741);
and U19463 (N_19463,N_18650,N_18545);
and U19464 (N_19464,N_18630,N_18646);
and U19465 (N_19465,N_18556,N_18521);
nand U19466 (N_19466,N_18953,N_18955);
nand U19467 (N_19467,N_18685,N_18773);
nor U19468 (N_19468,N_18815,N_18545);
nor U19469 (N_19469,N_18642,N_18626);
or U19470 (N_19470,N_18841,N_18639);
and U19471 (N_19471,N_18666,N_18594);
nand U19472 (N_19472,N_18814,N_18552);
or U19473 (N_19473,N_18706,N_18952);
xnor U19474 (N_19474,N_18521,N_18793);
or U19475 (N_19475,N_18578,N_18716);
and U19476 (N_19476,N_18773,N_18791);
nor U19477 (N_19477,N_18808,N_18908);
or U19478 (N_19478,N_18812,N_18714);
nor U19479 (N_19479,N_18597,N_18687);
and U19480 (N_19480,N_18507,N_18697);
xor U19481 (N_19481,N_18560,N_18726);
nor U19482 (N_19482,N_18669,N_18554);
and U19483 (N_19483,N_18794,N_18509);
nor U19484 (N_19484,N_18641,N_18598);
xnor U19485 (N_19485,N_18568,N_18529);
nor U19486 (N_19486,N_18549,N_18864);
and U19487 (N_19487,N_18763,N_18938);
or U19488 (N_19488,N_18571,N_18610);
or U19489 (N_19489,N_18697,N_18768);
nor U19490 (N_19490,N_18774,N_18542);
or U19491 (N_19491,N_18584,N_18897);
or U19492 (N_19492,N_18633,N_18624);
or U19493 (N_19493,N_18910,N_18697);
nor U19494 (N_19494,N_18604,N_18803);
nand U19495 (N_19495,N_18846,N_18565);
nand U19496 (N_19496,N_18901,N_18891);
nand U19497 (N_19497,N_18632,N_18956);
nor U19498 (N_19498,N_18526,N_18940);
xor U19499 (N_19499,N_18736,N_18657);
xnor U19500 (N_19500,N_19448,N_19494);
xor U19501 (N_19501,N_19053,N_19377);
nand U19502 (N_19502,N_19059,N_19165);
and U19503 (N_19503,N_19435,N_19299);
or U19504 (N_19504,N_19351,N_19347);
nand U19505 (N_19505,N_19392,N_19277);
nor U19506 (N_19506,N_19447,N_19117);
and U19507 (N_19507,N_19352,N_19330);
and U19508 (N_19508,N_19420,N_19144);
nor U19509 (N_19509,N_19453,N_19489);
xnor U19510 (N_19510,N_19413,N_19194);
nand U19511 (N_19511,N_19335,N_19212);
xnor U19512 (N_19512,N_19017,N_19444);
nand U19513 (N_19513,N_19309,N_19493);
nand U19514 (N_19514,N_19043,N_19090);
and U19515 (N_19515,N_19204,N_19026);
xnor U19516 (N_19516,N_19302,N_19081);
xnor U19517 (N_19517,N_19441,N_19062);
xnor U19518 (N_19518,N_19084,N_19037);
xnor U19519 (N_19519,N_19189,N_19180);
or U19520 (N_19520,N_19206,N_19146);
nand U19521 (N_19521,N_19230,N_19115);
or U19522 (N_19522,N_19310,N_19496);
nor U19523 (N_19523,N_19312,N_19305);
nand U19524 (N_19524,N_19170,N_19221);
nor U19525 (N_19525,N_19487,N_19054);
xnor U19526 (N_19526,N_19270,N_19429);
or U19527 (N_19527,N_19412,N_19105);
xnor U19528 (N_19528,N_19224,N_19161);
nand U19529 (N_19529,N_19152,N_19306);
xnor U19530 (N_19530,N_19032,N_19354);
and U19531 (N_19531,N_19148,N_19235);
nand U19532 (N_19532,N_19356,N_19359);
or U19533 (N_19533,N_19072,N_19050);
xnor U19534 (N_19534,N_19411,N_19488);
or U19535 (N_19535,N_19492,N_19385);
nor U19536 (N_19536,N_19193,N_19378);
nand U19537 (N_19537,N_19342,N_19329);
nand U19538 (N_19538,N_19045,N_19322);
nor U19539 (N_19539,N_19480,N_19005);
or U19540 (N_19540,N_19432,N_19314);
and U19541 (N_19541,N_19477,N_19091);
and U19542 (N_19542,N_19215,N_19058);
xnor U19543 (N_19543,N_19325,N_19135);
nand U19544 (N_19544,N_19225,N_19403);
nand U19545 (N_19545,N_19227,N_19339);
nand U19546 (N_19546,N_19001,N_19183);
nand U19547 (N_19547,N_19257,N_19009);
or U19548 (N_19548,N_19231,N_19121);
and U19549 (N_19549,N_19217,N_19308);
or U19550 (N_19550,N_19415,N_19141);
or U19551 (N_19551,N_19267,N_19401);
nor U19552 (N_19552,N_19426,N_19100);
and U19553 (N_19553,N_19164,N_19099);
nor U19554 (N_19554,N_19069,N_19210);
and U19555 (N_19555,N_19177,N_19458);
or U19556 (N_19556,N_19422,N_19056);
and U19557 (N_19557,N_19098,N_19174);
nor U19558 (N_19558,N_19338,N_19440);
or U19559 (N_19559,N_19218,N_19082);
and U19560 (N_19560,N_19355,N_19119);
xnor U19561 (N_19561,N_19387,N_19280);
and U19562 (N_19562,N_19243,N_19134);
and U19563 (N_19563,N_19162,N_19213);
xnor U19564 (N_19564,N_19349,N_19334);
and U19565 (N_19565,N_19048,N_19239);
or U19566 (N_19566,N_19394,N_19248);
or U19567 (N_19567,N_19229,N_19366);
nor U19568 (N_19568,N_19010,N_19168);
nor U19569 (N_19569,N_19083,N_19427);
and U19570 (N_19570,N_19110,N_19467);
or U19571 (N_19571,N_19129,N_19238);
or U19572 (N_19572,N_19195,N_19348);
nand U19573 (N_19573,N_19395,N_19102);
nand U19574 (N_19574,N_19317,N_19188);
nand U19575 (N_19575,N_19416,N_19262);
or U19576 (N_19576,N_19373,N_19002);
or U19577 (N_19577,N_19360,N_19311);
and U19578 (N_19578,N_19485,N_19143);
nand U19579 (N_19579,N_19240,N_19191);
xnor U19580 (N_19580,N_19469,N_19389);
xor U19581 (N_19581,N_19296,N_19085);
and U19582 (N_19582,N_19247,N_19086);
nor U19583 (N_19583,N_19220,N_19184);
and U19584 (N_19584,N_19236,N_19076);
nand U19585 (N_19585,N_19068,N_19479);
xnor U19586 (N_19586,N_19278,N_19003);
or U19587 (N_19587,N_19301,N_19285);
xnor U19588 (N_19588,N_19233,N_19434);
nand U19589 (N_19589,N_19315,N_19481);
and U19590 (N_19590,N_19078,N_19374);
xnor U19591 (N_19591,N_19461,N_19391);
xnor U19592 (N_19592,N_19020,N_19147);
nor U19593 (N_19593,N_19096,N_19067);
nand U19594 (N_19594,N_19261,N_19409);
nand U19595 (N_19595,N_19439,N_19042);
nand U19596 (N_19596,N_19297,N_19160);
nor U19597 (N_19597,N_19397,N_19064);
nor U19598 (N_19598,N_19242,N_19040);
or U19599 (N_19599,N_19071,N_19456);
and U19600 (N_19600,N_19203,N_19030);
or U19601 (N_19601,N_19476,N_19169);
and U19602 (N_19602,N_19109,N_19362);
nand U19603 (N_19603,N_19158,N_19404);
and U19604 (N_19604,N_19462,N_19122);
xnor U19605 (N_19605,N_19013,N_19087);
xnor U19606 (N_19606,N_19179,N_19150);
nor U19607 (N_19607,N_19414,N_19320);
or U19608 (N_19608,N_19331,N_19450);
and U19609 (N_19609,N_19120,N_19021);
nor U19610 (N_19610,N_19181,N_19323);
nor U19611 (N_19611,N_19118,N_19318);
and U19612 (N_19612,N_19430,N_19077);
and U19613 (N_19613,N_19445,N_19237);
and U19614 (N_19614,N_19190,N_19291);
nor U19615 (N_19615,N_19365,N_19128);
and U19616 (N_19616,N_19446,N_19149);
and U19617 (N_19617,N_19198,N_19419);
nor U19618 (N_19618,N_19127,N_19142);
xor U19619 (N_19619,N_19163,N_19222);
and U19620 (N_19620,N_19061,N_19327);
nor U19621 (N_19621,N_19324,N_19103);
xnor U19622 (N_19622,N_19490,N_19313);
nand U19623 (N_19623,N_19465,N_19421);
or U19624 (N_19624,N_19132,N_19358);
nand U19625 (N_19625,N_19264,N_19018);
xor U19626 (N_19626,N_19471,N_19497);
or U19627 (N_19627,N_19178,N_19151);
nor U19628 (N_19628,N_19350,N_19136);
and U19629 (N_19629,N_19024,N_19393);
nor U19630 (N_19630,N_19216,N_19341);
and U19631 (N_19631,N_19156,N_19486);
and U19632 (N_19632,N_19436,N_19316);
nand U19633 (N_19633,N_19271,N_19166);
xor U19634 (N_19634,N_19012,N_19396);
nor U19635 (N_19635,N_19140,N_19019);
and U19636 (N_19636,N_19408,N_19386);
xnor U19637 (N_19637,N_19281,N_19075);
xnor U19638 (N_19638,N_19113,N_19094);
nand U19639 (N_19639,N_19294,N_19182);
and U19640 (N_19640,N_19246,N_19367);
nand U19641 (N_19641,N_19375,N_19263);
or U19642 (N_19642,N_19259,N_19035);
and U19643 (N_19643,N_19390,N_19155);
nor U19644 (N_19644,N_19167,N_19258);
and U19645 (N_19645,N_19451,N_19423);
nor U19646 (N_19646,N_19343,N_19364);
nor U19647 (N_19647,N_19405,N_19251);
nand U19648 (N_19648,N_19474,N_19011);
and U19649 (N_19649,N_19014,N_19376);
and U19650 (N_19650,N_19292,N_19186);
nor U19651 (N_19651,N_19283,N_19382);
nand U19652 (N_19652,N_19379,N_19433);
or U19653 (N_19653,N_19000,N_19463);
and U19654 (N_19654,N_19326,N_19255);
nor U19655 (N_19655,N_19372,N_19250);
and U19656 (N_19656,N_19332,N_19455);
xnor U19657 (N_19657,N_19027,N_19368);
xor U19658 (N_19658,N_19266,N_19065);
and U19659 (N_19659,N_19004,N_19208);
and U19660 (N_19660,N_19388,N_19057);
or U19661 (N_19661,N_19498,N_19345);
xnor U19662 (N_19662,N_19399,N_19383);
xor U19663 (N_19663,N_19400,N_19052);
nand U19664 (N_19664,N_19093,N_19046);
or U19665 (N_19665,N_19293,N_19205);
xnor U19666 (N_19666,N_19049,N_19380);
and U19667 (N_19667,N_19060,N_19284);
nor U19668 (N_19668,N_19197,N_19101);
xor U19669 (N_19669,N_19256,N_19133);
or U19670 (N_19670,N_19464,N_19097);
or U19671 (N_19671,N_19276,N_19337);
xnor U19672 (N_19672,N_19066,N_19131);
nand U19673 (N_19673,N_19073,N_19457);
xnor U19674 (N_19674,N_19112,N_19279);
xnor U19675 (N_19675,N_19442,N_19344);
and U19676 (N_19676,N_19333,N_19398);
or U19677 (N_19677,N_19137,N_19176);
or U19678 (N_19678,N_19211,N_19468);
xnor U19679 (N_19679,N_19044,N_19138);
and U19680 (N_19680,N_19234,N_19371);
nand U19681 (N_19681,N_19123,N_19089);
nor U19682 (N_19682,N_19088,N_19039);
nor U19683 (N_19683,N_19023,N_19209);
nand U19684 (N_19684,N_19428,N_19286);
or U19685 (N_19685,N_19106,N_19438);
or U19686 (N_19686,N_19070,N_19241);
nand U19687 (N_19687,N_19370,N_19381);
xor U19688 (N_19688,N_19417,N_19307);
nor U19689 (N_19689,N_19475,N_19047);
nor U19690 (N_19690,N_19126,N_19092);
nor U19691 (N_19691,N_19406,N_19200);
xnor U19692 (N_19692,N_19300,N_19201);
xnor U19693 (N_19693,N_19029,N_19249);
nand U19694 (N_19694,N_19287,N_19478);
nor U19695 (N_19695,N_19491,N_19028);
nor U19696 (N_19696,N_19454,N_19016);
xnor U19697 (N_19697,N_19268,N_19402);
or U19698 (N_19698,N_19482,N_19063);
and U19699 (N_19699,N_19290,N_19095);
nor U19700 (N_19700,N_19288,N_19384);
and U19701 (N_19701,N_19431,N_19346);
or U19702 (N_19702,N_19175,N_19269);
or U19703 (N_19703,N_19449,N_19055);
or U19704 (N_19704,N_19172,N_19452);
or U19705 (N_19705,N_19304,N_19336);
nand U19706 (N_19706,N_19015,N_19226);
nand U19707 (N_19707,N_19499,N_19260);
nor U19708 (N_19708,N_19319,N_19145);
nor U19709 (N_19709,N_19252,N_19466);
xor U19710 (N_19710,N_19357,N_19187);
nand U19711 (N_19711,N_19116,N_19079);
and U19712 (N_19712,N_19298,N_19495);
or U19713 (N_19713,N_19130,N_19007);
and U19714 (N_19714,N_19080,N_19008);
nand U19715 (N_19715,N_19254,N_19223);
and U19716 (N_19716,N_19425,N_19111);
or U19717 (N_19717,N_19199,N_19038);
and U19718 (N_19718,N_19173,N_19036);
and U19719 (N_19719,N_19353,N_19185);
nand U19720 (N_19720,N_19041,N_19321);
and U19721 (N_19721,N_19274,N_19484);
nor U19722 (N_19722,N_19244,N_19153);
or U19723 (N_19723,N_19104,N_19369);
and U19724 (N_19724,N_19202,N_19033);
nand U19725 (N_19725,N_19214,N_19196);
xnor U19726 (N_19726,N_19157,N_19219);
and U19727 (N_19727,N_19124,N_19361);
nand U19728 (N_19728,N_19328,N_19407);
and U19729 (N_19729,N_19265,N_19025);
nor U19730 (N_19730,N_19034,N_19114);
xnor U19731 (N_19731,N_19272,N_19470);
and U19732 (N_19732,N_19022,N_19459);
xor U19733 (N_19733,N_19031,N_19154);
nand U19734 (N_19734,N_19282,N_19275);
xnor U19735 (N_19735,N_19289,N_19472);
nand U19736 (N_19736,N_19473,N_19171);
nand U19737 (N_19737,N_19303,N_19228);
nor U19738 (N_19738,N_19273,N_19051);
nor U19739 (N_19739,N_19125,N_19107);
nor U19740 (N_19740,N_19108,N_19232);
xor U19741 (N_19741,N_19245,N_19437);
nor U19742 (N_19742,N_19295,N_19443);
nor U19743 (N_19743,N_19363,N_19207);
nand U19744 (N_19744,N_19139,N_19192);
and U19745 (N_19745,N_19418,N_19424);
xnor U19746 (N_19746,N_19253,N_19460);
and U19747 (N_19747,N_19006,N_19483);
nor U19748 (N_19748,N_19159,N_19340);
xor U19749 (N_19749,N_19410,N_19074);
or U19750 (N_19750,N_19148,N_19122);
nor U19751 (N_19751,N_19308,N_19027);
nand U19752 (N_19752,N_19195,N_19130);
or U19753 (N_19753,N_19246,N_19450);
nor U19754 (N_19754,N_19281,N_19227);
nor U19755 (N_19755,N_19127,N_19223);
and U19756 (N_19756,N_19136,N_19316);
or U19757 (N_19757,N_19013,N_19285);
xnor U19758 (N_19758,N_19269,N_19457);
or U19759 (N_19759,N_19428,N_19053);
nor U19760 (N_19760,N_19304,N_19273);
or U19761 (N_19761,N_19457,N_19094);
nor U19762 (N_19762,N_19306,N_19223);
and U19763 (N_19763,N_19137,N_19128);
or U19764 (N_19764,N_19201,N_19496);
xor U19765 (N_19765,N_19482,N_19105);
and U19766 (N_19766,N_19344,N_19278);
nand U19767 (N_19767,N_19265,N_19335);
or U19768 (N_19768,N_19147,N_19319);
nor U19769 (N_19769,N_19460,N_19413);
nand U19770 (N_19770,N_19290,N_19315);
nor U19771 (N_19771,N_19354,N_19367);
or U19772 (N_19772,N_19086,N_19416);
nand U19773 (N_19773,N_19199,N_19343);
and U19774 (N_19774,N_19091,N_19385);
and U19775 (N_19775,N_19309,N_19050);
or U19776 (N_19776,N_19109,N_19108);
nor U19777 (N_19777,N_19376,N_19433);
nor U19778 (N_19778,N_19463,N_19069);
and U19779 (N_19779,N_19165,N_19110);
xor U19780 (N_19780,N_19236,N_19431);
nor U19781 (N_19781,N_19431,N_19305);
and U19782 (N_19782,N_19412,N_19132);
nor U19783 (N_19783,N_19401,N_19312);
xnor U19784 (N_19784,N_19029,N_19253);
nor U19785 (N_19785,N_19141,N_19041);
nand U19786 (N_19786,N_19108,N_19085);
or U19787 (N_19787,N_19080,N_19457);
nor U19788 (N_19788,N_19457,N_19389);
nor U19789 (N_19789,N_19218,N_19310);
xnor U19790 (N_19790,N_19259,N_19449);
nor U19791 (N_19791,N_19131,N_19057);
and U19792 (N_19792,N_19133,N_19458);
or U19793 (N_19793,N_19280,N_19291);
nand U19794 (N_19794,N_19246,N_19464);
nand U19795 (N_19795,N_19260,N_19012);
or U19796 (N_19796,N_19235,N_19354);
and U19797 (N_19797,N_19331,N_19355);
nand U19798 (N_19798,N_19137,N_19115);
and U19799 (N_19799,N_19143,N_19011);
xnor U19800 (N_19800,N_19014,N_19197);
nor U19801 (N_19801,N_19467,N_19390);
nand U19802 (N_19802,N_19274,N_19285);
nand U19803 (N_19803,N_19150,N_19331);
and U19804 (N_19804,N_19460,N_19157);
nor U19805 (N_19805,N_19204,N_19356);
xor U19806 (N_19806,N_19446,N_19329);
nand U19807 (N_19807,N_19063,N_19109);
nor U19808 (N_19808,N_19442,N_19169);
nand U19809 (N_19809,N_19440,N_19421);
xnor U19810 (N_19810,N_19284,N_19433);
nand U19811 (N_19811,N_19195,N_19328);
nand U19812 (N_19812,N_19237,N_19386);
nor U19813 (N_19813,N_19444,N_19275);
xnor U19814 (N_19814,N_19458,N_19152);
or U19815 (N_19815,N_19163,N_19391);
xor U19816 (N_19816,N_19029,N_19445);
xor U19817 (N_19817,N_19163,N_19030);
xor U19818 (N_19818,N_19221,N_19362);
or U19819 (N_19819,N_19354,N_19254);
nor U19820 (N_19820,N_19422,N_19397);
xnor U19821 (N_19821,N_19228,N_19341);
and U19822 (N_19822,N_19457,N_19453);
xor U19823 (N_19823,N_19098,N_19290);
xnor U19824 (N_19824,N_19297,N_19149);
nor U19825 (N_19825,N_19302,N_19409);
xor U19826 (N_19826,N_19067,N_19456);
nor U19827 (N_19827,N_19217,N_19280);
xor U19828 (N_19828,N_19237,N_19185);
and U19829 (N_19829,N_19488,N_19174);
nor U19830 (N_19830,N_19356,N_19415);
or U19831 (N_19831,N_19368,N_19248);
and U19832 (N_19832,N_19086,N_19459);
nor U19833 (N_19833,N_19240,N_19396);
and U19834 (N_19834,N_19313,N_19282);
nor U19835 (N_19835,N_19426,N_19198);
or U19836 (N_19836,N_19298,N_19405);
xor U19837 (N_19837,N_19411,N_19126);
or U19838 (N_19838,N_19371,N_19378);
nor U19839 (N_19839,N_19086,N_19136);
or U19840 (N_19840,N_19268,N_19308);
xnor U19841 (N_19841,N_19370,N_19235);
nand U19842 (N_19842,N_19441,N_19335);
nor U19843 (N_19843,N_19063,N_19058);
nor U19844 (N_19844,N_19045,N_19415);
or U19845 (N_19845,N_19190,N_19201);
nand U19846 (N_19846,N_19456,N_19015);
and U19847 (N_19847,N_19469,N_19299);
or U19848 (N_19848,N_19441,N_19488);
or U19849 (N_19849,N_19237,N_19086);
and U19850 (N_19850,N_19164,N_19306);
or U19851 (N_19851,N_19191,N_19305);
and U19852 (N_19852,N_19171,N_19297);
or U19853 (N_19853,N_19461,N_19265);
nor U19854 (N_19854,N_19294,N_19066);
nor U19855 (N_19855,N_19094,N_19239);
nor U19856 (N_19856,N_19477,N_19370);
nand U19857 (N_19857,N_19384,N_19485);
nor U19858 (N_19858,N_19085,N_19386);
xor U19859 (N_19859,N_19389,N_19032);
or U19860 (N_19860,N_19090,N_19386);
and U19861 (N_19861,N_19242,N_19284);
nor U19862 (N_19862,N_19028,N_19323);
nor U19863 (N_19863,N_19138,N_19233);
and U19864 (N_19864,N_19356,N_19219);
xor U19865 (N_19865,N_19369,N_19045);
xor U19866 (N_19866,N_19205,N_19357);
nand U19867 (N_19867,N_19430,N_19196);
nand U19868 (N_19868,N_19350,N_19192);
or U19869 (N_19869,N_19234,N_19184);
nand U19870 (N_19870,N_19165,N_19034);
and U19871 (N_19871,N_19221,N_19478);
nand U19872 (N_19872,N_19084,N_19066);
and U19873 (N_19873,N_19065,N_19137);
nor U19874 (N_19874,N_19387,N_19341);
xor U19875 (N_19875,N_19467,N_19202);
nor U19876 (N_19876,N_19457,N_19446);
nor U19877 (N_19877,N_19464,N_19044);
and U19878 (N_19878,N_19318,N_19328);
xnor U19879 (N_19879,N_19286,N_19245);
and U19880 (N_19880,N_19117,N_19246);
xor U19881 (N_19881,N_19253,N_19423);
nor U19882 (N_19882,N_19167,N_19464);
nand U19883 (N_19883,N_19467,N_19286);
nor U19884 (N_19884,N_19404,N_19377);
nand U19885 (N_19885,N_19324,N_19261);
nand U19886 (N_19886,N_19105,N_19350);
nand U19887 (N_19887,N_19365,N_19226);
xnor U19888 (N_19888,N_19478,N_19455);
and U19889 (N_19889,N_19269,N_19101);
or U19890 (N_19890,N_19498,N_19075);
nand U19891 (N_19891,N_19260,N_19444);
nor U19892 (N_19892,N_19002,N_19398);
and U19893 (N_19893,N_19101,N_19291);
nand U19894 (N_19894,N_19173,N_19231);
or U19895 (N_19895,N_19054,N_19402);
xor U19896 (N_19896,N_19122,N_19189);
or U19897 (N_19897,N_19420,N_19130);
nand U19898 (N_19898,N_19451,N_19158);
and U19899 (N_19899,N_19386,N_19069);
xor U19900 (N_19900,N_19298,N_19261);
nor U19901 (N_19901,N_19487,N_19448);
and U19902 (N_19902,N_19499,N_19391);
and U19903 (N_19903,N_19335,N_19457);
nand U19904 (N_19904,N_19060,N_19073);
nand U19905 (N_19905,N_19297,N_19394);
nor U19906 (N_19906,N_19046,N_19097);
nor U19907 (N_19907,N_19055,N_19429);
and U19908 (N_19908,N_19260,N_19203);
nand U19909 (N_19909,N_19031,N_19245);
xor U19910 (N_19910,N_19015,N_19075);
xnor U19911 (N_19911,N_19074,N_19131);
and U19912 (N_19912,N_19093,N_19281);
or U19913 (N_19913,N_19310,N_19415);
or U19914 (N_19914,N_19035,N_19105);
nor U19915 (N_19915,N_19202,N_19062);
nand U19916 (N_19916,N_19007,N_19107);
xor U19917 (N_19917,N_19392,N_19402);
or U19918 (N_19918,N_19079,N_19430);
and U19919 (N_19919,N_19250,N_19132);
nor U19920 (N_19920,N_19435,N_19478);
xnor U19921 (N_19921,N_19260,N_19386);
nor U19922 (N_19922,N_19445,N_19169);
xor U19923 (N_19923,N_19442,N_19341);
and U19924 (N_19924,N_19193,N_19317);
nand U19925 (N_19925,N_19106,N_19112);
xnor U19926 (N_19926,N_19491,N_19326);
xor U19927 (N_19927,N_19081,N_19343);
nand U19928 (N_19928,N_19328,N_19193);
or U19929 (N_19929,N_19044,N_19306);
or U19930 (N_19930,N_19168,N_19272);
or U19931 (N_19931,N_19107,N_19058);
nand U19932 (N_19932,N_19024,N_19319);
xnor U19933 (N_19933,N_19494,N_19390);
xor U19934 (N_19934,N_19447,N_19372);
nor U19935 (N_19935,N_19421,N_19186);
nand U19936 (N_19936,N_19121,N_19165);
and U19937 (N_19937,N_19383,N_19371);
or U19938 (N_19938,N_19216,N_19058);
nor U19939 (N_19939,N_19170,N_19059);
and U19940 (N_19940,N_19200,N_19466);
and U19941 (N_19941,N_19109,N_19048);
and U19942 (N_19942,N_19385,N_19333);
nor U19943 (N_19943,N_19478,N_19425);
or U19944 (N_19944,N_19479,N_19033);
nor U19945 (N_19945,N_19323,N_19384);
xnor U19946 (N_19946,N_19241,N_19276);
or U19947 (N_19947,N_19428,N_19254);
and U19948 (N_19948,N_19143,N_19470);
and U19949 (N_19949,N_19288,N_19260);
or U19950 (N_19950,N_19003,N_19102);
or U19951 (N_19951,N_19004,N_19276);
nand U19952 (N_19952,N_19372,N_19379);
and U19953 (N_19953,N_19428,N_19483);
or U19954 (N_19954,N_19324,N_19375);
or U19955 (N_19955,N_19280,N_19443);
or U19956 (N_19956,N_19499,N_19389);
or U19957 (N_19957,N_19014,N_19017);
nor U19958 (N_19958,N_19145,N_19483);
nand U19959 (N_19959,N_19369,N_19250);
or U19960 (N_19960,N_19436,N_19156);
or U19961 (N_19961,N_19205,N_19026);
and U19962 (N_19962,N_19218,N_19048);
nor U19963 (N_19963,N_19018,N_19209);
and U19964 (N_19964,N_19298,N_19422);
xnor U19965 (N_19965,N_19165,N_19290);
nor U19966 (N_19966,N_19144,N_19000);
xor U19967 (N_19967,N_19255,N_19253);
xor U19968 (N_19968,N_19038,N_19419);
nand U19969 (N_19969,N_19420,N_19380);
and U19970 (N_19970,N_19207,N_19237);
xor U19971 (N_19971,N_19396,N_19311);
nor U19972 (N_19972,N_19357,N_19068);
nand U19973 (N_19973,N_19056,N_19005);
nand U19974 (N_19974,N_19264,N_19498);
or U19975 (N_19975,N_19238,N_19165);
and U19976 (N_19976,N_19238,N_19270);
nand U19977 (N_19977,N_19163,N_19491);
nand U19978 (N_19978,N_19206,N_19411);
and U19979 (N_19979,N_19286,N_19223);
or U19980 (N_19980,N_19320,N_19490);
xnor U19981 (N_19981,N_19377,N_19093);
or U19982 (N_19982,N_19209,N_19288);
nand U19983 (N_19983,N_19121,N_19096);
or U19984 (N_19984,N_19282,N_19385);
xnor U19985 (N_19985,N_19161,N_19278);
and U19986 (N_19986,N_19495,N_19191);
nand U19987 (N_19987,N_19135,N_19193);
or U19988 (N_19988,N_19094,N_19245);
xor U19989 (N_19989,N_19458,N_19487);
xnor U19990 (N_19990,N_19439,N_19328);
xnor U19991 (N_19991,N_19232,N_19366);
nand U19992 (N_19992,N_19202,N_19268);
or U19993 (N_19993,N_19144,N_19286);
nor U19994 (N_19994,N_19444,N_19132);
xor U19995 (N_19995,N_19324,N_19140);
nor U19996 (N_19996,N_19157,N_19177);
and U19997 (N_19997,N_19210,N_19240);
nor U19998 (N_19998,N_19312,N_19420);
and U19999 (N_19999,N_19166,N_19373);
nand UO_0 (O_0,N_19686,N_19791);
or UO_1 (O_1,N_19871,N_19688);
nor UO_2 (O_2,N_19980,N_19519);
and UO_3 (O_3,N_19587,N_19925);
xnor UO_4 (O_4,N_19917,N_19597);
nor UO_5 (O_5,N_19785,N_19648);
xnor UO_6 (O_6,N_19713,N_19674);
nor UO_7 (O_7,N_19941,N_19699);
or UO_8 (O_8,N_19908,N_19976);
and UO_9 (O_9,N_19517,N_19650);
nand UO_10 (O_10,N_19526,N_19998);
and UO_11 (O_11,N_19865,N_19729);
xnor UO_12 (O_12,N_19877,N_19876);
xor UO_13 (O_13,N_19863,N_19851);
nor UO_14 (O_14,N_19602,N_19987);
or UO_15 (O_15,N_19751,N_19770);
or UO_16 (O_16,N_19986,N_19533);
and UO_17 (O_17,N_19920,N_19773);
or UO_18 (O_18,N_19826,N_19681);
nand UO_19 (O_19,N_19833,N_19937);
nand UO_20 (O_20,N_19895,N_19717);
xor UO_21 (O_21,N_19961,N_19931);
nand UO_22 (O_22,N_19616,N_19809);
and UO_23 (O_23,N_19520,N_19854);
nand UO_24 (O_24,N_19513,N_19595);
xor UO_25 (O_25,N_19757,N_19693);
nand UO_26 (O_26,N_19657,N_19868);
and UO_27 (O_27,N_19952,N_19535);
xnor UO_28 (O_28,N_19913,N_19608);
xnor UO_29 (O_29,N_19636,N_19735);
nor UO_30 (O_30,N_19839,N_19905);
xnor UO_31 (O_31,N_19601,N_19823);
nand UO_32 (O_32,N_19655,N_19704);
and UO_33 (O_33,N_19822,N_19645);
nor UO_34 (O_34,N_19829,N_19666);
nand UO_35 (O_35,N_19607,N_19664);
nand UO_36 (O_36,N_19754,N_19623);
and UO_37 (O_37,N_19971,N_19642);
nand UO_38 (O_38,N_19893,N_19700);
xnor UO_39 (O_39,N_19599,N_19677);
nor UO_40 (O_40,N_19705,N_19724);
xnor UO_41 (O_41,N_19989,N_19953);
nand UO_42 (O_42,N_19879,N_19631);
nor UO_43 (O_43,N_19887,N_19988);
nand UO_44 (O_44,N_19618,N_19944);
and UO_45 (O_45,N_19656,N_19716);
and UO_46 (O_46,N_19514,N_19529);
xor UO_47 (O_47,N_19641,N_19512);
nor UO_48 (O_48,N_19779,N_19938);
and UO_49 (O_49,N_19983,N_19834);
and UO_50 (O_50,N_19995,N_19906);
and UO_51 (O_51,N_19878,N_19554);
nor UO_52 (O_52,N_19584,N_19840);
or UO_53 (O_53,N_19510,N_19565);
nor UO_54 (O_54,N_19993,N_19598);
xor UO_55 (O_55,N_19538,N_19718);
or UO_56 (O_56,N_19847,N_19721);
nor UO_57 (O_57,N_19778,N_19614);
nand UO_58 (O_58,N_19794,N_19996);
nor UO_59 (O_59,N_19892,N_19685);
or UO_60 (O_60,N_19540,N_19860);
or UO_61 (O_61,N_19578,N_19982);
nor UO_62 (O_62,N_19518,N_19985);
xor UO_63 (O_63,N_19504,N_19991);
and UO_64 (O_64,N_19821,N_19886);
nor UO_65 (O_65,N_19555,N_19621);
nand UO_66 (O_66,N_19796,N_19615);
or UO_67 (O_67,N_19814,N_19680);
and UO_68 (O_68,N_19815,N_19710);
nand UO_69 (O_69,N_19869,N_19737);
nand UO_70 (O_70,N_19562,N_19795);
nor UO_71 (O_71,N_19684,N_19901);
nand UO_72 (O_72,N_19671,N_19675);
nand UO_73 (O_73,N_19975,N_19738);
nor UO_74 (O_74,N_19932,N_19862);
nand UO_75 (O_75,N_19997,N_19760);
nand UO_76 (O_76,N_19611,N_19654);
or UO_77 (O_77,N_19808,N_19954);
nand UO_78 (O_78,N_19825,N_19872);
nor UO_79 (O_79,N_19947,N_19544);
xnor UO_80 (O_80,N_19845,N_19748);
nor UO_81 (O_81,N_19707,N_19850);
or UO_82 (O_82,N_19593,N_19790);
xnor UO_83 (O_83,N_19969,N_19743);
or UO_84 (O_84,N_19950,N_19559);
or UO_85 (O_85,N_19768,N_19665);
nor UO_86 (O_86,N_19668,N_19816);
xnor UO_87 (O_87,N_19832,N_19509);
or UO_88 (O_88,N_19900,N_19697);
nor UO_89 (O_89,N_19817,N_19919);
nand UO_90 (O_90,N_19723,N_19525);
nand UO_91 (O_91,N_19708,N_19864);
or UO_92 (O_92,N_19807,N_19927);
and UO_93 (O_93,N_19506,N_19591);
nand UO_94 (O_94,N_19805,N_19867);
nor UO_95 (O_95,N_19799,N_19861);
xnor UO_96 (O_96,N_19866,N_19683);
or UO_97 (O_97,N_19739,N_19889);
or UO_98 (O_98,N_19965,N_19573);
nand UO_99 (O_99,N_19874,N_19740);
and UO_100 (O_100,N_19682,N_19962);
xor UO_101 (O_101,N_19522,N_19663);
nand UO_102 (O_102,N_19942,N_19719);
or UO_103 (O_103,N_19722,N_19726);
and UO_104 (O_104,N_19628,N_19911);
and UO_105 (O_105,N_19534,N_19767);
nor UO_106 (O_106,N_19973,N_19609);
xnor UO_107 (O_107,N_19756,N_19764);
xor UO_108 (O_108,N_19549,N_19928);
or UO_109 (O_109,N_19630,N_19945);
xor UO_110 (O_110,N_19955,N_19541);
or UO_111 (O_111,N_19776,N_19881);
or UO_112 (O_112,N_19563,N_19659);
nand UO_113 (O_113,N_19596,N_19553);
xnor UO_114 (O_114,N_19620,N_19612);
and UO_115 (O_115,N_19963,N_19909);
and UO_116 (O_116,N_19979,N_19643);
and UO_117 (O_117,N_19798,N_19736);
or UO_118 (O_118,N_19706,N_19936);
nor UO_119 (O_119,N_19896,N_19516);
and UO_120 (O_120,N_19940,N_19968);
xor UO_121 (O_121,N_19843,N_19557);
and UO_122 (O_122,N_19669,N_19780);
nand UO_123 (O_123,N_19692,N_19855);
nand UO_124 (O_124,N_19577,N_19552);
nand UO_125 (O_125,N_19752,N_19714);
and UO_126 (O_126,N_19503,N_19632);
or UO_127 (O_127,N_19701,N_19568);
or UO_128 (O_128,N_19781,N_19603);
xor UO_129 (O_129,N_19747,N_19546);
or UO_130 (O_130,N_19758,N_19922);
nor UO_131 (O_131,N_19613,N_19586);
nor UO_132 (O_132,N_19914,N_19592);
or UO_133 (O_133,N_19830,N_19806);
and UO_134 (O_134,N_19803,N_19951);
and UO_135 (O_135,N_19572,N_19766);
nor UO_136 (O_136,N_19782,N_19550);
nand UO_137 (O_137,N_19652,N_19560);
nor UO_138 (O_138,N_19696,N_19571);
or UO_139 (O_139,N_19753,N_19921);
and UO_140 (O_140,N_19731,N_19551);
and UO_141 (O_141,N_19977,N_19788);
nand UO_142 (O_142,N_19858,N_19957);
nor UO_143 (O_143,N_19500,N_19888);
xor UO_144 (O_144,N_19644,N_19604);
and UO_145 (O_145,N_19966,N_19967);
nand UO_146 (O_146,N_19810,N_19728);
nor UO_147 (O_147,N_19856,N_19994);
and UO_148 (O_148,N_19800,N_19742);
or UO_149 (O_149,N_19793,N_19838);
or UO_150 (O_150,N_19897,N_19567);
xnor UO_151 (O_151,N_19750,N_19831);
or UO_152 (O_152,N_19819,N_19884);
nand UO_153 (O_153,N_19580,N_19575);
xnor UO_154 (O_154,N_19733,N_19882);
xor UO_155 (O_155,N_19600,N_19916);
and UO_156 (O_156,N_19543,N_19576);
nor UO_157 (O_157,N_19992,N_19585);
and UO_158 (O_158,N_19762,N_19626);
nor UO_159 (O_159,N_19777,N_19531);
or UO_160 (O_160,N_19948,N_19691);
nand UO_161 (O_161,N_19569,N_19883);
nand UO_162 (O_162,N_19870,N_19676);
nor UO_163 (O_163,N_19918,N_19857);
nor UO_164 (O_164,N_19970,N_19617);
nor UO_165 (O_165,N_19813,N_19960);
or UO_166 (O_166,N_19670,N_19507);
xnor UO_167 (O_167,N_19828,N_19537);
nand UO_168 (O_168,N_19933,N_19959);
xor UO_169 (O_169,N_19712,N_19627);
and UO_170 (O_170,N_19761,N_19658);
nand UO_171 (O_171,N_19698,N_19702);
and UO_172 (O_172,N_19873,N_19846);
nand UO_173 (O_173,N_19605,N_19783);
xnor UO_174 (O_174,N_19859,N_19622);
and UO_175 (O_175,N_19589,N_19672);
nand UO_176 (O_176,N_19812,N_19899);
nor UO_177 (O_177,N_19974,N_19619);
and UO_178 (O_178,N_19527,N_19787);
xor UO_179 (O_179,N_19852,N_19792);
and UO_180 (O_180,N_19651,N_19934);
and UO_181 (O_181,N_19594,N_19678);
xor UO_182 (O_182,N_19749,N_19885);
and UO_183 (O_183,N_19949,N_19635);
nand UO_184 (O_184,N_19763,N_19990);
xor UO_185 (O_185,N_19842,N_19695);
or UO_186 (O_186,N_19528,N_19755);
nor UO_187 (O_187,N_19590,N_19946);
nand UO_188 (O_188,N_19924,N_19775);
and UO_189 (O_189,N_19802,N_19853);
nand UO_190 (O_190,N_19912,N_19907);
xnor UO_191 (O_191,N_19801,N_19505);
nor UO_192 (O_192,N_19709,N_19765);
nand UO_193 (O_193,N_19624,N_19849);
nor UO_194 (O_194,N_19910,N_19978);
xor UO_195 (O_195,N_19715,N_19894);
xnor UO_196 (O_196,N_19511,N_19759);
nand UO_197 (O_197,N_19732,N_19774);
xnor UO_198 (O_198,N_19521,N_19542);
or UO_199 (O_199,N_19502,N_19771);
or UO_200 (O_200,N_19653,N_19744);
xor UO_201 (O_201,N_19579,N_19661);
or UO_202 (O_202,N_19646,N_19923);
nand UO_203 (O_203,N_19848,N_19547);
and UO_204 (O_204,N_19539,N_19581);
nand UO_205 (O_205,N_19898,N_19915);
nand UO_206 (O_206,N_19902,N_19679);
and UO_207 (O_207,N_19633,N_19610);
and UO_208 (O_208,N_19935,N_19964);
xnor UO_209 (O_209,N_19556,N_19804);
nor UO_210 (O_210,N_19588,N_19958);
nor UO_211 (O_211,N_19981,N_19582);
or UO_212 (O_212,N_19694,N_19926);
or UO_213 (O_213,N_19637,N_19720);
nand UO_214 (O_214,N_19574,N_19772);
and UO_215 (O_215,N_19984,N_19903);
xor UO_216 (O_216,N_19561,N_19689);
and UO_217 (O_217,N_19956,N_19508);
xnor UO_218 (O_218,N_19818,N_19673);
and UO_219 (O_219,N_19649,N_19880);
or UO_220 (O_220,N_19524,N_19972);
nor UO_221 (O_221,N_19844,N_19904);
nand UO_222 (O_222,N_19746,N_19835);
and UO_223 (O_223,N_19583,N_19741);
and UO_224 (O_224,N_19939,N_19625);
nor UO_225 (O_225,N_19837,N_19536);
nand UO_226 (O_226,N_19523,N_19570);
nor UO_227 (O_227,N_19930,N_19558);
or UO_228 (O_228,N_19545,N_19789);
nor UO_229 (O_229,N_19784,N_19530);
and UO_230 (O_230,N_19827,N_19727);
nor UO_231 (O_231,N_19841,N_19891);
or UO_232 (O_232,N_19634,N_19999);
nor UO_233 (O_233,N_19725,N_19564);
and UO_234 (O_234,N_19667,N_19769);
nand UO_235 (O_235,N_19929,N_19820);
and UO_236 (O_236,N_19745,N_19662);
xnor UO_237 (O_237,N_19566,N_19690);
xnor UO_238 (O_238,N_19824,N_19797);
xnor UO_239 (O_239,N_19532,N_19647);
nor UO_240 (O_240,N_19687,N_19836);
nand UO_241 (O_241,N_19943,N_19501);
or UO_242 (O_242,N_19639,N_19730);
or UO_243 (O_243,N_19548,N_19811);
or UO_244 (O_244,N_19515,N_19606);
nor UO_245 (O_245,N_19875,N_19703);
nor UO_246 (O_246,N_19629,N_19734);
nand UO_247 (O_247,N_19640,N_19660);
and UO_248 (O_248,N_19638,N_19890);
and UO_249 (O_249,N_19786,N_19711);
and UO_250 (O_250,N_19914,N_19730);
or UO_251 (O_251,N_19567,N_19784);
nor UO_252 (O_252,N_19800,N_19861);
or UO_253 (O_253,N_19943,N_19762);
xnor UO_254 (O_254,N_19895,N_19751);
or UO_255 (O_255,N_19508,N_19721);
nor UO_256 (O_256,N_19738,N_19681);
or UO_257 (O_257,N_19502,N_19845);
nor UO_258 (O_258,N_19781,N_19688);
nor UO_259 (O_259,N_19549,N_19683);
nor UO_260 (O_260,N_19739,N_19750);
or UO_261 (O_261,N_19512,N_19849);
xnor UO_262 (O_262,N_19880,N_19893);
or UO_263 (O_263,N_19621,N_19995);
xor UO_264 (O_264,N_19871,N_19528);
nor UO_265 (O_265,N_19658,N_19627);
nand UO_266 (O_266,N_19944,N_19524);
xor UO_267 (O_267,N_19944,N_19742);
xor UO_268 (O_268,N_19717,N_19707);
and UO_269 (O_269,N_19990,N_19929);
and UO_270 (O_270,N_19865,N_19721);
nor UO_271 (O_271,N_19839,N_19790);
nor UO_272 (O_272,N_19537,N_19658);
nor UO_273 (O_273,N_19580,N_19788);
nand UO_274 (O_274,N_19721,N_19510);
and UO_275 (O_275,N_19565,N_19501);
and UO_276 (O_276,N_19930,N_19621);
nand UO_277 (O_277,N_19803,N_19866);
nand UO_278 (O_278,N_19611,N_19814);
nand UO_279 (O_279,N_19533,N_19918);
nor UO_280 (O_280,N_19674,N_19997);
and UO_281 (O_281,N_19582,N_19529);
nor UO_282 (O_282,N_19562,N_19748);
and UO_283 (O_283,N_19670,N_19772);
xnor UO_284 (O_284,N_19620,N_19721);
xor UO_285 (O_285,N_19928,N_19618);
xor UO_286 (O_286,N_19978,N_19686);
nand UO_287 (O_287,N_19723,N_19683);
or UO_288 (O_288,N_19586,N_19898);
and UO_289 (O_289,N_19831,N_19848);
or UO_290 (O_290,N_19840,N_19514);
or UO_291 (O_291,N_19721,N_19934);
nand UO_292 (O_292,N_19601,N_19581);
or UO_293 (O_293,N_19992,N_19625);
nor UO_294 (O_294,N_19773,N_19568);
or UO_295 (O_295,N_19820,N_19705);
nand UO_296 (O_296,N_19639,N_19846);
and UO_297 (O_297,N_19721,N_19626);
and UO_298 (O_298,N_19515,N_19891);
or UO_299 (O_299,N_19926,N_19741);
or UO_300 (O_300,N_19729,N_19984);
or UO_301 (O_301,N_19968,N_19916);
nor UO_302 (O_302,N_19931,N_19594);
and UO_303 (O_303,N_19852,N_19943);
or UO_304 (O_304,N_19563,N_19952);
xnor UO_305 (O_305,N_19651,N_19730);
or UO_306 (O_306,N_19570,N_19502);
and UO_307 (O_307,N_19979,N_19584);
nand UO_308 (O_308,N_19593,N_19536);
xnor UO_309 (O_309,N_19540,N_19898);
xnor UO_310 (O_310,N_19666,N_19635);
and UO_311 (O_311,N_19883,N_19985);
nand UO_312 (O_312,N_19733,N_19605);
nand UO_313 (O_313,N_19978,N_19993);
nor UO_314 (O_314,N_19596,N_19593);
nand UO_315 (O_315,N_19511,N_19633);
and UO_316 (O_316,N_19598,N_19587);
or UO_317 (O_317,N_19892,N_19586);
xor UO_318 (O_318,N_19992,N_19902);
or UO_319 (O_319,N_19574,N_19704);
nand UO_320 (O_320,N_19728,N_19884);
nand UO_321 (O_321,N_19933,N_19745);
or UO_322 (O_322,N_19936,N_19524);
nand UO_323 (O_323,N_19925,N_19679);
nand UO_324 (O_324,N_19984,N_19770);
nand UO_325 (O_325,N_19729,N_19850);
xnor UO_326 (O_326,N_19653,N_19683);
xor UO_327 (O_327,N_19871,N_19758);
or UO_328 (O_328,N_19812,N_19648);
or UO_329 (O_329,N_19611,N_19588);
and UO_330 (O_330,N_19874,N_19702);
or UO_331 (O_331,N_19801,N_19869);
and UO_332 (O_332,N_19730,N_19519);
nor UO_333 (O_333,N_19657,N_19727);
or UO_334 (O_334,N_19821,N_19901);
or UO_335 (O_335,N_19543,N_19961);
and UO_336 (O_336,N_19804,N_19765);
nor UO_337 (O_337,N_19524,N_19814);
nor UO_338 (O_338,N_19639,N_19802);
xor UO_339 (O_339,N_19963,N_19560);
nand UO_340 (O_340,N_19764,N_19901);
and UO_341 (O_341,N_19982,N_19536);
and UO_342 (O_342,N_19736,N_19941);
and UO_343 (O_343,N_19655,N_19692);
or UO_344 (O_344,N_19954,N_19725);
and UO_345 (O_345,N_19514,N_19575);
nand UO_346 (O_346,N_19738,N_19955);
nor UO_347 (O_347,N_19857,N_19665);
and UO_348 (O_348,N_19825,N_19813);
nor UO_349 (O_349,N_19782,N_19878);
xor UO_350 (O_350,N_19578,N_19612);
xnor UO_351 (O_351,N_19810,N_19642);
and UO_352 (O_352,N_19963,N_19890);
nand UO_353 (O_353,N_19771,N_19663);
nand UO_354 (O_354,N_19509,N_19784);
or UO_355 (O_355,N_19787,N_19934);
and UO_356 (O_356,N_19704,N_19575);
and UO_357 (O_357,N_19997,N_19695);
xor UO_358 (O_358,N_19632,N_19793);
or UO_359 (O_359,N_19822,N_19955);
and UO_360 (O_360,N_19722,N_19731);
nor UO_361 (O_361,N_19771,N_19854);
nand UO_362 (O_362,N_19892,N_19710);
nor UO_363 (O_363,N_19751,N_19730);
nand UO_364 (O_364,N_19605,N_19881);
xnor UO_365 (O_365,N_19829,N_19696);
nor UO_366 (O_366,N_19682,N_19634);
nor UO_367 (O_367,N_19950,N_19808);
nor UO_368 (O_368,N_19964,N_19745);
and UO_369 (O_369,N_19743,N_19597);
or UO_370 (O_370,N_19580,N_19675);
xor UO_371 (O_371,N_19886,N_19657);
and UO_372 (O_372,N_19503,N_19842);
and UO_373 (O_373,N_19830,N_19582);
nand UO_374 (O_374,N_19597,N_19666);
nand UO_375 (O_375,N_19890,N_19907);
xor UO_376 (O_376,N_19588,N_19722);
and UO_377 (O_377,N_19770,N_19691);
and UO_378 (O_378,N_19904,N_19966);
and UO_379 (O_379,N_19602,N_19975);
or UO_380 (O_380,N_19866,N_19767);
xor UO_381 (O_381,N_19659,N_19517);
nand UO_382 (O_382,N_19946,N_19657);
or UO_383 (O_383,N_19647,N_19803);
nand UO_384 (O_384,N_19723,N_19867);
or UO_385 (O_385,N_19792,N_19880);
nand UO_386 (O_386,N_19661,N_19810);
nand UO_387 (O_387,N_19992,N_19731);
and UO_388 (O_388,N_19677,N_19579);
and UO_389 (O_389,N_19581,N_19608);
nand UO_390 (O_390,N_19781,N_19575);
and UO_391 (O_391,N_19878,N_19918);
nand UO_392 (O_392,N_19626,N_19529);
or UO_393 (O_393,N_19818,N_19883);
or UO_394 (O_394,N_19716,N_19683);
and UO_395 (O_395,N_19675,N_19747);
nand UO_396 (O_396,N_19836,N_19863);
or UO_397 (O_397,N_19712,N_19520);
nand UO_398 (O_398,N_19530,N_19501);
nand UO_399 (O_399,N_19811,N_19880);
or UO_400 (O_400,N_19544,N_19808);
or UO_401 (O_401,N_19918,N_19566);
or UO_402 (O_402,N_19794,N_19535);
and UO_403 (O_403,N_19693,N_19776);
xnor UO_404 (O_404,N_19534,N_19594);
or UO_405 (O_405,N_19852,N_19544);
and UO_406 (O_406,N_19704,N_19841);
xnor UO_407 (O_407,N_19545,N_19523);
xor UO_408 (O_408,N_19735,N_19773);
nand UO_409 (O_409,N_19694,N_19995);
and UO_410 (O_410,N_19970,N_19919);
nor UO_411 (O_411,N_19669,N_19685);
nor UO_412 (O_412,N_19830,N_19846);
nand UO_413 (O_413,N_19758,N_19564);
nand UO_414 (O_414,N_19518,N_19582);
and UO_415 (O_415,N_19586,N_19951);
xnor UO_416 (O_416,N_19798,N_19869);
nand UO_417 (O_417,N_19961,N_19774);
xor UO_418 (O_418,N_19648,N_19568);
or UO_419 (O_419,N_19664,N_19767);
nand UO_420 (O_420,N_19550,N_19852);
or UO_421 (O_421,N_19703,N_19795);
and UO_422 (O_422,N_19681,N_19617);
or UO_423 (O_423,N_19976,N_19865);
nand UO_424 (O_424,N_19920,N_19555);
and UO_425 (O_425,N_19789,N_19928);
nor UO_426 (O_426,N_19683,N_19863);
nor UO_427 (O_427,N_19875,N_19934);
nand UO_428 (O_428,N_19763,N_19688);
xnor UO_429 (O_429,N_19616,N_19820);
xnor UO_430 (O_430,N_19773,N_19810);
xnor UO_431 (O_431,N_19976,N_19629);
and UO_432 (O_432,N_19981,N_19640);
and UO_433 (O_433,N_19689,N_19630);
and UO_434 (O_434,N_19613,N_19782);
xor UO_435 (O_435,N_19892,N_19558);
xor UO_436 (O_436,N_19882,N_19619);
and UO_437 (O_437,N_19978,N_19651);
nand UO_438 (O_438,N_19680,N_19608);
or UO_439 (O_439,N_19691,N_19794);
nand UO_440 (O_440,N_19512,N_19810);
nand UO_441 (O_441,N_19893,N_19602);
or UO_442 (O_442,N_19913,N_19696);
or UO_443 (O_443,N_19815,N_19746);
nand UO_444 (O_444,N_19583,N_19658);
or UO_445 (O_445,N_19693,N_19723);
xor UO_446 (O_446,N_19753,N_19733);
xnor UO_447 (O_447,N_19514,N_19928);
or UO_448 (O_448,N_19819,N_19906);
and UO_449 (O_449,N_19875,N_19546);
nor UO_450 (O_450,N_19888,N_19533);
or UO_451 (O_451,N_19776,N_19510);
or UO_452 (O_452,N_19588,N_19703);
or UO_453 (O_453,N_19872,N_19657);
and UO_454 (O_454,N_19925,N_19943);
or UO_455 (O_455,N_19826,N_19531);
xor UO_456 (O_456,N_19792,N_19500);
and UO_457 (O_457,N_19573,N_19886);
nor UO_458 (O_458,N_19923,N_19558);
or UO_459 (O_459,N_19649,N_19932);
nor UO_460 (O_460,N_19899,N_19807);
or UO_461 (O_461,N_19795,N_19651);
or UO_462 (O_462,N_19524,N_19558);
xnor UO_463 (O_463,N_19893,N_19617);
and UO_464 (O_464,N_19640,N_19518);
xnor UO_465 (O_465,N_19550,N_19938);
xor UO_466 (O_466,N_19702,N_19826);
or UO_467 (O_467,N_19733,N_19876);
nor UO_468 (O_468,N_19996,N_19581);
xor UO_469 (O_469,N_19777,N_19811);
nor UO_470 (O_470,N_19506,N_19934);
xnor UO_471 (O_471,N_19560,N_19832);
or UO_472 (O_472,N_19828,N_19602);
nand UO_473 (O_473,N_19923,N_19653);
and UO_474 (O_474,N_19646,N_19861);
nand UO_475 (O_475,N_19889,N_19845);
or UO_476 (O_476,N_19615,N_19647);
and UO_477 (O_477,N_19551,N_19700);
xnor UO_478 (O_478,N_19799,N_19995);
xor UO_479 (O_479,N_19936,N_19629);
or UO_480 (O_480,N_19658,N_19871);
or UO_481 (O_481,N_19520,N_19813);
xor UO_482 (O_482,N_19822,N_19995);
or UO_483 (O_483,N_19912,N_19766);
nand UO_484 (O_484,N_19810,N_19591);
xnor UO_485 (O_485,N_19557,N_19904);
nor UO_486 (O_486,N_19872,N_19708);
nor UO_487 (O_487,N_19790,N_19569);
nand UO_488 (O_488,N_19818,N_19750);
nor UO_489 (O_489,N_19871,N_19954);
or UO_490 (O_490,N_19691,N_19813);
and UO_491 (O_491,N_19513,N_19644);
nor UO_492 (O_492,N_19850,N_19937);
nor UO_493 (O_493,N_19888,N_19932);
or UO_494 (O_494,N_19689,N_19832);
nand UO_495 (O_495,N_19636,N_19580);
nor UO_496 (O_496,N_19986,N_19702);
nor UO_497 (O_497,N_19609,N_19648);
and UO_498 (O_498,N_19635,N_19627);
and UO_499 (O_499,N_19557,N_19957);
nor UO_500 (O_500,N_19793,N_19575);
nand UO_501 (O_501,N_19870,N_19713);
nor UO_502 (O_502,N_19976,N_19709);
nand UO_503 (O_503,N_19779,N_19945);
nand UO_504 (O_504,N_19609,N_19553);
nor UO_505 (O_505,N_19969,N_19623);
nor UO_506 (O_506,N_19692,N_19830);
or UO_507 (O_507,N_19945,N_19905);
nand UO_508 (O_508,N_19597,N_19595);
nand UO_509 (O_509,N_19738,N_19610);
nand UO_510 (O_510,N_19746,N_19652);
or UO_511 (O_511,N_19807,N_19514);
or UO_512 (O_512,N_19796,N_19927);
and UO_513 (O_513,N_19709,N_19665);
nand UO_514 (O_514,N_19661,N_19734);
or UO_515 (O_515,N_19650,N_19526);
nor UO_516 (O_516,N_19502,N_19679);
nand UO_517 (O_517,N_19611,N_19964);
nor UO_518 (O_518,N_19593,N_19687);
nor UO_519 (O_519,N_19521,N_19924);
nor UO_520 (O_520,N_19990,N_19649);
and UO_521 (O_521,N_19577,N_19900);
or UO_522 (O_522,N_19762,N_19559);
or UO_523 (O_523,N_19592,N_19791);
and UO_524 (O_524,N_19761,N_19672);
xor UO_525 (O_525,N_19989,N_19561);
and UO_526 (O_526,N_19728,N_19613);
nor UO_527 (O_527,N_19975,N_19777);
nand UO_528 (O_528,N_19614,N_19929);
nand UO_529 (O_529,N_19947,N_19684);
or UO_530 (O_530,N_19887,N_19616);
and UO_531 (O_531,N_19864,N_19731);
nand UO_532 (O_532,N_19599,N_19732);
nor UO_533 (O_533,N_19511,N_19906);
and UO_534 (O_534,N_19838,N_19895);
and UO_535 (O_535,N_19793,N_19871);
xnor UO_536 (O_536,N_19976,N_19620);
xnor UO_537 (O_537,N_19979,N_19942);
and UO_538 (O_538,N_19579,N_19942);
or UO_539 (O_539,N_19858,N_19536);
xnor UO_540 (O_540,N_19520,N_19800);
nand UO_541 (O_541,N_19882,N_19801);
nor UO_542 (O_542,N_19548,N_19770);
and UO_543 (O_543,N_19604,N_19832);
xor UO_544 (O_544,N_19695,N_19907);
or UO_545 (O_545,N_19626,N_19562);
xnor UO_546 (O_546,N_19711,N_19585);
or UO_547 (O_547,N_19578,N_19560);
nand UO_548 (O_548,N_19652,N_19520);
or UO_549 (O_549,N_19931,N_19712);
xor UO_550 (O_550,N_19885,N_19960);
nor UO_551 (O_551,N_19971,N_19774);
or UO_552 (O_552,N_19988,N_19778);
or UO_553 (O_553,N_19800,N_19690);
xnor UO_554 (O_554,N_19534,N_19791);
nor UO_555 (O_555,N_19624,N_19536);
nor UO_556 (O_556,N_19726,N_19983);
and UO_557 (O_557,N_19972,N_19856);
nand UO_558 (O_558,N_19567,N_19800);
and UO_559 (O_559,N_19596,N_19579);
nand UO_560 (O_560,N_19819,N_19638);
xor UO_561 (O_561,N_19956,N_19911);
nor UO_562 (O_562,N_19633,N_19864);
nand UO_563 (O_563,N_19609,N_19513);
nand UO_564 (O_564,N_19848,N_19970);
or UO_565 (O_565,N_19636,N_19593);
nor UO_566 (O_566,N_19680,N_19631);
and UO_567 (O_567,N_19707,N_19547);
or UO_568 (O_568,N_19589,N_19601);
nor UO_569 (O_569,N_19687,N_19652);
xor UO_570 (O_570,N_19923,N_19760);
xor UO_571 (O_571,N_19617,N_19531);
nor UO_572 (O_572,N_19865,N_19556);
nand UO_573 (O_573,N_19623,N_19851);
nand UO_574 (O_574,N_19733,N_19746);
xnor UO_575 (O_575,N_19668,N_19759);
nand UO_576 (O_576,N_19888,N_19722);
or UO_577 (O_577,N_19963,N_19608);
nand UO_578 (O_578,N_19931,N_19510);
xnor UO_579 (O_579,N_19724,N_19684);
or UO_580 (O_580,N_19998,N_19905);
nand UO_581 (O_581,N_19894,N_19801);
and UO_582 (O_582,N_19640,N_19950);
nand UO_583 (O_583,N_19630,N_19855);
or UO_584 (O_584,N_19733,N_19720);
xor UO_585 (O_585,N_19750,N_19982);
xnor UO_586 (O_586,N_19763,N_19891);
and UO_587 (O_587,N_19556,N_19812);
and UO_588 (O_588,N_19637,N_19915);
and UO_589 (O_589,N_19938,N_19628);
and UO_590 (O_590,N_19596,N_19800);
xnor UO_591 (O_591,N_19961,N_19549);
and UO_592 (O_592,N_19720,N_19950);
and UO_593 (O_593,N_19980,N_19732);
or UO_594 (O_594,N_19643,N_19869);
and UO_595 (O_595,N_19576,N_19694);
and UO_596 (O_596,N_19906,N_19796);
xor UO_597 (O_597,N_19554,N_19536);
and UO_598 (O_598,N_19610,N_19540);
and UO_599 (O_599,N_19955,N_19596);
or UO_600 (O_600,N_19822,N_19842);
nand UO_601 (O_601,N_19582,N_19689);
nor UO_602 (O_602,N_19557,N_19739);
or UO_603 (O_603,N_19814,N_19607);
and UO_604 (O_604,N_19754,N_19524);
nand UO_605 (O_605,N_19897,N_19889);
nor UO_606 (O_606,N_19780,N_19931);
nor UO_607 (O_607,N_19768,N_19859);
nor UO_608 (O_608,N_19772,N_19798);
and UO_609 (O_609,N_19940,N_19505);
xnor UO_610 (O_610,N_19512,N_19721);
xor UO_611 (O_611,N_19588,N_19693);
xor UO_612 (O_612,N_19944,N_19928);
or UO_613 (O_613,N_19908,N_19864);
nand UO_614 (O_614,N_19833,N_19888);
or UO_615 (O_615,N_19997,N_19970);
and UO_616 (O_616,N_19528,N_19832);
xor UO_617 (O_617,N_19543,N_19518);
nor UO_618 (O_618,N_19747,N_19637);
nand UO_619 (O_619,N_19510,N_19521);
and UO_620 (O_620,N_19968,N_19701);
nand UO_621 (O_621,N_19636,N_19648);
nand UO_622 (O_622,N_19772,N_19572);
nand UO_623 (O_623,N_19550,N_19610);
xor UO_624 (O_624,N_19935,N_19984);
and UO_625 (O_625,N_19651,N_19519);
nor UO_626 (O_626,N_19522,N_19628);
and UO_627 (O_627,N_19784,N_19524);
nand UO_628 (O_628,N_19735,N_19924);
xnor UO_629 (O_629,N_19605,N_19702);
nor UO_630 (O_630,N_19733,N_19842);
and UO_631 (O_631,N_19812,N_19505);
nor UO_632 (O_632,N_19800,N_19552);
or UO_633 (O_633,N_19699,N_19857);
xor UO_634 (O_634,N_19970,N_19758);
or UO_635 (O_635,N_19858,N_19857);
nand UO_636 (O_636,N_19592,N_19569);
or UO_637 (O_637,N_19690,N_19508);
and UO_638 (O_638,N_19622,N_19878);
or UO_639 (O_639,N_19879,N_19837);
or UO_640 (O_640,N_19514,N_19714);
or UO_641 (O_641,N_19579,N_19912);
nand UO_642 (O_642,N_19750,N_19808);
or UO_643 (O_643,N_19966,N_19734);
nor UO_644 (O_644,N_19733,N_19891);
nor UO_645 (O_645,N_19820,N_19801);
nor UO_646 (O_646,N_19778,N_19979);
nor UO_647 (O_647,N_19982,N_19937);
xnor UO_648 (O_648,N_19991,N_19772);
xnor UO_649 (O_649,N_19864,N_19607);
and UO_650 (O_650,N_19760,N_19670);
nand UO_651 (O_651,N_19959,N_19575);
and UO_652 (O_652,N_19922,N_19854);
nand UO_653 (O_653,N_19605,N_19999);
or UO_654 (O_654,N_19628,N_19884);
xnor UO_655 (O_655,N_19636,N_19630);
or UO_656 (O_656,N_19914,N_19688);
and UO_657 (O_657,N_19819,N_19863);
and UO_658 (O_658,N_19748,N_19710);
or UO_659 (O_659,N_19823,N_19936);
and UO_660 (O_660,N_19894,N_19531);
or UO_661 (O_661,N_19887,N_19768);
nand UO_662 (O_662,N_19535,N_19956);
nor UO_663 (O_663,N_19552,N_19505);
nor UO_664 (O_664,N_19790,N_19726);
and UO_665 (O_665,N_19509,N_19964);
or UO_666 (O_666,N_19913,N_19633);
xor UO_667 (O_667,N_19866,N_19796);
xor UO_668 (O_668,N_19549,N_19657);
nand UO_669 (O_669,N_19832,N_19974);
nand UO_670 (O_670,N_19841,N_19933);
and UO_671 (O_671,N_19765,N_19878);
and UO_672 (O_672,N_19954,N_19589);
nor UO_673 (O_673,N_19727,N_19687);
nor UO_674 (O_674,N_19594,N_19716);
xor UO_675 (O_675,N_19624,N_19576);
nand UO_676 (O_676,N_19814,N_19726);
or UO_677 (O_677,N_19526,N_19614);
or UO_678 (O_678,N_19927,N_19959);
nand UO_679 (O_679,N_19842,N_19941);
xor UO_680 (O_680,N_19922,N_19720);
nor UO_681 (O_681,N_19979,N_19746);
xnor UO_682 (O_682,N_19727,N_19867);
xor UO_683 (O_683,N_19880,N_19664);
and UO_684 (O_684,N_19770,N_19906);
nor UO_685 (O_685,N_19510,N_19574);
xor UO_686 (O_686,N_19505,N_19882);
nand UO_687 (O_687,N_19519,N_19540);
nand UO_688 (O_688,N_19745,N_19582);
and UO_689 (O_689,N_19611,N_19764);
nor UO_690 (O_690,N_19537,N_19504);
and UO_691 (O_691,N_19504,N_19708);
and UO_692 (O_692,N_19696,N_19503);
and UO_693 (O_693,N_19641,N_19932);
nand UO_694 (O_694,N_19750,N_19733);
nand UO_695 (O_695,N_19799,N_19803);
and UO_696 (O_696,N_19654,N_19777);
nand UO_697 (O_697,N_19573,N_19869);
or UO_698 (O_698,N_19769,N_19607);
xor UO_699 (O_699,N_19938,N_19976);
or UO_700 (O_700,N_19690,N_19655);
xnor UO_701 (O_701,N_19693,N_19533);
or UO_702 (O_702,N_19865,N_19815);
nor UO_703 (O_703,N_19908,N_19517);
nand UO_704 (O_704,N_19848,N_19732);
or UO_705 (O_705,N_19508,N_19817);
xor UO_706 (O_706,N_19968,N_19608);
nor UO_707 (O_707,N_19592,N_19651);
or UO_708 (O_708,N_19948,N_19937);
and UO_709 (O_709,N_19885,N_19991);
and UO_710 (O_710,N_19888,N_19703);
and UO_711 (O_711,N_19818,N_19978);
and UO_712 (O_712,N_19505,N_19617);
or UO_713 (O_713,N_19716,N_19581);
and UO_714 (O_714,N_19568,N_19915);
xnor UO_715 (O_715,N_19734,N_19876);
or UO_716 (O_716,N_19918,N_19742);
and UO_717 (O_717,N_19677,N_19671);
or UO_718 (O_718,N_19758,N_19890);
nor UO_719 (O_719,N_19708,N_19764);
nand UO_720 (O_720,N_19569,N_19502);
and UO_721 (O_721,N_19880,N_19814);
or UO_722 (O_722,N_19522,N_19793);
or UO_723 (O_723,N_19939,N_19869);
nand UO_724 (O_724,N_19529,N_19894);
and UO_725 (O_725,N_19635,N_19976);
and UO_726 (O_726,N_19958,N_19566);
or UO_727 (O_727,N_19834,N_19724);
nor UO_728 (O_728,N_19779,N_19525);
and UO_729 (O_729,N_19838,N_19999);
and UO_730 (O_730,N_19846,N_19990);
or UO_731 (O_731,N_19533,N_19919);
nor UO_732 (O_732,N_19732,N_19853);
nor UO_733 (O_733,N_19684,N_19591);
nand UO_734 (O_734,N_19859,N_19980);
xor UO_735 (O_735,N_19621,N_19993);
xor UO_736 (O_736,N_19847,N_19903);
and UO_737 (O_737,N_19702,N_19870);
or UO_738 (O_738,N_19891,N_19980);
and UO_739 (O_739,N_19561,N_19891);
xor UO_740 (O_740,N_19942,N_19682);
and UO_741 (O_741,N_19953,N_19945);
and UO_742 (O_742,N_19982,N_19527);
nand UO_743 (O_743,N_19666,N_19773);
nor UO_744 (O_744,N_19567,N_19795);
xor UO_745 (O_745,N_19851,N_19732);
and UO_746 (O_746,N_19683,N_19996);
and UO_747 (O_747,N_19605,N_19714);
or UO_748 (O_748,N_19648,N_19999);
xnor UO_749 (O_749,N_19730,N_19839);
and UO_750 (O_750,N_19688,N_19894);
and UO_751 (O_751,N_19971,N_19873);
nor UO_752 (O_752,N_19922,N_19592);
or UO_753 (O_753,N_19805,N_19970);
and UO_754 (O_754,N_19787,N_19562);
and UO_755 (O_755,N_19639,N_19996);
and UO_756 (O_756,N_19578,N_19658);
or UO_757 (O_757,N_19958,N_19664);
or UO_758 (O_758,N_19500,N_19514);
nand UO_759 (O_759,N_19903,N_19775);
or UO_760 (O_760,N_19898,N_19767);
xnor UO_761 (O_761,N_19759,N_19947);
nand UO_762 (O_762,N_19897,N_19689);
or UO_763 (O_763,N_19966,N_19836);
xor UO_764 (O_764,N_19992,N_19606);
or UO_765 (O_765,N_19632,N_19825);
and UO_766 (O_766,N_19929,N_19655);
or UO_767 (O_767,N_19949,N_19817);
and UO_768 (O_768,N_19504,N_19649);
xnor UO_769 (O_769,N_19943,N_19648);
nand UO_770 (O_770,N_19540,N_19756);
nor UO_771 (O_771,N_19740,N_19914);
xor UO_772 (O_772,N_19575,N_19780);
nand UO_773 (O_773,N_19984,N_19835);
and UO_774 (O_774,N_19803,N_19540);
and UO_775 (O_775,N_19828,N_19610);
or UO_776 (O_776,N_19934,N_19765);
nor UO_777 (O_777,N_19852,N_19770);
xnor UO_778 (O_778,N_19594,N_19997);
nand UO_779 (O_779,N_19635,N_19785);
or UO_780 (O_780,N_19811,N_19919);
xnor UO_781 (O_781,N_19646,N_19831);
or UO_782 (O_782,N_19804,N_19571);
xnor UO_783 (O_783,N_19800,N_19509);
xor UO_784 (O_784,N_19838,N_19780);
nor UO_785 (O_785,N_19984,N_19979);
xnor UO_786 (O_786,N_19881,N_19503);
nand UO_787 (O_787,N_19574,N_19699);
xnor UO_788 (O_788,N_19978,N_19529);
and UO_789 (O_789,N_19926,N_19871);
nand UO_790 (O_790,N_19767,N_19665);
nand UO_791 (O_791,N_19807,N_19519);
nand UO_792 (O_792,N_19895,N_19932);
nor UO_793 (O_793,N_19567,N_19524);
and UO_794 (O_794,N_19933,N_19697);
xnor UO_795 (O_795,N_19685,N_19767);
nor UO_796 (O_796,N_19537,N_19531);
nor UO_797 (O_797,N_19719,N_19876);
xor UO_798 (O_798,N_19957,N_19905);
and UO_799 (O_799,N_19503,N_19713);
and UO_800 (O_800,N_19640,N_19910);
or UO_801 (O_801,N_19671,N_19923);
nand UO_802 (O_802,N_19688,N_19954);
and UO_803 (O_803,N_19553,N_19587);
or UO_804 (O_804,N_19690,N_19674);
xnor UO_805 (O_805,N_19767,N_19835);
and UO_806 (O_806,N_19707,N_19542);
nand UO_807 (O_807,N_19663,N_19646);
nor UO_808 (O_808,N_19532,N_19758);
xor UO_809 (O_809,N_19519,N_19579);
nor UO_810 (O_810,N_19648,N_19929);
and UO_811 (O_811,N_19642,N_19680);
xor UO_812 (O_812,N_19869,N_19706);
nand UO_813 (O_813,N_19769,N_19900);
nor UO_814 (O_814,N_19621,N_19853);
or UO_815 (O_815,N_19829,N_19513);
and UO_816 (O_816,N_19659,N_19871);
and UO_817 (O_817,N_19892,N_19624);
or UO_818 (O_818,N_19819,N_19568);
nand UO_819 (O_819,N_19554,N_19746);
and UO_820 (O_820,N_19865,N_19656);
or UO_821 (O_821,N_19599,N_19950);
xnor UO_822 (O_822,N_19974,N_19730);
nor UO_823 (O_823,N_19692,N_19671);
xor UO_824 (O_824,N_19746,N_19593);
and UO_825 (O_825,N_19770,N_19600);
or UO_826 (O_826,N_19717,N_19712);
or UO_827 (O_827,N_19747,N_19814);
nand UO_828 (O_828,N_19883,N_19754);
xnor UO_829 (O_829,N_19759,N_19732);
or UO_830 (O_830,N_19574,N_19886);
nor UO_831 (O_831,N_19853,N_19885);
and UO_832 (O_832,N_19674,N_19744);
nand UO_833 (O_833,N_19715,N_19702);
nand UO_834 (O_834,N_19805,N_19600);
nand UO_835 (O_835,N_19989,N_19616);
nand UO_836 (O_836,N_19871,N_19975);
and UO_837 (O_837,N_19579,N_19512);
or UO_838 (O_838,N_19533,N_19698);
nor UO_839 (O_839,N_19698,N_19873);
nor UO_840 (O_840,N_19989,N_19792);
nor UO_841 (O_841,N_19977,N_19581);
xor UO_842 (O_842,N_19593,N_19800);
and UO_843 (O_843,N_19586,N_19814);
and UO_844 (O_844,N_19746,N_19745);
or UO_845 (O_845,N_19513,N_19956);
or UO_846 (O_846,N_19705,N_19758);
xor UO_847 (O_847,N_19597,N_19570);
xor UO_848 (O_848,N_19593,N_19932);
xor UO_849 (O_849,N_19837,N_19514);
or UO_850 (O_850,N_19734,N_19820);
xnor UO_851 (O_851,N_19760,N_19675);
xor UO_852 (O_852,N_19578,N_19584);
or UO_853 (O_853,N_19861,N_19745);
xnor UO_854 (O_854,N_19913,N_19771);
and UO_855 (O_855,N_19612,N_19957);
and UO_856 (O_856,N_19920,N_19811);
nor UO_857 (O_857,N_19911,N_19887);
nand UO_858 (O_858,N_19616,N_19966);
xor UO_859 (O_859,N_19761,N_19934);
xor UO_860 (O_860,N_19663,N_19926);
or UO_861 (O_861,N_19964,N_19851);
or UO_862 (O_862,N_19523,N_19816);
xnor UO_863 (O_863,N_19710,N_19642);
and UO_864 (O_864,N_19663,N_19742);
nor UO_865 (O_865,N_19991,N_19635);
nand UO_866 (O_866,N_19982,N_19864);
xor UO_867 (O_867,N_19512,N_19785);
nor UO_868 (O_868,N_19944,N_19694);
nor UO_869 (O_869,N_19802,N_19553);
nor UO_870 (O_870,N_19753,N_19844);
and UO_871 (O_871,N_19580,N_19811);
nor UO_872 (O_872,N_19988,N_19812);
and UO_873 (O_873,N_19928,N_19699);
or UO_874 (O_874,N_19688,N_19730);
nor UO_875 (O_875,N_19692,N_19577);
xor UO_876 (O_876,N_19911,N_19933);
and UO_877 (O_877,N_19541,N_19888);
nor UO_878 (O_878,N_19962,N_19716);
and UO_879 (O_879,N_19840,N_19686);
nand UO_880 (O_880,N_19532,N_19739);
xnor UO_881 (O_881,N_19964,N_19975);
and UO_882 (O_882,N_19552,N_19657);
or UO_883 (O_883,N_19571,N_19745);
or UO_884 (O_884,N_19957,N_19598);
xnor UO_885 (O_885,N_19891,N_19867);
nand UO_886 (O_886,N_19649,N_19884);
or UO_887 (O_887,N_19928,N_19817);
nand UO_888 (O_888,N_19702,N_19888);
xor UO_889 (O_889,N_19724,N_19837);
xnor UO_890 (O_890,N_19713,N_19977);
nor UO_891 (O_891,N_19814,N_19853);
nand UO_892 (O_892,N_19966,N_19540);
nor UO_893 (O_893,N_19541,N_19564);
and UO_894 (O_894,N_19576,N_19590);
and UO_895 (O_895,N_19758,N_19519);
and UO_896 (O_896,N_19904,N_19563);
nand UO_897 (O_897,N_19692,N_19656);
xnor UO_898 (O_898,N_19898,N_19776);
and UO_899 (O_899,N_19652,N_19730);
nor UO_900 (O_900,N_19980,N_19591);
or UO_901 (O_901,N_19907,N_19952);
nor UO_902 (O_902,N_19880,N_19868);
xnor UO_903 (O_903,N_19961,N_19605);
nor UO_904 (O_904,N_19957,N_19959);
or UO_905 (O_905,N_19563,N_19896);
or UO_906 (O_906,N_19742,N_19698);
xnor UO_907 (O_907,N_19853,N_19675);
nor UO_908 (O_908,N_19743,N_19846);
nor UO_909 (O_909,N_19700,N_19699);
nor UO_910 (O_910,N_19618,N_19932);
nor UO_911 (O_911,N_19912,N_19926);
xor UO_912 (O_912,N_19847,N_19609);
or UO_913 (O_913,N_19945,N_19877);
or UO_914 (O_914,N_19884,N_19814);
nand UO_915 (O_915,N_19928,N_19966);
or UO_916 (O_916,N_19924,N_19580);
nand UO_917 (O_917,N_19860,N_19763);
or UO_918 (O_918,N_19993,N_19933);
nand UO_919 (O_919,N_19799,N_19759);
or UO_920 (O_920,N_19520,N_19877);
or UO_921 (O_921,N_19877,N_19824);
and UO_922 (O_922,N_19714,N_19623);
xor UO_923 (O_923,N_19605,N_19713);
nor UO_924 (O_924,N_19719,N_19626);
nand UO_925 (O_925,N_19895,N_19927);
nand UO_926 (O_926,N_19774,N_19778);
and UO_927 (O_927,N_19907,N_19989);
or UO_928 (O_928,N_19596,N_19533);
nor UO_929 (O_929,N_19974,N_19805);
and UO_930 (O_930,N_19996,N_19713);
nor UO_931 (O_931,N_19949,N_19782);
and UO_932 (O_932,N_19677,N_19981);
xor UO_933 (O_933,N_19942,N_19633);
and UO_934 (O_934,N_19595,N_19976);
nand UO_935 (O_935,N_19508,N_19840);
or UO_936 (O_936,N_19796,N_19647);
nor UO_937 (O_937,N_19630,N_19517);
nor UO_938 (O_938,N_19711,N_19764);
and UO_939 (O_939,N_19723,N_19903);
nor UO_940 (O_940,N_19697,N_19734);
or UO_941 (O_941,N_19831,N_19872);
and UO_942 (O_942,N_19862,N_19640);
nor UO_943 (O_943,N_19880,N_19817);
and UO_944 (O_944,N_19811,N_19657);
nor UO_945 (O_945,N_19609,N_19556);
and UO_946 (O_946,N_19550,N_19828);
nand UO_947 (O_947,N_19873,N_19786);
or UO_948 (O_948,N_19770,N_19904);
xor UO_949 (O_949,N_19624,N_19877);
xnor UO_950 (O_950,N_19774,N_19947);
nor UO_951 (O_951,N_19918,N_19687);
and UO_952 (O_952,N_19720,N_19662);
and UO_953 (O_953,N_19664,N_19832);
nor UO_954 (O_954,N_19623,N_19968);
nor UO_955 (O_955,N_19796,N_19654);
xnor UO_956 (O_956,N_19897,N_19869);
nor UO_957 (O_957,N_19900,N_19973);
nand UO_958 (O_958,N_19603,N_19519);
nor UO_959 (O_959,N_19813,N_19729);
and UO_960 (O_960,N_19691,N_19781);
nand UO_961 (O_961,N_19882,N_19835);
or UO_962 (O_962,N_19683,N_19567);
and UO_963 (O_963,N_19993,N_19926);
and UO_964 (O_964,N_19661,N_19555);
or UO_965 (O_965,N_19897,N_19950);
and UO_966 (O_966,N_19762,N_19551);
and UO_967 (O_967,N_19681,N_19519);
nor UO_968 (O_968,N_19927,N_19723);
nand UO_969 (O_969,N_19930,N_19753);
nand UO_970 (O_970,N_19507,N_19831);
and UO_971 (O_971,N_19732,N_19598);
xor UO_972 (O_972,N_19565,N_19834);
nand UO_973 (O_973,N_19536,N_19950);
nor UO_974 (O_974,N_19940,N_19979);
nor UO_975 (O_975,N_19555,N_19972);
nand UO_976 (O_976,N_19514,N_19919);
xnor UO_977 (O_977,N_19826,N_19845);
and UO_978 (O_978,N_19814,N_19565);
xnor UO_979 (O_979,N_19827,N_19550);
nand UO_980 (O_980,N_19795,N_19825);
nand UO_981 (O_981,N_19522,N_19728);
nor UO_982 (O_982,N_19778,N_19574);
or UO_983 (O_983,N_19984,N_19623);
xor UO_984 (O_984,N_19512,N_19837);
nand UO_985 (O_985,N_19881,N_19662);
nand UO_986 (O_986,N_19690,N_19500);
and UO_987 (O_987,N_19932,N_19952);
and UO_988 (O_988,N_19577,N_19886);
or UO_989 (O_989,N_19582,N_19903);
and UO_990 (O_990,N_19836,N_19866);
xor UO_991 (O_991,N_19733,N_19832);
and UO_992 (O_992,N_19872,N_19551);
nand UO_993 (O_993,N_19949,N_19762);
or UO_994 (O_994,N_19635,N_19756);
nor UO_995 (O_995,N_19846,N_19603);
nor UO_996 (O_996,N_19529,N_19889);
and UO_997 (O_997,N_19780,N_19748);
nor UO_998 (O_998,N_19843,N_19865);
or UO_999 (O_999,N_19553,N_19503);
xnor UO_1000 (O_1000,N_19610,N_19850);
nor UO_1001 (O_1001,N_19927,N_19675);
xnor UO_1002 (O_1002,N_19901,N_19847);
and UO_1003 (O_1003,N_19879,N_19537);
and UO_1004 (O_1004,N_19507,N_19676);
or UO_1005 (O_1005,N_19760,N_19800);
nand UO_1006 (O_1006,N_19863,N_19839);
and UO_1007 (O_1007,N_19568,N_19762);
xnor UO_1008 (O_1008,N_19647,N_19864);
nand UO_1009 (O_1009,N_19961,N_19655);
xor UO_1010 (O_1010,N_19580,N_19592);
nand UO_1011 (O_1011,N_19553,N_19594);
nor UO_1012 (O_1012,N_19589,N_19683);
nor UO_1013 (O_1013,N_19917,N_19834);
nor UO_1014 (O_1014,N_19843,N_19763);
nand UO_1015 (O_1015,N_19514,N_19627);
nor UO_1016 (O_1016,N_19649,N_19572);
nor UO_1017 (O_1017,N_19684,N_19821);
nor UO_1018 (O_1018,N_19884,N_19501);
and UO_1019 (O_1019,N_19502,N_19741);
or UO_1020 (O_1020,N_19853,N_19859);
xnor UO_1021 (O_1021,N_19974,N_19980);
nor UO_1022 (O_1022,N_19830,N_19701);
xor UO_1023 (O_1023,N_19515,N_19943);
nand UO_1024 (O_1024,N_19842,N_19788);
or UO_1025 (O_1025,N_19712,N_19522);
xnor UO_1026 (O_1026,N_19773,N_19585);
or UO_1027 (O_1027,N_19923,N_19836);
xnor UO_1028 (O_1028,N_19827,N_19862);
xor UO_1029 (O_1029,N_19732,N_19625);
xnor UO_1030 (O_1030,N_19689,N_19556);
xor UO_1031 (O_1031,N_19891,N_19886);
or UO_1032 (O_1032,N_19551,N_19740);
nor UO_1033 (O_1033,N_19914,N_19591);
or UO_1034 (O_1034,N_19894,N_19522);
xnor UO_1035 (O_1035,N_19790,N_19912);
nand UO_1036 (O_1036,N_19741,N_19513);
and UO_1037 (O_1037,N_19891,N_19632);
nor UO_1038 (O_1038,N_19627,N_19992);
and UO_1039 (O_1039,N_19790,N_19890);
xor UO_1040 (O_1040,N_19963,N_19868);
or UO_1041 (O_1041,N_19735,N_19961);
nor UO_1042 (O_1042,N_19934,N_19534);
and UO_1043 (O_1043,N_19648,N_19694);
nand UO_1044 (O_1044,N_19573,N_19526);
and UO_1045 (O_1045,N_19927,N_19680);
and UO_1046 (O_1046,N_19809,N_19885);
nor UO_1047 (O_1047,N_19787,N_19577);
or UO_1048 (O_1048,N_19580,N_19667);
or UO_1049 (O_1049,N_19676,N_19823);
nand UO_1050 (O_1050,N_19796,N_19879);
and UO_1051 (O_1051,N_19728,N_19955);
or UO_1052 (O_1052,N_19624,N_19610);
nor UO_1053 (O_1053,N_19733,N_19547);
nand UO_1054 (O_1054,N_19758,N_19827);
nand UO_1055 (O_1055,N_19829,N_19761);
or UO_1056 (O_1056,N_19567,N_19866);
xnor UO_1057 (O_1057,N_19822,N_19859);
nand UO_1058 (O_1058,N_19851,N_19829);
and UO_1059 (O_1059,N_19930,N_19591);
or UO_1060 (O_1060,N_19712,N_19572);
nor UO_1061 (O_1061,N_19866,N_19657);
or UO_1062 (O_1062,N_19872,N_19797);
nor UO_1063 (O_1063,N_19928,N_19623);
nor UO_1064 (O_1064,N_19718,N_19717);
or UO_1065 (O_1065,N_19984,N_19600);
nor UO_1066 (O_1066,N_19612,N_19962);
nand UO_1067 (O_1067,N_19783,N_19963);
xnor UO_1068 (O_1068,N_19671,N_19755);
or UO_1069 (O_1069,N_19684,N_19746);
xor UO_1070 (O_1070,N_19786,N_19903);
nand UO_1071 (O_1071,N_19802,N_19680);
nand UO_1072 (O_1072,N_19767,N_19891);
xor UO_1073 (O_1073,N_19874,N_19606);
nand UO_1074 (O_1074,N_19569,N_19508);
and UO_1075 (O_1075,N_19784,N_19702);
and UO_1076 (O_1076,N_19539,N_19502);
or UO_1077 (O_1077,N_19696,N_19603);
xor UO_1078 (O_1078,N_19517,N_19544);
nand UO_1079 (O_1079,N_19864,N_19932);
xor UO_1080 (O_1080,N_19634,N_19898);
and UO_1081 (O_1081,N_19528,N_19730);
xnor UO_1082 (O_1082,N_19549,N_19942);
or UO_1083 (O_1083,N_19641,N_19557);
xnor UO_1084 (O_1084,N_19552,N_19936);
nor UO_1085 (O_1085,N_19980,N_19907);
or UO_1086 (O_1086,N_19801,N_19502);
xnor UO_1087 (O_1087,N_19968,N_19808);
xnor UO_1088 (O_1088,N_19885,N_19548);
nor UO_1089 (O_1089,N_19774,N_19978);
xnor UO_1090 (O_1090,N_19544,N_19710);
xnor UO_1091 (O_1091,N_19953,N_19584);
xor UO_1092 (O_1092,N_19806,N_19539);
and UO_1093 (O_1093,N_19997,N_19851);
xnor UO_1094 (O_1094,N_19919,N_19983);
xor UO_1095 (O_1095,N_19864,N_19947);
nor UO_1096 (O_1096,N_19815,N_19873);
nor UO_1097 (O_1097,N_19814,N_19998);
or UO_1098 (O_1098,N_19777,N_19828);
and UO_1099 (O_1099,N_19974,N_19774);
nor UO_1100 (O_1100,N_19676,N_19682);
nor UO_1101 (O_1101,N_19728,N_19762);
xor UO_1102 (O_1102,N_19963,N_19836);
or UO_1103 (O_1103,N_19873,N_19790);
or UO_1104 (O_1104,N_19678,N_19866);
or UO_1105 (O_1105,N_19702,N_19600);
and UO_1106 (O_1106,N_19626,N_19917);
or UO_1107 (O_1107,N_19807,N_19969);
xor UO_1108 (O_1108,N_19796,N_19820);
xor UO_1109 (O_1109,N_19700,N_19609);
or UO_1110 (O_1110,N_19573,N_19934);
and UO_1111 (O_1111,N_19757,N_19913);
xnor UO_1112 (O_1112,N_19546,N_19835);
xnor UO_1113 (O_1113,N_19717,N_19723);
nand UO_1114 (O_1114,N_19830,N_19534);
xnor UO_1115 (O_1115,N_19665,N_19792);
nor UO_1116 (O_1116,N_19613,N_19744);
xor UO_1117 (O_1117,N_19597,N_19899);
nor UO_1118 (O_1118,N_19931,N_19603);
nor UO_1119 (O_1119,N_19980,N_19991);
and UO_1120 (O_1120,N_19844,N_19896);
nor UO_1121 (O_1121,N_19771,N_19612);
nor UO_1122 (O_1122,N_19868,N_19951);
and UO_1123 (O_1123,N_19745,N_19767);
or UO_1124 (O_1124,N_19988,N_19691);
or UO_1125 (O_1125,N_19830,N_19733);
or UO_1126 (O_1126,N_19556,N_19988);
xor UO_1127 (O_1127,N_19976,N_19843);
or UO_1128 (O_1128,N_19940,N_19853);
or UO_1129 (O_1129,N_19863,N_19901);
xor UO_1130 (O_1130,N_19893,N_19500);
xnor UO_1131 (O_1131,N_19542,N_19841);
nand UO_1132 (O_1132,N_19511,N_19813);
or UO_1133 (O_1133,N_19785,N_19958);
or UO_1134 (O_1134,N_19976,N_19772);
and UO_1135 (O_1135,N_19728,N_19630);
xor UO_1136 (O_1136,N_19589,N_19534);
nand UO_1137 (O_1137,N_19783,N_19820);
nor UO_1138 (O_1138,N_19995,N_19827);
nand UO_1139 (O_1139,N_19581,N_19817);
or UO_1140 (O_1140,N_19587,N_19542);
xor UO_1141 (O_1141,N_19929,N_19677);
and UO_1142 (O_1142,N_19679,N_19509);
or UO_1143 (O_1143,N_19527,N_19941);
and UO_1144 (O_1144,N_19526,N_19759);
and UO_1145 (O_1145,N_19934,N_19566);
xnor UO_1146 (O_1146,N_19651,N_19688);
or UO_1147 (O_1147,N_19655,N_19781);
nor UO_1148 (O_1148,N_19733,N_19933);
nand UO_1149 (O_1149,N_19736,N_19915);
and UO_1150 (O_1150,N_19591,N_19601);
and UO_1151 (O_1151,N_19502,N_19750);
xnor UO_1152 (O_1152,N_19838,N_19509);
nor UO_1153 (O_1153,N_19648,N_19904);
and UO_1154 (O_1154,N_19558,N_19977);
xor UO_1155 (O_1155,N_19694,N_19587);
and UO_1156 (O_1156,N_19846,N_19849);
nand UO_1157 (O_1157,N_19538,N_19851);
or UO_1158 (O_1158,N_19704,N_19606);
nand UO_1159 (O_1159,N_19905,N_19721);
and UO_1160 (O_1160,N_19634,N_19914);
nand UO_1161 (O_1161,N_19932,N_19559);
or UO_1162 (O_1162,N_19855,N_19879);
and UO_1163 (O_1163,N_19860,N_19971);
nand UO_1164 (O_1164,N_19632,N_19695);
xor UO_1165 (O_1165,N_19981,N_19968);
or UO_1166 (O_1166,N_19544,N_19525);
and UO_1167 (O_1167,N_19831,N_19696);
and UO_1168 (O_1168,N_19924,N_19626);
and UO_1169 (O_1169,N_19589,N_19526);
nand UO_1170 (O_1170,N_19834,N_19566);
xnor UO_1171 (O_1171,N_19839,N_19741);
or UO_1172 (O_1172,N_19812,N_19635);
nand UO_1173 (O_1173,N_19723,N_19729);
and UO_1174 (O_1174,N_19648,N_19891);
or UO_1175 (O_1175,N_19782,N_19722);
and UO_1176 (O_1176,N_19845,N_19592);
nor UO_1177 (O_1177,N_19755,N_19757);
or UO_1178 (O_1178,N_19833,N_19829);
and UO_1179 (O_1179,N_19791,N_19945);
or UO_1180 (O_1180,N_19686,N_19582);
nor UO_1181 (O_1181,N_19589,N_19751);
or UO_1182 (O_1182,N_19547,N_19622);
nor UO_1183 (O_1183,N_19744,N_19772);
xor UO_1184 (O_1184,N_19747,N_19515);
nor UO_1185 (O_1185,N_19511,N_19964);
xor UO_1186 (O_1186,N_19821,N_19559);
nor UO_1187 (O_1187,N_19904,N_19905);
and UO_1188 (O_1188,N_19747,N_19711);
or UO_1189 (O_1189,N_19565,N_19735);
xnor UO_1190 (O_1190,N_19998,N_19845);
or UO_1191 (O_1191,N_19749,N_19595);
and UO_1192 (O_1192,N_19501,N_19849);
nand UO_1193 (O_1193,N_19753,N_19929);
nand UO_1194 (O_1194,N_19583,N_19922);
or UO_1195 (O_1195,N_19931,N_19718);
or UO_1196 (O_1196,N_19654,N_19958);
nor UO_1197 (O_1197,N_19557,N_19728);
xor UO_1198 (O_1198,N_19928,N_19859);
nand UO_1199 (O_1199,N_19920,N_19535);
or UO_1200 (O_1200,N_19803,N_19889);
nand UO_1201 (O_1201,N_19870,N_19751);
xor UO_1202 (O_1202,N_19500,N_19920);
nand UO_1203 (O_1203,N_19652,N_19668);
nor UO_1204 (O_1204,N_19998,N_19579);
nand UO_1205 (O_1205,N_19975,N_19841);
nor UO_1206 (O_1206,N_19874,N_19727);
xnor UO_1207 (O_1207,N_19916,N_19937);
and UO_1208 (O_1208,N_19500,N_19695);
or UO_1209 (O_1209,N_19532,N_19883);
and UO_1210 (O_1210,N_19900,N_19668);
nor UO_1211 (O_1211,N_19591,N_19567);
or UO_1212 (O_1212,N_19849,N_19806);
xor UO_1213 (O_1213,N_19912,N_19917);
nand UO_1214 (O_1214,N_19968,N_19983);
xnor UO_1215 (O_1215,N_19991,N_19829);
xor UO_1216 (O_1216,N_19911,N_19799);
and UO_1217 (O_1217,N_19870,N_19908);
nor UO_1218 (O_1218,N_19526,N_19956);
xnor UO_1219 (O_1219,N_19589,N_19518);
and UO_1220 (O_1220,N_19516,N_19530);
nor UO_1221 (O_1221,N_19602,N_19896);
and UO_1222 (O_1222,N_19912,N_19723);
nand UO_1223 (O_1223,N_19592,N_19974);
and UO_1224 (O_1224,N_19572,N_19747);
and UO_1225 (O_1225,N_19976,N_19685);
xor UO_1226 (O_1226,N_19784,N_19770);
and UO_1227 (O_1227,N_19778,N_19741);
nand UO_1228 (O_1228,N_19514,N_19704);
nand UO_1229 (O_1229,N_19628,N_19823);
xor UO_1230 (O_1230,N_19519,N_19504);
or UO_1231 (O_1231,N_19952,N_19761);
xor UO_1232 (O_1232,N_19555,N_19809);
nor UO_1233 (O_1233,N_19800,N_19920);
and UO_1234 (O_1234,N_19924,N_19565);
nand UO_1235 (O_1235,N_19822,N_19682);
and UO_1236 (O_1236,N_19913,N_19887);
or UO_1237 (O_1237,N_19852,N_19856);
or UO_1238 (O_1238,N_19832,N_19885);
or UO_1239 (O_1239,N_19606,N_19565);
and UO_1240 (O_1240,N_19982,N_19581);
xnor UO_1241 (O_1241,N_19824,N_19622);
or UO_1242 (O_1242,N_19746,N_19532);
nand UO_1243 (O_1243,N_19796,N_19576);
nand UO_1244 (O_1244,N_19555,N_19577);
or UO_1245 (O_1245,N_19844,N_19891);
and UO_1246 (O_1246,N_19788,N_19866);
nand UO_1247 (O_1247,N_19531,N_19622);
or UO_1248 (O_1248,N_19742,N_19634);
nor UO_1249 (O_1249,N_19720,N_19516);
nor UO_1250 (O_1250,N_19605,N_19978);
xor UO_1251 (O_1251,N_19965,N_19836);
or UO_1252 (O_1252,N_19672,N_19908);
and UO_1253 (O_1253,N_19654,N_19879);
nor UO_1254 (O_1254,N_19678,N_19536);
nand UO_1255 (O_1255,N_19797,N_19799);
and UO_1256 (O_1256,N_19687,N_19795);
or UO_1257 (O_1257,N_19656,N_19588);
nor UO_1258 (O_1258,N_19964,N_19982);
nor UO_1259 (O_1259,N_19674,N_19624);
and UO_1260 (O_1260,N_19841,N_19562);
xor UO_1261 (O_1261,N_19971,N_19520);
nor UO_1262 (O_1262,N_19824,N_19937);
nor UO_1263 (O_1263,N_19758,N_19787);
or UO_1264 (O_1264,N_19867,N_19638);
nand UO_1265 (O_1265,N_19996,N_19583);
or UO_1266 (O_1266,N_19868,N_19540);
nor UO_1267 (O_1267,N_19500,N_19586);
and UO_1268 (O_1268,N_19549,N_19624);
nand UO_1269 (O_1269,N_19577,N_19810);
and UO_1270 (O_1270,N_19883,N_19980);
nand UO_1271 (O_1271,N_19877,N_19923);
and UO_1272 (O_1272,N_19529,N_19567);
nor UO_1273 (O_1273,N_19978,N_19519);
nor UO_1274 (O_1274,N_19764,N_19911);
xor UO_1275 (O_1275,N_19525,N_19503);
xnor UO_1276 (O_1276,N_19707,N_19846);
and UO_1277 (O_1277,N_19501,N_19710);
and UO_1278 (O_1278,N_19865,N_19573);
nor UO_1279 (O_1279,N_19653,N_19610);
xnor UO_1280 (O_1280,N_19595,N_19504);
and UO_1281 (O_1281,N_19946,N_19922);
or UO_1282 (O_1282,N_19989,N_19928);
nor UO_1283 (O_1283,N_19975,N_19813);
and UO_1284 (O_1284,N_19858,N_19671);
nand UO_1285 (O_1285,N_19657,N_19760);
or UO_1286 (O_1286,N_19698,N_19523);
or UO_1287 (O_1287,N_19775,N_19709);
xor UO_1288 (O_1288,N_19973,N_19992);
nor UO_1289 (O_1289,N_19959,N_19848);
or UO_1290 (O_1290,N_19750,N_19519);
xor UO_1291 (O_1291,N_19695,N_19640);
and UO_1292 (O_1292,N_19550,N_19569);
or UO_1293 (O_1293,N_19856,N_19882);
and UO_1294 (O_1294,N_19689,N_19539);
nor UO_1295 (O_1295,N_19911,N_19615);
and UO_1296 (O_1296,N_19927,N_19551);
nor UO_1297 (O_1297,N_19675,N_19709);
xnor UO_1298 (O_1298,N_19631,N_19690);
nor UO_1299 (O_1299,N_19949,N_19835);
xor UO_1300 (O_1300,N_19662,N_19822);
xnor UO_1301 (O_1301,N_19510,N_19513);
nand UO_1302 (O_1302,N_19809,N_19920);
nand UO_1303 (O_1303,N_19974,N_19743);
and UO_1304 (O_1304,N_19880,N_19779);
and UO_1305 (O_1305,N_19630,N_19648);
nor UO_1306 (O_1306,N_19586,N_19527);
nand UO_1307 (O_1307,N_19684,N_19619);
or UO_1308 (O_1308,N_19949,N_19958);
nor UO_1309 (O_1309,N_19690,N_19982);
nor UO_1310 (O_1310,N_19538,N_19586);
and UO_1311 (O_1311,N_19749,N_19520);
nor UO_1312 (O_1312,N_19501,N_19907);
and UO_1313 (O_1313,N_19527,N_19580);
xor UO_1314 (O_1314,N_19825,N_19903);
nor UO_1315 (O_1315,N_19935,N_19627);
nand UO_1316 (O_1316,N_19922,N_19990);
nor UO_1317 (O_1317,N_19597,N_19868);
or UO_1318 (O_1318,N_19601,N_19558);
or UO_1319 (O_1319,N_19665,N_19790);
nand UO_1320 (O_1320,N_19589,N_19643);
xnor UO_1321 (O_1321,N_19670,N_19735);
nor UO_1322 (O_1322,N_19908,N_19993);
nor UO_1323 (O_1323,N_19647,N_19616);
nor UO_1324 (O_1324,N_19799,N_19502);
nand UO_1325 (O_1325,N_19982,N_19641);
nor UO_1326 (O_1326,N_19896,N_19867);
and UO_1327 (O_1327,N_19704,N_19568);
nand UO_1328 (O_1328,N_19754,N_19611);
nand UO_1329 (O_1329,N_19860,N_19715);
xnor UO_1330 (O_1330,N_19950,N_19885);
and UO_1331 (O_1331,N_19550,N_19979);
nand UO_1332 (O_1332,N_19571,N_19931);
and UO_1333 (O_1333,N_19688,N_19556);
xnor UO_1334 (O_1334,N_19541,N_19762);
nand UO_1335 (O_1335,N_19559,N_19576);
xnor UO_1336 (O_1336,N_19508,N_19834);
nor UO_1337 (O_1337,N_19619,N_19824);
and UO_1338 (O_1338,N_19531,N_19718);
and UO_1339 (O_1339,N_19810,N_19559);
nor UO_1340 (O_1340,N_19682,N_19601);
or UO_1341 (O_1341,N_19881,N_19625);
xor UO_1342 (O_1342,N_19623,N_19810);
and UO_1343 (O_1343,N_19615,N_19510);
or UO_1344 (O_1344,N_19682,N_19878);
and UO_1345 (O_1345,N_19983,N_19990);
and UO_1346 (O_1346,N_19827,N_19902);
and UO_1347 (O_1347,N_19917,N_19923);
or UO_1348 (O_1348,N_19846,N_19900);
and UO_1349 (O_1349,N_19575,N_19950);
xor UO_1350 (O_1350,N_19824,N_19958);
nor UO_1351 (O_1351,N_19653,N_19629);
nand UO_1352 (O_1352,N_19978,N_19681);
or UO_1353 (O_1353,N_19903,N_19604);
or UO_1354 (O_1354,N_19690,N_19940);
or UO_1355 (O_1355,N_19759,N_19915);
nand UO_1356 (O_1356,N_19703,N_19889);
nand UO_1357 (O_1357,N_19984,N_19965);
nand UO_1358 (O_1358,N_19751,N_19520);
or UO_1359 (O_1359,N_19951,N_19649);
or UO_1360 (O_1360,N_19501,N_19640);
or UO_1361 (O_1361,N_19906,N_19952);
nor UO_1362 (O_1362,N_19788,N_19581);
nor UO_1363 (O_1363,N_19877,N_19994);
nor UO_1364 (O_1364,N_19789,N_19782);
and UO_1365 (O_1365,N_19768,N_19996);
nand UO_1366 (O_1366,N_19960,N_19673);
nor UO_1367 (O_1367,N_19591,N_19987);
or UO_1368 (O_1368,N_19648,N_19552);
and UO_1369 (O_1369,N_19523,N_19702);
nor UO_1370 (O_1370,N_19759,N_19903);
nor UO_1371 (O_1371,N_19778,N_19724);
xor UO_1372 (O_1372,N_19960,N_19808);
nor UO_1373 (O_1373,N_19820,N_19671);
xnor UO_1374 (O_1374,N_19795,N_19869);
or UO_1375 (O_1375,N_19838,N_19843);
nor UO_1376 (O_1376,N_19516,N_19641);
nor UO_1377 (O_1377,N_19786,N_19662);
nand UO_1378 (O_1378,N_19800,N_19729);
nor UO_1379 (O_1379,N_19949,N_19945);
and UO_1380 (O_1380,N_19863,N_19970);
xor UO_1381 (O_1381,N_19556,N_19852);
nand UO_1382 (O_1382,N_19988,N_19827);
xor UO_1383 (O_1383,N_19972,N_19965);
nand UO_1384 (O_1384,N_19716,N_19661);
nand UO_1385 (O_1385,N_19635,N_19575);
or UO_1386 (O_1386,N_19505,N_19968);
or UO_1387 (O_1387,N_19925,N_19565);
and UO_1388 (O_1388,N_19549,N_19933);
and UO_1389 (O_1389,N_19974,N_19954);
or UO_1390 (O_1390,N_19960,N_19874);
and UO_1391 (O_1391,N_19674,N_19548);
nand UO_1392 (O_1392,N_19816,N_19683);
xor UO_1393 (O_1393,N_19568,N_19501);
and UO_1394 (O_1394,N_19583,N_19888);
and UO_1395 (O_1395,N_19835,N_19607);
xor UO_1396 (O_1396,N_19793,N_19962);
and UO_1397 (O_1397,N_19656,N_19712);
xnor UO_1398 (O_1398,N_19695,N_19736);
xor UO_1399 (O_1399,N_19879,N_19736);
nand UO_1400 (O_1400,N_19887,N_19557);
or UO_1401 (O_1401,N_19871,N_19811);
or UO_1402 (O_1402,N_19905,N_19574);
nand UO_1403 (O_1403,N_19868,N_19709);
xnor UO_1404 (O_1404,N_19987,N_19662);
and UO_1405 (O_1405,N_19940,N_19952);
and UO_1406 (O_1406,N_19504,N_19919);
and UO_1407 (O_1407,N_19893,N_19655);
or UO_1408 (O_1408,N_19689,N_19935);
or UO_1409 (O_1409,N_19505,N_19780);
nand UO_1410 (O_1410,N_19690,N_19934);
and UO_1411 (O_1411,N_19916,N_19757);
xor UO_1412 (O_1412,N_19567,N_19978);
or UO_1413 (O_1413,N_19773,N_19890);
nand UO_1414 (O_1414,N_19767,N_19792);
xnor UO_1415 (O_1415,N_19815,N_19697);
or UO_1416 (O_1416,N_19586,N_19996);
nor UO_1417 (O_1417,N_19723,N_19772);
and UO_1418 (O_1418,N_19954,N_19928);
nor UO_1419 (O_1419,N_19812,N_19914);
nand UO_1420 (O_1420,N_19665,N_19855);
nand UO_1421 (O_1421,N_19797,N_19753);
nor UO_1422 (O_1422,N_19913,N_19672);
and UO_1423 (O_1423,N_19605,N_19504);
nor UO_1424 (O_1424,N_19505,N_19989);
or UO_1425 (O_1425,N_19766,N_19707);
and UO_1426 (O_1426,N_19884,N_19567);
nor UO_1427 (O_1427,N_19788,N_19980);
nor UO_1428 (O_1428,N_19994,N_19648);
and UO_1429 (O_1429,N_19646,N_19825);
or UO_1430 (O_1430,N_19719,N_19753);
xnor UO_1431 (O_1431,N_19620,N_19982);
and UO_1432 (O_1432,N_19830,N_19660);
xnor UO_1433 (O_1433,N_19785,N_19730);
nor UO_1434 (O_1434,N_19661,N_19664);
or UO_1435 (O_1435,N_19680,N_19595);
or UO_1436 (O_1436,N_19781,N_19876);
xnor UO_1437 (O_1437,N_19600,N_19725);
and UO_1438 (O_1438,N_19988,N_19815);
nand UO_1439 (O_1439,N_19857,N_19871);
and UO_1440 (O_1440,N_19571,N_19952);
and UO_1441 (O_1441,N_19802,N_19765);
nor UO_1442 (O_1442,N_19875,N_19931);
or UO_1443 (O_1443,N_19674,N_19630);
nor UO_1444 (O_1444,N_19980,N_19525);
or UO_1445 (O_1445,N_19832,N_19660);
nand UO_1446 (O_1446,N_19964,N_19764);
or UO_1447 (O_1447,N_19882,N_19646);
nand UO_1448 (O_1448,N_19592,N_19756);
nor UO_1449 (O_1449,N_19706,N_19766);
and UO_1450 (O_1450,N_19574,N_19650);
and UO_1451 (O_1451,N_19995,N_19885);
and UO_1452 (O_1452,N_19887,N_19508);
xor UO_1453 (O_1453,N_19567,N_19708);
nor UO_1454 (O_1454,N_19990,N_19679);
or UO_1455 (O_1455,N_19735,N_19892);
and UO_1456 (O_1456,N_19751,N_19897);
nand UO_1457 (O_1457,N_19818,N_19655);
or UO_1458 (O_1458,N_19599,N_19997);
xnor UO_1459 (O_1459,N_19536,N_19900);
xnor UO_1460 (O_1460,N_19940,N_19631);
nor UO_1461 (O_1461,N_19710,N_19532);
and UO_1462 (O_1462,N_19977,N_19503);
nor UO_1463 (O_1463,N_19732,N_19607);
nand UO_1464 (O_1464,N_19853,N_19666);
nor UO_1465 (O_1465,N_19629,N_19591);
nor UO_1466 (O_1466,N_19923,N_19777);
or UO_1467 (O_1467,N_19885,N_19561);
nand UO_1468 (O_1468,N_19861,N_19723);
nor UO_1469 (O_1469,N_19757,N_19978);
or UO_1470 (O_1470,N_19559,N_19714);
or UO_1471 (O_1471,N_19602,N_19752);
nor UO_1472 (O_1472,N_19778,N_19949);
or UO_1473 (O_1473,N_19852,N_19818);
xnor UO_1474 (O_1474,N_19643,N_19966);
nand UO_1475 (O_1475,N_19965,N_19842);
and UO_1476 (O_1476,N_19746,N_19519);
or UO_1477 (O_1477,N_19528,N_19724);
nor UO_1478 (O_1478,N_19988,N_19714);
nand UO_1479 (O_1479,N_19728,N_19517);
or UO_1480 (O_1480,N_19628,N_19629);
and UO_1481 (O_1481,N_19597,N_19540);
nand UO_1482 (O_1482,N_19920,N_19798);
nor UO_1483 (O_1483,N_19528,N_19978);
xor UO_1484 (O_1484,N_19791,N_19910);
nand UO_1485 (O_1485,N_19670,N_19974);
or UO_1486 (O_1486,N_19562,N_19612);
nand UO_1487 (O_1487,N_19962,N_19772);
or UO_1488 (O_1488,N_19882,N_19584);
or UO_1489 (O_1489,N_19819,N_19915);
and UO_1490 (O_1490,N_19656,N_19807);
or UO_1491 (O_1491,N_19715,N_19893);
nand UO_1492 (O_1492,N_19644,N_19957);
or UO_1493 (O_1493,N_19999,N_19661);
and UO_1494 (O_1494,N_19971,N_19527);
or UO_1495 (O_1495,N_19650,N_19623);
nand UO_1496 (O_1496,N_19644,N_19782);
nand UO_1497 (O_1497,N_19619,N_19557);
or UO_1498 (O_1498,N_19822,N_19899);
xnor UO_1499 (O_1499,N_19734,N_19578);
nand UO_1500 (O_1500,N_19711,N_19572);
nor UO_1501 (O_1501,N_19548,N_19599);
xnor UO_1502 (O_1502,N_19717,N_19607);
and UO_1503 (O_1503,N_19727,N_19562);
xnor UO_1504 (O_1504,N_19561,N_19810);
xnor UO_1505 (O_1505,N_19653,N_19534);
nor UO_1506 (O_1506,N_19846,N_19928);
xor UO_1507 (O_1507,N_19789,N_19623);
nand UO_1508 (O_1508,N_19751,N_19706);
nor UO_1509 (O_1509,N_19896,N_19833);
nand UO_1510 (O_1510,N_19997,N_19781);
or UO_1511 (O_1511,N_19734,N_19672);
and UO_1512 (O_1512,N_19678,N_19683);
or UO_1513 (O_1513,N_19537,N_19931);
xor UO_1514 (O_1514,N_19968,N_19694);
and UO_1515 (O_1515,N_19683,N_19509);
xnor UO_1516 (O_1516,N_19573,N_19938);
and UO_1517 (O_1517,N_19941,N_19740);
nand UO_1518 (O_1518,N_19834,N_19594);
nand UO_1519 (O_1519,N_19986,N_19703);
and UO_1520 (O_1520,N_19757,N_19577);
nand UO_1521 (O_1521,N_19732,N_19770);
or UO_1522 (O_1522,N_19613,N_19696);
nand UO_1523 (O_1523,N_19529,N_19980);
nor UO_1524 (O_1524,N_19610,N_19862);
or UO_1525 (O_1525,N_19704,N_19733);
nand UO_1526 (O_1526,N_19552,N_19964);
xnor UO_1527 (O_1527,N_19532,N_19774);
or UO_1528 (O_1528,N_19749,N_19647);
nand UO_1529 (O_1529,N_19668,N_19511);
nor UO_1530 (O_1530,N_19608,N_19507);
or UO_1531 (O_1531,N_19910,N_19892);
or UO_1532 (O_1532,N_19943,N_19621);
and UO_1533 (O_1533,N_19547,N_19667);
and UO_1534 (O_1534,N_19592,N_19897);
and UO_1535 (O_1535,N_19947,N_19912);
or UO_1536 (O_1536,N_19878,N_19542);
xnor UO_1537 (O_1537,N_19900,N_19908);
xnor UO_1538 (O_1538,N_19665,N_19656);
xor UO_1539 (O_1539,N_19853,N_19874);
nand UO_1540 (O_1540,N_19679,N_19783);
xnor UO_1541 (O_1541,N_19655,N_19751);
and UO_1542 (O_1542,N_19997,N_19962);
or UO_1543 (O_1543,N_19800,N_19642);
nand UO_1544 (O_1544,N_19639,N_19653);
nand UO_1545 (O_1545,N_19549,N_19901);
nand UO_1546 (O_1546,N_19661,N_19752);
nand UO_1547 (O_1547,N_19809,N_19765);
nand UO_1548 (O_1548,N_19701,N_19686);
and UO_1549 (O_1549,N_19858,N_19898);
or UO_1550 (O_1550,N_19547,N_19952);
nor UO_1551 (O_1551,N_19680,N_19711);
nand UO_1552 (O_1552,N_19661,N_19970);
nor UO_1553 (O_1553,N_19868,N_19565);
and UO_1554 (O_1554,N_19568,N_19539);
and UO_1555 (O_1555,N_19504,N_19500);
xor UO_1556 (O_1556,N_19693,N_19675);
nand UO_1557 (O_1557,N_19523,N_19612);
nor UO_1558 (O_1558,N_19558,N_19695);
nor UO_1559 (O_1559,N_19958,N_19575);
and UO_1560 (O_1560,N_19546,N_19755);
nand UO_1561 (O_1561,N_19943,N_19682);
or UO_1562 (O_1562,N_19993,N_19717);
and UO_1563 (O_1563,N_19546,N_19820);
xnor UO_1564 (O_1564,N_19753,N_19739);
nand UO_1565 (O_1565,N_19671,N_19750);
nor UO_1566 (O_1566,N_19691,N_19707);
and UO_1567 (O_1567,N_19614,N_19587);
nor UO_1568 (O_1568,N_19508,N_19974);
nor UO_1569 (O_1569,N_19813,N_19718);
nand UO_1570 (O_1570,N_19749,N_19785);
nand UO_1571 (O_1571,N_19940,N_19957);
nor UO_1572 (O_1572,N_19863,N_19602);
nor UO_1573 (O_1573,N_19713,N_19904);
or UO_1574 (O_1574,N_19806,N_19863);
and UO_1575 (O_1575,N_19977,N_19627);
xnor UO_1576 (O_1576,N_19999,N_19898);
xor UO_1577 (O_1577,N_19956,N_19788);
nand UO_1578 (O_1578,N_19924,N_19882);
nor UO_1579 (O_1579,N_19954,N_19588);
nand UO_1580 (O_1580,N_19580,N_19815);
and UO_1581 (O_1581,N_19584,N_19877);
nand UO_1582 (O_1582,N_19897,N_19545);
nor UO_1583 (O_1583,N_19623,N_19841);
xor UO_1584 (O_1584,N_19611,N_19945);
xor UO_1585 (O_1585,N_19605,N_19773);
or UO_1586 (O_1586,N_19575,N_19698);
or UO_1587 (O_1587,N_19791,N_19868);
xor UO_1588 (O_1588,N_19576,N_19911);
and UO_1589 (O_1589,N_19914,N_19940);
and UO_1590 (O_1590,N_19949,N_19550);
and UO_1591 (O_1591,N_19564,N_19861);
xor UO_1592 (O_1592,N_19976,N_19946);
nor UO_1593 (O_1593,N_19760,N_19849);
and UO_1594 (O_1594,N_19986,N_19536);
and UO_1595 (O_1595,N_19914,N_19865);
xnor UO_1596 (O_1596,N_19895,N_19683);
xor UO_1597 (O_1597,N_19642,N_19713);
or UO_1598 (O_1598,N_19608,N_19877);
nor UO_1599 (O_1599,N_19628,N_19555);
xor UO_1600 (O_1600,N_19817,N_19555);
and UO_1601 (O_1601,N_19903,N_19670);
nor UO_1602 (O_1602,N_19509,N_19966);
xnor UO_1603 (O_1603,N_19925,N_19921);
nand UO_1604 (O_1604,N_19538,N_19909);
and UO_1605 (O_1605,N_19602,N_19751);
nand UO_1606 (O_1606,N_19613,N_19730);
and UO_1607 (O_1607,N_19592,N_19738);
xnor UO_1608 (O_1608,N_19748,N_19671);
and UO_1609 (O_1609,N_19576,N_19625);
xor UO_1610 (O_1610,N_19591,N_19798);
xnor UO_1611 (O_1611,N_19879,N_19964);
and UO_1612 (O_1612,N_19527,N_19733);
or UO_1613 (O_1613,N_19538,N_19526);
and UO_1614 (O_1614,N_19914,N_19697);
nand UO_1615 (O_1615,N_19779,N_19819);
nor UO_1616 (O_1616,N_19508,N_19976);
nor UO_1617 (O_1617,N_19814,N_19915);
xor UO_1618 (O_1618,N_19615,N_19870);
xor UO_1619 (O_1619,N_19790,N_19885);
and UO_1620 (O_1620,N_19974,N_19831);
nand UO_1621 (O_1621,N_19759,N_19679);
and UO_1622 (O_1622,N_19574,N_19957);
nor UO_1623 (O_1623,N_19727,N_19696);
nand UO_1624 (O_1624,N_19845,N_19782);
xor UO_1625 (O_1625,N_19815,N_19937);
nor UO_1626 (O_1626,N_19698,N_19926);
xnor UO_1627 (O_1627,N_19839,N_19705);
nand UO_1628 (O_1628,N_19515,N_19545);
nand UO_1629 (O_1629,N_19704,N_19586);
nor UO_1630 (O_1630,N_19646,N_19922);
nor UO_1631 (O_1631,N_19955,N_19766);
xnor UO_1632 (O_1632,N_19718,N_19631);
or UO_1633 (O_1633,N_19967,N_19611);
or UO_1634 (O_1634,N_19744,N_19526);
nand UO_1635 (O_1635,N_19505,N_19651);
nand UO_1636 (O_1636,N_19940,N_19672);
nor UO_1637 (O_1637,N_19708,N_19576);
and UO_1638 (O_1638,N_19661,N_19899);
nor UO_1639 (O_1639,N_19588,N_19679);
nor UO_1640 (O_1640,N_19628,N_19689);
nor UO_1641 (O_1641,N_19898,N_19721);
and UO_1642 (O_1642,N_19556,N_19555);
nor UO_1643 (O_1643,N_19737,N_19703);
nor UO_1644 (O_1644,N_19928,N_19647);
nand UO_1645 (O_1645,N_19510,N_19842);
and UO_1646 (O_1646,N_19540,N_19891);
xnor UO_1647 (O_1647,N_19751,N_19906);
nand UO_1648 (O_1648,N_19687,N_19863);
or UO_1649 (O_1649,N_19540,N_19548);
and UO_1650 (O_1650,N_19935,N_19968);
nand UO_1651 (O_1651,N_19952,N_19861);
and UO_1652 (O_1652,N_19576,N_19951);
and UO_1653 (O_1653,N_19785,N_19760);
nand UO_1654 (O_1654,N_19504,N_19798);
nand UO_1655 (O_1655,N_19508,N_19632);
or UO_1656 (O_1656,N_19683,N_19784);
or UO_1657 (O_1657,N_19756,N_19874);
or UO_1658 (O_1658,N_19811,N_19652);
or UO_1659 (O_1659,N_19841,N_19749);
nand UO_1660 (O_1660,N_19897,N_19565);
and UO_1661 (O_1661,N_19938,N_19578);
xnor UO_1662 (O_1662,N_19966,N_19647);
nand UO_1663 (O_1663,N_19932,N_19906);
nand UO_1664 (O_1664,N_19775,N_19716);
nand UO_1665 (O_1665,N_19950,N_19972);
nor UO_1666 (O_1666,N_19917,N_19532);
nand UO_1667 (O_1667,N_19801,N_19531);
nand UO_1668 (O_1668,N_19528,N_19987);
xnor UO_1669 (O_1669,N_19999,N_19876);
nor UO_1670 (O_1670,N_19887,N_19732);
or UO_1671 (O_1671,N_19762,N_19507);
and UO_1672 (O_1672,N_19555,N_19580);
nand UO_1673 (O_1673,N_19598,N_19731);
nor UO_1674 (O_1674,N_19878,N_19726);
nor UO_1675 (O_1675,N_19645,N_19787);
xor UO_1676 (O_1676,N_19735,N_19757);
nor UO_1677 (O_1677,N_19804,N_19589);
nor UO_1678 (O_1678,N_19879,N_19902);
or UO_1679 (O_1679,N_19669,N_19932);
nor UO_1680 (O_1680,N_19615,N_19517);
and UO_1681 (O_1681,N_19619,N_19972);
or UO_1682 (O_1682,N_19846,N_19711);
and UO_1683 (O_1683,N_19614,N_19761);
or UO_1684 (O_1684,N_19678,N_19798);
and UO_1685 (O_1685,N_19895,N_19768);
xnor UO_1686 (O_1686,N_19659,N_19956);
nand UO_1687 (O_1687,N_19661,N_19715);
and UO_1688 (O_1688,N_19532,N_19586);
nand UO_1689 (O_1689,N_19653,N_19929);
xor UO_1690 (O_1690,N_19739,N_19686);
nor UO_1691 (O_1691,N_19855,N_19773);
and UO_1692 (O_1692,N_19729,N_19924);
or UO_1693 (O_1693,N_19987,N_19541);
xnor UO_1694 (O_1694,N_19798,N_19709);
nand UO_1695 (O_1695,N_19590,N_19582);
or UO_1696 (O_1696,N_19795,N_19663);
or UO_1697 (O_1697,N_19624,N_19964);
nand UO_1698 (O_1698,N_19861,N_19995);
nand UO_1699 (O_1699,N_19623,N_19959);
or UO_1700 (O_1700,N_19984,N_19671);
nor UO_1701 (O_1701,N_19763,N_19753);
xor UO_1702 (O_1702,N_19617,N_19903);
and UO_1703 (O_1703,N_19838,N_19535);
xnor UO_1704 (O_1704,N_19760,N_19754);
xnor UO_1705 (O_1705,N_19798,N_19987);
and UO_1706 (O_1706,N_19775,N_19907);
nand UO_1707 (O_1707,N_19837,N_19558);
xnor UO_1708 (O_1708,N_19566,N_19868);
or UO_1709 (O_1709,N_19540,N_19704);
xnor UO_1710 (O_1710,N_19797,N_19813);
or UO_1711 (O_1711,N_19831,N_19802);
and UO_1712 (O_1712,N_19618,N_19561);
and UO_1713 (O_1713,N_19701,N_19561);
or UO_1714 (O_1714,N_19882,N_19691);
nand UO_1715 (O_1715,N_19754,N_19515);
nor UO_1716 (O_1716,N_19934,N_19984);
or UO_1717 (O_1717,N_19693,N_19726);
nor UO_1718 (O_1718,N_19783,N_19975);
or UO_1719 (O_1719,N_19647,N_19972);
xor UO_1720 (O_1720,N_19610,N_19705);
and UO_1721 (O_1721,N_19757,N_19504);
and UO_1722 (O_1722,N_19896,N_19566);
and UO_1723 (O_1723,N_19595,N_19788);
nor UO_1724 (O_1724,N_19952,N_19680);
nor UO_1725 (O_1725,N_19811,N_19683);
and UO_1726 (O_1726,N_19646,N_19644);
xnor UO_1727 (O_1727,N_19545,N_19530);
and UO_1728 (O_1728,N_19735,N_19978);
or UO_1729 (O_1729,N_19733,N_19592);
or UO_1730 (O_1730,N_19536,N_19640);
xnor UO_1731 (O_1731,N_19853,N_19768);
or UO_1732 (O_1732,N_19731,N_19670);
or UO_1733 (O_1733,N_19737,N_19604);
nor UO_1734 (O_1734,N_19666,N_19647);
nand UO_1735 (O_1735,N_19845,N_19746);
nor UO_1736 (O_1736,N_19898,N_19856);
nand UO_1737 (O_1737,N_19945,N_19909);
nor UO_1738 (O_1738,N_19760,N_19627);
or UO_1739 (O_1739,N_19611,N_19607);
nand UO_1740 (O_1740,N_19723,N_19982);
nand UO_1741 (O_1741,N_19818,N_19617);
nand UO_1742 (O_1742,N_19988,N_19929);
nor UO_1743 (O_1743,N_19533,N_19747);
nand UO_1744 (O_1744,N_19923,N_19981);
and UO_1745 (O_1745,N_19611,N_19928);
nand UO_1746 (O_1746,N_19549,N_19699);
nand UO_1747 (O_1747,N_19799,N_19967);
xor UO_1748 (O_1748,N_19841,N_19538);
nor UO_1749 (O_1749,N_19740,N_19674);
xor UO_1750 (O_1750,N_19612,N_19936);
or UO_1751 (O_1751,N_19537,N_19707);
xnor UO_1752 (O_1752,N_19873,N_19782);
and UO_1753 (O_1753,N_19808,N_19736);
nor UO_1754 (O_1754,N_19930,N_19588);
nor UO_1755 (O_1755,N_19695,N_19560);
nor UO_1756 (O_1756,N_19827,N_19617);
nor UO_1757 (O_1757,N_19519,N_19861);
xnor UO_1758 (O_1758,N_19934,N_19609);
nor UO_1759 (O_1759,N_19528,N_19788);
and UO_1760 (O_1760,N_19759,N_19625);
or UO_1761 (O_1761,N_19925,N_19751);
or UO_1762 (O_1762,N_19754,N_19726);
xor UO_1763 (O_1763,N_19923,N_19862);
or UO_1764 (O_1764,N_19758,N_19544);
nand UO_1765 (O_1765,N_19816,N_19895);
nor UO_1766 (O_1766,N_19888,N_19849);
and UO_1767 (O_1767,N_19784,N_19863);
and UO_1768 (O_1768,N_19726,N_19925);
and UO_1769 (O_1769,N_19515,N_19840);
xor UO_1770 (O_1770,N_19938,N_19545);
nor UO_1771 (O_1771,N_19864,N_19670);
xnor UO_1772 (O_1772,N_19681,N_19952);
nand UO_1773 (O_1773,N_19985,N_19741);
xnor UO_1774 (O_1774,N_19864,N_19739);
nand UO_1775 (O_1775,N_19935,N_19879);
xnor UO_1776 (O_1776,N_19892,N_19818);
xnor UO_1777 (O_1777,N_19642,N_19979);
or UO_1778 (O_1778,N_19620,N_19822);
xnor UO_1779 (O_1779,N_19549,N_19580);
and UO_1780 (O_1780,N_19542,N_19896);
or UO_1781 (O_1781,N_19707,N_19695);
xnor UO_1782 (O_1782,N_19686,N_19859);
and UO_1783 (O_1783,N_19848,N_19768);
nand UO_1784 (O_1784,N_19814,N_19943);
nand UO_1785 (O_1785,N_19502,N_19866);
nor UO_1786 (O_1786,N_19628,N_19751);
xor UO_1787 (O_1787,N_19916,N_19560);
and UO_1788 (O_1788,N_19825,N_19576);
nor UO_1789 (O_1789,N_19835,N_19686);
or UO_1790 (O_1790,N_19571,N_19936);
and UO_1791 (O_1791,N_19541,N_19597);
or UO_1792 (O_1792,N_19869,N_19620);
nor UO_1793 (O_1793,N_19867,N_19918);
or UO_1794 (O_1794,N_19880,N_19635);
or UO_1795 (O_1795,N_19934,N_19986);
xor UO_1796 (O_1796,N_19970,N_19513);
nor UO_1797 (O_1797,N_19896,N_19752);
xor UO_1798 (O_1798,N_19929,N_19520);
xnor UO_1799 (O_1799,N_19717,N_19804);
or UO_1800 (O_1800,N_19861,N_19898);
or UO_1801 (O_1801,N_19572,N_19610);
and UO_1802 (O_1802,N_19758,N_19775);
nand UO_1803 (O_1803,N_19534,N_19743);
xor UO_1804 (O_1804,N_19538,N_19726);
xor UO_1805 (O_1805,N_19872,N_19673);
and UO_1806 (O_1806,N_19861,N_19891);
xor UO_1807 (O_1807,N_19693,N_19642);
nand UO_1808 (O_1808,N_19735,N_19538);
or UO_1809 (O_1809,N_19982,N_19745);
or UO_1810 (O_1810,N_19788,N_19759);
or UO_1811 (O_1811,N_19899,N_19515);
xnor UO_1812 (O_1812,N_19533,N_19526);
xnor UO_1813 (O_1813,N_19516,N_19735);
or UO_1814 (O_1814,N_19577,N_19966);
nand UO_1815 (O_1815,N_19702,N_19817);
nand UO_1816 (O_1816,N_19547,N_19865);
nand UO_1817 (O_1817,N_19751,N_19726);
or UO_1818 (O_1818,N_19839,N_19649);
or UO_1819 (O_1819,N_19802,N_19707);
and UO_1820 (O_1820,N_19873,N_19690);
xnor UO_1821 (O_1821,N_19809,N_19808);
nand UO_1822 (O_1822,N_19620,N_19594);
nand UO_1823 (O_1823,N_19608,N_19741);
nand UO_1824 (O_1824,N_19656,N_19559);
or UO_1825 (O_1825,N_19783,N_19921);
nor UO_1826 (O_1826,N_19796,N_19917);
nor UO_1827 (O_1827,N_19546,N_19898);
nand UO_1828 (O_1828,N_19851,N_19802);
and UO_1829 (O_1829,N_19611,N_19575);
nand UO_1830 (O_1830,N_19938,N_19993);
and UO_1831 (O_1831,N_19640,N_19626);
and UO_1832 (O_1832,N_19939,N_19730);
or UO_1833 (O_1833,N_19711,N_19718);
xnor UO_1834 (O_1834,N_19651,N_19776);
nor UO_1835 (O_1835,N_19544,N_19609);
xor UO_1836 (O_1836,N_19956,N_19803);
nor UO_1837 (O_1837,N_19806,N_19727);
nand UO_1838 (O_1838,N_19933,N_19863);
or UO_1839 (O_1839,N_19696,N_19943);
nor UO_1840 (O_1840,N_19726,N_19845);
xnor UO_1841 (O_1841,N_19731,N_19898);
nor UO_1842 (O_1842,N_19648,N_19966);
and UO_1843 (O_1843,N_19532,N_19699);
and UO_1844 (O_1844,N_19819,N_19548);
nand UO_1845 (O_1845,N_19500,N_19708);
or UO_1846 (O_1846,N_19849,N_19664);
and UO_1847 (O_1847,N_19796,N_19809);
or UO_1848 (O_1848,N_19500,N_19646);
xor UO_1849 (O_1849,N_19580,N_19503);
and UO_1850 (O_1850,N_19899,N_19954);
xor UO_1851 (O_1851,N_19522,N_19631);
nor UO_1852 (O_1852,N_19767,N_19712);
or UO_1853 (O_1853,N_19958,N_19930);
and UO_1854 (O_1854,N_19791,N_19727);
xnor UO_1855 (O_1855,N_19971,N_19705);
and UO_1856 (O_1856,N_19676,N_19582);
and UO_1857 (O_1857,N_19694,N_19789);
nor UO_1858 (O_1858,N_19802,N_19848);
nand UO_1859 (O_1859,N_19660,N_19657);
nand UO_1860 (O_1860,N_19578,N_19793);
xor UO_1861 (O_1861,N_19848,N_19747);
xnor UO_1862 (O_1862,N_19967,N_19797);
and UO_1863 (O_1863,N_19892,N_19718);
xnor UO_1864 (O_1864,N_19897,N_19691);
or UO_1865 (O_1865,N_19903,N_19896);
nand UO_1866 (O_1866,N_19859,N_19535);
xor UO_1867 (O_1867,N_19865,N_19501);
nor UO_1868 (O_1868,N_19915,N_19563);
nor UO_1869 (O_1869,N_19757,N_19512);
and UO_1870 (O_1870,N_19812,N_19837);
xnor UO_1871 (O_1871,N_19694,N_19528);
nor UO_1872 (O_1872,N_19825,N_19855);
nand UO_1873 (O_1873,N_19662,N_19926);
nand UO_1874 (O_1874,N_19594,N_19995);
nor UO_1875 (O_1875,N_19780,N_19676);
nand UO_1876 (O_1876,N_19819,N_19984);
nand UO_1877 (O_1877,N_19535,N_19700);
xnor UO_1878 (O_1878,N_19588,N_19593);
xnor UO_1879 (O_1879,N_19598,N_19515);
and UO_1880 (O_1880,N_19580,N_19926);
xnor UO_1881 (O_1881,N_19720,N_19781);
xor UO_1882 (O_1882,N_19754,N_19604);
and UO_1883 (O_1883,N_19782,N_19710);
nor UO_1884 (O_1884,N_19925,N_19688);
nand UO_1885 (O_1885,N_19978,N_19859);
and UO_1886 (O_1886,N_19767,N_19556);
xor UO_1887 (O_1887,N_19673,N_19603);
or UO_1888 (O_1888,N_19702,N_19573);
xor UO_1889 (O_1889,N_19662,N_19883);
and UO_1890 (O_1890,N_19553,N_19560);
xnor UO_1891 (O_1891,N_19845,N_19671);
or UO_1892 (O_1892,N_19608,N_19535);
nand UO_1893 (O_1893,N_19602,N_19960);
xor UO_1894 (O_1894,N_19770,N_19503);
xor UO_1895 (O_1895,N_19987,N_19795);
and UO_1896 (O_1896,N_19900,N_19847);
or UO_1897 (O_1897,N_19978,N_19871);
or UO_1898 (O_1898,N_19809,N_19595);
nand UO_1899 (O_1899,N_19662,N_19941);
and UO_1900 (O_1900,N_19916,N_19511);
xor UO_1901 (O_1901,N_19912,N_19669);
xnor UO_1902 (O_1902,N_19828,N_19906);
nor UO_1903 (O_1903,N_19552,N_19848);
nand UO_1904 (O_1904,N_19633,N_19609);
and UO_1905 (O_1905,N_19660,N_19623);
or UO_1906 (O_1906,N_19908,N_19619);
nand UO_1907 (O_1907,N_19580,N_19653);
nor UO_1908 (O_1908,N_19806,N_19703);
nand UO_1909 (O_1909,N_19786,N_19845);
and UO_1910 (O_1910,N_19814,N_19847);
or UO_1911 (O_1911,N_19570,N_19794);
or UO_1912 (O_1912,N_19965,N_19542);
and UO_1913 (O_1913,N_19941,N_19687);
and UO_1914 (O_1914,N_19924,N_19658);
and UO_1915 (O_1915,N_19634,N_19799);
nor UO_1916 (O_1916,N_19710,N_19682);
nand UO_1917 (O_1917,N_19678,N_19827);
and UO_1918 (O_1918,N_19514,N_19661);
nor UO_1919 (O_1919,N_19829,N_19953);
nand UO_1920 (O_1920,N_19950,N_19999);
nor UO_1921 (O_1921,N_19813,N_19784);
or UO_1922 (O_1922,N_19579,N_19827);
or UO_1923 (O_1923,N_19919,N_19685);
or UO_1924 (O_1924,N_19851,N_19749);
or UO_1925 (O_1925,N_19610,N_19889);
nor UO_1926 (O_1926,N_19898,N_19901);
xor UO_1927 (O_1927,N_19767,N_19946);
nand UO_1928 (O_1928,N_19817,N_19568);
or UO_1929 (O_1929,N_19772,N_19639);
or UO_1930 (O_1930,N_19827,N_19938);
nor UO_1931 (O_1931,N_19944,N_19858);
nor UO_1932 (O_1932,N_19542,N_19977);
nand UO_1933 (O_1933,N_19857,N_19715);
or UO_1934 (O_1934,N_19761,N_19776);
xor UO_1935 (O_1935,N_19763,N_19677);
nand UO_1936 (O_1936,N_19689,N_19714);
xor UO_1937 (O_1937,N_19987,N_19974);
nand UO_1938 (O_1938,N_19718,N_19609);
nand UO_1939 (O_1939,N_19818,N_19709);
nor UO_1940 (O_1940,N_19907,N_19868);
nand UO_1941 (O_1941,N_19866,N_19544);
nor UO_1942 (O_1942,N_19911,N_19510);
nand UO_1943 (O_1943,N_19617,N_19804);
nand UO_1944 (O_1944,N_19900,N_19860);
nor UO_1945 (O_1945,N_19602,N_19658);
xnor UO_1946 (O_1946,N_19513,N_19889);
nand UO_1947 (O_1947,N_19580,N_19863);
xnor UO_1948 (O_1948,N_19970,N_19550);
xor UO_1949 (O_1949,N_19976,N_19835);
xor UO_1950 (O_1950,N_19880,N_19828);
xnor UO_1951 (O_1951,N_19516,N_19847);
or UO_1952 (O_1952,N_19634,N_19921);
nand UO_1953 (O_1953,N_19928,N_19984);
nand UO_1954 (O_1954,N_19888,N_19829);
nand UO_1955 (O_1955,N_19740,N_19664);
nand UO_1956 (O_1956,N_19993,N_19996);
nand UO_1957 (O_1957,N_19807,N_19594);
nor UO_1958 (O_1958,N_19816,N_19690);
and UO_1959 (O_1959,N_19930,N_19518);
xor UO_1960 (O_1960,N_19736,N_19673);
xor UO_1961 (O_1961,N_19565,N_19853);
or UO_1962 (O_1962,N_19941,N_19869);
nand UO_1963 (O_1963,N_19859,N_19667);
or UO_1964 (O_1964,N_19660,N_19600);
nor UO_1965 (O_1965,N_19606,N_19522);
nor UO_1966 (O_1966,N_19537,N_19902);
nor UO_1967 (O_1967,N_19606,N_19946);
nor UO_1968 (O_1968,N_19683,N_19909);
xor UO_1969 (O_1969,N_19574,N_19701);
nand UO_1970 (O_1970,N_19987,N_19647);
nand UO_1971 (O_1971,N_19669,N_19588);
nor UO_1972 (O_1972,N_19730,N_19801);
nand UO_1973 (O_1973,N_19805,N_19640);
or UO_1974 (O_1974,N_19958,N_19540);
or UO_1975 (O_1975,N_19985,N_19849);
or UO_1976 (O_1976,N_19936,N_19718);
or UO_1977 (O_1977,N_19809,N_19981);
nor UO_1978 (O_1978,N_19512,N_19869);
nor UO_1979 (O_1979,N_19879,N_19647);
or UO_1980 (O_1980,N_19930,N_19819);
or UO_1981 (O_1981,N_19801,N_19771);
nor UO_1982 (O_1982,N_19683,N_19556);
nand UO_1983 (O_1983,N_19912,N_19632);
nor UO_1984 (O_1984,N_19695,N_19685);
or UO_1985 (O_1985,N_19847,N_19985);
xor UO_1986 (O_1986,N_19861,N_19578);
and UO_1987 (O_1987,N_19968,N_19567);
or UO_1988 (O_1988,N_19931,N_19868);
nand UO_1989 (O_1989,N_19933,N_19578);
and UO_1990 (O_1990,N_19953,N_19796);
nor UO_1991 (O_1991,N_19788,N_19987);
xor UO_1992 (O_1992,N_19899,N_19626);
or UO_1993 (O_1993,N_19978,N_19665);
and UO_1994 (O_1994,N_19914,N_19911);
nor UO_1995 (O_1995,N_19974,N_19971);
nand UO_1996 (O_1996,N_19703,N_19989);
nand UO_1997 (O_1997,N_19883,N_19877);
and UO_1998 (O_1998,N_19685,N_19984);
and UO_1999 (O_1999,N_19551,N_19867);
nor UO_2000 (O_2000,N_19911,N_19525);
or UO_2001 (O_2001,N_19948,N_19832);
nor UO_2002 (O_2002,N_19845,N_19683);
and UO_2003 (O_2003,N_19816,N_19676);
xnor UO_2004 (O_2004,N_19904,N_19633);
nand UO_2005 (O_2005,N_19937,N_19557);
nand UO_2006 (O_2006,N_19983,N_19642);
nor UO_2007 (O_2007,N_19572,N_19576);
xor UO_2008 (O_2008,N_19892,N_19521);
nor UO_2009 (O_2009,N_19955,N_19993);
xnor UO_2010 (O_2010,N_19929,N_19918);
and UO_2011 (O_2011,N_19941,N_19514);
xor UO_2012 (O_2012,N_19735,N_19775);
and UO_2013 (O_2013,N_19823,N_19581);
and UO_2014 (O_2014,N_19848,N_19823);
xnor UO_2015 (O_2015,N_19721,N_19704);
and UO_2016 (O_2016,N_19523,N_19891);
and UO_2017 (O_2017,N_19527,N_19658);
xor UO_2018 (O_2018,N_19769,N_19674);
xor UO_2019 (O_2019,N_19751,N_19838);
and UO_2020 (O_2020,N_19916,N_19684);
nand UO_2021 (O_2021,N_19768,N_19938);
xor UO_2022 (O_2022,N_19547,N_19729);
and UO_2023 (O_2023,N_19548,N_19541);
nor UO_2024 (O_2024,N_19615,N_19989);
and UO_2025 (O_2025,N_19558,N_19839);
xnor UO_2026 (O_2026,N_19571,N_19798);
or UO_2027 (O_2027,N_19889,N_19814);
xor UO_2028 (O_2028,N_19793,N_19954);
nand UO_2029 (O_2029,N_19620,N_19627);
xor UO_2030 (O_2030,N_19878,N_19727);
and UO_2031 (O_2031,N_19508,N_19744);
or UO_2032 (O_2032,N_19564,N_19963);
nor UO_2033 (O_2033,N_19836,N_19621);
nor UO_2034 (O_2034,N_19696,N_19693);
and UO_2035 (O_2035,N_19582,N_19993);
nand UO_2036 (O_2036,N_19846,N_19966);
or UO_2037 (O_2037,N_19752,N_19697);
nor UO_2038 (O_2038,N_19502,N_19762);
xnor UO_2039 (O_2039,N_19863,N_19879);
nor UO_2040 (O_2040,N_19512,N_19822);
or UO_2041 (O_2041,N_19736,N_19567);
or UO_2042 (O_2042,N_19857,N_19965);
nand UO_2043 (O_2043,N_19527,N_19502);
nor UO_2044 (O_2044,N_19568,N_19599);
or UO_2045 (O_2045,N_19559,N_19724);
or UO_2046 (O_2046,N_19525,N_19722);
nand UO_2047 (O_2047,N_19566,N_19989);
or UO_2048 (O_2048,N_19658,N_19712);
or UO_2049 (O_2049,N_19978,N_19766);
nor UO_2050 (O_2050,N_19614,N_19897);
and UO_2051 (O_2051,N_19642,N_19880);
or UO_2052 (O_2052,N_19515,N_19709);
nand UO_2053 (O_2053,N_19920,N_19793);
nand UO_2054 (O_2054,N_19754,N_19821);
and UO_2055 (O_2055,N_19861,N_19879);
nand UO_2056 (O_2056,N_19848,N_19536);
or UO_2057 (O_2057,N_19651,N_19520);
nand UO_2058 (O_2058,N_19877,N_19754);
and UO_2059 (O_2059,N_19526,N_19667);
or UO_2060 (O_2060,N_19781,N_19700);
nor UO_2061 (O_2061,N_19888,N_19726);
nor UO_2062 (O_2062,N_19619,N_19811);
and UO_2063 (O_2063,N_19626,N_19805);
nand UO_2064 (O_2064,N_19931,N_19598);
nand UO_2065 (O_2065,N_19986,N_19597);
and UO_2066 (O_2066,N_19696,N_19811);
xor UO_2067 (O_2067,N_19852,N_19545);
and UO_2068 (O_2068,N_19532,N_19501);
nand UO_2069 (O_2069,N_19837,N_19538);
xnor UO_2070 (O_2070,N_19879,N_19844);
and UO_2071 (O_2071,N_19808,N_19729);
and UO_2072 (O_2072,N_19928,N_19709);
nor UO_2073 (O_2073,N_19972,N_19919);
nor UO_2074 (O_2074,N_19758,N_19746);
nor UO_2075 (O_2075,N_19597,N_19807);
and UO_2076 (O_2076,N_19993,N_19780);
nor UO_2077 (O_2077,N_19746,N_19856);
nand UO_2078 (O_2078,N_19788,N_19941);
and UO_2079 (O_2079,N_19868,N_19506);
or UO_2080 (O_2080,N_19858,N_19860);
nor UO_2081 (O_2081,N_19599,N_19754);
nand UO_2082 (O_2082,N_19545,N_19749);
nor UO_2083 (O_2083,N_19971,N_19700);
nand UO_2084 (O_2084,N_19618,N_19633);
nand UO_2085 (O_2085,N_19821,N_19715);
xnor UO_2086 (O_2086,N_19916,N_19981);
nand UO_2087 (O_2087,N_19678,N_19919);
or UO_2088 (O_2088,N_19786,N_19582);
nor UO_2089 (O_2089,N_19882,N_19774);
nor UO_2090 (O_2090,N_19642,N_19500);
nand UO_2091 (O_2091,N_19590,N_19842);
nand UO_2092 (O_2092,N_19883,N_19791);
nand UO_2093 (O_2093,N_19894,N_19817);
nand UO_2094 (O_2094,N_19621,N_19852);
xor UO_2095 (O_2095,N_19730,N_19812);
xor UO_2096 (O_2096,N_19825,N_19522);
xor UO_2097 (O_2097,N_19686,N_19905);
nand UO_2098 (O_2098,N_19796,N_19881);
or UO_2099 (O_2099,N_19685,N_19513);
or UO_2100 (O_2100,N_19503,N_19645);
nand UO_2101 (O_2101,N_19529,N_19882);
xor UO_2102 (O_2102,N_19720,N_19925);
or UO_2103 (O_2103,N_19915,N_19799);
xnor UO_2104 (O_2104,N_19631,N_19932);
or UO_2105 (O_2105,N_19525,N_19631);
nand UO_2106 (O_2106,N_19849,N_19601);
and UO_2107 (O_2107,N_19597,N_19609);
and UO_2108 (O_2108,N_19917,N_19740);
nand UO_2109 (O_2109,N_19988,N_19879);
or UO_2110 (O_2110,N_19666,N_19541);
nor UO_2111 (O_2111,N_19527,N_19846);
and UO_2112 (O_2112,N_19582,N_19840);
or UO_2113 (O_2113,N_19737,N_19994);
nor UO_2114 (O_2114,N_19936,N_19828);
xnor UO_2115 (O_2115,N_19872,N_19637);
xor UO_2116 (O_2116,N_19587,N_19753);
and UO_2117 (O_2117,N_19668,N_19821);
or UO_2118 (O_2118,N_19976,N_19923);
and UO_2119 (O_2119,N_19706,N_19740);
or UO_2120 (O_2120,N_19831,N_19943);
and UO_2121 (O_2121,N_19543,N_19685);
xnor UO_2122 (O_2122,N_19948,N_19926);
nand UO_2123 (O_2123,N_19888,N_19685);
xnor UO_2124 (O_2124,N_19729,N_19896);
or UO_2125 (O_2125,N_19875,N_19821);
nor UO_2126 (O_2126,N_19524,N_19714);
nor UO_2127 (O_2127,N_19916,N_19851);
and UO_2128 (O_2128,N_19927,N_19565);
nor UO_2129 (O_2129,N_19529,N_19728);
nand UO_2130 (O_2130,N_19713,N_19553);
nor UO_2131 (O_2131,N_19597,N_19892);
or UO_2132 (O_2132,N_19678,N_19644);
xor UO_2133 (O_2133,N_19955,N_19854);
xnor UO_2134 (O_2134,N_19549,N_19778);
and UO_2135 (O_2135,N_19806,N_19660);
and UO_2136 (O_2136,N_19570,N_19643);
xnor UO_2137 (O_2137,N_19516,N_19767);
xnor UO_2138 (O_2138,N_19761,N_19643);
and UO_2139 (O_2139,N_19867,N_19566);
and UO_2140 (O_2140,N_19715,N_19807);
and UO_2141 (O_2141,N_19545,N_19858);
or UO_2142 (O_2142,N_19625,N_19788);
and UO_2143 (O_2143,N_19812,N_19629);
xor UO_2144 (O_2144,N_19597,N_19801);
xnor UO_2145 (O_2145,N_19518,N_19580);
nand UO_2146 (O_2146,N_19911,N_19631);
xor UO_2147 (O_2147,N_19720,N_19943);
xnor UO_2148 (O_2148,N_19664,N_19631);
and UO_2149 (O_2149,N_19512,N_19668);
and UO_2150 (O_2150,N_19818,N_19771);
nand UO_2151 (O_2151,N_19927,N_19967);
xnor UO_2152 (O_2152,N_19683,N_19625);
or UO_2153 (O_2153,N_19613,N_19874);
nand UO_2154 (O_2154,N_19719,N_19687);
nor UO_2155 (O_2155,N_19712,N_19663);
xor UO_2156 (O_2156,N_19598,N_19624);
nor UO_2157 (O_2157,N_19759,N_19669);
nor UO_2158 (O_2158,N_19813,N_19860);
nor UO_2159 (O_2159,N_19854,N_19785);
and UO_2160 (O_2160,N_19799,N_19674);
xor UO_2161 (O_2161,N_19548,N_19557);
nand UO_2162 (O_2162,N_19580,N_19574);
xnor UO_2163 (O_2163,N_19922,N_19962);
nor UO_2164 (O_2164,N_19536,N_19718);
nor UO_2165 (O_2165,N_19541,N_19999);
nor UO_2166 (O_2166,N_19525,N_19762);
or UO_2167 (O_2167,N_19601,N_19784);
or UO_2168 (O_2168,N_19617,N_19648);
nand UO_2169 (O_2169,N_19649,N_19597);
nand UO_2170 (O_2170,N_19582,N_19777);
xnor UO_2171 (O_2171,N_19636,N_19575);
nor UO_2172 (O_2172,N_19772,N_19819);
nand UO_2173 (O_2173,N_19794,N_19919);
or UO_2174 (O_2174,N_19964,N_19695);
nor UO_2175 (O_2175,N_19717,N_19799);
nor UO_2176 (O_2176,N_19724,N_19842);
or UO_2177 (O_2177,N_19630,N_19738);
or UO_2178 (O_2178,N_19938,N_19908);
and UO_2179 (O_2179,N_19728,N_19794);
or UO_2180 (O_2180,N_19630,N_19547);
nor UO_2181 (O_2181,N_19918,N_19653);
and UO_2182 (O_2182,N_19969,N_19794);
nand UO_2183 (O_2183,N_19848,N_19974);
nor UO_2184 (O_2184,N_19657,N_19742);
or UO_2185 (O_2185,N_19842,N_19980);
xnor UO_2186 (O_2186,N_19832,N_19521);
nand UO_2187 (O_2187,N_19761,N_19717);
or UO_2188 (O_2188,N_19993,N_19683);
nand UO_2189 (O_2189,N_19765,N_19739);
and UO_2190 (O_2190,N_19602,N_19703);
or UO_2191 (O_2191,N_19543,N_19587);
nand UO_2192 (O_2192,N_19700,N_19540);
nand UO_2193 (O_2193,N_19873,N_19854);
nor UO_2194 (O_2194,N_19767,N_19701);
xor UO_2195 (O_2195,N_19634,N_19946);
or UO_2196 (O_2196,N_19571,N_19575);
and UO_2197 (O_2197,N_19970,N_19764);
and UO_2198 (O_2198,N_19892,N_19938);
nor UO_2199 (O_2199,N_19929,N_19517);
nand UO_2200 (O_2200,N_19562,N_19633);
nand UO_2201 (O_2201,N_19957,N_19775);
or UO_2202 (O_2202,N_19959,N_19729);
and UO_2203 (O_2203,N_19681,N_19784);
or UO_2204 (O_2204,N_19810,N_19521);
xor UO_2205 (O_2205,N_19968,N_19752);
xor UO_2206 (O_2206,N_19924,N_19690);
or UO_2207 (O_2207,N_19651,N_19920);
or UO_2208 (O_2208,N_19840,N_19975);
xor UO_2209 (O_2209,N_19911,N_19643);
nor UO_2210 (O_2210,N_19601,N_19647);
or UO_2211 (O_2211,N_19914,N_19742);
xnor UO_2212 (O_2212,N_19848,N_19960);
nand UO_2213 (O_2213,N_19624,N_19850);
nor UO_2214 (O_2214,N_19705,N_19851);
and UO_2215 (O_2215,N_19576,N_19695);
and UO_2216 (O_2216,N_19908,N_19812);
and UO_2217 (O_2217,N_19671,N_19512);
xnor UO_2218 (O_2218,N_19608,N_19537);
and UO_2219 (O_2219,N_19617,N_19643);
xor UO_2220 (O_2220,N_19614,N_19932);
xnor UO_2221 (O_2221,N_19973,N_19864);
and UO_2222 (O_2222,N_19587,N_19595);
nor UO_2223 (O_2223,N_19779,N_19979);
xor UO_2224 (O_2224,N_19685,N_19943);
or UO_2225 (O_2225,N_19858,N_19969);
nand UO_2226 (O_2226,N_19557,N_19733);
or UO_2227 (O_2227,N_19902,N_19874);
or UO_2228 (O_2228,N_19979,N_19890);
xnor UO_2229 (O_2229,N_19734,N_19942);
xnor UO_2230 (O_2230,N_19702,N_19845);
and UO_2231 (O_2231,N_19901,N_19521);
and UO_2232 (O_2232,N_19736,N_19854);
nand UO_2233 (O_2233,N_19634,N_19821);
and UO_2234 (O_2234,N_19701,N_19707);
nor UO_2235 (O_2235,N_19990,N_19842);
and UO_2236 (O_2236,N_19597,N_19958);
and UO_2237 (O_2237,N_19509,N_19533);
nor UO_2238 (O_2238,N_19949,N_19578);
nor UO_2239 (O_2239,N_19939,N_19984);
xnor UO_2240 (O_2240,N_19620,N_19819);
nor UO_2241 (O_2241,N_19560,N_19817);
nor UO_2242 (O_2242,N_19706,N_19986);
nand UO_2243 (O_2243,N_19853,N_19507);
xor UO_2244 (O_2244,N_19679,N_19548);
xnor UO_2245 (O_2245,N_19623,N_19951);
nor UO_2246 (O_2246,N_19565,N_19863);
and UO_2247 (O_2247,N_19932,N_19740);
nand UO_2248 (O_2248,N_19603,N_19505);
or UO_2249 (O_2249,N_19995,N_19817);
nand UO_2250 (O_2250,N_19907,N_19963);
nor UO_2251 (O_2251,N_19836,N_19676);
or UO_2252 (O_2252,N_19596,N_19563);
xnor UO_2253 (O_2253,N_19670,N_19537);
and UO_2254 (O_2254,N_19656,N_19596);
and UO_2255 (O_2255,N_19858,N_19924);
or UO_2256 (O_2256,N_19890,N_19784);
xnor UO_2257 (O_2257,N_19568,N_19838);
nand UO_2258 (O_2258,N_19654,N_19544);
or UO_2259 (O_2259,N_19956,N_19554);
xnor UO_2260 (O_2260,N_19545,N_19842);
and UO_2261 (O_2261,N_19559,N_19738);
nand UO_2262 (O_2262,N_19665,N_19812);
and UO_2263 (O_2263,N_19979,N_19532);
nand UO_2264 (O_2264,N_19765,N_19821);
or UO_2265 (O_2265,N_19986,N_19585);
nand UO_2266 (O_2266,N_19863,N_19800);
or UO_2267 (O_2267,N_19575,N_19548);
nand UO_2268 (O_2268,N_19958,N_19698);
and UO_2269 (O_2269,N_19777,N_19929);
nor UO_2270 (O_2270,N_19926,N_19505);
nand UO_2271 (O_2271,N_19950,N_19860);
xnor UO_2272 (O_2272,N_19615,N_19727);
or UO_2273 (O_2273,N_19966,N_19953);
or UO_2274 (O_2274,N_19672,N_19930);
xor UO_2275 (O_2275,N_19945,N_19772);
nor UO_2276 (O_2276,N_19741,N_19937);
nor UO_2277 (O_2277,N_19961,N_19554);
nor UO_2278 (O_2278,N_19573,N_19637);
nand UO_2279 (O_2279,N_19798,N_19906);
nor UO_2280 (O_2280,N_19906,N_19832);
nor UO_2281 (O_2281,N_19565,N_19914);
xnor UO_2282 (O_2282,N_19670,N_19971);
xor UO_2283 (O_2283,N_19804,N_19895);
nor UO_2284 (O_2284,N_19878,N_19532);
nand UO_2285 (O_2285,N_19611,N_19618);
or UO_2286 (O_2286,N_19863,N_19620);
xor UO_2287 (O_2287,N_19686,N_19733);
nor UO_2288 (O_2288,N_19593,N_19758);
or UO_2289 (O_2289,N_19940,N_19799);
xnor UO_2290 (O_2290,N_19529,N_19780);
nand UO_2291 (O_2291,N_19711,N_19516);
or UO_2292 (O_2292,N_19537,N_19559);
and UO_2293 (O_2293,N_19762,N_19639);
nand UO_2294 (O_2294,N_19697,N_19514);
nand UO_2295 (O_2295,N_19742,N_19896);
and UO_2296 (O_2296,N_19819,N_19870);
nand UO_2297 (O_2297,N_19570,N_19675);
xor UO_2298 (O_2298,N_19608,N_19545);
xnor UO_2299 (O_2299,N_19628,N_19921);
nor UO_2300 (O_2300,N_19607,N_19705);
or UO_2301 (O_2301,N_19794,N_19631);
xor UO_2302 (O_2302,N_19856,N_19914);
nand UO_2303 (O_2303,N_19587,N_19834);
xor UO_2304 (O_2304,N_19852,N_19968);
and UO_2305 (O_2305,N_19672,N_19926);
nor UO_2306 (O_2306,N_19964,N_19865);
xor UO_2307 (O_2307,N_19508,N_19670);
or UO_2308 (O_2308,N_19970,N_19953);
or UO_2309 (O_2309,N_19669,N_19566);
nand UO_2310 (O_2310,N_19834,N_19681);
nand UO_2311 (O_2311,N_19759,N_19674);
nor UO_2312 (O_2312,N_19736,N_19805);
nor UO_2313 (O_2313,N_19828,N_19948);
and UO_2314 (O_2314,N_19957,N_19567);
or UO_2315 (O_2315,N_19834,N_19544);
or UO_2316 (O_2316,N_19729,N_19794);
or UO_2317 (O_2317,N_19756,N_19932);
and UO_2318 (O_2318,N_19666,N_19538);
nor UO_2319 (O_2319,N_19817,N_19749);
xor UO_2320 (O_2320,N_19863,N_19543);
nand UO_2321 (O_2321,N_19696,N_19714);
or UO_2322 (O_2322,N_19746,N_19839);
and UO_2323 (O_2323,N_19819,N_19701);
nor UO_2324 (O_2324,N_19607,N_19870);
and UO_2325 (O_2325,N_19858,N_19964);
nor UO_2326 (O_2326,N_19676,N_19910);
nor UO_2327 (O_2327,N_19825,N_19720);
xnor UO_2328 (O_2328,N_19825,N_19500);
xnor UO_2329 (O_2329,N_19559,N_19839);
or UO_2330 (O_2330,N_19872,N_19615);
nand UO_2331 (O_2331,N_19981,N_19544);
and UO_2332 (O_2332,N_19849,N_19721);
xor UO_2333 (O_2333,N_19781,N_19860);
nand UO_2334 (O_2334,N_19681,N_19778);
or UO_2335 (O_2335,N_19871,N_19508);
or UO_2336 (O_2336,N_19715,N_19515);
nor UO_2337 (O_2337,N_19874,N_19690);
and UO_2338 (O_2338,N_19929,N_19685);
nand UO_2339 (O_2339,N_19546,N_19979);
or UO_2340 (O_2340,N_19816,N_19902);
or UO_2341 (O_2341,N_19581,N_19839);
and UO_2342 (O_2342,N_19685,N_19860);
or UO_2343 (O_2343,N_19810,N_19954);
and UO_2344 (O_2344,N_19621,N_19847);
or UO_2345 (O_2345,N_19505,N_19911);
xnor UO_2346 (O_2346,N_19959,N_19585);
nor UO_2347 (O_2347,N_19534,N_19860);
and UO_2348 (O_2348,N_19751,N_19567);
or UO_2349 (O_2349,N_19651,N_19901);
xor UO_2350 (O_2350,N_19787,N_19908);
nor UO_2351 (O_2351,N_19893,N_19919);
or UO_2352 (O_2352,N_19946,N_19537);
or UO_2353 (O_2353,N_19569,N_19628);
and UO_2354 (O_2354,N_19776,N_19595);
or UO_2355 (O_2355,N_19773,N_19712);
xor UO_2356 (O_2356,N_19837,N_19894);
nor UO_2357 (O_2357,N_19768,N_19775);
and UO_2358 (O_2358,N_19527,N_19681);
nand UO_2359 (O_2359,N_19821,N_19999);
and UO_2360 (O_2360,N_19983,N_19810);
and UO_2361 (O_2361,N_19816,N_19711);
and UO_2362 (O_2362,N_19830,N_19663);
nor UO_2363 (O_2363,N_19869,N_19536);
xnor UO_2364 (O_2364,N_19787,N_19665);
nand UO_2365 (O_2365,N_19506,N_19563);
nand UO_2366 (O_2366,N_19629,N_19674);
nor UO_2367 (O_2367,N_19625,N_19513);
and UO_2368 (O_2368,N_19989,N_19993);
nand UO_2369 (O_2369,N_19826,N_19544);
or UO_2370 (O_2370,N_19632,N_19709);
and UO_2371 (O_2371,N_19970,N_19606);
and UO_2372 (O_2372,N_19730,N_19757);
xor UO_2373 (O_2373,N_19992,N_19862);
and UO_2374 (O_2374,N_19595,N_19661);
or UO_2375 (O_2375,N_19607,N_19552);
nand UO_2376 (O_2376,N_19505,N_19763);
nand UO_2377 (O_2377,N_19684,N_19667);
xor UO_2378 (O_2378,N_19703,N_19923);
or UO_2379 (O_2379,N_19945,N_19886);
or UO_2380 (O_2380,N_19881,N_19838);
or UO_2381 (O_2381,N_19562,N_19641);
and UO_2382 (O_2382,N_19937,N_19687);
xor UO_2383 (O_2383,N_19691,N_19504);
xnor UO_2384 (O_2384,N_19865,N_19833);
or UO_2385 (O_2385,N_19631,N_19669);
xor UO_2386 (O_2386,N_19623,N_19973);
xnor UO_2387 (O_2387,N_19869,N_19597);
or UO_2388 (O_2388,N_19630,N_19583);
nor UO_2389 (O_2389,N_19698,N_19633);
and UO_2390 (O_2390,N_19839,N_19926);
nand UO_2391 (O_2391,N_19685,N_19809);
or UO_2392 (O_2392,N_19519,N_19524);
xnor UO_2393 (O_2393,N_19958,N_19942);
nand UO_2394 (O_2394,N_19981,N_19795);
nand UO_2395 (O_2395,N_19763,N_19599);
or UO_2396 (O_2396,N_19752,N_19516);
nor UO_2397 (O_2397,N_19731,N_19602);
xnor UO_2398 (O_2398,N_19770,N_19696);
and UO_2399 (O_2399,N_19944,N_19578);
nor UO_2400 (O_2400,N_19911,N_19833);
and UO_2401 (O_2401,N_19982,N_19845);
nor UO_2402 (O_2402,N_19895,N_19616);
and UO_2403 (O_2403,N_19856,N_19516);
or UO_2404 (O_2404,N_19632,N_19794);
and UO_2405 (O_2405,N_19612,N_19629);
nor UO_2406 (O_2406,N_19574,N_19845);
or UO_2407 (O_2407,N_19913,N_19554);
nand UO_2408 (O_2408,N_19587,N_19907);
nor UO_2409 (O_2409,N_19912,N_19647);
nor UO_2410 (O_2410,N_19681,N_19633);
or UO_2411 (O_2411,N_19615,N_19651);
and UO_2412 (O_2412,N_19862,N_19781);
xnor UO_2413 (O_2413,N_19869,N_19652);
and UO_2414 (O_2414,N_19870,N_19542);
xor UO_2415 (O_2415,N_19932,N_19717);
nor UO_2416 (O_2416,N_19897,N_19566);
xor UO_2417 (O_2417,N_19579,N_19726);
or UO_2418 (O_2418,N_19905,N_19545);
xor UO_2419 (O_2419,N_19879,N_19530);
nor UO_2420 (O_2420,N_19593,N_19621);
xor UO_2421 (O_2421,N_19538,N_19658);
and UO_2422 (O_2422,N_19891,N_19671);
nor UO_2423 (O_2423,N_19581,N_19774);
nor UO_2424 (O_2424,N_19846,N_19610);
or UO_2425 (O_2425,N_19692,N_19553);
nand UO_2426 (O_2426,N_19869,N_19898);
xnor UO_2427 (O_2427,N_19703,N_19757);
nand UO_2428 (O_2428,N_19633,N_19993);
or UO_2429 (O_2429,N_19954,N_19607);
nand UO_2430 (O_2430,N_19864,N_19895);
nor UO_2431 (O_2431,N_19666,N_19709);
and UO_2432 (O_2432,N_19898,N_19525);
and UO_2433 (O_2433,N_19936,N_19880);
and UO_2434 (O_2434,N_19910,N_19566);
nand UO_2435 (O_2435,N_19619,N_19982);
xor UO_2436 (O_2436,N_19959,N_19920);
nand UO_2437 (O_2437,N_19971,N_19927);
xnor UO_2438 (O_2438,N_19658,N_19724);
nor UO_2439 (O_2439,N_19521,N_19589);
nand UO_2440 (O_2440,N_19967,N_19932);
nor UO_2441 (O_2441,N_19702,N_19576);
nand UO_2442 (O_2442,N_19946,N_19867);
xnor UO_2443 (O_2443,N_19886,N_19545);
or UO_2444 (O_2444,N_19891,N_19812);
and UO_2445 (O_2445,N_19856,N_19786);
or UO_2446 (O_2446,N_19834,N_19580);
nor UO_2447 (O_2447,N_19697,N_19687);
and UO_2448 (O_2448,N_19662,N_19944);
nor UO_2449 (O_2449,N_19853,N_19550);
xnor UO_2450 (O_2450,N_19766,N_19612);
and UO_2451 (O_2451,N_19862,N_19607);
nand UO_2452 (O_2452,N_19827,N_19765);
and UO_2453 (O_2453,N_19898,N_19880);
nor UO_2454 (O_2454,N_19750,N_19809);
nor UO_2455 (O_2455,N_19535,N_19812);
and UO_2456 (O_2456,N_19594,N_19825);
and UO_2457 (O_2457,N_19900,N_19605);
or UO_2458 (O_2458,N_19816,N_19957);
nand UO_2459 (O_2459,N_19640,N_19761);
nand UO_2460 (O_2460,N_19586,N_19516);
nor UO_2461 (O_2461,N_19792,N_19724);
nor UO_2462 (O_2462,N_19535,N_19770);
and UO_2463 (O_2463,N_19729,N_19985);
nand UO_2464 (O_2464,N_19607,N_19528);
or UO_2465 (O_2465,N_19846,N_19892);
nand UO_2466 (O_2466,N_19893,N_19693);
or UO_2467 (O_2467,N_19574,N_19835);
or UO_2468 (O_2468,N_19665,N_19734);
nor UO_2469 (O_2469,N_19541,N_19706);
xnor UO_2470 (O_2470,N_19781,N_19699);
or UO_2471 (O_2471,N_19600,N_19747);
nand UO_2472 (O_2472,N_19708,N_19573);
nand UO_2473 (O_2473,N_19716,N_19849);
nor UO_2474 (O_2474,N_19518,N_19680);
nor UO_2475 (O_2475,N_19569,N_19676);
xnor UO_2476 (O_2476,N_19538,N_19730);
and UO_2477 (O_2477,N_19710,N_19595);
nand UO_2478 (O_2478,N_19893,N_19896);
nor UO_2479 (O_2479,N_19989,N_19876);
or UO_2480 (O_2480,N_19861,N_19539);
nor UO_2481 (O_2481,N_19662,N_19946);
nand UO_2482 (O_2482,N_19989,N_19601);
and UO_2483 (O_2483,N_19789,N_19647);
xnor UO_2484 (O_2484,N_19648,N_19705);
xnor UO_2485 (O_2485,N_19505,N_19742);
nor UO_2486 (O_2486,N_19772,N_19561);
nand UO_2487 (O_2487,N_19753,N_19656);
nand UO_2488 (O_2488,N_19849,N_19737);
and UO_2489 (O_2489,N_19971,N_19747);
xnor UO_2490 (O_2490,N_19848,N_19836);
and UO_2491 (O_2491,N_19624,N_19519);
and UO_2492 (O_2492,N_19757,N_19768);
and UO_2493 (O_2493,N_19995,N_19847);
xor UO_2494 (O_2494,N_19687,N_19639);
and UO_2495 (O_2495,N_19525,N_19790);
nor UO_2496 (O_2496,N_19595,N_19782);
nand UO_2497 (O_2497,N_19619,N_19766);
nand UO_2498 (O_2498,N_19854,N_19998);
nand UO_2499 (O_2499,N_19946,N_19805);
endmodule