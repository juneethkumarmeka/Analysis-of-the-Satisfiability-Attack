module basic_2000_20000_2500_50_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1120,In_1708);
nor U1 (N_1,In_830,In_1875);
nor U2 (N_2,In_1350,In_461);
nor U3 (N_3,In_1726,In_1964);
nor U4 (N_4,In_1476,In_482);
xor U5 (N_5,In_692,In_255);
nor U6 (N_6,In_1075,In_242);
and U7 (N_7,In_1689,In_1683);
xor U8 (N_8,In_349,In_391);
and U9 (N_9,In_1157,In_1381);
xnor U10 (N_10,In_1042,In_1436);
and U11 (N_11,In_173,In_1405);
xnor U12 (N_12,In_164,In_406);
nand U13 (N_13,In_535,In_593);
nor U14 (N_14,In_1718,In_12);
nand U15 (N_15,In_1428,In_1010);
nor U16 (N_16,In_656,In_1859);
and U17 (N_17,In_1809,In_452);
nor U18 (N_18,In_1071,In_329);
nor U19 (N_19,In_390,In_1206);
and U20 (N_20,In_757,In_202);
nand U21 (N_21,In_106,In_923);
nand U22 (N_22,In_1679,In_1722);
nor U23 (N_23,In_1976,In_1560);
xor U24 (N_24,In_1985,In_849);
and U25 (N_25,In_243,In_895);
xor U26 (N_26,In_416,In_1946);
nand U27 (N_27,In_1914,In_1880);
and U28 (N_28,In_1303,In_909);
and U29 (N_29,In_1281,In_1558);
or U30 (N_30,In_940,In_1314);
and U31 (N_31,In_1928,In_170);
nand U32 (N_32,In_401,In_1612);
or U33 (N_33,In_301,In_181);
xnor U34 (N_34,In_687,In_1421);
and U35 (N_35,In_1944,In_98);
xor U36 (N_36,In_1721,In_525);
and U37 (N_37,In_477,In_1579);
or U38 (N_38,In_671,In_1838);
xnor U39 (N_39,In_344,In_1854);
nor U40 (N_40,In_90,In_604);
nand U41 (N_41,In_1248,In_572);
xor U42 (N_42,In_1299,In_1237);
nor U43 (N_43,In_858,In_882);
nand U44 (N_44,In_26,In_188);
or U45 (N_45,In_1796,In_1040);
and U46 (N_46,In_1929,In_967);
xor U47 (N_47,In_1063,In_636);
nand U48 (N_48,In_1592,In_786);
xnor U49 (N_49,In_373,In_705);
nor U50 (N_50,In_558,In_1007);
or U51 (N_51,In_1958,In_567);
and U52 (N_52,In_532,In_1141);
nor U53 (N_53,In_1639,In_163);
or U54 (N_54,In_330,In_854);
and U55 (N_55,In_733,In_1348);
nand U56 (N_56,In_1247,In_856);
and U57 (N_57,In_260,In_1296);
nor U58 (N_58,In_1834,In_1680);
xor U59 (N_59,In_1054,In_1917);
nor U60 (N_60,In_792,In_1511);
xnor U61 (N_61,In_1886,In_1410);
nor U62 (N_62,In_1474,In_156);
xnor U63 (N_63,In_337,In_198);
xor U64 (N_64,In_980,In_884);
or U65 (N_65,In_965,In_500);
and U66 (N_66,In_113,In_916);
or U67 (N_67,In_75,In_828);
xnor U68 (N_68,In_353,In_54);
or U69 (N_69,In_1670,In_1764);
xnor U70 (N_70,In_1083,In_1619);
nor U71 (N_71,In_1665,In_1218);
xor U72 (N_72,In_1242,In_1530);
and U73 (N_73,In_1290,In_928);
nor U74 (N_74,In_1549,In_455);
or U75 (N_75,In_777,In_1351);
nor U76 (N_76,In_1598,In_1266);
and U77 (N_77,In_1447,In_1938);
and U78 (N_78,In_819,In_859);
or U79 (N_79,In_1165,In_1635);
and U80 (N_80,In_1261,In_30);
and U81 (N_81,In_1467,In_627);
nand U82 (N_82,In_1224,In_1481);
nor U83 (N_83,In_538,In_938);
xnor U84 (N_84,In_1401,In_557);
xor U85 (N_85,In_683,In_708);
and U86 (N_86,In_1716,In_738);
nor U87 (N_87,In_465,In_1170);
nand U88 (N_88,In_1438,In_843);
nor U89 (N_89,In_643,In_1426);
nor U90 (N_90,In_1647,In_620);
nand U91 (N_91,In_1143,In_237);
xnor U92 (N_92,In_1995,In_56);
nor U93 (N_93,In_1545,In_597);
and U94 (N_94,In_817,In_1738);
or U95 (N_95,In_1264,In_1115);
xor U96 (N_96,In_1769,In_224);
nand U97 (N_97,In_1110,In_363);
nand U98 (N_98,In_1860,In_1927);
or U99 (N_99,In_1525,In_565);
nand U100 (N_100,In_219,In_440);
and U101 (N_101,In_1576,In_1099);
and U102 (N_102,In_991,In_985);
xor U103 (N_103,In_324,In_721);
nor U104 (N_104,In_483,In_434);
or U105 (N_105,In_481,In_1562);
or U106 (N_106,In_602,In_1373);
xor U107 (N_107,In_1111,In_639);
nor U108 (N_108,In_901,In_334);
and U109 (N_109,In_507,In_713);
nand U110 (N_110,In_1888,In_670);
nor U111 (N_111,In_111,In_123);
xnor U112 (N_112,In_1383,In_1203);
xor U113 (N_113,In_262,In_1118);
nand U114 (N_114,In_1319,In_1459);
and U115 (N_115,In_1295,In_40);
and U116 (N_116,In_1322,In_1035);
and U117 (N_117,In_1747,In_1941);
or U118 (N_118,In_99,In_728);
nor U119 (N_119,In_216,In_47);
and U120 (N_120,In_1551,In_821);
xnor U121 (N_121,In_1152,In_190);
or U122 (N_122,In_1105,In_1523);
xnor U123 (N_123,In_1496,In_1030);
nand U124 (N_124,In_1832,In_339);
or U125 (N_125,In_1559,In_448);
nor U126 (N_126,In_905,In_1826);
xnor U127 (N_127,In_199,In_1807);
or U128 (N_128,In_1498,In_1342);
xnor U129 (N_129,In_1900,In_1666);
and U130 (N_130,In_62,In_1116);
or U131 (N_131,In_157,In_1706);
and U132 (N_132,In_1113,In_962);
or U133 (N_133,In_139,In_1132);
or U134 (N_134,In_800,In_1013);
nand U135 (N_135,In_2,In_506);
or U136 (N_136,In_801,In_802);
or U137 (N_137,In_1315,In_679);
and U138 (N_138,In_1090,In_1480);
xor U139 (N_139,In_1869,In_135);
nand U140 (N_140,In_400,In_1114);
nand U141 (N_141,In_1049,In_89);
or U142 (N_142,In_539,In_931);
xnor U143 (N_143,In_114,In_1603);
xor U144 (N_144,In_1181,In_1509);
nor U145 (N_145,In_887,In_1973);
or U146 (N_146,In_575,In_678);
or U147 (N_147,In_1044,In_1258);
or U148 (N_148,In_1901,In_1389);
nand U149 (N_149,In_529,In_1778);
or U150 (N_150,In_630,In_1332);
xor U151 (N_151,In_1257,In_1624);
xnor U152 (N_152,In_823,In_1546);
or U153 (N_153,In_1978,In_1338);
nand U154 (N_154,In_841,In_881);
nor U155 (N_155,In_1800,In_212);
nor U156 (N_156,In_1024,In_453);
nor U157 (N_157,In_977,In_537);
nor U158 (N_158,In_1799,In_205);
and U159 (N_159,In_327,In_1423);
xnor U160 (N_160,In_193,In_1210);
xnor U161 (N_161,In_1171,In_356);
nor U162 (N_162,In_16,In_807);
or U163 (N_163,In_1164,In_394);
nand U164 (N_164,In_1411,In_183);
nor U165 (N_165,In_1448,In_6);
nand U166 (N_166,In_1297,In_1369);
nand U167 (N_167,In_291,In_1824);
nand U168 (N_168,In_1121,In_893);
or U169 (N_169,In_421,In_1513);
xnor U170 (N_170,In_1067,In_1821);
or U171 (N_171,In_1653,In_1881);
xnor U172 (N_172,In_1632,In_413);
nor U173 (N_173,In_848,In_367);
nor U174 (N_174,In_4,In_542);
xor U175 (N_175,In_694,In_1001);
nor U176 (N_176,In_1790,In_340);
nor U177 (N_177,In_1943,In_1623);
or U178 (N_178,In_1845,In_1034);
nand U179 (N_179,In_274,In_302);
or U180 (N_180,In_1980,In_459);
or U181 (N_181,In_1056,In_997);
xnor U182 (N_182,In_1762,In_517);
xor U183 (N_183,In_96,In_1740);
nand U184 (N_184,In_1966,In_982);
and U185 (N_185,In_343,In_571);
nand U186 (N_186,In_499,In_1503);
or U187 (N_187,In_601,In_298);
nor U188 (N_188,In_650,In_402);
nand U189 (N_189,In_215,In_812);
and U190 (N_190,In_1804,In_596);
nand U191 (N_191,In_1555,In_904);
nor U192 (N_192,In_407,In_58);
and U193 (N_193,In_1074,In_1020);
xnor U194 (N_194,In_1419,In_418);
or U195 (N_195,In_171,In_1873);
xnor U196 (N_196,In_303,In_225);
nor U197 (N_197,In_1434,In_1540);
or U198 (N_198,In_559,In_690);
xor U199 (N_199,In_1737,In_700);
nor U200 (N_200,In_1674,In_689);
or U201 (N_201,In_924,In_534);
and U202 (N_202,In_871,In_1940);
xnor U203 (N_203,In_1457,In_1746);
nand U204 (N_204,In_763,In_674);
or U205 (N_205,In_617,In_1771);
xor U206 (N_206,In_1720,In_1786);
nand U207 (N_207,In_1285,In_370);
nand U208 (N_208,In_179,In_1884);
xor U209 (N_209,In_1077,In_1570);
or U210 (N_210,In_119,In_994);
or U211 (N_211,In_1002,In_1173);
xor U212 (N_212,In_844,In_1505);
or U213 (N_213,In_633,In_1161);
nor U214 (N_214,In_1490,In_1777);
or U215 (N_215,In_933,In_1375);
nand U216 (N_216,In_1455,In_257);
nor U217 (N_217,In_974,In_651);
nand U218 (N_218,In_1798,In_1376);
or U219 (N_219,In_874,In_1912);
xnor U220 (N_220,In_1211,In_1705);
nor U221 (N_221,In_839,In_231);
nor U222 (N_222,In_326,In_1953);
and U223 (N_223,In_1649,In_1866);
or U224 (N_224,In_403,In_361);
or U225 (N_225,In_42,In_1844);
xor U226 (N_226,In_1580,In_1364);
or U227 (N_227,In_1877,In_986);
xnor U228 (N_228,In_1420,In_1403);
xor U229 (N_229,In_1318,In_1533);
nand U230 (N_230,In_1456,In_1);
or U231 (N_231,In_714,In_1117);
nand U232 (N_232,In_1156,In_1794);
or U233 (N_233,In_1065,In_1552);
or U234 (N_234,In_5,In_299);
xor U235 (N_235,In_582,In_926);
nor U236 (N_236,In_1500,In_946);
nand U237 (N_237,In_1991,In_1899);
nor U238 (N_238,In_1204,In_153);
or U239 (N_239,In_374,In_1365);
and U240 (N_240,In_1196,In_644);
xnor U241 (N_241,In_655,In_1305);
nand U242 (N_242,In_616,In_1739);
xor U243 (N_243,In_1385,In_1217);
or U244 (N_244,In_428,In_146);
nand U245 (N_245,In_1023,In_509);
and U246 (N_246,In_1353,In_1341);
and U247 (N_247,In_248,In_1952);
and U248 (N_248,In_1774,In_1471);
nor U249 (N_249,In_732,In_1671);
nand U250 (N_250,In_993,In_79);
nor U251 (N_251,In_959,In_140);
nor U252 (N_252,In_1312,In_1249);
nor U253 (N_253,In_1849,In_1803);
or U254 (N_254,In_824,In_625);
or U255 (N_255,In_1634,In_1714);
nor U256 (N_256,In_233,In_427);
or U257 (N_257,In_165,In_1184);
or U258 (N_258,In_491,In_1855);
xnor U259 (N_259,In_463,In_186);
nand U260 (N_260,In_1223,In_1862);
nor U261 (N_261,In_1387,In_355);
nor U262 (N_262,In_116,In_1645);
xnor U263 (N_263,In_781,In_1177);
nand U264 (N_264,In_1470,In_804);
or U265 (N_265,In_868,In_1038);
or U266 (N_266,In_1997,In_1836);
nand U267 (N_267,In_1956,In_835);
xnor U268 (N_268,In_555,In_1144);
xor U269 (N_269,In_531,In_1047);
xor U270 (N_270,In_1911,In_372);
xor U271 (N_271,In_1775,In_587);
nor U272 (N_272,In_725,In_232);
nor U273 (N_273,In_1695,In_570);
or U274 (N_274,In_471,In_270);
or U275 (N_275,In_1112,In_825);
nand U276 (N_276,In_345,In_191);
nor U277 (N_277,In_957,In_386);
nand U278 (N_278,In_1232,In_1835);
nand U279 (N_279,In_1098,In_942);
nor U280 (N_280,In_115,In_1395);
nand U281 (N_281,In_1982,In_654);
and U282 (N_282,In_1532,In_1106);
xnor U283 (N_283,In_1394,In_1374);
nand U284 (N_284,In_1274,In_609);
nand U285 (N_285,In_1402,In_1022);
nand U286 (N_286,In_1923,In_666);
xor U287 (N_287,In_853,In_381);
or U288 (N_288,In_1427,In_1759);
xnor U289 (N_289,In_766,In_1648);
nand U290 (N_290,In_594,In_1664);
nor U291 (N_291,In_328,In_1230);
or U292 (N_292,In_1949,In_9);
and U293 (N_293,In_50,In_1614);
or U294 (N_294,In_1783,In_1418);
and U295 (N_295,In_104,In_863);
or U296 (N_296,In_1898,In_1335);
xnor U297 (N_297,In_526,In_266);
xor U298 (N_298,In_910,In_756);
nor U299 (N_299,In_278,In_1518);
nand U300 (N_300,In_1477,In_1445);
nand U301 (N_301,In_972,In_1306);
and U302 (N_302,In_852,In_624);
xnor U303 (N_303,In_1754,In_1753);
xnor U304 (N_304,In_1602,In_131);
xnor U305 (N_305,In_380,In_1617);
nand U306 (N_306,In_322,In_1735);
xnor U307 (N_307,In_1006,In_684);
nor U308 (N_308,In_1377,In_20);
or U309 (N_309,In_968,In_917);
or U310 (N_310,In_496,In_1717);
or U311 (N_311,In_426,In_321);
or U312 (N_312,In_1086,In_513);
nand U313 (N_313,In_1323,In_672);
nor U314 (N_314,In_251,In_1846);
or U315 (N_315,In_1704,In_1048);
xor U316 (N_316,In_1748,In_945);
and U317 (N_317,In_446,In_1301);
or U318 (N_318,In_281,In_1610);
or U319 (N_319,In_474,In_1159);
xor U320 (N_320,In_488,In_1703);
nand U321 (N_321,In_1693,In_934);
nor U322 (N_322,In_1588,In_1234);
or U323 (N_323,In_1349,In_680);
nand U324 (N_324,In_53,In_1425);
or U325 (N_325,In_1175,In_387);
or U326 (N_326,In_1287,In_80);
or U327 (N_327,In_57,In_1108);
and U328 (N_328,In_192,In_1308);
or U329 (N_329,In_1362,In_516);
or U330 (N_330,In_1524,In_816);
or U331 (N_331,In_1767,In_1616);
or U332 (N_332,In_1300,In_1519);
nor U333 (N_333,In_182,In_127);
xnor U334 (N_334,In_544,In_331);
nand U335 (N_335,In_1586,In_1885);
or U336 (N_336,In_836,In_494);
nand U337 (N_337,In_540,In_1069);
nor U338 (N_338,In_445,In_84);
and U339 (N_339,In_398,In_970);
nand U340 (N_340,In_1864,In_806);
nor U341 (N_341,In_943,In_1270);
or U342 (N_342,In_1221,In_914);
nor U343 (N_343,In_29,In_1313);
and U344 (N_344,In_23,In_748);
nor U345 (N_345,In_15,In_34);
nand U346 (N_346,In_1492,In_1765);
nand U347 (N_347,In_1463,In_336);
xor U348 (N_348,In_1092,In_1220);
nand U349 (N_349,In_950,In_667);
nor U350 (N_350,In_546,In_92);
or U351 (N_351,In_333,In_818);
and U352 (N_352,In_1892,In_285);
or U353 (N_353,In_681,In_1043);
nand U354 (N_354,In_85,In_1137);
xnor U355 (N_355,In_214,In_1730);
and U356 (N_356,In_1605,In_234);
nor U357 (N_357,In_457,In_776);
nor U358 (N_358,In_447,In_1651);
or U359 (N_359,In_963,In_207);
nor U360 (N_360,In_574,In_796);
or U361 (N_361,In_1903,In_1734);
nor U362 (N_362,In_731,In_287);
nand U363 (N_363,In_1593,In_1488);
nand U364 (N_364,In_168,In_898);
nand U365 (N_365,In_605,In_1019);
xor U366 (N_366,In_1930,In_1660);
nor U367 (N_367,In_1228,In_1346);
or U368 (N_368,In_13,In_1667);
xor U369 (N_369,In_1397,In_1378);
nand U370 (N_370,In_133,In_1238);
nand U371 (N_371,In_1131,In_851);
xnor U372 (N_372,In_711,In_951);
nor U373 (N_373,In_675,In_105);
and U374 (N_374,In_1517,In_1025);
xnor U375 (N_375,In_1856,In_1851);
or U376 (N_376,In_1003,In_409);
and U377 (N_377,In_1008,In_989);
nor U378 (N_378,In_809,In_1621);
nor U379 (N_379,In_1727,In_1413);
or U380 (N_380,In_282,In_846);
or U381 (N_381,In_726,In_1850);
nor U382 (N_382,In_696,In_1469);
and U383 (N_383,In_470,In_1415);
and U384 (N_384,In_1878,In_1102);
nand U385 (N_385,In_958,In_1936);
and U386 (N_386,In_1014,In_740);
xor U387 (N_387,In_729,In_896);
nor U388 (N_388,In_919,In_987);
and U389 (N_389,In_318,In_288);
or U390 (N_390,In_1863,In_1449);
nand U391 (N_391,In_1205,In_1654);
nand U392 (N_392,In_867,In_289);
and U393 (N_393,In_912,In_1882);
nor U394 (N_394,In_1245,In_1412);
nand U395 (N_395,In_1999,In_753);
nand U396 (N_396,In_1789,In_1333);
nand U397 (N_397,In_279,In_1133);
nor U398 (N_398,In_276,In_883);
xnor U399 (N_399,In_1416,In_798);
nand U400 (N_400,In_1399,N_358);
xor U401 (N_401,N_143,In_1784);
nand U402 (N_402,N_344,In_621);
or U403 (N_403,In_210,In_1696);
and U404 (N_404,N_13,In_1104);
and U405 (N_405,In_1556,In_1078);
and U406 (N_406,In_177,In_1197);
nand U407 (N_407,In_1363,In_1325);
xor U408 (N_408,In_522,In_1163);
xnor U409 (N_409,In_1534,In_915);
nand U410 (N_410,In_1430,In_1129);
xor U411 (N_411,N_204,In_235);
or U412 (N_412,In_990,In_699);
xnor U413 (N_413,In_787,In_1386);
nor U414 (N_414,In_1435,N_229);
nand U415 (N_415,In_109,In_554);
xnor U416 (N_416,In_27,In_108);
nand U417 (N_417,N_206,In_585);
and U418 (N_418,In_306,In_1847);
nand U419 (N_419,In_595,N_233);
and U420 (N_420,In_1316,In_1613);
xnor U421 (N_421,In_22,In_626);
nor U422 (N_422,In_1987,In_1569);
nor U423 (N_423,N_242,In_1583);
xnor U424 (N_424,In_1870,N_125);
nand U425 (N_425,In_117,In_46);
nand U426 (N_426,In_501,N_222);
nand U427 (N_427,In_1633,In_947);
or U428 (N_428,N_217,In_414);
xor U429 (N_429,N_212,In_805);
or U430 (N_430,N_215,In_311);
and U431 (N_431,In_885,In_1214);
nor U432 (N_432,In_519,In_1712);
and U433 (N_433,In_875,In_249);
nor U434 (N_434,N_5,N_368);
or U435 (N_435,In_87,In_775);
nor U436 (N_436,In_749,N_36);
nor U437 (N_437,N_196,In_869);
nand U438 (N_438,In_1841,N_210);
or U439 (N_439,N_178,In_1140);
and U440 (N_440,In_1622,In_451);
and U441 (N_441,In_907,In_1213);
or U442 (N_442,In_761,In_460);
nand U443 (N_443,In_722,In_1146);
or U444 (N_444,In_992,In_154);
or U445 (N_445,N_145,In_64);
or U446 (N_446,In_669,In_196);
xor U447 (N_447,N_320,N_12);
nand U448 (N_448,In_61,N_188);
nand U449 (N_449,N_237,In_1994);
nand U450 (N_450,In_388,N_235);
or U451 (N_451,In_1574,In_1975);
and U452 (N_452,In_1100,In_141);
and U453 (N_453,N_124,In_1162);
or U454 (N_454,In_988,N_275);
nand U455 (N_455,N_68,In_658);
or U456 (N_456,In_454,N_2);
nor U457 (N_457,In_468,In_780);
nor U458 (N_458,In_1950,In_1857);
or U459 (N_459,In_1921,In_112);
nor U460 (N_460,In_63,In_1382);
nor U461 (N_461,In_1637,In_1016);
xor U462 (N_462,In_1813,N_132);
nand U463 (N_463,In_48,In_528);
nor U464 (N_464,N_397,In_1125);
nand U465 (N_465,In_512,N_158);
or U466 (N_466,In_1631,N_243);
nand U467 (N_467,N_246,In_737);
nand U468 (N_468,In_1185,In_1066);
or U469 (N_469,N_153,In_784);
and U470 (N_470,In_208,In_313);
or U471 (N_471,In_1404,N_174);
and U472 (N_472,In_797,In_217);
nand U473 (N_473,In_668,In_855);
and U474 (N_474,In_1755,In_1169);
xnor U475 (N_475,In_879,In_73);
and U476 (N_476,In_866,In_1292);
nor U477 (N_477,In_110,N_234);
or U478 (N_478,In_1852,In_312);
nor U479 (N_479,N_219,In_1240);
nor U480 (N_480,In_1276,In_1393);
or U481 (N_481,In_1988,N_388);
and U482 (N_482,In_894,N_35);
nand U483 (N_483,N_272,In_419);
nand U484 (N_484,In_573,In_503);
nand U485 (N_485,In_1183,In_560);
nor U486 (N_486,In_1178,N_106);
xnor U487 (N_487,In_1189,In_1629);
nand U488 (N_488,In_1097,In_1677);
nor U489 (N_489,In_432,In_60);
and U490 (N_490,In_1101,In_1176);
nand U491 (N_491,In_1909,In_1578);
and U492 (N_492,N_49,N_342);
nor U493 (N_493,In_1920,In_395);
nand U494 (N_494,In_147,In_996);
xnor U495 (N_495,In_1906,N_61);
and U496 (N_496,In_1179,In_264);
or U497 (N_497,In_1277,In_456);
nand U498 (N_498,In_1628,N_87);
nor U499 (N_499,In_1585,In_1391);
and U500 (N_500,N_159,N_67);
and U501 (N_501,N_323,N_302);
nand U502 (N_502,In_1760,In_490);
or U503 (N_503,In_1029,N_144);
xnor U504 (N_504,In_677,N_346);
nor U505 (N_505,In_1926,In_976);
nand U506 (N_506,In_1792,N_269);
and U507 (N_507,In_789,In_1497);
and U508 (N_508,N_352,In_1758);
or U509 (N_509,N_288,In_1707);
or U510 (N_510,In_783,In_1051);
nand U511 (N_511,In_178,In_551);
nand U512 (N_512,In_1662,In_1079);
nand U513 (N_513,N_102,In_1808);
or U514 (N_514,In_1000,In_724);
nand U515 (N_515,N_110,In_747);
and U516 (N_516,N_384,N_250);
xor U517 (N_517,In_1293,In_1352);
nand U518 (N_518,N_189,In_376);
and U519 (N_519,In_1887,In_1479);
and U520 (N_520,In_1934,N_83);
xnor U521 (N_521,In_498,In_1145);
nor U522 (N_522,In_385,N_252);
and U523 (N_523,In_1883,N_297);
or U524 (N_524,In_1298,In_1453);
nand U525 (N_525,In_736,In_795);
or U526 (N_526,In_1690,In_1575);
nor U527 (N_527,In_1937,In_1192);
nand U528 (N_528,In_1968,In_1360);
nand U529 (N_529,In_1354,In_1268);
and U530 (N_530,In_1334,In_861);
nor U531 (N_531,N_111,In_286);
and U532 (N_532,In_541,In_1697);
xor U533 (N_533,In_508,In_315);
and U534 (N_534,N_396,In_1491);
xor U535 (N_535,In_239,In_1607);
nor U536 (N_536,In_1309,In_91);
nor U537 (N_537,In_1050,In_1954);
nor U538 (N_538,In_1581,N_199);
and U539 (N_539,In_1499,In_1782);
nand U540 (N_540,N_54,In_1489);
xor U541 (N_541,In_97,N_322);
or U542 (N_542,In_415,In_1731);
or U543 (N_543,N_371,In_142);
nor U544 (N_544,In_622,In_364);
and U545 (N_545,In_102,In_1267);
and U546 (N_546,In_1408,In_833);
nor U547 (N_547,N_301,In_891);
nor U548 (N_548,In_1636,In_1068);
or U549 (N_549,In_269,In_1522);
or U550 (N_550,In_1082,N_184);
and U551 (N_551,In_810,In_935);
nand U552 (N_552,In_1414,In_701);
nand U553 (N_553,N_361,N_249);
nor U554 (N_554,In_533,In_608);
nand U555 (N_555,In_383,N_126);
and U556 (N_556,In_815,In_172);
nand U557 (N_557,In_1681,In_1828);
and U558 (N_558,N_340,In_230);
nand U559 (N_559,In_1253,In_351);
or U560 (N_560,In_1273,In_1904);
and U561 (N_561,In_1510,In_101);
or U562 (N_562,In_295,In_148);
nor U563 (N_563,In_384,N_1);
or U564 (N_564,In_1330,N_218);
nor U565 (N_565,In_41,N_65);
or U566 (N_566,N_202,In_150);
nand U567 (N_567,N_45,In_143);
nand U568 (N_568,In_1494,N_90);
or U569 (N_569,In_325,In_1924);
nand U570 (N_570,In_1723,In_1366);
and U571 (N_571,In_118,N_27);
or U572 (N_572,In_1766,In_209);
nand U573 (N_573,N_387,In_1931);
and U574 (N_574,In_1640,N_334);
nor U575 (N_575,In_284,In_19);
or U576 (N_576,In_1126,In_1327);
or U577 (N_577,In_475,In_1951);
nor U578 (N_578,In_1304,In_969);
or U579 (N_579,In_1871,In_1465);
xor U580 (N_580,In_1933,In_107);
or U581 (N_581,N_389,In_1542);
or U582 (N_582,In_38,N_282);
xnor U583 (N_583,In_752,N_382);
or U584 (N_584,N_205,In_1908);
or U585 (N_585,In_1033,In_424);
and U586 (N_586,In_158,In_1970);
nand U587 (N_587,N_283,In_1802);
nand U588 (N_588,In_659,In_1544);
and U589 (N_589,N_0,In_1959);
nor U590 (N_590,In_1998,N_123);
and U591 (N_591,In_180,In_1874);
xnor U592 (N_592,N_84,N_34);
nor U593 (N_593,In_760,N_70);
nor U594 (N_594,N_325,In_1122);
and U595 (N_595,In_462,In_857);
and U596 (N_596,N_316,N_353);
nor U597 (N_597,In_1919,In_1830);
and U598 (N_598,N_308,N_117);
nand U599 (N_599,N_268,In_834);
nand U600 (N_600,In_1945,In_273);
nand U601 (N_601,In_920,N_4);
nor U602 (N_602,N_367,In_831);
nand U603 (N_603,In_827,In_1910);
and U604 (N_604,In_1361,In_1625);
and U605 (N_605,In_1191,In_1321);
or U606 (N_606,In_1339,In_566);
or U607 (N_607,In_998,In_1529);
or U608 (N_608,In_1537,N_214);
or U609 (N_609,In_1535,N_228);
nor U610 (N_610,In_359,N_133);
and U611 (N_611,N_239,In_1872);
nor U612 (N_612,N_24,In_521);
nor U613 (N_613,In_1606,In_1195);
nor U614 (N_614,In_720,In_66);
or U615 (N_615,In_185,In_259);
xor U616 (N_616,In_155,In_67);
and U617 (N_617,In_1827,In_228);
nand U618 (N_618,In_1443,In_258);
and U619 (N_619,In_1922,In_712);
and U620 (N_620,In_348,In_404);
nand U621 (N_621,In_1565,In_1107);
or U622 (N_622,In_377,In_1468);
or U623 (N_623,N_94,N_134);
nor U624 (N_624,In_548,N_52);
nor U625 (N_625,In_1539,N_162);
xor U626 (N_626,N_339,N_195);
nor U627 (N_627,N_20,In_1993);
or U628 (N_628,In_176,In_779);
xor U629 (N_629,N_163,In_1252);
nor U630 (N_630,In_1207,In_1925);
xor U631 (N_631,N_277,N_171);
or U632 (N_632,N_377,In_586);
nand U633 (N_633,In_1139,In_556);
and U634 (N_634,N_309,N_37);
xnor U635 (N_635,N_50,In_607);
or U636 (N_636,N_224,N_72);
nor U637 (N_637,In_1406,In_1109);
and U638 (N_638,In_569,In_1781);
or U639 (N_639,In_657,In_695);
nand U640 (N_640,N_185,In_1398);
nand U641 (N_641,In_1004,N_292);
xor U642 (N_642,In_1039,N_136);
xnor U643 (N_643,In_614,In_431);
xnor U644 (N_644,N_303,In_648);
xnor U645 (N_645,In_1698,In_1780);
nand U646 (N_646,N_262,In_581);
xor U647 (N_647,In_623,In_510);
xor U648 (N_648,In_226,In_562);
nand U649 (N_649,N_293,N_348);
xnor U650 (N_650,In_222,N_22);
nor U651 (N_651,In_1582,In_598);
nand U652 (N_652,In_820,In_1563);
nand U653 (N_653,In_1070,In_71);
nand U654 (N_654,In_1130,In_750);
or U655 (N_655,In_1757,In_536);
nor U656 (N_656,In_618,N_241);
and U657 (N_657,In_254,In_492);
or U658 (N_658,In_878,N_129);
nand U659 (N_659,N_394,In_1543);
xnor U660 (N_660,In_1868,In_305);
nand U661 (N_661,In_1446,In_1093);
nor U662 (N_662,N_75,In_1045);
nand U663 (N_663,N_107,In_144);
nor U664 (N_664,In_1501,In_229);
nand U665 (N_665,In_441,N_81);
nor U666 (N_666,N_326,N_265);
or U667 (N_667,In_1091,In_832);
nor U668 (N_668,N_370,In_790);
or U669 (N_669,In_435,In_444);
and U670 (N_670,In_51,In_1166);
and U671 (N_671,In_175,In_36);
and U672 (N_672,In_371,In_1840);
nand U673 (N_673,In_35,In_888);
nor U674 (N_674,N_177,N_286);
nor U675 (N_675,In_467,In_1329);
and U676 (N_676,In_277,N_91);
xnor U677 (N_677,In_1288,In_1466);
and U678 (N_678,In_662,In_1160);
and U679 (N_679,In_0,In_1620);
nand U680 (N_680,In_925,In_1052);
nor U681 (N_681,N_236,In_1271);
nor U682 (N_682,In_872,In_203);
nor U683 (N_683,In_1442,In_1187);
or U684 (N_684,In_1461,In_1685);
and U685 (N_685,In_1359,In_1302);
or U686 (N_686,In_860,N_335);
xor U687 (N_687,In_944,N_99);
xor U688 (N_688,In_1429,In_1915);
or U689 (N_689,In_723,N_137);
xnor U690 (N_690,N_357,In_717);
and U691 (N_691,In_1198,In_1810);
xor U692 (N_692,N_170,In_877);
and U693 (N_693,N_66,In_245);
or U694 (N_694,In_201,In_10);
nor U695 (N_695,In_1154,In_673);
or U696 (N_696,In_1599,In_160);
xor U697 (N_697,In_1669,In_1076);
or U698 (N_698,N_284,In_132);
xnor U699 (N_699,N_381,In_267);
or U700 (N_700,In_310,In_1831);
nor U701 (N_701,In_1967,In_1939);
nor U702 (N_702,N_393,In_1284);
and U703 (N_703,In_316,N_317);
or U704 (N_704,In_1822,N_191);
xnor U705 (N_705,In_81,In_1719);
nand U706 (N_706,In_1155,In_1032);
xnor U707 (N_707,In_999,In_850);
and U708 (N_708,In_1750,In_1027);
nand U709 (N_709,In_1009,In_411);
xnor U710 (N_710,In_649,In_1745);
or U711 (N_711,In_1788,In_953);
and U712 (N_712,In_1675,In_927);
or U713 (N_713,In_1700,N_43);
nand U714 (N_714,In_1590,In_1514);
nand U715 (N_715,In_122,In_960);
xor U716 (N_716,In_697,In_676);
xnor U717 (N_717,In_1554,In_1202);
and U718 (N_718,In_1370,In_1891);
nor U719 (N_719,In_1907,In_1749);
and U720 (N_720,In_1225,N_32);
nand U721 (N_721,N_167,In_811);
and U722 (N_722,In_1894,In_1779);
nor U723 (N_723,In_1787,In_1761);
nand U724 (N_724,In_984,In_838);
and U725 (N_725,In_847,In_1095);
and U726 (N_726,In_1260,N_349);
and U727 (N_727,In_773,In_1017);
and U728 (N_728,In_552,In_954);
nand U729 (N_729,In_1630,In_1324);
and U730 (N_730,In_1229,N_63);
nand U731 (N_731,In_1743,N_386);
nor U732 (N_732,In_873,In_1283);
nor U733 (N_733,N_330,In_584);
or U734 (N_734,In_606,N_121);
nand U735 (N_735,In_1269,N_115);
nand U736 (N_736,In_335,In_1948);
nor U737 (N_737,In_755,N_255);
or U738 (N_738,N_363,N_337);
or U739 (N_739,In_1059,In_936);
and U740 (N_740,In_754,In_1733);
or U741 (N_741,N_294,In_293);
and U742 (N_742,In_1021,In_706);
xnor U743 (N_743,In_1134,In_771);
or U744 (N_744,N_372,N_208);
nor U745 (N_745,N_360,N_324);
and U746 (N_746,In_1572,N_160);
xor U747 (N_747,In_793,In_1174);
and U748 (N_748,In_1506,In_1699);
and U749 (N_749,In_78,N_276);
and U750 (N_750,In_1974,In_323);
and U751 (N_751,In_707,In_1963);
or U752 (N_752,In_693,In_685);
and U753 (N_753,In_762,In_688);
nand U754 (N_754,In_590,In_1701);
nand U755 (N_755,In_1962,In_665);
nor U756 (N_756,N_221,In_603);
or U757 (N_757,N_19,In_1103);
nand U758 (N_758,N_141,N_179);
xor U759 (N_759,N_364,In_49);
or U760 (N_760,N_299,In_978);
nand U761 (N_761,In_1215,In_252);
or U762 (N_762,In_1969,In_653);
and U763 (N_763,In_1694,In_250);
or U764 (N_764,In_1642,N_46);
and U765 (N_765,In_1977,In_1736);
and U766 (N_766,In_495,In_1600);
or U767 (N_767,In_1981,In_1262);
nand U768 (N_768,In_746,In_1123);
nand U769 (N_769,In_21,In_829);
nor U770 (N_770,N_101,In_1072);
xnor U771 (N_771,In_354,In_292);
and U772 (N_772,In_1752,In_640);
nor U773 (N_773,In_1597,In_709);
or U774 (N_774,In_375,N_93);
nor U775 (N_775,In_218,N_8);
nor U776 (N_776,In_1557,In_930);
nor U777 (N_777,In_1233,In_1168);
or U778 (N_778,In_28,In_1843);
nand U779 (N_779,N_114,In_1379);
and U780 (N_780,In_458,In_949);
and U781 (N_781,In_922,N_148);
nor U782 (N_782,In_33,In_664);
xor U783 (N_783,In_1684,N_310);
xnor U784 (N_784,In_76,In_1128);
or U785 (N_785,In_342,N_347);
and U786 (N_786,N_258,N_259);
and U787 (N_787,In_449,In_1538);
and U788 (N_788,In_484,In_187);
nand U789 (N_789,In_918,In_8);
and U790 (N_790,In_1702,In_1905);
nor U791 (N_791,In_660,In_1655);
nand U792 (N_792,N_383,In_1200);
or U793 (N_793,N_29,In_837);
and U794 (N_794,In_130,In_941);
or U795 (N_795,In_100,In_1094);
xor U796 (N_796,In_317,In_1279);
nor U797 (N_797,In_524,In_1652);
nand U798 (N_798,N_392,In_159);
nand U799 (N_799,In_466,In_1331);
nand U800 (N_800,N_720,In_523);
and U801 (N_801,N_686,N_534);
nor U802 (N_802,N_327,N_527);
or U803 (N_803,N_714,In_346);
xor U804 (N_804,N_745,In_1482);
nand U805 (N_805,N_580,N_742);
and U806 (N_806,N_548,In_515);
nand U807 (N_807,In_502,N_157);
or U808 (N_808,N_355,In_1460);
nor U809 (N_809,N_571,N_662);
or U810 (N_810,N_155,In_473);
and U811 (N_811,N_223,N_227);
and U812 (N_812,N_456,N_118);
and U813 (N_813,In_1037,In_981);
xor U814 (N_814,N_405,N_425);
and U815 (N_815,N_567,In_1340);
and U816 (N_816,In_1188,N_427);
and U817 (N_817,In_1244,N_176);
or U818 (N_818,N_120,In_1136);
and U819 (N_819,N_664,N_260);
nor U820 (N_820,N_560,N_271);
nor U821 (N_821,N_207,N_640);
nor U822 (N_822,N_577,N_7);
and U823 (N_823,In_1439,In_822);
nor U824 (N_824,N_616,In_1682);
xnor U825 (N_825,N_165,In_1550);
or U826 (N_826,N_407,In_1236);
and U827 (N_827,N_267,N_95);
or U828 (N_828,In_1259,N_748);
nor U829 (N_829,N_703,N_569);
nand U830 (N_830,N_216,N_558);
nor U831 (N_831,N_274,N_590);
or U832 (N_832,In_663,In_890);
nand U833 (N_833,N_51,N_541);
nor U834 (N_834,N_89,N_417);
nand U835 (N_835,In_530,N_775);
nand U836 (N_836,In_1979,N_182);
nor U837 (N_837,In_223,In_410);
nor U838 (N_838,N_575,In_1058);
or U839 (N_839,In_88,In_1367);
nor U840 (N_840,In_1643,N_477);
and U841 (N_841,N_792,In_1686);
nand U842 (N_842,In_365,In_1742);
or U843 (N_843,N_203,N_333);
xnor U844 (N_844,N_418,In_1265);
nand U845 (N_845,In_1450,In_686);
or U846 (N_846,N_365,N_98);
nor U847 (N_847,In_1709,N_671);
xor U848 (N_848,In_1732,In_189);
nor U849 (N_849,In_1741,In_1454);
xnor U850 (N_850,N_47,In_341);
or U851 (N_851,N_298,N_92);
nand U852 (N_852,N_147,N_3);
nor U853 (N_853,N_149,N_247);
nor U854 (N_854,N_669,In_1358);
xor U855 (N_855,In_129,In_332);
or U856 (N_856,N_404,N_192);
nand U857 (N_857,N_231,N_401);
nand U858 (N_858,In_1180,N_109);
and U859 (N_859,N_506,In_265);
nor U860 (N_860,In_360,In_1493);
and U861 (N_861,N_62,N_463);
nand U862 (N_862,In_1485,In_283);
or U863 (N_863,N_402,In_1848);
xnor U864 (N_864,In_770,N_266);
xnor U865 (N_865,N_790,In_768);
nand U866 (N_866,N_770,In_921);
or U867 (N_867,N_794,N_173);
and U868 (N_868,In_1326,In_1515);
and U869 (N_869,N_369,N_305);
and U870 (N_870,N_668,In_1371);
nor U871 (N_871,N_650,N_416);
nand U872 (N_872,N_306,N_706);
and U873 (N_873,N_476,N_747);
nand U874 (N_874,N_778,In_1057);
and U875 (N_875,In_1291,In_1595);
and U876 (N_876,N_380,In_1820);
xnor U877 (N_877,In_589,N_354);
nor U878 (N_878,N_660,In_1986);
or U879 (N_879,In_568,In_1641);
nand U880 (N_880,N_731,In_1356);
and U881 (N_881,In_788,N_69);
nand U882 (N_882,In_782,In_619);
nand U883 (N_883,In_641,In_489);
and U884 (N_884,N_673,N_688);
and U885 (N_885,In_1250,In_504);
xnor U886 (N_886,In_1064,N_116);
or U887 (N_887,N_700,In_1842);
nand U888 (N_888,In_638,N_281);
nor U889 (N_889,N_619,N_586);
xnor U890 (N_890,N_257,N_435);
nand U891 (N_891,In_751,N_679);
and U892 (N_892,In_138,N_643);
or U893 (N_893,In_550,In_358);
nor U894 (N_894,In_1594,In_1201);
and U895 (N_895,N_798,In_611);
or U896 (N_896,N_783,N_760);
nor U897 (N_897,In_631,In_1611);
or U898 (N_898,In_1814,N_491);
nand U899 (N_899,N_452,N_359);
and U900 (N_900,In_1390,N_683);
xor U901 (N_901,N_79,In_1528);
xor U902 (N_902,N_728,N_493);
nor U903 (N_903,In_44,N_180);
nor U904 (N_904,In_379,In_774);
xnor U905 (N_905,N_403,In_1823);
and U906 (N_906,In_955,N_385);
and U907 (N_907,N_475,N_433);
or U908 (N_908,N_723,N_540);
xor U909 (N_909,In_576,N_749);
nand U910 (N_910,In_1433,In_1417);
nand U911 (N_911,N_18,In_767);
nor U912 (N_912,N_535,In_1478);
or U913 (N_913,In_889,In_197);
and U914 (N_914,N_759,N_736);
and U915 (N_915,N_56,N_716);
and U916 (N_916,N_727,In_1564);
xor U917 (N_917,In_1893,In_1687);
xor U918 (N_918,In_1504,In_1148);
nand U919 (N_919,N_374,In_120);
xor U920 (N_920,N_6,In_870);
or U921 (N_921,N_119,N_543);
and U922 (N_922,In_1984,N_413);
or U923 (N_923,N_240,In_1658);
or U924 (N_924,In_392,N_395);
nor U925 (N_925,In_1829,In_1957);
nand U926 (N_926,N_366,In_813);
nand U927 (N_927,N_645,In_1955);
nand U928 (N_928,N_345,In_86);
and U929 (N_929,N_434,N_496);
nand U930 (N_930,N_270,N_429);
nor U931 (N_931,N_568,N_724);
nand U932 (N_932,N_28,In_1158);
nor U933 (N_933,N_538,N_694);
or U934 (N_934,N_787,N_251);
or U935 (N_935,N_423,In_1663);
nor U936 (N_936,N_722,In_645);
nor U937 (N_937,In_319,N_140);
or U938 (N_938,In_31,In_1902);
nand U939 (N_939,In_485,In_549);
xnor U940 (N_940,In_211,N_633);
and U941 (N_941,In_1989,N_691);
nand U942 (N_942,In_45,In_1571);
nor U943 (N_943,In_983,N_139);
nor U944 (N_944,In_247,N_626);
nor U945 (N_945,N_530,In_1710);
nor U946 (N_946,In_438,N_515);
or U947 (N_947,N_419,In_1046);
nand U948 (N_948,In_408,In_545);
nor U949 (N_949,In_1199,In_1536);
or U950 (N_950,N_398,In_1520);
nor U951 (N_951,In_83,N_638);
nor U952 (N_952,In_1656,N_200);
and U953 (N_953,In_577,In_647);
or U954 (N_954,N_458,N_528);
nand U955 (N_955,N_629,In_1526);
nor U956 (N_956,N_647,N_786);
or U957 (N_957,In_1026,N_168);
xnor U958 (N_958,In_579,In_307);
nor U959 (N_959,In_702,N_85);
and U960 (N_960,N_484,In_1672);
and U961 (N_961,N_750,N_701);
or U962 (N_962,N_753,N_78);
nand U963 (N_963,N_112,N_410);
and U964 (N_964,N_597,In_615);
and U965 (N_965,N_44,N_409);
and U966 (N_966,N_651,N_646);
nand U967 (N_967,In_1896,N_667);
nor U968 (N_968,In_1715,In_588);
nand U969 (N_969,N_127,In_74);
nand U970 (N_970,N_156,N_279);
nand U971 (N_971,In_1768,N_744);
and U972 (N_972,In_1384,N_594);
nor U973 (N_973,In_308,N_244);
or U974 (N_974,In_1055,In_1502);
or U975 (N_975,N_555,In_995);
and U976 (N_976,N_482,In_93);
xnor U977 (N_977,In_1531,N_627);
and U978 (N_978,N_473,N_245);
or U979 (N_979,In_1776,N_80);
nor U980 (N_980,N_104,N_319);
or U981 (N_981,N_97,N_554);
nand U982 (N_982,In_1473,N_539);
nor U983 (N_983,In_1328,In_1472);
xnor U984 (N_984,N_307,N_767);
nor U985 (N_985,N_332,In_1527);
or U986 (N_986,In_24,N_261);
xnor U987 (N_987,In_1618,In_1889);
nor U988 (N_988,N_25,In_1227);
and U989 (N_989,N_725,In_527);
and U990 (N_990,In_423,In_1062);
nand U991 (N_991,N_642,In_1566);
xor U992 (N_992,In_1729,N_30);
or U993 (N_993,N_411,In_125);
or U994 (N_994,In_704,N_287);
nor U995 (N_995,In_476,N_142);
and U996 (N_996,N_547,N_479);
or U997 (N_997,N_451,N_776);
nand U998 (N_998,In_1441,N_489);
xnor U999 (N_999,In_195,N_754);
nor U1000 (N_1000,In_320,In_14);
nor U1001 (N_1001,N_296,In_1772);
nand U1002 (N_1002,N_454,N_225);
nand U1003 (N_1003,In_1475,In_1816);
and U1004 (N_1004,N_130,In_1320);
nand U1005 (N_1005,In_975,In_59);
nor U1006 (N_1006,N_755,In_378);
or U1007 (N_1007,In_1096,N_523);
nor U1008 (N_1008,In_443,N_608);
nor U1009 (N_1009,N_278,N_9);
and U1010 (N_1010,In_715,N_620);
or U1011 (N_1011,N_467,In_1638);
or U1012 (N_1012,In_1615,N_634);
or U1013 (N_1013,N_248,N_441);
and U1014 (N_1014,In_382,In_1825);
nor U1015 (N_1015,In_18,N_280);
nor U1016 (N_1016,In_814,N_376);
xnor U1017 (N_1017,In_1396,N_752);
nand U1018 (N_1018,N_552,N_438);
nand U1019 (N_1019,N_485,In_1793);
nand U1020 (N_1020,In_1407,N_161);
xnor U1021 (N_1021,In_433,N_58);
or U1022 (N_1022,In_162,In_52);
xor U1023 (N_1023,In_1725,In_487);
nand U1024 (N_1024,In_1791,N_338);
nor U1025 (N_1025,N_693,In_1005);
nor U1026 (N_1026,N_687,In_1785);
and U1027 (N_1027,N_593,N_655);
or U1028 (N_1028,N_730,In_124);
nor U1029 (N_1029,In_1182,N_644);
and U1030 (N_1030,In_304,N_77);
nand U1031 (N_1031,N_312,N_625);
and U1032 (N_1032,N_64,In_366);
nor U1033 (N_1033,N_583,In_719);
nand U1034 (N_1034,In_137,In_352);
nand U1035 (N_1035,N_682,In_450);
or U1036 (N_1036,In_698,In_803);
nand U1037 (N_1037,N_211,In_1879);
nand U1038 (N_1038,In_240,N_735);
and U1039 (N_1039,In_1960,In_1138);
nand U1040 (N_1040,In_591,In_1278);
xor U1041 (N_1041,In_393,N_661);
nor U1042 (N_1042,In_1996,N_582);
or U1043 (N_1043,In_253,N_505);
xnor U1044 (N_1044,N_793,In_886);
xor U1045 (N_1045,N_737,In_1343);
nor U1046 (N_1046,In_632,In_167);
nor U1047 (N_1047,In_17,In_1011);
or U1048 (N_1048,In_1819,In_161);
nor U1049 (N_1049,In_691,In_635);
or U1050 (N_1050,In_1345,N_400);
xor U1051 (N_1051,N_588,N_412);
or U1052 (N_1052,N_88,N_445);
xnor U1053 (N_1053,N_578,N_378);
nor U1054 (N_1054,In_437,N_391);
nand U1055 (N_1055,In_1372,In_1495);
or U1056 (N_1056,In_1084,N_331);
nand U1057 (N_1057,N_612,In_1573);
xnor U1058 (N_1058,In_227,In_1932);
nor U1059 (N_1059,In_1226,N_304);
nand U1060 (N_1060,In_439,N_631);
nor U1061 (N_1061,N_596,N_665);
nor U1062 (N_1062,N_677,In_973);
and U1063 (N_1063,N_73,In_599);
or U1064 (N_1064,In_396,In_661);
and U1065 (N_1065,In_39,N_295);
or U1066 (N_1066,N_719,In_25);
nand U1067 (N_1067,In_948,In_1918);
nor U1068 (N_1068,N_526,N_41);
nor U1069 (N_1069,N_470,In_280);
and U1070 (N_1070,In_1073,In_1061);
or U1071 (N_1071,N_455,N_15);
nand U1072 (N_1072,In_1012,In_1853);
nand U1073 (N_1073,In_412,In_436);
or U1074 (N_1074,N_757,In_1437);
nand U1075 (N_1075,N_220,In_149);
and U1076 (N_1076,In_629,N_517);
xor U1077 (N_1077,In_1015,In_1194);
and U1078 (N_1078,In_1149,In_842);
and U1079 (N_1079,In_1243,In_741);
nand U1080 (N_1080,N_613,In_1422);
or U1081 (N_1081,N_678,In_1235);
and U1082 (N_1082,N_630,N_514);
nand U1083 (N_1083,In_1041,In_911);
and U1084 (N_1084,In_1275,N_498);
xnor U1085 (N_1085,N_510,In_417);
xor U1086 (N_1086,In_1251,In_309);
or U1087 (N_1087,In_563,In_1368);
or U1088 (N_1088,In_1935,N_421);
nor U1089 (N_1089,N_457,In_479);
and U1090 (N_1090,In_634,In_642);
and U1091 (N_1091,In_1548,N_733);
xnor U1092 (N_1092,In_405,In_1521);
nand U1093 (N_1093,N_238,N_453);
nor U1094 (N_1094,In_845,N_618);
nand U1095 (N_1095,N_264,In_1604);
nand U1096 (N_1096,In_880,N_313);
and U1097 (N_1097,N_740,N_289);
nand U1098 (N_1098,In_1744,N_636);
or U1099 (N_1099,N_772,N_799);
and U1100 (N_1100,In_952,N_273);
or U1101 (N_1101,N_784,N_623);
nand U1102 (N_1102,N_599,In_213);
nor U1103 (N_1103,In_1763,In_1392);
or U1104 (N_1104,In_718,N_321);
nand U1105 (N_1105,N_60,In_1724);
or U1106 (N_1106,In_486,In_1608);
nand U1107 (N_1107,N_172,In_628);
nand U1108 (N_1108,N_226,In_772);
or U1109 (N_1109,N_420,N_652);
nand U1110 (N_1110,In_1713,N_663);
nor U1111 (N_1111,N_551,N_96);
xor U1112 (N_1112,N_717,In_1239);
xnor U1113 (N_1113,N_190,In_1646);
nand U1114 (N_1114,N_589,N_771);
nand U1115 (N_1115,In_32,N_461);
and U1116 (N_1116,N_138,In_979);
xnor U1117 (N_1117,In_1124,In_908);
xnor U1118 (N_1118,N_641,N_708);
nand U1119 (N_1119,In_964,In_1508);
or U1120 (N_1120,In_271,N_676);
and U1121 (N_1121,N_587,In_1272);
xor U1122 (N_1122,N_584,N_718);
or U1123 (N_1123,In_369,N_533);
nand U1124 (N_1124,N_42,N_542);
nand U1125 (N_1125,N_573,N_544);
xor U1126 (N_1126,N_739,In_1668);
and U1127 (N_1127,In_1797,In_1018);
or U1128 (N_1128,In_1971,N_656);
or U1129 (N_1129,N_622,In_1596);
or U1130 (N_1130,N_426,In_1609);
and U1131 (N_1131,In_1400,N_711);
or U1132 (N_1132,N_617,N_702);
nand U1133 (N_1133,N_615,In_1773);
and U1134 (N_1134,N_574,N_488);
nand U1135 (N_1135,N_328,N_637);
nand U1136 (N_1136,In_3,In_493);
or U1137 (N_1137,N_576,N_193);
and U1138 (N_1138,In_1028,N_648);
xor U1139 (N_1139,In_1627,In_1246);
nand U1140 (N_1140,N_486,In_1591);
or U1141 (N_1141,N_713,In_785);
nor U1142 (N_1142,In_764,N_194);
xor U1143 (N_1143,N_290,N_670);
or U1144 (N_1144,In_275,In_1440);
nor U1145 (N_1145,In_1678,In_580);
nand U1146 (N_1146,N_572,N_406);
or U1147 (N_1147,N_565,N_186);
xnor U1148 (N_1148,N_14,N_495);
and U1149 (N_1149,In_505,In_430);
nand U1150 (N_1150,In_902,In_1053);
and U1151 (N_1151,In_1587,In_652);
nor U1152 (N_1152,N_379,N_483);
xor U1153 (N_1153,N_734,In_1577);
xor U1154 (N_1154,In_389,N_743);
nand U1155 (N_1155,In_1913,In_578);
or U1156 (N_1156,N_761,In_900);
xnor U1157 (N_1157,In_200,N_300);
and U1158 (N_1158,N_462,N_82);
nor U1159 (N_1159,In_1190,N_518);
nor U1160 (N_1160,In_511,In_1085);
and U1161 (N_1161,N_490,N_442);
or U1162 (N_1162,N_756,In_1081);
nor U1163 (N_1163,N_256,In_238);
or U1164 (N_1164,N_785,In_263);
and U1165 (N_1165,N_253,In_338);
nor U1166 (N_1166,N_666,In_1867);
and U1167 (N_1167,N_697,In_1151);
nand U1168 (N_1168,N_628,In_399);
nand U1169 (N_1169,In_1770,In_1805);
nand U1170 (N_1170,N_632,In_520);
xnor U1171 (N_1171,N_469,In_971);
or U1172 (N_1172,N_356,N_524);
nand U1173 (N_1173,In_1409,In_903);
and U1174 (N_1174,N_213,N_675);
nor U1175 (N_1175,In_77,N_390);
nor U1176 (N_1176,N_796,In_7);
or U1177 (N_1177,N_672,In_478);
nor U1178 (N_1178,N_497,N_424);
and U1179 (N_1179,In_1172,N_698);
nand U1180 (N_1180,In_932,In_497);
xor U1181 (N_1181,In_1817,N_152);
and U1182 (N_1182,N_773,N_26);
and U1183 (N_1183,N_154,In_730);
nor U1184 (N_1184,In_561,N_546);
nand U1185 (N_1185,N_689,In_1965);
and U1186 (N_1186,N_55,In_514);
or U1187 (N_1187,N_710,In_1216);
or U1188 (N_1188,In_1222,N_658);
and U1189 (N_1189,N_492,In_1676);
nand U1190 (N_1190,In_68,N_183);
xor U1191 (N_1191,In_758,N_21);
and U1192 (N_1192,N_314,In_480);
nor U1193 (N_1193,In_794,In_862);
xor U1194 (N_1194,In_1286,In_1983);
or U1195 (N_1195,In_600,N_570);
nand U1196 (N_1196,In_1280,N_151);
or U1197 (N_1197,In_43,In_1452);
xor U1198 (N_1198,N_38,In_1294);
nor U1199 (N_1199,N_692,In_1691);
nand U1200 (N_1200,N_997,N_881);
xor U1201 (N_1201,N_1132,In_1487);
and U1202 (N_1202,N_955,In_1357);
nor U1203 (N_1203,N_765,N_1169);
and U1204 (N_1204,N_1172,N_817);
and U1205 (N_1205,N_864,N_1099);
xor U1206 (N_1206,N_811,N_850);
nand U1207 (N_1207,N_851,In_966);
xnor U1208 (N_1208,N_910,N_649);
xnor U1209 (N_1209,N_1005,N_842);
nor U1210 (N_1210,In_778,In_1568);
xnor U1211 (N_1211,N_621,In_1890);
or U1212 (N_1212,N_503,N_128);
and U1213 (N_1213,N_685,In_472);
or U1214 (N_1214,In_769,In_808);
or U1215 (N_1215,N_595,N_925);
and U1216 (N_1216,N_865,N_1146);
and U1217 (N_1217,N_1123,In_1311);
nand U1218 (N_1218,N_603,In_65);
nand U1219 (N_1219,In_1916,In_1310);
or U1220 (N_1220,N_820,N_1142);
or U1221 (N_1221,N_566,N_885);
and U1222 (N_1222,N_1092,N_520);
xor U1223 (N_1223,N_1156,N_1010);
or U1224 (N_1224,N_466,N_1018);
xor U1225 (N_1225,N_909,N_443);
and U1226 (N_1226,N_819,N_444);
nand U1227 (N_1227,N_408,In_1547);
nor U1228 (N_1228,N_1152,In_1858);
and U1229 (N_1229,In_469,N_1014);
or U1230 (N_1230,N_150,N_553);
or U1231 (N_1231,N_870,N_521);
xnor U1232 (N_1232,N_1098,N_841);
nand U1233 (N_1233,N_39,N_1042);
nand U1234 (N_1234,N_902,N_1175);
or U1235 (N_1235,N_1177,N_831);
xnor U1236 (N_1236,N_1120,In_1811);
and U1237 (N_1237,N_624,N_911);
nand U1238 (N_1238,N_1199,In_206);
nor U1239 (N_1239,N_977,In_865);
or U1240 (N_1240,N_695,N_906);
xor U1241 (N_1241,In_420,In_1897);
or U1242 (N_1242,N_797,N_465);
xnor U1243 (N_1243,N_919,N_336);
xnor U1244 (N_1244,N_1102,In_220);
nand U1245 (N_1245,In_745,N_53);
nand U1246 (N_1246,N_874,In_136);
nor U1247 (N_1247,In_1692,N_537);
and U1248 (N_1248,N_812,N_741);
nor U1249 (N_1249,In_425,In_1080);
nand U1250 (N_1250,N_887,In_1688);
and U1251 (N_1251,N_879,N_1197);
nand U1252 (N_1252,N_949,In_1812);
or U1253 (N_1253,N_1007,N_1016);
nor U1254 (N_1254,N_965,N_886);
or U1255 (N_1255,N_614,In_1432);
or U1256 (N_1256,N_900,N_875);
nor U1257 (N_1257,N_653,N_782);
and U1258 (N_1258,N_896,N_164);
and U1259 (N_1259,In_876,N_904);
nor U1260 (N_1260,N_76,N_813);
nand U1261 (N_1261,N_769,N_892);
and U1262 (N_1262,N_839,N_1054);
and U1263 (N_1263,N_1151,N_974);
nor U1264 (N_1264,In_1424,In_956);
nor U1265 (N_1265,N_1067,N_854);
nand U1266 (N_1266,N_1166,N_460);
nor U1267 (N_1267,N_780,In_1147);
nand U1268 (N_1268,N_945,N_709);
and U1269 (N_1269,N_1101,In_1282);
nor U1270 (N_1270,In_1153,N_1047);
xnor U1271 (N_1271,In_1512,N_876);
nand U1272 (N_1272,In_1584,In_1484);
nor U1273 (N_1273,N_894,N_1052);
xnor U1274 (N_1274,N_592,In_543);
nand U1275 (N_1275,N_818,N_113);
nand U1276 (N_1276,In_1961,N_732);
or U1277 (N_1277,N_607,N_922);
and U1278 (N_1278,N_1012,N_1040);
or U1279 (N_1279,N_10,N_549);
nor U1280 (N_1280,N_23,In_1644);
nand U1281 (N_1281,N_729,N_779);
nor U1282 (N_1282,N_1073,In_1601);
or U1283 (N_1283,N_209,N_480);
xor U1284 (N_1284,N_918,N_511);
nand U1285 (N_1285,In_290,N_1097);
xor U1286 (N_1286,N_1159,N_311);
and U1287 (N_1287,N_862,N_1056);
nand U1288 (N_1288,N_814,N_715);
nand U1289 (N_1289,N_895,N_830);
nand U1290 (N_1290,N_964,N_992);
or U1291 (N_1291,N_1160,N_1195);
nand U1292 (N_1292,N_880,N_1060);
and U1293 (N_1293,In_300,N_1028);
xor U1294 (N_1294,N_916,N_789);
nor U1295 (N_1295,In_791,N_1031);
nand U1296 (N_1296,N_459,N_604);
nor U1297 (N_1297,N_849,In_1801);
xnor U1298 (N_1298,N_1112,In_1255);
or U1299 (N_1299,In_221,N_169);
nor U1300 (N_1300,N_1191,N_802);
xnor U1301 (N_1301,In_1127,N_1037);
xor U1302 (N_1302,N_912,N_175);
xor U1303 (N_1303,N_635,In_1942);
xnor U1304 (N_1304,N_559,N_1050);
or U1305 (N_1305,In_1307,N_351);
xor U1306 (N_1306,In_256,N_1189);
nor U1307 (N_1307,N_329,N_888);
or U1308 (N_1308,N_468,N_1011);
and U1309 (N_1309,N_838,N_956);
nand U1310 (N_1310,In_1256,N_940);
and U1311 (N_1311,N_986,N_958);
and U1312 (N_1312,N_801,In_564);
xnor U1313 (N_1313,N_826,N_1184);
nor U1314 (N_1314,N_1088,N_920);
xor U1315 (N_1315,In_1507,In_145);
nor U1316 (N_1316,N_1164,N_882);
or U1317 (N_1317,N_1017,N_254);
xnor U1318 (N_1318,In_422,N_1036);
nand U1319 (N_1319,N_699,In_518);
xor U1320 (N_1320,N_201,N_531);
nand U1321 (N_1321,N_996,In_1464);
xor U1322 (N_1322,N_821,In_1541);
xor U1323 (N_1323,In_151,In_72);
and U1324 (N_1324,N_696,N_913);
nand U1325 (N_1325,N_674,N_1162);
and U1326 (N_1326,In_347,In_734);
and U1327 (N_1327,N_832,N_1070);
and U1328 (N_1328,In_1795,N_993);
nand U1329 (N_1329,N_263,N_509);
nor U1330 (N_1330,N_987,N_861);
xnor U1331 (N_1331,N_1090,In_1186);
or U1332 (N_1332,N_501,In_1193);
and U1333 (N_1333,N_513,In_1947);
nor U1334 (N_1334,N_835,N_350);
or U1335 (N_1335,N_17,N_1178);
xor U1336 (N_1336,In_11,In_204);
nor U1337 (N_1337,In_134,In_1135);
nand U1338 (N_1338,N_933,In_553);
nand U1339 (N_1339,In_765,N_848);
or U1340 (N_1340,N_763,N_1062);
nand U1341 (N_1341,N_581,N_1026);
and U1342 (N_1342,N_857,N_478);
and U1343 (N_1343,In_1036,N_950);
nand U1344 (N_1344,N_11,In_1876);
nor U1345 (N_1345,In_1347,N_502);
xor U1346 (N_1346,N_1114,N_1126);
nand U1347 (N_1347,N_1105,In_357);
or U1348 (N_1348,N_901,N_705);
or U1349 (N_1349,N_908,N_970);
and U1350 (N_1350,In_1388,N_598);
xnor U1351 (N_1351,N_285,N_1034);
nor U1352 (N_1352,In_464,N_878);
nor U1353 (N_1353,N_1173,N_1004);
and U1354 (N_1354,N_1119,N_1168);
and U1355 (N_1355,N_437,N_1188);
xnor U1356 (N_1356,N_1121,N_1183);
nand U1357 (N_1357,N_939,N_606);
or U1358 (N_1358,In_350,In_743);
nor U1359 (N_1359,N_1187,In_152);
or U1360 (N_1360,N_721,In_1673);
and U1361 (N_1361,N_198,N_375);
nand U1362 (N_1362,N_1117,In_121);
nand U1363 (N_1363,N_1131,In_1751);
or U1364 (N_1364,N_991,In_261);
nand U1365 (N_1365,N_74,N_943);
and U1366 (N_1366,N_1024,N_988);
or U1367 (N_1367,N_957,N_1051);
and U1368 (N_1368,In_583,N_1025);
or U1369 (N_1369,N_40,In_55);
nor U1370 (N_1370,In_913,N_1193);
nand U1371 (N_1371,N_318,N_464);
nand U1372 (N_1372,In_1451,N_1138);
and U1373 (N_1373,N_450,N_654);
xnor U1374 (N_1374,In_744,N_758);
nor U1375 (N_1375,N_942,N_1167);
and U1376 (N_1376,N_815,N_1063);
or U1377 (N_1377,N_941,In_1650);
and U1378 (N_1378,N_746,N_808);
nor U1379 (N_1379,N_971,In_174);
xnor U1380 (N_1380,N_166,In_961);
and U1381 (N_1381,N_1104,N_825);
xor U1382 (N_1382,N_609,N_1076);
xor U1383 (N_1383,In_703,In_1231);
or U1384 (N_1384,N_579,In_184);
nor U1385 (N_1385,N_1049,N_422);
and U1386 (N_1386,N_822,N_439);
and U1387 (N_1387,In_1208,N_108);
and U1388 (N_1388,N_791,N_432);
nand U1389 (N_1389,N_1094,N_436);
xor U1390 (N_1390,N_1192,N_768);
or U1391 (N_1391,N_105,N_959);
nor U1392 (N_1392,N_545,N_872);
or U1393 (N_1393,N_1032,N_1100);
and U1394 (N_1394,N_499,N_1078);
nor U1395 (N_1395,N_1041,N_834);
nor U1396 (N_1396,In_1553,N_1161);
and U1397 (N_1397,N_1150,N_982);
or U1398 (N_1398,N_1174,N_1030);
nor U1399 (N_1399,N_487,N_928);
nor U1400 (N_1400,N_187,In_710);
or U1401 (N_1401,N_59,N_446);
or U1402 (N_1402,N_1127,In_1561);
xnor U1403 (N_1403,N_829,In_429);
nor U1404 (N_1404,N_777,N_795);
nor U1405 (N_1405,N_1015,N_843);
nor U1406 (N_1406,N_751,In_1711);
nand U1407 (N_1407,In_272,N_1155);
or U1408 (N_1408,N_1071,In_1990);
nor U1409 (N_1409,N_602,N_522);
and U1410 (N_1410,In_236,N_952);
nor U1411 (N_1411,N_690,N_1038);
and U1412 (N_1412,N_893,N_968);
nor U1413 (N_1413,N_855,N_1103);
and U1414 (N_1414,N_341,N_1129);
nor U1415 (N_1415,In_1142,N_707);
or U1416 (N_1416,N_471,In_929);
nor U1417 (N_1417,In_1728,N_135);
xor U1418 (N_1418,N_525,In_314);
nor U1419 (N_1419,In_1254,In_296);
xnor U1420 (N_1420,N_863,In_1567);
xnor U1421 (N_1421,N_962,N_1048);
and U1422 (N_1422,N_999,N_428);
xor U1423 (N_1423,N_1057,In_1837);
or U1424 (N_1424,N_979,In_1241);
xnor U1425 (N_1425,N_181,N_873);
and U1426 (N_1426,N_1080,In_1263);
nand U1427 (N_1427,In_612,In_1380);
or U1428 (N_1428,N_1198,N_704);
nand U1429 (N_1429,N_905,In_1972);
and U1430 (N_1430,In_1119,In_1815);
or U1431 (N_1431,N_447,N_712);
xor U1432 (N_1432,N_1053,N_990);
xor U1433 (N_1433,N_1134,N_1140);
or U1434 (N_1434,In_94,N_1109);
nand U1435 (N_1435,N_512,N_146);
and U1436 (N_1436,N_508,In_1839);
nand U1437 (N_1437,N_953,N_877);
nor U1438 (N_1438,N_963,N_921);
or U1439 (N_1439,N_1035,N_903);
xor U1440 (N_1440,N_899,N_591);
and U1441 (N_1441,N_975,N_824);
or U1442 (N_1442,N_373,In_294);
nand U1443 (N_1443,In_37,N_914);
and U1444 (N_1444,In_1444,N_866);
and U1445 (N_1445,N_600,N_926);
xnor U1446 (N_1446,N_230,N_103);
and U1447 (N_1447,N_847,N_516);
nor U1448 (N_1448,N_890,N_657);
nor U1449 (N_1449,N_684,N_1106);
nand U1450 (N_1450,N_1002,N_1125);
or U1451 (N_1451,In_95,N_859);
or U1452 (N_1452,N_932,N_1157);
nor U1453 (N_1453,N_1074,N_1045);
and U1454 (N_1454,N_845,N_972);
and U1455 (N_1455,N_856,N_1085);
nor U1456 (N_1456,N_1081,N_1194);
xnor U1457 (N_1457,N_915,N_122);
nor U1458 (N_1458,In_735,In_1150);
and U1459 (N_1459,N_1069,N_1093);
nand U1460 (N_1460,In_1818,N_961);
or U1461 (N_1461,N_440,N_1182);
and U1462 (N_1462,N_936,N_871);
nor U1463 (N_1463,In_362,In_1431);
and U1464 (N_1464,N_1066,N_494);
or U1465 (N_1465,N_883,N_1165);
and U1466 (N_1466,N_998,N_966);
or U1467 (N_1467,N_762,N_931);
or U1468 (N_1468,N_519,In_70);
or U1469 (N_1469,In_82,N_1158);
nand U1470 (N_1470,N_1163,In_1060);
and U1471 (N_1471,N_803,N_1027);
and U1472 (N_1472,N_1082,N_827);
and U1473 (N_1473,In_547,In_1861);
or U1474 (N_1474,N_1128,In_103);
or U1475 (N_1475,N_1137,N_1064);
nor U1476 (N_1476,N_1124,N_924);
or U1477 (N_1477,N_1145,N_852);
or U1478 (N_1478,N_927,In_1336);
xnor U1479 (N_1479,N_967,N_929);
xor U1480 (N_1480,N_1180,N_781);
and U1481 (N_1481,In_69,N_1089);
nand U1482 (N_1482,In_610,N_1059);
nor U1483 (N_1483,In_1661,In_1317);
or U1484 (N_1484,N_532,In_906);
nor U1485 (N_1485,N_994,In_1626);
xor U1486 (N_1486,N_938,N_415);
or U1487 (N_1487,In_840,N_867);
xor U1488 (N_1488,In_297,N_948);
nand U1489 (N_1489,In_397,N_960);
nand U1490 (N_1490,N_995,In_937);
or U1491 (N_1491,In_899,N_738);
nand U1492 (N_1492,N_1008,N_71);
and U1493 (N_1493,N_788,In_742);
and U1494 (N_1494,N_1022,N_1003);
nor U1495 (N_1495,N_1144,N_1122);
and U1496 (N_1496,In_727,N_1154);
nor U1497 (N_1497,N_1068,N_564);
xor U1498 (N_1498,N_1147,N_610);
nor U1499 (N_1499,N_557,N_889);
and U1500 (N_1500,N_937,N_907);
or U1501 (N_1501,N_985,N_844);
nand U1502 (N_1502,N_504,N_858);
or U1503 (N_1503,N_100,N_1029);
xor U1504 (N_1504,N_976,N_563);
or U1505 (N_1505,In_268,In_1589);
xnor U1506 (N_1506,N_601,In_128);
nand U1507 (N_1507,N_1176,N_681);
and U1508 (N_1508,N_291,N_836);
nand U1509 (N_1509,N_766,N_536);
and U1510 (N_1510,In_1458,N_507);
xnor U1511 (N_1511,N_1072,In_592);
and U1512 (N_1512,N_605,N_806);
or U1513 (N_1513,In_759,N_561);
xnor U1514 (N_1514,In_799,N_131);
nor U1515 (N_1515,In_826,N_884);
nand U1516 (N_1516,N_1141,N_946);
or U1517 (N_1517,In_646,N_934);
or U1518 (N_1518,In_1895,N_935);
xnor U1519 (N_1519,N_983,N_897);
or U1520 (N_1520,N_774,N_57);
or U1521 (N_1521,N_1149,In_682);
and U1522 (N_1522,N_1115,N_1113);
and U1523 (N_1523,In_1087,In_739);
nand U1524 (N_1524,N_828,N_1043);
or U1525 (N_1525,In_1209,N_1075);
and U1526 (N_1526,N_197,N_556);
or U1527 (N_1527,In_1483,In_716);
nand U1528 (N_1528,N_930,N_898);
nor U1529 (N_1529,N_807,N_550);
nor U1530 (N_1530,N_981,In_368);
xnor U1531 (N_1531,In_613,N_232);
and U1532 (N_1532,N_448,In_897);
or U1533 (N_1533,N_1086,N_1111);
nand U1534 (N_1534,N_1116,N_809);
or U1535 (N_1535,N_1077,N_984);
xnor U1536 (N_1536,N_1186,In_1462);
xnor U1537 (N_1537,In_1992,N_969);
nor U1538 (N_1538,N_1044,N_1013);
or U1539 (N_1539,In_1516,N_16);
and U1540 (N_1540,In_939,N_1181);
or U1541 (N_1541,N_1058,N_399);
nor U1542 (N_1542,In_1031,N_1136);
and U1543 (N_1543,N_529,N_1055);
or U1544 (N_1544,N_804,N_1001);
nand U1545 (N_1545,N_680,N_1000);
and U1546 (N_1546,N_810,N_1065);
and U1547 (N_1547,N_1021,In_194);
and U1548 (N_1548,N_1108,N_989);
or U1549 (N_1549,N_837,N_823);
nor U1550 (N_1550,N_31,N_1118);
or U1551 (N_1551,N_805,In_166);
nand U1552 (N_1552,In_637,In_169);
and U1553 (N_1553,In_1219,N_1179);
or U1554 (N_1554,N_1096,N_474);
xor U1555 (N_1555,In_241,N_1185);
nand U1556 (N_1556,N_978,N_923);
or U1557 (N_1557,In_1806,N_726);
or U1558 (N_1558,N_1033,In_1212);
and U1559 (N_1559,In_892,N_1023);
or U1560 (N_1560,N_1087,In_1659);
nand U1561 (N_1561,In_1344,N_816);
nor U1562 (N_1562,N_430,N_1171);
or U1563 (N_1563,N_1020,N_860);
nor U1564 (N_1564,N_315,N_414);
xnor U1565 (N_1565,In_246,N_1039);
and U1566 (N_1566,N_951,N_585);
nor U1567 (N_1567,N_1110,N_944);
nor U1568 (N_1568,In_1833,N_840);
xnor U1569 (N_1569,N_1170,N_980);
nand U1570 (N_1570,N_1148,In_864);
and U1571 (N_1571,In_126,N_868);
xnor U1572 (N_1572,In_1337,In_1167);
nand U1573 (N_1573,N_1091,N_1079);
nand U1574 (N_1574,N_764,N_1196);
or U1575 (N_1575,In_1089,N_846);
xor U1576 (N_1576,N_800,N_1107);
nor U1577 (N_1577,In_1756,N_500);
nor U1578 (N_1578,N_917,In_1355);
nand U1579 (N_1579,N_481,N_562);
nand U1580 (N_1580,In_1486,In_1657);
and U1581 (N_1581,In_1088,N_343);
nand U1582 (N_1582,N_1046,N_1153);
or U1583 (N_1583,N_659,N_1135);
nor U1584 (N_1584,In_1865,In_1289);
xnor U1585 (N_1585,N_431,N_1143);
xor U1586 (N_1586,N_853,N_869);
or U1587 (N_1587,N_1190,N_891);
nor U1588 (N_1588,N_833,N_1009);
nor U1589 (N_1589,N_1006,N_1083);
or U1590 (N_1590,N_1019,N_449);
or U1591 (N_1591,N_1139,N_639);
nor U1592 (N_1592,N_472,N_1061);
nor U1593 (N_1593,N_1084,N_954);
and U1594 (N_1594,N_947,N_611);
nand U1595 (N_1595,N_973,N_1095);
and U1596 (N_1596,N_362,N_86);
or U1597 (N_1597,N_1133,N_1130);
and U1598 (N_1598,In_442,N_48);
xor U1599 (N_1599,N_33,In_244);
xor U1600 (N_1600,N_1414,N_1533);
nor U1601 (N_1601,N_1489,N_1265);
nand U1602 (N_1602,N_1376,N_1571);
nor U1603 (N_1603,N_1536,N_1517);
or U1604 (N_1604,N_1526,N_1227);
nand U1605 (N_1605,N_1587,N_1486);
xor U1606 (N_1606,N_1301,N_1535);
nand U1607 (N_1607,N_1212,N_1213);
xnor U1608 (N_1608,N_1454,N_1239);
or U1609 (N_1609,N_1396,N_1360);
or U1610 (N_1610,N_1322,N_1328);
nand U1611 (N_1611,N_1589,N_1218);
nor U1612 (N_1612,N_1488,N_1427);
or U1613 (N_1613,N_1594,N_1498);
nand U1614 (N_1614,N_1283,N_1547);
xnor U1615 (N_1615,N_1599,N_1242);
and U1616 (N_1616,N_1302,N_1300);
nor U1617 (N_1617,N_1553,N_1584);
or U1618 (N_1618,N_1275,N_1453);
xnor U1619 (N_1619,N_1209,N_1469);
nor U1620 (N_1620,N_1515,N_1542);
or U1621 (N_1621,N_1519,N_1540);
and U1622 (N_1622,N_1443,N_1492);
nor U1623 (N_1623,N_1309,N_1422);
nand U1624 (N_1624,N_1428,N_1579);
nand U1625 (N_1625,N_1387,N_1431);
nand U1626 (N_1626,N_1267,N_1389);
or U1627 (N_1627,N_1577,N_1470);
xnor U1628 (N_1628,N_1485,N_1397);
nand U1629 (N_1629,N_1590,N_1202);
xnor U1630 (N_1630,N_1429,N_1537);
nor U1631 (N_1631,N_1262,N_1543);
xor U1632 (N_1632,N_1316,N_1381);
or U1633 (N_1633,N_1296,N_1366);
xnor U1634 (N_1634,N_1356,N_1436);
nand U1635 (N_1635,N_1230,N_1483);
and U1636 (N_1636,N_1529,N_1509);
or U1637 (N_1637,N_1355,N_1413);
nor U1638 (N_1638,N_1285,N_1345);
or U1639 (N_1639,N_1390,N_1347);
nor U1640 (N_1640,N_1228,N_1541);
or U1641 (N_1641,N_1588,N_1578);
and U1642 (N_1642,N_1208,N_1241);
and U1643 (N_1643,N_1286,N_1277);
and U1644 (N_1644,N_1544,N_1268);
xor U1645 (N_1645,N_1290,N_1511);
nor U1646 (N_1646,N_1557,N_1260);
or U1647 (N_1647,N_1339,N_1531);
nor U1648 (N_1648,N_1391,N_1555);
nor U1649 (N_1649,N_1474,N_1365);
and U1650 (N_1650,N_1304,N_1507);
nand U1651 (N_1651,N_1246,N_1516);
nand U1652 (N_1652,N_1452,N_1580);
nor U1653 (N_1653,N_1412,N_1505);
nand U1654 (N_1654,N_1307,N_1289);
and U1655 (N_1655,N_1269,N_1565);
and U1656 (N_1656,N_1224,N_1459);
nor U1657 (N_1657,N_1359,N_1266);
nor U1658 (N_1658,N_1274,N_1513);
nor U1659 (N_1659,N_1203,N_1528);
and U1660 (N_1660,N_1424,N_1582);
xor U1661 (N_1661,N_1503,N_1433);
and U1662 (N_1662,N_1225,N_1221);
nor U1663 (N_1663,N_1477,N_1217);
nand U1664 (N_1664,N_1336,N_1320);
and U1665 (N_1665,N_1367,N_1292);
xnor U1666 (N_1666,N_1563,N_1349);
nand U1667 (N_1667,N_1313,N_1377);
nand U1668 (N_1668,N_1238,N_1575);
or U1669 (N_1669,N_1534,N_1506);
nand U1670 (N_1670,N_1251,N_1201);
nor U1671 (N_1671,N_1306,N_1423);
or U1672 (N_1672,N_1373,N_1403);
or U1673 (N_1673,N_1352,N_1402);
nand U1674 (N_1674,N_1530,N_1279);
nand U1675 (N_1675,N_1430,N_1438);
and U1676 (N_1676,N_1259,N_1244);
nor U1677 (N_1677,N_1338,N_1548);
and U1678 (N_1678,N_1404,N_1325);
nand U1679 (N_1679,N_1288,N_1445);
xnor U1680 (N_1680,N_1401,N_1425);
and U1681 (N_1681,N_1257,N_1372);
nand U1682 (N_1682,N_1234,N_1282);
nor U1683 (N_1683,N_1354,N_1434);
and U1684 (N_1684,N_1409,N_1329);
nor U1685 (N_1685,N_1346,N_1295);
nor U1686 (N_1686,N_1293,N_1466);
and U1687 (N_1687,N_1546,N_1441);
and U1688 (N_1688,N_1226,N_1362);
xor U1689 (N_1689,N_1576,N_1500);
nor U1690 (N_1690,N_1552,N_1214);
and U1691 (N_1691,N_1597,N_1585);
nor U1692 (N_1692,N_1432,N_1554);
nor U1693 (N_1693,N_1258,N_1421);
nor U1694 (N_1694,N_1574,N_1393);
xor U1695 (N_1695,N_1216,N_1596);
xnor U1696 (N_1696,N_1384,N_1317);
xnor U1697 (N_1697,N_1235,N_1512);
and U1698 (N_1698,N_1471,N_1406);
xor U1699 (N_1699,N_1375,N_1514);
xor U1700 (N_1700,N_1254,N_1206);
and U1701 (N_1701,N_1276,N_1399);
or U1702 (N_1702,N_1567,N_1368);
nand U1703 (N_1703,N_1324,N_1314);
nand U1704 (N_1704,N_1358,N_1457);
or U1705 (N_1705,N_1237,N_1508);
and U1706 (N_1706,N_1473,N_1504);
xnor U1707 (N_1707,N_1463,N_1523);
xnor U1708 (N_1708,N_1308,N_1250);
nor U1709 (N_1709,N_1478,N_1570);
and U1710 (N_1710,N_1363,N_1524);
nor U1711 (N_1711,N_1200,N_1331);
xnor U1712 (N_1712,N_1298,N_1545);
nor U1713 (N_1713,N_1326,N_1558);
and U1714 (N_1714,N_1497,N_1521);
nor U1715 (N_1715,N_1371,N_1484);
or U1716 (N_1716,N_1518,N_1245);
xnor U1717 (N_1717,N_1278,N_1207);
and U1718 (N_1718,N_1496,N_1353);
nand U1719 (N_1719,N_1499,N_1487);
and U1720 (N_1720,N_1568,N_1479);
nand U1721 (N_1721,N_1598,N_1291);
nor U1722 (N_1722,N_1551,N_1416);
and U1723 (N_1723,N_1231,N_1595);
nand U1724 (N_1724,N_1481,N_1229);
and U1725 (N_1725,N_1204,N_1591);
or U1726 (N_1726,N_1270,N_1476);
xnor U1727 (N_1727,N_1440,N_1380);
or U1728 (N_1728,N_1348,N_1319);
and U1729 (N_1729,N_1253,N_1263);
nand U1730 (N_1730,N_1586,N_1520);
nand U1731 (N_1731,N_1223,N_1573);
or U1732 (N_1732,N_1420,N_1388);
nand U1733 (N_1733,N_1233,N_1556);
or U1734 (N_1734,N_1252,N_1323);
and U1735 (N_1735,N_1446,N_1394);
or U1736 (N_1736,N_1462,N_1383);
and U1737 (N_1737,N_1386,N_1205);
or U1738 (N_1738,N_1550,N_1572);
or U1739 (N_1739,N_1418,N_1593);
nand U1740 (N_1740,N_1315,N_1311);
nand U1741 (N_1741,N_1344,N_1439);
nand U1742 (N_1742,N_1232,N_1340);
nor U1743 (N_1743,N_1456,N_1458);
nor U1744 (N_1744,N_1256,N_1379);
xor U1745 (N_1745,N_1482,N_1261);
and U1746 (N_1746,N_1271,N_1303);
nor U1747 (N_1747,N_1312,N_1475);
xor U1748 (N_1748,N_1243,N_1211);
xnor U1749 (N_1749,N_1564,N_1335);
nor U1750 (N_1750,N_1215,N_1334);
nor U1751 (N_1751,N_1467,N_1342);
xnor U1752 (N_1752,N_1549,N_1447);
or U1753 (N_1753,N_1330,N_1273);
nand U1754 (N_1754,N_1501,N_1451);
xor U1755 (N_1755,N_1392,N_1248);
nor U1756 (N_1756,N_1357,N_1294);
and U1757 (N_1757,N_1461,N_1464);
nand U1758 (N_1758,N_1411,N_1510);
xor U1759 (N_1759,N_1210,N_1272);
or U1760 (N_1760,N_1249,N_1341);
or U1761 (N_1761,N_1236,N_1494);
nor U1762 (N_1762,N_1332,N_1562);
nand U1763 (N_1763,N_1539,N_1343);
nor U1764 (N_1764,N_1310,N_1351);
and U1765 (N_1765,N_1240,N_1280);
or U1766 (N_1766,N_1378,N_1472);
nand U1767 (N_1767,N_1287,N_1415);
or U1768 (N_1768,N_1222,N_1491);
or U1769 (N_1769,N_1395,N_1321);
or U1770 (N_1770,N_1264,N_1468);
and U1771 (N_1771,N_1398,N_1495);
nand U1772 (N_1772,N_1449,N_1493);
or U1773 (N_1773,N_1361,N_1437);
nor U1774 (N_1774,N_1281,N_1370);
nand U1775 (N_1775,N_1581,N_1559);
nand U1776 (N_1776,N_1538,N_1299);
and U1777 (N_1777,N_1566,N_1400);
xor U1778 (N_1778,N_1364,N_1480);
xor U1779 (N_1779,N_1318,N_1460);
nor U1780 (N_1780,N_1444,N_1220);
and U1781 (N_1781,N_1369,N_1407);
xnor U1782 (N_1782,N_1527,N_1442);
xor U1783 (N_1783,N_1455,N_1465);
xnor U1784 (N_1784,N_1385,N_1522);
xnor U1785 (N_1785,N_1333,N_1382);
or U1786 (N_1786,N_1417,N_1525);
or U1787 (N_1787,N_1305,N_1561);
and U1788 (N_1788,N_1327,N_1490);
nor U1789 (N_1789,N_1374,N_1247);
and U1790 (N_1790,N_1560,N_1419);
nor U1791 (N_1791,N_1448,N_1337);
xor U1792 (N_1792,N_1255,N_1350);
and U1793 (N_1793,N_1450,N_1405);
or U1794 (N_1794,N_1284,N_1502);
and U1795 (N_1795,N_1408,N_1435);
nor U1796 (N_1796,N_1583,N_1219);
nor U1797 (N_1797,N_1569,N_1297);
xor U1798 (N_1798,N_1410,N_1532);
nor U1799 (N_1799,N_1592,N_1426);
nor U1800 (N_1800,N_1230,N_1470);
nor U1801 (N_1801,N_1326,N_1249);
or U1802 (N_1802,N_1283,N_1430);
or U1803 (N_1803,N_1479,N_1400);
xnor U1804 (N_1804,N_1259,N_1439);
and U1805 (N_1805,N_1281,N_1237);
nand U1806 (N_1806,N_1394,N_1598);
and U1807 (N_1807,N_1240,N_1289);
and U1808 (N_1808,N_1222,N_1231);
nand U1809 (N_1809,N_1233,N_1483);
and U1810 (N_1810,N_1541,N_1549);
nand U1811 (N_1811,N_1235,N_1449);
or U1812 (N_1812,N_1589,N_1526);
nor U1813 (N_1813,N_1327,N_1537);
nand U1814 (N_1814,N_1405,N_1246);
nor U1815 (N_1815,N_1593,N_1507);
or U1816 (N_1816,N_1235,N_1406);
xnor U1817 (N_1817,N_1540,N_1423);
and U1818 (N_1818,N_1336,N_1402);
and U1819 (N_1819,N_1252,N_1320);
and U1820 (N_1820,N_1348,N_1298);
nor U1821 (N_1821,N_1502,N_1201);
or U1822 (N_1822,N_1529,N_1208);
nor U1823 (N_1823,N_1236,N_1543);
and U1824 (N_1824,N_1420,N_1402);
and U1825 (N_1825,N_1271,N_1217);
nor U1826 (N_1826,N_1366,N_1297);
and U1827 (N_1827,N_1520,N_1427);
and U1828 (N_1828,N_1599,N_1260);
nor U1829 (N_1829,N_1555,N_1428);
nand U1830 (N_1830,N_1332,N_1554);
xor U1831 (N_1831,N_1213,N_1467);
xnor U1832 (N_1832,N_1546,N_1511);
xor U1833 (N_1833,N_1274,N_1394);
nor U1834 (N_1834,N_1479,N_1516);
or U1835 (N_1835,N_1573,N_1485);
nand U1836 (N_1836,N_1473,N_1233);
xor U1837 (N_1837,N_1545,N_1444);
xnor U1838 (N_1838,N_1499,N_1304);
or U1839 (N_1839,N_1433,N_1284);
or U1840 (N_1840,N_1587,N_1327);
xor U1841 (N_1841,N_1563,N_1356);
xor U1842 (N_1842,N_1545,N_1212);
nand U1843 (N_1843,N_1413,N_1568);
xor U1844 (N_1844,N_1513,N_1542);
xnor U1845 (N_1845,N_1496,N_1520);
nand U1846 (N_1846,N_1496,N_1360);
and U1847 (N_1847,N_1334,N_1489);
nor U1848 (N_1848,N_1252,N_1326);
nand U1849 (N_1849,N_1570,N_1409);
xnor U1850 (N_1850,N_1291,N_1562);
nand U1851 (N_1851,N_1436,N_1382);
nand U1852 (N_1852,N_1367,N_1584);
and U1853 (N_1853,N_1246,N_1374);
xnor U1854 (N_1854,N_1562,N_1231);
nor U1855 (N_1855,N_1278,N_1248);
and U1856 (N_1856,N_1303,N_1306);
and U1857 (N_1857,N_1500,N_1369);
or U1858 (N_1858,N_1566,N_1554);
and U1859 (N_1859,N_1316,N_1300);
nand U1860 (N_1860,N_1373,N_1430);
or U1861 (N_1861,N_1403,N_1585);
and U1862 (N_1862,N_1536,N_1331);
nand U1863 (N_1863,N_1482,N_1258);
or U1864 (N_1864,N_1423,N_1428);
nor U1865 (N_1865,N_1246,N_1570);
or U1866 (N_1866,N_1211,N_1345);
or U1867 (N_1867,N_1231,N_1201);
nand U1868 (N_1868,N_1543,N_1367);
xor U1869 (N_1869,N_1380,N_1540);
or U1870 (N_1870,N_1261,N_1362);
and U1871 (N_1871,N_1372,N_1311);
and U1872 (N_1872,N_1495,N_1450);
xor U1873 (N_1873,N_1460,N_1305);
and U1874 (N_1874,N_1431,N_1398);
or U1875 (N_1875,N_1325,N_1595);
nand U1876 (N_1876,N_1369,N_1395);
nand U1877 (N_1877,N_1391,N_1368);
xor U1878 (N_1878,N_1538,N_1537);
or U1879 (N_1879,N_1284,N_1324);
and U1880 (N_1880,N_1290,N_1544);
nor U1881 (N_1881,N_1261,N_1416);
nand U1882 (N_1882,N_1428,N_1279);
nand U1883 (N_1883,N_1367,N_1432);
nand U1884 (N_1884,N_1519,N_1507);
nor U1885 (N_1885,N_1245,N_1487);
or U1886 (N_1886,N_1299,N_1412);
nor U1887 (N_1887,N_1270,N_1577);
or U1888 (N_1888,N_1265,N_1270);
xnor U1889 (N_1889,N_1327,N_1238);
xor U1890 (N_1890,N_1327,N_1368);
xor U1891 (N_1891,N_1230,N_1451);
nand U1892 (N_1892,N_1586,N_1577);
and U1893 (N_1893,N_1481,N_1216);
nand U1894 (N_1894,N_1228,N_1547);
and U1895 (N_1895,N_1543,N_1478);
nor U1896 (N_1896,N_1275,N_1309);
and U1897 (N_1897,N_1576,N_1462);
and U1898 (N_1898,N_1389,N_1208);
nor U1899 (N_1899,N_1325,N_1459);
nor U1900 (N_1900,N_1349,N_1573);
and U1901 (N_1901,N_1210,N_1390);
nand U1902 (N_1902,N_1328,N_1411);
xor U1903 (N_1903,N_1453,N_1398);
and U1904 (N_1904,N_1260,N_1479);
and U1905 (N_1905,N_1450,N_1356);
or U1906 (N_1906,N_1362,N_1231);
nand U1907 (N_1907,N_1405,N_1334);
nand U1908 (N_1908,N_1381,N_1238);
and U1909 (N_1909,N_1344,N_1272);
nor U1910 (N_1910,N_1423,N_1514);
and U1911 (N_1911,N_1322,N_1412);
xor U1912 (N_1912,N_1565,N_1394);
nor U1913 (N_1913,N_1367,N_1561);
nor U1914 (N_1914,N_1211,N_1314);
and U1915 (N_1915,N_1269,N_1554);
xnor U1916 (N_1916,N_1404,N_1343);
and U1917 (N_1917,N_1271,N_1428);
nor U1918 (N_1918,N_1450,N_1553);
nand U1919 (N_1919,N_1233,N_1478);
or U1920 (N_1920,N_1264,N_1347);
and U1921 (N_1921,N_1560,N_1401);
xnor U1922 (N_1922,N_1580,N_1565);
and U1923 (N_1923,N_1542,N_1317);
or U1924 (N_1924,N_1483,N_1298);
xnor U1925 (N_1925,N_1420,N_1499);
nand U1926 (N_1926,N_1295,N_1490);
nand U1927 (N_1927,N_1579,N_1395);
or U1928 (N_1928,N_1496,N_1519);
xor U1929 (N_1929,N_1443,N_1580);
xor U1930 (N_1930,N_1249,N_1505);
nand U1931 (N_1931,N_1270,N_1279);
and U1932 (N_1932,N_1410,N_1528);
nand U1933 (N_1933,N_1459,N_1532);
and U1934 (N_1934,N_1303,N_1215);
and U1935 (N_1935,N_1231,N_1246);
nand U1936 (N_1936,N_1597,N_1259);
nor U1937 (N_1937,N_1507,N_1209);
nand U1938 (N_1938,N_1543,N_1389);
or U1939 (N_1939,N_1289,N_1525);
xor U1940 (N_1940,N_1217,N_1556);
nand U1941 (N_1941,N_1276,N_1254);
xnor U1942 (N_1942,N_1331,N_1546);
and U1943 (N_1943,N_1256,N_1331);
and U1944 (N_1944,N_1575,N_1209);
xor U1945 (N_1945,N_1351,N_1462);
and U1946 (N_1946,N_1381,N_1389);
nand U1947 (N_1947,N_1474,N_1589);
nand U1948 (N_1948,N_1470,N_1232);
or U1949 (N_1949,N_1552,N_1338);
and U1950 (N_1950,N_1514,N_1220);
xor U1951 (N_1951,N_1574,N_1241);
xor U1952 (N_1952,N_1211,N_1546);
nor U1953 (N_1953,N_1568,N_1344);
xnor U1954 (N_1954,N_1467,N_1325);
or U1955 (N_1955,N_1369,N_1541);
nand U1956 (N_1956,N_1395,N_1576);
nand U1957 (N_1957,N_1435,N_1318);
and U1958 (N_1958,N_1535,N_1581);
xnor U1959 (N_1959,N_1449,N_1599);
and U1960 (N_1960,N_1436,N_1594);
or U1961 (N_1961,N_1268,N_1215);
or U1962 (N_1962,N_1281,N_1224);
xnor U1963 (N_1963,N_1389,N_1548);
nand U1964 (N_1964,N_1374,N_1323);
nor U1965 (N_1965,N_1559,N_1578);
and U1966 (N_1966,N_1403,N_1239);
or U1967 (N_1967,N_1265,N_1323);
xnor U1968 (N_1968,N_1296,N_1292);
and U1969 (N_1969,N_1250,N_1409);
or U1970 (N_1970,N_1503,N_1561);
or U1971 (N_1971,N_1365,N_1242);
or U1972 (N_1972,N_1270,N_1441);
and U1973 (N_1973,N_1362,N_1567);
xnor U1974 (N_1974,N_1506,N_1447);
or U1975 (N_1975,N_1580,N_1537);
and U1976 (N_1976,N_1201,N_1495);
or U1977 (N_1977,N_1358,N_1212);
and U1978 (N_1978,N_1263,N_1307);
and U1979 (N_1979,N_1255,N_1488);
xor U1980 (N_1980,N_1320,N_1563);
or U1981 (N_1981,N_1360,N_1345);
nand U1982 (N_1982,N_1268,N_1252);
or U1983 (N_1983,N_1201,N_1348);
xnor U1984 (N_1984,N_1387,N_1549);
nor U1985 (N_1985,N_1434,N_1326);
xor U1986 (N_1986,N_1536,N_1409);
or U1987 (N_1987,N_1371,N_1238);
nor U1988 (N_1988,N_1390,N_1460);
xor U1989 (N_1989,N_1462,N_1371);
xnor U1990 (N_1990,N_1465,N_1514);
nor U1991 (N_1991,N_1496,N_1511);
and U1992 (N_1992,N_1496,N_1264);
nor U1993 (N_1993,N_1301,N_1588);
nor U1994 (N_1994,N_1473,N_1346);
or U1995 (N_1995,N_1430,N_1218);
or U1996 (N_1996,N_1443,N_1378);
or U1997 (N_1997,N_1261,N_1512);
xor U1998 (N_1998,N_1452,N_1599);
nand U1999 (N_1999,N_1374,N_1464);
nand U2000 (N_2000,N_1962,N_1921);
xnor U2001 (N_2001,N_1854,N_1663);
xor U2002 (N_2002,N_1658,N_1701);
or U2003 (N_2003,N_1636,N_1847);
nor U2004 (N_2004,N_1771,N_1920);
nor U2005 (N_2005,N_1896,N_1774);
xnor U2006 (N_2006,N_1825,N_1932);
nand U2007 (N_2007,N_1633,N_1722);
xor U2008 (N_2008,N_1787,N_1839);
and U2009 (N_2009,N_1826,N_1754);
nand U2010 (N_2010,N_1634,N_1809);
nor U2011 (N_2011,N_1657,N_1866);
xor U2012 (N_2012,N_1968,N_1939);
and U2013 (N_2013,N_1845,N_1645);
nor U2014 (N_2014,N_1913,N_1652);
nand U2015 (N_2015,N_1943,N_1702);
xor U2016 (N_2016,N_1791,N_1621);
nand U2017 (N_2017,N_1819,N_1990);
or U2018 (N_2018,N_1830,N_1811);
xnor U2019 (N_2019,N_1800,N_1924);
or U2020 (N_2020,N_1869,N_1901);
xor U2021 (N_2021,N_1824,N_1646);
and U2022 (N_2022,N_1688,N_1742);
and U2023 (N_2023,N_1915,N_1952);
nand U2024 (N_2024,N_1833,N_1785);
nand U2025 (N_2025,N_1991,N_1971);
nand U2026 (N_2026,N_1929,N_1673);
and U2027 (N_2027,N_1680,N_1834);
and U2028 (N_2028,N_1773,N_1922);
nand U2029 (N_2029,N_1644,N_1649);
nor U2030 (N_2030,N_1606,N_1998);
or U2031 (N_2031,N_1697,N_1717);
nor U2032 (N_2032,N_1861,N_1882);
and U2033 (N_2033,N_1863,N_1605);
xor U2034 (N_2034,N_1797,N_1953);
xnor U2035 (N_2035,N_1788,N_1611);
nor U2036 (N_2036,N_1950,N_1677);
nand U2037 (N_2037,N_1767,N_1617);
nor U2038 (N_2038,N_1978,N_1986);
or U2039 (N_2039,N_1955,N_1622);
nor U2040 (N_2040,N_1959,N_1779);
xnor U2041 (N_2041,N_1996,N_1780);
and U2042 (N_2042,N_1711,N_1739);
xnor U2043 (N_2043,N_1719,N_1887);
xnor U2044 (N_2044,N_1619,N_1841);
xor U2045 (N_2045,N_1855,N_1620);
xor U2046 (N_2046,N_1661,N_1917);
or U2047 (N_2047,N_1683,N_1975);
or U2048 (N_2048,N_1879,N_1902);
xnor U2049 (N_2049,N_1851,N_1713);
and U2050 (N_2050,N_1789,N_1935);
and U2051 (N_2051,N_1815,N_1752);
nor U2052 (N_2052,N_1691,N_1642);
nor U2053 (N_2053,N_1656,N_1686);
nand U2054 (N_2054,N_1872,N_1653);
and U2055 (N_2055,N_1625,N_1793);
xnor U2056 (N_2056,N_1602,N_1897);
or U2057 (N_2057,N_1980,N_1958);
nand U2058 (N_2058,N_1660,N_1731);
nand U2059 (N_2059,N_1782,N_1893);
nand U2060 (N_2060,N_1796,N_1669);
nor U2061 (N_2061,N_1670,N_1799);
nand U2062 (N_2062,N_1940,N_1890);
nand U2063 (N_2063,N_1807,N_1836);
xnor U2064 (N_2064,N_1979,N_1770);
and U2065 (N_2065,N_1601,N_1792);
nor U2066 (N_2066,N_1886,N_1698);
nand U2067 (N_2067,N_1870,N_1741);
nand U2068 (N_2068,N_1969,N_1842);
or U2069 (N_2069,N_1676,N_1694);
and U2070 (N_2070,N_1600,N_1678);
xor U2071 (N_2071,N_1786,N_1639);
nand U2072 (N_2072,N_1899,N_1727);
and U2073 (N_2073,N_1864,N_1859);
and U2074 (N_2074,N_1818,N_1994);
xnor U2075 (N_2075,N_1945,N_1710);
or U2076 (N_2076,N_1848,N_1999);
nand U2077 (N_2077,N_1726,N_1734);
or U2078 (N_2078,N_1755,N_1838);
xor U2079 (N_2079,N_1972,N_1712);
or U2080 (N_2080,N_1884,N_1610);
nor U2081 (N_2081,N_1984,N_1725);
nor U2082 (N_2082,N_1853,N_1757);
xor U2083 (N_2083,N_1703,N_1812);
and U2084 (N_2084,N_1808,N_1758);
nand U2085 (N_2085,N_1695,N_1720);
nor U2086 (N_2086,N_1748,N_1876);
or U2087 (N_2087,N_1696,N_1831);
and U2088 (N_2088,N_1988,N_1928);
nor U2089 (N_2089,N_1987,N_1765);
or U2090 (N_2090,N_1735,N_1655);
and U2091 (N_2091,N_1860,N_1936);
xnor U2092 (N_2092,N_1946,N_1967);
and U2093 (N_2093,N_1918,N_1730);
and U2094 (N_2094,N_1751,N_1806);
xnor U2095 (N_2095,N_1608,N_1891);
nor U2096 (N_2096,N_1700,N_1689);
nor U2097 (N_2097,N_1750,N_1692);
and U2098 (N_2098,N_1919,N_1867);
and U2099 (N_2099,N_1927,N_1900);
or U2100 (N_2100,N_1822,N_1963);
and U2101 (N_2101,N_1760,N_1715);
or U2102 (N_2102,N_1966,N_1837);
nand U2103 (N_2103,N_1829,N_1895);
nand U2104 (N_2104,N_1934,N_1856);
nor U2105 (N_2105,N_1944,N_1613);
nor U2106 (N_2106,N_1714,N_1965);
nand U2107 (N_2107,N_1981,N_1883);
or U2108 (N_2108,N_1708,N_1705);
and U2109 (N_2109,N_1684,N_1664);
nor U2110 (N_2110,N_1964,N_1740);
nand U2111 (N_2111,N_1828,N_1623);
xor U2112 (N_2112,N_1704,N_1805);
or U2113 (N_2113,N_1628,N_1736);
and U2114 (N_2114,N_1762,N_1948);
nand U2115 (N_2115,N_1681,N_1777);
nor U2116 (N_2116,N_1641,N_1629);
or U2117 (N_2117,N_1744,N_1763);
and U2118 (N_2118,N_1654,N_1849);
or U2119 (N_2119,N_1668,N_1888);
and U2120 (N_2120,N_1904,N_1956);
nand U2121 (N_2121,N_1857,N_1905);
nand U2122 (N_2122,N_1685,N_1630);
nor U2123 (N_2123,N_1638,N_1938);
and U2124 (N_2124,N_1976,N_1894);
nand U2125 (N_2125,N_1759,N_1775);
or U2126 (N_2126,N_1862,N_1603);
nor U2127 (N_2127,N_1957,N_1880);
nand U2128 (N_2128,N_1690,N_1724);
or U2129 (N_2129,N_1970,N_1781);
xor U2130 (N_2130,N_1618,N_1709);
and U2131 (N_2131,N_1733,N_1674);
and U2132 (N_2132,N_1877,N_1865);
xnor U2133 (N_2133,N_1973,N_1868);
nand U2134 (N_2134,N_1844,N_1954);
or U2135 (N_2135,N_1672,N_1648);
nand U2136 (N_2136,N_1614,N_1827);
or U2137 (N_2137,N_1840,N_1616);
or U2138 (N_2138,N_1647,N_1982);
or U2139 (N_2139,N_1804,N_1640);
and U2140 (N_2140,N_1749,N_1776);
xnor U2141 (N_2141,N_1914,N_1995);
nand U2142 (N_2142,N_1931,N_1667);
nand U2143 (N_2143,N_1783,N_1960);
nor U2144 (N_2144,N_1993,N_1632);
and U2145 (N_2145,N_1659,N_1949);
and U2146 (N_2146,N_1768,N_1743);
or U2147 (N_2147,N_1983,N_1843);
and U2148 (N_2148,N_1937,N_1769);
and U2149 (N_2149,N_1912,N_1989);
nor U2150 (N_2150,N_1604,N_1974);
or U2151 (N_2151,N_1930,N_1790);
and U2152 (N_2152,N_1977,N_1612);
and U2153 (N_2153,N_1687,N_1832);
or U2154 (N_2154,N_1728,N_1816);
or U2155 (N_2155,N_1772,N_1911);
nand U2156 (N_2156,N_1784,N_1666);
or U2157 (N_2157,N_1651,N_1801);
or U2158 (N_2158,N_1846,N_1803);
and U2159 (N_2159,N_1675,N_1906);
and U2160 (N_2160,N_1795,N_1814);
and U2161 (N_2161,N_1820,N_1881);
and U2162 (N_2162,N_1761,N_1745);
xnor U2163 (N_2163,N_1650,N_1794);
and U2164 (N_2164,N_1941,N_1933);
or U2165 (N_2165,N_1961,N_1738);
nand U2166 (N_2166,N_1823,N_1707);
nand U2167 (N_2167,N_1908,N_1753);
and U2168 (N_2168,N_1637,N_1671);
xnor U2169 (N_2169,N_1732,N_1873);
or U2170 (N_2170,N_1746,N_1643);
nand U2171 (N_2171,N_1992,N_1892);
nand U2172 (N_2172,N_1723,N_1871);
nor U2173 (N_2173,N_1665,N_1898);
xnor U2174 (N_2174,N_1721,N_1766);
or U2175 (N_2175,N_1852,N_1615);
nand U2176 (N_2176,N_1798,N_1903);
xnor U2177 (N_2177,N_1682,N_1909);
nand U2178 (N_2178,N_1885,N_1607);
nor U2179 (N_2179,N_1624,N_1858);
and U2180 (N_2180,N_1916,N_1942);
and U2181 (N_2181,N_1718,N_1627);
xnor U2182 (N_2182,N_1889,N_1821);
xor U2183 (N_2183,N_1875,N_1631);
nand U2184 (N_2184,N_1810,N_1878);
nand U2185 (N_2185,N_1835,N_1716);
xnor U2186 (N_2186,N_1626,N_1850);
nand U2187 (N_2187,N_1706,N_1756);
xnor U2188 (N_2188,N_1817,N_1778);
nor U2189 (N_2189,N_1737,N_1729);
nand U2190 (N_2190,N_1947,N_1609);
nand U2191 (N_2191,N_1699,N_1951);
xnor U2192 (N_2192,N_1662,N_1693);
and U2193 (N_2193,N_1813,N_1802);
nand U2194 (N_2194,N_1926,N_1747);
nand U2195 (N_2195,N_1874,N_1985);
or U2196 (N_2196,N_1635,N_1923);
nor U2197 (N_2197,N_1907,N_1997);
nand U2198 (N_2198,N_1764,N_1910);
and U2199 (N_2199,N_1925,N_1679);
nand U2200 (N_2200,N_1622,N_1797);
and U2201 (N_2201,N_1898,N_1940);
nand U2202 (N_2202,N_1982,N_1748);
or U2203 (N_2203,N_1638,N_1724);
nand U2204 (N_2204,N_1850,N_1872);
nor U2205 (N_2205,N_1994,N_1781);
or U2206 (N_2206,N_1861,N_1851);
or U2207 (N_2207,N_1853,N_1726);
and U2208 (N_2208,N_1744,N_1680);
nand U2209 (N_2209,N_1861,N_1884);
xnor U2210 (N_2210,N_1788,N_1741);
and U2211 (N_2211,N_1964,N_1878);
and U2212 (N_2212,N_1880,N_1695);
and U2213 (N_2213,N_1855,N_1682);
or U2214 (N_2214,N_1609,N_1729);
and U2215 (N_2215,N_1937,N_1831);
and U2216 (N_2216,N_1771,N_1615);
or U2217 (N_2217,N_1630,N_1942);
nor U2218 (N_2218,N_1756,N_1882);
nand U2219 (N_2219,N_1886,N_1884);
and U2220 (N_2220,N_1717,N_1945);
or U2221 (N_2221,N_1925,N_1901);
nand U2222 (N_2222,N_1885,N_1770);
or U2223 (N_2223,N_1770,N_1957);
or U2224 (N_2224,N_1788,N_1822);
or U2225 (N_2225,N_1912,N_1920);
and U2226 (N_2226,N_1816,N_1908);
nor U2227 (N_2227,N_1654,N_1662);
nor U2228 (N_2228,N_1853,N_1905);
nand U2229 (N_2229,N_1956,N_1746);
nor U2230 (N_2230,N_1918,N_1799);
and U2231 (N_2231,N_1876,N_1925);
or U2232 (N_2232,N_1985,N_1818);
nand U2233 (N_2233,N_1616,N_1605);
nand U2234 (N_2234,N_1656,N_1675);
nand U2235 (N_2235,N_1887,N_1952);
xor U2236 (N_2236,N_1991,N_1956);
xnor U2237 (N_2237,N_1708,N_1825);
nand U2238 (N_2238,N_1750,N_1904);
xnor U2239 (N_2239,N_1987,N_1928);
nor U2240 (N_2240,N_1718,N_1820);
nor U2241 (N_2241,N_1736,N_1803);
nand U2242 (N_2242,N_1960,N_1691);
or U2243 (N_2243,N_1993,N_1883);
nand U2244 (N_2244,N_1928,N_1912);
xnor U2245 (N_2245,N_1966,N_1683);
or U2246 (N_2246,N_1815,N_1789);
nor U2247 (N_2247,N_1977,N_1987);
or U2248 (N_2248,N_1772,N_1765);
and U2249 (N_2249,N_1935,N_1681);
and U2250 (N_2250,N_1756,N_1739);
or U2251 (N_2251,N_1958,N_1866);
nor U2252 (N_2252,N_1773,N_1655);
xnor U2253 (N_2253,N_1729,N_1628);
nor U2254 (N_2254,N_1988,N_1828);
nor U2255 (N_2255,N_1938,N_1701);
xnor U2256 (N_2256,N_1776,N_1681);
or U2257 (N_2257,N_1610,N_1615);
xnor U2258 (N_2258,N_1919,N_1753);
nor U2259 (N_2259,N_1840,N_1806);
xnor U2260 (N_2260,N_1631,N_1849);
or U2261 (N_2261,N_1629,N_1875);
nand U2262 (N_2262,N_1790,N_1764);
xor U2263 (N_2263,N_1833,N_1673);
nor U2264 (N_2264,N_1627,N_1699);
and U2265 (N_2265,N_1766,N_1775);
nand U2266 (N_2266,N_1692,N_1854);
and U2267 (N_2267,N_1899,N_1793);
nand U2268 (N_2268,N_1770,N_1888);
and U2269 (N_2269,N_1905,N_1631);
xor U2270 (N_2270,N_1774,N_1935);
nor U2271 (N_2271,N_1831,N_1971);
or U2272 (N_2272,N_1804,N_1646);
and U2273 (N_2273,N_1816,N_1849);
nand U2274 (N_2274,N_1964,N_1856);
or U2275 (N_2275,N_1823,N_1993);
xnor U2276 (N_2276,N_1841,N_1981);
nand U2277 (N_2277,N_1833,N_1936);
nor U2278 (N_2278,N_1853,N_1983);
nor U2279 (N_2279,N_1960,N_1871);
xnor U2280 (N_2280,N_1745,N_1731);
nor U2281 (N_2281,N_1985,N_1765);
nor U2282 (N_2282,N_1808,N_1681);
xor U2283 (N_2283,N_1655,N_1794);
nor U2284 (N_2284,N_1839,N_1684);
or U2285 (N_2285,N_1652,N_1979);
nor U2286 (N_2286,N_1849,N_1903);
nand U2287 (N_2287,N_1976,N_1678);
xor U2288 (N_2288,N_1934,N_1965);
and U2289 (N_2289,N_1652,N_1644);
nand U2290 (N_2290,N_1947,N_1867);
nor U2291 (N_2291,N_1729,N_1856);
xor U2292 (N_2292,N_1814,N_1738);
or U2293 (N_2293,N_1667,N_1840);
xor U2294 (N_2294,N_1761,N_1849);
xor U2295 (N_2295,N_1950,N_1976);
nor U2296 (N_2296,N_1649,N_1672);
xnor U2297 (N_2297,N_1984,N_1768);
or U2298 (N_2298,N_1998,N_1695);
or U2299 (N_2299,N_1643,N_1763);
xor U2300 (N_2300,N_1721,N_1817);
xor U2301 (N_2301,N_1677,N_1973);
nor U2302 (N_2302,N_1832,N_1803);
xor U2303 (N_2303,N_1655,N_1861);
and U2304 (N_2304,N_1995,N_1783);
xnor U2305 (N_2305,N_1994,N_1886);
or U2306 (N_2306,N_1884,N_1679);
nand U2307 (N_2307,N_1732,N_1945);
and U2308 (N_2308,N_1935,N_1876);
xor U2309 (N_2309,N_1708,N_1796);
or U2310 (N_2310,N_1922,N_1813);
xnor U2311 (N_2311,N_1781,N_1759);
or U2312 (N_2312,N_1704,N_1647);
xor U2313 (N_2313,N_1643,N_1632);
and U2314 (N_2314,N_1951,N_1933);
nand U2315 (N_2315,N_1849,N_1706);
or U2316 (N_2316,N_1767,N_1721);
or U2317 (N_2317,N_1689,N_1682);
xnor U2318 (N_2318,N_1959,N_1924);
and U2319 (N_2319,N_1829,N_1894);
or U2320 (N_2320,N_1604,N_1816);
or U2321 (N_2321,N_1732,N_1793);
nor U2322 (N_2322,N_1624,N_1842);
or U2323 (N_2323,N_1821,N_1923);
and U2324 (N_2324,N_1986,N_1676);
and U2325 (N_2325,N_1706,N_1654);
xnor U2326 (N_2326,N_1601,N_1655);
or U2327 (N_2327,N_1783,N_1935);
xnor U2328 (N_2328,N_1867,N_1862);
nor U2329 (N_2329,N_1877,N_1626);
xnor U2330 (N_2330,N_1814,N_1711);
nor U2331 (N_2331,N_1674,N_1726);
and U2332 (N_2332,N_1963,N_1682);
xnor U2333 (N_2333,N_1989,N_1624);
nand U2334 (N_2334,N_1662,N_1674);
xor U2335 (N_2335,N_1636,N_1620);
and U2336 (N_2336,N_1665,N_1743);
or U2337 (N_2337,N_1657,N_1602);
xor U2338 (N_2338,N_1771,N_1726);
nand U2339 (N_2339,N_1766,N_1718);
or U2340 (N_2340,N_1753,N_1639);
and U2341 (N_2341,N_1915,N_1614);
xor U2342 (N_2342,N_1709,N_1652);
or U2343 (N_2343,N_1676,N_1687);
and U2344 (N_2344,N_1848,N_1846);
xor U2345 (N_2345,N_1609,N_1850);
and U2346 (N_2346,N_1986,N_1902);
nor U2347 (N_2347,N_1905,N_1635);
xor U2348 (N_2348,N_1626,N_1894);
and U2349 (N_2349,N_1618,N_1891);
or U2350 (N_2350,N_1902,N_1675);
and U2351 (N_2351,N_1855,N_1829);
and U2352 (N_2352,N_1894,N_1778);
nor U2353 (N_2353,N_1773,N_1615);
nand U2354 (N_2354,N_1683,N_1672);
and U2355 (N_2355,N_1903,N_1843);
and U2356 (N_2356,N_1981,N_1705);
nor U2357 (N_2357,N_1989,N_1800);
or U2358 (N_2358,N_1740,N_1844);
xnor U2359 (N_2359,N_1779,N_1663);
nor U2360 (N_2360,N_1823,N_1627);
and U2361 (N_2361,N_1737,N_1760);
nand U2362 (N_2362,N_1763,N_1766);
and U2363 (N_2363,N_1956,N_1803);
nor U2364 (N_2364,N_1832,N_1669);
and U2365 (N_2365,N_1699,N_1807);
or U2366 (N_2366,N_1749,N_1845);
nand U2367 (N_2367,N_1867,N_1870);
and U2368 (N_2368,N_1832,N_1891);
and U2369 (N_2369,N_1616,N_1765);
and U2370 (N_2370,N_1661,N_1992);
nand U2371 (N_2371,N_1911,N_1830);
nand U2372 (N_2372,N_1991,N_1634);
nor U2373 (N_2373,N_1979,N_1782);
xnor U2374 (N_2374,N_1794,N_1843);
or U2375 (N_2375,N_1686,N_1877);
xor U2376 (N_2376,N_1951,N_1740);
nand U2377 (N_2377,N_1729,N_1806);
nand U2378 (N_2378,N_1640,N_1738);
and U2379 (N_2379,N_1931,N_1870);
and U2380 (N_2380,N_1783,N_1831);
xnor U2381 (N_2381,N_1802,N_1866);
and U2382 (N_2382,N_1917,N_1872);
or U2383 (N_2383,N_1957,N_1866);
and U2384 (N_2384,N_1838,N_1771);
xor U2385 (N_2385,N_1604,N_1815);
nand U2386 (N_2386,N_1886,N_1705);
nand U2387 (N_2387,N_1910,N_1909);
or U2388 (N_2388,N_1848,N_1694);
and U2389 (N_2389,N_1811,N_1687);
and U2390 (N_2390,N_1963,N_1968);
and U2391 (N_2391,N_1858,N_1970);
nand U2392 (N_2392,N_1677,N_1929);
or U2393 (N_2393,N_1941,N_1749);
nor U2394 (N_2394,N_1690,N_1876);
nor U2395 (N_2395,N_1682,N_1799);
nand U2396 (N_2396,N_1704,N_1910);
nor U2397 (N_2397,N_1892,N_1744);
and U2398 (N_2398,N_1612,N_1793);
nor U2399 (N_2399,N_1782,N_1846);
nor U2400 (N_2400,N_2251,N_2127);
and U2401 (N_2401,N_2057,N_2096);
nor U2402 (N_2402,N_2001,N_2334);
xor U2403 (N_2403,N_2182,N_2067);
nand U2404 (N_2404,N_2044,N_2064);
nor U2405 (N_2405,N_2019,N_2119);
nor U2406 (N_2406,N_2071,N_2260);
or U2407 (N_2407,N_2364,N_2207);
and U2408 (N_2408,N_2295,N_2277);
nor U2409 (N_2409,N_2206,N_2314);
or U2410 (N_2410,N_2220,N_2125);
nor U2411 (N_2411,N_2023,N_2013);
nand U2412 (N_2412,N_2045,N_2035);
and U2413 (N_2413,N_2340,N_2323);
and U2414 (N_2414,N_2238,N_2253);
and U2415 (N_2415,N_2075,N_2215);
nand U2416 (N_2416,N_2326,N_2050);
or U2417 (N_2417,N_2192,N_2305);
and U2418 (N_2418,N_2382,N_2298);
and U2419 (N_2419,N_2136,N_2068);
nor U2420 (N_2420,N_2325,N_2353);
and U2421 (N_2421,N_2155,N_2357);
and U2422 (N_2422,N_2370,N_2210);
nand U2423 (N_2423,N_2093,N_2331);
nor U2424 (N_2424,N_2265,N_2299);
nand U2425 (N_2425,N_2065,N_2287);
nor U2426 (N_2426,N_2386,N_2002);
and U2427 (N_2427,N_2393,N_2072);
or U2428 (N_2428,N_2313,N_2154);
xor U2429 (N_2429,N_2367,N_2303);
and U2430 (N_2430,N_2095,N_2279);
nand U2431 (N_2431,N_2368,N_2244);
or U2432 (N_2432,N_2134,N_2015);
xor U2433 (N_2433,N_2389,N_2376);
nor U2434 (N_2434,N_2232,N_2229);
xnor U2435 (N_2435,N_2103,N_2297);
or U2436 (N_2436,N_2217,N_2166);
xor U2437 (N_2437,N_2214,N_2087);
xnor U2438 (N_2438,N_2219,N_2234);
or U2439 (N_2439,N_2077,N_2117);
or U2440 (N_2440,N_2165,N_2373);
and U2441 (N_2441,N_2324,N_2026);
or U2442 (N_2442,N_2145,N_2218);
nand U2443 (N_2443,N_2164,N_2131);
nor U2444 (N_2444,N_2092,N_2054);
nor U2445 (N_2445,N_2375,N_2167);
nor U2446 (N_2446,N_2129,N_2395);
nand U2447 (N_2447,N_2080,N_2171);
nor U2448 (N_2448,N_2174,N_2098);
and U2449 (N_2449,N_2085,N_2014);
nand U2450 (N_2450,N_2149,N_2342);
or U2451 (N_2451,N_2005,N_2390);
nor U2452 (N_2452,N_2181,N_2073);
xnor U2453 (N_2453,N_2038,N_2300);
and U2454 (N_2454,N_2350,N_2000);
nand U2455 (N_2455,N_2285,N_2255);
and U2456 (N_2456,N_2027,N_2309);
xor U2457 (N_2457,N_2090,N_2320);
or U2458 (N_2458,N_2004,N_2282);
nor U2459 (N_2459,N_2191,N_2256);
or U2460 (N_2460,N_2083,N_2335);
nand U2461 (N_2461,N_2036,N_2147);
and U2462 (N_2462,N_2337,N_2143);
nor U2463 (N_2463,N_2017,N_2222);
nand U2464 (N_2464,N_2058,N_2195);
or U2465 (N_2465,N_2094,N_2341);
nand U2466 (N_2466,N_2158,N_2345);
or U2467 (N_2467,N_2359,N_2043);
nand U2468 (N_2468,N_2223,N_2266);
or U2469 (N_2469,N_2268,N_2230);
xor U2470 (N_2470,N_2264,N_2152);
and U2471 (N_2471,N_2120,N_2258);
xor U2472 (N_2472,N_2193,N_2302);
nand U2473 (N_2473,N_2304,N_2076);
nor U2474 (N_2474,N_2184,N_2024);
xnor U2475 (N_2475,N_2235,N_2301);
or U2476 (N_2476,N_2040,N_2059);
nor U2477 (N_2477,N_2063,N_2025);
or U2478 (N_2478,N_2237,N_2208);
and U2479 (N_2479,N_2316,N_2037);
nor U2480 (N_2480,N_2248,N_2088);
xor U2481 (N_2481,N_2079,N_2257);
or U2482 (N_2482,N_2178,N_2346);
xor U2483 (N_2483,N_2197,N_2365);
or U2484 (N_2484,N_2204,N_2113);
nand U2485 (N_2485,N_2306,N_2396);
and U2486 (N_2486,N_2159,N_2042);
xor U2487 (N_2487,N_2176,N_2332);
xnor U2488 (N_2488,N_2006,N_2212);
and U2489 (N_2489,N_2273,N_2362);
nor U2490 (N_2490,N_2078,N_2126);
or U2491 (N_2491,N_2318,N_2189);
nor U2492 (N_2492,N_2275,N_2209);
or U2493 (N_2493,N_2137,N_2177);
xor U2494 (N_2494,N_2007,N_2226);
nor U2495 (N_2495,N_2196,N_2378);
or U2496 (N_2496,N_2055,N_2199);
nand U2497 (N_2497,N_2116,N_2151);
nor U2498 (N_2498,N_2061,N_2211);
xnor U2499 (N_2499,N_2358,N_2106);
nor U2500 (N_2500,N_2122,N_2352);
or U2501 (N_2501,N_2089,N_2172);
and U2502 (N_2502,N_2239,N_2354);
xnor U2503 (N_2503,N_2377,N_2246);
nor U2504 (N_2504,N_2046,N_2278);
or U2505 (N_2505,N_2105,N_2101);
and U2506 (N_2506,N_2049,N_2289);
and U2507 (N_2507,N_2292,N_2086);
and U2508 (N_2508,N_2082,N_2010);
or U2509 (N_2509,N_2141,N_2188);
nand U2510 (N_2510,N_2062,N_2018);
nor U2511 (N_2511,N_2236,N_2311);
and U2512 (N_2512,N_2020,N_2048);
nor U2513 (N_2513,N_2163,N_2100);
or U2514 (N_2514,N_2109,N_2274);
nand U2515 (N_2515,N_2319,N_2271);
xnor U2516 (N_2516,N_2081,N_2240);
nor U2517 (N_2517,N_2228,N_2112);
nand U2518 (N_2518,N_2021,N_2203);
nand U2519 (N_2519,N_2130,N_2333);
nor U2520 (N_2520,N_2392,N_2315);
nand U2521 (N_2521,N_2347,N_2329);
nand U2522 (N_2522,N_2132,N_2138);
nor U2523 (N_2523,N_2280,N_2241);
nor U2524 (N_2524,N_2388,N_2157);
or U2525 (N_2525,N_2121,N_2231);
or U2526 (N_2526,N_2254,N_2194);
xnor U2527 (N_2527,N_2286,N_2374);
nor U2528 (N_2528,N_2224,N_2307);
nor U2529 (N_2529,N_2011,N_2221);
nand U2530 (N_2530,N_2108,N_2183);
xnor U2531 (N_2531,N_2169,N_2162);
and U2532 (N_2532,N_2160,N_2385);
or U2533 (N_2533,N_2366,N_2028);
or U2534 (N_2534,N_2270,N_2327);
xnor U2535 (N_2535,N_2102,N_2139);
xnor U2536 (N_2536,N_2281,N_2016);
and U2537 (N_2537,N_2118,N_2186);
and U2538 (N_2538,N_2115,N_2371);
nor U2539 (N_2539,N_2262,N_2384);
nand U2540 (N_2540,N_2267,N_2198);
and U2541 (N_2541,N_2175,N_2110);
nand U2542 (N_2542,N_2276,N_2394);
nand U2543 (N_2543,N_2124,N_2259);
nand U2544 (N_2544,N_2107,N_2336);
nand U2545 (N_2545,N_2012,N_2069);
and U2546 (N_2546,N_2047,N_2030);
or U2547 (N_2547,N_2097,N_2247);
nand U2548 (N_2548,N_2104,N_2056);
xor U2549 (N_2549,N_2363,N_2070);
or U2550 (N_2550,N_2140,N_2312);
and U2551 (N_2551,N_2387,N_2156);
nand U2552 (N_2552,N_2170,N_2032);
and U2553 (N_2553,N_2201,N_2398);
and U2554 (N_2554,N_2216,N_2084);
nor U2555 (N_2555,N_2243,N_2269);
xor U2556 (N_2556,N_2344,N_2383);
or U2557 (N_2557,N_2009,N_2135);
and U2558 (N_2558,N_2074,N_2338);
or U2559 (N_2559,N_2294,N_2272);
nand U2560 (N_2560,N_2252,N_2379);
or U2561 (N_2561,N_2039,N_2200);
or U2562 (N_2562,N_2249,N_2008);
nor U2563 (N_2563,N_2291,N_2099);
and U2564 (N_2564,N_2052,N_2111);
and U2565 (N_2565,N_2351,N_2205);
nor U2566 (N_2566,N_2356,N_2242);
and U2567 (N_2567,N_2369,N_2187);
and U2568 (N_2568,N_2173,N_2399);
or U2569 (N_2569,N_2033,N_2148);
nor U2570 (N_2570,N_2202,N_2348);
and U2571 (N_2571,N_2361,N_2179);
or U2572 (N_2572,N_2168,N_2322);
nand U2573 (N_2573,N_2381,N_2308);
nand U2574 (N_2574,N_2293,N_2128);
nor U2575 (N_2575,N_2330,N_2190);
nor U2576 (N_2576,N_2034,N_2284);
nor U2577 (N_2577,N_2349,N_2343);
xor U2578 (N_2578,N_2060,N_2360);
nand U2579 (N_2579,N_2161,N_2029);
nor U2580 (N_2580,N_2031,N_2397);
xor U2581 (N_2581,N_2317,N_2051);
nor U2582 (N_2582,N_2144,N_2261);
or U2583 (N_2583,N_2142,N_2123);
and U2584 (N_2584,N_2022,N_2233);
nor U2585 (N_2585,N_2372,N_2225);
or U2586 (N_2586,N_2146,N_2283);
and U2587 (N_2587,N_2355,N_2321);
nor U2588 (N_2588,N_2213,N_2185);
xnor U2589 (N_2589,N_2091,N_2133);
and U2590 (N_2590,N_2288,N_2290);
nand U2591 (N_2591,N_2227,N_2180);
or U2592 (N_2592,N_2114,N_2310);
xor U2593 (N_2593,N_2053,N_2153);
nor U2594 (N_2594,N_2328,N_2250);
and U2595 (N_2595,N_2003,N_2150);
or U2596 (N_2596,N_2380,N_2245);
or U2597 (N_2597,N_2296,N_2339);
xnor U2598 (N_2598,N_2066,N_2391);
nor U2599 (N_2599,N_2041,N_2263);
and U2600 (N_2600,N_2187,N_2184);
xnor U2601 (N_2601,N_2116,N_2287);
nand U2602 (N_2602,N_2189,N_2296);
nand U2603 (N_2603,N_2313,N_2103);
xor U2604 (N_2604,N_2341,N_2180);
xor U2605 (N_2605,N_2198,N_2049);
xnor U2606 (N_2606,N_2186,N_2153);
xnor U2607 (N_2607,N_2065,N_2308);
nand U2608 (N_2608,N_2382,N_2098);
nand U2609 (N_2609,N_2132,N_2214);
xnor U2610 (N_2610,N_2065,N_2263);
nor U2611 (N_2611,N_2380,N_2362);
nand U2612 (N_2612,N_2353,N_2087);
xnor U2613 (N_2613,N_2235,N_2046);
xor U2614 (N_2614,N_2330,N_2127);
or U2615 (N_2615,N_2312,N_2064);
nor U2616 (N_2616,N_2243,N_2012);
and U2617 (N_2617,N_2146,N_2003);
nand U2618 (N_2618,N_2216,N_2201);
or U2619 (N_2619,N_2193,N_2274);
nor U2620 (N_2620,N_2091,N_2046);
xnor U2621 (N_2621,N_2083,N_2387);
xor U2622 (N_2622,N_2323,N_2035);
and U2623 (N_2623,N_2354,N_2228);
nand U2624 (N_2624,N_2086,N_2346);
nand U2625 (N_2625,N_2001,N_2379);
xnor U2626 (N_2626,N_2384,N_2398);
nand U2627 (N_2627,N_2377,N_2375);
xnor U2628 (N_2628,N_2054,N_2183);
and U2629 (N_2629,N_2086,N_2080);
xnor U2630 (N_2630,N_2173,N_2058);
xor U2631 (N_2631,N_2309,N_2058);
or U2632 (N_2632,N_2269,N_2085);
xor U2633 (N_2633,N_2112,N_2150);
or U2634 (N_2634,N_2069,N_2293);
and U2635 (N_2635,N_2069,N_2295);
nand U2636 (N_2636,N_2061,N_2052);
nor U2637 (N_2637,N_2324,N_2097);
nor U2638 (N_2638,N_2269,N_2072);
and U2639 (N_2639,N_2160,N_2113);
nor U2640 (N_2640,N_2283,N_2233);
or U2641 (N_2641,N_2333,N_2092);
xnor U2642 (N_2642,N_2090,N_2316);
and U2643 (N_2643,N_2286,N_2204);
or U2644 (N_2644,N_2074,N_2108);
nor U2645 (N_2645,N_2077,N_2203);
xor U2646 (N_2646,N_2059,N_2027);
xor U2647 (N_2647,N_2189,N_2172);
and U2648 (N_2648,N_2005,N_2251);
nand U2649 (N_2649,N_2104,N_2022);
or U2650 (N_2650,N_2142,N_2361);
xor U2651 (N_2651,N_2102,N_2152);
xnor U2652 (N_2652,N_2042,N_2177);
nand U2653 (N_2653,N_2043,N_2259);
xnor U2654 (N_2654,N_2397,N_2051);
and U2655 (N_2655,N_2052,N_2114);
xnor U2656 (N_2656,N_2192,N_2376);
xor U2657 (N_2657,N_2337,N_2346);
or U2658 (N_2658,N_2127,N_2157);
nand U2659 (N_2659,N_2235,N_2335);
and U2660 (N_2660,N_2277,N_2368);
nand U2661 (N_2661,N_2086,N_2095);
and U2662 (N_2662,N_2184,N_2099);
and U2663 (N_2663,N_2160,N_2174);
or U2664 (N_2664,N_2152,N_2114);
and U2665 (N_2665,N_2179,N_2157);
xnor U2666 (N_2666,N_2382,N_2019);
nor U2667 (N_2667,N_2264,N_2386);
or U2668 (N_2668,N_2344,N_2063);
xnor U2669 (N_2669,N_2027,N_2293);
or U2670 (N_2670,N_2149,N_2161);
nor U2671 (N_2671,N_2011,N_2134);
or U2672 (N_2672,N_2186,N_2028);
nor U2673 (N_2673,N_2139,N_2170);
and U2674 (N_2674,N_2334,N_2005);
and U2675 (N_2675,N_2029,N_2238);
nor U2676 (N_2676,N_2053,N_2107);
nor U2677 (N_2677,N_2135,N_2132);
and U2678 (N_2678,N_2141,N_2080);
nor U2679 (N_2679,N_2111,N_2195);
xnor U2680 (N_2680,N_2008,N_2269);
nor U2681 (N_2681,N_2109,N_2087);
xnor U2682 (N_2682,N_2148,N_2248);
and U2683 (N_2683,N_2223,N_2037);
nor U2684 (N_2684,N_2338,N_2354);
and U2685 (N_2685,N_2051,N_2114);
nor U2686 (N_2686,N_2254,N_2097);
or U2687 (N_2687,N_2031,N_2220);
or U2688 (N_2688,N_2332,N_2266);
nor U2689 (N_2689,N_2281,N_2048);
and U2690 (N_2690,N_2221,N_2371);
nand U2691 (N_2691,N_2369,N_2085);
nor U2692 (N_2692,N_2203,N_2269);
and U2693 (N_2693,N_2217,N_2120);
xor U2694 (N_2694,N_2270,N_2062);
nor U2695 (N_2695,N_2125,N_2368);
nand U2696 (N_2696,N_2224,N_2328);
nor U2697 (N_2697,N_2054,N_2038);
or U2698 (N_2698,N_2265,N_2011);
and U2699 (N_2699,N_2289,N_2148);
nor U2700 (N_2700,N_2335,N_2023);
nor U2701 (N_2701,N_2120,N_2068);
xnor U2702 (N_2702,N_2383,N_2047);
or U2703 (N_2703,N_2008,N_2044);
or U2704 (N_2704,N_2322,N_2226);
and U2705 (N_2705,N_2015,N_2227);
or U2706 (N_2706,N_2254,N_2102);
xor U2707 (N_2707,N_2207,N_2336);
nor U2708 (N_2708,N_2194,N_2038);
or U2709 (N_2709,N_2229,N_2150);
or U2710 (N_2710,N_2304,N_2325);
nand U2711 (N_2711,N_2203,N_2043);
or U2712 (N_2712,N_2304,N_2251);
nand U2713 (N_2713,N_2068,N_2053);
nor U2714 (N_2714,N_2168,N_2289);
xor U2715 (N_2715,N_2313,N_2353);
nor U2716 (N_2716,N_2107,N_2297);
nor U2717 (N_2717,N_2272,N_2285);
nand U2718 (N_2718,N_2182,N_2021);
nand U2719 (N_2719,N_2089,N_2278);
nor U2720 (N_2720,N_2310,N_2008);
nand U2721 (N_2721,N_2133,N_2311);
xor U2722 (N_2722,N_2061,N_2175);
and U2723 (N_2723,N_2267,N_2322);
nor U2724 (N_2724,N_2378,N_2030);
xor U2725 (N_2725,N_2372,N_2349);
nand U2726 (N_2726,N_2137,N_2046);
and U2727 (N_2727,N_2244,N_2000);
xor U2728 (N_2728,N_2262,N_2046);
xnor U2729 (N_2729,N_2110,N_2099);
xor U2730 (N_2730,N_2020,N_2170);
nor U2731 (N_2731,N_2240,N_2396);
xnor U2732 (N_2732,N_2061,N_2091);
and U2733 (N_2733,N_2038,N_2395);
nor U2734 (N_2734,N_2303,N_2386);
xnor U2735 (N_2735,N_2358,N_2323);
and U2736 (N_2736,N_2356,N_2148);
nor U2737 (N_2737,N_2250,N_2393);
xor U2738 (N_2738,N_2282,N_2310);
xor U2739 (N_2739,N_2281,N_2389);
and U2740 (N_2740,N_2136,N_2222);
or U2741 (N_2741,N_2203,N_2333);
and U2742 (N_2742,N_2339,N_2039);
or U2743 (N_2743,N_2042,N_2007);
nand U2744 (N_2744,N_2280,N_2131);
and U2745 (N_2745,N_2067,N_2295);
nor U2746 (N_2746,N_2109,N_2102);
nor U2747 (N_2747,N_2299,N_2365);
and U2748 (N_2748,N_2276,N_2025);
xnor U2749 (N_2749,N_2340,N_2284);
or U2750 (N_2750,N_2309,N_2259);
nand U2751 (N_2751,N_2390,N_2149);
and U2752 (N_2752,N_2161,N_2200);
xnor U2753 (N_2753,N_2386,N_2015);
nor U2754 (N_2754,N_2190,N_2168);
or U2755 (N_2755,N_2182,N_2072);
xnor U2756 (N_2756,N_2270,N_2129);
nand U2757 (N_2757,N_2212,N_2029);
nor U2758 (N_2758,N_2252,N_2176);
and U2759 (N_2759,N_2196,N_2153);
nor U2760 (N_2760,N_2104,N_2210);
nor U2761 (N_2761,N_2215,N_2347);
xor U2762 (N_2762,N_2330,N_2151);
and U2763 (N_2763,N_2260,N_2085);
nand U2764 (N_2764,N_2207,N_2236);
nand U2765 (N_2765,N_2286,N_2135);
xnor U2766 (N_2766,N_2132,N_2043);
nand U2767 (N_2767,N_2238,N_2154);
nor U2768 (N_2768,N_2010,N_2084);
nor U2769 (N_2769,N_2064,N_2018);
xor U2770 (N_2770,N_2247,N_2103);
xnor U2771 (N_2771,N_2126,N_2164);
xnor U2772 (N_2772,N_2234,N_2023);
and U2773 (N_2773,N_2375,N_2280);
xor U2774 (N_2774,N_2326,N_2013);
nand U2775 (N_2775,N_2262,N_2313);
and U2776 (N_2776,N_2161,N_2081);
nand U2777 (N_2777,N_2150,N_2278);
or U2778 (N_2778,N_2065,N_2382);
nand U2779 (N_2779,N_2149,N_2132);
and U2780 (N_2780,N_2236,N_2322);
or U2781 (N_2781,N_2262,N_2094);
xnor U2782 (N_2782,N_2055,N_2306);
nand U2783 (N_2783,N_2068,N_2192);
and U2784 (N_2784,N_2002,N_2106);
or U2785 (N_2785,N_2029,N_2305);
xnor U2786 (N_2786,N_2218,N_2229);
or U2787 (N_2787,N_2168,N_2158);
nand U2788 (N_2788,N_2018,N_2236);
nand U2789 (N_2789,N_2020,N_2208);
xor U2790 (N_2790,N_2367,N_2006);
nand U2791 (N_2791,N_2198,N_2300);
nand U2792 (N_2792,N_2084,N_2267);
nor U2793 (N_2793,N_2225,N_2067);
and U2794 (N_2794,N_2260,N_2190);
nor U2795 (N_2795,N_2389,N_2367);
xor U2796 (N_2796,N_2237,N_2027);
and U2797 (N_2797,N_2111,N_2304);
xnor U2798 (N_2798,N_2137,N_2289);
and U2799 (N_2799,N_2101,N_2196);
and U2800 (N_2800,N_2537,N_2559);
nor U2801 (N_2801,N_2725,N_2628);
xnor U2802 (N_2802,N_2756,N_2616);
nor U2803 (N_2803,N_2498,N_2463);
or U2804 (N_2804,N_2694,N_2752);
and U2805 (N_2805,N_2760,N_2609);
or U2806 (N_2806,N_2758,N_2736);
and U2807 (N_2807,N_2768,N_2749);
xor U2808 (N_2808,N_2702,N_2605);
and U2809 (N_2809,N_2792,N_2751);
nor U2810 (N_2810,N_2481,N_2594);
nor U2811 (N_2811,N_2447,N_2483);
nor U2812 (N_2812,N_2429,N_2693);
nor U2813 (N_2813,N_2545,N_2626);
and U2814 (N_2814,N_2610,N_2458);
xor U2815 (N_2815,N_2492,N_2524);
nor U2816 (N_2816,N_2465,N_2689);
nand U2817 (N_2817,N_2477,N_2421);
nand U2818 (N_2818,N_2419,N_2434);
and U2819 (N_2819,N_2522,N_2620);
and U2820 (N_2820,N_2675,N_2454);
nand U2821 (N_2821,N_2474,N_2427);
xnor U2822 (N_2822,N_2707,N_2523);
nor U2823 (N_2823,N_2517,N_2782);
or U2824 (N_2824,N_2645,N_2794);
xor U2825 (N_2825,N_2512,N_2568);
and U2826 (N_2826,N_2646,N_2740);
or U2827 (N_2827,N_2491,N_2406);
and U2828 (N_2828,N_2764,N_2676);
or U2829 (N_2829,N_2759,N_2569);
xor U2830 (N_2830,N_2667,N_2437);
xnor U2831 (N_2831,N_2402,N_2521);
nand U2832 (N_2832,N_2453,N_2621);
nand U2833 (N_2833,N_2767,N_2473);
xnor U2834 (N_2834,N_2542,N_2634);
xor U2835 (N_2835,N_2507,N_2556);
nor U2836 (N_2836,N_2573,N_2576);
nor U2837 (N_2837,N_2662,N_2661);
xnor U2838 (N_2838,N_2600,N_2433);
xnor U2839 (N_2839,N_2618,N_2533);
or U2840 (N_2840,N_2709,N_2684);
xnor U2841 (N_2841,N_2774,N_2765);
nand U2842 (N_2842,N_2485,N_2452);
xor U2843 (N_2843,N_2762,N_2753);
and U2844 (N_2844,N_2698,N_2670);
nand U2845 (N_2845,N_2510,N_2410);
and U2846 (N_2846,N_2435,N_2557);
nand U2847 (N_2847,N_2722,N_2497);
xor U2848 (N_2848,N_2478,N_2417);
xnor U2849 (N_2849,N_2641,N_2532);
xnor U2850 (N_2850,N_2459,N_2785);
xnor U2851 (N_2851,N_2549,N_2494);
nand U2852 (N_2852,N_2595,N_2401);
nor U2853 (N_2853,N_2691,N_2450);
and U2854 (N_2854,N_2598,N_2743);
or U2855 (N_2855,N_2688,N_2761);
and U2856 (N_2856,N_2627,N_2731);
or U2857 (N_2857,N_2713,N_2791);
or U2858 (N_2858,N_2674,N_2490);
or U2859 (N_2859,N_2516,N_2714);
xor U2860 (N_2860,N_2565,N_2416);
nor U2861 (N_2861,N_2505,N_2680);
or U2862 (N_2862,N_2581,N_2747);
nand U2863 (N_2863,N_2525,N_2509);
and U2864 (N_2864,N_2672,N_2701);
or U2865 (N_2865,N_2639,N_2415);
or U2866 (N_2866,N_2708,N_2527);
xor U2867 (N_2867,N_2658,N_2487);
nand U2868 (N_2868,N_2718,N_2504);
nor U2869 (N_2869,N_2561,N_2738);
and U2870 (N_2870,N_2480,N_2467);
nor U2871 (N_2871,N_2409,N_2783);
and U2872 (N_2872,N_2440,N_2717);
nor U2873 (N_2873,N_2563,N_2624);
and U2874 (N_2874,N_2457,N_2651);
nor U2875 (N_2875,N_2597,N_2750);
or U2876 (N_2876,N_2479,N_2536);
nor U2877 (N_2877,N_2786,N_2404);
xnor U2878 (N_2878,N_2547,N_2793);
nand U2879 (N_2879,N_2499,N_2574);
xor U2880 (N_2880,N_2625,N_2766);
nand U2881 (N_2881,N_2654,N_2660);
nand U2882 (N_2882,N_2408,N_2629);
nand U2883 (N_2883,N_2413,N_2789);
or U2884 (N_2884,N_2451,N_2471);
nand U2885 (N_2885,N_2704,N_2682);
or U2886 (N_2886,N_2461,N_2443);
nor U2887 (N_2887,N_2608,N_2588);
nand U2888 (N_2888,N_2612,N_2712);
and U2889 (N_2889,N_2486,N_2601);
and U2890 (N_2890,N_2687,N_2585);
and U2891 (N_2891,N_2548,N_2772);
xor U2892 (N_2892,N_2613,N_2464);
nand U2893 (N_2893,N_2664,N_2622);
and U2894 (N_2894,N_2703,N_2795);
nor U2895 (N_2895,N_2614,N_2784);
xnor U2896 (N_2896,N_2649,N_2446);
nand U2897 (N_2897,N_2679,N_2528);
and U2898 (N_2898,N_2403,N_2518);
and U2899 (N_2899,N_2539,N_2638);
and U2900 (N_2900,N_2721,N_2636);
nor U2901 (N_2901,N_2754,N_2642);
nand U2902 (N_2902,N_2592,N_2673);
and U2903 (N_2903,N_2432,N_2666);
and U2904 (N_2904,N_2602,N_2445);
or U2905 (N_2905,N_2583,N_2637);
nor U2906 (N_2906,N_2551,N_2781);
or U2907 (N_2907,N_2554,N_2790);
xnor U2908 (N_2908,N_2582,N_2650);
nor U2909 (N_2909,N_2733,N_2562);
nand U2910 (N_2910,N_2630,N_2719);
nor U2911 (N_2911,N_2570,N_2644);
xor U2912 (N_2912,N_2534,N_2449);
nand U2913 (N_2913,N_2502,N_2773);
or U2914 (N_2914,N_2729,N_2577);
and U2915 (N_2915,N_2716,N_2411);
and U2916 (N_2916,N_2705,N_2572);
nor U2917 (N_2917,N_2737,N_2586);
nand U2918 (N_2918,N_2739,N_2423);
or U2919 (N_2919,N_2631,N_2500);
xnor U2920 (N_2920,N_2476,N_2589);
nand U2921 (N_2921,N_2466,N_2599);
xor U2922 (N_2922,N_2770,N_2558);
or U2923 (N_2923,N_2414,N_2787);
or U2924 (N_2924,N_2441,N_2428);
nand U2925 (N_2925,N_2635,N_2697);
and U2926 (N_2926,N_2741,N_2696);
and U2927 (N_2927,N_2734,N_2550);
nor U2928 (N_2928,N_2514,N_2615);
and U2929 (N_2929,N_2515,N_2460);
or U2930 (N_2930,N_2438,N_2796);
and U2931 (N_2931,N_2724,N_2643);
nand U2932 (N_2932,N_2591,N_2665);
nand U2933 (N_2933,N_2555,N_2677);
nand U2934 (N_2934,N_2678,N_2590);
xnor U2935 (N_2935,N_2617,N_2671);
xor U2936 (N_2936,N_2543,N_2611);
nor U2937 (N_2937,N_2744,N_2775);
xnor U2938 (N_2938,N_2526,N_2412);
and U2939 (N_2939,N_2560,N_2779);
and U2940 (N_2940,N_2400,N_2771);
and U2941 (N_2941,N_2553,N_2407);
nor U2942 (N_2942,N_2567,N_2720);
nor U2943 (N_2943,N_2493,N_2587);
nor U2944 (N_2944,N_2552,N_2640);
nand U2945 (N_2945,N_2462,N_2788);
xor U2946 (N_2946,N_2619,N_2439);
nand U2947 (N_2947,N_2541,N_2706);
xor U2948 (N_2948,N_2578,N_2520);
xor U2949 (N_2949,N_2746,N_2424);
or U2950 (N_2950,N_2444,N_2663);
and U2951 (N_2951,N_2659,N_2531);
or U2952 (N_2952,N_2472,N_2436);
xnor U2953 (N_2953,N_2544,N_2503);
or U2954 (N_2954,N_2727,N_2495);
or U2955 (N_2955,N_2657,N_2603);
and U2956 (N_2956,N_2763,N_2575);
nand U2957 (N_2957,N_2695,N_2469);
xor U2958 (N_2958,N_2606,N_2732);
nand U2959 (N_2959,N_2777,N_2797);
xor U2960 (N_2960,N_2431,N_2632);
nor U2961 (N_2961,N_2593,N_2692);
nor U2962 (N_2962,N_2425,N_2726);
nor U2963 (N_2963,N_2699,N_2508);
or U2964 (N_2964,N_2669,N_2535);
xnor U2965 (N_2965,N_2604,N_2776);
nand U2966 (N_2966,N_2488,N_2668);
and U2967 (N_2967,N_2579,N_2470);
and U2968 (N_2968,N_2418,N_2420);
nor U2969 (N_2969,N_2540,N_2489);
and U2970 (N_2970,N_2580,N_2501);
nor U2971 (N_2971,N_2506,N_2648);
or U2972 (N_2972,N_2455,N_2571);
xnor U2973 (N_2973,N_2742,N_2584);
or U2974 (N_2974,N_2513,N_2530);
nand U2975 (N_2975,N_2799,N_2769);
xnor U2976 (N_2976,N_2728,N_2442);
nand U2977 (N_2977,N_2652,N_2538);
or U2978 (N_2978,N_2656,N_2730);
or U2979 (N_2979,N_2685,N_2633);
xnor U2980 (N_2980,N_2647,N_2426);
nand U2981 (N_2981,N_2405,N_2482);
nor U2982 (N_2982,N_2422,N_2715);
nor U2983 (N_2983,N_2683,N_2519);
nand U2984 (N_2984,N_2484,N_2700);
and U2985 (N_2985,N_2757,N_2566);
xnor U2986 (N_2986,N_2745,N_2798);
or U2987 (N_2987,N_2529,N_2546);
or U2988 (N_2988,N_2755,N_2430);
nand U2989 (N_2989,N_2686,N_2456);
or U2990 (N_2990,N_2448,N_2723);
and U2991 (N_2991,N_2653,N_2690);
nand U2992 (N_2992,N_2511,N_2475);
nor U2993 (N_2993,N_2681,N_2711);
or U2994 (N_2994,N_2780,N_2748);
nand U2995 (N_2995,N_2710,N_2778);
nor U2996 (N_2996,N_2564,N_2468);
xor U2997 (N_2997,N_2655,N_2735);
nand U2998 (N_2998,N_2623,N_2596);
nand U2999 (N_2999,N_2607,N_2496);
nand U3000 (N_3000,N_2549,N_2634);
nor U3001 (N_3001,N_2675,N_2440);
and U3002 (N_3002,N_2700,N_2561);
nand U3003 (N_3003,N_2531,N_2526);
nand U3004 (N_3004,N_2500,N_2527);
xor U3005 (N_3005,N_2680,N_2755);
nor U3006 (N_3006,N_2618,N_2792);
xnor U3007 (N_3007,N_2502,N_2582);
or U3008 (N_3008,N_2527,N_2675);
or U3009 (N_3009,N_2764,N_2695);
nand U3010 (N_3010,N_2654,N_2778);
and U3011 (N_3011,N_2479,N_2475);
and U3012 (N_3012,N_2687,N_2633);
nor U3013 (N_3013,N_2574,N_2534);
nand U3014 (N_3014,N_2727,N_2493);
xnor U3015 (N_3015,N_2451,N_2550);
nor U3016 (N_3016,N_2610,N_2511);
nor U3017 (N_3017,N_2522,N_2564);
or U3018 (N_3018,N_2757,N_2565);
nand U3019 (N_3019,N_2514,N_2461);
nand U3020 (N_3020,N_2747,N_2692);
nand U3021 (N_3021,N_2559,N_2487);
xor U3022 (N_3022,N_2465,N_2755);
nand U3023 (N_3023,N_2486,N_2675);
nor U3024 (N_3024,N_2659,N_2624);
and U3025 (N_3025,N_2664,N_2788);
nand U3026 (N_3026,N_2477,N_2666);
nand U3027 (N_3027,N_2472,N_2473);
nand U3028 (N_3028,N_2429,N_2469);
xor U3029 (N_3029,N_2577,N_2794);
nor U3030 (N_3030,N_2545,N_2738);
and U3031 (N_3031,N_2616,N_2628);
and U3032 (N_3032,N_2442,N_2410);
xor U3033 (N_3033,N_2627,N_2478);
xor U3034 (N_3034,N_2744,N_2785);
and U3035 (N_3035,N_2486,N_2506);
xnor U3036 (N_3036,N_2625,N_2485);
nand U3037 (N_3037,N_2730,N_2426);
and U3038 (N_3038,N_2516,N_2401);
nand U3039 (N_3039,N_2541,N_2650);
and U3040 (N_3040,N_2442,N_2691);
and U3041 (N_3041,N_2467,N_2677);
and U3042 (N_3042,N_2526,N_2728);
nor U3043 (N_3043,N_2511,N_2606);
or U3044 (N_3044,N_2438,N_2427);
or U3045 (N_3045,N_2768,N_2514);
or U3046 (N_3046,N_2461,N_2689);
or U3047 (N_3047,N_2463,N_2642);
or U3048 (N_3048,N_2728,N_2759);
or U3049 (N_3049,N_2462,N_2410);
xnor U3050 (N_3050,N_2672,N_2555);
xor U3051 (N_3051,N_2734,N_2501);
xnor U3052 (N_3052,N_2400,N_2538);
xnor U3053 (N_3053,N_2543,N_2659);
or U3054 (N_3054,N_2508,N_2456);
nor U3055 (N_3055,N_2557,N_2753);
nor U3056 (N_3056,N_2783,N_2797);
nor U3057 (N_3057,N_2737,N_2726);
and U3058 (N_3058,N_2733,N_2491);
xor U3059 (N_3059,N_2560,N_2487);
or U3060 (N_3060,N_2761,N_2522);
nor U3061 (N_3061,N_2661,N_2764);
xor U3062 (N_3062,N_2561,N_2478);
nand U3063 (N_3063,N_2573,N_2675);
or U3064 (N_3064,N_2626,N_2585);
or U3065 (N_3065,N_2717,N_2612);
xor U3066 (N_3066,N_2665,N_2695);
or U3067 (N_3067,N_2638,N_2469);
nor U3068 (N_3068,N_2512,N_2403);
nand U3069 (N_3069,N_2611,N_2513);
nand U3070 (N_3070,N_2470,N_2560);
nor U3071 (N_3071,N_2495,N_2779);
xnor U3072 (N_3072,N_2465,N_2717);
nor U3073 (N_3073,N_2659,N_2577);
or U3074 (N_3074,N_2720,N_2535);
or U3075 (N_3075,N_2577,N_2461);
nand U3076 (N_3076,N_2498,N_2468);
or U3077 (N_3077,N_2619,N_2620);
or U3078 (N_3078,N_2662,N_2412);
xor U3079 (N_3079,N_2605,N_2585);
or U3080 (N_3080,N_2495,N_2545);
and U3081 (N_3081,N_2554,N_2755);
nor U3082 (N_3082,N_2762,N_2522);
nor U3083 (N_3083,N_2680,N_2782);
nor U3084 (N_3084,N_2427,N_2434);
nand U3085 (N_3085,N_2403,N_2732);
nor U3086 (N_3086,N_2729,N_2462);
nand U3087 (N_3087,N_2459,N_2718);
nor U3088 (N_3088,N_2731,N_2599);
and U3089 (N_3089,N_2736,N_2756);
nand U3090 (N_3090,N_2708,N_2634);
xor U3091 (N_3091,N_2739,N_2778);
xnor U3092 (N_3092,N_2530,N_2622);
and U3093 (N_3093,N_2684,N_2743);
nor U3094 (N_3094,N_2403,N_2704);
xnor U3095 (N_3095,N_2717,N_2541);
and U3096 (N_3096,N_2454,N_2682);
or U3097 (N_3097,N_2492,N_2442);
or U3098 (N_3098,N_2550,N_2464);
nor U3099 (N_3099,N_2416,N_2707);
xnor U3100 (N_3100,N_2421,N_2570);
or U3101 (N_3101,N_2767,N_2406);
or U3102 (N_3102,N_2421,N_2696);
nor U3103 (N_3103,N_2678,N_2405);
xnor U3104 (N_3104,N_2766,N_2582);
or U3105 (N_3105,N_2715,N_2686);
nand U3106 (N_3106,N_2665,N_2766);
nand U3107 (N_3107,N_2632,N_2600);
and U3108 (N_3108,N_2783,N_2658);
nor U3109 (N_3109,N_2578,N_2582);
nor U3110 (N_3110,N_2511,N_2631);
or U3111 (N_3111,N_2634,N_2566);
nor U3112 (N_3112,N_2503,N_2479);
or U3113 (N_3113,N_2599,N_2682);
nand U3114 (N_3114,N_2639,N_2612);
nand U3115 (N_3115,N_2473,N_2510);
nand U3116 (N_3116,N_2657,N_2462);
xnor U3117 (N_3117,N_2720,N_2731);
or U3118 (N_3118,N_2525,N_2654);
nand U3119 (N_3119,N_2406,N_2550);
xnor U3120 (N_3120,N_2555,N_2618);
xor U3121 (N_3121,N_2530,N_2563);
nor U3122 (N_3122,N_2542,N_2606);
and U3123 (N_3123,N_2596,N_2614);
xnor U3124 (N_3124,N_2507,N_2746);
and U3125 (N_3125,N_2791,N_2567);
nand U3126 (N_3126,N_2665,N_2749);
xor U3127 (N_3127,N_2464,N_2483);
or U3128 (N_3128,N_2428,N_2481);
nand U3129 (N_3129,N_2723,N_2407);
xor U3130 (N_3130,N_2653,N_2461);
and U3131 (N_3131,N_2639,N_2504);
or U3132 (N_3132,N_2429,N_2493);
nor U3133 (N_3133,N_2477,N_2423);
xnor U3134 (N_3134,N_2442,N_2638);
and U3135 (N_3135,N_2447,N_2777);
nand U3136 (N_3136,N_2581,N_2436);
and U3137 (N_3137,N_2629,N_2497);
and U3138 (N_3138,N_2479,N_2612);
nor U3139 (N_3139,N_2479,N_2643);
nand U3140 (N_3140,N_2559,N_2776);
xnor U3141 (N_3141,N_2718,N_2426);
nand U3142 (N_3142,N_2774,N_2635);
and U3143 (N_3143,N_2487,N_2770);
and U3144 (N_3144,N_2536,N_2676);
or U3145 (N_3145,N_2530,N_2727);
xor U3146 (N_3146,N_2594,N_2619);
nand U3147 (N_3147,N_2419,N_2572);
and U3148 (N_3148,N_2512,N_2675);
and U3149 (N_3149,N_2672,N_2463);
nor U3150 (N_3150,N_2626,N_2692);
nor U3151 (N_3151,N_2475,N_2728);
xnor U3152 (N_3152,N_2471,N_2626);
xnor U3153 (N_3153,N_2438,N_2636);
and U3154 (N_3154,N_2794,N_2522);
nand U3155 (N_3155,N_2710,N_2579);
or U3156 (N_3156,N_2407,N_2604);
nand U3157 (N_3157,N_2439,N_2403);
xnor U3158 (N_3158,N_2451,N_2467);
or U3159 (N_3159,N_2434,N_2469);
nand U3160 (N_3160,N_2640,N_2644);
or U3161 (N_3161,N_2431,N_2576);
nor U3162 (N_3162,N_2673,N_2590);
nor U3163 (N_3163,N_2685,N_2519);
or U3164 (N_3164,N_2598,N_2531);
nand U3165 (N_3165,N_2540,N_2493);
xor U3166 (N_3166,N_2649,N_2434);
xnor U3167 (N_3167,N_2584,N_2738);
and U3168 (N_3168,N_2649,N_2792);
nand U3169 (N_3169,N_2661,N_2496);
xor U3170 (N_3170,N_2590,N_2459);
nand U3171 (N_3171,N_2757,N_2573);
xnor U3172 (N_3172,N_2419,N_2452);
xor U3173 (N_3173,N_2786,N_2739);
nor U3174 (N_3174,N_2722,N_2732);
or U3175 (N_3175,N_2569,N_2418);
nand U3176 (N_3176,N_2632,N_2525);
xor U3177 (N_3177,N_2407,N_2528);
nand U3178 (N_3178,N_2508,N_2729);
or U3179 (N_3179,N_2653,N_2720);
xnor U3180 (N_3180,N_2449,N_2487);
nand U3181 (N_3181,N_2788,N_2415);
nand U3182 (N_3182,N_2576,N_2772);
xnor U3183 (N_3183,N_2639,N_2749);
or U3184 (N_3184,N_2420,N_2724);
nand U3185 (N_3185,N_2437,N_2785);
or U3186 (N_3186,N_2432,N_2463);
and U3187 (N_3187,N_2495,N_2460);
or U3188 (N_3188,N_2517,N_2520);
xnor U3189 (N_3189,N_2476,N_2603);
or U3190 (N_3190,N_2687,N_2796);
nand U3191 (N_3191,N_2738,N_2656);
nand U3192 (N_3192,N_2592,N_2737);
and U3193 (N_3193,N_2677,N_2692);
xor U3194 (N_3194,N_2723,N_2468);
or U3195 (N_3195,N_2663,N_2431);
and U3196 (N_3196,N_2767,N_2414);
nand U3197 (N_3197,N_2752,N_2667);
xor U3198 (N_3198,N_2412,N_2675);
xnor U3199 (N_3199,N_2612,N_2413);
nor U3200 (N_3200,N_3097,N_3031);
nand U3201 (N_3201,N_3147,N_3002);
xor U3202 (N_3202,N_3039,N_2992);
and U3203 (N_3203,N_2895,N_2869);
xor U3204 (N_3204,N_3077,N_2945);
nor U3205 (N_3205,N_3128,N_2814);
xor U3206 (N_3206,N_2836,N_3114);
or U3207 (N_3207,N_2861,N_3119);
and U3208 (N_3208,N_3134,N_2952);
nor U3209 (N_3209,N_2975,N_2838);
or U3210 (N_3210,N_2829,N_3028);
xor U3211 (N_3211,N_2854,N_3071);
or U3212 (N_3212,N_2845,N_2976);
or U3213 (N_3213,N_3197,N_2894);
nand U3214 (N_3214,N_2913,N_2847);
xor U3215 (N_3215,N_3172,N_2928);
nand U3216 (N_3216,N_3030,N_2809);
or U3217 (N_3217,N_3116,N_2818);
nand U3218 (N_3218,N_2853,N_3088);
nand U3219 (N_3219,N_2973,N_3008);
xnor U3220 (N_3220,N_3064,N_3146);
and U3221 (N_3221,N_2817,N_3016);
xor U3222 (N_3222,N_3098,N_3100);
nor U3223 (N_3223,N_3165,N_3003);
and U3224 (N_3224,N_2848,N_2994);
nand U3225 (N_3225,N_3163,N_2984);
nor U3226 (N_3226,N_3032,N_2842);
nand U3227 (N_3227,N_3007,N_3140);
xnor U3228 (N_3228,N_3096,N_2939);
xnor U3229 (N_3229,N_3051,N_3173);
nand U3230 (N_3230,N_2918,N_3045);
and U3231 (N_3231,N_2806,N_2880);
xnor U3232 (N_3232,N_3168,N_3170);
xnor U3233 (N_3233,N_3084,N_2926);
or U3234 (N_3234,N_2942,N_3018);
nand U3235 (N_3235,N_3118,N_2911);
xnor U3236 (N_3236,N_2860,N_2832);
and U3237 (N_3237,N_2959,N_3179);
nor U3238 (N_3238,N_2866,N_2948);
nand U3239 (N_3239,N_2883,N_2999);
and U3240 (N_3240,N_3113,N_3171);
nor U3241 (N_3241,N_3136,N_3060);
or U3242 (N_3242,N_3117,N_3034);
or U3243 (N_3243,N_2953,N_3185);
xnor U3244 (N_3244,N_3042,N_2985);
and U3245 (N_3245,N_2901,N_3055);
and U3246 (N_3246,N_3001,N_2978);
nand U3247 (N_3247,N_2982,N_3157);
nor U3248 (N_3248,N_2937,N_2826);
and U3249 (N_3249,N_3017,N_3049);
or U3250 (N_3250,N_3063,N_2987);
nor U3251 (N_3251,N_3048,N_2864);
nand U3252 (N_3252,N_2872,N_3069);
or U3253 (N_3253,N_3065,N_2819);
nor U3254 (N_3254,N_3198,N_2950);
xor U3255 (N_3255,N_2882,N_2896);
xnor U3256 (N_3256,N_2962,N_2917);
and U3257 (N_3257,N_3152,N_2825);
nor U3258 (N_3258,N_3068,N_2892);
and U3259 (N_3259,N_2820,N_3075);
nor U3260 (N_3260,N_3059,N_3108);
nor U3261 (N_3261,N_3046,N_3036);
or U3262 (N_3262,N_3021,N_3133);
nand U3263 (N_3263,N_3043,N_2961);
or U3264 (N_3264,N_3109,N_2830);
nand U3265 (N_3265,N_2904,N_2824);
or U3266 (N_3266,N_2977,N_2803);
and U3267 (N_3267,N_2821,N_2972);
and U3268 (N_3268,N_3177,N_3105);
xnor U3269 (N_3269,N_3126,N_3131);
nand U3270 (N_3270,N_2859,N_2938);
and U3271 (N_3271,N_3085,N_2857);
nand U3272 (N_3272,N_3006,N_2890);
xnor U3273 (N_3273,N_2943,N_3111);
xor U3274 (N_3274,N_3190,N_3082);
nor U3275 (N_3275,N_2876,N_3101);
and U3276 (N_3276,N_2893,N_3011);
and U3277 (N_3277,N_2902,N_2899);
or U3278 (N_3278,N_3066,N_2989);
nor U3279 (N_3279,N_3089,N_2881);
xor U3280 (N_3280,N_3115,N_3141);
nand U3281 (N_3281,N_2931,N_2849);
and U3282 (N_3282,N_2967,N_2908);
xnor U3283 (N_3283,N_3103,N_2903);
and U3284 (N_3284,N_2960,N_2851);
xnor U3285 (N_3285,N_3005,N_3073);
nor U3286 (N_3286,N_3056,N_2879);
xor U3287 (N_3287,N_3015,N_3010);
or U3288 (N_3288,N_3013,N_3174);
xor U3289 (N_3289,N_3132,N_2981);
or U3290 (N_3290,N_3162,N_2875);
or U3291 (N_3291,N_2862,N_2888);
nand U3292 (N_3292,N_2884,N_2839);
and U3293 (N_3293,N_3033,N_3070);
xnor U3294 (N_3294,N_3023,N_3182);
or U3295 (N_3295,N_3192,N_3058);
or U3296 (N_3296,N_3154,N_3166);
xor U3297 (N_3297,N_2877,N_3112);
or U3298 (N_3298,N_2850,N_3090);
or U3299 (N_3299,N_2891,N_3142);
nand U3300 (N_3300,N_2927,N_3078);
xor U3301 (N_3301,N_2833,N_2886);
and U3302 (N_3302,N_2801,N_3139);
and U3303 (N_3303,N_2963,N_2980);
nor U3304 (N_3304,N_2807,N_2993);
or U3305 (N_3305,N_2921,N_3095);
nor U3306 (N_3306,N_3135,N_2951);
nor U3307 (N_3307,N_2954,N_3176);
and U3308 (N_3308,N_2919,N_3040);
or U3309 (N_3309,N_2843,N_2885);
nor U3310 (N_3310,N_3037,N_2815);
and U3311 (N_3311,N_2970,N_3199);
or U3312 (N_3312,N_2871,N_2924);
or U3313 (N_3313,N_3067,N_3129);
xor U3314 (N_3314,N_2949,N_2856);
xnor U3315 (N_3315,N_3153,N_3180);
nor U3316 (N_3316,N_3193,N_2898);
and U3317 (N_3317,N_2957,N_3127);
and U3318 (N_3318,N_2906,N_2841);
and U3319 (N_3319,N_2813,N_2935);
nor U3320 (N_3320,N_3124,N_3035);
xor U3321 (N_3321,N_2965,N_2909);
nor U3322 (N_3322,N_2812,N_2823);
xnor U3323 (N_3323,N_2944,N_3062);
and U3324 (N_3324,N_2956,N_2916);
nor U3325 (N_3325,N_3123,N_3004);
nor U3326 (N_3326,N_3050,N_3164);
xor U3327 (N_3327,N_3187,N_3029);
or U3328 (N_3328,N_2997,N_2805);
or U3329 (N_3329,N_2922,N_2932);
nor U3330 (N_3330,N_3091,N_2983);
nand U3331 (N_3331,N_2878,N_2912);
xor U3332 (N_3332,N_3102,N_3158);
nor U3333 (N_3333,N_3191,N_3175);
xor U3334 (N_3334,N_2971,N_2936);
xor U3335 (N_3335,N_3188,N_2867);
or U3336 (N_3336,N_2868,N_2827);
nand U3337 (N_3337,N_2974,N_3161);
xor U3338 (N_3338,N_3189,N_3110);
and U3339 (N_3339,N_2910,N_2889);
xor U3340 (N_3340,N_3019,N_3107);
nand U3341 (N_3341,N_2905,N_2811);
and U3342 (N_3342,N_3009,N_3057);
nor U3343 (N_3343,N_3086,N_2874);
or U3344 (N_3344,N_3130,N_2933);
and U3345 (N_3345,N_2947,N_3106);
or U3346 (N_3346,N_3194,N_2907);
xnor U3347 (N_3347,N_3052,N_2966);
nand U3348 (N_3348,N_3186,N_2995);
and U3349 (N_3349,N_3020,N_3053);
nor U3350 (N_3350,N_3022,N_3122);
nand U3351 (N_3351,N_3026,N_3155);
xor U3352 (N_3352,N_3083,N_2855);
nor U3353 (N_3353,N_3150,N_2969);
xnor U3354 (N_3354,N_2930,N_2923);
or U3355 (N_3355,N_2998,N_3094);
nor U3356 (N_3356,N_3167,N_2914);
nand U3357 (N_3357,N_2946,N_2844);
and U3358 (N_3358,N_2900,N_2979);
nand U3359 (N_3359,N_3178,N_2915);
or U3360 (N_3360,N_2858,N_3138);
nor U3361 (N_3361,N_2837,N_3061);
and U3362 (N_3362,N_3014,N_2840);
nand U3363 (N_3363,N_3145,N_3076);
and U3364 (N_3364,N_3169,N_3080);
nand U3365 (N_3365,N_2941,N_2990);
nor U3366 (N_3366,N_2808,N_3027);
and U3367 (N_3367,N_3093,N_2940);
nand U3368 (N_3368,N_3047,N_2929);
nor U3369 (N_3369,N_3143,N_2988);
nor U3370 (N_3370,N_3099,N_2865);
or U3371 (N_3371,N_3024,N_2958);
and U3372 (N_3372,N_3137,N_3181);
nor U3373 (N_3373,N_2991,N_2870);
or U3374 (N_3374,N_3012,N_3120);
or U3375 (N_3375,N_2920,N_3148);
or U3376 (N_3376,N_2800,N_2831);
and U3377 (N_3377,N_3151,N_3041);
nand U3378 (N_3378,N_3079,N_3195);
nand U3379 (N_3379,N_3000,N_3160);
or U3380 (N_3380,N_2986,N_2802);
nor U3381 (N_3381,N_3184,N_3044);
or U3382 (N_3382,N_2968,N_2873);
xor U3383 (N_3383,N_2816,N_3054);
or U3384 (N_3384,N_2846,N_3092);
nor U3385 (N_3385,N_2834,N_3149);
nand U3386 (N_3386,N_3121,N_3144);
or U3387 (N_3387,N_2804,N_3156);
and U3388 (N_3388,N_3038,N_2897);
xnor U3389 (N_3389,N_2863,N_3125);
or U3390 (N_3390,N_2996,N_2852);
nand U3391 (N_3391,N_2822,N_2934);
xnor U3392 (N_3392,N_3183,N_3025);
nand U3393 (N_3393,N_3104,N_3081);
nand U3394 (N_3394,N_2964,N_2828);
or U3395 (N_3395,N_2810,N_3074);
nor U3396 (N_3396,N_2887,N_2925);
or U3397 (N_3397,N_3196,N_3072);
or U3398 (N_3398,N_3159,N_2835);
xnor U3399 (N_3399,N_3087,N_2955);
and U3400 (N_3400,N_3199,N_2973);
nor U3401 (N_3401,N_3184,N_2931);
and U3402 (N_3402,N_2999,N_3145);
xor U3403 (N_3403,N_2919,N_3197);
or U3404 (N_3404,N_2979,N_3032);
or U3405 (N_3405,N_2969,N_3009);
xor U3406 (N_3406,N_2944,N_3136);
xnor U3407 (N_3407,N_2920,N_3030);
nand U3408 (N_3408,N_2822,N_3092);
nand U3409 (N_3409,N_2926,N_2976);
or U3410 (N_3410,N_3006,N_2885);
nor U3411 (N_3411,N_2929,N_3073);
nor U3412 (N_3412,N_3194,N_3098);
xor U3413 (N_3413,N_2854,N_3042);
nand U3414 (N_3414,N_2814,N_3072);
nand U3415 (N_3415,N_3006,N_2978);
and U3416 (N_3416,N_2941,N_2962);
nor U3417 (N_3417,N_2928,N_3099);
or U3418 (N_3418,N_3063,N_2931);
nor U3419 (N_3419,N_3046,N_2989);
and U3420 (N_3420,N_2906,N_3087);
nand U3421 (N_3421,N_3104,N_2844);
and U3422 (N_3422,N_3159,N_3012);
nor U3423 (N_3423,N_2856,N_3026);
xnor U3424 (N_3424,N_3130,N_3081);
nor U3425 (N_3425,N_3154,N_3056);
nor U3426 (N_3426,N_2907,N_2876);
and U3427 (N_3427,N_2914,N_2916);
xnor U3428 (N_3428,N_2830,N_2929);
nor U3429 (N_3429,N_2979,N_3169);
nor U3430 (N_3430,N_2832,N_2990);
or U3431 (N_3431,N_3147,N_2835);
or U3432 (N_3432,N_3037,N_3058);
nor U3433 (N_3433,N_3099,N_2836);
and U3434 (N_3434,N_3136,N_2947);
nor U3435 (N_3435,N_3097,N_3068);
nor U3436 (N_3436,N_2878,N_2866);
nor U3437 (N_3437,N_3121,N_2881);
nor U3438 (N_3438,N_3192,N_3186);
nor U3439 (N_3439,N_2879,N_2819);
nor U3440 (N_3440,N_3193,N_2896);
and U3441 (N_3441,N_2838,N_3174);
nor U3442 (N_3442,N_3013,N_3066);
nand U3443 (N_3443,N_3051,N_3107);
or U3444 (N_3444,N_2817,N_2945);
or U3445 (N_3445,N_3118,N_3070);
nand U3446 (N_3446,N_2935,N_2811);
xnor U3447 (N_3447,N_3168,N_3006);
and U3448 (N_3448,N_2849,N_2825);
nand U3449 (N_3449,N_2807,N_3090);
nand U3450 (N_3450,N_2984,N_2940);
nand U3451 (N_3451,N_2919,N_3122);
nand U3452 (N_3452,N_3016,N_2886);
xor U3453 (N_3453,N_3088,N_2932);
nand U3454 (N_3454,N_2962,N_3099);
xnor U3455 (N_3455,N_2944,N_3000);
nor U3456 (N_3456,N_2978,N_2975);
nor U3457 (N_3457,N_3066,N_3122);
and U3458 (N_3458,N_2895,N_2845);
xor U3459 (N_3459,N_2881,N_3023);
or U3460 (N_3460,N_3126,N_2928);
nand U3461 (N_3461,N_2856,N_2889);
and U3462 (N_3462,N_3133,N_3117);
xnor U3463 (N_3463,N_3164,N_2904);
nand U3464 (N_3464,N_2839,N_3100);
xor U3465 (N_3465,N_3175,N_2897);
nor U3466 (N_3466,N_2872,N_2813);
nor U3467 (N_3467,N_3166,N_3081);
nand U3468 (N_3468,N_2986,N_3174);
and U3469 (N_3469,N_2933,N_2804);
xnor U3470 (N_3470,N_2934,N_2946);
and U3471 (N_3471,N_3189,N_2870);
or U3472 (N_3472,N_3038,N_2963);
nor U3473 (N_3473,N_2848,N_2881);
or U3474 (N_3474,N_2957,N_2979);
and U3475 (N_3475,N_2998,N_3139);
and U3476 (N_3476,N_3047,N_3172);
or U3477 (N_3477,N_2818,N_3142);
or U3478 (N_3478,N_2878,N_3084);
and U3479 (N_3479,N_2856,N_3002);
nor U3480 (N_3480,N_2981,N_2827);
xnor U3481 (N_3481,N_3068,N_2935);
or U3482 (N_3482,N_2822,N_3177);
and U3483 (N_3483,N_3159,N_2863);
nand U3484 (N_3484,N_3113,N_3100);
or U3485 (N_3485,N_2977,N_2992);
or U3486 (N_3486,N_2836,N_3034);
nor U3487 (N_3487,N_3076,N_2992);
xnor U3488 (N_3488,N_3045,N_3113);
xnor U3489 (N_3489,N_3161,N_3192);
or U3490 (N_3490,N_3160,N_2956);
and U3491 (N_3491,N_2836,N_3105);
and U3492 (N_3492,N_2919,N_2924);
xor U3493 (N_3493,N_2989,N_3017);
xor U3494 (N_3494,N_2975,N_3085);
or U3495 (N_3495,N_2849,N_3149);
xnor U3496 (N_3496,N_2839,N_2992);
or U3497 (N_3497,N_2916,N_3129);
xnor U3498 (N_3498,N_2823,N_2875);
nand U3499 (N_3499,N_2967,N_3075);
and U3500 (N_3500,N_2947,N_2873);
xnor U3501 (N_3501,N_2992,N_2893);
nor U3502 (N_3502,N_3171,N_2918);
nor U3503 (N_3503,N_2885,N_2904);
and U3504 (N_3504,N_3032,N_2815);
or U3505 (N_3505,N_2993,N_2848);
nor U3506 (N_3506,N_2815,N_2972);
nor U3507 (N_3507,N_2906,N_3126);
or U3508 (N_3508,N_2947,N_2997);
nand U3509 (N_3509,N_3164,N_3099);
or U3510 (N_3510,N_2861,N_3081);
nand U3511 (N_3511,N_2856,N_3099);
and U3512 (N_3512,N_3097,N_2962);
nor U3513 (N_3513,N_3180,N_2965);
nor U3514 (N_3514,N_2808,N_2927);
nand U3515 (N_3515,N_2934,N_2955);
xor U3516 (N_3516,N_2928,N_2914);
nand U3517 (N_3517,N_3179,N_2889);
or U3518 (N_3518,N_2904,N_2827);
nand U3519 (N_3519,N_2955,N_2959);
and U3520 (N_3520,N_3029,N_2877);
nand U3521 (N_3521,N_2941,N_3114);
nand U3522 (N_3522,N_3187,N_3004);
nand U3523 (N_3523,N_3028,N_3163);
or U3524 (N_3524,N_3133,N_3100);
and U3525 (N_3525,N_2921,N_2810);
and U3526 (N_3526,N_3084,N_3053);
or U3527 (N_3527,N_2964,N_3178);
nor U3528 (N_3528,N_3035,N_3027);
xor U3529 (N_3529,N_3171,N_2963);
or U3530 (N_3530,N_2939,N_3174);
and U3531 (N_3531,N_3190,N_3076);
nand U3532 (N_3532,N_3152,N_3156);
nand U3533 (N_3533,N_3049,N_2988);
or U3534 (N_3534,N_3036,N_2843);
nor U3535 (N_3535,N_3089,N_3052);
or U3536 (N_3536,N_3145,N_3059);
nor U3537 (N_3537,N_2803,N_3067);
and U3538 (N_3538,N_2954,N_3079);
and U3539 (N_3539,N_2809,N_2842);
or U3540 (N_3540,N_3116,N_2942);
nor U3541 (N_3541,N_3040,N_2908);
or U3542 (N_3542,N_2941,N_3140);
xnor U3543 (N_3543,N_2986,N_3193);
nand U3544 (N_3544,N_2954,N_2825);
or U3545 (N_3545,N_2800,N_2865);
nand U3546 (N_3546,N_2872,N_2852);
or U3547 (N_3547,N_3021,N_2861);
and U3548 (N_3548,N_2986,N_2942);
nor U3549 (N_3549,N_3094,N_3054);
or U3550 (N_3550,N_3104,N_3089);
and U3551 (N_3551,N_3043,N_2817);
and U3552 (N_3552,N_3098,N_3123);
nor U3553 (N_3553,N_3034,N_2987);
or U3554 (N_3554,N_2938,N_3142);
xor U3555 (N_3555,N_2942,N_2919);
or U3556 (N_3556,N_2839,N_2849);
nor U3557 (N_3557,N_3194,N_3020);
or U3558 (N_3558,N_3082,N_3023);
nor U3559 (N_3559,N_3194,N_2852);
xnor U3560 (N_3560,N_2804,N_3132);
or U3561 (N_3561,N_3154,N_2952);
or U3562 (N_3562,N_3078,N_2816);
nand U3563 (N_3563,N_3129,N_2969);
nand U3564 (N_3564,N_3097,N_2872);
and U3565 (N_3565,N_3161,N_3109);
and U3566 (N_3566,N_3087,N_3085);
nand U3567 (N_3567,N_2926,N_3150);
xnor U3568 (N_3568,N_2946,N_2909);
or U3569 (N_3569,N_2906,N_2853);
and U3570 (N_3570,N_2881,N_2897);
nor U3571 (N_3571,N_2847,N_3190);
and U3572 (N_3572,N_3195,N_3130);
nand U3573 (N_3573,N_3083,N_2937);
nand U3574 (N_3574,N_2828,N_3077);
nand U3575 (N_3575,N_2855,N_3102);
nor U3576 (N_3576,N_3176,N_2922);
xnor U3577 (N_3577,N_3105,N_3145);
or U3578 (N_3578,N_2810,N_2802);
and U3579 (N_3579,N_2995,N_2972);
xor U3580 (N_3580,N_3089,N_2986);
xnor U3581 (N_3581,N_3116,N_3063);
nor U3582 (N_3582,N_2804,N_3044);
xnor U3583 (N_3583,N_3019,N_3029);
or U3584 (N_3584,N_3171,N_2947);
or U3585 (N_3585,N_2987,N_2968);
and U3586 (N_3586,N_2899,N_2884);
nand U3587 (N_3587,N_2919,N_3052);
nand U3588 (N_3588,N_3040,N_2978);
xor U3589 (N_3589,N_3149,N_3155);
nor U3590 (N_3590,N_2830,N_3046);
and U3591 (N_3591,N_2993,N_2868);
nor U3592 (N_3592,N_3049,N_2892);
nor U3593 (N_3593,N_3031,N_2822);
and U3594 (N_3594,N_2804,N_3141);
nand U3595 (N_3595,N_3188,N_3166);
nor U3596 (N_3596,N_3022,N_3060);
or U3597 (N_3597,N_2995,N_3072);
nand U3598 (N_3598,N_3133,N_2885);
nand U3599 (N_3599,N_3033,N_2887);
xor U3600 (N_3600,N_3594,N_3246);
and U3601 (N_3601,N_3519,N_3560);
nand U3602 (N_3602,N_3523,N_3331);
nand U3603 (N_3603,N_3505,N_3529);
nor U3604 (N_3604,N_3209,N_3296);
and U3605 (N_3605,N_3319,N_3305);
nor U3606 (N_3606,N_3596,N_3348);
nor U3607 (N_3607,N_3547,N_3432);
nand U3608 (N_3608,N_3537,N_3384);
or U3609 (N_3609,N_3201,N_3288);
nand U3610 (N_3610,N_3369,N_3234);
xnor U3611 (N_3611,N_3309,N_3585);
xnor U3612 (N_3612,N_3409,N_3395);
nand U3613 (N_3613,N_3407,N_3251);
xor U3614 (N_3614,N_3219,N_3487);
and U3615 (N_3615,N_3490,N_3206);
xnor U3616 (N_3616,N_3279,N_3474);
or U3617 (N_3617,N_3464,N_3308);
nand U3618 (N_3618,N_3479,N_3303);
and U3619 (N_3619,N_3412,N_3447);
and U3620 (N_3620,N_3315,N_3227);
xor U3621 (N_3621,N_3549,N_3451);
and U3622 (N_3622,N_3586,N_3530);
xnor U3623 (N_3623,N_3563,N_3415);
nor U3624 (N_3624,N_3213,N_3354);
nor U3625 (N_3625,N_3438,N_3420);
nor U3626 (N_3626,N_3581,N_3345);
xnor U3627 (N_3627,N_3245,N_3314);
xnor U3628 (N_3628,N_3427,N_3244);
nand U3629 (N_3629,N_3297,N_3332);
xnor U3630 (N_3630,N_3437,N_3365);
nor U3631 (N_3631,N_3590,N_3439);
and U3632 (N_3632,N_3231,N_3295);
or U3633 (N_3633,N_3250,N_3272);
nor U3634 (N_3634,N_3265,N_3401);
nand U3635 (N_3635,N_3214,N_3429);
and U3636 (N_3636,N_3321,N_3249);
and U3637 (N_3637,N_3564,N_3471);
nand U3638 (N_3638,N_3504,N_3416);
nand U3639 (N_3639,N_3388,N_3204);
and U3640 (N_3640,N_3285,N_3258);
nor U3641 (N_3641,N_3255,N_3459);
and U3642 (N_3642,N_3476,N_3382);
nand U3643 (N_3643,N_3521,N_3466);
nor U3644 (N_3644,N_3394,N_3240);
nor U3645 (N_3645,N_3210,N_3555);
and U3646 (N_3646,N_3557,N_3327);
and U3647 (N_3647,N_3374,N_3402);
xnor U3648 (N_3648,N_3253,N_3575);
and U3649 (N_3649,N_3270,N_3486);
nor U3650 (N_3650,N_3310,N_3511);
or U3651 (N_3651,N_3299,N_3572);
xor U3652 (N_3652,N_3228,N_3524);
xnor U3653 (N_3653,N_3243,N_3443);
or U3654 (N_3654,N_3462,N_3280);
and U3655 (N_3655,N_3503,N_3478);
and U3656 (N_3656,N_3358,N_3460);
and U3657 (N_3657,N_3455,N_3533);
xor U3658 (N_3658,N_3597,N_3329);
or U3659 (N_3659,N_3256,N_3263);
and U3660 (N_3660,N_3553,N_3411);
nor U3661 (N_3661,N_3540,N_3337);
xor U3662 (N_3662,N_3525,N_3262);
and U3663 (N_3663,N_3452,N_3548);
nand U3664 (N_3664,N_3498,N_3220);
nand U3665 (N_3665,N_3458,N_3284);
or U3666 (N_3666,N_3495,N_3569);
and U3667 (N_3667,N_3221,N_3283);
and U3668 (N_3668,N_3208,N_3287);
and U3669 (N_3669,N_3326,N_3468);
and U3670 (N_3670,N_3440,N_3494);
and U3671 (N_3671,N_3334,N_3323);
or U3672 (N_3672,N_3376,N_3304);
nand U3673 (N_3673,N_3517,N_3482);
and U3674 (N_3674,N_3344,N_3398);
nand U3675 (N_3675,N_3470,N_3215);
xnor U3676 (N_3676,N_3424,N_3218);
nand U3677 (N_3677,N_3264,N_3377);
xnor U3678 (N_3678,N_3268,N_3343);
xnor U3679 (N_3679,N_3306,N_3472);
and U3680 (N_3680,N_3535,N_3276);
or U3681 (N_3681,N_3469,N_3252);
xnor U3682 (N_3682,N_3266,N_3274);
nand U3683 (N_3683,N_3532,N_3372);
or U3684 (N_3684,N_3527,N_3520);
and U3685 (N_3685,N_3502,N_3399);
nor U3686 (N_3686,N_3313,N_3580);
and U3687 (N_3687,N_3408,N_3387);
or U3688 (N_3688,N_3294,N_3561);
or U3689 (N_3689,N_3342,N_3328);
and U3690 (N_3690,N_3538,N_3271);
or U3691 (N_3691,N_3480,N_3542);
or U3692 (N_3692,N_3577,N_3446);
and U3693 (N_3693,N_3457,N_3592);
and U3694 (N_3694,N_3587,N_3428);
or U3695 (N_3695,N_3426,N_3477);
and U3696 (N_3696,N_3422,N_3225);
nand U3697 (N_3697,N_3565,N_3257);
nor U3698 (N_3698,N_3442,N_3423);
nor U3699 (N_3699,N_3551,N_3397);
or U3700 (N_3700,N_3340,N_3510);
or U3701 (N_3701,N_3320,N_3403);
xor U3702 (N_3702,N_3237,N_3368);
and U3703 (N_3703,N_3559,N_3355);
nand U3704 (N_3704,N_3599,N_3230);
nor U3705 (N_3705,N_3278,N_3324);
and U3706 (N_3706,N_3545,N_3336);
and U3707 (N_3707,N_3335,N_3341);
and U3708 (N_3708,N_3373,N_3291);
or U3709 (N_3709,N_3558,N_3528);
and U3710 (N_3710,N_3473,N_3531);
nand U3711 (N_3711,N_3302,N_3353);
and U3712 (N_3712,N_3364,N_3570);
and U3713 (N_3713,N_3410,N_3346);
or U3714 (N_3714,N_3212,N_3259);
and U3715 (N_3715,N_3307,N_3582);
and U3716 (N_3716,N_3400,N_3325);
xor U3717 (N_3717,N_3450,N_3444);
nor U3718 (N_3718,N_3514,N_3200);
nand U3719 (N_3719,N_3235,N_3456);
xor U3720 (N_3720,N_3496,N_3431);
and U3721 (N_3721,N_3216,N_3367);
xnor U3722 (N_3722,N_3534,N_3539);
xnor U3723 (N_3723,N_3406,N_3571);
nand U3724 (N_3724,N_3544,N_3293);
and U3725 (N_3725,N_3485,N_3390);
nand U3726 (N_3726,N_3391,N_3556);
xnor U3727 (N_3727,N_3238,N_3361);
xor U3728 (N_3728,N_3589,N_3389);
nand U3729 (N_3729,N_3573,N_3425);
xor U3730 (N_3730,N_3393,N_3404);
and U3731 (N_3731,N_3375,N_3378);
xnor U3732 (N_3732,N_3546,N_3317);
and U3733 (N_3733,N_3300,N_3366);
nor U3734 (N_3734,N_3435,N_3461);
nand U3735 (N_3735,N_3499,N_3386);
nand U3736 (N_3736,N_3260,N_3261);
xnor U3737 (N_3737,N_3493,N_3282);
and U3738 (N_3738,N_3509,N_3554);
nand U3739 (N_3739,N_3475,N_3232);
xnor U3740 (N_3740,N_3226,N_3311);
nor U3741 (N_3741,N_3491,N_3506);
or U3742 (N_3742,N_3449,N_3363);
or U3743 (N_3743,N_3593,N_3352);
or U3744 (N_3744,N_3383,N_3417);
or U3745 (N_3745,N_3360,N_3500);
and U3746 (N_3746,N_3465,N_3489);
or U3747 (N_3747,N_3350,N_3513);
and U3748 (N_3748,N_3568,N_3298);
xnor U3749 (N_3749,N_3598,N_3351);
xor U3750 (N_3750,N_3567,N_3357);
nand U3751 (N_3751,N_3413,N_3522);
and U3752 (N_3752,N_3508,N_3543);
and U3753 (N_3753,N_3380,N_3405);
nand U3754 (N_3754,N_3217,N_3359);
nand U3755 (N_3755,N_3205,N_3541);
nand U3756 (N_3756,N_3290,N_3267);
nand U3757 (N_3757,N_3281,N_3515);
or U3758 (N_3758,N_3552,N_3497);
nand U3759 (N_3759,N_3301,N_3211);
and U3760 (N_3760,N_3289,N_3233);
or U3761 (N_3761,N_3436,N_3379);
and U3762 (N_3762,N_3418,N_3441);
xor U3763 (N_3763,N_3536,N_3322);
nor U3764 (N_3764,N_3339,N_3488);
nor U3765 (N_3765,N_3516,N_3241);
xnor U3766 (N_3766,N_3316,N_3562);
and U3767 (N_3767,N_3445,N_3578);
and U3768 (N_3768,N_3349,N_3242);
xor U3769 (N_3769,N_3338,N_3588);
xnor U3770 (N_3770,N_3518,N_3275);
or U3771 (N_3771,N_3421,N_3254);
or U3772 (N_3772,N_3392,N_3236);
or U3773 (N_3773,N_3484,N_3453);
xor U3774 (N_3774,N_3370,N_3448);
xor U3775 (N_3775,N_3584,N_3318);
and U3776 (N_3776,N_3574,N_3330);
xor U3777 (N_3777,N_3396,N_3371);
or U3778 (N_3778,N_3381,N_3433);
xor U3779 (N_3779,N_3434,N_3222);
and U3780 (N_3780,N_3454,N_3347);
and U3781 (N_3781,N_3286,N_3483);
or U3782 (N_3782,N_3385,N_3223);
or U3783 (N_3783,N_3550,N_3481);
and U3784 (N_3784,N_3583,N_3566);
and U3785 (N_3785,N_3207,N_3202);
xor U3786 (N_3786,N_3224,N_3595);
or U3787 (N_3787,N_3247,N_3273);
and U3788 (N_3788,N_3492,N_3526);
and U3789 (N_3789,N_3248,N_3507);
nand U3790 (N_3790,N_3467,N_3269);
nand U3791 (N_3791,N_3312,N_3292);
or U3792 (N_3792,N_3229,N_3576);
nand U3793 (N_3793,N_3362,N_3356);
and U3794 (N_3794,N_3203,N_3591);
nand U3795 (N_3795,N_3430,N_3333);
and U3796 (N_3796,N_3414,N_3463);
nand U3797 (N_3797,N_3579,N_3501);
nor U3798 (N_3798,N_3419,N_3239);
nor U3799 (N_3799,N_3512,N_3277);
nor U3800 (N_3800,N_3593,N_3503);
and U3801 (N_3801,N_3473,N_3454);
or U3802 (N_3802,N_3335,N_3312);
nor U3803 (N_3803,N_3268,N_3496);
nand U3804 (N_3804,N_3303,N_3313);
xnor U3805 (N_3805,N_3599,N_3248);
and U3806 (N_3806,N_3328,N_3397);
and U3807 (N_3807,N_3545,N_3458);
nor U3808 (N_3808,N_3353,N_3357);
or U3809 (N_3809,N_3529,N_3565);
or U3810 (N_3810,N_3451,N_3320);
or U3811 (N_3811,N_3509,N_3401);
xnor U3812 (N_3812,N_3314,N_3531);
nand U3813 (N_3813,N_3294,N_3524);
or U3814 (N_3814,N_3483,N_3423);
xor U3815 (N_3815,N_3279,N_3276);
or U3816 (N_3816,N_3555,N_3228);
nand U3817 (N_3817,N_3595,N_3300);
nand U3818 (N_3818,N_3277,N_3359);
xnor U3819 (N_3819,N_3331,N_3323);
nor U3820 (N_3820,N_3235,N_3527);
nand U3821 (N_3821,N_3565,N_3231);
nor U3822 (N_3822,N_3429,N_3550);
nor U3823 (N_3823,N_3444,N_3355);
nand U3824 (N_3824,N_3347,N_3462);
nand U3825 (N_3825,N_3402,N_3593);
or U3826 (N_3826,N_3315,N_3421);
nor U3827 (N_3827,N_3221,N_3428);
nor U3828 (N_3828,N_3373,N_3344);
xnor U3829 (N_3829,N_3510,N_3203);
xnor U3830 (N_3830,N_3237,N_3378);
nor U3831 (N_3831,N_3224,N_3322);
or U3832 (N_3832,N_3387,N_3420);
nor U3833 (N_3833,N_3447,N_3430);
xnor U3834 (N_3834,N_3322,N_3462);
and U3835 (N_3835,N_3388,N_3505);
xor U3836 (N_3836,N_3536,N_3553);
nand U3837 (N_3837,N_3523,N_3416);
xnor U3838 (N_3838,N_3325,N_3225);
xor U3839 (N_3839,N_3332,N_3262);
and U3840 (N_3840,N_3277,N_3351);
xor U3841 (N_3841,N_3384,N_3507);
and U3842 (N_3842,N_3412,N_3210);
or U3843 (N_3843,N_3512,N_3536);
xnor U3844 (N_3844,N_3461,N_3427);
xor U3845 (N_3845,N_3489,N_3434);
xnor U3846 (N_3846,N_3342,N_3324);
and U3847 (N_3847,N_3270,N_3364);
xnor U3848 (N_3848,N_3491,N_3593);
nand U3849 (N_3849,N_3443,N_3545);
nor U3850 (N_3850,N_3214,N_3441);
xor U3851 (N_3851,N_3312,N_3593);
nand U3852 (N_3852,N_3457,N_3489);
nand U3853 (N_3853,N_3542,N_3487);
nor U3854 (N_3854,N_3222,N_3392);
or U3855 (N_3855,N_3562,N_3354);
nand U3856 (N_3856,N_3415,N_3279);
or U3857 (N_3857,N_3486,N_3275);
and U3858 (N_3858,N_3446,N_3588);
or U3859 (N_3859,N_3451,N_3233);
nor U3860 (N_3860,N_3553,N_3523);
and U3861 (N_3861,N_3287,N_3568);
or U3862 (N_3862,N_3439,N_3487);
nand U3863 (N_3863,N_3321,N_3224);
nor U3864 (N_3864,N_3535,N_3591);
and U3865 (N_3865,N_3429,N_3565);
xor U3866 (N_3866,N_3597,N_3559);
and U3867 (N_3867,N_3563,N_3473);
nand U3868 (N_3868,N_3553,N_3422);
and U3869 (N_3869,N_3231,N_3554);
xor U3870 (N_3870,N_3315,N_3290);
or U3871 (N_3871,N_3395,N_3396);
nand U3872 (N_3872,N_3348,N_3273);
nor U3873 (N_3873,N_3251,N_3313);
xnor U3874 (N_3874,N_3271,N_3212);
or U3875 (N_3875,N_3575,N_3440);
nor U3876 (N_3876,N_3235,N_3578);
or U3877 (N_3877,N_3506,N_3369);
nand U3878 (N_3878,N_3220,N_3384);
nor U3879 (N_3879,N_3226,N_3481);
or U3880 (N_3880,N_3224,N_3298);
nor U3881 (N_3881,N_3476,N_3540);
or U3882 (N_3882,N_3537,N_3315);
or U3883 (N_3883,N_3514,N_3588);
or U3884 (N_3884,N_3416,N_3495);
nor U3885 (N_3885,N_3520,N_3311);
or U3886 (N_3886,N_3513,N_3389);
nand U3887 (N_3887,N_3247,N_3475);
xor U3888 (N_3888,N_3424,N_3309);
and U3889 (N_3889,N_3291,N_3289);
nand U3890 (N_3890,N_3303,N_3385);
xnor U3891 (N_3891,N_3286,N_3423);
or U3892 (N_3892,N_3225,N_3568);
nor U3893 (N_3893,N_3409,N_3279);
nand U3894 (N_3894,N_3252,N_3239);
nand U3895 (N_3895,N_3228,N_3331);
and U3896 (N_3896,N_3543,N_3364);
xor U3897 (N_3897,N_3212,N_3268);
and U3898 (N_3898,N_3228,N_3423);
nand U3899 (N_3899,N_3560,N_3237);
nand U3900 (N_3900,N_3323,N_3237);
nand U3901 (N_3901,N_3333,N_3473);
or U3902 (N_3902,N_3373,N_3343);
xor U3903 (N_3903,N_3383,N_3236);
nor U3904 (N_3904,N_3269,N_3585);
and U3905 (N_3905,N_3451,N_3278);
or U3906 (N_3906,N_3576,N_3426);
nor U3907 (N_3907,N_3523,N_3296);
nand U3908 (N_3908,N_3335,N_3207);
nor U3909 (N_3909,N_3467,N_3412);
nor U3910 (N_3910,N_3213,N_3503);
nand U3911 (N_3911,N_3522,N_3431);
nor U3912 (N_3912,N_3418,N_3273);
nand U3913 (N_3913,N_3294,N_3445);
and U3914 (N_3914,N_3400,N_3426);
xnor U3915 (N_3915,N_3478,N_3425);
and U3916 (N_3916,N_3422,N_3589);
and U3917 (N_3917,N_3445,N_3385);
or U3918 (N_3918,N_3599,N_3535);
nand U3919 (N_3919,N_3415,N_3449);
nand U3920 (N_3920,N_3301,N_3572);
nand U3921 (N_3921,N_3331,N_3271);
nor U3922 (N_3922,N_3520,N_3561);
xnor U3923 (N_3923,N_3397,N_3599);
nor U3924 (N_3924,N_3251,N_3278);
nand U3925 (N_3925,N_3571,N_3366);
and U3926 (N_3926,N_3249,N_3580);
or U3927 (N_3927,N_3325,N_3561);
nand U3928 (N_3928,N_3218,N_3406);
nand U3929 (N_3929,N_3438,N_3519);
xnor U3930 (N_3930,N_3422,N_3330);
nand U3931 (N_3931,N_3509,N_3237);
nand U3932 (N_3932,N_3366,N_3223);
nor U3933 (N_3933,N_3388,N_3200);
or U3934 (N_3934,N_3479,N_3205);
and U3935 (N_3935,N_3212,N_3217);
xor U3936 (N_3936,N_3524,N_3499);
nor U3937 (N_3937,N_3346,N_3275);
and U3938 (N_3938,N_3290,N_3489);
nor U3939 (N_3939,N_3408,N_3205);
nor U3940 (N_3940,N_3377,N_3459);
and U3941 (N_3941,N_3447,N_3468);
and U3942 (N_3942,N_3440,N_3587);
nand U3943 (N_3943,N_3543,N_3336);
nor U3944 (N_3944,N_3511,N_3246);
and U3945 (N_3945,N_3378,N_3497);
or U3946 (N_3946,N_3389,N_3286);
nand U3947 (N_3947,N_3447,N_3359);
nand U3948 (N_3948,N_3537,N_3253);
xnor U3949 (N_3949,N_3596,N_3315);
and U3950 (N_3950,N_3527,N_3484);
and U3951 (N_3951,N_3309,N_3293);
or U3952 (N_3952,N_3267,N_3416);
xor U3953 (N_3953,N_3469,N_3341);
and U3954 (N_3954,N_3493,N_3326);
or U3955 (N_3955,N_3272,N_3241);
and U3956 (N_3956,N_3209,N_3510);
nand U3957 (N_3957,N_3449,N_3528);
nand U3958 (N_3958,N_3335,N_3259);
nor U3959 (N_3959,N_3479,N_3432);
xor U3960 (N_3960,N_3417,N_3223);
nor U3961 (N_3961,N_3367,N_3217);
or U3962 (N_3962,N_3263,N_3352);
and U3963 (N_3963,N_3550,N_3360);
nand U3964 (N_3964,N_3238,N_3264);
or U3965 (N_3965,N_3451,N_3413);
or U3966 (N_3966,N_3318,N_3570);
and U3967 (N_3967,N_3222,N_3557);
or U3968 (N_3968,N_3550,N_3332);
xnor U3969 (N_3969,N_3270,N_3594);
or U3970 (N_3970,N_3255,N_3305);
or U3971 (N_3971,N_3219,N_3580);
xor U3972 (N_3972,N_3493,N_3582);
nor U3973 (N_3973,N_3371,N_3208);
nand U3974 (N_3974,N_3462,N_3281);
and U3975 (N_3975,N_3564,N_3398);
nand U3976 (N_3976,N_3204,N_3476);
nand U3977 (N_3977,N_3268,N_3225);
or U3978 (N_3978,N_3505,N_3561);
or U3979 (N_3979,N_3593,N_3327);
or U3980 (N_3980,N_3223,N_3426);
or U3981 (N_3981,N_3496,N_3378);
nand U3982 (N_3982,N_3261,N_3267);
xor U3983 (N_3983,N_3446,N_3570);
or U3984 (N_3984,N_3254,N_3577);
or U3985 (N_3985,N_3332,N_3450);
nor U3986 (N_3986,N_3290,N_3467);
and U3987 (N_3987,N_3207,N_3237);
nand U3988 (N_3988,N_3393,N_3429);
and U3989 (N_3989,N_3431,N_3490);
nor U3990 (N_3990,N_3249,N_3528);
xnor U3991 (N_3991,N_3576,N_3334);
xor U3992 (N_3992,N_3218,N_3202);
or U3993 (N_3993,N_3595,N_3246);
nor U3994 (N_3994,N_3564,N_3309);
and U3995 (N_3995,N_3420,N_3576);
xor U3996 (N_3996,N_3561,N_3328);
xnor U3997 (N_3997,N_3529,N_3479);
nor U3998 (N_3998,N_3377,N_3534);
nor U3999 (N_3999,N_3592,N_3500);
and U4000 (N_4000,N_3859,N_3804);
nand U4001 (N_4001,N_3778,N_3767);
and U4002 (N_4002,N_3784,N_3770);
nor U4003 (N_4003,N_3895,N_3671);
or U4004 (N_4004,N_3818,N_3891);
nand U4005 (N_4005,N_3983,N_3606);
and U4006 (N_4006,N_3824,N_3880);
or U4007 (N_4007,N_3973,N_3688);
xnor U4008 (N_4008,N_3947,N_3650);
xnor U4009 (N_4009,N_3972,N_3939);
or U4010 (N_4010,N_3788,N_3633);
xnor U4011 (N_4011,N_3902,N_3833);
and U4012 (N_4012,N_3830,N_3709);
and U4013 (N_4013,N_3917,N_3635);
xor U4014 (N_4014,N_3748,N_3812);
or U4015 (N_4015,N_3881,N_3660);
nand U4016 (N_4016,N_3847,N_3640);
xnor U4017 (N_4017,N_3716,N_3913);
xnor U4018 (N_4018,N_3747,N_3900);
xnor U4019 (N_4019,N_3736,N_3651);
xnor U4020 (N_4020,N_3740,N_3791);
or U4021 (N_4021,N_3643,N_3874);
nor U4022 (N_4022,N_3673,N_3738);
or U4023 (N_4023,N_3906,N_3963);
or U4024 (N_4024,N_3867,N_3836);
xor U4025 (N_4025,N_3618,N_3607);
nor U4026 (N_4026,N_3807,N_3990);
nor U4027 (N_4027,N_3999,N_3863);
xnor U4028 (N_4028,N_3931,N_3619);
nor U4029 (N_4029,N_3893,N_3873);
xor U4030 (N_4030,N_3670,N_3711);
or U4031 (N_4031,N_3745,N_3879);
nor U4032 (N_4032,N_3678,N_3706);
and U4033 (N_4033,N_3734,N_3666);
or U4034 (N_4034,N_3679,N_3687);
and U4035 (N_4035,N_3732,N_3754);
xor U4036 (N_4036,N_3890,N_3831);
and U4037 (N_4037,N_3882,N_3652);
nor U4038 (N_4038,N_3970,N_3855);
nor U4039 (N_4039,N_3760,N_3667);
and U4040 (N_4040,N_3648,N_3968);
nand U4041 (N_4041,N_3612,N_3665);
or U4042 (N_4042,N_3783,N_3878);
nand U4043 (N_4043,N_3842,N_3759);
xnor U4044 (N_4044,N_3884,N_3914);
or U4045 (N_4045,N_3676,N_3712);
nand U4046 (N_4046,N_3845,N_3720);
nand U4047 (N_4047,N_3866,N_3800);
nand U4048 (N_4048,N_3647,N_3657);
and U4049 (N_4049,N_3953,N_3834);
and U4050 (N_4050,N_3645,N_3802);
nor U4051 (N_4051,N_3739,N_3725);
and U4052 (N_4052,N_3871,N_3792);
nor U4053 (N_4053,N_3630,N_3659);
and U4054 (N_4054,N_3785,N_3623);
and U4055 (N_4055,N_3624,N_3625);
nand U4056 (N_4056,N_3769,N_3705);
nor U4057 (N_4057,N_3786,N_3954);
or U4058 (N_4058,N_3961,N_3932);
xnor U4059 (N_4059,N_3975,N_3974);
and U4060 (N_4060,N_3951,N_3865);
nor U4061 (N_4061,N_3699,N_3813);
and U4062 (N_4062,N_3929,N_3952);
or U4063 (N_4063,N_3921,N_3779);
nand U4064 (N_4064,N_3762,N_3795);
nand U4065 (N_4065,N_3735,N_3780);
nor U4066 (N_4066,N_3924,N_3823);
nor U4067 (N_4067,N_3835,N_3996);
or U4068 (N_4068,N_3885,N_3985);
nor U4069 (N_4069,N_3601,N_3971);
nand U4070 (N_4070,N_3819,N_3799);
nand U4071 (N_4071,N_3946,N_3909);
and U4072 (N_4072,N_3758,N_3658);
or U4073 (N_4073,N_3628,N_3926);
and U4074 (N_4074,N_3677,N_3701);
nor U4075 (N_4075,N_3627,N_3771);
xor U4076 (N_4076,N_3850,N_3982);
xnor U4077 (N_4077,N_3825,N_3768);
nor U4078 (N_4078,N_3984,N_3719);
and U4079 (N_4079,N_3856,N_3753);
nand U4080 (N_4080,N_3776,N_3989);
and U4081 (N_4081,N_3896,N_3663);
nand U4082 (N_4082,N_3948,N_3827);
nand U4083 (N_4083,N_3629,N_3899);
and U4084 (N_4084,N_3700,N_3993);
nor U4085 (N_4085,N_3763,N_3694);
xor U4086 (N_4086,N_3641,N_3892);
nor U4087 (N_4087,N_3978,N_3730);
nor U4088 (N_4088,N_3649,N_3870);
or U4089 (N_4089,N_3904,N_3756);
xnor U4090 (N_4090,N_3793,N_3668);
and U4091 (N_4091,N_3944,N_3696);
xor U4092 (N_4092,N_3962,N_3684);
or U4093 (N_4093,N_3811,N_3689);
nor U4094 (N_4094,N_3790,N_3883);
or U4095 (N_4095,N_3622,N_3693);
or U4096 (N_4096,N_3614,N_3654);
or U4097 (N_4097,N_3782,N_3702);
xnor U4098 (N_4098,N_3981,N_3814);
or U4099 (N_4099,N_3936,N_3897);
or U4100 (N_4100,N_3639,N_3766);
nor U4101 (N_4101,N_3949,N_3774);
xnor U4102 (N_4102,N_3682,N_3940);
xnor U4103 (N_4103,N_3632,N_3886);
nor U4104 (N_4104,N_3937,N_3726);
nand U4105 (N_4105,N_3631,N_3761);
nand U4106 (N_4106,N_3826,N_3964);
xnor U4107 (N_4107,N_3731,N_3988);
xor U4108 (N_4108,N_3898,N_3894);
nor U4109 (N_4109,N_3801,N_3777);
nand U4110 (N_4110,N_3656,N_3805);
or U4111 (N_4111,N_3943,N_3644);
and U4112 (N_4112,N_3848,N_3822);
or U4113 (N_4113,N_3728,N_3752);
nor U4114 (N_4114,N_3724,N_3608);
nor U4115 (N_4115,N_3765,N_3723);
nand U4116 (N_4116,N_3683,N_3789);
nor U4117 (N_4117,N_3621,N_3613);
nand U4118 (N_4118,N_3957,N_3797);
or U4119 (N_4119,N_3945,N_3849);
or U4120 (N_4120,N_3923,N_3710);
xor U4121 (N_4121,N_3887,N_3987);
nor U4122 (N_4122,N_3979,N_3672);
nor U4123 (N_4123,N_3888,N_3815);
nand U4124 (N_4124,N_3857,N_3718);
nor U4125 (N_4125,N_3609,N_3994);
or U4126 (N_4126,N_3832,N_3603);
nor U4127 (N_4127,N_3992,N_3746);
nand U4128 (N_4128,N_3794,N_3916);
xnor U4129 (N_4129,N_3956,N_3772);
nor U4130 (N_4130,N_3602,N_3717);
nor U4131 (N_4131,N_3600,N_3860);
and U4132 (N_4132,N_3773,N_3715);
nand U4133 (N_4133,N_3828,N_3869);
xor U4134 (N_4134,N_3820,N_3912);
nor U4135 (N_4135,N_3862,N_3617);
or U4136 (N_4136,N_3919,N_3675);
nand U4137 (N_4137,N_3809,N_3707);
nor U4138 (N_4138,N_3955,N_3755);
xor U4139 (N_4139,N_3930,N_3729);
xnor U4140 (N_4140,N_3674,N_3685);
nand U4141 (N_4141,N_3959,N_3941);
nand U4142 (N_4142,N_3965,N_3751);
or U4143 (N_4143,N_3889,N_3634);
xnor U4144 (N_4144,N_3703,N_3698);
xnor U4145 (N_4145,N_3911,N_3669);
xor U4146 (N_4146,N_3872,N_3655);
nor U4147 (N_4147,N_3722,N_3977);
nor U4148 (N_4148,N_3966,N_3744);
and U4149 (N_4149,N_3796,N_3781);
or U4150 (N_4150,N_3713,N_3838);
and U4151 (N_4151,N_3920,N_3803);
and U4152 (N_4152,N_3611,N_3806);
xor U4153 (N_4153,N_3626,N_3829);
xnor U4154 (N_4154,N_3901,N_3976);
nand U4155 (N_4155,N_3757,N_3750);
and U4156 (N_4156,N_3697,N_3733);
and U4157 (N_4157,N_3817,N_3810);
and U4158 (N_4158,N_3997,N_3816);
nand U4159 (N_4159,N_3910,N_3664);
or U4160 (N_4160,N_3737,N_3708);
nand U4161 (N_4161,N_3868,N_3915);
and U4162 (N_4162,N_3935,N_3605);
and U4163 (N_4163,N_3653,N_3636);
and U4164 (N_4164,N_3616,N_3995);
or U4165 (N_4165,N_3690,N_3852);
or U4166 (N_4166,N_3714,N_3704);
and U4167 (N_4167,N_3692,N_3695);
nand U4168 (N_4168,N_3918,N_3908);
or U4169 (N_4169,N_3604,N_3749);
nand U4170 (N_4170,N_3637,N_3840);
nand U4171 (N_4171,N_3691,N_3903);
and U4172 (N_4172,N_3743,N_3686);
or U4173 (N_4173,N_3986,N_3875);
nand U4174 (N_4174,N_3764,N_3933);
or U4175 (N_4175,N_3876,N_3798);
or U4176 (N_4176,N_3938,N_3681);
xor U4177 (N_4177,N_3821,N_3727);
xnor U4178 (N_4178,N_3922,N_3980);
nand U4179 (N_4179,N_3960,N_3646);
xor U4180 (N_4180,N_3925,N_3851);
nor U4181 (N_4181,N_3905,N_3638);
nor U4182 (N_4182,N_3839,N_3844);
nand U4183 (N_4183,N_3864,N_3843);
nand U4184 (N_4184,N_3958,N_3969);
xor U4185 (N_4185,N_3642,N_3928);
nand U4186 (N_4186,N_3787,N_3854);
xor U4187 (N_4187,N_3991,N_3927);
or U4188 (N_4188,N_3662,N_3610);
and U4189 (N_4189,N_3808,N_3934);
nor U4190 (N_4190,N_3967,N_3877);
nand U4191 (N_4191,N_3620,N_3742);
nand U4192 (N_4192,N_3907,N_3861);
or U4193 (N_4193,N_3837,N_3721);
xor U4194 (N_4194,N_3942,N_3661);
nand U4195 (N_4195,N_3858,N_3775);
nand U4196 (N_4196,N_3841,N_3846);
nor U4197 (N_4197,N_3615,N_3998);
nor U4198 (N_4198,N_3741,N_3853);
or U4199 (N_4199,N_3950,N_3680);
and U4200 (N_4200,N_3876,N_3746);
and U4201 (N_4201,N_3700,N_3965);
nor U4202 (N_4202,N_3962,N_3644);
and U4203 (N_4203,N_3636,N_3906);
and U4204 (N_4204,N_3868,N_3717);
nor U4205 (N_4205,N_3948,N_3946);
nand U4206 (N_4206,N_3940,N_3901);
nand U4207 (N_4207,N_3810,N_3702);
or U4208 (N_4208,N_3663,N_3676);
or U4209 (N_4209,N_3756,N_3702);
or U4210 (N_4210,N_3997,N_3905);
xnor U4211 (N_4211,N_3653,N_3668);
nand U4212 (N_4212,N_3697,N_3816);
xnor U4213 (N_4213,N_3901,N_3855);
nand U4214 (N_4214,N_3785,N_3679);
or U4215 (N_4215,N_3796,N_3982);
xor U4216 (N_4216,N_3699,N_3659);
nor U4217 (N_4217,N_3770,N_3875);
or U4218 (N_4218,N_3801,N_3868);
nor U4219 (N_4219,N_3691,N_3661);
and U4220 (N_4220,N_3922,N_3710);
or U4221 (N_4221,N_3797,N_3784);
and U4222 (N_4222,N_3759,N_3941);
nand U4223 (N_4223,N_3761,N_3847);
nand U4224 (N_4224,N_3954,N_3976);
and U4225 (N_4225,N_3631,N_3610);
nor U4226 (N_4226,N_3646,N_3680);
xor U4227 (N_4227,N_3868,N_3795);
and U4228 (N_4228,N_3948,N_3688);
xnor U4229 (N_4229,N_3931,N_3873);
and U4230 (N_4230,N_3690,N_3996);
or U4231 (N_4231,N_3897,N_3801);
nor U4232 (N_4232,N_3976,N_3673);
xor U4233 (N_4233,N_3868,N_3931);
or U4234 (N_4234,N_3695,N_3976);
nand U4235 (N_4235,N_3994,N_3651);
xor U4236 (N_4236,N_3980,N_3622);
and U4237 (N_4237,N_3704,N_3762);
nor U4238 (N_4238,N_3925,N_3723);
xor U4239 (N_4239,N_3991,N_3926);
xor U4240 (N_4240,N_3704,N_3702);
or U4241 (N_4241,N_3941,N_3775);
or U4242 (N_4242,N_3766,N_3715);
xnor U4243 (N_4243,N_3678,N_3954);
and U4244 (N_4244,N_3872,N_3878);
or U4245 (N_4245,N_3866,N_3637);
or U4246 (N_4246,N_3656,N_3616);
nor U4247 (N_4247,N_3683,N_3710);
and U4248 (N_4248,N_3910,N_3984);
and U4249 (N_4249,N_3965,N_3959);
or U4250 (N_4250,N_3600,N_3604);
or U4251 (N_4251,N_3937,N_3700);
xnor U4252 (N_4252,N_3902,N_3659);
and U4253 (N_4253,N_3829,N_3673);
nor U4254 (N_4254,N_3991,N_3625);
and U4255 (N_4255,N_3797,N_3665);
xor U4256 (N_4256,N_3691,N_3803);
xor U4257 (N_4257,N_3733,N_3896);
or U4258 (N_4258,N_3885,N_3767);
or U4259 (N_4259,N_3904,N_3613);
or U4260 (N_4260,N_3898,N_3735);
nor U4261 (N_4261,N_3891,N_3977);
xor U4262 (N_4262,N_3924,N_3997);
or U4263 (N_4263,N_3682,N_3728);
nand U4264 (N_4264,N_3924,N_3859);
nand U4265 (N_4265,N_3843,N_3996);
xnor U4266 (N_4266,N_3927,N_3767);
xnor U4267 (N_4267,N_3823,N_3665);
nand U4268 (N_4268,N_3784,N_3767);
or U4269 (N_4269,N_3699,N_3644);
nor U4270 (N_4270,N_3677,N_3721);
nand U4271 (N_4271,N_3993,N_3881);
nor U4272 (N_4272,N_3826,N_3916);
xnor U4273 (N_4273,N_3737,N_3803);
or U4274 (N_4274,N_3946,N_3961);
nor U4275 (N_4275,N_3943,N_3804);
and U4276 (N_4276,N_3710,N_3602);
nor U4277 (N_4277,N_3821,N_3932);
nand U4278 (N_4278,N_3666,N_3692);
or U4279 (N_4279,N_3832,N_3960);
xnor U4280 (N_4280,N_3836,N_3754);
xor U4281 (N_4281,N_3982,N_3701);
or U4282 (N_4282,N_3670,N_3997);
xor U4283 (N_4283,N_3778,N_3652);
nand U4284 (N_4284,N_3632,N_3833);
or U4285 (N_4285,N_3694,N_3917);
or U4286 (N_4286,N_3884,N_3828);
or U4287 (N_4287,N_3810,N_3801);
nor U4288 (N_4288,N_3619,N_3643);
nand U4289 (N_4289,N_3656,N_3689);
xor U4290 (N_4290,N_3926,N_3728);
nand U4291 (N_4291,N_3614,N_3813);
xnor U4292 (N_4292,N_3719,N_3628);
nor U4293 (N_4293,N_3849,N_3961);
and U4294 (N_4294,N_3758,N_3948);
nor U4295 (N_4295,N_3631,N_3968);
nand U4296 (N_4296,N_3609,N_3966);
xnor U4297 (N_4297,N_3707,N_3652);
nand U4298 (N_4298,N_3676,N_3875);
nand U4299 (N_4299,N_3902,N_3629);
xor U4300 (N_4300,N_3768,N_3887);
nand U4301 (N_4301,N_3974,N_3862);
nand U4302 (N_4302,N_3658,N_3724);
xor U4303 (N_4303,N_3693,N_3983);
xnor U4304 (N_4304,N_3989,N_3870);
nand U4305 (N_4305,N_3669,N_3980);
nand U4306 (N_4306,N_3886,N_3728);
xnor U4307 (N_4307,N_3867,N_3740);
xor U4308 (N_4308,N_3908,N_3776);
nor U4309 (N_4309,N_3687,N_3827);
and U4310 (N_4310,N_3818,N_3784);
or U4311 (N_4311,N_3818,N_3888);
nor U4312 (N_4312,N_3878,N_3738);
and U4313 (N_4313,N_3686,N_3784);
or U4314 (N_4314,N_3764,N_3958);
xor U4315 (N_4315,N_3682,N_3621);
or U4316 (N_4316,N_3870,N_3896);
or U4317 (N_4317,N_3804,N_3603);
nand U4318 (N_4318,N_3995,N_3679);
nand U4319 (N_4319,N_3804,N_3744);
xnor U4320 (N_4320,N_3696,N_3798);
nor U4321 (N_4321,N_3788,N_3997);
nor U4322 (N_4322,N_3608,N_3916);
nand U4323 (N_4323,N_3915,N_3691);
or U4324 (N_4324,N_3963,N_3856);
nand U4325 (N_4325,N_3733,N_3812);
xor U4326 (N_4326,N_3723,N_3763);
and U4327 (N_4327,N_3912,N_3682);
or U4328 (N_4328,N_3656,N_3804);
nand U4329 (N_4329,N_3796,N_3777);
nand U4330 (N_4330,N_3824,N_3893);
nand U4331 (N_4331,N_3997,N_3715);
and U4332 (N_4332,N_3703,N_3981);
nor U4333 (N_4333,N_3872,N_3961);
and U4334 (N_4334,N_3729,N_3979);
nor U4335 (N_4335,N_3823,N_3636);
and U4336 (N_4336,N_3706,N_3764);
and U4337 (N_4337,N_3985,N_3864);
nand U4338 (N_4338,N_3776,N_3739);
xor U4339 (N_4339,N_3918,N_3816);
nand U4340 (N_4340,N_3677,N_3833);
nor U4341 (N_4341,N_3666,N_3647);
or U4342 (N_4342,N_3884,N_3832);
and U4343 (N_4343,N_3972,N_3935);
nand U4344 (N_4344,N_3802,N_3639);
nand U4345 (N_4345,N_3700,N_3881);
and U4346 (N_4346,N_3885,N_3772);
or U4347 (N_4347,N_3928,N_3874);
nor U4348 (N_4348,N_3606,N_3745);
nand U4349 (N_4349,N_3778,N_3937);
and U4350 (N_4350,N_3870,N_3654);
nor U4351 (N_4351,N_3760,N_3621);
or U4352 (N_4352,N_3800,N_3775);
nor U4353 (N_4353,N_3875,N_3790);
nor U4354 (N_4354,N_3703,N_3625);
xor U4355 (N_4355,N_3931,N_3635);
nand U4356 (N_4356,N_3701,N_3868);
and U4357 (N_4357,N_3811,N_3610);
nand U4358 (N_4358,N_3615,N_3708);
nand U4359 (N_4359,N_3606,N_3982);
nor U4360 (N_4360,N_3890,N_3690);
nor U4361 (N_4361,N_3823,N_3694);
or U4362 (N_4362,N_3932,N_3872);
nand U4363 (N_4363,N_3707,N_3828);
nor U4364 (N_4364,N_3625,N_3949);
nor U4365 (N_4365,N_3649,N_3846);
or U4366 (N_4366,N_3736,N_3889);
xnor U4367 (N_4367,N_3681,N_3964);
and U4368 (N_4368,N_3651,N_3774);
nor U4369 (N_4369,N_3801,N_3974);
or U4370 (N_4370,N_3641,N_3815);
or U4371 (N_4371,N_3819,N_3991);
and U4372 (N_4372,N_3946,N_3697);
nand U4373 (N_4373,N_3820,N_3986);
nor U4374 (N_4374,N_3698,N_3970);
nor U4375 (N_4375,N_3781,N_3696);
and U4376 (N_4376,N_3874,N_3636);
xnor U4377 (N_4377,N_3855,N_3682);
xor U4378 (N_4378,N_3772,N_3692);
or U4379 (N_4379,N_3840,N_3627);
or U4380 (N_4380,N_3874,N_3953);
nor U4381 (N_4381,N_3963,N_3900);
nand U4382 (N_4382,N_3816,N_3748);
nor U4383 (N_4383,N_3719,N_3906);
nand U4384 (N_4384,N_3802,N_3671);
nand U4385 (N_4385,N_3938,N_3929);
or U4386 (N_4386,N_3837,N_3977);
nand U4387 (N_4387,N_3687,N_3885);
and U4388 (N_4388,N_3984,N_3972);
or U4389 (N_4389,N_3819,N_3648);
and U4390 (N_4390,N_3830,N_3668);
or U4391 (N_4391,N_3737,N_3659);
nor U4392 (N_4392,N_3722,N_3620);
or U4393 (N_4393,N_3617,N_3642);
and U4394 (N_4394,N_3972,N_3937);
or U4395 (N_4395,N_3642,N_3673);
nand U4396 (N_4396,N_3654,N_3774);
nor U4397 (N_4397,N_3732,N_3889);
nor U4398 (N_4398,N_3976,N_3888);
xnor U4399 (N_4399,N_3602,N_3999);
nor U4400 (N_4400,N_4243,N_4042);
nand U4401 (N_4401,N_4156,N_4031);
nor U4402 (N_4402,N_4365,N_4111);
and U4403 (N_4403,N_4226,N_4179);
and U4404 (N_4404,N_4159,N_4232);
nand U4405 (N_4405,N_4324,N_4277);
xor U4406 (N_4406,N_4257,N_4102);
and U4407 (N_4407,N_4290,N_4353);
or U4408 (N_4408,N_4104,N_4278);
nor U4409 (N_4409,N_4009,N_4192);
and U4410 (N_4410,N_4266,N_4363);
xor U4411 (N_4411,N_4237,N_4040);
or U4412 (N_4412,N_4078,N_4381);
xnor U4413 (N_4413,N_4044,N_4183);
nor U4414 (N_4414,N_4119,N_4005);
xor U4415 (N_4415,N_4215,N_4197);
and U4416 (N_4416,N_4173,N_4082);
xnor U4417 (N_4417,N_4108,N_4316);
nand U4418 (N_4418,N_4357,N_4045);
nor U4419 (N_4419,N_4331,N_4393);
nand U4420 (N_4420,N_4354,N_4137);
nor U4421 (N_4421,N_4304,N_4050);
xnor U4422 (N_4422,N_4340,N_4129);
or U4423 (N_4423,N_4067,N_4329);
nand U4424 (N_4424,N_4010,N_4072);
or U4425 (N_4425,N_4207,N_4367);
nor U4426 (N_4426,N_4372,N_4326);
xnor U4427 (N_4427,N_4306,N_4016);
or U4428 (N_4428,N_4336,N_4268);
or U4429 (N_4429,N_4396,N_4246);
or U4430 (N_4430,N_4214,N_4348);
xnor U4431 (N_4431,N_4384,N_4064);
xor U4432 (N_4432,N_4099,N_4377);
xnor U4433 (N_4433,N_4253,N_4218);
xnor U4434 (N_4434,N_4101,N_4039);
nor U4435 (N_4435,N_4149,N_4241);
xnor U4436 (N_4436,N_4299,N_4341);
or U4437 (N_4437,N_4053,N_4093);
xor U4438 (N_4438,N_4202,N_4355);
nor U4439 (N_4439,N_4171,N_4162);
nand U4440 (N_4440,N_4014,N_4313);
nand U4441 (N_4441,N_4032,N_4375);
xor U4442 (N_4442,N_4100,N_4066);
nor U4443 (N_4443,N_4398,N_4263);
and U4444 (N_4444,N_4325,N_4164);
xor U4445 (N_4445,N_4323,N_4081);
nor U4446 (N_4446,N_4392,N_4086);
nor U4447 (N_4447,N_4302,N_4186);
nand U4448 (N_4448,N_4388,N_4228);
nand U4449 (N_4449,N_4395,N_4017);
nor U4450 (N_4450,N_4062,N_4151);
xor U4451 (N_4451,N_4288,N_4110);
nor U4452 (N_4452,N_4131,N_4085);
and U4453 (N_4453,N_4293,N_4282);
or U4454 (N_4454,N_4090,N_4153);
nor U4455 (N_4455,N_4168,N_4223);
nor U4456 (N_4456,N_4285,N_4198);
or U4457 (N_4457,N_4008,N_4115);
and U4458 (N_4458,N_4335,N_4224);
nand U4459 (N_4459,N_4125,N_4112);
and U4460 (N_4460,N_4056,N_4175);
and U4461 (N_4461,N_4387,N_4206);
xor U4462 (N_4462,N_4296,N_4004);
nand U4463 (N_4463,N_4035,N_4174);
nand U4464 (N_4464,N_4264,N_4330);
nor U4465 (N_4465,N_4244,N_4318);
and U4466 (N_4466,N_4087,N_4034);
nand U4467 (N_4467,N_4126,N_4231);
nand U4468 (N_4468,N_4194,N_4320);
xor U4469 (N_4469,N_4158,N_4128);
nand U4470 (N_4470,N_4369,N_4059);
xnor U4471 (N_4471,N_4201,N_4233);
or U4472 (N_4472,N_4028,N_4091);
nor U4473 (N_4473,N_4127,N_4216);
nor U4474 (N_4474,N_4310,N_4200);
nand U4475 (N_4475,N_4250,N_4184);
nand U4476 (N_4476,N_4176,N_4230);
xnor U4477 (N_4477,N_4238,N_4141);
and U4478 (N_4478,N_4148,N_4006);
nor U4479 (N_4479,N_4220,N_4178);
nor U4480 (N_4480,N_4360,N_4023);
and U4481 (N_4481,N_4029,N_4261);
or U4482 (N_4482,N_4182,N_4048);
or U4483 (N_4483,N_4358,N_4275);
xnor U4484 (N_4484,N_4350,N_4265);
nand U4485 (N_4485,N_4113,N_4105);
nor U4486 (N_4486,N_4322,N_4297);
xnor U4487 (N_4487,N_4181,N_4037);
and U4488 (N_4488,N_4152,N_4366);
and U4489 (N_4489,N_4361,N_4191);
or U4490 (N_4490,N_4076,N_4060);
or U4491 (N_4491,N_4143,N_4254);
and U4492 (N_4492,N_4150,N_4189);
xnor U4493 (N_4493,N_4002,N_4283);
nor U4494 (N_4494,N_4052,N_4321);
xor U4495 (N_4495,N_4287,N_4356);
nor U4496 (N_4496,N_4172,N_4041);
or U4497 (N_4497,N_4196,N_4139);
and U4498 (N_4498,N_4227,N_4291);
nor U4499 (N_4499,N_4209,N_4012);
and U4500 (N_4500,N_4077,N_4258);
nor U4501 (N_4501,N_4373,N_4122);
nor U4502 (N_4502,N_4222,N_4269);
and U4503 (N_4503,N_4272,N_4145);
nand U4504 (N_4504,N_4146,N_4364);
nand U4505 (N_4505,N_4003,N_4276);
or U4506 (N_4506,N_4020,N_4382);
nor U4507 (N_4507,N_4133,N_4368);
or U4508 (N_4508,N_4301,N_4177);
or U4509 (N_4509,N_4300,N_4051);
nand U4510 (N_4510,N_4088,N_4245);
xnor U4511 (N_4511,N_4351,N_4021);
and U4512 (N_4512,N_4347,N_4147);
xor U4513 (N_4513,N_4309,N_4225);
or U4514 (N_4514,N_4134,N_4057);
or U4515 (N_4515,N_4095,N_4007);
xor U4516 (N_4516,N_4397,N_4024);
nand U4517 (N_4517,N_4074,N_4080);
or U4518 (N_4518,N_4109,N_4235);
xor U4519 (N_4519,N_4312,N_4289);
or U4520 (N_4520,N_4180,N_4219);
xor U4521 (N_4521,N_4170,N_4036);
or U4522 (N_4522,N_4294,N_4308);
or U4523 (N_4523,N_4063,N_4169);
nor U4524 (N_4524,N_4157,N_4092);
nor U4525 (N_4525,N_4383,N_4185);
or U4526 (N_4526,N_4025,N_4096);
xor U4527 (N_4527,N_4305,N_4259);
nand U4528 (N_4528,N_4281,N_4135);
or U4529 (N_4529,N_4061,N_4075);
xor U4530 (N_4530,N_4339,N_4187);
and U4531 (N_4531,N_4089,N_4084);
nand U4532 (N_4532,N_4103,N_4199);
nand U4533 (N_4533,N_4252,N_4116);
or U4534 (N_4534,N_4352,N_4047);
and U4535 (N_4535,N_4274,N_4097);
or U4536 (N_4536,N_4251,N_4391);
xnor U4537 (N_4537,N_4120,N_4065);
nor U4538 (N_4538,N_4279,N_4247);
nand U4539 (N_4539,N_4132,N_4221);
xor U4540 (N_4540,N_4188,N_4195);
nand U4541 (N_4541,N_4190,N_4026);
nor U4542 (N_4542,N_4015,N_4155);
or U4543 (N_4543,N_4255,N_4121);
or U4544 (N_4544,N_4140,N_4208);
nand U4545 (N_4545,N_4114,N_4362);
or U4546 (N_4546,N_4046,N_4205);
xnor U4547 (N_4547,N_4163,N_4071);
nor U4548 (N_4548,N_4385,N_4286);
or U4549 (N_4549,N_4033,N_4271);
xnor U4550 (N_4550,N_4142,N_4314);
nor U4551 (N_4551,N_4079,N_4055);
and U4552 (N_4552,N_4211,N_4049);
xor U4553 (N_4553,N_4248,N_4166);
nand U4554 (N_4554,N_4043,N_4013);
xor U4555 (N_4555,N_4107,N_4344);
and U4556 (N_4556,N_4027,N_4068);
nor U4557 (N_4557,N_4193,N_4307);
xnor U4558 (N_4558,N_4019,N_4386);
nand U4559 (N_4559,N_4073,N_4338);
nand U4560 (N_4560,N_4349,N_4117);
xor U4561 (N_4561,N_4160,N_4379);
nand U4562 (N_4562,N_4001,N_4124);
nand U4563 (N_4563,N_4376,N_4240);
xor U4564 (N_4564,N_4203,N_4311);
nand U4565 (N_4565,N_4022,N_4298);
nor U4566 (N_4566,N_4249,N_4260);
or U4567 (N_4567,N_4346,N_4378);
and U4568 (N_4568,N_4236,N_4242);
nand U4569 (N_4569,N_4371,N_4030);
nor U4570 (N_4570,N_4123,N_4167);
or U4571 (N_4571,N_4210,N_4234);
and U4572 (N_4572,N_4018,N_4038);
nand U4573 (N_4573,N_4327,N_4098);
and U4574 (N_4574,N_4267,N_4273);
nor U4575 (N_4575,N_4165,N_4239);
nand U4576 (N_4576,N_4328,N_4334);
or U4577 (N_4577,N_4144,N_4058);
xor U4578 (N_4578,N_4292,N_4136);
nor U4579 (N_4579,N_4317,N_4342);
nor U4580 (N_4580,N_4399,N_4315);
nand U4581 (N_4581,N_4161,N_4343);
and U4582 (N_4582,N_4070,N_4106);
nand U4583 (N_4583,N_4295,N_4138);
nand U4584 (N_4584,N_4332,N_4212);
xnor U4585 (N_4585,N_4000,N_4213);
or U4586 (N_4586,N_4094,N_4130);
xnor U4587 (N_4587,N_4204,N_4270);
or U4588 (N_4588,N_4256,N_4217);
and U4589 (N_4589,N_4069,N_4374);
nor U4590 (N_4590,N_4118,N_4389);
or U4591 (N_4591,N_4345,N_4280);
and U4592 (N_4592,N_4337,N_4333);
or U4593 (N_4593,N_4303,N_4359);
xnor U4594 (N_4594,N_4319,N_4083);
nand U4595 (N_4595,N_4284,N_4390);
nor U4596 (N_4596,N_4262,N_4011);
and U4597 (N_4597,N_4054,N_4154);
or U4598 (N_4598,N_4370,N_4394);
and U4599 (N_4599,N_4229,N_4380);
and U4600 (N_4600,N_4326,N_4285);
and U4601 (N_4601,N_4345,N_4105);
and U4602 (N_4602,N_4060,N_4168);
xnor U4603 (N_4603,N_4345,N_4352);
and U4604 (N_4604,N_4065,N_4207);
nand U4605 (N_4605,N_4370,N_4072);
nand U4606 (N_4606,N_4068,N_4113);
xor U4607 (N_4607,N_4330,N_4333);
nor U4608 (N_4608,N_4233,N_4085);
nor U4609 (N_4609,N_4056,N_4378);
nand U4610 (N_4610,N_4105,N_4098);
nor U4611 (N_4611,N_4274,N_4207);
and U4612 (N_4612,N_4365,N_4094);
xor U4613 (N_4613,N_4066,N_4106);
nand U4614 (N_4614,N_4308,N_4149);
xnor U4615 (N_4615,N_4288,N_4139);
xor U4616 (N_4616,N_4351,N_4062);
nor U4617 (N_4617,N_4256,N_4258);
nand U4618 (N_4618,N_4277,N_4362);
and U4619 (N_4619,N_4083,N_4344);
xnor U4620 (N_4620,N_4206,N_4398);
and U4621 (N_4621,N_4255,N_4366);
nor U4622 (N_4622,N_4132,N_4164);
or U4623 (N_4623,N_4306,N_4252);
nand U4624 (N_4624,N_4004,N_4209);
and U4625 (N_4625,N_4101,N_4246);
xnor U4626 (N_4626,N_4265,N_4299);
nand U4627 (N_4627,N_4233,N_4126);
and U4628 (N_4628,N_4163,N_4328);
xor U4629 (N_4629,N_4316,N_4154);
and U4630 (N_4630,N_4059,N_4164);
or U4631 (N_4631,N_4295,N_4343);
and U4632 (N_4632,N_4327,N_4083);
nor U4633 (N_4633,N_4192,N_4282);
and U4634 (N_4634,N_4042,N_4127);
nor U4635 (N_4635,N_4199,N_4283);
xor U4636 (N_4636,N_4030,N_4104);
nor U4637 (N_4637,N_4042,N_4360);
nor U4638 (N_4638,N_4173,N_4061);
and U4639 (N_4639,N_4060,N_4086);
nor U4640 (N_4640,N_4028,N_4058);
xor U4641 (N_4641,N_4379,N_4251);
or U4642 (N_4642,N_4339,N_4261);
nand U4643 (N_4643,N_4207,N_4063);
and U4644 (N_4644,N_4085,N_4368);
or U4645 (N_4645,N_4298,N_4381);
and U4646 (N_4646,N_4109,N_4388);
nor U4647 (N_4647,N_4001,N_4174);
xnor U4648 (N_4648,N_4177,N_4299);
xor U4649 (N_4649,N_4205,N_4271);
nand U4650 (N_4650,N_4053,N_4092);
nor U4651 (N_4651,N_4344,N_4182);
nand U4652 (N_4652,N_4069,N_4079);
nor U4653 (N_4653,N_4379,N_4105);
nand U4654 (N_4654,N_4349,N_4307);
and U4655 (N_4655,N_4040,N_4096);
and U4656 (N_4656,N_4232,N_4391);
nor U4657 (N_4657,N_4366,N_4003);
nor U4658 (N_4658,N_4214,N_4216);
nand U4659 (N_4659,N_4363,N_4359);
xor U4660 (N_4660,N_4387,N_4081);
nor U4661 (N_4661,N_4313,N_4230);
or U4662 (N_4662,N_4369,N_4392);
or U4663 (N_4663,N_4245,N_4204);
and U4664 (N_4664,N_4144,N_4298);
nand U4665 (N_4665,N_4311,N_4362);
nor U4666 (N_4666,N_4212,N_4314);
or U4667 (N_4667,N_4175,N_4124);
or U4668 (N_4668,N_4063,N_4205);
nand U4669 (N_4669,N_4279,N_4059);
nand U4670 (N_4670,N_4027,N_4245);
or U4671 (N_4671,N_4385,N_4089);
nor U4672 (N_4672,N_4127,N_4093);
or U4673 (N_4673,N_4309,N_4179);
nor U4674 (N_4674,N_4227,N_4354);
nand U4675 (N_4675,N_4332,N_4186);
nand U4676 (N_4676,N_4246,N_4382);
and U4677 (N_4677,N_4279,N_4232);
and U4678 (N_4678,N_4280,N_4306);
or U4679 (N_4679,N_4176,N_4059);
nand U4680 (N_4680,N_4011,N_4241);
and U4681 (N_4681,N_4310,N_4090);
xnor U4682 (N_4682,N_4316,N_4130);
nand U4683 (N_4683,N_4136,N_4285);
nand U4684 (N_4684,N_4352,N_4073);
nand U4685 (N_4685,N_4313,N_4036);
or U4686 (N_4686,N_4113,N_4352);
xnor U4687 (N_4687,N_4122,N_4382);
nand U4688 (N_4688,N_4367,N_4301);
nor U4689 (N_4689,N_4384,N_4241);
and U4690 (N_4690,N_4027,N_4137);
nand U4691 (N_4691,N_4291,N_4212);
nand U4692 (N_4692,N_4227,N_4050);
nand U4693 (N_4693,N_4375,N_4022);
nor U4694 (N_4694,N_4113,N_4297);
nand U4695 (N_4695,N_4263,N_4187);
nor U4696 (N_4696,N_4331,N_4042);
xor U4697 (N_4697,N_4113,N_4003);
xnor U4698 (N_4698,N_4256,N_4146);
nor U4699 (N_4699,N_4388,N_4334);
xnor U4700 (N_4700,N_4282,N_4261);
xnor U4701 (N_4701,N_4396,N_4017);
nor U4702 (N_4702,N_4005,N_4234);
xnor U4703 (N_4703,N_4177,N_4307);
nand U4704 (N_4704,N_4036,N_4271);
or U4705 (N_4705,N_4322,N_4254);
or U4706 (N_4706,N_4120,N_4079);
and U4707 (N_4707,N_4384,N_4317);
xor U4708 (N_4708,N_4190,N_4119);
and U4709 (N_4709,N_4040,N_4346);
nor U4710 (N_4710,N_4268,N_4247);
xor U4711 (N_4711,N_4079,N_4285);
or U4712 (N_4712,N_4171,N_4167);
nand U4713 (N_4713,N_4125,N_4244);
nand U4714 (N_4714,N_4292,N_4087);
and U4715 (N_4715,N_4359,N_4156);
nor U4716 (N_4716,N_4231,N_4009);
and U4717 (N_4717,N_4177,N_4098);
nor U4718 (N_4718,N_4308,N_4329);
xnor U4719 (N_4719,N_4240,N_4160);
nor U4720 (N_4720,N_4035,N_4086);
nor U4721 (N_4721,N_4332,N_4358);
nor U4722 (N_4722,N_4288,N_4042);
nand U4723 (N_4723,N_4084,N_4332);
nor U4724 (N_4724,N_4174,N_4387);
xnor U4725 (N_4725,N_4389,N_4114);
xor U4726 (N_4726,N_4145,N_4118);
or U4727 (N_4727,N_4105,N_4299);
nor U4728 (N_4728,N_4392,N_4376);
and U4729 (N_4729,N_4155,N_4217);
or U4730 (N_4730,N_4158,N_4223);
nor U4731 (N_4731,N_4337,N_4080);
or U4732 (N_4732,N_4304,N_4220);
xnor U4733 (N_4733,N_4122,N_4236);
nand U4734 (N_4734,N_4122,N_4144);
or U4735 (N_4735,N_4289,N_4069);
xnor U4736 (N_4736,N_4067,N_4391);
and U4737 (N_4737,N_4035,N_4278);
or U4738 (N_4738,N_4086,N_4209);
xor U4739 (N_4739,N_4152,N_4242);
nor U4740 (N_4740,N_4015,N_4237);
and U4741 (N_4741,N_4278,N_4024);
nor U4742 (N_4742,N_4189,N_4132);
nor U4743 (N_4743,N_4364,N_4116);
nor U4744 (N_4744,N_4247,N_4397);
nand U4745 (N_4745,N_4352,N_4194);
xnor U4746 (N_4746,N_4077,N_4351);
or U4747 (N_4747,N_4342,N_4259);
nor U4748 (N_4748,N_4225,N_4226);
xor U4749 (N_4749,N_4286,N_4156);
nand U4750 (N_4750,N_4251,N_4042);
xnor U4751 (N_4751,N_4050,N_4060);
nor U4752 (N_4752,N_4182,N_4188);
or U4753 (N_4753,N_4323,N_4056);
or U4754 (N_4754,N_4141,N_4047);
and U4755 (N_4755,N_4164,N_4099);
and U4756 (N_4756,N_4148,N_4250);
and U4757 (N_4757,N_4388,N_4071);
xor U4758 (N_4758,N_4068,N_4152);
nor U4759 (N_4759,N_4042,N_4060);
nand U4760 (N_4760,N_4036,N_4175);
or U4761 (N_4761,N_4014,N_4324);
nor U4762 (N_4762,N_4022,N_4010);
and U4763 (N_4763,N_4090,N_4003);
xor U4764 (N_4764,N_4206,N_4092);
or U4765 (N_4765,N_4267,N_4042);
nand U4766 (N_4766,N_4026,N_4123);
nor U4767 (N_4767,N_4359,N_4308);
nor U4768 (N_4768,N_4061,N_4086);
and U4769 (N_4769,N_4125,N_4153);
nand U4770 (N_4770,N_4348,N_4390);
nor U4771 (N_4771,N_4288,N_4038);
or U4772 (N_4772,N_4265,N_4201);
xor U4773 (N_4773,N_4268,N_4019);
nor U4774 (N_4774,N_4337,N_4096);
and U4775 (N_4775,N_4206,N_4178);
nor U4776 (N_4776,N_4138,N_4077);
or U4777 (N_4777,N_4110,N_4359);
or U4778 (N_4778,N_4199,N_4154);
or U4779 (N_4779,N_4110,N_4014);
or U4780 (N_4780,N_4033,N_4029);
nand U4781 (N_4781,N_4147,N_4050);
nor U4782 (N_4782,N_4388,N_4235);
xor U4783 (N_4783,N_4306,N_4305);
or U4784 (N_4784,N_4311,N_4027);
nand U4785 (N_4785,N_4234,N_4023);
xnor U4786 (N_4786,N_4230,N_4165);
nand U4787 (N_4787,N_4049,N_4271);
nand U4788 (N_4788,N_4136,N_4383);
nand U4789 (N_4789,N_4363,N_4178);
nand U4790 (N_4790,N_4337,N_4338);
nor U4791 (N_4791,N_4317,N_4059);
nand U4792 (N_4792,N_4311,N_4210);
or U4793 (N_4793,N_4255,N_4010);
nor U4794 (N_4794,N_4033,N_4344);
nor U4795 (N_4795,N_4141,N_4261);
nand U4796 (N_4796,N_4150,N_4332);
nand U4797 (N_4797,N_4386,N_4084);
xor U4798 (N_4798,N_4067,N_4342);
and U4799 (N_4799,N_4315,N_4244);
nand U4800 (N_4800,N_4640,N_4685);
nor U4801 (N_4801,N_4686,N_4474);
xnor U4802 (N_4802,N_4653,N_4597);
xor U4803 (N_4803,N_4538,N_4529);
and U4804 (N_4804,N_4795,N_4649);
or U4805 (N_4805,N_4794,N_4603);
nand U4806 (N_4806,N_4576,N_4430);
xnor U4807 (N_4807,N_4413,N_4532);
and U4808 (N_4808,N_4674,N_4728);
or U4809 (N_4809,N_4475,N_4444);
and U4810 (N_4810,N_4664,N_4652);
xor U4811 (N_4811,N_4406,N_4564);
nand U4812 (N_4812,N_4676,N_4735);
nor U4813 (N_4813,N_4566,N_4447);
xor U4814 (N_4814,N_4672,N_4575);
xor U4815 (N_4815,N_4446,N_4691);
and U4816 (N_4816,N_4524,N_4675);
and U4817 (N_4817,N_4680,N_4767);
nand U4818 (N_4818,N_4527,N_4762);
or U4819 (N_4819,N_4556,N_4561);
xor U4820 (N_4820,N_4559,N_4707);
xnor U4821 (N_4821,N_4678,N_4623);
xnor U4822 (N_4822,N_4695,N_4582);
nor U4823 (N_4823,N_4421,N_4694);
nand U4824 (N_4824,N_4687,N_4494);
nor U4825 (N_4825,N_4468,N_4470);
nor U4826 (N_4826,N_4791,N_4591);
and U4827 (N_4827,N_4534,N_4551);
or U4828 (N_4828,N_4788,N_4454);
and U4829 (N_4829,N_4429,N_4688);
nor U4830 (N_4830,N_4585,N_4417);
nand U4831 (N_4831,N_4528,N_4700);
nor U4832 (N_4832,N_4544,N_4659);
nand U4833 (N_4833,N_4478,N_4477);
nand U4834 (N_4834,N_4753,N_4658);
and U4835 (N_4835,N_4772,N_4626);
nor U4836 (N_4836,N_4628,N_4606);
or U4837 (N_4837,N_4655,N_4460);
nand U4838 (N_4838,N_4441,N_4634);
xor U4839 (N_4839,N_4755,N_4630);
nand U4840 (N_4840,N_4706,N_4761);
and U4841 (N_4841,N_4732,N_4537);
nand U4842 (N_4842,N_4426,N_4458);
nand U4843 (N_4843,N_4504,N_4785);
xor U4844 (N_4844,N_4784,N_4642);
nor U4845 (N_4845,N_4765,N_4701);
nand U4846 (N_4846,N_4486,N_4774);
xnor U4847 (N_4847,N_4496,N_4693);
nand U4848 (N_4848,N_4547,N_4548);
xor U4849 (N_4849,N_4799,N_4609);
xor U4850 (N_4850,N_4500,N_4648);
nand U4851 (N_4851,N_4433,N_4667);
and U4852 (N_4852,N_4673,N_4565);
and U4853 (N_4853,N_4419,N_4773);
or U4854 (N_4854,N_4593,N_4711);
xor U4855 (N_4855,N_4793,N_4736);
xor U4856 (N_4856,N_4594,N_4748);
nor U4857 (N_4857,N_4646,N_4714);
nand U4858 (N_4858,N_4572,N_4747);
nor U4859 (N_4859,N_4465,N_4440);
or U4860 (N_4860,N_4432,N_4487);
nor U4861 (N_4861,N_4668,N_4493);
nor U4862 (N_4862,N_4407,N_4450);
nand U4863 (N_4863,N_4490,N_4457);
or U4864 (N_4864,N_4567,N_4595);
or U4865 (N_4865,N_4756,N_4438);
nor U4866 (N_4866,N_4560,N_4779);
nor U4867 (N_4867,N_4611,N_4645);
nor U4868 (N_4868,N_4778,N_4553);
and U4869 (N_4869,N_4427,N_4546);
nand U4870 (N_4870,N_4671,N_4545);
xnor U4871 (N_4871,N_4550,N_4428);
nor U4872 (N_4872,N_4453,N_4643);
xnor U4873 (N_4873,N_4589,N_4635);
nor U4874 (N_4874,N_4758,N_4618);
nand U4875 (N_4875,N_4411,N_4510);
nor U4876 (N_4876,N_4592,N_4746);
nand U4877 (N_4877,N_4776,N_4709);
xnor U4878 (N_4878,N_4400,N_4721);
and U4879 (N_4879,N_4627,N_4768);
xnor U4880 (N_4880,N_4763,N_4410);
and U4881 (N_4881,N_4555,N_4401);
xnor U4882 (N_4882,N_4525,N_4690);
xor U4883 (N_4883,N_4702,N_4608);
or U4884 (N_4884,N_4583,N_4506);
nor U4885 (N_4885,N_4614,N_4734);
nor U4886 (N_4886,N_4619,N_4631);
nor U4887 (N_4887,N_4462,N_4482);
nor U4888 (N_4888,N_4509,N_4770);
nand U4889 (N_4889,N_4459,N_4574);
xor U4890 (N_4890,N_4657,N_4639);
or U4891 (N_4891,N_4666,N_4786);
or U4892 (N_4892,N_4442,N_4577);
xor U4893 (N_4893,N_4520,N_4481);
or U4894 (N_4894,N_4514,N_4483);
nor U4895 (N_4895,N_4604,N_4415);
xor U4896 (N_4896,N_4472,N_4515);
or U4897 (N_4897,N_4435,N_4543);
and U4898 (N_4898,N_4656,N_4495);
nand U4899 (N_4899,N_4719,N_4420);
nand U4900 (N_4900,N_4796,N_4581);
nor U4901 (N_4901,N_4436,N_4650);
xnor U4902 (N_4902,N_4601,N_4713);
nand U4903 (N_4903,N_4610,N_4769);
nor U4904 (N_4904,N_4681,N_4424);
xnor U4905 (N_4905,N_4573,N_4503);
or U4906 (N_4906,N_4705,N_4452);
and U4907 (N_4907,N_4451,N_4729);
nand U4908 (N_4908,N_4521,N_4488);
and U4909 (N_4909,N_4683,N_4703);
xnor U4910 (N_4910,N_4744,N_4530);
nor U4911 (N_4911,N_4775,N_4501);
xor U4912 (N_4912,N_4715,N_4792);
nand U4913 (N_4913,N_4638,N_4743);
and U4914 (N_4914,N_4661,N_4513);
nor U4915 (N_4915,N_4412,N_4760);
or U4916 (N_4916,N_4549,N_4570);
or U4917 (N_4917,N_4689,N_4697);
nor U4918 (N_4918,N_4710,N_4404);
nor U4919 (N_4919,N_4456,N_4605);
or U4920 (N_4920,N_4699,N_4726);
xnor U4921 (N_4921,N_4662,N_4740);
xor U4922 (N_4922,N_4704,N_4751);
nand U4923 (N_4923,N_4600,N_4539);
nand U4924 (N_4924,N_4750,N_4598);
nor U4925 (N_4925,N_4616,N_4737);
nand U4926 (N_4926,N_4716,N_4562);
nor U4927 (N_4927,N_4422,N_4665);
or U4928 (N_4928,N_4781,N_4588);
nand U4929 (N_4929,N_4502,N_4620);
or U4930 (N_4930,N_4654,N_4522);
nand U4931 (N_4931,N_4759,N_4731);
or U4932 (N_4932,N_4677,N_4787);
nand U4933 (N_4933,N_4612,N_4409);
and U4934 (N_4934,N_4479,N_4484);
and U4935 (N_4935,N_4632,N_4586);
xor U4936 (N_4936,N_4443,N_4717);
nand U4937 (N_4937,N_4679,N_4511);
or U4938 (N_4938,N_4669,N_4599);
nand U4939 (N_4939,N_4602,N_4584);
nand U4940 (N_4940,N_4523,N_4738);
or U4941 (N_4941,N_4449,N_4663);
and U4942 (N_4942,N_4579,N_4590);
or U4943 (N_4943,N_4437,N_4568);
nand U4944 (N_4944,N_4418,N_4749);
and U4945 (N_4945,N_4526,N_4414);
or U4946 (N_4946,N_4764,N_4403);
nor U4947 (N_4947,N_4448,N_4622);
nor U4948 (N_4948,N_4730,N_4464);
xor U4949 (N_4949,N_4512,N_4651);
or U4950 (N_4950,N_4471,N_4423);
nand U4951 (N_4951,N_4624,N_4508);
xnor U4952 (N_4952,N_4480,N_4613);
nor U4953 (N_4953,N_4636,N_4644);
or U4954 (N_4954,N_4402,N_4542);
nand U4955 (N_4955,N_4498,N_4517);
nor U4956 (N_4956,N_4554,N_4684);
xor U4957 (N_4957,N_4596,N_4798);
and U4958 (N_4958,N_4789,N_4416);
nand U4959 (N_4959,N_4754,N_4516);
nand U4960 (N_4960,N_4757,N_4558);
or U4961 (N_4961,N_4629,N_4431);
and U4962 (N_4962,N_4535,N_4797);
nand U4963 (N_4963,N_4720,N_4587);
nor U4964 (N_4964,N_4518,N_4718);
nand U4965 (N_4965,N_4708,N_4557);
and U4966 (N_4966,N_4473,N_4682);
or U4967 (N_4967,N_4445,N_4647);
or U4968 (N_4968,N_4625,N_4771);
nor U4969 (N_4969,N_4461,N_4439);
nor U4970 (N_4970,N_4745,N_4569);
nand U4971 (N_4971,N_4563,N_4497);
and U4972 (N_4972,N_4540,N_4782);
nor U4973 (N_4973,N_4692,N_4742);
nand U4974 (N_4974,N_4466,N_4780);
or U4975 (N_4975,N_4722,N_4507);
nand U4976 (N_4976,N_4536,N_4752);
and U4977 (N_4977,N_4425,N_4790);
nor U4978 (N_4978,N_4485,N_4783);
and U4979 (N_4979,N_4578,N_4476);
and U4980 (N_4980,N_4712,N_4405);
and U4981 (N_4981,N_4660,N_4492);
and U4982 (N_4982,N_4724,N_4725);
and U4983 (N_4983,N_4641,N_4723);
nor U4984 (N_4984,N_4489,N_4607);
nand U4985 (N_4985,N_4615,N_4727);
xor U4986 (N_4986,N_4696,N_4777);
xnor U4987 (N_4987,N_4733,N_4533);
xnor U4988 (N_4988,N_4580,N_4463);
xor U4989 (N_4989,N_4637,N_4467);
or U4990 (N_4990,N_4455,N_4617);
nand U4991 (N_4991,N_4434,N_4698);
nand U4992 (N_4992,N_4571,N_4505);
nor U4993 (N_4993,N_4541,N_4741);
or U4994 (N_4994,N_4633,N_4552);
and U4995 (N_4995,N_4408,N_4739);
and U4996 (N_4996,N_4499,N_4469);
or U4997 (N_4997,N_4766,N_4670);
and U4998 (N_4998,N_4621,N_4519);
or U4999 (N_4999,N_4491,N_4531);
nand U5000 (N_5000,N_4630,N_4561);
nor U5001 (N_5001,N_4426,N_4730);
nand U5002 (N_5002,N_4493,N_4573);
nor U5003 (N_5003,N_4641,N_4758);
nor U5004 (N_5004,N_4521,N_4668);
xnor U5005 (N_5005,N_4749,N_4642);
or U5006 (N_5006,N_4492,N_4468);
xnor U5007 (N_5007,N_4694,N_4707);
nand U5008 (N_5008,N_4566,N_4717);
or U5009 (N_5009,N_4781,N_4443);
nand U5010 (N_5010,N_4564,N_4427);
or U5011 (N_5011,N_4774,N_4648);
nor U5012 (N_5012,N_4666,N_4728);
or U5013 (N_5013,N_4565,N_4483);
nand U5014 (N_5014,N_4606,N_4769);
and U5015 (N_5015,N_4448,N_4763);
or U5016 (N_5016,N_4682,N_4462);
and U5017 (N_5017,N_4562,N_4758);
xnor U5018 (N_5018,N_4404,N_4644);
and U5019 (N_5019,N_4536,N_4534);
nand U5020 (N_5020,N_4770,N_4698);
or U5021 (N_5021,N_4759,N_4525);
nor U5022 (N_5022,N_4401,N_4661);
and U5023 (N_5023,N_4550,N_4632);
and U5024 (N_5024,N_4569,N_4495);
and U5025 (N_5025,N_4598,N_4558);
or U5026 (N_5026,N_4690,N_4418);
or U5027 (N_5027,N_4742,N_4690);
nor U5028 (N_5028,N_4708,N_4499);
or U5029 (N_5029,N_4624,N_4433);
nand U5030 (N_5030,N_4701,N_4461);
or U5031 (N_5031,N_4700,N_4440);
nor U5032 (N_5032,N_4512,N_4603);
nor U5033 (N_5033,N_4606,N_4705);
nor U5034 (N_5034,N_4689,N_4508);
and U5035 (N_5035,N_4721,N_4502);
nor U5036 (N_5036,N_4542,N_4701);
nor U5037 (N_5037,N_4673,N_4738);
or U5038 (N_5038,N_4788,N_4511);
nor U5039 (N_5039,N_4540,N_4757);
xnor U5040 (N_5040,N_4719,N_4795);
nor U5041 (N_5041,N_4750,N_4544);
nand U5042 (N_5042,N_4616,N_4623);
and U5043 (N_5043,N_4700,N_4681);
or U5044 (N_5044,N_4657,N_4401);
nand U5045 (N_5045,N_4768,N_4796);
nand U5046 (N_5046,N_4602,N_4686);
or U5047 (N_5047,N_4516,N_4717);
nor U5048 (N_5048,N_4454,N_4709);
and U5049 (N_5049,N_4761,N_4541);
xor U5050 (N_5050,N_4692,N_4756);
nand U5051 (N_5051,N_4587,N_4487);
and U5052 (N_5052,N_4693,N_4688);
xor U5053 (N_5053,N_4797,N_4571);
or U5054 (N_5054,N_4434,N_4713);
or U5055 (N_5055,N_4453,N_4579);
and U5056 (N_5056,N_4753,N_4610);
and U5057 (N_5057,N_4476,N_4426);
nand U5058 (N_5058,N_4483,N_4411);
or U5059 (N_5059,N_4614,N_4584);
nand U5060 (N_5060,N_4601,N_4563);
xnor U5061 (N_5061,N_4729,N_4420);
nand U5062 (N_5062,N_4426,N_4793);
nor U5063 (N_5063,N_4700,N_4728);
nor U5064 (N_5064,N_4684,N_4426);
or U5065 (N_5065,N_4608,N_4596);
or U5066 (N_5066,N_4623,N_4438);
and U5067 (N_5067,N_4447,N_4730);
nor U5068 (N_5068,N_4529,N_4676);
nor U5069 (N_5069,N_4410,N_4602);
or U5070 (N_5070,N_4527,N_4606);
xor U5071 (N_5071,N_4468,N_4687);
and U5072 (N_5072,N_4672,N_4693);
nand U5073 (N_5073,N_4738,N_4685);
nand U5074 (N_5074,N_4522,N_4722);
or U5075 (N_5075,N_4763,N_4701);
or U5076 (N_5076,N_4618,N_4585);
nand U5077 (N_5077,N_4600,N_4502);
nand U5078 (N_5078,N_4417,N_4522);
xnor U5079 (N_5079,N_4763,N_4685);
nor U5080 (N_5080,N_4598,N_4536);
or U5081 (N_5081,N_4665,N_4400);
nor U5082 (N_5082,N_4733,N_4568);
and U5083 (N_5083,N_4680,N_4540);
and U5084 (N_5084,N_4630,N_4451);
xnor U5085 (N_5085,N_4528,N_4750);
nor U5086 (N_5086,N_4506,N_4695);
or U5087 (N_5087,N_4623,N_4533);
or U5088 (N_5088,N_4721,N_4706);
and U5089 (N_5089,N_4557,N_4788);
xor U5090 (N_5090,N_4778,N_4638);
or U5091 (N_5091,N_4414,N_4600);
nor U5092 (N_5092,N_4564,N_4516);
nor U5093 (N_5093,N_4652,N_4559);
or U5094 (N_5094,N_4774,N_4558);
and U5095 (N_5095,N_4612,N_4514);
nor U5096 (N_5096,N_4565,N_4461);
nand U5097 (N_5097,N_4587,N_4712);
xnor U5098 (N_5098,N_4610,N_4634);
xor U5099 (N_5099,N_4564,N_4694);
or U5100 (N_5100,N_4416,N_4675);
xnor U5101 (N_5101,N_4470,N_4705);
and U5102 (N_5102,N_4509,N_4624);
xnor U5103 (N_5103,N_4466,N_4557);
xnor U5104 (N_5104,N_4439,N_4484);
xnor U5105 (N_5105,N_4607,N_4428);
nand U5106 (N_5106,N_4510,N_4690);
and U5107 (N_5107,N_4786,N_4466);
or U5108 (N_5108,N_4543,N_4606);
xor U5109 (N_5109,N_4730,N_4598);
nand U5110 (N_5110,N_4646,N_4612);
or U5111 (N_5111,N_4500,N_4613);
xor U5112 (N_5112,N_4763,N_4645);
and U5113 (N_5113,N_4716,N_4436);
and U5114 (N_5114,N_4667,N_4462);
nand U5115 (N_5115,N_4464,N_4525);
or U5116 (N_5116,N_4565,N_4581);
nand U5117 (N_5117,N_4425,N_4543);
nor U5118 (N_5118,N_4657,N_4527);
nor U5119 (N_5119,N_4505,N_4647);
and U5120 (N_5120,N_4782,N_4766);
and U5121 (N_5121,N_4684,N_4670);
and U5122 (N_5122,N_4778,N_4449);
xnor U5123 (N_5123,N_4536,N_4469);
or U5124 (N_5124,N_4635,N_4527);
or U5125 (N_5125,N_4431,N_4505);
nor U5126 (N_5126,N_4651,N_4726);
and U5127 (N_5127,N_4771,N_4420);
xor U5128 (N_5128,N_4632,N_4626);
or U5129 (N_5129,N_4622,N_4579);
xor U5130 (N_5130,N_4489,N_4513);
nor U5131 (N_5131,N_4582,N_4458);
or U5132 (N_5132,N_4567,N_4404);
nor U5133 (N_5133,N_4504,N_4534);
or U5134 (N_5134,N_4652,N_4404);
nand U5135 (N_5135,N_4715,N_4520);
and U5136 (N_5136,N_4761,N_4532);
nand U5137 (N_5137,N_4555,N_4413);
and U5138 (N_5138,N_4739,N_4411);
nand U5139 (N_5139,N_4742,N_4707);
nor U5140 (N_5140,N_4491,N_4612);
and U5141 (N_5141,N_4542,N_4405);
nand U5142 (N_5142,N_4460,N_4427);
or U5143 (N_5143,N_4518,N_4748);
xnor U5144 (N_5144,N_4667,N_4736);
nor U5145 (N_5145,N_4438,N_4609);
and U5146 (N_5146,N_4582,N_4405);
nor U5147 (N_5147,N_4532,N_4522);
xnor U5148 (N_5148,N_4687,N_4733);
and U5149 (N_5149,N_4516,N_4683);
nor U5150 (N_5150,N_4419,N_4705);
nor U5151 (N_5151,N_4506,N_4796);
and U5152 (N_5152,N_4666,N_4510);
or U5153 (N_5153,N_4463,N_4445);
xnor U5154 (N_5154,N_4570,N_4441);
or U5155 (N_5155,N_4474,N_4774);
nor U5156 (N_5156,N_4700,N_4763);
nor U5157 (N_5157,N_4661,N_4462);
nor U5158 (N_5158,N_4506,N_4624);
nand U5159 (N_5159,N_4765,N_4689);
or U5160 (N_5160,N_4563,N_4627);
or U5161 (N_5161,N_4794,N_4447);
or U5162 (N_5162,N_4588,N_4661);
nand U5163 (N_5163,N_4673,N_4746);
nand U5164 (N_5164,N_4481,N_4612);
or U5165 (N_5165,N_4581,N_4781);
and U5166 (N_5166,N_4488,N_4589);
and U5167 (N_5167,N_4790,N_4764);
nor U5168 (N_5168,N_4535,N_4412);
nand U5169 (N_5169,N_4580,N_4460);
xor U5170 (N_5170,N_4644,N_4547);
nand U5171 (N_5171,N_4438,N_4619);
and U5172 (N_5172,N_4616,N_4518);
or U5173 (N_5173,N_4730,N_4655);
nand U5174 (N_5174,N_4723,N_4408);
and U5175 (N_5175,N_4643,N_4543);
or U5176 (N_5176,N_4716,N_4480);
nor U5177 (N_5177,N_4574,N_4401);
or U5178 (N_5178,N_4544,N_4640);
xor U5179 (N_5179,N_4549,N_4458);
nand U5180 (N_5180,N_4628,N_4715);
and U5181 (N_5181,N_4683,N_4783);
or U5182 (N_5182,N_4520,N_4429);
or U5183 (N_5183,N_4644,N_4687);
nand U5184 (N_5184,N_4663,N_4675);
and U5185 (N_5185,N_4650,N_4706);
xor U5186 (N_5186,N_4406,N_4560);
or U5187 (N_5187,N_4608,N_4511);
xnor U5188 (N_5188,N_4745,N_4664);
nand U5189 (N_5189,N_4677,N_4641);
nor U5190 (N_5190,N_4460,N_4799);
and U5191 (N_5191,N_4714,N_4532);
nor U5192 (N_5192,N_4786,N_4714);
nand U5193 (N_5193,N_4738,N_4407);
xor U5194 (N_5194,N_4710,N_4719);
xor U5195 (N_5195,N_4407,N_4510);
or U5196 (N_5196,N_4420,N_4529);
or U5197 (N_5197,N_4659,N_4489);
nand U5198 (N_5198,N_4701,N_4716);
and U5199 (N_5199,N_4592,N_4755);
nand U5200 (N_5200,N_4923,N_5198);
and U5201 (N_5201,N_5113,N_4869);
or U5202 (N_5202,N_4878,N_5065);
nand U5203 (N_5203,N_5045,N_4986);
nand U5204 (N_5204,N_4973,N_4945);
nor U5205 (N_5205,N_4944,N_4839);
and U5206 (N_5206,N_5023,N_5024);
or U5207 (N_5207,N_5064,N_4803);
xor U5208 (N_5208,N_4913,N_5136);
and U5209 (N_5209,N_5121,N_4958);
and U5210 (N_5210,N_5173,N_5193);
and U5211 (N_5211,N_4881,N_4863);
or U5212 (N_5212,N_4963,N_4883);
and U5213 (N_5213,N_4821,N_4954);
xnor U5214 (N_5214,N_5016,N_4903);
nor U5215 (N_5215,N_4998,N_4802);
and U5216 (N_5216,N_4955,N_5127);
or U5217 (N_5217,N_5048,N_4801);
nand U5218 (N_5218,N_4942,N_5177);
xnor U5219 (N_5219,N_5165,N_4933);
or U5220 (N_5220,N_5194,N_5109);
xnor U5221 (N_5221,N_5091,N_5036);
nand U5222 (N_5222,N_4897,N_4912);
nor U5223 (N_5223,N_5152,N_5139);
or U5224 (N_5224,N_4867,N_4800);
or U5225 (N_5225,N_4895,N_5178);
and U5226 (N_5226,N_4979,N_5015);
nor U5227 (N_5227,N_4815,N_5179);
xnor U5228 (N_5228,N_5108,N_4814);
xor U5229 (N_5229,N_4907,N_5143);
nor U5230 (N_5230,N_4843,N_4980);
xnor U5231 (N_5231,N_4823,N_5039);
xor U5232 (N_5232,N_4994,N_4834);
or U5233 (N_5233,N_5078,N_4949);
nand U5234 (N_5234,N_5050,N_4857);
nand U5235 (N_5235,N_4808,N_4953);
nor U5236 (N_5236,N_5086,N_5115);
nor U5237 (N_5237,N_4888,N_5058);
or U5238 (N_5238,N_4886,N_5103);
nand U5239 (N_5239,N_5020,N_5159);
or U5240 (N_5240,N_4899,N_4946);
nand U5241 (N_5241,N_5180,N_5038);
nor U5242 (N_5242,N_4941,N_5129);
nand U5243 (N_5243,N_5160,N_4995);
nand U5244 (N_5244,N_4860,N_5014);
nor U5245 (N_5245,N_5126,N_5144);
nor U5246 (N_5246,N_4844,N_5049);
xor U5247 (N_5247,N_5120,N_4951);
xnor U5248 (N_5248,N_5057,N_4876);
nand U5249 (N_5249,N_4935,N_4922);
and U5250 (N_5250,N_4837,N_4835);
nand U5251 (N_5251,N_5138,N_4943);
and U5252 (N_5252,N_4921,N_4969);
nor U5253 (N_5253,N_5034,N_5080);
and U5254 (N_5254,N_4905,N_5021);
nor U5255 (N_5255,N_4915,N_4950);
and U5256 (N_5256,N_5124,N_4931);
xor U5257 (N_5257,N_4926,N_5122);
nor U5258 (N_5258,N_4990,N_4822);
nor U5259 (N_5259,N_4929,N_5140);
xnor U5260 (N_5260,N_4819,N_4978);
nand U5261 (N_5261,N_5006,N_5189);
nand U5262 (N_5262,N_4902,N_4810);
nand U5263 (N_5263,N_5102,N_5009);
nor U5264 (N_5264,N_4987,N_4811);
and U5265 (N_5265,N_4974,N_4812);
xnor U5266 (N_5266,N_5040,N_5069);
or U5267 (N_5267,N_5118,N_5134);
nand U5268 (N_5268,N_5051,N_4882);
nor U5269 (N_5269,N_4893,N_4825);
xnor U5270 (N_5270,N_5031,N_5079);
xnor U5271 (N_5271,N_5155,N_4924);
nand U5272 (N_5272,N_5005,N_4846);
nand U5273 (N_5273,N_5030,N_5043);
and U5274 (N_5274,N_4999,N_4804);
nand U5275 (N_5275,N_5183,N_4900);
and U5276 (N_5276,N_5184,N_4865);
and U5277 (N_5277,N_5104,N_5157);
nor U5278 (N_5278,N_5167,N_5135);
or U5279 (N_5279,N_5137,N_4925);
nand U5280 (N_5280,N_5084,N_5077);
nor U5281 (N_5281,N_5114,N_5082);
nand U5282 (N_5282,N_5085,N_4866);
or U5283 (N_5283,N_5192,N_5092);
or U5284 (N_5284,N_5187,N_4845);
or U5285 (N_5285,N_5076,N_5029);
xor U5286 (N_5286,N_4809,N_5170);
nor U5287 (N_5287,N_4909,N_4805);
and U5288 (N_5288,N_5149,N_4827);
nand U5289 (N_5289,N_4849,N_5055);
nor U5290 (N_5290,N_4920,N_5164);
xor U5291 (N_5291,N_4864,N_4874);
xnor U5292 (N_5292,N_4828,N_5075);
nor U5293 (N_5293,N_5105,N_4989);
nor U5294 (N_5294,N_5188,N_4936);
xor U5295 (N_5295,N_5003,N_5071);
nor U5296 (N_5296,N_5095,N_5096);
or U5297 (N_5297,N_4964,N_4960);
nor U5298 (N_5298,N_5141,N_5146);
nand U5299 (N_5299,N_5035,N_5081);
and U5300 (N_5300,N_4873,N_5119);
nor U5301 (N_5301,N_5161,N_5190);
or U5302 (N_5302,N_5197,N_4813);
nor U5303 (N_5303,N_4908,N_4879);
nor U5304 (N_5304,N_5088,N_4894);
or U5305 (N_5305,N_5151,N_5002);
and U5306 (N_5306,N_5195,N_4996);
nor U5307 (N_5307,N_5169,N_5072);
and U5308 (N_5308,N_5060,N_5117);
and U5309 (N_5309,N_4967,N_5001);
or U5310 (N_5310,N_4901,N_4847);
nor U5311 (N_5311,N_4852,N_4887);
nor U5312 (N_5312,N_5054,N_4896);
xnor U5313 (N_5313,N_5008,N_4928);
and U5314 (N_5314,N_4972,N_4914);
nand U5315 (N_5315,N_5162,N_5019);
and U5316 (N_5316,N_4861,N_4890);
and U5317 (N_5317,N_4991,N_5130);
or U5318 (N_5318,N_5099,N_4956);
or U5319 (N_5319,N_5196,N_4842);
nand U5320 (N_5320,N_4836,N_4853);
and U5321 (N_5321,N_5176,N_4970);
nor U5322 (N_5322,N_4976,N_4993);
nor U5323 (N_5323,N_4971,N_4820);
or U5324 (N_5324,N_4961,N_5100);
xor U5325 (N_5325,N_5111,N_4947);
nor U5326 (N_5326,N_5110,N_4871);
nor U5327 (N_5327,N_5112,N_5094);
xor U5328 (N_5328,N_5182,N_5017);
xor U5329 (N_5329,N_5063,N_4984);
nor U5330 (N_5330,N_5090,N_4807);
xnor U5331 (N_5331,N_4982,N_5172);
nor U5332 (N_5332,N_4851,N_5000);
and U5333 (N_5333,N_5107,N_4959);
nand U5334 (N_5334,N_5007,N_5083);
nand U5335 (N_5335,N_4848,N_4877);
xor U5336 (N_5336,N_4997,N_5133);
or U5337 (N_5337,N_5010,N_4981);
nor U5338 (N_5338,N_5101,N_5047);
nand U5339 (N_5339,N_4833,N_4930);
nor U5340 (N_5340,N_5061,N_5056);
nor U5341 (N_5341,N_4831,N_5046);
and U5342 (N_5342,N_4816,N_4911);
xor U5343 (N_5343,N_4832,N_4937);
nand U5344 (N_5344,N_5145,N_4917);
nand U5345 (N_5345,N_5116,N_5154);
xor U5346 (N_5346,N_5106,N_5153);
and U5347 (N_5347,N_5018,N_5168);
or U5348 (N_5348,N_4906,N_4932);
nor U5349 (N_5349,N_4884,N_5181);
and U5350 (N_5350,N_4966,N_4919);
nor U5351 (N_5351,N_5191,N_5053);
nand U5352 (N_5352,N_5186,N_4855);
or U5353 (N_5353,N_4988,N_5026);
nand U5354 (N_5354,N_5132,N_4918);
or U5355 (N_5355,N_5059,N_5166);
xnor U5356 (N_5356,N_5087,N_5013);
or U5357 (N_5357,N_4939,N_4858);
or U5358 (N_5358,N_5022,N_5074);
or U5359 (N_5359,N_5011,N_5163);
nand U5360 (N_5360,N_5070,N_4885);
nand U5361 (N_5361,N_5052,N_4806);
nor U5362 (N_5362,N_5148,N_4904);
nand U5363 (N_5363,N_4948,N_5185);
nand U5364 (N_5364,N_4870,N_4898);
xnor U5365 (N_5365,N_5171,N_4891);
xnor U5366 (N_5366,N_5073,N_5033);
xnor U5367 (N_5367,N_4940,N_5093);
xor U5368 (N_5368,N_5044,N_4826);
xnor U5369 (N_5369,N_5175,N_5012);
xor U5370 (N_5370,N_4952,N_4985);
and U5371 (N_5371,N_4838,N_5027);
nand U5372 (N_5372,N_4818,N_5068);
nand U5373 (N_5373,N_4934,N_4892);
nand U5374 (N_5374,N_4862,N_4859);
and U5375 (N_5375,N_5131,N_4830);
xor U5376 (N_5376,N_5125,N_5042);
xor U5377 (N_5377,N_4975,N_5025);
xnor U5378 (N_5378,N_5089,N_4824);
nor U5379 (N_5379,N_5062,N_4916);
xnor U5380 (N_5380,N_4817,N_4880);
nand U5381 (N_5381,N_4965,N_5123);
nand U5382 (N_5382,N_5041,N_5098);
and U5383 (N_5383,N_5199,N_4856);
or U5384 (N_5384,N_4910,N_4840);
or U5385 (N_5385,N_5004,N_5147);
xnor U5386 (N_5386,N_4889,N_4977);
nand U5387 (N_5387,N_4854,N_4829);
nand U5388 (N_5388,N_4968,N_4957);
or U5389 (N_5389,N_5150,N_5067);
and U5390 (N_5390,N_4841,N_4872);
xnor U5391 (N_5391,N_4850,N_5174);
nor U5392 (N_5392,N_5066,N_5028);
nor U5393 (N_5393,N_4983,N_5037);
xnor U5394 (N_5394,N_4962,N_5097);
or U5395 (N_5395,N_4938,N_4868);
nor U5396 (N_5396,N_4992,N_4927);
nand U5397 (N_5397,N_5142,N_5032);
or U5398 (N_5398,N_5158,N_5156);
or U5399 (N_5399,N_5128,N_4875);
or U5400 (N_5400,N_5027,N_5028);
or U5401 (N_5401,N_4880,N_5163);
or U5402 (N_5402,N_5125,N_4856);
or U5403 (N_5403,N_5114,N_4813);
and U5404 (N_5404,N_4878,N_5051);
nor U5405 (N_5405,N_4867,N_4871);
and U5406 (N_5406,N_5098,N_4846);
or U5407 (N_5407,N_4856,N_4930);
nor U5408 (N_5408,N_5060,N_4840);
or U5409 (N_5409,N_4964,N_4880);
or U5410 (N_5410,N_5027,N_5147);
or U5411 (N_5411,N_4953,N_5039);
nor U5412 (N_5412,N_4868,N_5180);
or U5413 (N_5413,N_4868,N_5079);
and U5414 (N_5414,N_5004,N_4820);
or U5415 (N_5415,N_5002,N_5192);
nand U5416 (N_5416,N_4966,N_5016);
or U5417 (N_5417,N_4966,N_4892);
or U5418 (N_5418,N_5189,N_5180);
or U5419 (N_5419,N_5043,N_4970);
and U5420 (N_5420,N_5137,N_4834);
and U5421 (N_5421,N_4877,N_5127);
xnor U5422 (N_5422,N_4920,N_4938);
nor U5423 (N_5423,N_5039,N_4848);
and U5424 (N_5424,N_4813,N_4826);
or U5425 (N_5425,N_4950,N_4905);
nand U5426 (N_5426,N_4932,N_4852);
or U5427 (N_5427,N_4821,N_5045);
xnor U5428 (N_5428,N_4899,N_4920);
nand U5429 (N_5429,N_5194,N_4995);
xor U5430 (N_5430,N_4822,N_4853);
nand U5431 (N_5431,N_5060,N_5155);
xor U5432 (N_5432,N_5086,N_4918);
or U5433 (N_5433,N_5166,N_4993);
nand U5434 (N_5434,N_4828,N_5004);
nand U5435 (N_5435,N_5114,N_5167);
nor U5436 (N_5436,N_4806,N_4906);
and U5437 (N_5437,N_4878,N_4979);
nand U5438 (N_5438,N_4937,N_4996);
nand U5439 (N_5439,N_4930,N_4837);
or U5440 (N_5440,N_4946,N_5024);
xnor U5441 (N_5441,N_5016,N_4958);
xor U5442 (N_5442,N_5190,N_5052);
or U5443 (N_5443,N_5141,N_4996);
or U5444 (N_5444,N_4982,N_5004);
and U5445 (N_5445,N_5163,N_4996);
or U5446 (N_5446,N_4925,N_4982);
nand U5447 (N_5447,N_4972,N_5050);
nand U5448 (N_5448,N_4965,N_4860);
or U5449 (N_5449,N_4906,N_4955);
xnor U5450 (N_5450,N_4906,N_5095);
nand U5451 (N_5451,N_4821,N_5175);
and U5452 (N_5452,N_5077,N_4880);
nor U5453 (N_5453,N_5179,N_4889);
xor U5454 (N_5454,N_4805,N_5123);
nand U5455 (N_5455,N_5113,N_5165);
and U5456 (N_5456,N_4998,N_5065);
xor U5457 (N_5457,N_4848,N_5163);
nand U5458 (N_5458,N_4864,N_5095);
and U5459 (N_5459,N_5073,N_4875);
and U5460 (N_5460,N_5069,N_5169);
nand U5461 (N_5461,N_5111,N_5016);
or U5462 (N_5462,N_5100,N_5120);
xor U5463 (N_5463,N_4874,N_5166);
xnor U5464 (N_5464,N_5176,N_5041);
xnor U5465 (N_5465,N_4981,N_4837);
nor U5466 (N_5466,N_4840,N_5103);
nand U5467 (N_5467,N_4833,N_5151);
and U5468 (N_5468,N_5145,N_5122);
xor U5469 (N_5469,N_4847,N_5133);
nand U5470 (N_5470,N_5034,N_5031);
and U5471 (N_5471,N_5181,N_4900);
and U5472 (N_5472,N_4979,N_5125);
xnor U5473 (N_5473,N_4942,N_5117);
or U5474 (N_5474,N_4930,N_5184);
xnor U5475 (N_5475,N_5114,N_5078);
or U5476 (N_5476,N_4819,N_4810);
or U5477 (N_5477,N_5089,N_5005);
nor U5478 (N_5478,N_5066,N_4962);
or U5479 (N_5479,N_4832,N_5147);
xnor U5480 (N_5480,N_5020,N_4854);
xnor U5481 (N_5481,N_5165,N_4846);
xnor U5482 (N_5482,N_4898,N_4892);
xnor U5483 (N_5483,N_4857,N_5059);
nand U5484 (N_5484,N_4810,N_4907);
or U5485 (N_5485,N_5051,N_4922);
xnor U5486 (N_5486,N_4907,N_5171);
xor U5487 (N_5487,N_5082,N_4857);
nand U5488 (N_5488,N_5085,N_5157);
nand U5489 (N_5489,N_5187,N_4902);
nand U5490 (N_5490,N_4866,N_5194);
and U5491 (N_5491,N_4938,N_5011);
or U5492 (N_5492,N_4905,N_4877);
nor U5493 (N_5493,N_4802,N_4869);
or U5494 (N_5494,N_4898,N_4927);
xor U5495 (N_5495,N_4831,N_4948);
nor U5496 (N_5496,N_5068,N_5135);
or U5497 (N_5497,N_5017,N_5183);
xnor U5498 (N_5498,N_4879,N_5141);
xnor U5499 (N_5499,N_4953,N_4850);
nand U5500 (N_5500,N_4857,N_5034);
nor U5501 (N_5501,N_4852,N_4938);
xnor U5502 (N_5502,N_5132,N_5042);
and U5503 (N_5503,N_5115,N_4915);
xnor U5504 (N_5504,N_4849,N_4886);
and U5505 (N_5505,N_5128,N_4983);
xor U5506 (N_5506,N_4860,N_5156);
nand U5507 (N_5507,N_5049,N_4921);
nand U5508 (N_5508,N_4901,N_5001);
xnor U5509 (N_5509,N_4988,N_5073);
nand U5510 (N_5510,N_4914,N_5033);
or U5511 (N_5511,N_5135,N_4882);
nand U5512 (N_5512,N_5135,N_4961);
nand U5513 (N_5513,N_4942,N_5154);
xnor U5514 (N_5514,N_4951,N_5137);
nand U5515 (N_5515,N_4929,N_4945);
nand U5516 (N_5516,N_5177,N_4921);
nor U5517 (N_5517,N_4932,N_5134);
or U5518 (N_5518,N_5123,N_5125);
and U5519 (N_5519,N_5158,N_4942);
nand U5520 (N_5520,N_5178,N_4878);
nand U5521 (N_5521,N_5156,N_5074);
nand U5522 (N_5522,N_4876,N_4815);
xnor U5523 (N_5523,N_5041,N_5013);
xnor U5524 (N_5524,N_4874,N_5122);
and U5525 (N_5525,N_4834,N_4801);
nor U5526 (N_5526,N_5094,N_4839);
and U5527 (N_5527,N_4889,N_4873);
nor U5528 (N_5528,N_5152,N_4987);
xnor U5529 (N_5529,N_5012,N_5084);
nor U5530 (N_5530,N_5174,N_4861);
xor U5531 (N_5531,N_4878,N_4835);
and U5532 (N_5532,N_4929,N_4907);
xor U5533 (N_5533,N_4877,N_4852);
xor U5534 (N_5534,N_5116,N_5120);
or U5535 (N_5535,N_4977,N_4892);
xnor U5536 (N_5536,N_4816,N_4991);
and U5537 (N_5537,N_5117,N_5126);
or U5538 (N_5538,N_5039,N_5149);
and U5539 (N_5539,N_5062,N_5146);
and U5540 (N_5540,N_5146,N_5152);
and U5541 (N_5541,N_5133,N_5188);
and U5542 (N_5542,N_5112,N_4913);
and U5543 (N_5543,N_5185,N_5035);
xor U5544 (N_5544,N_5183,N_5165);
xnor U5545 (N_5545,N_4909,N_4994);
and U5546 (N_5546,N_4875,N_4996);
or U5547 (N_5547,N_5084,N_5093);
or U5548 (N_5548,N_4867,N_4933);
or U5549 (N_5549,N_4963,N_5170);
nand U5550 (N_5550,N_5142,N_4919);
nand U5551 (N_5551,N_4863,N_5145);
nor U5552 (N_5552,N_4954,N_5158);
nand U5553 (N_5553,N_4967,N_5167);
and U5554 (N_5554,N_5139,N_4912);
and U5555 (N_5555,N_4806,N_4869);
and U5556 (N_5556,N_5036,N_5188);
nand U5557 (N_5557,N_4933,N_5193);
and U5558 (N_5558,N_5147,N_4915);
nor U5559 (N_5559,N_5010,N_4912);
xor U5560 (N_5560,N_4883,N_5174);
nand U5561 (N_5561,N_4884,N_4978);
xor U5562 (N_5562,N_5194,N_4996);
or U5563 (N_5563,N_4952,N_4920);
nand U5564 (N_5564,N_5194,N_4914);
nand U5565 (N_5565,N_5138,N_4864);
nor U5566 (N_5566,N_4882,N_4820);
or U5567 (N_5567,N_5193,N_5177);
and U5568 (N_5568,N_4837,N_4917);
nor U5569 (N_5569,N_4987,N_5188);
or U5570 (N_5570,N_4981,N_4810);
xnor U5571 (N_5571,N_4863,N_5118);
and U5572 (N_5572,N_4865,N_4805);
nor U5573 (N_5573,N_4840,N_5004);
xnor U5574 (N_5574,N_5091,N_5092);
nor U5575 (N_5575,N_4860,N_5170);
and U5576 (N_5576,N_5004,N_4941);
or U5577 (N_5577,N_4899,N_5176);
nand U5578 (N_5578,N_4949,N_5031);
xnor U5579 (N_5579,N_4844,N_4917);
xor U5580 (N_5580,N_5044,N_4858);
xor U5581 (N_5581,N_4954,N_5022);
or U5582 (N_5582,N_5151,N_4928);
nand U5583 (N_5583,N_4871,N_4899);
xnor U5584 (N_5584,N_5165,N_5091);
nand U5585 (N_5585,N_5018,N_5166);
nand U5586 (N_5586,N_4887,N_5039);
nand U5587 (N_5587,N_4915,N_4826);
nand U5588 (N_5588,N_5129,N_4943);
or U5589 (N_5589,N_4816,N_5086);
xor U5590 (N_5590,N_5108,N_5095);
nand U5591 (N_5591,N_5012,N_4866);
xnor U5592 (N_5592,N_5166,N_4915);
and U5593 (N_5593,N_4958,N_4942);
or U5594 (N_5594,N_4921,N_5025);
xor U5595 (N_5595,N_4990,N_5068);
nand U5596 (N_5596,N_5058,N_4835);
nand U5597 (N_5597,N_5050,N_5154);
xor U5598 (N_5598,N_4931,N_4949);
and U5599 (N_5599,N_4919,N_5131);
xnor U5600 (N_5600,N_5576,N_5565);
nand U5601 (N_5601,N_5235,N_5424);
nand U5602 (N_5602,N_5457,N_5237);
xnor U5603 (N_5603,N_5242,N_5384);
nor U5604 (N_5604,N_5543,N_5439);
or U5605 (N_5605,N_5426,N_5532);
nand U5606 (N_5606,N_5541,N_5560);
nand U5607 (N_5607,N_5420,N_5452);
nor U5608 (N_5608,N_5526,N_5524);
and U5609 (N_5609,N_5364,N_5536);
xor U5610 (N_5610,N_5370,N_5594);
and U5611 (N_5611,N_5510,N_5398);
nor U5612 (N_5612,N_5337,N_5278);
xor U5613 (N_5613,N_5486,N_5280);
nand U5614 (N_5614,N_5395,N_5417);
xor U5615 (N_5615,N_5512,N_5517);
and U5616 (N_5616,N_5302,N_5238);
or U5617 (N_5617,N_5497,N_5410);
nor U5618 (N_5618,N_5401,N_5249);
xnor U5619 (N_5619,N_5202,N_5305);
xnor U5620 (N_5620,N_5312,N_5492);
or U5621 (N_5621,N_5411,N_5393);
and U5622 (N_5622,N_5349,N_5493);
or U5623 (N_5623,N_5385,N_5256);
nor U5624 (N_5624,N_5529,N_5422);
and U5625 (N_5625,N_5366,N_5599);
nand U5626 (N_5626,N_5458,N_5483);
nor U5627 (N_5627,N_5352,N_5453);
nor U5628 (N_5628,N_5261,N_5380);
or U5629 (N_5629,N_5511,N_5584);
xnor U5630 (N_5630,N_5583,N_5437);
nor U5631 (N_5631,N_5563,N_5266);
or U5632 (N_5632,N_5234,N_5327);
nor U5633 (N_5633,N_5525,N_5389);
xnor U5634 (N_5634,N_5315,N_5468);
or U5635 (N_5635,N_5431,N_5329);
nand U5636 (N_5636,N_5471,N_5296);
or U5637 (N_5637,N_5204,N_5416);
nand U5638 (N_5638,N_5503,N_5341);
nor U5639 (N_5639,N_5523,N_5519);
or U5640 (N_5640,N_5274,N_5252);
nor U5641 (N_5641,N_5430,N_5592);
nor U5642 (N_5642,N_5507,N_5250);
and U5643 (N_5643,N_5570,N_5295);
xnor U5644 (N_5644,N_5338,N_5396);
and U5645 (N_5645,N_5284,N_5449);
xnor U5646 (N_5646,N_5262,N_5243);
or U5647 (N_5647,N_5432,N_5596);
xnor U5648 (N_5648,N_5546,N_5551);
nand U5649 (N_5649,N_5224,N_5264);
and U5650 (N_5650,N_5346,N_5566);
nor U5651 (N_5651,N_5530,N_5419);
nand U5652 (N_5652,N_5595,N_5253);
nand U5653 (N_5653,N_5292,N_5217);
or U5654 (N_5654,N_5372,N_5404);
or U5655 (N_5655,N_5323,N_5581);
or U5656 (N_5656,N_5528,N_5455);
and U5657 (N_5657,N_5265,N_5228);
nor U5658 (N_5658,N_5454,N_5520);
or U5659 (N_5659,N_5226,N_5379);
or U5660 (N_5660,N_5571,N_5498);
nor U5661 (N_5661,N_5374,N_5462);
nand U5662 (N_5662,N_5300,N_5553);
or U5663 (N_5663,N_5209,N_5218);
xor U5664 (N_5664,N_5445,N_5232);
and U5665 (N_5665,N_5347,N_5239);
nor U5666 (N_5666,N_5531,N_5298);
nand U5667 (N_5667,N_5499,N_5459);
and U5668 (N_5668,N_5527,N_5506);
or U5669 (N_5669,N_5255,N_5388);
nand U5670 (N_5670,N_5474,N_5588);
xnor U5671 (N_5671,N_5465,N_5200);
xnor U5672 (N_5672,N_5476,N_5310);
nand U5673 (N_5673,N_5211,N_5326);
xor U5674 (N_5674,N_5275,N_5277);
xnor U5675 (N_5675,N_5537,N_5350);
nor U5676 (N_5676,N_5436,N_5362);
nor U5677 (N_5677,N_5263,N_5518);
nand U5678 (N_5678,N_5301,N_5285);
nor U5679 (N_5679,N_5375,N_5590);
nand U5680 (N_5680,N_5438,N_5478);
and U5681 (N_5681,N_5267,N_5308);
nand U5682 (N_5682,N_5258,N_5355);
nor U5683 (N_5683,N_5585,N_5221);
and U5684 (N_5684,N_5552,N_5399);
nand U5685 (N_5685,N_5522,N_5429);
nand U5686 (N_5686,N_5297,N_5535);
nor U5687 (N_5687,N_5466,N_5593);
or U5688 (N_5688,N_5539,N_5540);
xnor U5689 (N_5689,N_5282,N_5409);
or U5690 (N_5690,N_5397,N_5490);
nor U5691 (N_5691,N_5472,N_5387);
nor U5692 (N_5692,N_5214,N_5494);
or U5693 (N_5693,N_5351,N_5544);
or U5694 (N_5694,N_5365,N_5291);
or U5695 (N_5695,N_5545,N_5220);
nor U5696 (N_5696,N_5271,N_5331);
and U5697 (N_5697,N_5574,N_5319);
xnor U5698 (N_5698,N_5394,N_5367);
nand U5699 (N_5699,N_5236,N_5230);
nand U5700 (N_5700,N_5477,N_5550);
nor U5701 (N_5701,N_5373,N_5270);
nor U5702 (N_5702,N_5360,N_5555);
nand U5703 (N_5703,N_5304,N_5371);
nor U5704 (N_5704,N_5359,N_5335);
and U5705 (N_5705,N_5533,N_5484);
nand U5706 (N_5706,N_5311,N_5402);
and U5707 (N_5707,N_5582,N_5336);
nor U5708 (N_5708,N_5299,N_5421);
or U5709 (N_5709,N_5475,N_5223);
nand U5710 (N_5710,N_5377,N_5485);
and U5711 (N_5711,N_5245,N_5279);
xnor U5712 (N_5712,N_5248,N_5491);
nor U5713 (N_5713,N_5502,N_5244);
nand U5714 (N_5714,N_5440,N_5521);
nand U5715 (N_5715,N_5559,N_5568);
or U5716 (N_5716,N_5227,N_5461);
or U5717 (N_5717,N_5504,N_5333);
and U5718 (N_5718,N_5446,N_5213);
or U5719 (N_5719,N_5460,N_5339);
nand U5720 (N_5720,N_5408,N_5210);
or U5721 (N_5721,N_5231,N_5442);
xnor U5722 (N_5722,N_5547,N_5317);
xor U5723 (N_5723,N_5342,N_5293);
and U5724 (N_5724,N_5233,N_5260);
nor U5725 (N_5725,N_5240,N_5448);
nand U5726 (N_5726,N_5515,N_5434);
or U5727 (N_5727,N_5463,N_5324);
or U5728 (N_5728,N_5586,N_5273);
nor U5729 (N_5729,N_5573,N_5225);
or U5730 (N_5730,N_5307,N_5325);
or U5731 (N_5731,N_5363,N_5215);
or U5732 (N_5732,N_5514,N_5314);
xnor U5733 (N_5733,N_5435,N_5320);
nand U5734 (N_5734,N_5356,N_5358);
and U5735 (N_5735,N_5340,N_5201);
nand U5736 (N_5736,N_5470,N_5309);
and U5737 (N_5737,N_5538,N_5428);
nor U5738 (N_5738,N_5212,N_5423);
nor U5739 (N_5739,N_5257,N_5332);
nand U5740 (N_5740,N_5381,N_5208);
nand U5741 (N_5741,N_5246,N_5287);
nand U5742 (N_5742,N_5508,N_5316);
nand U5743 (N_5743,N_5286,N_5534);
xnor U5744 (N_5744,N_5561,N_5578);
xor U5745 (N_5745,N_5587,N_5572);
xnor U5746 (N_5746,N_5569,N_5501);
and U5747 (N_5747,N_5254,N_5405);
nand U5748 (N_5748,N_5318,N_5294);
or U5749 (N_5749,N_5283,N_5591);
and U5750 (N_5750,N_5353,N_5496);
nor U5751 (N_5751,N_5361,N_5412);
or U5752 (N_5752,N_5383,N_5216);
nor U5753 (N_5753,N_5345,N_5334);
nand U5754 (N_5754,N_5473,N_5391);
xor U5755 (N_5755,N_5597,N_5589);
nand U5756 (N_5756,N_5480,N_5281);
and U5757 (N_5757,N_5328,N_5427);
nand U5758 (N_5758,N_5450,N_5382);
or U5759 (N_5759,N_5418,N_5269);
or U5760 (N_5760,N_5577,N_5203);
and U5761 (N_5761,N_5415,N_5441);
or U5762 (N_5762,N_5500,N_5481);
xor U5763 (N_5763,N_5313,N_5272);
nand U5764 (N_5764,N_5376,N_5580);
and U5765 (N_5765,N_5425,N_5549);
and U5766 (N_5766,N_5557,N_5344);
xnor U5767 (N_5767,N_5343,N_5456);
or U5768 (N_5768,N_5489,N_5403);
or U5769 (N_5769,N_5505,N_5241);
or U5770 (N_5770,N_5447,N_5479);
nand U5771 (N_5771,N_5564,N_5369);
or U5772 (N_5772,N_5205,N_5259);
and U5773 (N_5773,N_5368,N_5414);
nor U5774 (N_5774,N_5251,N_5321);
nor U5775 (N_5775,N_5206,N_5451);
nor U5776 (N_5776,N_5464,N_5219);
or U5777 (N_5777,N_5378,N_5390);
nand U5778 (N_5778,N_5407,N_5598);
xnor U5779 (N_5779,N_5579,N_5433);
or U5780 (N_5780,N_5354,N_5567);
or U5781 (N_5781,N_5229,N_5276);
nor U5782 (N_5782,N_5207,N_5556);
or U5783 (N_5783,N_5495,N_5268);
nor U5784 (N_5784,N_5575,N_5290);
or U5785 (N_5785,N_5558,N_5322);
nand U5786 (N_5786,N_5444,N_5406);
and U5787 (N_5787,N_5357,N_5487);
nand U5788 (N_5788,N_5222,N_5289);
and U5789 (N_5789,N_5413,N_5288);
nand U5790 (N_5790,N_5348,N_5554);
or U5791 (N_5791,N_5247,N_5392);
nand U5792 (N_5792,N_5303,N_5513);
xnor U5793 (N_5793,N_5562,N_5516);
or U5794 (N_5794,N_5548,N_5400);
or U5795 (N_5795,N_5386,N_5542);
nand U5796 (N_5796,N_5482,N_5330);
and U5797 (N_5797,N_5467,N_5469);
nand U5798 (N_5798,N_5488,N_5306);
xnor U5799 (N_5799,N_5509,N_5443);
or U5800 (N_5800,N_5475,N_5538);
nand U5801 (N_5801,N_5528,N_5276);
nand U5802 (N_5802,N_5499,N_5447);
or U5803 (N_5803,N_5577,N_5297);
nand U5804 (N_5804,N_5314,N_5379);
or U5805 (N_5805,N_5377,N_5267);
nor U5806 (N_5806,N_5375,N_5450);
nand U5807 (N_5807,N_5457,N_5363);
and U5808 (N_5808,N_5229,N_5523);
or U5809 (N_5809,N_5516,N_5445);
and U5810 (N_5810,N_5300,N_5560);
or U5811 (N_5811,N_5380,N_5228);
and U5812 (N_5812,N_5466,N_5486);
and U5813 (N_5813,N_5345,N_5501);
nor U5814 (N_5814,N_5569,N_5258);
xor U5815 (N_5815,N_5267,N_5369);
or U5816 (N_5816,N_5575,N_5499);
nand U5817 (N_5817,N_5259,N_5408);
nor U5818 (N_5818,N_5290,N_5511);
xor U5819 (N_5819,N_5217,N_5280);
and U5820 (N_5820,N_5490,N_5576);
and U5821 (N_5821,N_5523,N_5535);
nor U5822 (N_5822,N_5399,N_5400);
xor U5823 (N_5823,N_5350,N_5561);
xor U5824 (N_5824,N_5570,N_5437);
xnor U5825 (N_5825,N_5588,N_5525);
xnor U5826 (N_5826,N_5307,N_5300);
nor U5827 (N_5827,N_5232,N_5204);
and U5828 (N_5828,N_5237,N_5530);
or U5829 (N_5829,N_5571,N_5457);
or U5830 (N_5830,N_5558,N_5218);
nand U5831 (N_5831,N_5388,N_5398);
xnor U5832 (N_5832,N_5544,N_5337);
nand U5833 (N_5833,N_5283,N_5580);
xnor U5834 (N_5834,N_5462,N_5450);
or U5835 (N_5835,N_5336,N_5300);
xnor U5836 (N_5836,N_5528,N_5274);
nor U5837 (N_5837,N_5382,N_5538);
or U5838 (N_5838,N_5239,N_5467);
nand U5839 (N_5839,N_5328,N_5593);
xnor U5840 (N_5840,N_5244,N_5326);
nand U5841 (N_5841,N_5456,N_5235);
nand U5842 (N_5842,N_5433,N_5253);
nor U5843 (N_5843,N_5272,N_5559);
or U5844 (N_5844,N_5459,N_5224);
xor U5845 (N_5845,N_5366,N_5328);
nor U5846 (N_5846,N_5270,N_5335);
or U5847 (N_5847,N_5496,N_5432);
and U5848 (N_5848,N_5406,N_5276);
xnor U5849 (N_5849,N_5353,N_5204);
xnor U5850 (N_5850,N_5331,N_5318);
xor U5851 (N_5851,N_5457,N_5250);
and U5852 (N_5852,N_5331,N_5463);
and U5853 (N_5853,N_5475,N_5590);
or U5854 (N_5854,N_5569,N_5272);
nor U5855 (N_5855,N_5341,N_5336);
nor U5856 (N_5856,N_5419,N_5200);
xor U5857 (N_5857,N_5355,N_5392);
xnor U5858 (N_5858,N_5252,N_5250);
nor U5859 (N_5859,N_5276,N_5562);
xnor U5860 (N_5860,N_5577,N_5236);
nand U5861 (N_5861,N_5540,N_5235);
or U5862 (N_5862,N_5563,N_5551);
xor U5863 (N_5863,N_5402,N_5493);
nor U5864 (N_5864,N_5318,N_5513);
xor U5865 (N_5865,N_5438,N_5264);
and U5866 (N_5866,N_5282,N_5239);
nand U5867 (N_5867,N_5383,N_5407);
nor U5868 (N_5868,N_5237,N_5560);
xor U5869 (N_5869,N_5257,N_5234);
and U5870 (N_5870,N_5230,N_5457);
or U5871 (N_5871,N_5592,N_5232);
xnor U5872 (N_5872,N_5222,N_5460);
nand U5873 (N_5873,N_5414,N_5302);
nand U5874 (N_5874,N_5485,N_5531);
nand U5875 (N_5875,N_5496,N_5395);
or U5876 (N_5876,N_5479,N_5358);
xnor U5877 (N_5877,N_5220,N_5494);
nand U5878 (N_5878,N_5467,N_5254);
xnor U5879 (N_5879,N_5302,N_5552);
or U5880 (N_5880,N_5460,N_5249);
nor U5881 (N_5881,N_5305,N_5432);
nand U5882 (N_5882,N_5346,N_5382);
nand U5883 (N_5883,N_5488,N_5356);
nand U5884 (N_5884,N_5501,N_5249);
or U5885 (N_5885,N_5274,N_5365);
xor U5886 (N_5886,N_5377,N_5341);
xnor U5887 (N_5887,N_5432,N_5371);
and U5888 (N_5888,N_5482,N_5557);
and U5889 (N_5889,N_5319,N_5313);
and U5890 (N_5890,N_5245,N_5388);
nand U5891 (N_5891,N_5260,N_5513);
xnor U5892 (N_5892,N_5581,N_5318);
xnor U5893 (N_5893,N_5519,N_5578);
or U5894 (N_5894,N_5508,N_5539);
and U5895 (N_5895,N_5566,N_5576);
nand U5896 (N_5896,N_5538,N_5328);
xor U5897 (N_5897,N_5255,N_5243);
nand U5898 (N_5898,N_5548,N_5422);
and U5899 (N_5899,N_5285,N_5247);
and U5900 (N_5900,N_5413,N_5395);
or U5901 (N_5901,N_5457,N_5516);
xnor U5902 (N_5902,N_5558,N_5317);
nor U5903 (N_5903,N_5487,N_5410);
nor U5904 (N_5904,N_5476,N_5528);
or U5905 (N_5905,N_5527,N_5554);
nor U5906 (N_5906,N_5303,N_5202);
nor U5907 (N_5907,N_5580,N_5294);
xnor U5908 (N_5908,N_5383,N_5302);
or U5909 (N_5909,N_5327,N_5475);
xnor U5910 (N_5910,N_5595,N_5568);
xor U5911 (N_5911,N_5370,N_5258);
nand U5912 (N_5912,N_5588,N_5244);
and U5913 (N_5913,N_5553,N_5314);
nand U5914 (N_5914,N_5567,N_5206);
and U5915 (N_5915,N_5446,N_5398);
nand U5916 (N_5916,N_5225,N_5339);
xor U5917 (N_5917,N_5348,N_5511);
xnor U5918 (N_5918,N_5523,N_5568);
and U5919 (N_5919,N_5296,N_5478);
and U5920 (N_5920,N_5334,N_5229);
and U5921 (N_5921,N_5466,N_5502);
and U5922 (N_5922,N_5414,N_5441);
and U5923 (N_5923,N_5574,N_5283);
nor U5924 (N_5924,N_5248,N_5305);
or U5925 (N_5925,N_5468,N_5414);
nor U5926 (N_5926,N_5201,N_5242);
nand U5927 (N_5927,N_5411,N_5499);
nor U5928 (N_5928,N_5514,N_5422);
xnor U5929 (N_5929,N_5525,N_5386);
xnor U5930 (N_5930,N_5489,N_5370);
nand U5931 (N_5931,N_5555,N_5206);
nor U5932 (N_5932,N_5361,N_5505);
xor U5933 (N_5933,N_5305,N_5587);
xnor U5934 (N_5934,N_5431,N_5412);
xor U5935 (N_5935,N_5438,N_5417);
nor U5936 (N_5936,N_5256,N_5327);
nor U5937 (N_5937,N_5565,N_5389);
and U5938 (N_5938,N_5573,N_5296);
or U5939 (N_5939,N_5521,N_5361);
nand U5940 (N_5940,N_5496,N_5412);
and U5941 (N_5941,N_5444,N_5358);
xor U5942 (N_5942,N_5388,N_5396);
and U5943 (N_5943,N_5278,N_5438);
or U5944 (N_5944,N_5245,N_5260);
xor U5945 (N_5945,N_5357,N_5222);
or U5946 (N_5946,N_5512,N_5583);
nor U5947 (N_5947,N_5473,N_5479);
xor U5948 (N_5948,N_5586,N_5361);
nand U5949 (N_5949,N_5228,N_5406);
nor U5950 (N_5950,N_5320,N_5234);
nor U5951 (N_5951,N_5210,N_5207);
or U5952 (N_5952,N_5438,N_5539);
nand U5953 (N_5953,N_5245,N_5263);
nand U5954 (N_5954,N_5425,N_5330);
nand U5955 (N_5955,N_5466,N_5330);
and U5956 (N_5956,N_5512,N_5540);
or U5957 (N_5957,N_5591,N_5370);
nand U5958 (N_5958,N_5563,N_5376);
xor U5959 (N_5959,N_5419,N_5389);
or U5960 (N_5960,N_5403,N_5513);
nor U5961 (N_5961,N_5237,N_5517);
and U5962 (N_5962,N_5292,N_5455);
xnor U5963 (N_5963,N_5351,N_5529);
xnor U5964 (N_5964,N_5599,N_5530);
nand U5965 (N_5965,N_5303,N_5593);
nor U5966 (N_5966,N_5519,N_5288);
or U5967 (N_5967,N_5490,N_5258);
or U5968 (N_5968,N_5204,N_5312);
and U5969 (N_5969,N_5207,N_5254);
nor U5970 (N_5970,N_5366,N_5338);
nand U5971 (N_5971,N_5443,N_5525);
nor U5972 (N_5972,N_5420,N_5213);
or U5973 (N_5973,N_5402,N_5542);
or U5974 (N_5974,N_5227,N_5575);
nand U5975 (N_5975,N_5577,N_5531);
nand U5976 (N_5976,N_5287,N_5587);
xor U5977 (N_5977,N_5370,N_5519);
nand U5978 (N_5978,N_5277,N_5556);
xor U5979 (N_5979,N_5456,N_5508);
and U5980 (N_5980,N_5403,N_5583);
and U5981 (N_5981,N_5404,N_5362);
and U5982 (N_5982,N_5207,N_5419);
nand U5983 (N_5983,N_5461,N_5500);
or U5984 (N_5984,N_5526,N_5269);
and U5985 (N_5985,N_5516,N_5530);
nor U5986 (N_5986,N_5345,N_5305);
nor U5987 (N_5987,N_5561,N_5362);
or U5988 (N_5988,N_5520,N_5553);
and U5989 (N_5989,N_5585,N_5281);
nand U5990 (N_5990,N_5225,N_5464);
or U5991 (N_5991,N_5562,N_5214);
and U5992 (N_5992,N_5331,N_5513);
nor U5993 (N_5993,N_5456,N_5419);
nor U5994 (N_5994,N_5250,N_5555);
nor U5995 (N_5995,N_5401,N_5575);
xor U5996 (N_5996,N_5490,N_5387);
nor U5997 (N_5997,N_5528,N_5579);
nor U5998 (N_5998,N_5220,N_5330);
and U5999 (N_5999,N_5571,N_5468);
nand U6000 (N_6000,N_5748,N_5713);
xor U6001 (N_6001,N_5891,N_5699);
and U6002 (N_6002,N_5808,N_5636);
xor U6003 (N_6003,N_5942,N_5710);
xor U6004 (N_6004,N_5773,N_5766);
nand U6005 (N_6005,N_5859,N_5733);
nand U6006 (N_6006,N_5805,N_5902);
nor U6007 (N_6007,N_5620,N_5921);
or U6008 (N_6008,N_5867,N_5819);
xnor U6009 (N_6009,N_5799,N_5789);
xnor U6010 (N_6010,N_5793,N_5880);
and U6011 (N_6011,N_5760,N_5953);
xor U6012 (N_6012,N_5745,N_5767);
nand U6013 (N_6013,N_5944,N_5955);
nor U6014 (N_6014,N_5926,N_5654);
nor U6015 (N_6015,N_5976,N_5701);
or U6016 (N_6016,N_5833,N_5885);
xnor U6017 (N_6017,N_5650,N_5844);
nand U6018 (N_6018,N_5632,N_5837);
nand U6019 (N_6019,N_5898,N_5712);
nor U6020 (N_6020,N_5879,N_5858);
and U6021 (N_6021,N_5659,N_5915);
nor U6022 (N_6022,N_5616,N_5769);
nor U6023 (N_6023,N_5897,N_5910);
and U6024 (N_6024,N_5857,N_5903);
xnor U6025 (N_6025,N_5887,N_5978);
xnor U6026 (N_6026,N_5724,N_5652);
xor U6027 (N_6027,N_5801,N_5983);
nand U6028 (N_6028,N_5618,N_5909);
nand U6029 (N_6029,N_5900,N_5992);
xor U6030 (N_6030,N_5875,N_5817);
nor U6031 (N_6031,N_5856,N_5969);
and U6032 (N_6032,N_5706,N_5991);
or U6033 (N_6033,N_5619,N_5904);
nor U6034 (N_6034,N_5623,N_5873);
and U6035 (N_6035,N_5923,N_5684);
nand U6036 (N_6036,N_5762,N_5695);
nor U6037 (N_6037,N_5912,N_5931);
nand U6038 (N_6038,N_5606,N_5839);
and U6039 (N_6039,N_5641,N_5602);
xor U6040 (N_6040,N_5664,N_5899);
nor U6041 (N_6041,N_5917,N_5611);
xnor U6042 (N_6042,N_5711,N_5657);
xnor U6043 (N_6043,N_5826,N_5963);
nand U6044 (N_6044,N_5780,N_5845);
nor U6045 (N_6045,N_5673,N_5852);
xor U6046 (N_6046,N_5696,N_5802);
nor U6047 (N_6047,N_5851,N_5661);
or U6048 (N_6048,N_5613,N_5718);
and U6049 (N_6049,N_5959,N_5646);
or U6050 (N_6050,N_5688,N_5896);
or U6051 (N_6051,N_5700,N_5964);
nor U6052 (N_6052,N_5617,N_5601);
or U6053 (N_6053,N_5866,N_5888);
xor U6054 (N_6054,N_5849,N_5776);
nand U6055 (N_6055,N_5807,N_5989);
nor U6056 (N_6056,N_5750,N_5666);
xor U6057 (N_6057,N_5968,N_5810);
nor U6058 (N_6058,N_5994,N_5665);
xor U6059 (N_6059,N_5631,N_5947);
nand U6060 (N_6060,N_5816,N_5850);
nor U6061 (N_6061,N_5941,N_5907);
nand U6062 (N_6062,N_5752,N_5691);
nor U6063 (N_6063,N_5723,N_5615);
xor U6064 (N_6064,N_5894,N_5985);
nand U6065 (N_6065,N_5999,N_5715);
and U6066 (N_6066,N_5779,N_5952);
xnor U6067 (N_6067,N_5981,N_5627);
xnor U6068 (N_6068,N_5677,N_5756);
and U6069 (N_6069,N_5672,N_5694);
xnor U6070 (N_6070,N_5751,N_5683);
xnor U6071 (N_6071,N_5922,N_5640);
or U6072 (N_6072,N_5737,N_5932);
nand U6073 (N_6073,N_5872,N_5704);
nand U6074 (N_6074,N_5772,N_5739);
xnor U6075 (N_6075,N_5831,N_5809);
and U6076 (N_6076,N_5972,N_5609);
nor U6077 (N_6077,N_5720,N_5645);
or U6078 (N_6078,N_5693,N_5804);
nand U6079 (N_6079,N_5884,N_5823);
nor U6080 (N_6080,N_5697,N_5919);
and U6081 (N_6081,N_5945,N_5876);
xnor U6082 (N_6082,N_5729,N_5689);
nand U6083 (N_6083,N_5814,N_5763);
nand U6084 (N_6084,N_5675,N_5916);
xnor U6085 (N_6085,N_5822,N_5800);
nand U6086 (N_6086,N_5956,N_5803);
nor U6087 (N_6087,N_5768,N_5868);
and U6088 (N_6088,N_5883,N_5993);
nand U6089 (N_6089,N_5795,N_5753);
xor U6090 (N_6090,N_5749,N_5946);
and U6091 (N_6091,N_5667,N_5626);
xnor U6092 (N_6092,N_5863,N_5882);
or U6093 (N_6093,N_5893,N_5997);
nor U6094 (N_6094,N_5927,N_5854);
nor U6095 (N_6095,N_5797,N_5920);
nand U6096 (N_6096,N_5928,N_5629);
or U6097 (N_6097,N_5612,N_5986);
xor U6098 (N_6098,N_5977,N_5658);
nor U6099 (N_6099,N_5950,N_5744);
nor U6100 (N_6100,N_5643,N_5990);
nand U6101 (N_6101,N_5965,N_5791);
nor U6102 (N_6102,N_5934,N_5975);
nor U6103 (N_6103,N_5624,N_5656);
nand U6104 (N_6104,N_5818,N_5727);
or U6105 (N_6105,N_5841,N_5958);
or U6106 (N_6106,N_5832,N_5638);
or U6107 (N_6107,N_5970,N_5600);
or U6108 (N_6108,N_5951,N_5735);
xor U6109 (N_6109,N_5628,N_5625);
nor U6110 (N_6110,N_5703,N_5669);
and U6111 (N_6111,N_5709,N_5871);
xnor U6112 (N_6112,N_5930,N_5778);
nor U6113 (N_6113,N_5954,N_5686);
xor U6114 (N_6114,N_5905,N_5812);
nor U6115 (N_6115,N_5614,N_5639);
and U6116 (N_6116,N_5821,N_5878);
nand U6117 (N_6117,N_5716,N_5906);
or U6118 (N_6118,N_5813,N_5864);
and U6119 (N_6119,N_5676,N_5651);
xor U6120 (N_6120,N_5936,N_5792);
and U6121 (N_6121,N_5732,N_5759);
xor U6122 (N_6122,N_5662,N_5765);
xor U6123 (N_6123,N_5913,N_5847);
nor U6124 (N_6124,N_5815,N_5775);
and U6125 (N_6125,N_5860,N_5730);
xor U6126 (N_6126,N_5908,N_5787);
xnor U6127 (N_6127,N_5874,N_5770);
nand U6128 (N_6128,N_5848,N_5644);
nor U6129 (N_6129,N_5742,N_5961);
xor U6130 (N_6130,N_5634,N_5996);
or U6131 (N_6131,N_5734,N_5853);
xnor U6132 (N_6132,N_5731,N_5830);
nor U6133 (N_6133,N_5648,N_5929);
xnor U6134 (N_6134,N_5855,N_5726);
and U6135 (N_6135,N_5971,N_5877);
nand U6136 (N_6136,N_5973,N_5892);
xor U6137 (N_6137,N_5608,N_5834);
and U6138 (N_6138,N_5806,N_5870);
and U6139 (N_6139,N_5663,N_5987);
or U6140 (N_6140,N_5670,N_5924);
or U6141 (N_6141,N_5707,N_5796);
xor U6142 (N_6142,N_5777,N_5633);
nand U6143 (N_6143,N_5918,N_5988);
nand U6144 (N_6144,N_5842,N_5719);
and U6145 (N_6145,N_5869,N_5682);
or U6146 (N_6146,N_5743,N_5722);
or U6147 (N_6147,N_5943,N_5740);
and U6148 (N_6148,N_5714,N_5604);
or U6149 (N_6149,N_5671,N_5798);
nand U6150 (N_6150,N_5678,N_5702);
nand U6151 (N_6151,N_5690,N_5755);
xnor U6152 (N_6152,N_5785,N_5933);
xor U6153 (N_6153,N_5794,N_5736);
and U6154 (N_6154,N_5642,N_5914);
nand U6155 (N_6155,N_5980,N_5680);
and U6156 (N_6156,N_5825,N_5746);
xnor U6157 (N_6157,N_5901,N_5846);
xnor U6158 (N_6158,N_5966,N_5843);
nor U6159 (N_6159,N_5911,N_5962);
xnor U6160 (N_6160,N_5747,N_5705);
or U6161 (N_6161,N_5741,N_5895);
or U6162 (N_6162,N_5838,N_5948);
nor U6163 (N_6163,N_5786,N_5774);
and U6164 (N_6164,N_5649,N_5653);
nand U6165 (N_6165,N_5840,N_5984);
and U6166 (N_6166,N_5998,N_5610);
nand U6167 (N_6167,N_5674,N_5655);
and U6168 (N_6168,N_5783,N_5788);
nor U6169 (N_6169,N_5757,N_5647);
nor U6170 (N_6170,N_5728,N_5721);
nand U6171 (N_6171,N_5660,N_5949);
nand U6172 (N_6172,N_5865,N_5938);
xor U6173 (N_6173,N_5758,N_5824);
nand U6174 (N_6174,N_5708,N_5637);
and U6175 (N_6175,N_5764,N_5605);
and U6176 (N_6176,N_5681,N_5635);
xor U6177 (N_6177,N_5940,N_5754);
nor U6178 (N_6178,N_5861,N_5761);
and U6179 (N_6179,N_5607,N_5937);
or U6180 (N_6180,N_5811,N_5979);
xnor U6181 (N_6181,N_5828,N_5790);
and U6182 (N_6182,N_5630,N_5890);
nor U6183 (N_6183,N_5784,N_5925);
nor U6184 (N_6184,N_5881,N_5698);
xnor U6185 (N_6185,N_5622,N_5692);
nor U6186 (N_6186,N_5782,N_5668);
nor U6187 (N_6187,N_5960,N_5957);
and U6188 (N_6188,N_5781,N_5995);
or U6189 (N_6189,N_5725,N_5974);
nand U6190 (N_6190,N_5967,N_5679);
nor U6191 (N_6191,N_5835,N_5603);
and U6192 (N_6192,N_5687,N_5862);
nand U6193 (N_6193,N_5738,N_5820);
and U6194 (N_6194,N_5827,N_5982);
xnor U6195 (N_6195,N_5829,N_5717);
xnor U6196 (N_6196,N_5771,N_5939);
and U6197 (N_6197,N_5935,N_5886);
nand U6198 (N_6198,N_5685,N_5836);
nor U6199 (N_6199,N_5621,N_5889);
xor U6200 (N_6200,N_5755,N_5764);
and U6201 (N_6201,N_5916,N_5856);
xnor U6202 (N_6202,N_5615,N_5793);
nand U6203 (N_6203,N_5644,N_5716);
or U6204 (N_6204,N_5902,N_5875);
xnor U6205 (N_6205,N_5702,N_5906);
nor U6206 (N_6206,N_5856,N_5793);
or U6207 (N_6207,N_5944,N_5632);
or U6208 (N_6208,N_5894,N_5990);
or U6209 (N_6209,N_5729,N_5725);
or U6210 (N_6210,N_5862,N_5631);
nor U6211 (N_6211,N_5995,N_5680);
nand U6212 (N_6212,N_5687,N_5963);
nor U6213 (N_6213,N_5891,N_5617);
xor U6214 (N_6214,N_5980,N_5829);
and U6215 (N_6215,N_5818,N_5618);
xnor U6216 (N_6216,N_5759,N_5954);
xor U6217 (N_6217,N_5960,N_5764);
nand U6218 (N_6218,N_5897,N_5991);
xor U6219 (N_6219,N_5950,N_5837);
nor U6220 (N_6220,N_5811,N_5812);
nand U6221 (N_6221,N_5966,N_5975);
xnor U6222 (N_6222,N_5828,N_5937);
nand U6223 (N_6223,N_5818,N_5935);
or U6224 (N_6224,N_5786,N_5903);
and U6225 (N_6225,N_5818,N_5610);
or U6226 (N_6226,N_5893,N_5625);
or U6227 (N_6227,N_5646,N_5811);
nand U6228 (N_6228,N_5626,N_5831);
xnor U6229 (N_6229,N_5832,N_5962);
or U6230 (N_6230,N_5963,N_5673);
or U6231 (N_6231,N_5968,N_5768);
xnor U6232 (N_6232,N_5921,N_5683);
xnor U6233 (N_6233,N_5732,N_5895);
or U6234 (N_6234,N_5775,N_5738);
nor U6235 (N_6235,N_5878,N_5961);
nand U6236 (N_6236,N_5776,N_5744);
and U6237 (N_6237,N_5910,N_5886);
or U6238 (N_6238,N_5939,N_5602);
xnor U6239 (N_6239,N_5919,N_5724);
xor U6240 (N_6240,N_5891,N_5636);
and U6241 (N_6241,N_5752,N_5925);
and U6242 (N_6242,N_5772,N_5719);
or U6243 (N_6243,N_5826,N_5766);
and U6244 (N_6244,N_5763,N_5688);
nor U6245 (N_6245,N_5851,N_5933);
nand U6246 (N_6246,N_5658,N_5869);
and U6247 (N_6247,N_5951,N_5837);
nor U6248 (N_6248,N_5829,N_5786);
nand U6249 (N_6249,N_5686,N_5962);
or U6250 (N_6250,N_5834,N_5847);
xnor U6251 (N_6251,N_5835,N_5857);
and U6252 (N_6252,N_5754,N_5659);
nand U6253 (N_6253,N_5964,N_5888);
or U6254 (N_6254,N_5655,N_5753);
or U6255 (N_6255,N_5955,N_5981);
and U6256 (N_6256,N_5862,N_5886);
xnor U6257 (N_6257,N_5665,N_5802);
nor U6258 (N_6258,N_5923,N_5678);
and U6259 (N_6259,N_5699,N_5828);
and U6260 (N_6260,N_5941,N_5799);
nand U6261 (N_6261,N_5934,N_5616);
nor U6262 (N_6262,N_5888,N_5801);
nand U6263 (N_6263,N_5736,N_5757);
and U6264 (N_6264,N_5789,N_5614);
and U6265 (N_6265,N_5804,N_5835);
nand U6266 (N_6266,N_5618,N_5860);
nor U6267 (N_6267,N_5789,N_5617);
and U6268 (N_6268,N_5682,N_5841);
and U6269 (N_6269,N_5701,N_5734);
nand U6270 (N_6270,N_5834,N_5833);
or U6271 (N_6271,N_5723,N_5894);
or U6272 (N_6272,N_5978,N_5838);
nand U6273 (N_6273,N_5776,N_5730);
nor U6274 (N_6274,N_5792,N_5712);
and U6275 (N_6275,N_5723,N_5952);
xnor U6276 (N_6276,N_5851,N_5924);
xor U6277 (N_6277,N_5681,N_5751);
or U6278 (N_6278,N_5870,N_5654);
nor U6279 (N_6279,N_5617,N_5855);
xnor U6280 (N_6280,N_5828,N_5636);
and U6281 (N_6281,N_5698,N_5906);
and U6282 (N_6282,N_5698,N_5826);
and U6283 (N_6283,N_5682,N_5829);
and U6284 (N_6284,N_5786,N_5811);
nand U6285 (N_6285,N_5877,N_5886);
and U6286 (N_6286,N_5843,N_5780);
nand U6287 (N_6287,N_5948,N_5991);
nor U6288 (N_6288,N_5945,N_5858);
xnor U6289 (N_6289,N_5892,N_5622);
and U6290 (N_6290,N_5780,N_5761);
nand U6291 (N_6291,N_5770,N_5640);
or U6292 (N_6292,N_5905,N_5937);
or U6293 (N_6293,N_5827,N_5722);
nand U6294 (N_6294,N_5761,N_5887);
nor U6295 (N_6295,N_5736,N_5854);
nor U6296 (N_6296,N_5934,N_5872);
nor U6297 (N_6297,N_5882,N_5869);
xnor U6298 (N_6298,N_5777,N_5866);
and U6299 (N_6299,N_5619,N_5870);
or U6300 (N_6300,N_5754,N_5727);
and U6301 (N_6301,N_5653,N_5741);
or U6302 (N_6302,N_5979,N_5600);
and U6303 (N_6303,N_5782,N_5791);
xor U6304 (N_6304,N_5947,N_5887);
nor U6305 (N_6305,N_5658,N_5884);
and U6306 (N_6306,N_5757,N_5712);
and U6307 (N_6307,N_5698,N_5959);
and U6308 (N_6308,N_5621,N_5728);
and U6309 (N_6309,N_5995,N_5945);
and U6310 (N_6310,N_5608,N_5975);
nand U6311 (N_6311,N_5839,N_5703);
nor U6312 (N_6312,N_5857,N_5972);
and U6313 (N_6313,N_5848,N_5957);
xor U6314 (N_6314,N_5823,N_5968);
nor U6315 (N_6315,N_5982,N_5986);
xnor U6316 (N_6316,N_5800,N_5690);
xnor U6317 (N_6317,N_5710,N_5830);
nor U6318 (N_6318,N_5887,N_5928);
nor U6319 (N_6319,N_5960,N_5845);
and U6320 (N_6320,N_5968,N_5977);
xnor U6321 (N_6321,N_5973,N_5947);
and U6322 (N_6322,N_5899,N_5846);
and U6323 (N_6323,N_5734,N_5882);
nor U6324 (N_6324,N_5682,N_5717);
nor U6325 (N_6325,N_5743,N_5831);
nand U6326 (N_6326,N_5749,N_5904);
nor U6327 (N_6327,N_5983,N_5919);
nor U6328 (N_6328,N_5852,N_5666);
nor U6329 (N_6329,N_5814,N_5699);
or U6330 (N_6330,N_5797,N_5816);
nor U6331 (N_6331,N_5899,N_5853);
or U6332 (N_6332,N_5666,N_5987);
or U6333 (N_6333,N_5731,N_5900);
nor U6334 (N_6334,N_5747,N_5827);
xor U6335 (N_6335,N_5961,N_5698);
nand U6336 (N_6336,N_5798,N_5766);
nand U6337 (N_6337,N_5849,N_5708);
nand U6338 (N_6338,N_5931,N_5761);
and U6339 (N_6339,N_5793,N_5846);
nor U6340 (N_6340,N_5784,N_5960);
nand U6341 (N_6341,N_5992,N_5805);
and U6342 (N_6342,N_5807,N_5653);
nor U6343 (N_6343,N_5855,N_5804);
or U6344 (N_6344,N_5945,N_5809);
and U6345 (N_6345,N_5680,N_5749);
nor U6346 (N_6346,N_5747,N_5977);
nor U6347 (N_6347,N_5674,N_5699);
nor U6348 (N_6348,N_5657,N_5843);
nand U6349 (N_6349,N_5966,N_5625);
and U6350 (N_6350,N_5683,N_5790);
nor U6351 (N_6351,N_5874,N_5961);
nor U6352 (N_6352,N_5934,N_5750);
or U6353 (N_6353,N_5904,N_5628);
nor U6354 (N_6354,N_5662,N_5971);
nand U6355 (N_6355,N_5899,N_5952);
nor U6356 (N_6356,N_5958,N_5909);
xor U6357 (N_6357,N_5875,N_5870);
xnor U6358 (N_6358,N_5968,N_5692);
nor U6359 (N_6359,N_5672,N_5615);
nor U6360 (N_6360,N_5671,N_5761);
nand U6361 (N_6361,N_5635,N_5685);
or U6362 (N_6362,N_5961,N_5741);
xor U6363 (N_6363,N_5846,N_5983);
nor U6364 (N_6364,N_5763,N_5769);
nand U6365 (N_6365,N_5740,N_5718);
xor U6366 (N_6366,N_5795,N_5853);
nor U6367 (N_6367,N_5744,N_5717);
or U6368 (N_6368,N_5894,N_5675);
xnor U6369 (N_6369,N_5873,N_5676);
nor U6370 (N_6370,N_5791,N_5677);
xnor U6371 (N_6371,N_5904,N_5866);
xnor U6372 (N_6372,N_5969,N_5862);
nand U6373 (N_6373,N_5753,N_5684);
and U6374 (N_6374,N_5847,N_5765);
nand U6375 (N_6375,N_5709,N_5976);
nand U6376 (N_6376,N_5658,N_5848);
nor U6377 (N_6377,N_5636,N_5877);
xor U6378 (N_6378,N_5728,N_5852);
nand U6379 (N_6379,N_5988,N_5971);
or U6380 (N_6380,N_5940,N_5985);
and U6381 (N_6381,N_5744,N_5716);
xor U6382 (N_6382,N_5955,N_5692);
or U6383 (N_6383,N_5660,N_5850);
nand U6384 (N_6384,N_5838,N_5711);
xnor U6385 (N_6385,N_5841,N_5788);
or U6386 (N_6386,N_5649,N_5882);
and U6387 (N_6387,N_5788,N_5760);
or U6388 (N_6388,N_5893,N_5810);
nand U6389 (N_6389,N_5637,N_5890);
xnor U6390 (N_6390,N_5740,N_5683);
nor U6391 (N_6391,N_5773,N_5799);
or U6392 (N_6392,N_5914,N_5751);
nand U6393 (N_6393,N_5821,N_5775);
or U6394 (N_6394,N_5667,N_5841);
and U6395 (N_6395,N_5885,N_5988);
and U6396 (N_6396,N_5992,N_5936);
xnor U6397 (N_6397,N_5651,N_5936);
xnor U6398 (N_6398,N_5961,N_5845);
and U6399 (N_6399,N_5873,N_5643);
and U6400 (N_6400,N_6296,N_6215);
nor U6401 (N_6401,N_6186,N_6279);
xnor U6402 (N_6402,N_6132,N_6046);
and U6403 (N_6403,N_6115,N_6317);
nor U6404 (N_6404,N_6360,N_6056);
xnor U6405 (N_6405,N_6208,N_6345);
and U6406 (N_6406,N_6103,N_6228);
xnor U6407 (N_6407,N_6098,N_6383);
nand U6408 (N_6408,N_6151,N_6323);
and U6409 (N_6409,N_6124,N_6045);
and U6410 (N_6410,N_6367,N_6162);
xnor U6411 (N_6411,N_6169,N_6100);
and U6412 (N_6412,N_6220,N_6280);
and U6413 (N_6413,N_6313,N_6200);
nand U6414 (N_6414,N_6356,N_6217);
xor U6415 (N_6415,N_6000,N_6222);
or U6416 (N_6416,N_6157,N_6051);
xor U6417 (N_6417,N_6391,N_6010);
nor U6418 (N_6418,N_6156,N_6246);
nand U6419 (N_6419,N_6226,N_6073);
nor U6420 (N_6420,N_6030,N_6096);
and U6421 (N_6421,N_6397,N_6389);
xnor U6422 (N_6422,N_6348,N_6372);
nand U6423 (N_6423,N_6362,N_6193);
and U6424 (N_6424,N_6231,N_6335);
xnor U6425 (N_6425,N_6137,N_6057);
and U6426 (N_6426,N_6190,N_6181);
or U6427 (N_6427,N_6330,N_6252);
nor U6428 (N_6428,N_6387,N_6080);
nor U6429 (N_6429,N_6067,N_6224);
xor U6430 (N_6430,N_6159,N_6202);
or U6431 (N_6431,N_6072,N_6239);
xor U6432 (N_6432,N_6150,N_6248);
nand U6433 (N_6433,N_6295,N_6095);
or U6434 (N_6434,N_6020,N_6061);
nand U6435 (N_6435,N_6087,N_6235);
nand U6436 (N_6436,N_6140,N_6089);
nand U6437 (N_6437,N_6354,N_6049);
or U6438 (N_6438,N_6039,N_6191);
or U6439 (N_6439,N_6188,N_6034);
and U6440 (N_6440,N_6017,N_6244);
xor U6441 (N_6441,N_6309,N_6301);
or U6442 (N_6442,N_6324,N_6086);
nor U6443 (N_6443,N_6138,N_6171);
or U6444 (N_6444,N_6349,N_6319);
xnor U6445 (N_6445,N_6037,N_6161);
and U6446 (N_6446,N_6303,N_6371);
or U6447 (N_6447,N_6281,N_6163);
nand U6448 (N_6448,N_6021,N_6343);
nor U6449 (N_6449,N_6198,N_6154);
xnor U6450 (N_6450,N_6088,N_6366);
xor U6451 (N_6451,N_6311,N_6358);
nand U6452 (N_6452,N_6338,N_6192);
xor U6453 (N_6453,N_6376,N_6218);
xnor U6454 (N_6454,N_6363,N_6275);
xnor U6455 (N_6455,N_6286,N_6346);
nand U6456 (N_6456,N_6395,N_6238);
xnor U6457 (N_6457,N_6187,N_6052);
or U6458 (N_6458,N_6143,N_6083);
nor U6459 (N_6459,N_6111,N_6055);
and U6460 (N_6460,N_6204,N_6022);
nand U6461 (N_6461,N_6031,N_6069);
and U6462 (N_6462,N_6084,N_6318);
nor U6463 (N_6463,N_6347,N_6002);
or U6464 (N_6464,N_6058,N_6274);
nor U6465 (N_6465,N_6093,N_6199);
and U6466 (N_6466,N_6108,N_6203);
xnor U6467 (N_6467,N_6266,N_6306);
nor U6468 (N_6468,N_6062,N_6234);
xnor U6469 (N_6469,N_6079,N_6059);
and U6470 (N_6470,N_6283,N_6113);
nand U6471 (N_6471,N_6129,N_6265);
nor U6472 (N_6472,N_6322,N_6101);
and U6473 (N_6473,N_6142,N_6160);
nor U6474 (N_6474,N_6178,N_6305);
nor U6475 (N_6475,N_6044,N_6126);
or U6476 (N_6476,N_6141,N_6382);
xor U6477 (N_6477,N_6078,N_6085);
nand U6478 (N_6478,N_6251,N_6229);
or U6479 (N_6479,N_6119,N_6260);
or U6480 (N_6480,N_6380,N_6298);
nand U6481 (N_6481,N_6024,N_6291);
and U6482 (N_6482,N_6247,N_6201);
and U6483 (N_6483,N_6352,N_6353);
xor U6484 (N_6484,N_6092,N_6091);
xor U6485 (N_6485,N_6326,N_6120);
nor U6486 (N_6486,N_6219,N_6174);
xor U6487 (N_6487,N_6134,N_6048);
xnor U6488 (N_6488,N_6253,N_6036);
nor U6489 (N_6489,N_6249,N_6003);
nor U6490 (N_6490,N_6015,N_6148);
xor U6491 (N_6491,N_6336,N_6107);
and U6492 (N_6492,N_6340,N_6370);
nor U6493 (N_6493,N_6018,N_6118);
nor U6494 (N_6494,N_6077,N_6212);
nand U6495 (N_6495,N_6355,N_6243);
nand U6496 (N_6496,N_6026,N_6070);
nand U6497 (N_6497,N_6339,N_6043);
nor U6498 (N_6498,N_6232,N_6384);
nand U6499 (N_6499,N_6377,N_6144);
xnor U6500 (N_6500,N_6292,N_6196);
or U6501 (N_6501,N_6385,N_6230);
and U6502 (N_6502,N_6344,N_6005);
xor U6503 (N_6503,N_6259,N_6104);
nand U6504 (N_6504,N_6158,N_6097);
nor U6505 (N_6505,N_6105,N_6206);
or U6506 (N_6506,N_6315,N_6109);
nor U6507 (N_6507,N_6040,N_6165);
and U6508 (N_6508,N_6331,N_6236);
nand U6509 (N_6509,N_6321,N_6237);
nand U6510 (N_6510,N_6012,N_6288);
nor U6511 (N_6511,N_6378,N_6361);
nor U6512 (N_6512,N_6271,N_6337);
or U6513 (N_6513,N_6241,N_6147);
nand U6514 (N_6514,N_6130,N_6307);
or U6515 (N_6515,N_6168,N_6155);
xnor U6516 (N_6516,N_6145,N_6262);
xnor U6517 (N_6517,N_6197,N_6029);
or U6518 (N_6518,N_6233,N_6110);
nor U6519 (N_6519,N_6270,N_6277);
xnor U6520 (N_6520,N_6175,N_6250);
nand U6521 (N_6521,N_6304,N_6269);
nand U6522 (N_6522,N_6257,N_6334);
or U6523 (N_6523,N_6261,N_6006);
and U6524 (N_6524,N_6060,N_6041);
or U6525 (N_6525,N_6013,N_6146);
xor U6526 (N_6526,N_6106,N_6364);
or U6527 (N_6527,N_6112,N_6254);
nor U6528 (N_6528,N_6068,N_6133);
xor U6529 (N_6529,N_6374,N_6082);
nand U6530 (N_6530,N_6267,N_6263);
nand U6531 (N_6531,N_6293,N_6242);
nor U6532 (N_6532,N_6127,N_6221);
or U6533 (N_6533,N_6170,N_6121);
and U6534 (N_6534,N_6302,N_6278);
xor U6535 (N_6535,N_6185,N_6205);
xnor U6536 (N_6536,N_6167,N_6123);
xnor U6537 (N_6537,N_6179,N_6054);
nor U6538 (N_6538,N_6365,N_6064);
xor U6539 (N_6539,N_6042,N_6063);
xnor U6540 (N_6540,N_6379,N_6125);
xor U6541 (N_6541,N_6182,N_6194);
or U6542 (N_6542,N_6299,N_6386);
nor U6543 (N_6543,N_6394,N_6001);
and U6544 (N_6544,N_6038,N_6240);
or U6545 (N_6545,N_6223,N_6189);
nor U6546 (N_6546,N_6327,N_6245);
nand U6547 (N_6547,N_6350,N_6359);
xor U6548 (N_6548,N_6272,N_6164);
or U6549 (N_6549,N_6341,N_6053);
or U6550 (N_6550,N_6268,N_6128);
nand U6551 (N_6551,N_6312,N_6396);
nor U6552 (N_6552,N_6342,N_6008);
nand U6553 (N_6553,N_6289,N_6153);
or U6554 (N_6554,N_6183,N_6195);
or U6555 (N_6555,N_6284,N_6264);
or U6556 (N_6556,N_6066,N_6149);
nor U6557 (N_6557,N_6300,N_6290);
nor U6558 (N_6558,N_6294,N_6357);
xor U6559 (N_6559,N_6392,N_6102);
nor U6560 (N_6560,N_6116,N_6035);
xnor U6561 (N_6561,N_6032,N_6025);
and U6562 (N_6562,N_6375,N_6173);
xor U6563 (N_6563,N_6065,N_6177);
and U6564 (N_6564,N_6152,N_6393);
nand U6565 (N_6565,N_6213,N_6381);
nand U6566 (N_6566,N_6273,N_6282);
and U6567 (N_6567,N_6076,N_6184);
nand U6568 (N_6568,N_6297,N_6131);
xor U6569 (N_6569,N_6004,N_6325);
and U6570 (N_6570,N_6287,N_6332);
or U6571 (N_6571,N_6074,N_6207);
nand U6572 (N_6572,N_6211,N_6176);
or U6573 (N_6573,N_6023,N_6047);
and U6574 (N_6574,N_6310,N_6314);
and U6575 (N_6575,N_6050,N_6368);
xnor U6576 (N_6576,N_6216,N_6373);
nand U6577 (N_6577,N_6014,N_6320);
nor U6578 (N_6578,N_6210,N_6328);
or U6579 (N_6579,N_6090,N_6081);
or U6580 (N_6580,N_6136,N_6390);
nor U6581 (N_6581,N_6258,N_6028);
nor U6582 (N_6582,N_6369,N_6316);
xnor U6583 (N_6583,N_6007,N_6308);
and U6584 (N_6584,N_6094,N_6256);
xor U6585 (N_6585,N_6399,N_6180);
and U6586 (N_6586,N_6333,N_6099);
or U6587 (N_6587,N_6135,N_6075);
xnor U6588 (N_6588,N_6114,N_6172);
and U6589 (N_6589,N_6209,N_6388);
nand U6590 (N_6590,N_6016,N_6329);
and U6591 (N_6591,N_6227,N_6276);
or U6592 (N_6592,N_6166,N_6011);
nor U6593 (N_6593,N_6139,N_6351);
nand U6594 (N_6594,N_6122,N_6225);
nand U6595 (N_6595,N_6398,N_6019);
and U6596 (N_6596,N_6009,N_6285);
xor U6597 (N_6597,N_6071,N_6117);
or U6598 (N_6598,N_6027,N_6033);
nand U6599 (N_6599,N_6214,N_6255);
nor U6600 (N_6600,N_6088,N_6305);
or U6601 (N_6601,N_6158,N_6247);
and U6602 (N_6602,N_6351,N_6021);
nand U6603 (N_6603,N_6230,N_6368);
or U6604 (N_6604,N_6093,N_6390);
nor U6605 (N_6605,N_6003,N_6099);
xnor U6606 (N_6606,N_6040,N_6366);
nand U6607 (N_6607,N_6189,N_6067);
nand U6608 (N_6608,N_6104,N_6091);
xor U6609 (N_6609,N_6388,N_6195);
nand U6610 (N_6610,N_6054,N_6234);
nand U6611 (N_6611,N_6313,N_6358);
xor U6612 (N_6612,N_6271,N_6381);
nor U6613 (N_6613,N_6062,N_6095);
nor U6614 (N_6614,N_6062,N_6236);
or U6615 (N_6615,N_6229,N_6033);
xor U6616 (N_6616,N_6208,N_6210);
nand U6617 (N_6617,N_6233,N_6192);
xnor U6618 (N_6618,N_6282,N_6295);
nand U6619 (N_6619,N_6043,N_6038);
xnor U6620 (N_6620,N_6009,N_6357);
and U6621 (N_6621,N_6044,N_6196);
or U6622 (N_6622,N_6062,N_6219);
and U6623 (N_6623,N_6242,N_6047);
nor U6624 (N_6624,N_6012,N_6016);
and U6625 (N_6625,N_6347,N_6159);
nor U6626 (N_6626,N_6313,N_6213);
and U6627 (N_6627,N_6316,N_6212);
nor U6628 (N_6628,N_6077,N_6377);
or U6629 (N_6629,N_6112,N_6014);
or U6630 (N_6630,N_6292,N_6076);
xor U6631 (N_6631,N_6383,N_6376);
or U6632 (N_6632,N_6122,N_6350);
nand U6633 (N_6633,N_6140,N_6238);
xor U6634 (N_6634,N_6187,N_6129);
or U6635 (N_6635,N_6338,N_6288);
nor U6636 (N_6636,N_6340,N_6048);
and U6637 (N_6637,N_6392,N_6071);
and U6638 (N_6638,N_6265,N_6226);
nand U6639 (N_6639,N_6306,N_6357);
xnor U6640 (N_6640,N_6215,N_6247);
nor U6641 (N_6641,N_6103,N_6182);
or U6642 (N_6642,N_6243,N_6232);
or U6643 (N_6643,N_6013,N_6056);
nor U6644 (N_6644,N_6322,N_6227);
and U6645 (N_6645,N_6284,N_6322);
or U6646 (N_6646,N_6150,N_6353);
nand U6647 (N_6647,N_6029,N_6295);
nor U6648 (N_6648,N_6043,N_6099);
or U6649 (N_6649,N_6372,N_6046);
and U6650 (N_6650,N_6089,N_6064);
xnor U6651 (N_6651,N_6150,N_6169);
xnor U6652 (N_6652,N_6304,N_6205);
nand U6653 (N_6653,N_6163,N_6055);
nand U6654 (N_6654,N_6153,N_6333);
nor U6655 (N_6655,N_6204,N_6300);
nand U6656 (N_6656,N_6309,N_6267);
or U6657 (N_6657,N_6199,N_6145);
nor U6658 (N_6658,N_6119,N_6125);
xor U6659 (N_6659,N_6250,N_6261);
and U6660 (N_6660,N_6152,N_6391);
nand U6661 (N_6661,N_6209,N_6160);
xnor U6662 (N_6662,N_6258,N_6336);
or U6663 (N_6663,N_6109,N_6311);
and U6664 (N_6664,N_6277,N_6252);
nor U6665 (N_6665,N_6364,N_6235);
and U6666 (N_6666,N_6289,N_6148);
or U6667 (N_6667,N_6285,N_6203);
nand U6668 (N_6668,N_6042,N_6318);
and U6669 (N_6669,N_6205,N_6394);
nor U6670 (N_6670,N_6368,N_6206);
or U6671 (N_6671,N_6351,N_6123);
nand U6672 (N_6672,N_6030,N_6203);
nor U6673 (N_6673,N_6038,N_6254);
nor U6674 (N_6674,N_6221,N_6210);
and U6675 (N_6675,N_6262,N_6283);
xnor U6676 (N_6676,N_6077,N_6256);
and U6677 (N_6677,N_6277,N_6249);
xnor U6678 (N_6678,N_6043,N_6311);
or U6679 (N_6679,N_6341,N_6041);
nand U6680 (N_6680,N_6368,N_6021);
nor U6681 (N_6681,N_6113,N_6134);
nor U6682 (N_6682,N_6205,N_6082);
xnor U6683 (N_6683,N_6064,N_6284);
xor U6684 (N_6684,N_6162,N_6117);
nor U6685 (N_6685,N_6372,N_6226);
or U6686 (N_6686,N_6054,N_6364);
or U6687 (N_6687,N_6053,N_6067);
nor U6688 (N_6688,N_6258,N_6223);
or U6689 (N_6689,N_6227,N_6105);
or U6690 (N_6690,N_6355,N_6312);
xnor U6691 (N_6691,N_6208,N_6028);
nand U6692 (N_6692,N_6153,N_6079);
nor U6693 (N_6693,N_6217,N_6338);
xnor U6694 (N_6694,N_6160,N_6324);
nor U6695 (N_6695,N_6088,N_6091);
or U6696 (N_6696,N_6165,N_6385);
or U6697 (N_6697,N_6273,N_6081);
and U6698 (N_6698,N_6234,N_6214);
xnor U6699 (N_6699,N_6193,N_6376);
nor U6700 (N_6700,N_6103,N_6058);
xor U6701 (N_6701,N_6392,N_6105);
or U6702 (N_6702,N_6376,N_6186);
nor U6703 (N_6703,N_6088,N_6370);
nand U6704 (N_6704,N_6168,N_6025);
or U6705 (N_6705,N_6386,N_6280);
nor U6706 (N_6706,N_6328,N_6179);
and U6707 (N_6707,N_6099,N_6204);
nor U6708 (N_6708,N_6360,N_6195);
nor U6709 (N_6709,N_6212,N_6051);
xor U6710 (N_6710,N_6193,N_6130);
and U6711 (N_6711,N_6160,N_6195);
nand U6712 (N_6712,N_6349,N_6326);
nor U6713 (N_6713,N_6032,N_6333);
xnor U6714 (N_6714,N_6306,N_6137);
nor U6715 (N_6715,N_6163,N_6293);
nor U6716 (N_6716,N_6039,N_6038);
xor U6717 (N_6717,N_6209,N_6115);
xnor U6718 (N_6718,N_6152,N_6330);
nor U6719 (N_6719,N_6068,N_6151);
xnor U6720 (N_6720,N_6381,N_6375);
nand U6721 (N_6721,N_6302,N_6164);
nor U6722 (N_6722,N_6061,N_6353);
nand U6723 (N_6723,N_6133,N_6173);
nor U6724 (N_6724,N_6271,N_6179);
xor U6725 (N_6725,N_6165,N_6246);
xnor U6726 (N_6726,N_6144,N_6049);
nor U6727 (N_6727,N_6256,N_6092);
and U6728 (N_6728,N_6149,N_6344);
nor U6729 (N_6729,N_6188,N_6109);
nand U6730 (N_6730,N_6240,N_6374);
nand U6731 (N_6731,N_6329,N_6076);
xor U6732 (N_6732,N_6399,N_6308);
nand U6733 (N_6733,N_6009,N_6265);
nand U6734 (N_6734,N_6011,N_6306);
or U6735 (N_6735,N_6315,N_6001);
nor U6736 (N_6736,N_6195,N_6381);
nand U6737 (N_6737,N_6237,N_6369);
and U6738 (N_6738,N_6294,N_6001);
nand U6739 (N_6739,N_6179,N_6350);
nor U6740 (N_6740,N_6351,N_6003);
nand U6741 (N_6741,N_6061,N_6324);
nor U6742 (N_6742,N_6259,N_6054);
and U6743 (N_6743,N_6327,N_6203);
and U6744 (N_6744,N_6150,N_6335);
nor U6745 (N_6745,N_6118,N_6199);
nor U6746 (N_6746,N_6374,N_6032);
xnor U6747 (N_6747,N_6250,N_6235);
nor U6748 (N_6748,N_6270,N_6130);
nor U6749 (N_6749,N_6017,N_6373);
nand U6750 (N_6750,N_6058,N_6145);
nor U6751 (N_6751,N_6241,N_6368);
xnor U6752 (N_6752,N_6355,N_6039);
and U6753 (N_6753,N_6337,N_6354);
and U6754 (N_6754,N_6350,N_6157);
or U6755 (N_6755,N_6069,N_6180);
xnor U6756 (N_6756,N_6076,N_6204);
nand U6757 (N_6757,N_6147,N_6337);
and U6758 (N_6758,N_6081,N_6220);
xnor U6759 (N_6759,N_6164,N_6093);
nand U6760 (N_6760,N_6088,N_6120);
nor U6761 (N_6761,N_6003,N_6037);
and U6762 (N_6762,N_6050,N_6358);
xor U6763 (N_6763,N_6288,N_6317);
or U6764 (N_6764,N_6393,N_6335);
or U6765 (N_6765,N_6276,N_6108);
nand U6766 (N_6766,N_6285,N_6149);
nand U6767 (N_6767,N_6033,N_6248);
and U6768 (N_6768,N_6255,N_6187);
xnor U6769 (N_6769,N_6398,N_6364);
nand U6770 (N_6770,N_6266,N_6319);
xor U6771 (N_6771,N_6245,N_6382);
nand U6772 (N_6772,N_6366,N_6087);
nor U6773 (N_6773,N_6264,N_6194);
or U6774 (N_6774,N_6002,N_6167);
nand U6775 (N_6775,N_6246,N_6268);
or U6776 (N_6776,N_6162,N_6036);
nand U6777 (N_6777,N_6008,N_6113);
nor U6778 (N_6778,N_6089,N_6296);
xnor U6779 (N_6779,N_6297,N_6097);
and U6780 (N_6780,N_6381,N_6126);
and U6781 (N_6781,N_6340,N_6270);
xor U6782 (N_6782,N_6200,N_6051);
xor U6783 (N_6783,N_6070,N_6010);
or U6784 (N_6784,N_6152,N_6290);
xnor U6785 (N_6785,N_6088,N_6189);
nor U6786 (N_6786,N_6397,N_6324);
nand U6787 (N_6787,N_6175,N_6247);
xor U6788 (N_6788,N_6131,N_6324);
or U6789 (N_6789,N_6174,N_6125);
nor U6790 (N_6790,N_6057,N_6024);
or U6791 (N_6791,N_6272,N_6010);
nand U6792 (N_6792,N_6039,N_6015);
and U6793 (N_6793,N_6245,N_6087);
nand U6794 (N_6794,N_6206,N_6052);
nand U6795 (N_6795,N_6269,N_6247);
xor U6796 (N_6796,N_6253,N_6273);
and U6797 (N_6797,N_6025,N_6045);
nand U6798 (N_6798,N_6246,N_6063);
or U6799 (N_6799,N_6087,N_6232);
xnor U6800 (N_6800,N_6730,N_6495);
nor U6801 (N_6801,N_6517,N_6700);
xor U6802 (N_6802,N_6455,N_6512);
xor U6803 (N_6803,N_6647,N_6741);
and U6804 (N_6804,N_6651,N_6697);
nor U6805 (N_6805,N_6779,N_6487);
nor U6806 (N_6806,N_6702,N_6532);
nor U6807 (N_6807,N_6780,N_6614);
nor U6808 (N_6808,N_6719,N_6635);
or U6809 (N_6809,N_6688,N_6555);
nand U6810 (N_6810,N_6692,N_6563);
xnor U6811 (N_6811,N_6744,N_6416);
nand U6812 (N_6812,N_6794,N_6403);
nor U6813 (N_6813,N_6645,N_6498);
xnor U6814 (N_6814,N_6727,N_6690);
xnor U6815 (N_6815,N_6570,N_6504);
and U6816 (N_6816,N_6634,N_6765);
and U6817 (N_6817,N_6595,N_6400);
xnor U6818 (N_6818,N_6522,N_6511);
or U6819 (N_6819,N_6716,N_6772);
nand U6820 (N_6820,N_6592,N_6476);
or U6821 (N_6821,N_6432,N_6798);
nor U6822 (N_6822,N_6714,N_6444);
and U6823 (N_6823,N_6650,N_6593);
xnor U6824 (N_6824,N_6795,N_6457);
and U6825 (N_6825,N_6732,N_6435);
or U6826 (N_6826,N_6408,N_6470);
nand U6827 (N_6827,N_6685,N_6679);
nand U6828 (N_6828,N_6789,N_6648);
xor U6829 (N_6829,N_6499,N_6680);
nand U6830 (N_6830,N_6670,N_6740);
nand U6831 (N_6831,N_6469,N_6756);
xnor U6832 (N_6832,N_6754,N_6663);
nand U6833 (N_6833,N_6622,N_6747);
or U6834 (N_6834,N_6790,N_6673);
or U6835 (N_6835,N_6560,N_6567);
and U6836 (N_6836,N_6429,N_6607);
nor U6837 (N_6837,N_6462,N_6632);
nor U6838 (N_6838,N_6571,N_6610);
xnor U6839 (N_6839,N_6581,N_6646);
and U6840 (N_6840,N_6691,N_6753);
xnor U6841 (N_6841,N_6551,N_6694);
xnor U6842 (N_6842,N_6686,N_6676);
xnor U6843 (N_6843,N_6475,N_6681);
or U6844 (N_6844,N_6419,N_6778);
or U6845 (N_6845,N_6535,N_6643);
nand U6846 (N_6846,N_6599,N_6433);
nor U6847 (N_6847,N_6497,N_6750);
and U6848 (N_6848,N_6713,N_6710);
nand U6849 (N_6849,N_6451,N_6585);
and U6850 (N_6850,N_6545,N_6652);
nor U6851 (N_6851,N_6678,N_6482);
nor U6852 (N_6852,N_6709,N_6786);
or U6853 (N_6853,N_6547,N_6699);
nor U6854 (N_6854,N_6423,N_6496);
xor U6855 (N_6855,N_6401,N_6544);
nor U6856 (N_6856,N_6724,N_6683);
xor U6857 (N_6857,N_6549,N_6528);
nor U6858 (N_6858,N_6600,N_6757);
or U6859 (N_6859,N_6708,N_6565);
and U6860 (N_6860,N_6509,N_6474);
and U6861 (N_6861,N_6494,N_6760);
and U6862 (N_6862,N_6667,N_6738);
nand U6863 (N_6863,N_6630,N_6684);
or U6864 (N_6864,N_6717,N_6426);
nor U6865 (N_6865,N_6440,N_6589);
nor U6866 (N_6866,N_6639,N_6707);
xnor U6867 (N_6867,N_6471,N_6736);
nand U6868 (N_6868,N_6598,N_6442);
and U6869 (N_6869,N_6743,N_6566);
nor U6870 (N_6870,N_6590,N_6458);
or U6871 (N_6871,N_6460,N_6425);
xnor U6872 (N_6872,N_6576,N_6488);
nand U6873 (N_6873,N_6711,N_6613);
nand U6874 (N_6874,N_6568,N_6759);
xnor U6875 (N_6875,N_6627,N_6580);
nor U6876 (N_6876,N_6562,N_6529);
or U6877 (N_6877,N_6775,N_6594);
nand U6878 (N_6878,N_6503,N_6480);
xnor U6879 (N_6879,N_6749,N_6438);
or U6880 (N_6880,N_6505,N_6659);
and U6881 (N_6881,N_6418,N_6669);
nand U6882 (N_6882,N_6543,N_6409);
and U6883 (N_6883,N_6412,N_6611);
nor U6884 (N_6884,N_6490,N_6770);
xnor U6885 (N_6885,N_6797,N_6604);
or U6886 (N_6886,N_6771,N_6675);
or U6887 (N_6887,N_6703,N_6596);
and U6888 (N_6888,N_6665,N_6406);
xor U6889 (N_6889,N_6662,N_6661);
nand U6890 (N_6890,N_6453,N_6449);
nand U6891 (N_6891,N_6653,N_6636);
or U6892 (N_6892,N_6561,N_6620);
or U6893 (N_6893,N_6446,N_6784);
xor U6894 (N_6894,N_6459,N_6584);
or U6895 (N_6895,N_6542,N_6623);
or U6896 (N_6896,N_6410,N_6552);
xor U6897 (N_6897,N_6564,N_6452);
xnor U6898 (N_6898,N_6587,N_6486);
and U6899 (N_6899,N_6621,N_6417);
nand U6900 (N_6900,N_6510,N_6572);
and U6901 (N_6901,N_6658,N_6774);
or U6902 (N_6902,N_6725,N_6407);
nand U6903 (N_6903,N_6461,N_6722);
nor U6904 (N_6904,N_6721,N_6609);
nand U6905 (N_6905,N_6540,N_6637);
nand U6906 (N_6906,N_6484,N_6558);
nand U6907 (N_6907,N_6448,N_6728);
nor U6908 (N_6908,N_6715,N_6538);
or U6909 (N_6909,N_6640,N_6616);
nor U6910 (N_6910,N_6783,N_6421);
or U6911 (N_6911,N_6597,N_6657);
nor U6912 (N_6912,N_6633,N_6785);
xor U6913 (N_6913,N_6704,N_6631);
and U6914 (N_6914,N_6427,N_6641);
nand U6915 (N_6915,N_6649,N_6508);
nor U6916 (N_6916,N_6588,N_6574);
and U6917 (N_6917,N_6625,N_6553);
or U6918 (N_6918,N_6519,N_6521);
xnor U6919 (N_6919,N_6674,N_6537);
xnor U6920 (N_6920,N_6737,N_6660);
xnor U6921 (N_6921,N_6642,N_6726);
nor U6922 (N_6922,N_6735,N_6404);
nand U6923 (N_6923,N_6729,N_6533);
xnor U6924 (N_6924,N_6605,N_6733);
nor U6925 (N_6925,N_6677,N_6472);
nor U6926 (N_6926,N_6769,N_6437);
nor U6927 (N_6927,N_6734,N_6424);
nand U6928 (N_6928,N_6706,N_6513);
and U6929 (N_6929,N_6463,N_6582);
nand U6930 (N_6930,N_6550,N_6698);
xor U6931 (N_6931,N_6479,N_6671);
nand U6932 (N_6932,N_6693,N_6583);
nor U6933 (N_6933,N_6525,N_6602);
nand U6934 (N_6934,N_6799,N_6739);
and U6935 (N_6935,N_6477,N_6644);
or U6936 (N_6936,N_6447,N_6465);
or U6937 (N_6937,N_6422,N_6501);
and U6938 (N_6938,N_6468,N_6788);
and U6939 (N_6939,N_6420,N_6695);
xnor U6940 (N_6940,N_6485,N_6655);
nand U6941 (N_6941,N_6656,N_6742);
nor U6942 (N_6942,N_6762,N_6758);
nand U6943 (N_6943,N_6578,N_6626);
nand U6944 (N_6944,N_6405,N_6776);
and U6945 (N_6945,N_6518,N_6664);
nand U6946 (N_6946,N_6615,N_6624);
and U6947 (N_6947,N_6668,N_6763);
and U6948 (N_6948,N_6539,N_6767);
nand U6949 (N_6949,N_6450,N_6515);
nor U6950 (N_6950,N_6575,N_6516);
nor U6951 (N_6951,N_6434,N_6723);
and U6952 (N_6952,N_6573,N_6796);
nor U6953 (N_6953,N_6439,N_6415);
nand U6954 (N_6954,N_6531,N_6491);
nor U6955 (N_6955,N_6608,N_6687);
nand U6956 (N_6956,N_6617,N_6773);
and U6957 (N_6957,N_6428,N_6492);
nand U6958 (N_6958,N_6689,N_6793);
nand U6959 (N_6959,N_6791,N_6466);
nor U6960 (N_6960,N_6445,N_6530);
nor U6961 (N_6961,N_6523,N_6546);
and U6962 (N_6962,N_6441,N_6751);
nand U6963 (N_6963,N_6478,N_6705);
and U6964 (N_6964,N_6764,N_6654);
or U6965 (N_6965,N_6557,N_6554);
or U6966 (N_6966,N_6489,N_6507);
and U6967 (N_6967,N_6629,N_6638);
or U6968 (N_6968,N_6601,N_6493);
and U6969 (N_6969,N_6483,N_6748);
nand U6970 (N_6970,N_6586,N_6569);
xor U6971 (N_6971,N_6787,N_6527);
or U6972 (N_6972,N_6454,N_6752);
nor U6973 (N_6973,N_6520,N_6473);
xnor U6974 (N_6974,N_6696,N_6506);
or U6975 (N_6975,N_6536,N_6402);
xor U6976 (N_6976,N_6731,N_6792);
xnor U6977 (N_6977,N_6606,N_6712);
and U6978 (N_6978,N_6430,N_6718);
nand U6979 (N_6979,N_6618,N_6502);
or U6980 (N_6980,N_6526,N_6720);
and U6981 (N_6981,N_6746,N_6548);
and U6982 (N_6982,N_6591,N_6755);
xnor U6983 (N_6983,N_6514,N_6411);
nor U6984 (N_6984,N_6782,N_6436);
xnor U6985 (N_6985,N_6524,N_6414);
xor U6986 (N_6986,N_6761,N_6781);
xor U6987 (N_6987,N_6534,N_6766);
or U6988 (N_6988,N_6768,N_6431);
nor U6989 (N_6989,N_6559,N_6579);
nand U6990 (N_6990,N_6413,N_6464);
nor U6991 (N_6991,N_6577,N_6777);
xor U6992 (N_6992,N_6467,N_6672);
xnor U6993 (N_6993,N_6443,N_6619);
or U6994 (N_6994,N_6612,N_6456);
nor U6995 (N_6995,N_6541,N_6556);
or U6996 (N_6996,N_6682,N_6666);
or U6997 (N_6997,N_6603,N_6628);
or U6998 (N_6998,N_6701,N_6745);
nor U6999 (N_6999,N_6500,N_6481);
and U7000 (N_7000,N_6465,N_6758);
nor U7001 (N_7001,N_6593,N_6471);
or U7002 (N_7002,N_6666,N_6405);
and U7003 (N_7003,N_6767,N_6447);
or U7004 (N_7004,N_6769,N_6707);
and U7005 (N_7005,N_6416,N_6728);
or U7006 (N_7006,N_6636,N_6408);
and U7007 (N_7007,N_6571,N_6784);
and U7008 (N_7008,N_6757,N_6633);
xnor U7009 (N_7009,N_6734,N_6404);
and U7010 (N_7010,N_6658,N_6562);
or U7011 (N_7011,N_6482,N_6618);
nand U7012 (N_7012,N_6655,N_6593);
xnor U7013 (N_7013,N_6640,N_6674);
nor U7014 (N_7014,N_6735,N_6546);
xor U7015 (N_7015,N_6654,N_6758);
nand U7016 (N_7016,N_6779,N_6623);
nand U7017 (N_7017,N_6429,N_6441);
or U7018 (N_7018,N_6691,N_6680);
nor U7019 (N_7019,N_6501,N_6607);
xor U7020 (N_7020,N_6436,N_6478);
xor U7021 (N_7021,N_6659,N_6596);
or U7022 (N_7022,N_6498,N_6786);
nor U7023 (N_7023,N_6441,N_6767);
or U7024 (N_7024,N_6647,N_6500);
nor U7025 (N_7025,N_6432,N_6636);
or U7026 (N_7026,N_6524,N_6780);
nand U7027 (N_7027,N_6795,N_6638);
and U7028 (N_7028,N_6683,N_6674);
nor U7029 (N_7029,N_6612,N_6744);
xor U7030 (N_7030,N_6546,N_6633);
nand U7031 (N_7031,N_6418,N_6529);
xor U7032 (N_7032,N_6505,N_6775);
xnor U7033 (N_7033,N_6547,N_6632);
or U7034 (N_7034,N_6576,N_6626);
nor U7035 (N_7035,N_6526,N_6654);
nand U7036 (N_7036,N_6673,N_6468);
nand U7037 (N_7037,N_6611,N_6440);
nor U7038 (N_7038,N_6647,N_6798);
or U7039 (N_7039,N_6665,N_6485);
and U7040 (N_7040,N_6425,N_6431);
and U7041 (N_7041,N_6756,N_6586);
nor U7042 (N_7042,N_6408,N_6421);
or U7043 (N_7043,N_6408,N_6519);
and U7044 (N_7044,N_6579,N_6558);
xnor U7045 (N_7045,N_6463,N_6581);
xnor U7046 (N_7046,N_6772,N_6569);
nand U7047 (N_7047,N_6550,N_6407);
xnor U7048 (N_7048,N_6450,N_6704);
nor U7049 (N_7049,N_6476,N_6604);
nor U7050 (N_7050,N_6518,N_6513);
nand U7051 (N_7051,N_6470,N_6692);
nand U7052 (N_7052,N_6655,N_6521);
and U7053 (N_7053,N_6518,N_6738);
or U7054 (N_7054,N_6790,N_6752);
and U7055 (N_7055,N_6737,N_6512);
or U7056 (N_7056,N_6496,N_6788);
and U7057 (N_7057,N_6503,N_6605);
and U7058 (N_7058,N_6681,N_6467);
and U7059 (N_7059,N_6573,N_6517);
and U7060 (N_7060,N_6427,N_6760);
nand U7061 (N_7061,N_6793,N_6412);
or U7062 (N_7062,N_6469,N_6624);
nor U7063 (N_7063,N_6427,N_6587);
nor U7064 (N_7064,N_6530,N_6594);
and U7065 (N_7065,N_6710,N_6692);
xor U7066 (N_7066,N_6774,N_6489);
and U7067 (N_7067,N_6553,N_6498);
nor U7068 (N_7068,N_6679,N_6501);
and U7069 (N_7069,N_6725,N_6783);
and U7070 (N_7070,N_6452,N_6457);
or U7071 (N_7071,N_6408,N_6688);
or U7072 (N_7072,N_6542,N_6767);
nand U7073 (N_7073,N_6591,N_6425);
nand U7074 (N_7074,N_6651,N_6440);
or U7075 (N_7075,N_6746,N_6739);
or U7076 (N_7076,N_6435,N_6704);
nor U7077 (N_7077,N_6435,N_6727);
and U7078 (N_7078,N_6718,N_6588);
and U7079 (N_7079,N_6656,N_6743);
xnor U7080 (N_7080,N_6485,N_6719);
and U7081 (N_7081,N_6586,N_6615);
nor U7082 (N_7082,N_6539,N_6694);
and U7083 (N_7083,N_6639,N_6664);
and U7084 (N_7084,N_6616,N_6403);
and U7085 (N_7085,N_6491,N_6636);
or U7086 (N_7086,N_6700,N_6681);
or U7087 (N_7087,N_6478,N_6689);
xor U7088 (N_7088,N_6544,N_6526);
xor U7089 (N_7089,N_6419,N_6773);
or U7090 (N_7090,N_6754,N_6769);
nand U7091 (N_7091,N_6652,N_6442);
or U7092 (N_7092,N_6640,N_6594);
nor U7093 (N_7093,N_6477,N_6708);
nor U7094 (N_7094,N_6697,N_6788);
nand U7095 (N_7095,N_6780,N_6435);
xnor U7096 (N_7096,N_6631,N_6464);
and U7097 (N_7097,N_6638,N_6488);
nand U7098 (N_7098,N_6715,N_6719);
or U7099 (N_7099,N_6747,N_6573);
nand U7100 (N_7100,N_6743,N_6616);
and U7101 (N_7101,N_6676,N_6784);
nor U7102 (N_7102,N_6744,N_6737);
and U7103 (N_7103,N_6495,N_6714);
and U7104 (N_7104,N_6425,N_6437);
nor U7105 (N_7105,N_6734,N_6548);
xnor U7106 (N_7106,N_6597,N_6617);
nand U7107 (N_7107,N_6522,N_6675);
nand U7108 (N_7108,N_6556,N_6774);
nand U7109 (N_7109,N_6537,N_6554);
or U7110 (N_7110,N_6649,N_6619);
and U7111 (N_7111,N_6761,N_6740);
and U7112 (N_7112,N_6507,N_6482);
nand U7113 (N_7113,N_6683,N_6614);
nand U7114 (N_7114,N_6473,N_6527);
or U7115 (N_7115,N_6605,N_6593);
xor U7116 (N_7116,N_6590,N_6688);
nand U7117 (N_7117,N_6434,N_6762);
and U7118 (N_7118,N_6798,N_6795);
or U7119 (N_7119,N_6692,N_6722);
or U7120 (N_7120,N_6461,N_6630);
nor U7121 (N_7121,N_6425,N_6421);
nand U7122 (N_7122,N_6450,N_6430);
nor U7123 (N_7123,N_6506,N_6719);
xnor U7124 (N_7124,N_6449,N_6550);
or U7125 (N_7125,N_6478,N_6420);
xor U7126 (N_7126,N_6439,N_6642);
xor U7127 (N_7127,N_6442,N_6503);
xor U7128 (N_7128,N_6655,N_6543);
nor U7129 (N_7129,N_6421,N_6532);
nor U7130 (N_7130,N_6602,N_6544);
or U7131 (N_7131,N_6441,N_6753);
nand U7132 (N_7132,N_6626,N_6544);
nor U7133 (N_7133,N_6416,N_6606);
nor U7134 (N_7134,N_6431,N_6714);
or U7135 (N_7135,N_6754,N_6685);
and U7136 (N_7136,N_6521,N_6401);
or U7137 (N_7137,N_6766,N_6444);
nor U7138 (N_7138,N_6435,N_6565);
or U7139 (N_7139,N_6744,N_6734);
and U7140 (N_7140,N_6503,N_6798);
nand U7141 (N_7141,N_6706,N_6711);
nand U7142 (N_7142,N_6587,N_6657);
xnor U7143 (N_7143,N_6682,N_6764);
xor U7144 (N_7144,N_6486,N_6446);
xor U7145 (N_7145,N_6590,N_6674);
xor U7146 (N_7146,N_6455,N_6710);
nand U7147 (N_7147,N_6764,N_6404);
and U7148 (N_7148,N_6710,N_6473);
and U7149 (N_7149,N_6678,N_6743);
and U7150 (N_7150,N_6679,N_6723);
and U7151 (N_7151,N_6477,N_6769);
xnor U7152 (N_7152,N_6620,N_6419);
nor U7153 (N_7153,N_6581,N_6689);
and U7154 (N_7154,N_6534,N_6652);
or U7155 (N_7155,N_6513,N_6544);
nor U7156 (N_7156,N_6613,N_6707);
and U7157 (N_7157,N_6447,N_6701);
and U7158 (N_7158,N_6784,N_6452);
or U7159 (N_7159,N_6781,N_6775);
nand U7160 (N_7160,N_6579,N_6587);
or U7161 (N_7161,N_6699,N_6565);
or U7162 (N_7162,N_6755,N_6791);
and U7163 (N_7163,N_6695,N_6585);
nor U7164 (N_7164,N_6796,N_6640);
nor U7165 (N_7165,N_6422,N_6724);
nor U7166 (N_7166,N_6690,N_6537);
or U7167 (N_7167,N_6735,N_6650);
and U7168 (N_7168,N_6452,N_6586);
nand U7169 (N_7169,N_6457,N_6533);
or U7170 (N_7170,N_6764,N_6507);
xnor U7171 (N_7171,N_6447,N_6650);
nand U7172 (N_7172,N_6417,N_6495);
nor U7173 (N_7173,N_6598,N_6606);
nor U7174 (N_7174,N_6464,N_6727);
nor U7175 (N_7175,N_6693,N_6792);
xor U7176 (N_7176,N_6729,N_6421);
and U7177 (N_7177,N_6796,N_6448);
nor U7178 (N_7178,N_6423,N_6627);
or U7179 (N_7179,N_6529,N_6600);
or U7180 (N_7180,N_6527,N_6480);
xor U7181 (N_7181,N_6510,N_6486);
nor U7182 (N_7182,N_6766,N_6692);
nor U7183 (N_7183,N_6759,N_6716);
xor U7184 (N_7184,N_6791,N_6488);
xor U7185 (N_7185,N_6651,N_6511);
nor U7186 (N_7186,N_6665,N_6681);
or U7187 (N_7187,N_6623,N_6521);
and U7188 (N_7188,N_6726,N_6678);
nand U7189 (N_7189,N_6548,N_6583);
or U7190 (N_7190,N_6703,N_6563);
or U7191 (N_7191,N_6719,N_6626);
xor U7192 (N_7192,N_6754,N_6467);
and U7193 (N_7193,N_6706,N_6507);
nand U7194 (N_7194,N_6449,N_6749);
and U7195 (N_7195,N_6450,N_6579);
and U7196 (N_7196,N_6448,N_6698);
nor U7197 (N_7197,N_6427,N_6598);
nor U7198 (N_7198,N_6720,N_6541);
xor U7199 (N_7199,N_6411,N_6524);
xnor U7200 (N_7200,N_7174,N_7128);
nand U7201 (N_7201,N_6812,N_7161);
nor U7202 (N_7202,N_7119,N_7168);
or U7203 (N_7203,N_7077,N_6940);
or U7204 (N_7204,N_7156,N_6874);
and U7205 (N_7205,N_6868,N_6901);
xnor U7206 (N_7206,N_7023,N_6831);
nand U7207 (N_7207,N_6918,N_7140);
and U7208 (N_7208,N_6904,N_6991);
or U7209 (N_7209,N_7016,N_7052);
xnor U7210 (N_7210,N_7005,N_6948);
and U7211 (N_7211,N_6898,N_6866);
nand U7212 (N_7212,N_6951,N_7107);
and U7213 (N_7213,N_6969,N_6893);
or U7214 (N_7214,N_6808,N_6835);
and U7215 (N_7215,N_6900,N_7046);
or U7216 (N_7216,N_6955,N_6894);
xor U7217 (N_7217,N_7183,N_6859);
xor U7218 (N_7218,N_7059,N_6828);
xnor U7219 (N_7219,N_6892,N_6897);
xor U7220 (N_7220,N_7191,N_7143);
and U7221 (N_7221,N_7181,N_6838);
and U7222 (N_7222,N_7007,N_6875);
xnor U7223 (N_7223,N_7086,N_6978);
nand U7224 (N_7224,N_7083,N_7134);
nor U7225 (N_7225,N_6878,N_7159);
and U7226 (N_7226,N_7149,N_7045);
and U7227 (N_7227,N_6819,N_7067);
nand U7228 (N_7228,N_7188,N_7082);
nor U7229 (N_7229,N_6843,N_6881);
nand U7230 (N_7230,N_7163,N_7121);
nor U7231 (N_7231,N_6959,N_6864);
xor U7232 (N_7232,N_7173,N_6999);
nor U7233 (N_7233,N_7177,N_6899);
and U7234 (N_7234,N_7195,N_7003);
xnor U7235 (N_7235,N_6932,N_7141);
or U7236 (N_7236,N_7055,N_6954);
nor U7237 (N_7237,N_6925,N_6912);
and U7238 (N_7238,N_6994,N_6818);
xor U7239 (N_7239,N_6858,N_6852);
nor U7240 (N_7240,N_6891,N_6846);
nor U7241 (N_7241,N_7166,N_6884);
nor U7242 (N_7242,N_6889,N_7115);
and U7243 (N_7243,N_7095,N_7014);
and U7244 (N_7244,N_6847,N_6953);
nand U7245 (N_7245,N_7013,N_7085);
xnor U7246 (N_7246,N_7145,N_7006);
xor U7247 (N_7247,N_6957,N_6934);
xor U7248 (N_7248,N_7136,N_6807);
nand U7249 (N_7249,N_6865,N_7099);
xnor U7250 (N_7250,N_6817,N_6887);
and U7251 (N_7251,N_7147,N_6990);
xor U7252 (N_7252,N_6809,N_7030);
xor U7253 (N_7253,N_7132,N_7087);
nor U7254 (N_7254,N_6811,N_7127);
xnor U7255 (N_7255,N_7092,N_6933);
nor U7256 (N_7256,N_7196,N_6824);
and U7257 (N_7257,N_7021,N_7028);
or U7258 (N_7258,N_6802,N_7024);
or U7259 (N_7259,N_6939,N_7053);
nand U7260 (N_7260,N_6869,N_7084);
xnor U7261 (N_7261,N_6872,N_7144);
nor U7262 (N_7262,N_6930,N_7069);
xnor U7263 (N_7263,N_6942,N_7135);
and U7264 (N_7264,N_6801,N_7138);
or U7265 (N_7265,N_6924,N_6938);
or U7266 (N_7266,N_7043,N_6840);
nand U7267 (N_7267,N_6810,N_6814);
nand U7268 (N_7268,N_6982,N_6826);
or U7269 (N_7269,N_7039,N_6863);
or U7270 (N_7270,N_6946,N_7190);
nor U7271 (N_7271,N_6945,N_6970);
or U7272 (N_7272,N_7026,N_6806);
nor U7273 (N_7273,N_7027,N_7063);
or U7274 (N_7274,N_7198,N_7088);
xor U7275 (N_7275,N_7105,N_6989);
and U7276 (N_7276,N_6964,N_6979);
nand U7277 (N_7277,N_7098,N_6841);
xor U7278 (N_7278,N_7126,N_7194);
nand U7279 (N_7279,N_7012,N_7150);
xor U7280 (N_7280,N_7076,N_6913);
nand U7281 (N_7281,N_6935,N_7189);
xor U7282 (N_7282,N_6976,N_7186);
xnor U7283 (N_7283,N_7112,N_7050);
and U7284 (N_7284,N_6823,N_7057);
and U7285 (N_7285,N_6879,N_6856);
xnor U7286 (N_7286,N_7151,N_6839);
xnor U7287 (N_7287,N_7080,N_6848);
or U7288 (N_7288,N_7116,N_7049);
nand U7289 (N_7289,N_6820,N_6917);
xor U7290 (N_7290,N_6937,N_7068);
and U7291 (N_7291,N_7096,N_6877);
and U7292 (N_7292,N_7032,N_7022);
or U7293 (N_7293,N_7008,N_6963);
nor U7294 (N_7294,N_6803,N_7036);
xnor U7295 (N_7295,N_6886,N_6880);
nand U7296 (N_7296,N_6983,N_6950);
nand U7297 (N_7297,N_6860,N_7125);
and U7298 (N_7298,N_6830,N_7160);
or U7299 (N_7299,N_7172,N_7179);
nand U7300 (N_7300,N_7031,N_6927);
nand U7301 (N_7301,N_7010,N_6921);
nor U7302 (N_7302,N_6903,N_7169);
and U7303 (N_7303,N_7019,N_7009);
or U7304 (N_7304,N_7040,N_7101);
or U7305 (N_7305,N_7081,N_7062);
or U7306 (N_7306,N_6914,N_7109);
xor U7307 (N_7307,N_6958,N_7035);
nor U7308 (N_7308,N_7075,N_6853);
or U7309 (N_7309,N_7122,N_7180);
nor U7310 (N_7310,N_7018,N_6906);
xor U7311 (N_7311,N_6896,N_7094);
or U7312 (N_7312,N_6861,N_7090);
nor U7313 (N_7313,N_6873,N_6949);
nor U7314 (N_7314,N_7193,N_7142);
or U7315 (N_7315,N_7089,N_6973);
nor U7316 (N_7316,N_6952,N_6966);
and U7317 (N_7317,N_7114,N_7111);
and U7318 (N_7318,N_6908,N_6890);
nor U7319 (N_7319,N_6911,N_6975);
xor U7320 (N_7320,N_7029,N_7146);
nor U7321 (N_7321,N_7118,N_6922);
nand U7322 (N_7322,N_6876,N_6936);
or U7323 (N_7323,N_7041,N_6928);
or U7324 (N_7324,N_7167,N_6834);
nor U7325 (N_7325,N_6895,N_7165);
nor U7326 (N_7326,N_7154,N_6905);
and U7327 (N_7327,N_7102,N_7001);
or U7328 (N_7328,N_6915,N_7199);
and U7329 (N_7329,N_6816,N_7072);
nand U7330 (N_7330,N_6870,N_6855);
nand U7331 (N_7331,N_6832,N_7170);
xnor U7332 (N_7332,N_7171,N_6993);
and U7333 (N_7333,N_6800,N_7108);
xnor U7334 (N_7334,N_6998,N_6919);
nor U7335 (N_7335,N_6926,N_6995);
and U7336 (N_7336,N_7185,N_7056);
or U7337 (N_7337,N_7157,N_7162);
and U7338 (N_7338,N_7061,N_7131);
nand U7339 (N_7339,N_7164,N_7187);
or U7340 (N_7340,N_7123,N_6986);
and U7341 (N_7341,N_7079,N_6947);
nor U7342 (N_7342,N_7025,N_6943);
nor U7343 (N_7343,N_7197,N_7002);
xor U7344 (N_7344,N_6849,N_6837);
nand U7345 (N_7345,N_7033,N_7192);
and U7346 (N_7346,N_6965,N_6972);
nor U7347 (N_7347,N_6885,N_6821);
nor U7348 (N_7348,N_6845,N_6968);
and U7349 (N_7349,N_6804,N_7182);
xor U7350 (N_7350,N_6974,N_6854);
nand U7351 (N_7351,N_7106,N_7133);
xor U7352 (N_7352,N_6836,N_7065);
and U7353 (N_7353,N_6813,N_6844);
and U7354 (N_7354,N_6829,N_7139);
nand U7355 (N_7355,N_6850,N_6987);
nand U7356 (N_7356,N_6825,N_6827);
nand U7357 (N_7357,N_6851,N_7017);
and U7358 (N_7358,N_6977,N_7176);
and U7359 (N_7359,N_7037,N_7097);
or U7360 (N_7360,N_6882,N_6971);
xnor U7361 (N_7361,N_7048,N_7060);
nor U7362 (N_7362,N_7078,N_6902);
or U7363 (N_7363,N_7155,N_7070);
or U7364 (N_7364,N_7042,N_6862);
or U7365 (N_7365,N_7178,N_6984);
nand U7366 (N_7366,N_7093,N_7047);
or U7367 (N_7367,N_6920,N_6822);
and U7368 (N_7368,N_7104,N_6944);
nor U7369 (N_7369,N_6962,N_7038);
nand U7370 (N_7370,N_6929,N_6960);
and U7371 (N_7371,N_6871,N_7020);
nand U7372 (N_7372,N_6996,N_7015);
and U7373 (N_7373,N_6980,N_6923);
or U7374 (N_7374,N_7058,N_6857);
nand U7375 (N_7375,N_6985,N_6833);
nand U7376 (N_7376,N_7158,N_7175);
nand U7377 (N_7377,N_6910,N_7064);
or U7378 (N_7378,N_6956,N_7117);
xor U7379 (N_7379,N_7044,N_7100);
or U7380 (N_7380,N_6992,N_7113);
nand U7381 (N_7381,N_7110,N_7011);
nor U7382 (N_7382,N_6997,N_6888);
nand U7383 (N_7383,N_6931,N_6805);
and U7384 (N_7384,N_7054,N_6883);
xnor U7385 (N_7385,N_6988,N_6941);
xor U7386 (N_7386,N_6961,N_6916);
nand U7387 (N_7387,N_7034,N_7130);
and U7388 (N_7388,N_6909,N_7152);
or U7389 (N_7389,N_7004,N_6815);
nand U7390 (N_7390,N_7071,N_7184);
xnor U7391 (N_7391,N_7051,N_7074);
and U7392 (N_7392,N_7148,N_7091);
nor U7393 (N_7393,N_6907,N_7124);
xnor U7394 (N_7394,N_7073,N_7153);
xnor U7395 (N_7395,N_6981,N_6867);
nand U7396 (N_7396,N_7137,N_6967);
nand U7397 (N_7397,N_7103,N_7129);
nand U7398 (N_7398,N_7000,N_7066);
nor U7399 (N_7399,N_7120,N_6842);
and U7400 (N_7400,N_7061,N_7000);
nor U7401 (N_7401,N_6960,N_7143);
or U7402 (N_7402,N_7070,N_7118);
xor U7403 (N_7403,N_7068,N_7148);
or U7404 (N_7404,N_6934,N_7023);
nor U7405 (N_7405,N_7090,N_6893);
nand U7406 (N_7406,N_7059,N_6993);
nor U7407 (N_7407,N_6882,N_6943);
nand U7408 (N_7408,N_6902,N_6809);
xnor U7409 (N_7409,N_7127,N_7053);
nand U7410 (N_7410,N_6875,N_7010);
nor U7411 (N_7411,N_7076,N_7123);
nor U7412 (N_7412,N_6965,N_7133);
nand U7413 (N_7413,N_7195,N_6857);
nand U7414 (N_7414,N_6921,N_6804);
nand U7415 (N_7415,N_6932,N_6843);
xnor U7416 (N_7416,N_7053,N_6962);
nor U7417 (N_7417,N_7179,N_7057);
xor U7418 (N_7418,N_6873,N_7125);
or U7419 (N_7419,N_6999,N_7133);
or U7420 (N_7420,N_7107,N_7133);
nand U7421 (N_7421,N_6972,N_7062);
xnor U7422 (N_7422,N_7112,N_6813);
xnor U7423 (N_7423,N_6944,N_6838);
and U7424 (N_7424,N_7171,N_6835);
and U7425 (N_7425,N_6857,N_7021);
nand U7426 (N_7426,N_7046,N_7029);
nand U7427 (N_7427,N_6964,N_7059);
or U7428 (N_7428,N_7134,N_7010);
nand U7429 (N_7429,N_7153,N_7115);
or U7430 (N_7430,N_7146,N_6971);
or U7431 (N_7431,N_6832,N_7138);
and U7432 (N_7432,N_7165,N_6980);
and U7433 (N_7433,N_6815,N_6825);
nand U7434 (N_7434,N_6945,N_6904);
xor U7435 (N_7435,N_6942,N_7028);
nand U7436 (N_7436,N_6812,N_6844);
or U7437 (N_7437,N_7122,N_7134);
xnor U7438 (N_7438,N_7020,N_7188);
and U7439 (N_7439,N_7134,N_7006);
and U7440 (N_7440,N_7068,N_6856);
nand U7441 (N_7441,N_7125,N_7100);
or U7442 (N_7442,N_6904,N_6923);
and U7443 (N_7443,N_7156,N_6856);
nor U7444 (N_7444,N_7082,N_7150);
xor U7445 (N_7445,N_6863,N_6861);
xnor U7446 (N_7446,N_7028,N_7026);
and U7447 (N_7447,N_7046,N_6804);
and U7448 (N_7448,N_6811,N_7001);
xor U7449 (N_7449,N_6875,N_7084);
or U7450 (N_7450,N_7025,N_7081);
xnor U7451 (N_7451,N_6844,N_7079);
xnor U7452 (N_7452,N_7040,N_6806);
nor U7453 (N_7453,N_7109,N_6829);
nand U7454 (N_7454,N_6936,N_7082);
and U7455 (N_7455,N_6831,N_6928);
nand U7456 (N_7456,N_7186,N_7048);
and U7457 (N_7457,N_6869,N_6877);
nor U7458 (N_7458,N_6833,N_7134);
or U7459 (N_7459,N_7072,N_7160);
or U7460 (N_7460,N_6882,N_6982);
or U7461 (N_7461,N_6851,N_6917);
nor U7462 (N_7462,N_6867,N_7035);
xor U7463 (N_7463,N_6875,N_7173);
nor U7464 (N_7464,N_7169,N_7032);
xnor U7465 (N_7465,N_7053,N_6971);
and U7466 (N_7466,N_6956,N_6922);
xnor U7467 (N_7467,N_7068,N_6998);
and U7468 (N_7468,N_7055,N_7126);
xor U7469 (N_7469,N_6952,N_6954);
and U7470 (N_7470,N_6946,N_7037);
xnor U7471 (N_7471,N_7174,N_7102);
or U7472 (N_7472,N_6893,N_6935);
and U7473 (N_7473,N_7042,N_6895);
or U7474 (N_7474,N_6858,N_7144);
nand U7475 (N_7475,N_7040,N_7139);
nand U7476 (N_7476,N_6926,N_7191);
nand U7477 (N_7477,N_7040,N_7051);
or U7478 (N_7478,N_7012,N_6848);
and U7479 (N_7479,N_6967,N_7149);
and U7480 (N_7480,N_6888,N_7155);
nor U7481 (N_7481,N_6922,N_7016);
and U7482 (N_7482,N_6978,N_7085);
or U7483 (N_7483,N_6989,N_6990);
nor U7484 (N_7484,N_7104,N_6954);
nor U7485 (N_7485,N_7090,N_6830);
xor U7486 (N_7486,N_6808,N_6938);
nor U7487 (N_7487,N_7000,N_7128);
and U7488 (N_7488,N_7037,N_6927);
nor U7489 (N_7489,N_6853,N_7095);
xnor U7490 (N_7490,N_6821,N_7188);
nand U7491 (N_7491,N_6916,N_6960);
or U7492 (N_7492,N_7019,N_6949);
and U7493 (N_7493,N_7033,N_6920);
nand U7494 (N_7494,N_6870,N_6862);
nor U7495 (N_7495,N_7023,N_6845);
or U7496 (N_7496,N_6837,N_7170);
nor U7497 (N_7497,N_6854,N_7018);
nor U7498 (N_7498,N_7137,N_7069);
nand U7499 (N_7499,N_6958,N_6908);
xnor U7500 (N_7500,N_6941,N_6921);
nand U7501 (N_7501,N_6885,N_6811);
or U7502 (N_7502,N_6833,N_6963);
or U7503 (N_7503,N_6981,N_6938);
or U7504 (N_7504,N_6970,N_7142);
or U7505 (N_7505,N_7092,N_7198);
xor U7506 (N_7506,N_7076,N_6877);
or U7507 (N_7507,N_6972,N_7167);
or U7508 (N_7508,N_7019,N_6889);
xnor U7509 (N_7509,N_7051,N_7000);
or U7510 (N_7510,N_7180,N_6800);
and U7511 (N_7511,N_6901,N_6802);
xnor U7512 (N_7512,N_7196,N_6989);
nor U7513 (N_7513,N_7044,N_7179);
and U7514 (N_7514,N_7036,N_6815);
xnor U7515 (N_7515,N_6802,N_6801);
nand U7516 (N_7516,N_7162,N_7102);
or U7517 (N_7517,N_7105,N_7196);
xor U7518 (N_7518,N_6981,N_6861);
nor U7519 (N_7519,N_6969,N_6856);
nand U7520 (N_7520,N_7022,N_7168);
xnor U7521 (N_7521,N_7057,N_7008);
nand U7522 (N_7522,N_7129,N_6909);
xor U7523 (N_7523,N_7020,N_7023);
nand U7524 (N_7524,N_7147,N_6817);
or U7525 (N_7525,N_6891,N_7124);
xor U7526 (N_7526,N_6842,N_7010);
and U7527 (N_7527,N_7153,N_6932);
or U7528 (N_7528,N_7087,N_6922);
nor U7529 (N_7529,N_6951,N_7148);
nor U7530 (N_7530,N_6873,N_7109);
or U7531 (N_7531,N_6946,N_7188);
nand U7532 (N_7532,N_6887,N_6833);
or U7533 (N_7533,N_7163,N_6962);
and U7534 (N_7534,N_6980,N_6845);
nand U7535 (N_7535,N_7177,N_6833);
xnor U7536 (N_7536,N_7146,N_6888);
or U7537 (N_7537,N_7147,N_7065);
nand U7538 (N_7538,N_7144,N_6957);
and U7539 (N_7539,N_6848,N_7166);
nand U7540 (N_7540,N_6938,N_6897);
nand U7541 (N_7541,N_7197,N_7112);
or U7542 (N_7542,N_6854,N_6840);
or U7543 (N_7543,N_7166,N_7171);
and U7544 (N_7544,N_7183,N_7036);
xnor U7545 (N_7545,N_7170,N_7015);
nor U7546 (N_7546,N_6848,N_6867);
nor U7547 (N_7547,N_7059,N_6839);
nand U7548 (N_7548,N_7132,N_6876);
nand U7549 (N_7549,N_7195,N_6839);
nor U7550 (N_7550,N_7182,N_7051);
xnor U7551 (N_7551,N_7004,N_7127);
nor U7552 (N_7552,N_7169,N_6809);
and U7553 (N_7553,N_7173,N_6830);
and U7554 (N_7554,N_7016,N_6944);
nor U7555 (N_7555,N_7167,N_6917);
and U7556 (N_7556,N_7144,N_7145);
nor U7557 (N_7557,N_7103,N_6910);
or U7558 (N_7558,N_7044,N_7095);
nand U7559 (N_7559,N_6810,N_6828);
xnor U7560 (N_7560,N_7055,N_6834);
and U7561 (N_7561,N_6991,N_6937);
nor U7562 (N_7562,N_6891,N_6858);
nor U7563 (N_7563,N_6914,N_7099);
and U7564 (N_7564,N_7030,N_6917);
or U7565 (N_7565,N_6946,N_6918);
nand U7566 (N_7566,N_6997,N_7100);
and U7567 (N_7567,N_7021,N_7077);
xor U7568 (N_7568,N_7181,N_6952);
xnor U7569 (N_7569,N_7186,N_6972);
xor U7570 (N_7570,N_7132,N_7073);
and U7571 (N_7571,N_6965,N_7050);
or U7572 (N_7572,N_6833,N_6960);
nor U7573 (N_7573,N_6969,N_6837);
xnor U7574 (N_7574,N_6875,N_7021);
and U7575 (N_7575,N_6868,N_7061);
nor U7576 (N_7576,N_7187,N_6952);
and U7577 (N_7577,N_7179,N_7168);
nand U7578 (N_7578,N_7078,N_6831);
or U7579 (N_7579,N_7184,N_7099);
xor U7580 (N_7580,N_6947,N_7100);
or U7581 (N_7581,N_6898,N_7160);
and U7582 (N_7582,N_6862,N_6900);
or U7583 (N_7583,N_6927,N_7097);
nor U7584 (N_7584,N_7043,N_6856);
nand U7585 (N_7585,N_6923,N_7199);
xnor U7586 (N_7586,N_7186,N_7136);
xor U7587 (N_7587,N_6913,N_7188);
nor U7588 (N_7588,N_6813,N_7172);
xnor U7589 (N_7589,N_7032,N_6862);
and U7590 (N_7590,N_6826,N_7015);
nor U7591 (N_7591,N_7083,N_7001);
nor U7592 (N_7592,N_6805,N_7093);
and U7593 (N_7593,N_6882,N_7180);
and U7594 (N_7594,N_6859,N_7153);
nand U7595 (N_7595,N_7079,N_6942);
nor U7596 (N_7596,N_7170,N_7042);
nor U7597 (N_7597,N_7016,N_7015);
and U7598 (N_7598,N_7074,N_7196);
nand U7599 (N_7599,N_7197,N_7140);
or U7600 (N_7600,N_7429,N_7233);
and U7601 (N_7601,N_7359,N_7468);
nor U7602 (N_7602,N_7524,N_7386);
nand U7603 (N_7603,N_7383,N_7477);
nor U7604 (N_7604,N_7577,N_7217);
or U7605 (N_7605,N_7377,N_7462);
and U7606 (N_7606,N_7492,N_7450);
and U7607 (N_7607,N_7240,N_7581);
xor U7608 (N_7608,N_7270,N_7481);
and U7609 (N_7609,N_7466,N_7311);
and U7610 (N_7610,N_7419,N_7446);
and U7611 (N_7611,N_7500,N_7326);
and U7612 (N_7612,N_7455,N_7243);
xnor U7613 (N_7613,N_7398,N_7545);
and U7614 (N_7614,N_7300,N_7288);
and U7615 (N_7615,N_7510,N_7213);
nor U7616 (N_7616,N_7232,N_7474);
nor U7617 (N_7617,N_7593,N_7491);
and U7618 (N_7618,N_7422,N_7253);
xnor U7619 (N_7619,N_7327,N_7360);
xnor U7620 (N_7620,N_7478,N_7285);
nand U7621 (N_7621,N_7588,N_7442);
nand U7622 (N_7622,N_7210,N_7424);
nand U7623 (N_7623,N_7597,N_7259);
nand U7624 (N_7624,N_7564,N_7301);
and U7625 (N_7625,N_7458,N_7426);
and U7626 (N_7626,N_7527,N_7599);
nor U7627 (N_7627,N_7451,N_7313);
nand U7628 (N_7628,N_7428,N_7391);
nand U7629 (N_7629,N_7512,N_7539);
xor U7630 (N_7630,N_7309,N_7333);
and U7631 (N_7631,N_7282,N_7367);
and U7632 (N_7632,N_7228,N_7485);
xnor U7633 (N_7633,N_7330,N_7387);
and U7634 (N_7634,N_7591,N_7328);
and U7635 (N_7635,N_7552,N_7268);
xnor U7636 (N_7636,N_7308,N_7337);
or U7637 (N_7637,N_7515,N_7502);
and U7638 (N_7638,N_7408,N_7252);
xor U7639 (N_7639,N_7453,N_7236);
or U7640 (N_7640,N_7237,N_7412);
nor U7641 (N_7641,N_7304,N_7521);
nand U7642 (N_7642,N_7223,N_7522);
nand U7643 (N_7643,N_7574,N_7293);
nand U7644 (N_7644,N_7427,N_7441);
xnor U7645 (N_7645,N_7516,N_7399);
or U7646 (N_7646,N_7334,N_7310);
or U7647 (N_7647,N_7518,N_7467);
or U7648 (N_7648,N_7405,N_7350);
nand U7649 (N_7649,N_7266,N_7287);
nor U7650 (N_7650,N_7595,N_7353);
and U7651 (N_7651,N_7322,N_7421);
xor U7652 (N_7652,N_7508,N_7370);
or U7653 (N_7653,N_7269,N_7303);
nand U7654 (N_7654,N_7473,N_7385);
or U7655 (N_7655,N_7275,N_7224);
nand U7656 (N_7656,N_7498,N_7382);
nand U7657 (N_7657,N_7431,N_7482);
or U7658 (N_7658,N_7592,N_7530);
and U7659 (N_7659,N_7220,N_7561);
nor U7660 (N_7660,N_7406,N_7336);
nand U7661 (N_7661,N_7415,N_7461);
or U7662 (N_7662,N_7494,N_7340);
nand U7663 (N_7663,N_7245,N_7535);
and U7664 (N_7664,N_7251,N_7576);
nand U7665 (N_7665,N_7411,N_7277);
nor U7666 (N_7666,N_7487,N_7437);
xnor U7667 (N_7667,N_7476,N_7380);
nor U7668 (N_7668,N_7436,N_7459);
or U7669 (N_7669,N_7486,N_7395);
or U7670 (N_7670,N_7258,N_7571);
nand U7671 (N_7671,N_7529,N_7205);
nand U7672 (N_7672,N_7320,N_7263);
or U7673 (N_7673,N_7509,N_7208);
or U7674 (N_7674,N_7323,N_7338);
and U7675 (N_7675,N_7452,N_7554);
nor U7676 (N_7676,N_7244,N_7432);
and U7677 (N_7677,N_7291,N_7345);
nor U7678 (N_7678,N_7302,N_7578);
and U7679 (N_7679,N_7255,N_7586);
nor U7680 (N_7680,N_7257,N_7557);
nor U7681 (N_7681,N_7381,N_7517);
nand U7682 (N_7682,N_7507,N_7409);
xor U7683 (N_7683,N_7278,N_7348);
and U7684 (N_7684,N_7443,N_7307);
and U7685 (N_7685,N_7211,N_7563);
or U7686 (N_7686,N_7339,N_7202);
or U7687 (N_7687,N_7403,N_7559);
nand U7688 (N_7688,N_7358,N_7294);
or U7689 (N_7689,N_7575,N_7549);
and U7690 (N_7690,N_7324,N_7573);
or U7691 (N_7691,N_7388,N_7531);
or U7692 (N_7692,N_7449,N_7480);
or U7693 (N_7693,N_7495,N_7548);
xnor U7694 (N_7694,N_7425,N_7538);
nand U7695 (N_7695,N_7585,N_7447);
or U7696 (N_7696,N_7582,N_7393);
nor U7697 (N_7697,N_7534,N_7225);
xor U7698 (N_7698,N_7470,N_7318);
or U7699 (N_7699,N_7506,N_7265);
and U7700 (N_7700,N_7219,N_7204);
nor U7701 (N_7701,N_7212,N_7544);
nand U7702 (N_7702,N_7404,N_7596);
nand U7703 (N_7703,N_7580,N_7400);
or U7704 (N_7704,N_7594,N_7207);
and U7705 (N_7705,N_7361,N_7357);
or U7706 (N_7706,N_7389,N_7587);
nand U7707 (N_7707,N_7368,N_7471);
xor U7708 (N_7708,N_7335,N_7469);
nand U7709 (N_7709,N_7503,N_7222);
nand U7710 (N_7710,N_7261,N_7249);
and U7711 (N_7711,N_7499,N_7364);
nand U7712 (N_7712,N_7363,N_7221);
xor U7713 (N_7713,N_7344,N_7215);
nor U7714 (N_7714,N_7438,N_7297);
or U7715 (N_7715,N_7365,N_7295);
or U7716 (N_7716,N_7292,N_7465);
or U7717 (N_7717,N_7375,N_7250);
and U7718 (N_7718,N_7369,N_7519);
xor U7719 (N_7719,N_7513,N_7341);
nand U7720 (N_7720,N_7546,N_7543);
nor U7721 (N_7721,N_7355,N_7414);
or U7722 (N_7722,N_7394,N_7281);
nor U7723 (N_7723,N_7523,N_7540);
and U7724 (N_7724,N_7315,N_7342);
and U7725 (N_7725,N_7347,N_7346);
or U7726 (N_7726,N_7464,N_7460);
or U7727 (N_7727,N_7218,N_7475);
and U7728 (N_7728,N_7314,N_7384);
or U7729 (N_7729,N_7239,N_7298);
xor U7730 (N_7730,N_7351,N_7558);
nand U7731 (N_7731,N_7454,N_7201);
nor U7732 (N_7732,N_7290,N_7520);
xnor U7733 (N_7733,N_7214,N_7456);
nand U7734 (N_7734,N_7227,N_7484);
and U7735 (N_7735,N_7584,N_7241);
nor U7736 (N_7736,N_7271,N_7306);
or U7737 (N_7737,N_7550,N_7444);
nor U7738 (N_7738,N_7490,N_7483);
and U7739 (N_7739,N_7279,N_7254);
nand U7740 (N_7740,N_7349,N_7420);
nor U7741 (N_7741,N_7296,N_7248);
nor U7742 (N_7742,N_7579,N_7238);
nor U7743 (N_7743,N_7247,N_7463);
nor U7744 (N_7744,N_7407,N_7537);
nor U7745 (N_7745,N_7590,N_7390);
or U7746 (N_7746,N_7572,N_7372);
and U7747 (N_7747,N_7566,N_7329);
and U7748 (N_7748,N_7246,N_7283);
nor U7749 (N_7749,N_7264,N_7343);
xor U7750 (N_7750,N_7362,N_7206);
nor U7751 (N_7751,N_7541,N_7435);
xor U7752 (N_7752,N_7280,N_7373);
nand U7753 (N_7753,N_7504,N_7305);
nand U7754 (N_7754,N_7583,N_7231);
and U7755 (N_7755,N_7553,N_7440);
and U7756 (N_7756,N_7472,N_7433);
and U7757 (N_7757,N_7312,N_7423);
xnor U7758 (N_7758,N_7439,N_7589);
xnor U7759 (N_7759,N_7331,N_7274);
nand U7760 (N_7760,N_7514,N_7536);
nand U7761 (N_7761,N_7289,N_7366);
nor U7762 (N_7762,N_7505,N_7569);
xor U7763 (N_7763,N_7378,N_7262);
or U7764 (N_7764,N_7321,N_7560);
nand U7765 (N_7765,N_7260,N_7488);
nor U7766 (N_7766,N_7430,N_7316);
nand U7767 (N_7767,N_7493,N_7319);
and U7768 (N_7768,N_7286,N_7570);
or U7769 (N_7769,N_7525,N_7371);
xor U7770 (N_7770,N_7379,N_7413);
or U7771 (N_7771,N_7497,N_7533);
xnor U7772 (N_7772,N_7402,N_7376);
nor U7773 (N_7773,N_7417,N_7547);
or U7774 (N_7774,N_7511,N_7235);
nand U7775 (N_7775,N_7532,N_7397);
nor U7776 (N_7776,N_7273,N_7396);
nor U7777 (N_7777,N_7267,N_7445);
nor U7778 (N_7778,N_7489,N_7203);
nor U7779 (N_7779,N_7230,N_7496);
nand U7780 (N_7780,N_7256,N_7392);
nand U7781 (N_7781,N_7556,N_7299);
nor U7782 (N_7782,N_7410,N_7479);
nor U7783 (N_7783,N_7555,N_7374);
nor U7784 (N_7784,N_7272,N_7501);
and U7785 (N_7785,N_7416,N_7542);
nor U7786 (N_7786,N_7457,N_7325);
xnor U7787 (N_7787,N_7528,N_7356);
and U7788 (N_7788,N_7448,N_7562);
xnor U7789 (N_7789,N_7352,N_7317);
or U7790 (N_7790,N_7242,N_7354);
nor U7791 (N_7791,N_7565,N_7234);
and U7792 (N_7792,N_7401,N_7598);
xor U7793 (N_7793,N_7567,N_7568);
or U7794 (N_7794,N_7209,N_7200);
or U7795 (N_7795,N_7216,N_7229);
and U7796 (N_7796,N_7551,N_7284);
xnor U7797 (N_7797,N_7226,N_7526);
nand U7798 (N_7798,N_7332,N_7276);
or U7799 (N_7799,N_7418,N_7434);
or U7800 (N_7800,N_7472,N_7274);
nor U7801 (N_7801,N_7243,N_7323);
and U7802 (N_7802,N_7423,N_7349);
and U7803 (N_7803,N_7522,N_7209);
or U7804 (N_7804,N_7291,N_7516);
and U7805 (N_7805,N_7209,N_7397);
and U7806 (N_7806,N_7217,N_7548);
nor U7807 (N_7807,N_7490,N_7539);
or U7808 (N_7808,N_7223,N_7250);
xnor U7809 (N_7809,N_7249,N_7366);
or U7810 (N_7810,N_7395,N_7233);
xnor U7811 (N_7811,N_7440,N_7222);
and U7812 (N_7812,N_7551,N_7312);
xnor U7813 (N_7813,N_7280,N_7289);
nand U7814 (N_7814,N_7288,N_7478);
or U7815 (N_7815,N_7502,N_7411);
xor U7816 (N_7816,N_7580,N_7317);
xnor U7817 (N_7817,N_7579,N_7508);
nand U7818 (N_7818,N_7422,N_7213);
or U7819 (N_7819,N_7350,N_7534);
nand U7820 (N_7820,N_7220,N_7560);
xor U7821 (N_7821,N_7379,N_7414);
nor U7822 (N_7822,N_7550,N_7512);
or U7823 (N_7823,N_7395,N_7202);
xnor U7824 (N_7824,N_7429,N_7292);
nand U7825 (N_7825,N_7544,N_7483);
or U7826 (N_7826,N_7469,N_7566);
xor U7827 (N_7827,N_7375,N_7439);
and U7828 (N_7828,N_7264,N_7366);
nand U7829 (N_7829,N_7566,N_7251);
xnor U7830 (N_7830,N_7384,N_7457);
nand U7831 (N_7831,N_7547,N_7421);
nand U7832 (N_7832,N_7504,N_7417);
nor U7833 (N_7833,N_7376,N_7265);
or U7834 (N_7834,N_7269,N_7542);
nor U7835 (N_7835,N_7502,N_7406);
xor U7836 (N_7836,N_7415,N_7368);
nor U7837 (N_7837,N_7563,N_7485);
nor U7838 (N_7838,N_7382,N_7245);
xnor U7839 (N_7839,N_7504,N_7531);
nand U7840 (N_7840,N_7345,N_7553);
nor U7841 (N_7841,N_7366,N_7325);
nand U7842 (N_7842,N_7204,N_7252);
or U7843 (N_7843,N_7388,N_7372);
nor U7844 (N_7844,N_7457,N_7399);
nor U7845 (N_7845,N_7434,N_7363);
xnor U7846 (N_7846,N_7408,N_7267);
and U7847 (N_7847,N_7455,N_7431);
nor U7848 (N_7848,N_7505,N_7402);
or U7849 (N_7849,N_7313,N_7544);
nor U7850 (N_7850,N_7340,N_7586);
xnor U7851 (N_7851,N_7462,N_7445);
xnor U7852 (N_7852,N_7561,N_7235);
nand U7853 (N_7853,N_7569,N_7496);
nand U7854 (N_7854,N_7559,N_7568);
or U7855 (N_7855,N_7590,N_7291);
or U7856 (N_7856,N_7200,N_7422);
nor U7857 (N_7857,N_7513,N_7510);
nor U7858 (N_7858,N_7212,N_7506);
or U7859 (N_7859,N_7368,N_7512);
nand U7860 (N_7860,N_7589,N_7281);
nor U7861 (N_7861,N_7523,N_7582);
nand U7862 (N_7862,N_7580,N_7294);
nand U7863 (N_7863,N_7276,N_7362);
nor U7864 (N_7864,N_7236,N_7452);
or U7865 (N_7865,N_7429,N_7538);
xor U7866 (N_7866,N_7559,N_7313);
and U7867 (N_7867,N_7437,N_7330);
nand U7868 (N_7868,N_7351,N_7536);
xnor U7869 (N_7869,N_7410,N_7594);
xnor U7870 (N_7870,N_7479,N_7428);
nand U7871 (N_7871,N_7394,N_7321);
and U7872 (N_7872,N_7570,N_7400);
nand U7873 (N_7873,N_7281,N_7397);
or U7874 (N_7874,N_7290,N_7587);
nor U7875 (N_7875,N_7337,N_7487);
and U7876 (N_7876,N_7504,N_7358);
and U7877 (N_7877,N_7385,N_7548);
or U7878 (N_7878,N_7377,N_7235);
xor U7879 (N_7879,N_7425,N_7314);
nand U7880 (N_7880,N_7469,N_7543);
and U7881 (N_7881,N_7294,N_7419);
nor U7882 (N_7882,N_7516,N_7286);
nor U7883 (N_7883,N_7582,N_7347);
xor U7884 (N_7884,N_7214,N_7546);
and U7885 (N_7885,N_7307,N_7346);
nor U7886 (N_7886,N_7561,N_7525);
nor U7887 (N_7887,N_7387,N_7490);
or U7888 (N_7888,N_7381,N_7226);
and U7889 (N_7889,N_7465,N_7315);
nand U7890 (N_7890,N_7262,N_7288);
and U7891 (N_7891,N_7432,N_7467);
or U7892 (N_7892,N_7484,N_7466);
and U7893 (N_7893,N_7577,N_7517);
nor U7894 (N_7894,N_7257,N_7462);
nor U7895 (N_7895,N_7328,N_7325);
nor U7896 (N_7896,N_7387,N_7208);
and U7897 (N_7897,N_7473,N_7556);
or U7898 (N_7898,N_7263,N_7222);
nor U7899 (N_7899,N_7201,N_7521);
or U7900 (N_7900,N_7304,N_7225);
or U7901 (N_7901,N_7495,N_7468);
or U7902 (N_7902,N_7485,N_7502);
or U7903 (N_7903,N_7552,N_7426);
nand U7904 (N_7904,N_7491,N_7499);
nor U7905 (N_7905,N_7367,N_7575);
and U7906 (N_7906,N_7203,N_7320);
xnor U7907 (N_7907,N_7504,N_7497);
nand U7908 (N_7908,N_7377,N_7524);
xor U7909 (N_7909,N_7488,N_7462);
and U7910 (N_7910,N_7322,N_7471);
xnor U7911 (N_7911,N_7598,N_7586);
nand U7912 (N_7912,N_7242,N_7209);
and U7913 (N_7913,N_7459,N_7400);
nand U7914 (N_7914,N_7580,N_7405);
xor U7915 (N_7915,N_7466,N_7559);
nor U7916 (N_7916,N_7468,N_7504);
and U7917 (N_7917,N_7438,N_7251);
nand U7918 (N_7918,N_7313,N_7395);
or U7919 (N_7919,N_7539,N_7211);
xor U7920 (N_7920,N_7356,N_7354);
xor U7921 (N_7921,N_7292,N_7497);
and U7922 (N_7922,N_7345,N_7245);
and U7923 (N_7923,N_7510,N_7519);
or U7924 (N_7924,N_7277,N_7400);
xnor U7925 (N_7925,N_7470,N_7428);
and U7926 (N_7926,N_7309,N_7297);
xnor U7927 (N_7927,N_7485,N_7389);
nor U7928 (N_7928,N_7210,N_7463);
xor U7929 (N_7929,N_7265,N_7505);
and U7930 (N_7930,N_7345,N_7318);
and U7931 (N_7931,N_7316,N_7377);
xor U7932 (N_7932,N_7417,N_7439);
xor U7933 (N_7933,N_7515,N_7242);
and U7934 (N_7934,N_7346,N_7251);
xor U7935 (N_7935,N_7350,N_7557);
or U7936 (N_7936,N_7524,N_7490);
nor U7937 (N_7937,N_7420,N_7583);
nor U7938 (N_7938,N_7558,N_7597);
and U7939 (N_7939,N_7294,N_7261);
xnor U7940 (N_7940,N_7367,N_7528);
or U7941 (N_7941,N_7493,N_7409);
and U7942 (N_7942,N_7250,N_7231);
or U7943 (N_7943,N_7489,N_7316);
nand U7944 (N_7944,N_7364,N_7518);
or U7945 (N_7945,N_7214,N_7267);
nand U7946 (N_7946,N_7365,N_7245);
nand U7947 (N_7947,N_7492,N_7537);
or U7948 (N_7948,N_7311,N_7245);
and U7949 (N_7949,N_7439,N_7588);
nor U7950 (N_7950,N_7490,N_7356);
and U7951 (N_7951,N_7508,N_7254);
nand U7952 (N_7952,N_7393,N_7571);
nand U7953 (N_7953,N_7253,N_7497);
or U7954 (N_7954,N_7578,N_7501);
nand U7955 (N_7955,N_7508,N_7390);
or U7956 (N_7956,N_7308,N_7527);
or U7957 (N_7957,N_7377,N_7545);
nor U7958 (N_7958,N_7465,N_7270);
nor U7959 (N_7959,N_7575,N_7431);
nand U7960 (N_7960,N_7519,N_7544);
and U7961 (N_7961,N_7529,N_7517);
nor U7962 (N_7962,N_7311,N_7483);
nand U7963 (N_7963,N_7355,N_7593);
and U7964 (N_7964,N_7368,N_7215);
nand U7965 (N_7965,N_7404,N_7537);
and U7966 (N_7966,N_7308,N_7484);
nand U7967 (N_7967,N_7598,N_7284);
xnor U7968 (N_7968,N_7372,N_7287);
or U7969 (N_7969,N_7372,N_7221);
nor U7970 (N_7970,N_7208,N_7599);
or U7971 (N_7971,N_7484,N_7350);
or U7972 (N_7972,N_7586,N_7475);
and U7973 (N_7973,N_7368,N_7479);
nand U7974 (N_7974,N_7211,N_7215);
nand U7975 (N_7975,N_7333,N_7428);
xor U7976 (N_7976,N_7372,N_7535);
or U7977 (N_7977,N_7554,N_7549);
and U7978 (N_7978,N_7304,N_7444);
nor U7979 (N_7979,N_7282,N_7588);
xnor U7980 (N_7980,N_7385,N_7541);
or U7981 (N_7981,N_7253,N_7207);
and U7982 (N_7982,N_7581,N_7559);
xor U7983 (N_7983,N_7239,N_7346);
and U7984 (N_7984,N_7309,N_7400);
and U7985 (N_7985,N_7382,N_7296);
and U7986 (N_7986,N_7328,N_7568);
nand U7987 (N_7987,N_7577,N_7200);
or U7988 (N_7988,N_7301,N_7540);
and U7989 (N_7989,N_7544,N_7422);
nor U7990 (N_7990,N_7491,N_7264);
nor U7991 (N_7991,N_7270,N_7415);
and U7992 (N_7992,N_7323,N_7211);
xor U7993 (N_7993,N_7431,N_7501);
or U7994 (N_7994,N_7258,N_7230);
and U7995 (N_7995,N_7437,N_7243);
nand U7996 (N_7996,N_7332,N_7223);
nor U7997 (N_7997,N_7452,N_7444);
nand U7998 (N_7998,N_7271,N_7522);
or U7999 (N_7999,N_7301,N_7444);
nor U8000 (N_8000,N_7619,N_7810);
xnor U8001 (N_8001,N_7747,N_7988);
nand U8002 (N_8002,N_7622,N_7891);
nor U8003 (N_8003,N_7749,N_7805);
and U8004 (N_8004,N_7944,N_7853);
nand U8005 (N_8005,N_7842,N_7672);
nand U8006 (N_8006,N_7857,N_7973);
and U8007 (N_8007,N_7893,N_7949);
xor U8008 (N_8008,N_7728,N_7795);
nand U8009 (N_8009,N_7665,N_7854);
and U8010 (N_8010,N_7982,N_7678);
nor U8011 (N_8011,N_7715,N_7647);
nor U8012 (N_8012,N_7675,N_7606);
and U8013 (N_8013,N_7624,N_7866);
or U8014 (N_8014,N_7929,N_7762);
or U8015 (N_8015,N_7629,N_7708);
nor U8016 (N_8016,N_7938,N_7714);
xnor U8017 (N_8017,N_7947,N_7964);
or U8018 (N_8018,N_7943,N_7711);
nor U8019 (N_8019,N_7630,N_7743);
nor U8020 (N_8020,N_7803,N_7661);
or U8021 (N_8021,N_7781,N_7843);
nor U8022 (N_8022,N_7981,N_7607);
and U8023 (N_8023,N_7787,N_7908);
nand U8024 (N_8024,N_7816,N_7693);
or U8025 (N_8025,N_7636,N_7821);
or U8026 (N_8026,N_7748,N_7741);
and U8027 (N_8027,N_7727,N_7890);
or U8028 (N_8028,N_7742,N_7756);
nor U8029 (N_8029,N_7990,N_7862);
nand U8030 (N_8030,N_7915,N_7831);
or U8031 (N_8031,N_7820,N_7774);
or U8032 (N_8032,N_7924,N_7861);
xnor U8033 (N_8033,N_7783,N_7840);
xnor U8034 (N_8034,N_7836,N_7977);
xnor U8035 (N_8035,N_7666,N_7823);
nor U8036 (N_8036,N_7677,N_7645);
nor U8037 (N_8037,N_7612,N_7737);
and U8038 (N_8038,N_7919,N_7962);
xnor U8039 (N_8039,N_7791,N_7855);
nor U8040 (N_8040,N_7818,N_7758);
xnor U8041 (N_8041,N_7621,N_7692);
nand U8042 (N_8042,N_7730,N_7641);
or U8043 (N_8043,N_7697,N_7927);
nand U8044 (N_8044,N_7860,N_7999);
nand U8045 (N_8045,N_7910,N_7784);
and U8046 (N_8046,N_7948,N_7685);
nor U8047 (N_8047,N_7957,N_7751);
xor U8048 (N_8048,N_7614,N_7682);
xnor U8049 (N_8049,N_7766,N_7884);
or U8050 (N_8050,N_7811,N_7750);
nor U8051 (N_8051,N_7625,N_7768);
nor U8052 (N_8052,N_7709,N_7807);
nand U8053 (N_8053,N_7732,N_7705);
and U8054 (N_8054,N_7892,N_7806);
and U8055 (N_8055,N_7663,N_7907);
and U8056 (N_8056,N_7826,N_7897);
nand U8057 (N_8057,N_7965,N_7912);
nor U8058 (N_8058,N_7902,N_7695);
nor U8059 (N_8059,N_7968,N_7996);
nand U8060 (N_8060,N_7955,N_7769);
nand U8061 (N_8061,N_7946,N_7710);
nand U8062 (N_8062,N_7640,N_7833);
nor U8063 (N_8063,N_7754,N_7909);
xnor U8064 (N_8064,N_7802,N_7984);
nand U8065 (N_8065,N_7918,N_7815);
nor U8066 (N_8066,N_7713,N_7793);
and U8067 (N_8067,N_7706,N_7753);
or U8068 (N_8068,N_7601,N_7778);
and U8069 (N_8069,N_7814,N_7679);
nand U8070 (N_8070,N_7650,N_7755);
or U8071 (N_8071,N_7765,N_7933);
nor U8072 (N_8072,N_7790,N_7696);
and U8073 (N_8073,N_7637,N_7864);
nand U8074 (N_8074,N_7772,N_7789);
and U8075 (N_8075,N_7786,N_7992);
nand U8076 (N_8076,N_7746,N_7617);
or U8077 (N_8077,N_7659,N_7722);
xor U8078 (N_8078,N_7669,N_7881);
nand U8079 (N_8079,N_7654,N_7998);
or U8080 (N_8080,N_7880,N_7978);
or U8081 (N_8081,N_7940,N_7983);
or U8082 (N_8082,N_7604,N_7960);
nand U8083 (N_8083,N_7782,N_7761);
and U8084 (N_8084,N_7963,N_7951);
and U8085 (N_8085,N_7870,N_7632);
xnor U8086 (N_8086,N_7917,N_7904);
and U8087 (N_8087,N_7937,N_7877);
xnor U8088 (N_8088,N_7703,N_7876);
and U8089 (N_8089,N_7676,N_7898);
and U8090 (N_8090,N_7856,N_7792);
nand U8091 (N_8091,N_7633,N_7626);
or U8092 (N_8092,N_7616,N_7740);
or U8093 (N_8093,N_7812,N_7941);
nor U8094 (N_8094,N_7648,N_7716);
nand U8095 (N_8095,N_7916,N_7886);
nor U8096 (N_8096,N_7776,N_7667);
xor U8097 (N_8097,N_7660,N_7800);
xnor U8098 (N_8098,N_7674,N_7829);
nor U8099 (N_8099,N_7899,N_7993);
and U8100 (N_8100,N_7888,N_7689);
nor U8101 (N_8101,N_7618,N_7687);
nor U8102 (N_8102,N_7627,N_7723);
and U8103 (N_8103,N_7851,N_7798);
xnor U8104 (N_8104,N_7731,N_7980);
or U8105 (N_8105,N_7688,N_7920);
nand U8106 (N_8106,N_7738,N_7615);
and U8107 (N_8107,N_7869,N_7773);
nor U8108 (N_8108,N_7651,N_7808);
nor U8109 (N_8109,N_7871,N_7817);
nor U8110 (N_8110,N_7691,N_7889);
or U8111 (N_8111,N_7958,N_7736);
nor U8112 (N_8112,N_7646,N_7923);
xnor U8113 (N_8113,N_7926,N_7700);
and U8114 (N_8114,N_7610,N_7875);
and U8115 (N_8115,N_7763,N_7914);
or U8116 (N_8116,N_7739,N_7865);
xor U8117 (N_8117,N_7956,N_7759);
and U8118 (N_8118,N_7704,N_7882);
and U8119 (N_8119,N_7837,N_7702);
xor U8120 (N_8120,N_7945,N_7994);
nor U8121 (N_8121,N_7987,N_7760);
nor U8122 (N_8122,N_7989,N_7922);
nor U8123 (N_8123,N_7844,N_7794);
nor U8124 (N_8124,N_7657,N_7699);
and U8125 (N_8125,N_7906,N_7879);
nand U8126 (N_8126,N_7780,N_7639);
nand U8127 (N_8127,N_7901,N_7824);
or U8128 (N_8128,N_7967,N_7850);
nor U8129 (N_8129,N_7863,N_7995);
nor U8130 (N_8130,N_7690,N_7975);
xnor U8131 (N_8131,N_7859,N_7670);
nor U8132 (N_8132,N_7724,N_7734);
nand U8133 (N_8133,N_7848,N_7858);
or U8134 (N_8134,N_7623,N_7628);
xnor U8135 (N_8135,N_7834,N_7698);
nor U8136 (N_8136,N_7717,N_7830);
nor U8137 (N_8137,N_7643,N_7775);
nand U8138 (N_8138,N_7936,N_7652);
and U8139 (N_8139,N_7894,N_7720);
nor U8140 (N_8140,N_7744,N_7770);
and U8141 (N_8141,N_7966,N_7673);
nor U8142 (N_8142,N_7976,N_7779);
nand U8143 (N_8143,N_7868,N_7991);
and U8144 (N_8144,N_7997,N_7935);
xnor U8145 (N_8145,N_7939,N_7683);
nor U8146 (N_8146,N_7928,N_7913);
or U8147 (N_8147,N_7712,N_7986);
nand U8148 (N_8148,N_7934,N_7900);
and U8149 (N_8149,N_7681,N_7600);
and U8150 (N_8150,N_7671,N_7735);
nor U8151 (N_8151,N_7942,N_7804);
nand U8152 (N_8152,N_7930,N_7719);
or U8153 (N_8153,N_7668,N_7801);
xnor U8154 (N_8154,N_7635,N_7777);
and U8155 (N_8155,N_7733,N_7839);
xnor U8156 (N_8156,N_7608,N_7903);
xor U8157 (N_8157,N_7785,N_7662);
nand U8158 (N_8158,N_7985,N_7603);
nor U8159 (N_8159,N_7883,N_7634);
nand U8160 (N_8160,N_7655,N_7847);
or U8161 (N_8161,N_7680,N_7819);
nor U8162 (N_8162,N_7950,N_7664);
xor U8163 (N_8163,N_7809,N_7873);
nand U8164 (N_8164,N_7796,N_7799);
or U8165 (N_8165,N_7961,N_7813);
xor U8166 (N_8166,N_7620,N_7684);
or U8167 (N_8167,N_7925,N_7788);
nor U8168 (N_8168,N_7885,N_7718);
nand U8169 (N_8169,N_7974,N_7845);
nand U8170 (N_8170,N_7707,N_7931);
nor U8171 (N_8171,N_7686,N_7729);
xor U8172 (N_8172,N_7642,N_7832);
or U8173 (N_8173,N_7921,N_7822);
or U8174 (N_8174,N_7835,N_7952);
or U8175 (N_8175,N_7721,N_7605);
and U8176 (N_8176,N_7649,N_7609);
nand U8177 (N_8177,N_7849,N_7771);
or U8178 (N_8178,N_7896,N_7752);
or U8179 (N_8179,N_7828,N_7725);
xnor U8180 (N_8180,N_7767,N_7979);
or U8181 (N_8181,N_7701,N_7694);
nand U8182 (N_8182,N_7797,N_7841);
or U8183 (N_8183,N_7611,N_7932);
and U8184 (N_8184,N_7745,N_7631);
or U8185 (N_8185,N_7644,N_7638);
nand U8186 (N_8186,N_7971,N_7827);
nor U8187 (N_8187,N_7895,N_7653);
or U8188 (N_8188,N_7846,N_7959);
or U8189 (N_8189,N_7656,N_7726);
xnor U8190 (N_8190,N_7764,N_7613);
nor U8191 (N_8191,N_7838,N_7905);
and U8192 (N_8192,N_7872,N_7874);
or U8193 (N_8193,N_7658,N_7602);
nand U8194 (N_8194,N_7972,N_7954);
nand U8195 (N_8195,N_7887,N_7953);
xnor U8196 (N_8196,N_7911,N_7970);
nand U8197 (N_8197,N_7757,N_7867);
xor U8198 (N_8198,N_7825,N_7969);
and U8199 (N_8199,N_7852,N_7878);
and U8200 (N_8200,N_7651,N_7652);
nand U8201 (N_8201,N_7971,N_7931);
and U8202 (N_8202,N_7998,N_7766);
xor U8203 (N_8203,N_7774,N_7842);
xnor U8204 (N_8204,N_7868,N_7892);
nand U8205 (N_8205,N_7802,N_7665);
xnor U8206 (N_8206,N_7618,N_7938);
or U8207 (N_8207,N_7859,N_7601);
xor U8208 (N_8208,N_7607,N_7881);
and U8209 (N_8209,N_7873,N_7638);
or U8210 (N_8210,N_7972,N_7835);
or U8211 (N_8211,N_7708,N_7647);
nand U8212 (N_8212,N_7746,N_7772);
nand U8213 (N_8213,N_7701,N_7685);
nand U8214 (N_8214,N_7988,N_7949);
nand U8215 (N_8215,N_7625,N_7943);
nor U8216 (N_8216,N_7762,N_7777);
or U8217 (N_8217,N_7896,N_7857);
nand U8218 (N_8218,N_7757,N_7901);
nand U8219 (N_8219,N_7678,N_7918);
xnor U8220 (N_8220,N_7616,N_7678);
and U8221 (N_8221,N_7975,N_7681);
or U8222 (N_8222,N_7735,N_7603);
nor U8223 (N_8223,N_7807,N_7968);
xnor U8224 (N_8224,N_7962,N_7952);
nand U8225 (N_8225,N_7943,N_7829);
or U8226 (N_8226,N_7858,N_7825);
nand U8227 (N_8227,N_7640,N_7758);
nor U8228 (N_8228,N_7750,N_7746);
xnor U8229 (N_8229,N_7843,N_7741);
nand U8230 (N_8230,N_7724,N_7892);
and U8231 (N_8231,N_7707,N_7775);
nand U8232 (N_8232,N_7881,N_7645);
nand U8233 (N_8233,N_7615,N_7963);
nand U8234 (N_8234,N_7927,N_7797);
and U8235 (N_8235,N_7600,N_7811);
nand U8236 (N_8236,N_7873,N_7868);
or U8237 (N_8237,N_7628,N_7928);
or U8238 (N_8238,N_7965,N_7665);
or U8239 (N_8239,N_7945,N_7873);
nor U8240 (N_8240,N_7975,N_7809);
and U8241 (N_8241,N_7923,N_7746);
nor U8242 (N_8242,N_7782,N_7714);
xor U8243 (N_8243,N_7839,N_7989);
nor U8244 (N_8244,N_7641,N_7783);
nand U8245 (N_8245,N_7625,N_7743);
xnor U8246 (N_8246,N_7805,N_7889);
or U8247 (N_8247,N_7976,N_7826);
and U8248 (N_8248,N_7991,N_7851);
nor U8249 (N_8249,N_7899,N_7734);
xnor U8250 (N_8250,N_7944,N_7727);
nand U8251 (N_8251,N_7991,N_7914);
or U8252 (N_8252,N_7720,N_7997);
and U8253 (N_8253,N_7889,N_7897);
or U8254 (N_8254,N_7699,N_7782);
nor U8255 (N_8255,N_7773,N_7969);
nand U8256 (N_8256,N_7999,N_7676);
nand U8257 (N_8257,N_7904,N_7741);
nor U8258 (N_8258,N_7685,N_7825);
xnor U8259 (N_8259,N_7877,N_7802);
nand U8260 (N_8260,N_7764,N_7812);
or U8261 (N_8261,N_7751,N_7762);
or U8262 (N_8262,N_7955,N_7715);
xnor U8263 (N_8263,N_7789,N_7767);
xnor U8264 (N_8264,N_7887,N_7917);
nand U8265 (N_8265,N_7980,N_7667);
nand U8266 (N_8266,N_7627,N_7609);
nand U8267 (N_8267,N_7602,N_7889);
xor U8268 (N_8268,N_7988,N_7873);
or U8269 (N_8269,N_7634,N_7687);
or U8270 (N_8270,N_7842,N_7643);
nor U8271 (N_8271,N_7936,N_7657);
nor U8272 (N_8272,N_7684,N_7757);
xnor U8273 (N_8273,N_7795,N_7639);
or U8274 (N_8274,N_7692,N_7940);
nand U8275 (N_8275,N_7611,N_7947);
and U8276 (N_8276,N_7662,N_7753);
xnor U8277 (N_8277,N_7900,N_7834);
nor U8278 (N_8278,N_7795,N_7785);
nor U8279 (N_8279,N_7947,N_7662);
nand U8280 (N_8280,N_7768,N_7871);
nand U8281 (N_8281,N_7962,N_7881);
or U8282 (N_8282,N_7920,N_7687);
or U8283 (N_8283,N_7635,N_7855);
xor U8284 (N_8284,N_7752,N_7735);
or U8285 (N_8285,N_7992,N_7823);
nand U8286 (N_8286,N_7766,N_7634);
nor U8287 (N_8287,N_7922,N_7909);
nor U8288 (N_8288,N_7686,N_7675);
nand U8289 (N_8289,N_7621,N_7901);
nor U8290 (N_8290,N_7694,N_7945);
or U8291 (N_8291,N_7623,N_7797);
and U8292 (N_8292,N_7660,N_7688);
nor U8293 (N_8293,N_7670,N_7738);
or U8294 (N_8294,N_7835,N_7615);
xnor U8295 (N_8295,N_7715,N_7605);
xnor U8296 (N_8296,N_7837,N_7882);
and U8297 (N_8297,N_7653,N_7908);
or U8298 (N_8298,N_7616,N_7635);
nand U8299 (N_8299,N_7679,N_7651);
nand U8300 (N_8300,N_7999,N_7850);
and U8301 (N_8301,N_7632,N_7814);
or U8302 (N_8302,N_7673,N_7615);
xnor U8303 (N_8303,N_7748,N_7995);
or U8304 (N_8304,N_7634,N_7824);
or U8305 (N_8305,N_7848,N_7703);
or U8306 (N_8306,N_7845,N_7846);
nor U8307 (N_8307,N_7691,N_7620);
or U8308 (N_8308,N_7725,N_7605);
nand U8309 (N_8309,N_7953,N_7606);
and U8310 (N_8310,N_7936,N_7682);
nor U8311 (N_8311,N_7864,N_7760);
nor U8312 (N_8312,N_7891,N_7971);
and U8313 (N_8313,N_7721,N_7700);
nand U8314 (N_8314,N_7821,N_7793);
or U8315 (N_8315,N_7652,N_7780);
nand U8316 (N_8316,N_7883,N_7973);
and U8317 (N_8317,N_7710,N_7936);
xor U8318 (N_8318,N_7780,N_7625);
or U8319 (N_8319,N_7692,N_7701);
and U8320 (N_8320,N_7621,N_7770);
and U8321 (N_8321,N_7681,N_7716);
or U8322 (N_8322,N_7695,N_7898);
xnor U8323 (N_8323,N_7621,N_7780);
xnor U8324 (N_8324,N_7622,N_7672);
and U8325 (N_8325,N_7945,N_7619);
and U8326 (N_8326,N_7671,N_7795);
or U8327 (N_8327,N_7745,N_7689);
or U8328 (N_8328,N_7960,N_7691);
and U8329 (N_8329,N_7874,N_7663);
nor U8330 (N_8330,N_7956,N_7846);
xnor U8331 (N_8331,N_7981,N_7833);
or U8332 (N_8332,N_7813,N_7680);
or U8333 (N_8333,N_7681,N_7929);
xor U8334 (N_8334,N_7871,N_7730);
nor U8335 (N_8335,N_7923,N_7632);
nand U8336 (N_8336,N_7851,N_7987);
and U8337 (N_8337,N_7881,N_7782);
nor U8338 (N_8338,N_7666,N_7968);
and U8339 (N_8339,N_7977,N_7654);
and U8340 (N_8340,N_7822,N_7693);
xor U8341 (N_8341,N_7715,N_7870);
xnor U8342 (N_8342,N_7742,N_7905);
xnor U8343 (N_8343,N_7817,N_7803);
nor U8344 (N_8344,N_7669,N_7837);
or U8345 (N_8345,N_7686,N_7776);
nor U8346 (N_8346,N_7886,N_7896);
or U8347 (N_8347,N_7794,N_7808);
or U8348 (N_8348,N_7872,N_7927);
xnor U8349 (N_8349,N_7965,N_7806);
or U8350 (N_8350,N_7874,N_7845);
nand U8351 (N_8351,N_7765,N_7927);
nand U8352 (N_8352,N_7887,N_7980);
nand U8353 (N_8353,N_7970,N_7857);
or U8354 (N_8354,N_7719,N_7902);
nand U8355 (N_8355,N_7840,N_7630);
or U8356 (N_8356,N_7616,N_7949);
nor U8357 (N_8357,N_7629,N_7613);
or U8358 (N_8358,N_7906,N_7893);
xor U8359 (N_8359,N_7986,N_7646);
or U8360 (N_8360,N_7783,N_7863);
nand U8361 (N_8361,N_7767,N_7771);
and U8362 (N_8362,N_7875,N_7787);
or U8363 (N_8363,N_7823,N_7936);
or U8364 (N_8364,N_7983,N_7684);
or U8365 (N_8365,N_7626,N_7704);
nand U8366 (N_8366,N_7890,N_7813);
nand U8367 (N_8367,N_7862,N_7657);
or U8368 (N_8368,N_7707,N_7695);
nand U8369 (N_8369,N_7782,N_7855);
nor U8370 (N_8370,N_7777,N_7876);
nand U8371 (N_8371,N_7976,N_7893);
nand U8372 (N_8372,N_7918,N_7653);
and U8373 (N_8373,N_7972,N_7763);
nand U8374 (N_8374,N_7944,N_7687);
nor U8375 (N_8375,N_7924,N_7982);
nor U8376 (N_8376,N_7769,N_7967);
nand U8377 (N_8377,N_7928,N_7657);
nand U8378 (N_8378,N_7687,N_7813);
nor U8379 (N_8379,N_7992,N_7807);
nor U8380 (N_8380,N_7648,N_7611);
nor U8381 (N_8381,N_7677,N_7994);
nor U8382 (N_8382,N_7761,N_7622);
or U8383 (N_8383,N_7749,N_7835);
or U8384 (N_8384,N_7933,N_7901);
xor U8385 (N_8385,N_7921,N_7630);
nand U8386 (N_8386,N_7637,N_7655);
and U8387 (N_8387,N_7790,N_7984);
nor U8388 (N_8388,N_7936,N_7642);
nand U8389 (N_8389,N_7950,N_7969);
nand U8390 (N_8390,N_7867,N_7759);
nand U8391 (N_8391,N_7806,N_7674);
or U8392 (N_8392,N_7666,N_7601);
nand U8393 (N_8393,N_7710,N_7778);
and U8394 (N_8394,N_7742,N_7724);
xor U8395 (N_8395,N_7760,N_7829);
xnor U8396 (N_8396,N_7707,N_7700);
xnor U8397 (N_8397,N_7808,N_7993);
nand U8398 (N_8398,N_7729,N_7906);
nand U8399 (N_8399,N_7846,N_7686);
and U8400 (N_8400,N_8022,N_8187);
and U8401 (N_8401,N_8211,N_8209);
nand U8402 (N_8402,N_8267,N_8043);
nand U8403 (N_8403,N_8192,N_8333);
xor U8404 (N_8404,N_8232,N_8205);
and U8405 (N_8405,N_8372,N_8195);
or U8406 (N_8406,N_8093,N_8253);
nor U8407 (N_8407,N_8106,N_8304);
nor U8408 (N_8408,N_8008,N_8386);
nand U8409 (N_8409,N_8114,N_8025);
xnor U8410 (N_8410,N_8342,N_8256);
nor U8411 (N_8411,N_8111,N_8283);
nor U8412 (N_8412,N_8203,N_8359);
and U8413 (N_8413,N_8103,N_8049);
and U8414 (N_8414,N_8084,N_8269);
nor U8415 (N_8415,N_8235,N_8229);
or U8416 (N_8416,N_8319,N_8223);
xor U8417 (N_8417,N_8107,N_8110);
nor U8418 (N_8418,N_8099,N_8073);
and U8419 (N_8419,N_8344,N_8214);
or U8420 (N_8420,N_8348,N_8115);
xnor U8421 (N_8421,N_8332,N_8071);
or U8422 (N_8422,N_8280,N_8362);
nor U8423 (N_8423,N_8350,N_8385);
xnor U8424 (N_8424,N_8265,N_8054);
or U8425 (N_8425,N_8293,N_8230);
nor U8426 (N_8426,N_8009,N_8397);
xnor U8427 (N_8427,N_8081,N_8351);
nor U8428 (N_8428,N_8378,N_8045);
xnor U8429 (N_8429,N_8289,N_8090);
or U8430 (N_8430,N_8311,N_8198);
nor U8431 (N_8431,N_8142,N_8023);
nor U8432 (N_8432,N_8322,N_8382);
xor U8433 (N_8433,N_8001,N_8094);
nor U8434 (N_8434,N_8347,N_8238);
or U8435 (N_8435,N_8302,N_8301);
xnor U8436 (N_8436,N_8029,N_8307);
nor U8437 (N_8437,N_8006,N_8150);
or U8438 (N_8438,N_8053,N_8363);
nand U8439 (N_8439,N_8066,N_8276);
nand U8440 (N_8440,N_8091,N_8051);
or U8441 (N_8441,N_8037,N_8279);
nor U8442 (N_8442,N_8296,N_8297);
xnor U8443 (N_8443,N_8287,N_8180);
xnor U8444 (N_8444,N_8288,N_8096);
xor U8445 (N_8445,N_8075,N_8095);
nor U8446 (N_8446,N_8349,N_8334);
and U8447 (N_8447,N_8146,N_8018);
xnor U8448 (N_8448,N_8394,N_8373);
nor U8449 (N_8449,N_8316,N_8318);
nand U8450 (N_8450,N_8182,N_8219);
xor U8451 (N_8451,N_8188,N_8181);
xnor U8452 (N_8452,N_8005,N_8167);
nor U8453 (N_8453,N_8346,N_8149);
nand U8454 (N_8454,N_8021,N_8343);
and U8455 (N_8455,N_8245,N_8092);
and U8456 (N_8456,N_8208,N_8225);
or U8457 (N_8457,N_8166,N_8077);
nand U8458 (N_8458,N_8174,N_8058);
and U8459 (N_8459,N_8263,N_8104);
xnor U8460 (N_8460,N_8340,N_8282);
or U8461 (N_8461,N_8196,N_8159);
nor U8462 (N_8462,N_8113,N_8070);
xnor U8463 (N_8463,N_8171,N_8065);
nand U8464 (N_8464,N_8087,N_8185);
or U8465 (N_8465,N_8014,N_8273);
nor U8466 (N_8466,N_8120,N_8173);
and U8467 (N_8467,N_8312,N_8193);
or U8468 (N_8468,N_8160,N_8170);
or U8469 (N_8469,N_8147,N_8074);
or U8470 (N_8470,N_8278,N_8162);
nand U8471 (N_8471,N_8153,N_8286);
nor U8472 (N_8472,N_8161,N_8124);
nor U8473 (N_8473,N_8299,N_8345);
nand U8474 (N_8474,N_8169,N_8175);
nor U8475 (N_8475,N_8371,N_8375);
or U8476 (N_8476,N_8381,N_8121);
nand U8477 (N_8477,N_8308,N_8038);
xor U8478 (N_8478,N_8064,N_8369);
nand U8479 (N_8479,N_8285,N_8068);
xor U8480 (N_8480,N_8379,N_8341);
and U8481 (N_8481,N_8183,N_8041);
xor U8482 (N_8482,N_8031,N_8030);
nand U8483 (N_8483,N_8112,N_8080);
or U8484 (N_8484,N_8133,N_8295);
nand U8485 (N_8485,N_8251,N_8315);
xnor U8486 (N_8486,N_8108,N_8085);
or U8487 (N_8487,N_8360,N_8317);
xnor U8488 (N_8488,N_8306,N_8339);
and U8489 (N_8489,N_8290,N_8275);
nor U8490 (N_8490,N_8395,N_8059);
and U8491 (N_8491,N_8393,N_8168);
and U8492 (N_8492,N_8044,N_8189);
or U8493 (N_8493,N_8237,N_8067);
or U8494 (N_8494,N_8156,N_8220);
or U8495 (N_8495,N_8199,N_8262);
nand U8496 (N_8496,N_8097,N_8004);
xnor U8497 (N_8497,N_8206,N_8154);
and U8498 (N_8498,N_8165,N_8027);
and U8499 (N_8499,N_8191,N_8274);
nand U8500 (N_8500,N_8047,N_8069);
and U8501 (N_8501,N_8010,N_8258);
nor U8502 (N_8502,N_8144,N_8016);
nor U8503 (N_8503,N_8098,N_8123);
nand U8504 (N_8504,N_8329,N_8143);
nand U8505 (N_8505,N_8015,N_8152);
nor U8506 (N_8506,N_8366,N_8032);
nor U8507 (N_8507,N_8392,N_8186);
nand U8508 (N_8508,N_8358,N_8336);
xor U8509 (N_8509,N_8135,N_8052);
and U8510 (N_8510,N_8013,N_8255);
and U8511 (N_8511,N_8061,N_8204);
nor U8512 (N_8512,N_8079,N_8352);
xor U8513 (N_8513,N_8327,N_8228);
and U8514 (N_8514,N_8056,N_8226);
xor U8515 (N_8515,N_8017,N_8356);
nand U8516 (N_8516,N_8050,N_8261);
xnor U8517 (N_8517,N_8040,N_8270);
or U8518 (N_8518,N_8390,N_8155);
and U8519 (N_8519,N_8011,N_8179);
and U8520 (N_8520,N_8398,N_8158);
xor U8521 (N_8521,N_8042,N_8252);
and U8522 (N_8522,N_8361,N_8151);
xor U8523 (N_8523,N_8063,N_8020);
or U8524 (N_8524,N_8268,N_8239);
nand U8525 (N_8525,N_8355,N_8122);
xnor U8526 (N_8526,N_8046,N_8126);
or U8527 (N_8527,N_8243,N_8326);
and U8528 (N_8528,N_8197,N_8244);
xor U8529 (N_8529,N_8377,N_8222);
nand U8530 (N_8530,N_8164,N_8109);
and U8531 (N_8531,N_8200,N_8086);
or U8532 (N_8532,N_8019,N_8076);
xnor U8533 (N_8533,N_8257,N_8148);
xor U8534 (N_8534,N_8357,N_8088);
or U8535 (N_8535,N_8314,N_8310);
and U8536 (N_8536,N_8254,N_8003);
nor U8537 (N_8537,N_8119,N_8100);
and U8538 (N_8538,N_8082,N_8163);
nor U8539 (N_8539,N_8233,N_8337);
nand U8540 (N_8540,N_8324,N_8368);
nand U8541 (N_8541,N_8141,N_8083);
xnor U8542 (N_8542,N_8383,N_8231);
nor U8543 (N_8543,N_8399,N_8145);
xor U8544 (N_8544,N_8117,N_8241);
or U8545 (N_8545,N_8365,N_8264);
and U8546 (N_8546,N_8242,N_8331);
or U8547 (N_8547,N_8291,N_8136);
nand U8548 (N_8548,N_8260,N_8294);
and U8549 (N_8549,N_8134,N_8328);
and U8550 (N_8550,N_8078,N_8012);
or U8551 (N_8551,N_8137,N_8048);
nand U8552 (N_8552,N_8212,N_8125);
xnor U8553 (N_8553,N_8367,N_8374);
nand U8554 (N_8554,N_8202,N_8028);
and U8555 (N_8555,N_8177,N_8089);
nand U8556 (N_8556,N_8062,N_8236);
xor U8557 (N_8557,N_8323,N_8039);
nor U8558 (N_8558,N_8380,N_8303);
nor U8559 (N_8559,N_8221,N_8213);
nand U8560 (N_8560,N_8139,N_8128);
and U8561 (N_8561,N_8036,N_8246);
or U8562 (N_8562,N_8266,N_8207);
xor U8563 (N_8563,N_8157,N_8194);
nand U8564 (N_8564,N_8292,N_8224);
xnor U8565 (N_8565,N_8210,N_8396);
xnor U8566 (N_8566,N_8178,N_8118);
nand U8567 (N_8567,N_8300,N_8101);
or U8568 (N_8568,N_8000,N_8320);
xor U8569 (N_8569,N_8201,N_8057);
and U8570 (N_8570,N_8272,N_8184);
xnor U8571 (N_8571,N_8354,N_8140);
and U8572 (N_8572,N_8384,N_8387);
and U8573 (N_8573,N_8190,N_8227);
nand U8574 (N_8574,N_8321,N_8007);
nor U8575 (N_8575,N_8072,N_8055);
and U8576 (N_8576,N_8132,N_8364);
nor U8577 (N_8577,N_8138,N_8026);
nand U8578 (N_8578,N_8024,N_8127);
and U8579 (N_8579,N_8131,N_8060);
nand U8580 (N_8580,N_8313,N_8129);
nand U8581 (N_8581,N_8335,N_8172);
nand U8582 (N_8582,N_8249,N_8247);
and U8583 (N_8583,N_8116,N_8002);
nor U8584 (N_8584,N_8216,N_8176);
xor U8585 (N_8585,N_8105,N_8035);
nand U8586 (N_8586,N_8240,N_8391);
nand U8587 (N_8587,N_8389,N_8217);
nand U8588 (N_8588,N_8234,N_8248);
and U8589 (N_8589,N_8271,N_8218);
nor U8590 (N_8590,N_8305,N_8298);
nor U8591 (N_8591,N_8330,N_8376);
xor U8592 (N_8592,N_8215,N_8281);
or U8593 (N_8593,N_8370,N_8259);
nand U8594 (N_8594,N_8130,N_8388);
xor U8595 (N_8595,N_8309,N_8325);
or U8596 (N_8596,N_8277,N_8250);
nor U8597 (N_8597,N_8034,N_8338);
nand U8598 (N_8598,N_8102,N_8033);
or U8599 (N_8599,N_8353,N_8284);
or U8600 (N_8600,N_8221,N_8246);
xor U8601 (N_8601,N_8117,N_8178);
nor U8602 (N_8602,N_8073,N_8043);
and U8603 (N_8603,N_8184,N_8327);
nor U8604 (N_8604,N_8246,N_8266);
xor U8605 (N_8605,N_8054,N_8069);
and U8606 (N_8606,N_8111,N_8128);
nand U8607 (N_8607,N_8147,N_8321);
xnor U8608 (N_8608,N_8084,N_8221);
nor U8609 (N_8609,N_8029,N_8066);
nand U8610 (N_8610,N_8206,N_8172);
or U8611 (N_8611,N_8200,N_8115);
nand U8612 (N_8612,N_8312,N_8367);
xnor U8613 (N_8613,N_8277,N_8343);
and U8614 (N_8614,N_8228,N_8210);
xnor U8615 (N_8615,N_8275,N_8011);
nand U8616 (N_8616,N_8047,N_8188);
and U8617 (N_8617,N_8131,N_8064);
nand U8618 (N_8618,N_8321,N_8094);
nor U8619 (N_8619,N_8326,N_8024);
or U8620 (N_8620,N_8045,N_8214);
nand U8621 (N_8621,N_8022,N_8131);
xnor U8622 (N_8622,N_8200,N_8023);
and U8623 (N_8623,N_8010,N_8349);
nor U8624 (N_8624,N_8154,N_8126);
xor U8625 (N_8625,N_8075,N_8250);
or U8626 (N_8626,N_8193,N_8317);
or U8627 (N_8627,N_8078,N_8395);
xor U8628 (N_8628,N_8021,N_8329);
xnor U8629 (N_8629,N_8219,N_8295);
xor U8630 (N_8630,N_8291,N_8190);
or U8631 (N_8631,N_8254,N_8336);
and U8632 (N_8632,N_8062,N_8354);
nand U8633 (N_8633,N_8064,N_8027);
and U8634 (N_8634,N_8337,N_8013);
and U8635 (N_8635,N_8015,N_8328);
and U8636 (N_8636,N_8173,N_8115);
xnor U8637 (N_8637,N_8252,N_8263);
or U8638 (N_8638,N_8169,N_8145);
or U8639 (N_8639,N_8039,N_8171);
xnor U8640 (N_8640,N_8121,N_8223);
nor U8641 (N_8641,N_8106,N_8249);
and U8642 (N_8642,N_8130,N_8305);
nand U8643 (N_8643,N_8379,N_8268);
nor U8644 (N_8644,N_8297,N_8090);
and U8645 (N_8645,N_8037,N_8241);
nor U8646 (N_8646,N_8206,N_8253);
and U8647 (N_8647,N_8345,N_8045);
nor U8648 (N_8648,N_8038,N_8245);
nor U8649 (N_8649,N_8325,N_8310);
xnor U8650 (N_8650,N_8129,N_8346);
nor U8651 (N_8651,N_8165,N_8158);
or U8652 (N_8652,N_8180,N_8247);
or U8653 (N_8653,N_8390,N_8179);
xnor U8654 (N_8654,N_8214,N_8379);
nand U8655 (N_8655,N_8027,N_8045);
nor U8656 (N_8656,N_8198,N_8381);
and U8657 (N_8657,N_8174,N_8382);
and U8658 (N_8658,N_8001,N_8205);
and U8659 (N_8659,N_8370,N_8330);
xnor U8660 (N_8660,N_8320,N_8260);
xnor U8661 (N_8661,N_8082,N_8070);
or U8662 (N_8662,N_8354,N_8248);
xnor U8663 (N_8663,N_8150,N_8374);
or U8664 (N_8664,N_8351,N_8180);
xnor U8665 (N_8665,N_8349,N_8360);
nor U8666 (N_8666,N_8069,N_8012);
xor U8667 (N_8667,N_8034,N_8309);
and U8668 (N_8668,N_8197,N_8002);
nor U8669 (N_8669,N_8332,N_8003);
nor U8670 (N_8670,N_8104,N_8200);
nor U8671 (N_8671,N_8148,N_8220);
nor U8672 (N_8672,N_8089,N_8319);
nor U8673 (N_8673,N_8239,N_8083);
nand U8674 (N_8674,N_8201,N_8396);
nand U8675 (N_8675,N_8288,N_8136);
xor U8676 (N_8676,N_8314,N_8081);
or U8677 (N_8677,N_8191,N_8289);
xnor U8678 (N_8678,N_8350,N_8338);
and U8679 (N_8679,N_8377,N_8399);
or U8680 (N_8680,N_8121,N_8172);
or U8681 (N_8681,N_8113,N_8043);
nand U8682 (N_8682,N_8386,N_8077);
and U8683 (N_8683,N_8180,N_8086);
nor U8684 (N_8684,N_8098,N_8147);
xnor U8685 (N_8685,N_8061,N_8299);
nand U8686 (N_8686,N_8152,N_8310);
xor U8687 (N_8687,N_8155,N_8127);
and U8688 (N_8688,N_8085,N_8160);
xnor U8689 (N_8689,N_8306,N_8133);
nor U8690 (N_8690,N_8200,N_8063);
and U8691 (N_8691,N_8398,N_8261);
nor U8692 (N_8692,N_8301,N_8146);
nand U8693 (N_8693,N_8151,N_8076);
xor U8694 (N_8694,N_8236,N_8040);
nand U8695 (N_8695,N_8151,N_8259);
nor U8696 (N_8696,N_8132,N_8304);
and U8697 (N_8697,N_8067,N_8287);
and U8698 (N_8698,N_8363,N_8246);
nand U8699 (N_8699,N_8341,N_8006);
nand U8700 (N_8700,N_8242,N_8009);
or U8701 (N_8701,N_8322,N_8233);
or U8702 (N_8702,N_8123,N_8186);
xnor U8703 (N_8703,N_8217,N_8033);
nand U8704 (N_8704,N_8024,N_8027);
and U8705 (N_8705,N_8107,N_8299);
nor U8706 (N_8706,N_8203,N_8309);
xor U8707 (N_8707,N_8128,N_8178);
nand U8708 (N_8708,N_8177,N_8218);
and U8709 (N_8709,N_8210,N_8367);
nor U8710 (N_8710,N_8033,N_8386);
nor U8711 (N_8711,N_8132,N_8229);
nor U8712 (N_8712,N_8195,N_8084);
and U8713 (N_8713,N_8266,N_8176);
and U8714 (N_8714,N_8012,N_8075);
and U8715 (N_8715,N_8278,N_8019);
xor U8716 (N_8716,N_8088,N_8029);
nor U8717 (N_8717,N_8219,N_8375);
nor U8718 (N_8718,N_8054,N_8298);
xor U8719 (N_8719,N_8113,N_8180);
and U8720 (N_8720,N_8093,N_8220);
nor U8721 (N_8721,N_8033,N_8045);
or U8722 (N_8722,N_8311,N_8368);
and U8723 (N_8723,N_8387,N_8001);
nor U8724 (N_8724,N_8385,N_8046);
and U8725 (N_8725,N_8250,N_8076);
and U8726 (N_8726,N_8110,N_8070);
nor U8727 (N_8727,N_8219,N_8322);
or U8728 (N_8728,N_8130,N_8120);
nand U8729 (N_8729,N_8256,N_8242);
nor U8730 (N_8730,N_8317,N_8367);
nor U8731 (N_8731,N_8045,N_8325);
nor U8732 (N_8732,N_8283,N_8312);
or U8733 (N_8733,N_8068,N_8122);
and U8734 (N_8734,N_8377,N_8118);
nor U8735 (N_8735,N_8157,N_8102);
nor U8736 (N_8736,N_8159,N_8076);
nand U8737 (N_8737,N_8203,N_8215);
nand U8738 (N_8738,N_8101,N_8315);
and U8739 (N_8739,N_8155,N_8372);
and U8740 (N_8740,N_8260,N_8279);
and U8741 (N_8741,N_8284,N_8123);
and U8742 (N_8742,N_8387,N_8122);
nand U8743 (N_8743,N_8306,N_8175);
and U8744 (N_8744,N_8278,N_8000);
xor U8745 (N_8745,N_8038,N_8319);
nand U8746 (N_8746,N_8223,N_8283);
nor U8747 (N_8747,N_8016,N_8364);
and U8748 (N_8748,N_8108,N_8241);
and U8749 (N_8749,N_8277,N_8121);
nor U8750 (N_8750,N_8256,N_8235);
and U8751 (N_8751,N_8127,N_8003);
nor U8752 (N_8752,N_8225,N_8024);
or U8753 (N_8753,N_8043,N_8086);
nor U8754 (N_8754,N_8192,N_8061);
xnor U8755 (N_8755,N_8071,N_8350);
or U8756 (N_8756,N_8070,N_8215);
or U8757 (N_8757,N_8054,N_8190);
xnor U8758 (N_8758,N_8037,N_8178);
or U8759 (N_8759,N_8163,N_8149);
nor U8760 (N_8760,N_8012,N_8074);
or U8761 (N_8761,N_8024,N_8233);
nor U8762 (N_8762,N_8188,N_8324);
or U8763 (N_8763,N_8057,N_8218);
or U8764 (N_8764,N_8368,N_8078);
nor U8765 (N_8765,N_8391,N_8341);
nor U8766 (N_8766,N_8288,N_8249);
xor U8767 (N_8767,N_8261,N_8064);
and U8768 (N_8768,N_8200,N_8324);
or U8769 (N_8769,N_8071,N_8344);
and U8770 (N_8770,N_8087,N_8194);
nand U8771 (N_8771,N_8383,N_8065);
nand U8772 (N_8772,N_8214,N_8002);
nand U8773 (N_8773,N_8180,N_8350);
and U8774 (N_8774,N_8332,N_8008);
or U8775 (N_8775,N_8236,N_8175);
nand U8776 (N_8776,N_8261,N_8129);
or U8777 (N_8777,N_8375,N_8168);
or U8778 (N_8778,N_8045,N_8211);
nor U8779 (N_8779,N_8013,N_8133);
or U8780 (N_8780,N_8337,N_8025);
or U8781 (N_8781,N_8088,N_8363);
nand U8782 (N_8782,N_8361,N_8296);
xor U8783 (N_8783,N_8267,N_8233);
and U8784 (N_8784,N_8071,N_8204);
nor U8785 (N_8785,N_8212,N_8076);
nand U8786 (N_8786,N_8041,N_8023);
and U8787 (N_8787,N_8224,N_8092);
xnor U8788 (N_8788,N_8192,N_8213);
xor U8789 (N_8789,N_8308,N_8162);
xor U8790 (N_8790,N_8394,N_8242);
xnor U8791 (N_8791,N_8085,N_8042);
nand U8792 (N_8792,N_8049,N_8071);
xor U8793 (N_8793,N_8263,N_8325);
or U8794 (N_8794,N_8165,N_8080);
xnor U8795 (N_8795,N_8042,N_8322);
and U8796 (N_8796,N_8245,N_8241);
and U8797 (N_8797,N_8366,N_8374);
xnor U8798 (N_8798,N_8118,N_8112);
nand U8799 (N_8799,N_8324,N_8196);
nand U8800 (N_8800,N_8588,N_8696);
xor U8801 (N_8801,N_8748,N_8514);
nor U8802 (N_8802,N_8474,N_8591);
xor U8803 (N_8803,N_8475,N_8604);
nor U8804 (N_8804,N_8682,N_8651);
nand U8805 (N_8805,N_8614,N_8492);
xor U8806 (N_8806,N_8419,N_8733);
and U8807 (N_8807,N_8793,N_8573);
nor U8808 (N_8808,N_8508,N_8530);
nand U8809 (N_8809,N_8408,N_8473);
nor U8810 (N_8810,N_8746,N_8464);
xor U8811 (N_8811,N_8581,N_8586);
and U8812 (N_8812,N_8569,N_8714);
nand U8813 (N_8813,N_8520,N_8483);
nand U8814 (N_8814,N_8480,N_8669);
nand U8815 (N_8815,N_8570,N_8524);
xnor U8816 (N_8816,N_8576,N_8773);
xor U8817 (N_8817,N_8612,N_8684);
xnor U8818 (N_8818,N_8723,N_8704);
or U8819 (N_8819,N_8502,N_8525);
nor U8820 (N_8820,N_8797,N_8607);
nor U8821 (N_8821,N_8646,N_8499);
and U8822 (N_8822,N_8790,N_8517);
and U8823 (N_8823,N_8784,N_8407);
nor U8824 (N_8824,N_8726,N_8759);
or U8825 (N_8825,N_8565,N_8424);
and U8826 (N_8826,N_8645,N_8739);
xor U8827 (N_8827,N_8609,N_8467);
nor U8828 (N_8828,N_8495,N_8572);
nand U8829 (N_8829,N_8554,N_8453);
and U8830 (N_8830,N_8516,N_8425);
nand U8831 (N_8831,N_8428,N_8561);
nand U8832 (N_8832,N_8460,N_8452);
nand U8833 (N_8833,N_8724,N_8546);
nor U8834 (N_8834,N_8527,N_8403);
and U8835 (N_8835,N_8664,N_8519);
or U8836 (N_8836,N_8778,N_8788);
and U8837 (N_8837,N_8434,N_8789);
and U8838 (N_8838,N_8764,N_8648);
nand U8839 (N_8839,N_8549,N_8478);
xor U8840 (N_8840,N_8445,N_8537);
or U8841 (N_8841,N_8541,N_8463);
or U8842 (N_8842,N_8674,N_8738);
nor U8843 (N_8843,N_8550,N_8427);
and U8844 (N_8844,N_8617,N_8489);
xor U8845 (N_8845,N_8754,N_8484);
or U8846 (N_8846,N_8633,N_8639);
nand U8847 (N_8847,N_8566,N_8417);
nor U8848 (N_8848,N_8421,N_8433);
nor U8849 (N_8849,N_8681,N_8437);
xnor U8850 (N_8850,N_8785,N_8439);
nor U8851 (N_8851,N_8652,N_8624);
nor U8852 (N_8852,N_8683,N_8640);
or U8853 (N_8853,N_8486,N_8636);
nand U8854 (N_8854,N_8692,N_8736);
or U8855 (N_8855,N_8711,N_8623);
nand U8856 (N_8856,N_8718,N_8423);
or U8857 (N_8857,N_8757,N_8571);
or U8858 (N_8858,N_8481,N_8548);
and U8859 (N_8859,N_8575,N_8415);
xnor U8860 (N_8860,N_8668,N_8509);
nor U8861 (N_8861,N_8448,N_8606);
xor U8862 (N_8862,N_8765,N_8558);
nand U8863 (N_8863,N_8631,N_8485);
xnor U8864 (N_8864,N_8410,N_8597);
nor U8865 (N_8865,N_8698,N_8539);
or U8866 (N_8866,N_8488,N_8510);
xnor U8867 (N_8867,N_8563,N_8414);
nor U8868 (N_8868,N_8756,N_8659);
and U8869 (N_8869,N_8409,N_8479);
nand U8870 (N_8870,N_8552,N_8400);
nand U8871 (N_8871,N_8725,N_8647);
or U8872 (N_8872,N_8768,N_8740);
nand U8873 (N_8873,N_8616,N_8753);
nand U8874 (N_8874,N_8729,N_8441);
and U8875 (N_8875,N_8580,N_8625);
xnor U8876 (N_8876,N_8528,N_8432);
xnor U8877 (N_8877,N_8727,N_8670);
and U8878 (N_8878,N_8719,N_8534);
xnor U8879 (N_8879,N_8660,N_8611);
or U8880 (N_8880,N_8447,N_8717);
xor U8881 (N_8881,N_8654,N_8435);
and U8882 (N_8882,N_8406,N_8608);
and U8883 (N_8883,N_8587,N_8730);
xor U8884 (N_8884,N_8656,N_8713);
and U8885 (N_8885,N_8493,N_8701);
and U8886 (N_8886,N_8574,N_8497);
or U8887 (N_8887,N_8521,N_8705);
xor U8888 (N_8888,N_8796,N_8500);
or U8889 (N_8889,N_8413,N_8430);
or U8890 (N_8890,N_8637,N_8506);
and U8891 (N_8891,N_8540,N_8551);
or U8892 (N_8892,N_8622,N_8568);
nor U8893 (N_8893,N_8470,N_8661);
nand U8894 (N_8894,N_8672,N_8487);
and U8895 (N_8895,N_8629,N_8451);
xnor U8896 (N_8896,N_8578,N_8589);
nand U8897 (N_8897,N_8469,N_8583);
xor U8898 (N_8898,N_8700,N_8742);
nor U8899 (N_8899,N_8496,N_8596);
xor U8900 (N_8900,N_8777,N_8542);
xnor U8901 (N_8901,N_8728,N_8538);
or U8902 (N_8902,N_8787,N_8613);
nand U8903 (N_8903,N_8454,N_8456);
and U8904 (N_8904,N_8709,N_8544);
nor U8905 (N_8905,N_8455,N_8595);
nor U8906 (N_8906,N_8559,N_8721);
xor U8907 (N_8907,N_8676,N_8774);
nand U8908 (N_8908,N_8716,N_8515);
nand U8909 (N_8909,N_8780,N_8436);
or U8910 (N_8910,N_8642,N_8560);
or U8911 (N_8911,N_8644,N_8507);
nand U8912 (N_8912,N_8665,N_8501);
nor U8913 (N_8913,N_8511,N_8603);
nor U8914 (N_8914,N_8638,N_8786);
or U8915 (N_8915,N_8641,N_8649);
nor U8916 (N_8916,N_8752,N_8564);
xnor U8917 (N_8917,N_8402,N_8601);
nor U8918 (N_8918,N_8630,N_8533);
or U8919 (N_8919,N_8699,N_8518);
nor U8920 (N_8920,N_8468,N_8663);
and U8921 (N_8921,N_8476,N_8431);
nand U8922 (N_8922,N_8734,N_8689);
nand U8923 (N_8923,N_8771,N_8459);
or U8924 (N_8924,N_8535,N_8465);
and U8925 (N_8925,N_8557,N_8556);
and U8926 (N_8926,N_8593,N_8703);
or U8927 (N_8927,N_8671,N_8675);
or U8928 (N_8928,N_8599,N_8602);
nor U8929 (N_8929,N_8769,N_8767);
or U8930 (N_8930,N_8567,N_8662);
and U8931 (N_8931,N_8761,N_8776);
nand U8932 (N_8932,N_8781,N_8401);
xnor U8933 (N_8933,N_8526,N_8600);
nand U8934 (N_8934,N_8763,N_8693);
xor U8935 (N_8935,N_8498,N_8422);
xor U8936 (N_8936,N_8782,N_8655);
nor U8937 (N_8937,N_8582,N_8412);
nand U8938 (N_8938,N_8420,N_8450);
nand U8939 (N_8939,N_8505,N_8710);
or U8940 (N_8940,N_8536,N_8585);
nand U8941 (N_8941,N_8743,N_8504);
nand U8942 (N_8942,N_8594,N_8691);
nor U8943 (N_8943,N_8523,N_8513);
xnor U8944 (N_8944,N_8628,N_8418);
xor U8945 (N_8945,N_8720,N_8766);
nor U8946 (N_8946,N_8737,N_8695);
nor U8947 (N_8947,N_8694,N_8744);
and U8948 (N_8948,N_8758,N_8750);
xnor U8949 (N_8949,N_8678,N_8762);
nor U8950 (N_8950,N_8532,N_8482);
or U8951 (N_8951,N_8687,N_8531);
nor U8952 (N_8952,N_8547,N_8783);
and U8953 (N_8953,N_8735,N_8706);
xor U8954 (N_8954,N_8626,N_8477);
and U8955 (N_8955,N_8627,N_8795);
nor U8956 (N_8956,N_8775,N_8697);
and U8957 (N_8957,N_8794,N_8590);
or U8958 (N_8958,N_8555,N_8749);
xnor U8959 (N_8959,N_8650,N_8666);
nand U8960 (N_8960,N_8620,N_8471);
nand U8961 (N_8961,N_8619,N_8529);
xor U8962 (N_8962,N_8494,N_8449);
and U8963 (N_8963,N_8702,N_8598);
and U8964 (N_8964,N_8751,N_8690);
and U8965 (N_8965,N_8579,N_8466);
or U8966 (N_8966,N_8715,N_8426);
nor U8967 (N_8967,N_8444,N_8621);
or U8968 (N_8968,N_8722,N_8708);
xor U8969 (N_8969,N_8440,N_8462);
or U8970 (N_8970,N_8618,N_8686);
xor U8971 (N_8971,N_8405,N_8772);
nor U8972 (N_8972,N_8634,N_8677);
xor U8973 (N_8973,N_8792,N_8442);
or U8974 (N_8974,N_8438,N_8667);
nand U8975 (N_8975,N_8562,N_8741);
and U8976 (N_8976,N_8632,N_8472);
xor U8977 (N_8977,N_8457,N_8653);
xnor U8978 (N_8978,N_8635,N_8592);
or U8979 (N_8979,N_8461,N_8446);
xnor U8980 (N_8980,N_8490,N_8615);
nand U8981 (N_8981,N_8770,N_8799);
and U8982 (N_8982,N_8755,N_8658);
nor U8983 (N_8983,N_8503,N_8610);
nand U8984 (N_8984,N_8707,N_8512);
or U8985 (N_8985,N_8688,N_8679);
or U8986 (N_8986,N_8553,N_8543);
xor U8987 (N_8987,N_8411,N_8731);
nor U8988 (N_8988,N_8443,N_8673);
nor U8989 (N_8989,N_8643,N_8429);
xnor U8990 (N_8990,N_8712,N_8760);
or U8991 (N_8991,N_8404,N_8545);
and U8992 (N_8992,N_8791,N_8732);
nand U8993 (N_8993,N_8680,N_8745);
nand U8994 (N_8994,N_8657,N_8491);
or U8995 (N_8995,N_8458,N_8584);
nor U8996 (N_8996,N_8577,N_8798);
nor U8997 (N_8997,N_8779,N_8605);
and U8998 (N_8998,N_8522,N_8416);
or U8999 (N_8999,N_8685,N_8747);
nor U9000 (N_9000,N_8713,N_8526);
nor U9001 (N_9001,N_8583,N_8480);
nand U9002 (N_9002,N_8718,N_8619);
nor U9003 (N_9003,N_8609,N_8785);
nor U9004 (N_9004,N_8647,N_8485);
nor U9005 (N_9005,N_8749,N_8447);
xnor U9006 (N_9006,N_8522,N_8502);
nor U9007 (N_9007,N_8655,N_8578);
nand U9008 (N_9008,N_8606,N_8697);
and U9009 (N_9009,N_8528,N_8623);
xnor U9010 (N_9010,N_8631,N_8487);
nand U9011 (N_9011,N_8400,N_8468);
or U9012 (N_9012,N_8402,N_8495);
nand U9013 (N_9013,N_8703,N_8602);
and U9014 (N_9014,N_8663,N_8780);
or U9015 (N_9015,N_8633,N_8642);
xnor U9016 (N_9016,N_8542,N_8766);
nor U9017 (N_9017,N_8782,N_8609);
nor U9018 (N_9018,N_8787,N_8587);
and U9019 (N_9019,N_8719,N_8478);
xor U9020 (N_9020,N_8605,N_8530);
nand U9021 (N_9021,N_8471,N_8584);
and U9022 (N_9022,N_8657,N_8718);
xnor U9023 (N_9023,N_8641,N_8450);
or U9024 (N_9024,N_8786,N_8411);
nor U9025 (N_9025,N_8449,N_8451);
and U9026 (N_9026,N_8641,N_8501);
or U9027 (N_9027,N_8528,N_8762);
nand U9028 (N_9028,N_8502,N_8537);
or U9029 (N_9029,N_8635,N_8721);
and U9030 (N_9030,N_8524,N_8766);
nand U9031 (N_9031,N_8714,N_8535);
xor U9032 (N_9032,N_8724,N_8638);
xnor U9033 (N_9033,N_8672,N_8496);
or U9034 (N_9034,N_8437,N_8590);
nor U9035 (N_9035,N_8449,N_8578);
or U9036 (N_9036,N_8708,N_8660);
and U9037 (N_9037,N_8672,N_8483);
nand U9038 (N_9038,N_8504,N_8645);
xnor U9039 (N_9039,N_8706,N_8571);
xor U9040 (N_9040,N_8768,N_8479);
and U9041 (N_9041,N_8760,N_8783);
nand U9042 (N_9042,N_8564,N_8615);
or U9043 (N_9043,N_8688,N_8419);
and U9044 (N_9044,N_8717,N_8544);
nand U9045 (N_9045,N_8765,N_8665);
and U9046 (N_9046,N_8722,N_8669);
or U9047 (N_9047,N_8412,N_8473);
or U9048 (N_9048,N_8713,N_8495);
nand U9049 (N_9049,N_8436,N_8474);
and U9050 (N_9050,N_8583,N_8745);
xor U9051 (N_9051,N_8768,N_8608);
or U9052 (N_9052,N_8612,N_8408);
and U9053 (N_9053,N_8763,N_8699);
and U9054 (N_9054,N_8649,N_8687);
or U9055 (N_9055,N_8536,N_8441);
and U9056 (N_9056,N_8748,N_8799);
nor U9057 (N_9057,N_8772,N_8440);
xnor U9058 (N_9058,N_8799,N_8490);
xnor U9059 (N_9059,N_8780,N_8529);
and U9060 (N_9060,N_8650,N_8427);
xor U9061 (N_9061,N_8452,N_8463);
nand U9062 (N_9062,N_8526,N_8464);
nand U9063 (N_9063,N_8711,N_8766);
nand U9064 (N_9064,N_8460,N_8708);
or U9065 (N_9065,N_8701,N_8433);
or U9066 (N_9066,N_8488,N_8543);
nand U9067 (N_9067,N_8656,N_8582);
xnor U9068 (N_9068,N_8516,N_8573);
nand U9069 (N_9069,N_8584,N_8700);
and U9070 (N_9070,N_8692,N_8640);
xor U9071 (N_9071,N_8624,N_8416);
or U9072 (N_9072,N_8411,N_8645);
nor U9073 (N_9073,N_8608,N_8716);
or U9074 (N_9074,N_8457,N_8419);
nor U9075 (N_9075,N_8580,N_8787);
or U9076 (N_9076,N_8664,N_8457);
or U9077 (N_9077,N_8574,N_8436);
and U9078 (N_9078,N_8434,N_8422);
nor U9079 (N_9079,N_8778,N_8515);
xor U9080 (N_9080,N_8442,N_8551);
xor U9081 (N_9081,N_8639,N_8694);
xor U9082 (N_9082,N_8676,N_8762);
nand U9083 (N_9083,N_8642,N_8421);
and U9084 (N_9084,N_8743,N_8551);
or U9085 (N_9085,N_8766,N_8675);
or U9086 (N_9086,N_8796,N_8563);
or U9087 (N_9087,N_8730,N_8653);
xnor U9088 (N_9088,N_8789,N_8406);
or U9089 (N_9089,N_8785,N_8648);
nor U9090 (N_9090,N_8659,N_8629);
nor U9091 (N_9091,N_8594,N_8700);
xnor U9092 (N_9092,N_8662,N_8756);
nor U9093 (N_9093,N_8415,N_8761);
or U9094 (N_9094,N_8571,N_8694);
xnor U9095 (N_9095,N_8562,N_8744);
nand U9096 (N_9096,N_8409,N_8764);
or U9097 (N_9097,N_8538,N_8699);
or U9098 (N_9098,N_8489,N_8698);
nor U9099 (N_9099,N_8703,N_8608);
and U9100 (N_9100,N_8561,N_8710);
and U9101 (N_9101,N_8705,N_8529);
or U9102 (N_9102,N_8717,N_8521);
nand U9103 (N_9103,N_8637,N_8757);
and U9104 (N_9104,N_8460,N_8788);
nor U9105 (N_9105,N_8490,N_8732);
and U9106 (N_9106,N_8533,N_8797);
xnor U9107 (N_9107,N_8524,N_8568);
nand U9108 (N_9108,N_8702,N_8509);
and U9109 (N_9109,N_8692,N_8466);
and U9110 (N_9110,N_8579,N_8586);
or U9111 (N_9111,N_8507,N_8730);
xor U9112 (N_9112,N_8528,N_8533);
and U9113 (N_9113,N_8499,N_8708);
nor U9114 (N_9114,N_8472,N_8716);
and U9115 (N_9115,N_8695,N_8597);
and U9116 (N_9116,N_8483,N_8566);
nor U9117 (N_9117,N_8668,N_8681);
nand U9118 (N_9118,N_8453,N_8636);
or U9119 (N_9119,N_8512,N_8661);
and U9120 (N_9120,N_8616,N_8478);
xnor U9121 (N_9121,N_8413,N_8727);
xnor U9122 (N_9122,N_8672,N_8489);
nand U9123 (N_9123,N_8750,N_8531);
or U9124 (N_9124,N_8474,N_8737);
nor U9125 (N_9125,N_8797,N_8528);
or U9126 (N_9126,N_8509,N_8479);
nor U9127 (N_9127,N_8785,N_8783);
and U9128 (N_9128,N_8530,N_8460);
nand U9129 (N_9129,N_8501,N_8413);
and U9130 (N_9130,N_8580,N_8521);
nand U9131 (N_9131,N_8495,N_8490);
or U9132 (N_9132,N_8770,N_8533);
or U9133 (N_9133,N_8751,N_8582);
nand U9134 (N_9134,N_8502,N_8607);
nand U9135 (N_9135,N_8569,N_8469);
nand U9136 (N_9136,N_8604,N_8608);
nand U9137 (N_9137,N_8565,N_8582);
xnor U9138 (N_9138,N_8470,N_8529);
nor U9139 (N_9139,N_8596,N_8648);
xnor U9140 (N_9140,N_8472,N_8516);
xor U9141 (N_9141,N_8661,N_8697);
or U9142 (N_9142,N_8418,N_8710);
nand U9143 (N_9143,N_8744,N_8726);
nor U9144 (N_9144,N_8652,N_8531);
nor U9145 (N_9145,N_8510,N_8413);
and U9146 (N_9146,N_8499,N_8584);
xnor U9147 (N_9147,N_8721,N_8620);
nor U9148 (N_9148,N_8446,N_8752);
nor U9149 (N_9149,N_8436,N_8550);
or U9150 (N_9150,N_8696,N_8520);
and U9151 (N_9151,N_8455,N_8562);
nor U9152 (N_9152,N_8436,N_8691);
and U9153 (N_9153,N_8642,N_8500);
xnor U9154 (N_9154,N_8484,N_8526);
and U9155 (N_9155,N_8517,N_8780);
and U9156 (N_9156,N_8508,N_8539);
nor U9157 (N_9157,N_8661,N_8792);
or U9158 (N_9158,N_8575,N_8442);
xnor U9159 (N_9159,N_8691,N_8622);
xor U9160 (N_9160,N_8783,N_8537);
xor U9161 (N_9161,N_8629,N_8553);
xor U9162 (N_9162,N_8553,N_8602);
xor U9163 (N_9163,N_8531,N_8577);
nand U9164 (N_9164,N_8621,N_8633);
nor U9165 (N_9165,N_8797,N_8609);
nor U9166 (N_9166,N_8769,N_8527);
nor U9167 (N_9167,N_8567,N_8478);
nor U9168 (N_9168,N_8507,N_8722);
nand U9169 (N_9169,N_8618,N_8451);
and U9170 (N_9170,N_8763,N_8688);
nor U9171 (N_9171,N_8499,N_8529);
xnor U9172 (N_9172,N_8672,N_8690);
xnor U9173 (N_9173,N_8644,N_8557);
or U9174 (N_9174,N_8727,N_8633);
xor U9175 (N_9175,N_8605,N_8709);
xnor U9176 (N_9176,N_8470,N_8428);
xor U9177 (N_9177,N_8715,N_8671);
nand U9178 (N_9178,N_8560,N_8659);
xnor U9179 (N_9179,N_8622,N_8541);
and U9180 (N_9180,N_8651,N_8672);
xnor U9181 (N_9181,N_8431,N_8738);
nand U9182 (N_9182,N_8605,N_8705);
xnor U9183 (N_9183,N_8641,N_8789);
or U9184 (N_9184,N_8475,N_8668);
xnor U9185 (N_9185,N_8687,N_8660);
nor U9186 (N_9186,N_8790,N_8695);
or U9187 (N_9187,N_8597,N_8458);
and U9188 (N_9188,N_8438,N_8641);
and U9189 (N_9189,N_8475,N_8763);
and U9190 (N_9190,N_8679,N_8592);
xnor U9191 (N_9191,N_8678,N_8654);
and U9192 (N_9192,N_8721,N_8740);
and U9193 (N_9193,N_8438,N_8531);
or U9194 (N_9194,N_8768,N_8622);
or U9195 (N_9195,N_8597,N_8514);
or U9196 (N_9196,N_8671,N_8588);
nand U9197 (N_9197,N_8526,N_8538);
nor U9198 (N_9198,N_8530,N_8760);
or U9199 (N_9199,N_8482,N_8484);
or U9200 (N_9200,N_8971,N_8894);
or U9201 (N_9201,N_8978,N_8854);
nor U9202 (N_9202,N_9059,N_9150);
xnor U9203 (N_9203,N_8875,N_9137);
xor U9204 (N_9204,N_8960,N_9064);
or U9205 (N_9205,N_8891,N_9107);
and U9206 (N_9206,N_8956,N_9034);
nor U9207 (N_9207,N_9015,N_9177);
or U9208 (N_9208,N_9124,N_9099);
xnor U9209 (N_9209,N_9142,N_9032);
or U9210 (N_9210,N_9149,N_8982);
xor U9211 (N_9211,N_9069,N_8905);
xor U9212 (N_9212,N_8964,N_8916);
nand U9213 (N_9213,N_9006,N_8828);
nand U9214 (N_9214,N_8840,N_8924);
nand U9215 (N_9215,N_8803,N_8805);
or U9216 (N_9216,N_9085,N_9030);
nor U9217 (N_9217,N_8902,N_9089);
nor U9218 (N_9218,N_9072,N_8892);
nand U9219 (N_9219,N_8830,N_8896);
nand U9220 (N_9220,N_8808,N_8801);
or U9221 (N_9221,N_8913,N_9047);
nand U9222 (N_9222,N_8987,N_9160);
nor U9223 (N_9223,N_9174,N_8959);
xnor U9224 (N_9224,N_9037,N_8813);
nand U9225 (N_9225,N_8863,N_8999);
nand U9226 (N_9226,N_9018,N_9168);
nand U9227 (N_9227,N_8886,N_9139);
nor U9228 (N_9228,N_8867,N_8906);
and U9229 (N_9229,N_8893,N_8909);
nand U9230 (N_9230,N_8983,N_9082);
nand U9231 (N_9231,N_9170,N_9148);
nor U9232 (N_9232,N_9087,N_9046);
nor U9233 (N_9233,N_9054,N_8878);
xnor U9234 (N_9234,N_9005,N_9126);
or U9235 (N_9235,N_8991,N_9179);
and U9236 (N_9236,N_9144,N_9100);
nor U9237 (N_9237,N_8972,N_9039);
xor U9238 (N_9238,N_8915,N_8861);
or U9239 (N_9239,N_8953,N_8809);
nor U9240 (N_9240,N_8925,N_9128);
xnor U9241 (N_9241,N_9096,N_9033);
and U9242 (N_9242,N_8821,N_9029);
or U9243 (N_9243,N_8986,N_8997);
or U9244 (N_9244,N_9021,N_8988);
or U9245 (N_9245,N_8980,N_8873);
nor U9246 (N_9246,N_8818,N_8967);
nor U9247 (N_9247,N_8827,N_8900);
xor U9248 (N_9248,N_8898,N_8928);
xor U9249 (N_9249,N_9004,N_9116);
or U9250 (N_9250,N_9061,N_8974);
and U9251 (N_9251,N_8897,N_9023);
and U9252 (N_9252,N_8885,N_8831);
nand U9253 (N_9253,N_9080,N_8976);
or U9254 (N_9254,N_8984,N_9153);
xnor U9255 (N_9255,N_9156,N_9119);
nor U9256 (N_9256,N_9014,N_9191);
xor U9257 (N_9257,N_9042,N_8936);
or U9258 (N_9258,N_9196,N_9152);
and U9259 (N_9259,N_8910,N_9162);
nand U9260 (N_9260,N_8958,N_8853);
nor U9261 (N_9261,N_8911,N_8800);
xnor U9262 (N_9262,N_9008,N_8890);
or U9263 (N_9263,N_8825,N_8823);
xnor U9264 (N_9264,N_9075,N_8824);
nand U9265 (N_9265,N_9184,N_8946);
nor U9266 (N_9266,N_9133,N_9113);
xor U9267 (N_9267,N_9055,N_8804);
xnor U9268 (N_9268,N_8985,N_9165);
xor U9269 (N_9269,N_9026,N_9091);
xnor U9270 (N_9270,N_8942,N_8817);
and U9271 (N_9271,N_9172,N_8859);
nand U9272 (N_9272,N_9189,N_9105);
nor U9273 (N_9273,N_8865,N_9135);
nor U9274 (N_9274,N_8895,N_9171);
nor U9275 (N_9275,N_9058,N_8903);
xor U9276 (N_9276,N_9073,N_9114);
and U9277 (N_9277,N_8832,N_9199);
nand U9278 (N_9278,N_9195,N_9130);
nand U9279 (N_9279,N_9079,N_9163);
or U9280 (N_9280,N_8848,N_8837);
nor U9281 (N_9281,N_8917,N_8869);
nor U9282 (N_9282,N_8908,N_8949);
or U9283 (N_9283,N_9193,N_8922);
xor U9284 (N_9284,N_9118,N_8899);
and U9285 (N_9285,N_8802,N_8851);
xor U9286 (N_9286,N_9183,N_9088);
or U9287 (N_9287,N_9143,N_9090);
nor U9288 (N_9288,N_8981,N_9141);
nand U9289 (N_9289,N_8940,N_9093);
xor U9290 (N_9290,N_8975,N_8864);
nor U9291 (N_9291,N_8932,N_8935);
xor U9292 (N_9292,N_9041,N_9035);
or U9293 (N_9293,N_9062,N_9007);
nand U9294 (N_9294,N_8833,N_9036);
xor U9295 (N_9295,N_8874,N_9084);
nand U9296 (N_9296,N_9154,N_8994);
nor U9297 (N_9297,N_8965,N_9169);
nor U9298 (N_9298,N_9020,N_9031);
xnor U9299 (N_9299,N_8871,N_9098);
nand U9300 (N_9300,N_8839,N_8934);
and U9301 (N_9301,N_9051,N_8998);
xor U9302 (N_9302,N_8901,N_9001);
xnor U9303 (N_9303,N_9044,N_9028);
xor U9304 (N_9304,N_9186,N_8961);
xor U9305 (N_9305,N_9083,N_9104);
or U9306 (N_9306,N_9092,N_8927);
or U9307 (N_9307,N_8846,N_9131);
nand U9308 (N_9308,N_9145,N_8933);
or U9309 (N_9309,N_9159,N_8814);
and U9310 (N_9310,N_8847,N_8938);
xnor U9311 (N_9311,N_9158,N_8963);
or U9312 (N_9312,N_8968,N_9115);
and U9313 (N_9313,N_8844,N_9000);
and U9314 (N_9314,N_8877,N_9056);
xnor U9315 (N_9315,N_8931,N_8919);
and U9316 (N_9316,N_8941,N_9016);
nor U9317 (N_9317,N_9192,N_9017);
nor U9318 (N_9318,N_8856,N_9102);
and U9319 (N_9319,N_9147,N_9022);
xnor U9320 (N_9320,N_8841,N_9129);
or U9321 (N_9321,N_9040,N_9112);
xnor U9322 (N_9322,N_9038,N_8950);
nand U9323 (N_9323,N_9188,N_9178);
xor U9324 (N_9324,N_9002,N_9138);
nor U9325 (N_9325,N_9109,N_9157);
or U9326 (N_9326,N_9019,N_8970);
xnor U9327 (N_9327,N_9197,N_8929);
and U9328 (N_9328,N_8921,N_9164);
nand U9329 (N_9329,N_9187,N_8945);
xor U9330 (N_9330,N_8836,N_9048);
xnor U9331 (N_9331,N_9166,N_8834);
nor U9332 (N_9332,N_9194,N_9097);
nor U9333 (N_9333,N_8973,N_8845);
nor U9334 (N_9334,N_8862,N_9045);
and U9335 (N_9335,N_9111,N_9081);
and U9336 (N_9336,N_8904,N_9086);
nand U9337 (N_9337,N_8843,N_9103);
xor U9338 (N_9338,N_9185,N_9027);
and U9339 (N_9339,N_8948,N_8914);
or U9340 (N_9340,N_9101,N_8954);
xnor U9341 (N_9341,N_8868,N_9120);
and U9342 (N_9342,N_8951,N_9010);
nand U9343 (N_9343,N_9176,N_9127);
nor U9344 (N_9344,N_8822,N_9151);
or U9345 (N_9345,N_9060,N_9161);
xor U9346 (N_9346,N_8883,N_9173);
xnor U9347 (N_9347,N_8815,N_9198);
nand U9348 (N_9348,N_9180,N_8993);
nor U9349 (N_9349,N_8969,N_8850);
xnor U9350 (N_9350,N_9011,N_8912);
and U9351 (N_9351,N_9108,N_8955);
and U9352 (N_9352,N_9181,N_8855);
nand U9353 (N_9353,N_9063,N_8937);
nand U9354 (N_9354,N_8838,N_9125);
nor U9355 (N_9355,N_8879,N_9012);
and U9356 (N_9356,N_8889,N_8880);
nor U9357 (N_9357,N_8977,N_8872);
or U9358 (N_9358,N_9132,N_8952);
nand U9359 (N_9359,N_8966,N_8990);
nor U9360 (N_9360,N_8812,N_9009);
xor U9361 (N_9361,N_8829,N_9043);
nor U9362 (N_9362,N_8884,N_8826);
xor U9363 (N_9363,N_8939,N_8979);
nor U9364 (N_9364,N_9095,N_9146);
xor U9365 (N_9365,N_9053,N_8907);
nand U9366 (N_9366,N_9136,N_8811);
and U9367 (N_9367,N_8849,N_8870);
nor U9368 (N_9368,N_9067,N_8989);
nand U9369 (N_9369,N_9078,N_9025);
nor U9370 (N_9370,N_8920,N_9074);
nand U9371 (N_9371,N_8852,N_8819);
nor U9372 (N_9372,N_9122,N_9070);
xnor U9373 (N_9373,N_8887,N_9052);
or U9374 (N_9374,N_8881,N_9117);
or U9375 (N_9375,N_8996,N_9140);
nand U9376 (N_9376,N_9050,N_9182);
and U9377 (N_9377,N_9175,N_9071);
nand U9378 (N_9378,N_9123,N_8835);
and U9379 (N_9379,N_8926,N_9094);
nand U9380 (N_9380,N_8888,N_9121);
or U9381 (N_9381,N_8943,N_9077);
and U9382 (N_9382,N_8882,N_9076);
or U9383 (N_9383,N_8957,N_8947);
or U9384 (N_9384,N_9066,N_8860);
nor U9385 (N_9385,N_8816,N_8806);
nor U9386 (N_9386,N_8810,N_8918);
xor U9387 (N_9387,N_9167,N_8930);
nand U9388 (N_9388,N_8962,N_8820);
xor U9389 (N_9389,N_8992,N_9057);
nor U9390 (N_9390,N_8842,N_9106);
or U9391 (N_9391,N_9065,N_9110);
xor U9392 (N_9392,N_8944,N_9155);
and U9393 (N_9393,N_8866,N_9003);
xor U9394 (N_9394,N_9024,N_9049);
nand U9395 (N_9395,N_8858,N_8876);
or U9396 (N_9396,N_8807,N_9068);
or U9397 (N_9397,N_9013,N_8923);
xor U9398 (N_9398,N_9190,N_8857);
or U9399 (N_9399,N_8995,N_9134);
or U9400 (N_9400,N_9166,N_9050);
nand U9401 (N_9401,N_8954,N_9172);
nand U9402 (N_9402,N_9121,N_9031);
nor U9403 (N_9403,N_8999,N_9147);
nor U9404 (N_9404,N_8934,N_8954);
nor U9405 (N_9405,N_9103,N_9011);
xnor U9406 (N_9406,N_8833,N_9070);
and U9407 (N_9407,N_8920,N_9060);
and U9408 (N_9408,N_8816,N_9190);
or U9409 (N_9409,N_8931,N_9124);
nand U9410 (N_9410,N_9155,N_9045);
nand U9411 (N_9411,N_8841,N_9114);
and U9412 (N_9412,N_8944,N_8953);
nand U9413 (N_9413,N_9039,N_9005);
xor U9414 (N_9414,N_9139,N_8840);
or U9415 (N_9415,N_9191,N_9030);
xnor U9416 (N_9416,N_8892,N_8801);
xor U9417 (N_9417,N_8883,N_9110);
and U9418 (N_9418,N_9017,N_9184);
and U9419 (N_9419,N_8830,N_8979);
xnor U9420 (N_9420,N_8855,N_9148);
or U9421 (N_9421,N_9057,N_9194);
nor U9422 (N_9422,N_9198,N_8820);
and U9423 (N_9423,N_9182,N_8880);
nor U9424 (N_9424,N_9167,N_8929);
or U9425 (N_9425,N_9151,N_8900);
xor U9426 (N_9426,N_9083,N_9178);
and U9427 (N_9427,N_8987,N_8863);
or U9428 (N_9428,N_8823,N_8893);
xor U9429 (N_9429,N_9096,N_9179);
and U9430 (N_9430,N_9118,N_8801);
nor U9431 (N_9431,N_8829,N_8983);
nor U9432 (N_9432,N_9198,N_8901);
nand U9433 (N_9433,N_8951,N_8809);
nor U9434 (N_9434,N_9198,N_9020);
nor U9435 (N_9435,N_8928,N_8841);
nor U9436 (N_9436,N_9014,N_8963);
and U9437 (N_9437,N_9083,N_8987);
nand U9438 (N_9438,N_9053,N_9023);
xor U9439 (N_9439,N_9137,N_9083);
and U9440 (N_9440,N_9027,N_9044);
nand U9441 (N_9441,N_8957,N_8909);
and U9442 (N_9442,N_8810,N_9046);
or U9443 (N_9443,N_8855,N_8927);
xnor U9444 (N_9444,N_9036,N_9034);
xnor U9445 (N_9445,N_9006,N_8970);
or U9446 (N_9446,N_9081,N_8997);
nand U9447 (N_9447,N_8990,N_9169);
and U9448 (N_9448,N_8985,N_8823);
or U9449 (N_9449,N_9170,N_9122);
xor U9450 (N_9450,N_8874,N_8964);
and U9451 (N_9451,N_8926,N_8807);
xor U9452 (N_9452,N_9063,N_8891);
nand U9453 (N_9453,N_9072,N_9071);
nand U9454 (N_9454,N_8949,N_8904);
nor U9455 (N_9455,N_8967,N_8938);
nand U9456 (N_9456,N_9027,N_8860);
or U9457 (N_9457,N_9117,N_9108);
or U9458 (N_9458,N_9169,N_9053);
nor U9459 (N_9459,N_9018,N_9108);
or U9460 (N_9460,N_9171,N_8813);
or U9461 (N_9461,N_9082,N_8892);
xor U9462 (N_9462,N_9050,N_9151);
nand U9463 (N_9463,N_8940,N_8912);
or U9464 (N_9464,N_8829,N_9001);
and U9465 (N_9465,N_8954,N_8839);
or U9466 (N_9466,N_9004,N_9181);
nor U9467 (N_9467,N_9197,N_9002);
nor U9468 (N_9468,N_9045,N_9018);
nand U9469 (N_9469,N_8942,N_9166);
nand U9470 (N_9470,N_9063,N_8884);
xor U9471 (N_9471,N_9166,N_9067);
or U9472 (N_9472,N_8901,N_8939);
xnor U9473 (N_9473,N_9107,N_9105);
nand U9474 (N_9474,N_9095,N_9125);
nor U9475 (N_9475,N_8811,N_8915);
and U9476 (N_9476,N_9020,N_8902);
nand U9477 (N_9477,N_9141,N_9184);
xnor U9478 (N_9478,N_9127,N_9079);
xor U9479 (N_9479,N_8964,N_8859);
xnor U9480 (N_9480,N_9146,N_9191);
or U9481 (N_9481,N_8958,N_9097);
nand U9482 (N_9482,N_8926,N_8887);
nand U9483 (N_9483,N_9085,N_8823);
nor U9484 (N_9484,N_8833,N_9042);
nand U9485 (N_9485,N_8994,N_9084);
xnor U9486 (N_9486,N_8941,N_8968);
or U9487 (N_9487,N_9115,N_9024);
nand U9488 (N_9488,N_8842,N_8929);
nor U9489 (N_9489,N_9152,N_9082);
nor U9490 (N_9490,N_8846,N_9080);
and U9491 (N_9491,N_8994,N_9000);
nand U9492 (N_9492,N_8856,N_9001);
and U9493 (N_9493,N_9175,N_9086);
and U9494 (N_9494,N_8847,N_8916);
nor U9495 (N_9495,N_8852,N_9157);
and U9496 (N_9496,N_9076,N_8970);
and U9497 (N_9497,N_9175,N_9166);
and U9498 (N_9498,N_9156,N_8868);
or U9499 (N_9499,N_9160,N_8803);
nand U9500 (N_9500,N_8980,N_9154);
xor U9501 (N_9501,N_8974,N_8924);
nor U9502 (N_9502,N_8968,N_8834);
or U9503 (N_9503,N_8854,N_8813);
and U9504 (N_9504,N_8962,N_9061);
xor U9505 (N_9505,N_9170,N_8958);
and U9506 (N_9506,N_9056,N_9155);
and U9507 (N_9507,N_9031,N_9000);
nor U9508 (N_9508,N_9060,N_9028);
and U9509 (N_9509,N_9103,N_9198);
xnor U9510 (N_9510,N_8906,N_8880);
or U9511 (N_9511,N_8903,N_9116);
nand U9512 (N_9512,N_8945,N_9019);
xor U9513 (N_9513,N_9059,N_9054);
and U9514 (N_9514,N_8860,N_8843);
nor U9515 (N_9515,N_9013,N_8829);
nor U9516 (N_9516,N_8804,N_9086);
nor U9517 (N_9517,N_9002,N_8897);
nand U9518 (N_9518,N_9173,N_8982);
nand U9519 (N_9519,N_9067,N_9143);
xnor U9520 (N_9520,N_9110,N_9170);
nor U9521 (N_9521,N_9011,N_9126);
and U9522 (N_9522,N_8952,N_8935);
nor U9523 (N_9523,N_8920,N_9171);
and U9524 (N_9524,N_9125,N_9003);
nor U9525 (N_9525,N_8849,N_8972);
and U9526 (N_9526,N_8807,N_9165);
xor U9527 (N_9527,N_9199,N_8987);
or U9528 (N_9528,N_9147,N_8921);
nor U9529 (N_9529,N_9140,N_8923);
or U9530 (N_9530,N_8917,N_8902);
nor U9531 (N_9531,N_9184,N_8941);
and U9532 (N_9532,N_9017,N_8908);
nand U9533 (N_9533,N_8843,N_8879);
and U9534 (N_9534,N_9065,N_9102);
nand U9535 (N_9535,N_9117,N_9196);
nor U9536 (N_9536,N_8847,N_9037);
xor U9537 (N_9537,N_9146,N_9085);
xor U9538 (N_9538,N_9187,N_8917);
nor U9539 (N_9539,N_9069,N_8975);
nand U9540 (N_9540,N_8941,N_9035);
xor U9541 (N_9541,N_9194,N_9051);
nand U9542 (N_9542,N_8986,N_8853);
nand U9543 (N_9543,N_9073,N_9106);
or U9544 (N_9544,N_9138,N_9079);
nor U9545 (N_9545,N_9147,N_9102);
xnor U9546 (N_9546,N_8859,N_9153);
nand U9547 (N_9547,N_9064,N_8852);
nand U9548 (N_9548,N_9174,N_8911);
or U9549 (N_9549,N_8932,N_9120);
xnor U9550 (N_9550,N_9118,N_9090);
nand U9551 (N_9551,N_8883,N_8948);
and U9552 (N_9552,N_8973,N_9036);
nand U9553 (N_9553,N_8976,N_8919);
nor U9554 (N_9554,N_9133,N_8983);
nor U9555 (N_9555,N_9024,N_8946);
nor U9556 (N_9556,N_9039,N_8877);
nand U9557 (N_9557,N_9032,N_8839);
and U9558 (N_9558,N_9137,N_8988);
and U9559 (N_9559,N_9059,N_9029);
or U9560 (N_9560,N_8856,N_8989);
nor U9561 (N_9561,N_9090,N_8860);
or U9562 (N_9562,N_9118,N_8950);
and U9563 (N_9563,N_8873,N_9003);
and U9564 (N_9564,N_8805,N_8920);
xor U9565 (N_9565,N_9182,N_8970);
nand U9566 (N_9566,N_8914,N_8803);
nor U9567 (N_9567,N_8857,N_8838);
xnor U9568 (N_9568,N_8885,N_8976);
and U9569 (N_9569,N_8951,N_8873);
xnor U9570 (N_9570,N_8946,N_8878);
nor U9571 (N_9571,N_8842,N_9138);
nor U9572 (N_9572,N_9198,N_8860);
nand U9573 (N_9573,N_9153,N_8952);
and U9574 (N_9574,N_8977,N_8822);
xor U9575 (N_9575,N_9107,N_8900);
nand U9576 (N_9576,N_9135,N_8842);
xnor U9577 (N_9577,N_9039,N_9142);
xnor U9578 (N_9578,N_9051,N_9135);
nand U9579 (N_9579,N_9136,N_8952);
xnor U9580 (N_9580,N_8956,N_9128);
nor U9581 (N_9581,N_9008,N_8960);
nand U9582 (N_9582,N_9095,N_9150);
and U9583 (N_9583,N_8950,N_8930);
nand U9584 (N_9584,N_8802,N_8866);
nand U9585 (N_9585,N_8882,N_8905);
xor U9586 (N_9586,N_8936,N_8917);
nor U9587 (N_9587,N_8814,N_8914);
or U9588 (N_9588,N_8867,N_9180);
and U9589 (N_9589,N_8973,N_8943);
nand U9590 (N_9590,N_9040,N_9032);
or U9591 (N_9591,N_9156,N_9194);
nor U9592 (N_9592,N_8940,N_9039);
xnor U9593 (N_9593,N_8803,N_9108);
nand U9594 (N_9594,N_8928,N_8808);
and U9595 (N_9595,N_8942,N_8947);
nand U9596 (N_9596,N_8955,N_8999);
nand U9597 (N_9597,N_8963,N_8869);
nand U9598 (N_9598,N_9033,N_9177);
or U9599 (N_9599,N_9018,N_9025);
nand U9600 (N_9600,N_9582,N_9230);
xor U9601 (N_9601,N_9244,N_9229);
nor U9602 (N_9602,N_9518,N_9286);
and U9603 (N_9603,N_9246,N_9453);
nor U9604 (N_9604,N_9257,N_9381);
xor U9605 (N_9605,N_9420,N_9404);
nor U9606 (N_9606,N_9384,N_9468);
xnor U9607 (N_9607,N_9555,N_9342);
or U9608 (N_9608,N_9245,N_9587);
nand U9609 (N_9609,N_9238,N_9500);
nor U9610 (N_9610,N_9465,N_9336);
xnor U9611 (N_9611,N_9380,N_9217);
and U9612 (N_9612,N_9530,N_9202);
and U9613 (N_9613,N_9407,N_9337);
and U9614 (N_9614,N_9461,N_9451);
nor U9615 (N_9615,N_9452,N_9547);
xor U9616 (N_9616,N_9361,N_9548);
nand U9617 (N_9617,N_9466,N_9445);
and U9618 (N_9618,N_9426,N_9327);
nand U9619 (N_9619,N_9488,N_9273);
xnor U9620 (N_9620,N_9397,N_9583);
and U9621 (N_9621,N_9235,N_9302);
nor U9622 (N_9622,N_9540,N_9545);
or U9623 (N_9623,N_9522,N_9595);
or U9624 (N_9624,N_9262,N_9476);
nor U9625 (N_9625,N_9589,N_9306);
xnor U9626 (N_9626,N_9419,N_9362);
and U9627 (N_9627,N_9508,N_9299);
nand U9628 (N_9628,N_9350,N_9456);
nand U9629 (N_9629,N_9394,N_9467);
xnor U9630 (N_9630,N_9318,N_9218);
and U9631 (N_9631,N_9571,N_9275);
or U9632 (N_9632,N_9387,N_9501);
or U9633 (N_9633,N_9575,N_9359);
or U9634 (N_9634,N_9289,N_9374);
nand U9635 (N_9635,N_9566,N_9439);
or U9636 (N_9636,N_9416,N_9430);
nor U9637 (N_9637,N_9271,N_9509);
nor U9638 (N_9638,N_9484,N_9537);
nor U9639 (N_9639,N_9332,N_9323);
and U9640 (N_9640,N_9363,N_9528);
nand U9641 (N_9641,N_9523,N_9417);
xnor U9642 (N_9642,N_9499,N_9348);
nand U9643 (N_9643,N_9365,N_9581);
nand U9644 (N_9644,N_9267,N_9373);
nand U9645 (N_9645,N_9236,N_9534);
nand U9646 (N_9646,N_9335,N_9560);
nand U9647 (N_9647,N_9525,N_9242);
nor U9648 (N_9648,N_9584,N_9408);
nand U9649 (N_9649,N_9364,N_9211);
nand U9650 (N_9650,N_9446,N_9270);
xor U9651 (N_9651,N_9313,N_9551);
nand U9652 (N_9652,N_9305,N_9368);
and U9653 (N_9653,N_9248,N_9458);
nor U9654 (N_9654,N_9228,N_9303);
nor U9655 (N_9655,N_9330,N_9532);
nor U9656 (N_9656,N_9435,N_9564);
and U9657 (N_9657,N_9410,N_9539);
nor U9658 (N_9658,N_9475,N_9383);
nand U9659 (N_9659,N_9487,N_9317);
and U9660 (N_9660,N_9429,N_9207);
and U9661 (N_9661,N_9366,N_9599);
or U9662 (N_9662,N_9212,N_9382);
nor U9663 (N_9663,N_9208,N_9436);
and U9664 (N_9664,N_9215,N_9304);
xor U9665 (N_9665,N_9515,N_9514);
xor U9666 (N_9666,N_9422,N_9203);
nand U9667 (N_9667,N_9529,N_9541);
nand U9668 (N_9668,N_9353,N_9274);
xor U9669 (N_9669,N_9561,N_9240);
nand U9670 (N_9670,N_9320,N_9300);
nor U9671 (N_9671,N_9421,N_9285);
xnor U9672 (N_9672,N_9409,N_9224);
or U9673 (N_9673,N_9586,N_9553);
and U9674 (N_9674,N_9521,N_9495);
or U9675 (N_9675,N_9333,N_9249);
nand U9676 (N_9676,N_9315,N_9402);
nand U9677 (N_9677,N_9340,N_9276);
nand U9678 (N_9678,N_9434,N_9572);
and U9679 (N_9679,N_9231,N_9216);
nor U9680 (N_9680,N_9200,N_9293);
nand U9681 (N_9681,N_9570,N_9415);
and U9682 (N_9682,N_9550,N_9234);
and U9683 (N_9683,N_9290,N_9449);
xor U9684 (N_9684,N_9524,N_9357);
nand U9685 (N_9685,N_9232,N_9328);
and U9686 (N_9686,N_9369,N_9414);
xnor U9687 (N_9687,N_9279,N_9379);
xnor U9688 (N_9688,N_9356,N_9473);
or U9689 (N_9689,N_9204,N_9554);
and U9690 (N_9690,N_9574,N_9502);
and U9691 (N_9691,N_9527,N_9209);
nand U9692 (N_9692,N_9345,N_9351);
nand U9693 (N_9693,N_9423,N_9390);
or U9694 (N_9694,N_9296,N_9598);
and U9695 (N_9695,N_9510,N_9557);
or U9696 (N_9696,N_9597,N_9294);
or U9697 (N_9697,N_9210,N_9205);
nand U9698 (N_9698,N_9213,N_9310);
or U9699 (N_9699,N_9226,N_9386);
nor U9700 (N_9700,N_9312,N_9450);
nor U9701 (N_9701,N_9444,N_9459);
and U9702 (N_9702,N_9562,N_9341);
nand U9703 (N_9703,N_9399,N_9441);
xor U9704 (N_9704,N_9287,N_9371);
xor U9705 (N_9705,N_9385,N_9454);
nand U9706 (N_9706,N_9247,N_9580);
or U9707 (N_9707,N_9474,N_9222);
nand U9708 (N_9708,N_9505,N_9546);
xor U9709 (N_9709,N_9585,N_9412);
xnor U9710 (N_9710,N_9389,N_9406);
and U9711 (N_9711,N_9301,N_9490);
nor U9712 (N_9712,N_9588,N_9411);
xor U9713 (N_9713,N_9486,N_9259);
nor U9714 (N_9714,N_9201,N_9497);
xor U9715 (N_9715,N_9517,N_9269);
xor U9716 (N_9716,N_9513,N_9295);
nor U9717 (N_9717,N_9591,N_9573);
or U9718 (N_9718,N_9506,N_9291);
or U9719 (N_9719,N_9392,N_9214);
nand U9720 (N_9720,N_9442,N_9482);
nor U9721 (N_9721,N_9319,N_9349);
xor U9722 (N_9722,N_9241,N_9593);
nor U9723 (N_9723,N_9334,N_9258);
or U9724 (N_9724,N_9594,N_9526);
nor U9725 (N_9725,N_9280,N_9331);
and U9726 (N_9726,N_9481,N_9314);
nand U9727 (N_9727,N_9463,N_9223);
nor U9728 (N_9728,N_9346,N_9284);
or U9729 (N_9729,N_9489,N_9256);
or U9730 (N_9730,N_9512,N_9516);
or U9731 (N_9731,N_9272,N_9283);
and U9732 (N_9732,N_9533,N_9376);
nand U9733 (N_9733,N_9355,N_9316);
and U9734 (N_9734,N_9309,N_9478);
and U9735 (N_9735,N_9443,N_9344);
xor U9736 (N_9736,N_9297,N_9360);
nor U9737 (N_9737,N_9457,N_9464);
nand U9738 (N_9738,N_9396,N_9252);
nand U9739 (N_9739,N_9322,N_9233);
and U9740 (N_9740,N_9577,N_9221);
or U9741 (N_9741,N_9590,N_9326);
nor U9742 (N_9742,N_9433,N_9471);
nand U9743 (N_9743,N_9354,N_9496);
or U9744 (N_9744,N_9431,N_9579);
nor U9745 (N_9745,N_9455,N_9448);
nand U9746 (N_9746,N_9470,N_9325);
nand U9747 (N_9747,N_9329,N_9428);
or U9748 (N_9748,N_9219,N_9480);
nand U9749 (N_9749,N_9343,N_9485);
and U9750 (N_9750,N_9292,N_9375);
xnor U9751 (N_9751,N_9206,N_9403);
and U9752 (N_9752,N_9307,N_9378);
nand U9753 (N_9753,N_9298,N_9264);
nor U9754 (N_9754,N_9578,N_9388);
and U9755 (N_9755,N_9358,N_9479);
nand U9756 (N_9756,N_9253,N_9543);
xor U9757 (N_9757,N_9596,N_9437);
nor U9758 (N_9758,N_9237,N_9282);
xor U9759 (N_9759,N_9367,N_9401);
xor U9760 (N_9760,N_9372,N_9432);
and U9761 (N_9761,N_9427,N_9398);
nand U9762 (N_9762,N_9549,N_9251);
nand U9763 (N_9763,N_9592,N_9544);
nor U9764 (N_9764,N_9542,N_9324);
nand U9765 (N_9765,N_9552,N_9535);
and U9766 (N_9766,N_9483,N_9576);
xnor U9767 (N_9767,N_9347,N_9492);
and U9768 (N_9768,N_9377,N_9556);
nor U9769 (N_9769,N_9277,N_9393);
and U9770 (N_9770,N_9261,N_9503);
nand U9771 (N_9771,N_9268,N_9405);
nor U9772 (N_9772,N_9227,N_9425);
xor U9773 (N_9773,N_9338,N_9472);
or U9774 (N_9774,N_9447,N_9493);
nand U9775 (N_9775,N_9263,N_9536);
or U9776 (N_9776,N_9440,N_9568);
nor U9777 (N_9777,N_9477,N_9288);
and U9778 (N_9778,N_9559,N_9494);
nand U9779 (N_9779,N_9563,N_9260);
nand U9780 (N_9780,N_9531,N_9413);
nand U9781 (N_9781,N_9569,N_9400);
nand U9782 (N_9782,N_9438,N_9519);
nand U9783 (N_9783,N_9220,N_9538);
xnor U9784 (N_9784,N_9255,N_9491);
nor U9785 (N_9785,N_9462,N_9339);
xnor U9786 (N_9786,N_9239,N_9370);
nor U9787 (N_9787,N_9498,N_9504);
and U9788 (N_9788,N_9321,N_9507);
nand U9789 (N_9789,N_9308,N_9418);
nand U9790 (N_9790,N_9225,N_9352);
and U9791 (N_9791,N_9520,N_9391);
nand U9792 (N_9792,N_9567,N_9424);
nand U9793 (N_9793,N_9281,N_9278);
or U9794 (N_9794,N_9311,N_9243);
and U9795 (N_9795,N_9395,N_9265);
or U9796 (N_9796,N_9511,N_9266);
xnor U9797 (N_9797,N_9565,N_9250);
nand U9798 (N_9798,N_9469,N_9460);
nand U9799 (N_9799,N_9254,N_9558);
nor U9800 (N_9800,N_9274,N_9488);
xor U9801 (N_9801,N_9233,N_9425);
and U9802 (N_9802,N_9476,N_9437);
or U9803 (N_9803,N_9433,N_9317);
nor U9804 (N_9804,N_9578,N_9396);
nand U9805 (N_9805,N_9524,N_9325);
nor U9806 (N_9806,N_9263,N_9367);
or U9807 (N_9807,N_9396,N_9475);
nand U9808 (N_9808,N_9244,N_9369);
nand U9809 (N_9809,N_9399,N_9430);
nand U9810 (N_9810,N_9491,N_9404);
xnor U9811 (N_9811,N_9504,N_9425);
nand U9812 (N_9812,N_9288,N_9495);
or U9813 (N_9813,N_9273,N_9565);
xnor U9814 (N_9814,N_9488,N_9314);
and U9815 (N_9815,N_9406,N_9363);
or U9816 (N_9816,N_9354,N_9403);
nand U9817 (N_9817,N_9310,N_9575);
or U9818 (N_9818,N_9464,N_9268);
and U9819 (N_9819,N_9411,N_9424);
and U9820 (N_9820,N_9433,N_9459);
or U9821 (N_9821,N_9383,N_9225);
and U9822 (N_9822,N_9503,N_9549);
or U9823 (N_9823,N_9521,N_9467);
or U9824 (N_9824,N_9423,N_9598);
and U9825 (N_9825,N_9376,N_9587);
and U9826 (N_9826,N_9539,N_9382);
and U9827 (N_9827,N_9444,N_9505);
xnor U9828 (N_9828,N_9234,N_9515);
or U9829 (N_9829,N_9461,N_9556);
xnor U9830 (N_9830,N_9408,N_9303);
or U9831 (N_9831,N_9412,N_9540);
and U9832 (N_9832,N_9398,N_9499);
xor U9833 (N_9833,N_9348,N_9460);
or U9834 (N_9834,N_9290,N_9389);
nor U9835 (N_9835,N_9309,N_9502);
and U9836 (N_9836,N_9379,N_9465);
nand U9837 (N_9837,N_9301,N_9576);
xor U9838 (N_9838,N_9213,N_9296);
nand U9839 (N_9839,N_9295,N_9569);
and U9840 (N_9840,N_9377,N_9405);
nand U9841 (N_9841,N_9246,N_9308);
nand U9842 (N_9842,N_9437,N_9384);
nand U9843 (N_9843,N_9599,N_9227);
nand U9844 (N_9844,N_9457,N_9285);
nor U9845 (N_9845,N_9235,N_9253);
nand U9846 (N_9846,N_9293,N_9259);
and U9847 (N_9847,N_9390,N_9484);
and U9848 (N_9848,N_9593,N_9222);
and U9849 (N_9849,N_9240,N_9352);
xor U9850 (N_9850,N_9592,N_9455);
and U9851 (N_9851,N_9235,N_9210);
and U9852 (N_9852,N_9277,N_9562);
and U9853 (N_9853,N_9383,N_9422);
xnor U9854 (N_9854,N_9436,N_9319);
xor U9855 (N_9855,N_9344,N_9293);
or U9856 (N_9856,N_9248,N_9500);
and U9857 (N_9857,N_9240,N_9222);
xnor U9858 (N_9858,N_9306,N_9517);
nand U9859 (N_9859,N_9394,N_9542);
and U9860 (N_9860,N_9303,N_9599);
nand U9861 (N_9861,N_9414,N_9301);
nand U9862 (N_9862,N_9428,N_9441);
or U9863 (N_9863,N_9522,N_9437);
nand U9864 (N_9864,N_9341,N_9285);
and U9865 (N_9865,N_9581,N_9480);
nand U9866 (N_9866,N_9340,N_9444);
nor U9867 (N_9867,N_9359,N_9263);
and U9868 (N_9868,N_9531,N_9324);
and U9869 (N_9869,N_9518,N_9453);
nand U9870 (N_9870,N_9565,N_9212);
nand U9871 (N_9871,N_9342,N_9276);
nor U9872 (N_9872,N_9506,N_9512);
nor U9873 (N_9873,N_9580,N_9278);
nor U9874 (N_9874,N_9290,N_9516);
and U9875 (N_9875,N_9414,N_9568);
xnor U9876 (N_9876,N_9378,N_9547);
xor U9877 (N_9877,N_9427,N_9364);
nand U9878 (N_9878,N_9260,N_9236);
nand U9879 (N_9879,N_9530,N_9264);
and U9880 (N_9880,N_9591,N_9299);
or U9881 (N_9881,N_9597,N_9466);
xor U9882 (N_9882,N_9287,N_9510);
and U9883 (N_9883,N_9528,N_9399);
xor U9884 (N_9884,N_9546,N_9243);
nand U9885 (N_9885,N_9494,N_9294);
nor U9886 (N_9886,N_9514,N_9469);
and U9887 (N_9887,N_9406,N_9403);
and U9888 (N_9888,N_9239,N_9537);
or U9889 (N_9889,N_9225,N_9544);
and U9890 (N_9890,N_9468,N_9497);
and U9891 (N_9891,N_9594,N_9482);
xnor U9892 (N_9892,N_9543,N_9547);
xor U9893 (N_9893,N_9515,N_9344);
nand U9894 (N_9894,N_9205,N_9309);
nand U9895 (N_9895,N_9226,N_9242);
nor U9896 (N_9896,N_9514,N_9262);
and U9897 (N_9897,N_9520,N_9453);
and U9898 (N_9898,N_9538,N_9554);
or U9899 (N_9899,N_9259,N_9349);
nor U9900 (N_9900,N_9535,N_9566);
and U9901 (N_9901,N_9381,N_9321);
nor U9902 (N_9902,N_9394,N_9378);
nor U9903 (N_9903,N_9420,N_9474);
xor U9904 (N_9904,N_9533,N_9574);
and U9905 (N_9905,N_9560,N_9518);
nand U9906 (N_9906,N_9513,N_9496);
or U9907 (N_9907,N_9478,N_9304);
nand U9908 (N_9908,N_9442,N_9420);
nand U9909 (N_9909,N_9394,N_9502);
nand U9910 (N_9910,N_9352,N_9480);
or U9911 (N_9911,N_9280,N_9569);
and U9912 (N_9912,N_9451,N_9267);
nor U9913 (N_9913,N_9221,N_9225);
and U9914 (N_9914,N_9326,N_9345);
xnor U9915 (N_9915,N_9598,N_9327);
or U9916 (N_9916,N_9528,N_9348);
and U9917 (N_9917,N_9496,N_9200);
nor U9918 (N_9918,N_9313,N_9588);
and U9919 (N_9919,N_9502,N_9513);
xor U9920 (N_9920,N_9550,N_9201);
xor U9921 (N_9921,N_9545,N_9361);
or U9922 (N_9922,N_9502,N_9549);
nor U9923 (N_9923,N_9340,N_9533);
and U9924 (N_9924,N_9371,N_9365);
nor U9925 (N_9925,N_9326,N_9381);
and U9926 (N_9926,N_9397,N_9501);
xor U9927 (N_9927,N_9349,N_9418);
or U9928 (N_9928,N_9249,N_9334);
nand U9929 (N_9929,N_9345,N_9363);
or U9930 (N_9930,N_9306,N_9477);
and U9931 (N_9931,N_9312,N_9275);
nand U9932 (N_9932,N_9217,N_9205);
xor U9933 (N_9933,N_9404,N_9575);
or U9934 (N_9934,N_9250,N_9482);
xnor U9935 (N_9935,N_9377,N_9262);
xnor U9936 (N_9936,N_9579,N_9514);
nor U9937 (N_9937,N_9443,N_9411);
nor U9938 (N_9938,N_9360,N_9316);
nor U9939 (N_9939,N_9519,N_9554);
nor U9940 (N_9940,N_9388,N_9306);
or U9941 (N_9941,N_9287,N_9545);
or U9942 (N_9942,N_9537,N_9345);
or U9943 (N_9943,N_9538,N_9391);
xnor U9944 (N_9944,N_9308,N_9478);
xor U9945 (N_9945,N_9367,N_9390);
nand U9946 (N_9946,N_9299,N_9421);
nor U9947 (N_9947,N_9340,N_9478);
nand U9948 (N_9948,N_9458,N_9226);
xor U9949 (N_9949,N_9388,N_9392);
nor U9950 (N_9950,N_9373,N_9307);
xor U9951 (N_9951,N_9521,N_9237);
nand U9952 (N_9952,N_9531,N_9254);
nand U9953 (N_9953,N_9477,N_9386);
or U9954 (N_9954,N_9248,N_9589);
and U9955 (N_9955,N_9580,N_9537);
nor U9956 (N_9956,N_9391,N_9263);
nand U9957 (N_9957,N_9501,N_9550);
nand U9958 (N_9958,N_9438,N_9216);
xor U9959 (N_9959,N_9550,N_9484);
xor U9960 (N_9960,N_9360,N_9368);
nor U9961 (N_9961,N_9473,N_9491);
and U9962 (N_9962,N_9572,N_9547);
xnor U9963 (N_9963,N_9524,N_9217);
and U9964 (N_9964,N_9585,N_9524);
nand U9965 (N_9965,N_9253,N_9213);
nor U9966 (N_9966,N_9305,N_9578);
nor U9967 (N_9967,N_9555,N_9539);
or U9968 (N_9968,N_9301,N_9523);
xor U9969 (N_9969,N_9472,N_9467);
xor U9970 (N_9970,N_9508,N_9347);
nor U9971 (N_9971,N_9425,N_9477);
or U9972 (N_9972,N_9435,N_9434);
or U9973 (N_9973,N_9452,N_9579);
or U9974 (N_9974,N_9466,N_9440);
nand U9975 (N_9975,N_9581,N_9299);
and U9976 (N_9976,N_9467,N_9209);
or U9977 (N_9977,N_9218,N_9376);
nor U9978 (N_9978,N_9334,N_9594);
or U9979 (N_9979,N_9562,N_9355);
and U9980 (N_9980,N_9249,N_9487);
nor U9981 (N_9981,N_9301,N_9342);
nor U9982 (N_9982,N_9277,N_9422);
nand U9983 (N_9983,N_9459,N_9588);
nor U9984 (N_9984,N_9528,N_9361);
and U9985 (N_9985,N_9444,N_9428);
and U9986 (N_9986,N_9597,N_9397);
xor U9987 (N_9987,N_9555,N_9215);
or U9988 (N_9988,N_9421,N_9311);
nand U9989 (N_9989,N_9213,N_9383);
or U9990 (N_9990,N_9561,N_9223);
or U9991 (N_9991,N_9581,N_9270);
xnor U9992 (N_9992,N_9284,N_9310);
xnor U9993 (N_9993,N_9279,N_9266);
or U9994 (N_9994,N_9380,N_9473);
xnor U9995 (N_9995,N_9340,N_9569);
nor U9996 (N_9996,N_9550,N_9518);
xnor U9997 (N_9997,N_9350,N_9404);
nand U9998 (N_9998,N_9435,N_9310);
xor U9999 (N_9999,N_9256,N_9571);
xnor U10000 (N_10000,N_9733,N_9860);
xor U10001 (N_10001,N_9781,N_9937);
and U10002 (N_10002,N_9710,N_9983);
or U10003 (N_10003,N_9763,N_9767);
or U10004 (N_10004,N_9700,N_9955);
xor U10005 (N_10005,N_9887,N_9968);
nand U10006 (N_10006,N_9984,N_9689);
xor U10007 (N_10007,N_9637,N_9999);
or U10008 (N_10008,N_9635,N_9948);
or U10009 (N_10009,N_9656,N_9705);
nor U10010 (N_10010,N_9876,N_9838);
or U10011 (N_10011,N_9821,N_9819);
and U10012 (N_10012,N_9632,N_9771);
xnor U10013 (N_10013,N_9619,N_9663);
nand U10014 (N_10014,N_9963,N_9988);
nor U10015 (N_10015,N_9752,N_9659);
and U10016 (N_10016,N_9629,N_9929);
nand U10017 (N_10017,N_9823,N_9882);
and U10018 (N_10018,N_9897,N_9600);
xnor U10019 (N_10019,N_9861,N_9869);
or U10020 (N_10020,N_9920,N_9908);
xnor U10021 (N_10021,N_9830,N_9986);
nand U10022 (N_10022,N_9901,N_9972);
nor U10023 (N_10023,N_9630,N_9636);
nand U10024 (N_10024,N_9910,N_9765);
or U10025 (N_10025,N_9746,N_9673);
nand U10026 (N_10026,N_9660,N_9906);
nand U10027 (N_10027,N_9985,N_9727);
nand U10028 (N_10028,N_9745,N_9607);
nor U10029 (N_10029,N_9835,N_9758);
nand U10030 (N_10030,N_9616,N_9889);
or U10031 (N_10031,N_9777,N_9898);
and U10032 (N_10032,N_9859,N_9842);
xnor U10033 (N_10033,N_9828,N_9759);
nand U10034 (N_10034,N_9793,N_9631);
xor U10035 (N_10035,N_9831,N_9739);
xor U10036 (N_10036,N_9686,N_9750);
nor U10037 (N_10037,N_9715,N_9854);
or U10038 (N_10038,N_9847,N_9627);
nor U10039 (N_10039,N_9696,N_9722);
nor U10040 (N_10040,N_9928,N_9974);
xnor U10041 (N_10041,N_9617,N_9711);
nor U10042 (N_10042,N_9971,N_9792);
nor U10043 (N_10043,N_9824,N_9825);
xnor U10044 (N_10044,N_9601,N_9729);
or U10045 (N_10045,N_9938,N_9879);
nor U10046 (N_10046,N_9959,N_9678);
nand U10047 (N_10047,N_9926,N_9618);
and U10048 (N_10048,N_9837,N_9858);
and U10049 (N_10049,N_9989,N_9977);
nand U10050 (N_10050,N_9909,N_9975);
or U10051 (N_10051,N_9864,N_9947);
xnor U10052 (N_10052,N_9813,N_9776);
xor U10053 (N_10053,N_9878,N_9918);
and U10054 (N_10054,N_9851,N_9726);
xor U10055 (N_10055,N_9826,N_9880);
xnor U10056 (N_10056,N_9907,N_9679);
nand U10057 (N_10057,N_9870,N_9902);
xnor U10058 (N_10058,N_9704,N_9736);
or U10059 (N_10059,N_9961,N_9694);
or U10060 (N_10060,N_9766,N_9982);
nand U10061 (N_10061,N_9890,N_9872);
nand U10062 (N_10062,N_9784,N_9891);
or U10063 (N_10063,N_9931,N_9874);
xnor U10064 (N_10064,N_9922,N_9973);
xnor U10065 (N_10065,N_9956,N_9788);
or U10066 (N_10066,N_9952,N_9677);
nand U10067 (N_10067,N_9987,N_9644);
nor U10068 (N_10068,N_9743,N_9625);
or U10069 (N_10069,N_9899,N_9932);
xor U10070 (N_10070,N_9894,N_9723);
or U10071 (N_10071,N_9643,N_9693);
nand U10072 (N_10072,N_9939,N_9810);
or U10073 (N_10073,N_9913,N_9954);
xor U10074 (N_10074,N_9747,N_9805);
xnor U10075 (N_10075,N_9875,N_9709);
nor U10076 (N_10076,N_9642,N_9769);
xnor U10077 (N_10077,N_9681,N_9732);
nor U10078 (N_10078,N_9964,N_9841);
xnor U10079 (N_10079,N_9791,N_9924);
or U10080 (N_10080,N_9978,N_9967);
nand U10081 (N_10081,N_9900,N_9603);
nor U10082 (N_10082,N_9935,N_9740);
nor U10083 (N_10083,N_9965,N_9981);
and U10084 (N_10084,N_9707,N_9728);
and U10085 (N_10085,N_9957,N_9685);
and U10086 (N_10086,N_9998,N_9903);
nor U10087 (N_10087,N_9628,N_9741);
xnor U10088 (N_10088,N_9785,N_9773);
nand U10089 (N_10089,N_9832,N_9818);
xor U10090 (N_10090,N_9936,N_9754);
and U10091 (N_10091,N_9633,N_9916);
xor U10092 (N_10092,N_9638,N_9695);
or U10093 (N_10093,N_9812,N_9645);
nor U10094 (N_10094,N_9829,N_9782);
or U10095 (N_10095,N_9698,N_9666);
nand U10096 (N_10096,N_9995,N_9713);
and U10097 (N_10097,N_9647,N_9863);
nand U10098 (N_10098,N_9654,N_9760);
and U10099 (N_10099,N_9667,N_9622);
xnor U10100 (N_10100,N_9856,N_9775);
nand U10101 (N_10101,N_9702,N_9953);
xor U10102 (N_10102,N_9868,N_9850);
or U10103 (N_10103,N_9669,N_9640);
and U10104 (N_10104,N_9845,N_9650);
and U10105 (N_10105,N_9933,N_9811);
or U10106 (N_10106,N_9990,N_9881);
nand U10107 (N_10107,N_9605,N_9606);
and U10108 (N_10108,N_9840,N_9892);
or U10109 (N_10109,N_9621,N_9714);
nor U10110 (N_10110,N_9701,N_9820);
nand U10111 (N_10111,N_9712,N_9786);
nand U10112 (N_10112,N_9996,N_9944);
nor U10113 (N_10113,N_9783,N_9688);
xnor U10114 (N_10114,N_9737,N_9853);
nor U10115 (N_10115,N_9787,N_9799);
and U10116 (N_10116,N_9814,N_9646);
xor U10117 (N_10117,N_9604,N_9843);
nand U10118 (N_10118,N_9921,N_9833);
nand U10119 (N_10119,N_9839,N_9718);
and U10120 (N_10120,N_9960,N_9762);
xnor U10121 (N_10121,N_9730,N_9896);
nor U10122 (N_10122,N_9761,N_9676);
nand U10123 (N_10123,N_9862,N_9849);
or U10124 (N_10124,N_9612,N_9690);
and U10125 (N_10125,N_9958,N_9724);
nor U10126 (N_10126,N_9925,N_9940);
or U10127 (N_10127,N_9768,N_9742);
xnor U10128 (N_10128,N_9735,N_9962);
nand U10129 (N_10129,N_9668,N_9753);
nand U10130 (N_10130,N_9795,N_9914);
or U10131 (N_10131,N_9803,N_9992);
nor U10132 (N_10132,N_9751,N_9721);
nand U10133 (N_10133,N_9731,N_9934);
nand U10134 (N_10134,N_9748,N_9883);
nand U10135 (N_10135,N_9664,N_9822);
or U10136 (N_10136,N_9893,N_9764);
and U10137 (N_10137,N_9991,N_9969);
and U10138 (N_10138,N_9871,N_9915);
or U10139 (N_10139,N_9661,N_9602);
or U10140 (N_10140,N_9846,N_9855);
nand U10141 (N_10141,N_9634,N_9683);
and U10142 (N_10142,N_9888,N_9623);
nand U10143 (N_10143,N_9873,N_9717);
and U10144 (N_10144,N_9834,N_9993);
and U10145 (N_10145,N_9755,N_9895);
nand U10146 (N_10146,N_9657,N_9778);
or U10147 (N_10147,N_9798,N_9772);
and U10148 (N_10148,N_9946,N_9716);
nor U10149 (N_10149,N_9662,N_9749);
and U10150 (N_10150,N_9942,N_9608);
nand U10151 (N_10151,N_9951,N_9796);
xor U10152 (N_10152,N_9919,N_9658);
xnor U10153 (N_10153,N_9697,N_9912);
nand U10154 (N_10154,N_9852,N_9884);
nand U10155 (N_10155,N_9844,N_9980);
or U10156 (N_10156,N_9774,N_9809);
and U10157 (N_10157,N_9789,N_9665);
and U10158 (N_10158,N_9649,N_9651);
or U10159 (N_10159,N_9719,N_9807);
or U10160 (N_10160,N_9615,N_9613);
or U10161 (N_10161,N_9780,N_9744);
nor U10162 (N_10162,N_9610,N_9738);
and U10163 (N_10163,N_9725,N_9949);
nand U10164 (N_10164,N_9997,N_9917);
or U10165 (N_10165,N_9866,N_9757);
and U10166 (N_10166,N_9609,N_9671);
nor U10167 (N_10167,N_9779,N_9923);
xor U10168 (N_10168,N_9927,N_9684);
nor U10169 (N_10169,N_9804,N_9652);
nand U10170 (N_10170,N_9943,N_9808);
and U10171 (N_10171,N_9687,N_9905);
xor U10172 (N_10172,N_9970,N_9801);
nor U10173 (N_10173,N_9857,N_9626);
and U10174 (N_10174,N_9800,N_9836);
and U10175 (N_10175,N_9670,N_9682);
xor U10176 (N_10176,N_9911,N_9930);
xor U10177 (N_10177,N_9790,N_9877);
or U10178 (N_10178,N_9641,N_9806);
nor U10179 (N_10179,N_9706,N_9848);
or U10180 (N_10180,N_9966,N_9941);
and U10181 (N_10181,N_9692,N_9620);
xnor U10182 (N_10182,N_9885,N_9611);
nand U10183 (N_10183,N_9802,N_9797);
xor U10184 (N_10184,N_9708,N_9720);
nand U10185 (N_10185,N_9653,N_9827);
or U10186 (N_10186,N_9794,N_9675);
or U10187 (N_10187,N_9994,N_9703);
or U10188 (N_10188,N_9624,N_9655);
or U10189 (N_10189,N_9648,N_9816);
nand U10190 (N_10190,N_9672,N_9886);
and U10191 (N_10191,N_9945,N_9674);
or U10192 (N_10192,N_9691,N_9770);
nand U10193 (N_10193,N_9979,N_9867);
and U10194 (N_10194,N_9865,N_9699);
and U10195 (N_10195,N_9680,N_9815);
nor U10196 (N_10196,N_9976,N_9817);
xor U10197 (N_10197,N_9734,N_9756);
nand U10198 (N_10198,N_9950,N_9904);
xor U10199 (N_10199,N_9639,N_9614);
or U10200 (N_10200,N_9955,N_9631);
xnor U10201 (N_10201,N_9922,N_9951);
nand U10202 (N_10202,N_9979,N_9875);
nand U10203 (N_10203,N_9706,N_9943);
nand U10204 (N_10204,N_9948,N_9713);
nand U10205 (N_10205,N_9998,N_9904);
nand U10206 (N_10206,N_9677,N_9805);
nor U10207 (N_10207,N_9954,N_9931);
or U10208 (N_10208,N_9896,N_9643);
nand U10209 (N_10209,N_9740,N_9647);
nand U10210 (N_10210,N_9788,N_9604);
xnor U10211 (N_10211,N_9801,N_9862);
nor U10212 (N_10212,N_9837,N_9995);
xor U10213 (N_10213,N_9603,N_9919);
or U10214 (N_10214,N_9672,N_9604);
nor U10215 (N_10215,N_9917,N_9726);
or U10216 (N_10216,N_9789,N_9825);
nor U10217 (N_10217,N_9909,N_9876);
or U10218 (N_10218,N_9794,N_9716);
nor U10219 (N_10219,N_9973,N_9837);
xor U10220 (N_10220,N_9867,N_9802);
nand U10221 (N_10221,N_9961,N_9622);
and U10222 (N_10222,N_9624,N_9685);
nor U10223 (N_10223,N_9906,N_9772);
nor U10224 (N_10224,N_9887,N_9919);
nand U10225 (N_10225,N_9858,N_9901);
nand U10226 (N_10226,N_9847,N_9975);
nand U10227 (N_10227,N_9876,N_9644);
or U10228 (N_10228,N_9806,N_9933);
xor U10229 (N_10229,N_9915,N_9931);
xnor U10230 (N_10230,N_9792,N_9610);
nand U10231 (N_10231,N_9882,N_9781);
nor U10232 (N_10232,N_9894,N_9879);
and U10233 (N_10233,N_9928,N_9606);
or U10234 (N_10234,N_9655,N_9832);
and U10235 (N_10235,N_9648,N_9766);
nor U10236 (N_10236,N_9960,N_9688);
nand U10237 (N_10237,N_9678,N_9795);
or U10238 (N_10238,N_9949,N_9673);
and U10239 (N_10239,N_9998,N_9659);
or U10240 (N_10240,N_9630,N_9958);
or U10241 (N_10241,N_9618,N_9709);
xor U10242 (N_10242,N_9874,N_9674);
and U10243 (N_10243,N_9793,N_9708);
or U10244 (N_10244,N_9873,N_9814);
nand U10245 (N_10245,N_9989,N_9839);
nor U10246 (N_10246,N_9939,N_9883);
and U10247 (N_10247,N_9906,N_9755);
or U10248 (N_10248,N_9771,N_9606);
nand U10249 (N_10249,N_9848,N_9762);
and U10250 (N_10250,N_9824,N_9944);
xor U10251 (N_10251,N_9614,N_9691);
or U10252 (N_10252,N_9901,N_9836);
or U10253 (N_10253,N_9603,N_9682);
nand U10254 (N_10254,N_9804,N_9633);
xnor U10255 (N_10255,N_9925,N_9687);
nor U10256 (N_10256,N_9778,N_9962);
and U10257 (N_10257,N_9638,N_9601);
nor U10258 (N_10258,N_9628,N_9867);
xnor U10259 (N_10259,N_9790,N_9636);
nor U10260 (N_10260,N_9634,N_9878);
and U10261 (N_10261,N_9736,N_9899);
nand U10262 (N_10262,N_9992,N_9650);
nand U10263 (N_10263,N_9611,N_9860);
xnor U10264 (N_10264,N_9697,N_9705);
or U10265 (N_10265,N_9774,N_9715);
nand U10266 (N_10266,N_9945,N_9614);
or U10267 (N_10267,N_9958,N_9939);
nand U10268 (N_10268,N_9638,N_9648);
and U10269 (N_10269,N_9968,N_9771);
nand U10270 (N_10270,N_9970,N_9764);
nand U10271 (N_10271,N_9820,N_9688);
nand U10272 (N_10272,N_9678,N_9869);
nand U10273 (N_10273,N_9704,N_9884);
and U10274 (N_10274,N_9659,N_9670);
nor U10275 (N_10275,N_9765,N_9934);
nand U10276 (N_10276,N_9719,N_9885);
nor U10277 (N_10277,N_9710,N_9790);
or U10278 (N_10278,N_9809,N_9686);
xor U10279 (N_10279,N_9896,N_9874);
xnor U10280 (N_10280,N_9848,N_9698);
nand U10281 (N_10281,N_9729,N_9838);
xnor U10282 (N_10282,N_9707,N_9958);
and U10283 (N_10283,N_9863,N_9750);
nand U10284 (N_10284,N_9921,N_9819);
nand U10285 (N_10285,N_9860,N_9639);
xor U10286 (N_10286,N_9757,N_9840);
nand U10287 (N_10287,N_9963,N_9770);
nand U10288 (N_10288,N_9845,N_9776);
or U10289 (N_10289,N_9859,N_9943);
or U10290 (N_10290,N_9825,N_9916);
and U10291 (N_10291,N_9902,N_9600);
xnor U10292 (N_10292,N_9780,N_9987);
nand U10293 (N_10293,N_9874,N_9773);
and U10294 (N_10294,N_9815,N_9915);
and U10295 (N_10295,N_9821,N_9666);
nor U10296 (N_10296,N_9888,N_9944);
or U10297 (N_10297,N_9987,N_9830);
nand U10298 (N_10298,N_9700,N_9827);
and U10299 (N_10299,N_9962,N_9948);
nand U10300 (N_10300,N_9923,N_9660);
and U10301 (N_10301,N_9825,N_9922);
xnor U10302 (N_10302,N_9875,N_9935);
nand U10303 (N_10303,N_9731,N_9709);
and U10304 (N_10304,N_9859,N_9909);
xor U10305 (N_10305,N_9632,N_9728);
and U10306 (N_10306,N_9739,N_9887);
nand U10307 (N_10307,N_9933,N_9725);
xnor U10308 (N_10308,N_9822,N_9849);
nand U10309 (N_10309,N_9758,N_9737);
xor U10310 (N_10310,N_9801,N_9622);
nor U10311 (N_10311,N_9823,N_9698);
xnor U10312 (N_10312,N_9606,N_9779);
nor U10313 (N_10313,N_9914,N_9982);
or U10314 (N_10314,N_9654,N_9600);
xnor U10315 (N_10315,N_9827,N_9626);
or U10316 (N_10316,N_9854,N_9685);
or U10317 (N_10317,N_9824,N_9864);
or U10318 (N_10318,N_9698,N_9665);
or U10319 (N_10319,N_9859,N_9606);
nor U10320 (N_10320,N_9973,N_9767);
and U10321 (N_10321,N_9984,N_9651);
nor U10322 (N_10322,N_9789,N_9953);
and U10323 (N_10323,N_9909,N_9946);
or U10324 (N_10324,N_9703,N_9943);
and U10325 (N_10325,N_9715,N_9751);
and U10326 (N_10326,N_9808,N_9743);
or U10327 (N_10327,N_9942,N_9861);
nand U10328 (N_10328,N_9711,N_9762);
or U10329 (N_10329,N_9642,N_9970);
or U10330 (N_10330,N_9956,N_9973);
xnor U10331 (N_10331,N_9650,N_9825);
xnor U10332 (N_10332,N_9702,N_9668);
nor U10333 (N_10333,N_9700,N_9933);
or U10334 (N_10334,N_9785,N_9901);
and U10335 (N_10335,N_9604,N_9668);
or U10336 (N_10336,N_9654,N_9888);
xnor U10337 (N_10337,N_9652,N_9871);
nor U10338 (N_10338,N_9783,N_9860);
and U10339 (N_10339,N_9887,N_9712);
or U10340 (N_10340,N_9617,N_9972);
or U10341 (N_10341,N_9964,N_9784);
xor U10342 (N_10342,N_9890,N_9851);
nor U10343 (N_10343,N_9792,N_9690);
nand U10344 (N_10344,N_9796,N_9706);
xor U10345 (N_10345,N_9677,N_9774);
and U10346 (N_10346,N_9698,N_9759);
xnor U10347 (N_10347,N_9794,N_9910);
xnor U10348 (N_10348,N_9704,N_9793);
nor U10349 (N_10349,N_9989,N_9656);
or U10350 (N_10350,N_9752,N_9776);
or U10351 (N_10351,N_9823,N_9770);
or U10352 (N_10352,N_9714,N_9944);
nand U10353 (N_10353,N_9957,N_9836);
nor U10354 (N_10354,N_9927,N_9635);
nand U10355 (N_10355,N_9946,N_9744);
nand U10356 (N_10356,N_9993,N_9790);
and U10357 (N_10357,N_9905,N_9949);
nor U10358 (N_10358,N_9938,N_9608);
nor U10359 (N_10359,N_9986,N_9752);
or U10360 (N_10360,N_9983,N_9939);
and U10361 (N_10361,N_9603,N_9871);
nand U10362 (N_10362,N_9627,N_9795);
xor U10363 (N_10363,N_9850,N_9771);
and U10364 (N_10364,N_9738,N_9638);
xor U10365 (N_10365,N_9830,N_9627);
nand U10366 (N_10366,N_9939,N_9796);
and U10367 (N_10367,N_9954,N_9656);
or U10368 (N_10368,N_9829,N_9622);
xor U10369 (N_10369,N_9863,N_9861);
nor U10370 (N_10370,N_9801,N_9831);
and U10371 (N_10371,N_9615,N_9691);
and U10372 (N_10372,N_9883,N_9964);
nor U10373 (N_10373,N_9949,N_9682);
nor U10374 (N_10374,N_9836,N_9668);
and U10375 (N_10375,N_9643,N_9992);
or U10376 (N_10376,N_9634,N_9651);
or U10377 (N_10377,N_9684,N_9876);
nand U10378 (N_10378,N_9600,N_9911);
nor U10379 (N_10379,N_9754,N_9899);
nor U10380 (N_10380,N_9779,N_9933);
and U10381 (N_10381,N_9738,N_9617);
xor U10382 (N_10382,N_9880,N_9971);
and U10383 (N_10383,N_9659,N_9920);
or U10384 (N_10384,N_9896,N_9803);
nand U10385 (N_10385,N_9873,N_9723);
and U10386 (N_10386,N_9612,N_9945);
nand U10387 (N_10387,N_9963,N_9992);
and U10388 (N_10388,N_9998,N_9815);
and U10389 (N_10389,N_9999,N_9948);
and U10390 (N_10390,N_9934,N_9932);
nand U10391 (N_10391,N_9816,N_9748);
nand U10392 (N_10392,N_9626,N_9980);
or U10393 (N_10393,N_9790,N_9851);
xnor U10394 (N_10394,N_9648,N_9905);
or U10395 (N_10395,N_9790,N_9671);
nor U10396 (N_10396,N_9649,N_9628);
and U10397 (N_10397,N_9793,N_9895);
nor U10398 (N_10398,N_9601,N_9634);
nor U10399 (N_10399,N_9959,N_9680);
or U10400 (N_10400,N_10208,N_10362);
or U10401 (N_10401,N_10165,N_10129);
xor U10402 (N_10402,N_10137,N_10178);
xnor U10403 (N_10403,N_10278,N_10309);
xnor U10404 (N_10404,N_10265,N_10025);
or U10405 (N_10405,N_10079,N_10334);
nand U10406 (N_10406,N_10007,N_10193);
nand U10407 (N_10407,N_10160,N_10042);
and U10408 (N_10408,N_10266,N_10071);
and U10409 (N_10409,N_10107,N_10354);
or U10410 (N_10410,N_10269,N_10228);
nor U10411 (N_10411,N_10171,N_10324);
or U10412 (N_10412,N_10183,N_10316);
and U10413 (N_10413,N_10172,N_10031);
nor U10414 (N_10414,N_10388,N_10088);
nor U10415 (N_10415,N_10290,N_10030);
xnor U10416 (N_10416,N_10289,N_10006);
xor U10417 (N_10417,N_10340,N_10126);
and U10418 (N_10418,N_10268,N_10026);
nand U10419 (N_10419,N_10398,N_10052);
and U10420 (N_10420,N_10124,N_10242);
xnor U10421 (N_10421,N_10229,N_10247);
xor U10422 (N_10422,N_10190,N_10188);
nor U10423 (N_10423,N_10373,N_10147);
nand U10424 (N_10424,N_10196,N_10067);
nand U10425 (N_10425,N_10320,N_10297);
nand U10426 (N_10426,N_10282,N_10167);
xnor U10427 (N_10427,N_10146,N_10206);
and U10428 (N_10428,N_10224,N_10011);
xnor U10429 (N_10429,N_10032,N_10351);
nand U10430 (N_10430,N_10072,N_10382);
and U10431 (N_10431,N_10391,N_10363);
or U10432 (N_10432,N_10357,N_10083);
and U10433 (N_10433,N_10055,N_10399);
and U10434 (N_10434,N_10003,N_10081);
xor U10435 (N_10435,N_10315,N_10211);
xor U10436 (N_10436,N_10087,N_10029);
and U10437 (N_10437,N_10392,N_10018);
nor U10438 (N_10438,N_10037,N_10022);
nor U10439 (N_10439,N_10256,N_10001);
or U10440 (N_10440,N_10380,N_10213);
nand U10441 (N_10441,N_10306,N_10243);
xor U10442 (N_10442,N_10343,N_10075);
xor U10443 (N_10443,N_10186,N_10200);
nor U10444 (N_10444,N_10109,N_10150);
or U10445 (N_10445,N_10317,N_10258);
or U10446 (N_10446,N_10038,N_10017);
or U10447 (N_10447,N_10097,N_10285);
and U10448 (N_10448,N_10288,N_10198);
nand U10449 (N_10449,N_10326,N_10118);
or U10450 (N_10450,N_10267,N_10063);
nand U10451 (N_10451,N_10085,N_10093);
xor U10452 (N_10452,N_10130,N_10332);
xor U10453 (N_10453,N_10221,N_10368);
or U10454 (N_10454,N_10264,N_10176);
or U10455 (N_10455,N_10028,N_10084);
xnor U10456 (N_10456,N_10385,N_10323);
xnor U10457 (N_10457,N_10195,N_10134);
and U10458 (N_10458,N_10123,N_10179);
or U10459 (N_10459,N_10305,N_10074);
or U10460 (N_10460,N_10145,N_10260);
and U10461 (N_10461,N_10161,N_10394);
nor U10462 (N_10462,N_10045,N_10076);
nand U10463 (N_10463,N_10117,N_10240);
and U10464 (N_10464,N_10080,N_10249);
nand U10465 (N_10465,N_10027,N_10133);
xor U10466 (N_10466,N_10311,N_10155);
and U10467 (N_10467,N_10148,N_10149);
xor U10468 (N_10468,N_10387,N_10041);
and U10469 (N_10469,N_10180,N_10077);
and U10470 (N_10470,N_10222,N_10284);
and U10471 (N_10471,N_10371,N_10271);
and U10472 (N_10472,N_10291,N_10318);
nor U10473 (N_10473,N_10341,N_10102);
xnor U10474 (N_10474,N_10021,N_10319);
and U10475 (N_10475,N_10216,N_10300);
xnor U10476 (N_10476,N_10364,N_10152);
xnor U10477 (N_10477,N_10207,N_10372);
nor U10478 (N_10478,N_10230,N_10227);
xnor U10479 (N_10479,N_10287,N_10314);
nand U10480 (N_10480,N_10136,N_10068);
nor U10481 (N_10481,N_10330,N_10203);
and U10482 (N_10482,N_10000,N_10333);
and U10483 (N_10483,N_10389,N_10054);
xor U10484 (N_10484,N_10094,N_10131);
nand U10485 (N_10485,N_10255,N_10307);
nor U10486 (N_10486,N_10231,N_10008);
xnor U10487 (N_10487,N_10238,N_10367);
nand U10488 (N_10488,N_10159,N_10060);
nor U10489 (N_10489,N_10254,N_10349);
nand U10490 (N_10490,N_10012,N_10292);
and U10491 (N_10491,N_10336,N_10090);
or U10492 (N_10492,N_10245,N_10234);
or U10493 (N_10493,N_10144,N_10089);
nand U10494 (N_10494,N_10239,N_10331);
nor U10495 (N_10495,N_10009,N_10036);
or U10496 (N_10496,N_10047,N_10277);
or U10497 (N_10497,N_10162,N_10274);
nor U10498 (N_10498,N_10327,N_10177);
xnor U10499 (N_10499,N_10252,N_10158);
or U10500 (N_10500,N_10040,N_10112);
or U10501 (N_10501,N_10024,N_10023);
or U10502 (N_10502,N_10396,N_10393);
nor U10503 (N_10503,N_10064,N_10185);
or U10504 (N_10504,N_10381,N_10166);
xnor U10505 (N_10505,N_10376,N_10272);
or U10506 (N_10506,N_10053,N_10191);
nand U10507 (N_10507,N_10046,N_10283);
or U10508 (N_10508,N_10328,N_10105);
xnor U10509 (N_10509,N_10044,N_10066);
nor U10510 (N_10510,N_10168,N_10226);
nor U10511 (N_10511,N_10106,N_10169);
and U10512 (N_10512,N_10345,N_10270);
or U10513 (N_10513,N_10138,N_10236);
and U10514 (N_10514,N_10062,N_10369);
xnor U10515 (N_10515,N_10142,N_10209);
xnor U10516 (N_10516,N_10360,N_10344);
and U10517 (N_10517,N_10199,N_10005);
xor U10518 (N_10518,N_10163,N_10214);
or U10519 (N_10519,N_10154,N_10104);
nor U10520 (N_10520,N_10181,N_10135);
xnor U10521 (N_10521,N_10020,N_10127);
or U10522 (N_10522,N_10338,N_10065);
and U10523 (N_10523,N_10164,N_10061);
or U10524 (N_10524,N_10119,N_10335);
and U10525 (N_10525,N_10110,N_10212);
and U10526 (N_10526,N_10051,N_10099);
or U10527 (N_10527,N_10049,N_10321);
xor U10528 (N_10528,N_10220,N_10189);
nor U10529 (N_10529,N_10361,N_10174);
or U10530 (N_10530,N_10034,N_10359);
xnor U10531 (N_10531,N_10019,N_10375);
and U10532 (N_10532,N_10016,N_10069);
nor U10533 (N_10533,N_10275,N_10108);
or U10534 (N_10534,N_10141,N_10139);
xnor U10535 (N_10535,N_10241,N_10281);
xor U10536 (N_10536,N_10303,N_10201);
xnor U10537 (N_10537,N_10096,N_10346);
and U10538 (N_10538,N_10101,N_10050);
or U10539 (N_10539,N_10298,N_10013);
nor U10540 (N_10540,N_10313,N_10056);
or U10541 (N_10541,N_10325,N_10073);
or U10542 (N_10542,N_10153,N_10223);
and U10543 (N_10543,N_10033,N_10070);
nand U10544 (N_10544,N_10035,N_10157);
nand U10545 (N_10545,N_10312,N_10276);
or U10546 (N_10546,N_10175,N_10293);
or U10547 (N_10547,N_10286,N_10095);
or U10548 (N_10548,N_10347,N_10004);
or U10549 (N_10549,N_10002,N_10092);
or U10550 (N_10550,N_10352,N_10122);
nor U10551 (N_10551,N_10082,N_10111);
nand U10552 (N_10552,N_10010,N_10182);
nand U10553 (N_10553,N_10244,N_10114);
and U10554 (N_10554,N_10237,N_10366);
xnor U10555 (N_10555,N_10355,N_10246);
and U10556 (N_10556,N_10132,N_10308);
or U10557 (N_10557,N_10302,N_10337);
and U10558 (N_10558,N_10261,N_10262);
or U10559 (N_10559,N_10257,N_10120);
and U10560 (N_10560,N_10365,N_10232);
nor U10561 (N_10561,N_10370,N_10358);
nand U10562 (N_10562,N_10078,N_10348);
and U10563 (N_10563,N_10280,N_10116);
or U10564 (N_10564,N_10113,N_10386);
xnor U10565 (N_10565,N_10235,N_10250);
nor U10566 (N_10566,N_10140,N_10310);
or U10567 (N_10567,N_10210,N_10248);
or U10568 (N_10568,N_10128,N_10217);
and U10569 (N_10569,N_10205,N_10173);
or U10570 (N_10570,N_10014,N_10296);
nor U10571 (N_10571,N_10279,N_10294);
nand U10572 (N_10572,N_10395,N_10342);
nor U10573 (N_10573,N_10015,N_10197);
nand U10574 (N_10574,N_10125,N_10121);
or U10575 (N_10575,N_10263,N_10194);
and U10576 (N_10576,N_10259,N_10170);
nor U10577 (N_10577,N_10304,N_10299);
or U10578 (N_10578,N_10329,N_10301);
nand U10579 (N_10579,N_10039,N_10384);
xnor U10580 (N_10580,N_10273,N_10187);
nand U10581 (N_10581,N_10390,N_10048);
or U10582 (N_10582,N_10233,N_10151);
and U10583 (N_10583,N_10353,N_10397);
xnor U10584 (N_10584,N_10143,N_10204);
or U10585 (N_10585,N_10225,N_10215);
nand U10586 (N_10586,N_10098,N_10218);
nand U10587 (N_10587,N_10192,N_10184);
or U10588 (N_10588,N_10378,N_10043);
nand U10589 (N_10589,N_10086,N_10103);
xnor U10590 (N_10590,N_10377,N_10057);
or U10591 (N_10591,N_10350,N_10251);
nor U10592 (N_10592,N_10059,N_10322);
or U10593 (N_10593,N_10356,N_10156);
or U10594 (N_10594,N_10253,N_10383);
or U10595 (N_10595,N_10115,N_10339);
or U10596 (N_10596,N_10100,N_10219);
or U10597 (N_10597,N_10058,N_10091);
and U10598 (N_10598,N_10374,N_10202);
xor U10599 (N_10599,N_10379,N_10295);
xor U10600 (N_10600,N_10205,N_10317);
nand U10601 (N_10601,N_10070,N_10047);
nor U10602 (N_10602,N_10162,N_10130);
nand U10603 (N_10603,N_10257,N_10358);
or U10604 (N_10604,N_10339,N_10196);
nor U10605 (N_10605,N_10358,N_10380);
or U10606 (N_10606,N_10093,N_10168);
nand U10607 (N_10607,N_10014,N_10390);
nor U10608 (N_10608,N_10088,N_10060);
nor U10609 (N_10609,N_10109,N_10286);
nor U10610 (N_10610,N_10184,N_10275);
or U10611 (N_10611,N_10063,N_10105);
and U10612 (N_10612,N_10304,N_10290);
xor U10613 (N_10613,N_10135,N_10131);
nand U10614 (N_10614,N_10318,N_10239);
nand U10615 (N_10615,N_10240,N_10088);
nor U10616 (N_10616,N_10173,N_10371);
nor U10617 (N_10617,N_10184,N_10341);
nor U10618 (N_10618,N_10349,N_10221);
nor U10619 (N_10619,N_10104,N_10040);
nor U10620 (N_10620,N_10166,N_10109);
nor U10621 (N_10621,N_10011,N_10228);
or U10622 (N_10622,N_10152,N_10391);
or U10623 (N_10623,N_10130,N_10206);
and U10624 (N_10624,N_10358,N_10308);
and U10625 (N_10625,N_10092,N_10107);
nand U10626 (N_10626,N_10013,N_10072);
or U10627 (N_10627,N_10179,N_10054);
or U10628 (N_10628,N_10325,N_10312);
nand U10629 (N_10629,N_10358,N_10249);
and U10630 (N_10630,N_10013,N_10073);
nand U10631 (N_10631,N_10065,N_10120);
xnor U10632 (N_10632,N_10357,N_10071);
nor U10633 (N_10633,N_10239,N_10035);
and U10634 (N_10634,N_10214,N_10084);
nor U10635 (N_10635,N_10263,N_10163);
xnor U10636 (N_10636,N_10270,N_10039);
or U10637 (N_10637,N_10257,N_10341);
and U10638 (N_10638,N_10193,N_10397);
or U10639 (N_10639,N_10201,N_10322);
xor U10640 (N_10640,N_10281,N_10032);
nand U10641 (N_10641,N_10211,N_10309);
and U10642 (N_10642,N_10344,N_10012);
xnor U10643 (N_10643,N_10003,N_10138);
nor U10644 (N_10644,N_10192,N_10028);
nand U10645 (N_10645,N_10312,N_10141);
and U10646 (N_10646,N_10267,N_10385);
xor U10647 (N_10647,N_10036,N_10269);
nand U10648 (N_10648,N_10137,N_10017);
nor U10649 (N_10649,N_10021,N_10167);
and U10650 (N_10650,N_10272,N_10110);
nand U10651 (N_10651,N_10159,N_10351);
and U10652 (N_10652,N_10306,N_10298);
and U10653 (N_10653,N_10373,N_10292);
or U10654 (N_10654,N_10140,N_10315);
nand U10655 (N_10655,N_10131,N_10041);
nor U10656 (N_10656,N_10182,N_10104);
nor U10657 (N_10657,N_10149,N_10282);
or U10658 (N_10658,N_10388,N_10263);
nor U10659 (N_10659,N_10056,N_10334);
and U10660 (N_10660,N_10181,N_10093);
or U10661 (N_10661,N_10279,N_10397);
nor U10662 (N_10662,N_10312,N_10306);
or U10663 (N_10663,N_10094,N_10354);
and U10664 (N_10664,N_10331,N_10186);
nor U10665 (N_10665,N_10142,N_10057);
nand U10666 (N_10666,N_10107,N_10265);
nor U10667 (N_10667,N_10278,N_10075);
nand U10668 (N_10668,N_10044,N_10071);
nor U10669 (N_10669,N_10274,N_10127);
and U10670 (N_10670,N_10397,N_10201);
xnor U10671 (N_10671,N_10154,N_10241);
nand U10672 (N_10672,N_10274,N_10387);
nand U10673 (N_10673,N_10227,N_10098);
and U10674 (N_10674,N_10344,N_10396);
and U10675 (N_10675,N_10385,N_10032);
or U10676 (N_10676,N_10212,N_10101);
nand U10677 (N_10677,N_10008,N_10016);
xnor U10678 (N_10678,N_10310,N_10378);
xor U10679 (N_10679,N_10305,N_10059);
and U10680 (N_10680,N_10000,N_10200);
and U10681 (N_10681,N_10124,N_10165);
xor U10682 (N_10682,N_10317,N_10168);
or U10683 (N_10683,N_10392,N_10106);
nor U10684 (N_10684,N_10122,N_10237);
or U10685 (N_10685,N_10027,N_10287);
xnor U10686 (N_10686,N_10156,N_10255);
nand U10687 (N_10687,N_10137,N_10258);
nand U10688 (N_10688,N_10317,N_10004);
nor U10689 (N_10689,N_10273,N_10328);
nor U10690 (N_10690,N_10140,N_10216);
or U10691 (N_10691,N_10379,N_10307);
or U10692 (N_10692,N_10130,N_10132);
nor U10693 (N_10693,N_10099,N_10004);
or U10694 (N_10694,N_10127,N_10015);
nand U10695 (N_10695,N_10245,N_10257);
nand U10696 (N_10696,N_10143,N_10096);
or U10697 (N_10697,N_10218,N_10173);
xor U10698 (N_10698,N_10277,N_10343);
xor U10699 (N_10699,N_10023,N_10259);
nor U10700 (N_10700,N_10286,N_10101);
xnor U10701 (N_10701,N_10086,N_10005);
and U10702 (N_10702,N_10030,N_10214);
nor U10703 (N_10703,N_10191,N_10311);
nand U10704 (N_10704,N_10220,N_10149);
and U10705 (N_10705,N_10234,N_10089);
and U10706 (N_10706,N_10268,N_10298);
or U10707 (N_10707,N_10223,N_10116);
xnor U10708 (N_10708,N_10179,N_10194);
or U10709 (N_10709,N_10389,N_10218);
nor U10710 (N_10710,N_10068,N_10336);
or U10711 (N_10711,N_10293,N_10150);
nor U10712 (N_10712,N_10074,N_10388);
and U10713 (N_10713,N_10350,N_10143);
and U10714 (N_10714,N_10161,N_10040);
nand U10715 (N_10715,N_10380,N_10117);
nor U10716 (N_10716,N_10313,N_10074);
xor U10717 (N_10717,N_10255,N_10275);
or U10718 (N_10718,N_10347,N_10330);
nor U10719 (N_10719,N_10167,N_10364);
or U10720 (N_10720,N_10201,N_10000);
xor U10721 (N_10721,N_10052,N_10392);
xnor U10722 (N_10722,N_10194,N_10380);
and U10723 (N_10723,N_10296,N_10114);
xor U10724 (N_10724,N_10318,N_10171);
nand U10725 (N_10725,N_10238,N_10172);
nand U10726 (N_10726,N_10282,N_10250);
and U10727 (N_10727,N_10186,N_10346);
nor U10728 (N_10728,N_10018,N_10124);
nand U10729 (N_10729,N_10374,N_10035);
xor U10730 (N_10730,N_10291,N_10287);
nand U10731 (N_10731,N_10179,N_10047);
nor U10732 (N_10732,N_10313,N_10305);
xnor U10733 (N_10733,N_10114,N_10207);
xor U10734 (N_10734,N_10044,N_10383);
nor U10735 (N_10735,N_10084,N_10282);
nor U10736 (N_10736,N_10213,N_10258);
nand U10737 (N_10737,N_10259,N_10374);
and U10738 (N_10738,N_10241,N_10349);
nor U10739 (N_10739,N_10127,N_10146);
nand U10740 (N_10740,N_10032,N_10301);
xnor U10741 (N_10741,N_10279,N_10011);
or U10742 (N_10742,N_10128,N_10312);
xor U10743 (N_10743,N_10297,N_10048);
xor U10744 (N_10744,N_10166,N_10163);
xnor U10745 (N_10745,N_10033,N_10085);
nand U10746 (N_10746,N_10144,N_10272);
xor U10747 (N_10747,N_10379,N_10029);
nor U10748 (N_10748,N_10332,N_10170);
xnor U10749 (N_10749,N_10102,N_10075);
or U10750 (N_10750,N_10354,N_10093);
xnor U10751 (N_10751,N_10263,N_10032);
nand U10752 (N_10752,N_10190,N_10398);
and U10753 (N_10753,N_10322,N_10158);
or U10754 (N_10754,N_10279,N_10200);
nor U10755 (N_10755,N_10169,N_10133);
or U10756 (N_10756,N_10280,N_10297);
or U10757 (N_10757,N_10161,N_10299);
or U10758 (N_10758,N_10092,N_10064);
nor U10759 (N_10759,N_10334,N_10292);
nand U10760 (N_10760,N_10171,N_10136);
and U10761 (N_10761,N_10258,N_10395);
xnor U10762 (N_10762,N_10072,N_10380);
or U10763 (N_10763,N_10374,N_10350);
and U10764 (N_10764,N_10019,N_10009);
xnor U10765 (N_10765,N_10312,N_10247);
xnor U10766 (N_10766,N_10081,N_10158);
nand U10767 (N_10767,N_10327,N_10235);
nand U10768 (N_10768,N_10271,N_10079);
or U10769 (N_10769,N_10171,N_10150);
nand U10770 (N_10770,N_10211,N_10286);
xnor U10771 (N_10771,N_10077,N_10041);
and U10772 (N_10772,N_10039,N_10037);
or U10773 (N_10773,N_10212,N_10045);
nor U10774 (N_10774,N_10056,N_10225);
nand U10775 (N_10775,N_10372,N_10310);
nor U10776 (N_10776,N_10384,N_10087);
or U10777 (N_10777,N_10003,N_10274);
and U10778 (N_10778,N_10019,N_10070);
and U10779 (N_10779,N_10236,N_10263);
or U10780 (N_10780,N_10215,N_10030);
and U10781 (N_10781,N_10350,N_10214);
xor U10782 (N_10782,N_10015,N_10397);
nand U10783 (N_10783,N_10275,N_10344);
or U10784 (N_10784,N_10225,N_10219);
or U10785 (N_10785,N_10038,N_10397);
or U10786 (N_10786,N_10244,N_10387);
and U10787 (N_10787,N_10170,N_10230);
xor U10788 (N_10788,N_10304,N_10062);
and U10789 (N_10789,N_10340,N_10184);
and U10790 (N_10790,N_10391,N_10359);
or U10791 (N_10791,N_10284,N_10016);
xor U10792 (N_10792,N_10378,N_10261);
and U10793 (N_10793,N_10133,N_10200);
or U10794 (N_10794,N_10394,N_10307);
and U10795 (N_10795,N_10010,N_10153);
or U10796 (N_10796,N_10115,N_10219);
nor U10797 (N_10797,N_10176,N_10116);
xnor U10798 (N_10798,N_10115,N_10369);
xor U10799 (N_10799,N_10026,N_10140);
or U10800 (N_10800,N_10427,N_10784);
and U10801 (N_10801,N_10408,N_10471);
or U10802 (N_10802,N_10596,N_10787);
xor U10803 (N_10803,N_10790,N_10468);
or U10804 (N_10804,N_10490,N_10704);
nor U10805 (N_10805,N_10527,N_10572);
xor U10806 (N_10806,N_10440,N_10683);
or U10807 (N_10807,N_10518,N_10606);
xor U10808 (N_10808,N_10785,N_10480);
nor U10809 (N_10809,N_10594,N_10525);
or U10810 (N_10810,N_10515,N_10595);
nand U10811 (N_10811,N_10493,N_10432);
xnor U10812 (N_10812,N_10728,N_10653);
xnor U10813 (N_10813,N_10589,N_10489);
nor U10814 (N_10814,N_10508,N_10580);
xnor U10815 (N_10815,N_10757,N_10668);
nor U10816 (N_10816,N_10454,N_10610);
xnor U10817 (N_10817,N_10530,N_10667);
and U10818 (N_10818,N_10755,N_10529);
nand U10819 (N_10819,N_10738,N_10484);
xnor U10820 (N_10820,N_10776,N_10462);
nand U10821 (N_10821,N_10429,N_10777);
nand U10822 (N_10822,N_10442,N_10403);
or U10823 (N_10823,N_10762,N_10688);
nand U10824 (N_10824,N_10485,N_10754);
or U10825 (N_10825,N_10409,N_10513);
and U10826 (N_10826,N_10670,N_10693);
nand U10827 (N_10827,N_10449,N_10591);
nor U10828 (N_10828,N_10772,N_10565);
xor U10829 (N_10829,N_10569,N_10561);
and U10830 (N_10830,N_10548,N_10708);
and U10831 (N_10831,N_10458,N_10634);
and U10832 (N_10832,N_10647,N_10654);
xor U10833 (N_10833,N_10652,N_10577);
nand U10834 (N_10834,N_10737,N_10717);
nand U10835 (N_10835,N_10522,N_10694);
xor U10836 (N_10836,N_10732,N_10643);
nand U10837 (N_10837,N_10731,N_10472);
nand U10838 (N_10838,N_10450,N_10707);
and U10839 (N_10839,N_10638,N_10656);
nand U10840 (N_10840,N_10481,N_10494);
nand U10841 (N_10841,N_10767,N_10501);
and U10842 (N_10842,N_10506,N_10430);
or U10843 (N_10843,N_10526,N_10623);
or U10844 (N_10844,N_10794,N_10628);
and U10845 (N_10845,N_10697,N_10624);
or U10846 (N_10846,N_10400,N_10478);
nor U10847 (N_10847,N_10517,N_10404);
nor U10848 (N_10848,N_10679,N_10672);
nand U10849 (N_10849,N_10751,N_10648);
or U10850 (N_10850,N_10431,N_10415);
nand U10851 (N_10851,N_10632,N_10775);
or U10852 (N_10852,N_10464,N_10540);
or U10853 (N_10853,N_10781,N_10770);
nand U10854 (N_10854,N_10631,N_10786);
xor U10855 (N_10855,N_10741,N_10406);
xnor U10856 (N_10856,N_10742,N_10684);
and U10857 (N_10857,N_10663,N_10682);
nor U10858 (N_10858,N_10542,N_10523);
xor U10859 (N_10859,N_10676,N_10660);
xnor U10860 (N_10860,N_10753,N_10495);
nand U10861 (N_10861,N_10789,N_10605);
nand U10862 (N_10862,N_10763,N_10692);
xnor U10863 (N_10863,N_10657,N_10766);
xor U10864 (N_10864,N_10761,N_10460);
nand U10865 (N_10865,N_10743,N_10444);
nor U10866 (N_10866,N_10677,N_10756);
and U10867 (N_10867,N_10499,N_10538);
xor U10868 (N_10868,N_10712,N_10710);
nor U10869 (N_10869,N_10563,N_10510);
or U10870 (N_10870,N_10455,N_10503);
nand U10871 (N_10871,N_10553,N_10488);
and U10872 (N_10872,N_10607,N_10725);
nand U10873 (N_10873,N_10604,N_10441);
and U10874 (N_10874,N_10507,N_10718);
or U10875 (N_10875,N_10570,N_10615);
xnor U10876 (N_10876,N_10598,N_10410);
xor U10877 (N_10877,N_10476,N_10750);
xor U10878 (N_10878,N_10617,N_10782);
or U10879 (N_10879,N_10696,N_10706);
or U10880 (N_10880,N_10439,N_10419);
or U10881 (N_10881,N_10659,N_10630);
xnor U10882 (N_10882,N_10524,N_10603);
or U10883 (N_10883,N_10685,N_10407);
or U10884 (N_10884,N_10665,N_10649);
or U10885 (N_10885,N_10780,N_10560);
nor U10886 (N_10886,N_10747,N_10636);
or U10887 (N_10887,N_10774,N_10477);
nor U10888 (N_10888,N_10593,N_10740);
and U10889 (N_10889,N_10552,N_10555);
nand U10890 (N_10890,N_10711,N_10509);
nand U10891 (N_10891,N_10746,N_10673);
and U10892 (N_10892,N_10662,N_10461);
nand U10893 (N_10893,N_10719,N_10641);
and U10894 (N_10894,N_10412,N_10434);
nand U10895 (N_10895,N_10633,N_10744);
nor U10896 (N_10896,N_10535,N_10562);
or U10897 (N_10897,N_10613,N_10547);
xnor U10898 (N_10898,N_10414,N_10544);
and U10899 (N_10899,N_10532,N_10765);
or U10900 (N_10900,N_10578,N_10716);
and U10901 (N_10901,N_10534,N_10674);
and U10902 (N_10902,N_10799,N_10724);
xnor U10903 (N_10903,N_10511,N_10666);
nor U10904 (N_10904,N_10625,N_10498);
and U10905 (N_10905,N_10585,N_10793);
xor U10906 (N_10906,N_10729,N_10671);
nor U10907 (N_10907,N_10639,N_10587);
and U10908 (N_10908,N_10614,N_10635);
or U10909 (N_10909,N_10686,N_10436);
nor U10910 (N_10910,N_10459,N_10646);
or U10911 (N_10911,N_10637,N_10655);
xor U10912 (N_10912,N_10416,N_10512);
nand U10913 (N_10913,N_10690,N_10629);
or U10914 (N_10914,N_10497,N_10689);
or U10915 (N_10915,N_10764,N_10470);
or U10916 (N_10916,N_10675,N_10422);
xor U10917 (N_10917,N_10418,N_10733);
and U10918 (N_10918,N_10514,N_10680);
and U10919 (N_10919,N_10760,N_10622);
and U10920 (N_10920,N_10531,N_10723);
and U10921 (N_10921,N_10445,N_10730);
or U10922 (N_10922,N_10557,N_10588);
nand U10923 (N_10923,N_10448,N_10769);
nand U10924 (N_10924,N_10504,N_10681);
xor U10925 (N_10925,N_10752,N_10661);
xor U10926 (N_10926,N_10626,N_10465);
and U10927 (N_10927,N_10796,N_10437);
or U10928 (N_10928,N_10541,N_10564);
and U10929 (N_10929,N_10792,N_10620);
nand U10930 (N_10930,N_10483,N_10411);
and U10931 (N_10931,N_10745,N_10543);
or U10932 (N_10932,N_10658,N_10650);
nand U10933 (N_10933,N_10469,N_10550);
and U10934 (N_10934,N_10502,N_10642);
and U10935 (N_10935,N_10433,N_10519);
nor U10936 (N_10936,N_10616,N_10714);
or U10937 (N_10937,N_10748,N_10474);
xor U10938 (N_10938,N_10691,N_10584);
nand U10939 (N_10939,N_10453,N_10749);
and U10940 (N_10940,N_10703,N_10521);
and U10941 (N_10941,N_10758,N_10567);
nor U10942 (N_10942,N_10566,N_10621);
nor U10943 (N_10943,N_10558,N_10425);
nand U10944 (N_10944,N_10579,N_10401);
nor U10945 (N_10945,N_10701,N_10699);
nand U10946 (N_10946,N_10664,N_10612);
nor U10947 (N_10947,N_10486,N_10492);
xnor U10948 (N_10948,N_10651,N_10582);
nor U10949 (N_10949,N_10500,N_10736);
nor U10950 (N_10950,N_10735,N_10573);
and U10951 (N_10951,N_10487,N_10576);
and U10952 (N_10952,N_10788,N_10734);
nor U10953 (N_10953,N_10669,N_10739);
or U10954 (N_10954,N_10537,N_10452);
or U10955 (N_10955,N_10601,N_10705);
nand U10956 (N_10956,N_10554,N_10586);
xnor U10957 (N_10957,N_10597,N_10581);
nor U10958 (N_10958,N_10640,N_10491);
nor U10959 (N_10959,N_10721,N_10421);
or U10960 (N_10960,N_10443,N_10539);
nor U10961 (N_10961,N_10602,N_10795);
and U10962 (N_10962,N_10618,N_10768);
or U10963 (N_10963,N_10520,N_10644);
xnor U10964 (N_10964,N_10516,N_10466);
nand U10965 (N_10965,N_10559,N_10713);
or U10966 (N_10966,N_10759,N_10420);
nand U10967 (N_10967,N_10773,N_10467);
nand U10968 (N_10968,N_10592,N_10797);
and U10969 (N_10969,N_10702,N_10791);
or U10970 (N_10970,N_10426,N_10505);
or U10971 (N_10971,N_10798,N_10709);
nor U10972 (N_10972,N_10473,N_10778);
and U10973 (N_10973,N_10402,N_10599);
nor U10974 (N_10974,N_10727,N_10536);
and U10975 (N_10975,N_10771,N_10549);
nand U10976 (N_10976,N_10456,N_10545);
and U10977 (N_10977,N_10457,N_10575);
nor U10978 (N_10978,N_10463,N_10571);
nor U10979 (N_10979,N_10413,N_10574);
xnor U10980 (N_10980,N_10678,N_10627);
and U10981 (N_10981,N_10475,N_10551);
nand U10982 (N_10982,N_10423,N_10428);
nand U10983 (N_10983,N_10583,N_10687);
xnor U10984 (N_10984,N_10528,N_10611);
nand U10985 (N_10985,N_10568,N_10700);
nand U10986 (N_10986,N_10479,N_10783);
and U10987 (N_10987,N_10590,N_10405);
nand U10988 (N_10988,N_10619,N_10609);
and U10989 (N_10989,N_10726,N_10556);
xor U10990 (N_10990,N_10424,N_10438);
nor U10991 (N_10991,N_10533,N_10645);
nor U10992 (N_10992,N_10720,N_10600);
or U10993 (N_10993,N_10608,N_10779);
or U10994 (N_10994,N_10435,N_10451);
nor U10995 (N_10995,N_10446,N_10695);
and U10996 (N_10996,N_10417,N_10698);
nand U10997 (N_10997,N_10447,N_10482);
or U10998 (N_10998,N_10722,N_10715);
nand U10999 (N_10999,N_10546,N_10496);
nor U11000 (N_11000,N_10673,N_10446);
nand U11001 (N_11001,N_10706,N_10766);
and U11002 (N_11002,N_10403,N_10779);
nand U11003 (N_11003,N_10686,N_10596);
nor U11004 (N_11004,N_10459,N_10415);
or U11005 (N_11005,N_10735,N_10737);
nand U11006 (N_11006,N_10677,N_10636);
nor U11007 (N_11007,N_10780,N_10655);
and U11008 (N_11008,N_10774,N_10579);
xor U11009 (N_11009,N_10548,N_10704);
and U11010 (N_11010,N_10584,N_10629);
xor U11011 (N_11011,N_10725,N_10528);
and U11012 (N_11012,N_10712,N_10675);
nor U11013 (N_11013,N_10798,N_10460);
and U11014 (N_11014,N_10431,N_10653);
xor U11015 (N_11015,N_10617,N_10522);
or U11016 (N_11016,N_10786,N_10415);
nand U11017 (N_11017,N_10471,N_10747);
and U11018 (N_11018,N_10528,N_10762);
and U11019 (N_11019,N_10506,N_10461);
xor U11020 (N_11020,N_10433,N_10496);
xor U11021 (N_11021,N_10689,N_10411);
xnor U11022 (N_11022,N_10617,N_10703);
nor U11023 (N_11023,N_10536,N_10716);
nor U11024 (N_11024,N_10475,N_10784);
xnor U11025 (N_11025,N_10685,N_10413);
or U11026 (N_11026,N_10696,N_10713);
or U11027 (N_11027,N_10611,N_10525);
nor U11028 (N_11028,N_10697,N_10526);
and U11029 (N_11029,N_10568,N_10446);
nand U11030 (N_11030,N_10505,N_10580);
xor U11031 (N_11031,N_10406,N_10712);
nand U11032 (N_11032,N_10752,N_10479);
nand U11033 (N_11033,N_10561,N_10677);
nor U11034 (N_11034,N_10643,N_10532);
and U11035 (N_11035,N_10503,N_10714);
nand U11036 (N_11036,N_10781,N_10798);
nand U11037 (N_11037,N_10526,N_10768);
nand U11038 (N_11038,N_10570,N_10418);
nand U11039 (N_11039,N_10403,N_10714);
nand U11040 (N_11040,N_10491,N_10753);
nand U11041 (N_11041,N_10783,N_10527);
and U11042 (N_11042,N_10770,N_10528);
xor U11043 (N_11043,N_10658,N_10782);
xnor U11044 (N_11044,N_10412,N_10658);
xor U11045 (N_11045,N_10770,N_10718);
nand U11046 (N_11046,N_10727,N_10773);
or U11047 (N_11047,N_10534,N_10732);
and U11048 (N_11048,N_10790,N_10729);
nand U11049 (N_11049,N_10611,N_10589);
and U11050 (N_11050,N_10664,N_10509);
nand U11051 (N_11051,N_10724,N_10621);
nor U11052 (N_11052,N_10538,N_10480);
and U11053 (N_11053,N_10520,N_10681);
xnor U11054 (N_11054,N_10793,N_10569);
or U11055 (N_11055,N_10490,N_10614);
nand U11056 (N_11056,N_10631,N_10659);
and U11057 (N_11057,N_10767,N_10762);
nand U11058 (N_11058,N_10661,N_10623);
nor U11059 (N_11059,N_10548,N_10792);
nor U11060 (N_11060,N_10725,N_10774);
and U11061 (N_11061,N_10522,N_10533);
nand U11062 (N_11062,N_10400,N_10730);
nand U11063 (N_11063,N_10722,N_10436);
xnor U11064 (N_11064,N_10660,N_10536);
and U11065 (N_11065,N_10785,N_10408);
nand U11066 (N_11066,N_10499,N_10439);
and U11067 (N_11067,N_10412,N_10461);
and U11068 (N_11068,N_10463,N_10498);
nor U11069 (N_11069,N_10743,N_10768);
nor U11070 (N_11070,N_10712,N_10481);
and U11071 (N_11071,N_10444,N_10470);
or U11072 (N_11072,N_10473,N_10693);
nor U11073 (N_11073,N_10738,N_10590);
or U11074 (N_11074,N_10518,N_10623);
nand U11075 (N_11075,N_10751,N_10776);
and U11076 (N_11076,N_10478,N_10619);
and U11077 (N_11077,N_10687,N_10611);
nor U11078 (N_11078,N_10675,N_10444);
nand U11079 (N_11079,N_10495,N_10480);
or U11080 (N_11080,N_10591,N_10516);
nor U11081 (N_11081,N_10799,N_10699);
xor U11082 (N_11082,N_10543,N_10497);
nand U11083 (N_11083,N_10560,N_10683);
nand U11084 (N_11084,N_10569,N_10679);
or U11085 (N_11085,N_10487,N_10569);
nand U11086 (N_11086,N_10503,N_10651);
nand U11087 (N_11087,N_10539,N_10783);
or U11088 (N_11088,N_10761,N_10471);
or U11089 (N_11089,N_10607,N_10708);
nand U11090 (N_11090,N_10514,N_10679);
nor U11091 (N_11091,N_10673,N_10783);
and U11092 (N_11092,N_10488,N_10400);
nand U11093 (N_11093,N_10416,N_10568);
nor U11094 (N_11094,N_10599,N_10659);
nor U11095 (N_11095,N_10588,N_10764);
xnor U11096 (N_11096,N_10462,N_10777);
nand U11097 (N_11097,N_10474,N_10583);
xor U11098 (N_11098,N_10622,N_10677);
or U11099 (N_11099,N_10706,N_10774);
and U11100 (N_11100,N_10592,N_10736);
nand U11101 (N_11101,N_10592,N_10764);
xnor U11102 (N_11102,N_10558,N_10521);
nor U11103 (N_11103,N_10692,N_10762);
xor U11104 (N_11104,N_10590,N_10556);
xor U11105 (N_11105,N_10549,N_10737);
xnor U11106 (N_11106,N_10754,N_10467);
and U11107 (N_11107,N_10484,N_10565);
nor U11108 (N_11108,N_10486,N_10671);
or U11109 (N_11109,N_10699,N_10553);
nor U11110 (N_11110,N_10493,N_10655);
nor U11111 (N_11111,N_10552,N_10425);
nand U11112 (N_11112,N_10488,N_10570);
and U11113 (N_11113,N_10668,N_10678);
xor U11114 (N_11114,N_10742,N_10620);
nor U11115 (N_11115,N_10431,N_10596);
and U11116 (N_11116,N_10566,N_10742);
and U11117 (N_11117,N_10597,N_10546);
nand U11118 (N_11118,N_10494,N_10515);
or U11119 (N_11119,N_10741,N_10748);
or U11120 (N_11120,N_10554,N_10762);
xor U11121 (N_11121,N_10781,N_10753);
nand U11122 (N_11122,N_10776,N_10452);
xor U11123 (N_11123,N_10503,N_10751);
nor U11124 (N_11124,N_10522,N_10663);
nor U11125 (N_11125,N_10581,N_10424);
or U11126 (N_11126,N_10459,N_10542);
and U11127 (N_11127,N_10414,N_10595);
xnor U11128 (N_11128,N_10578,N_10584);
xnor U11129 (N_11129,N_10420,N_10751);
xnor U11130 (N_11130,N_10517,N_10523);
nand U11131 (N_11131,N_10649,N_10621);
xor U11132 (N_11132,N_10592,N_10645);
or U11133 (N_11133,N_10616,N_10490);
or U11134 (N_11134,N_10520,N_10676);
or U11135 (N_11135,N_10652,N_10616);
xnor U11136 (N_11136,N_10791,N_10515);
and U11137 (N_11137,N_10576,N_10758);
nor U11138 (N_11138,N_10606,N_10756);
or U11139 (N_11139,N_10609,N_10424);
xor U11140 (N_11140,N_10759,N_10435);
nand U11141 (N_11141,N_10727,N_10794);
nand U11142 (N_11142,N_10401,N_10723);
xnor U11143 (N_11143,N_10469,N_10548);
nor U11144 (N_11144,N_10617,N_10755);
and U11145 (N_11145,N_10578,N_10466);
and U11146 (N_11146,N_10691,N_10760);
xor U11147 (N_11147,N_10501,N_10774);
and U11148 (N_11148,N_10535,N_10557);
or U11149 (N_11149,N_10405,N_10415);
xor U11150 (N_11150,N_10423,N_10489);
xnor U11151 (N_11151,N_10676,N_10626);
or U11152 (N_11152,N_10723,N_10766);
nor U11153 (N_11153,N_10738,N_10441);
and U11154 (N_11154,N_10709,N_10506);
and U11155 (N_11155,N_10504,N_10676);
xor U11156 (N_11156,N_10473,N_10493);
or U11157 (N_11157,N_10771,N_10460);
xor U11158 (N_11158,N_10719,N_10464);
nor U11159 (N_11159,N_10725,N_10436);
xnor U11160 (N_11160,N_10785,N_10652);
nor U11161 (N_11161,N_10410,N_10573);
nand U11162 (N_11162,N_10691,N_10665);
or U11163 (N_11163,N_10542,N_10456);
nor U11164 (N_11164,N_10745,N_10765);
or U11165 (N_11165,N_10702,N_10695);
xnor U11166 (N_11166,N_10728,N_10723);
nand U11167 (N_11167,N_10637,N_10584);
or U11168 (N_11168,N_10753,N_10623);
xnor U11169 (N_11169,N_10673,N_10600);
nor U11170 (N_11170,N_10733,N_10628);
or U11171 (N_11171,N_10639,N_10684);
nor U11172 (N_11172,N_10545,N_10692);
nor U11173 (N_11173,N_10712,N_10652);
or U11174 (N_11174,N_10472,N_10651);
and U11175 (N_11175,N_10450,N_10483);
xnor U11176 (N_11176,N_10592,N_10760);
or U11177 (N_11177,N_10609,N_10671);
nor U11178 (N_11178,N_10400,N_10601);
nor U11179 (N_11179,N_10634,N_10607);
nor U11180 (N_11180,N_10556,N_10567);
nand U11181 (N_11181,N_10725,N_10427);
or U11182 (N_11182,N_10722,N_10656);
nor U11183 (N_11183,N_10518,N_10428);
nand U11184 (N_11184,N_10672,N_10473);
nand U11185 (N_11185,N_10595,N_10702);
nand U11186 (N_11186,N_10715,N_10713);
or U11187 (N_11187,N_10603,N_10749);
or U11188 (N_11188,N_10419,N_10741);
or U11189 (N_11189,N_10628,N_10683);
xnor U11190 (N_11190,N_10714,N_10567);
nor U11191 (N_11191,N_10631,N_10420);
nand U11192 (N_11192,N_10560,N_10503);
xor U11193 (N_11193,N_10755,N_10505);
xor U11194 (N_11194,N_10680,N_10428);
nand U11195 (N_11195,N_10596,N_10684);
xnor U11196 (N_11196,N_10618,N_10516);
xor U11197 (N_11197,N_10452,N_10495);
xor U11198 (N_11198,N_10604,N_10484);
and U11199 (N_11199,N_10796,N_10630);
or U11200 (N_11200,N_11053,N_10949);
and U11201 (N_11201,N_11024,N_10955);
xnor U11202 (N_11202,N_11152,N_11186);
nand U11203 (N_11203,N_11043,N_11123);
nor U11204 (N_11204,N_11182,N_11117);
or U11205 (N_11205,N_11107,N_11039);
nand U11206 (N_11206,N_10987,N_11002);
nand U11207 (N_11207,N_11108,N_11083);
and U11208 (N_11208,N_11138,N_10965);
nand U11209 (N_11209,N_10894,N_10856);
nand U11210 (N_11210,N_11170,N_11036);
and U11211 (N_11211,N_10883,N_10925);
nor U11212 (N_11212,N_10871,N_10834);
and U11213 (N_11213,N_10958,N_11047);
and U11214 (N_11214,N_10954,N_11173);
xnor U11215 (N_11215,N_10908,N_11062);
nand U11216 (N_11216,N_10988,N_11198);
or U11217 (N_11217,N_11081,N_11089);
nand U11218 (N_11218,N_10896,N_10811);
or U11219 (N_11219,N_10858,N_11038);
nor U11220 (N_11220,N_10808,N_10963);
nand U11221 (N_11221,N_10866,N_10930);
xor U11222 (N_11222,N_11011,N_11155);
and U11223 (N_11223,N_10975,N_10953);
xor U11224 (N_11224,N_10961,N_10861);
or U11225 (N_11225,N_10882,N_10997);
nand U11226 (N_11226,N_10990,N_11102);
nand U11227 (N_11227,N_11103,N_10960);
and U11228 (N_11228,N_10859,N_10815);
nand U11229 (N_11229,N_11183,N_11129);
or U11230 (N_11230,N_10819,N_11176);
and U11231 (N_11231,N_10804,N_11158);
and U11232 (N_11232,N_11013,N_10835);
and U11233 (N_11233,N_11063,N_11100);
or U11234 (N_11234,N_11082,N_11065);
xnor U11235 (N_11235,N_11190,N_11185);
nor U11236 (N_11236,N_11007,N_10853);
or U11237 (N_11237,N_11104,N_10909);
xnor U11238 (N_11238,N_10847,N_10971);
nand U11239 (N_11239,N_11092,N_11021);
nor U11240 (N_11240,N_10869,N_11044);
nor U11241 (N_11241,N_10889,N_10881);
and U11242 (N_11242,N_11090,N_10951);
nand U11243 (N_11243,N_11064,N_10974);
nor U11244 (N_11244,N_11077,N_10845);
xor U11245 (N_11245,N_10920,N_10812);
or U11246 (N_11246,N_11136,N_11048);
nor U11247 (N_11247,N_11005,N_11035);
xnor U11248 (N_11248,N_11033,N_11006);
xor U11249 (N_11249,N_10867,N_10982);
nand U11250 (N_11250,N_11160,N_11075);
and U11251 (N_11251,N_10814,N_10905);
nand U11252 (N_11252,N_10839,N_10966);
and U11253 (N_11253,N_11174,N_11093);
nor U11254 (N_11254,N_11040,N_10921);
and U11255 (N_11255,N_11150,N_11028);
xnor U11256 (N_11256,N_11025,N_10898);
and U11257 (N_11257,N_11073,N_10855);
and U11258 (N_11258,N_10843,N_10913);
xnor U11259 (N_11259,N_10902,N_11034);
nor U11260 (N_11260,N_10980,N_11042);
nor U11261 (N_11261,N_10891,N_10817);
or U11262 (N_11262,N_10849,N_11139);
xnor U11263 (N_11263,N_11131,N_10911);
nand U11264 (N_11264,N_11088,N_10984);
or U11265 (N_11265,N_11161,N_10876);
nand U11266 (N_11266,N_10977,N_11084);
and U11267 (N_11267,N_10886,N_11134);
xnor U11268 (N_11268,N_10995,N_11135);
or U11269 (N_11269,N_10936,N_10993);
xor U11270 (N_11270,N_11059,N_11116);
xnor U11271 (N_11271,N_10964,N_10848);
or U11272 (N_11272,N_11066,N_10810);
nand U11273 (N_11273,N_11001,N_11012);
nor U11274 (N_11274,N_10967,N_11106);
nor U11275 (N_11275,N_10873,N_11156);
and U11276 (N_11276,N_11056,N_10850);
and U11277 (N_11277,N_10991,N_11060);
nor U11278 (N_11278,N_11192,N_11140);
and U11279 (N_11279,N_10885,N_10901);
and U11280 (N_11280,N_10945,N_11019);
or U11281 (N_11281,N_10823,N_11175);
xor U11282 (N_11282,N_10938,N_11050);
or U11283 (N_11283,N_10892,N_11189);
xor U11284 (N_11284,N_10924,N_10926);
nor U11285 (N_11285,N_11097,N_11020);
nand U11286 (N_11286,N_10923,N_10900);
nor U11287 (N_11287,N_10922,N_11037);
nand U11288 (N_11288,N_10948,N_10985);
nor U11289 (N_11289,N_10822,N_10992);
nand U11290 (N_11290,N_11184,N_10956);
nand U11291 (N_11291,N_10880,N_11099);
xor U11292 (N_11292,N_11032,N_10842);
and U11293 (N_11293,N_10865,N_11162);
and U11294 (N_11294,N_11142,N_11143);
xnor U11295 (N_11295,N_10973,N_11127);
and U11296 (N_11296,N_11166,N_11027);
nand U11297 (N_11297,N_10820,N_11141);
nand U11298 (N_11298,N_10830,N_10903);
and U11299 (N_11299,N_11003,N_11031);
xor U11300 (N_11300,N_11008,N_10827);
nor U11301 (N_11301,N_11068,N_11159);
and U11302 (N_11302,N_10832,N_10904);
nand U11303 (N_11303,N_11074,N_10933);
xor U11304 (N_11304,N_10844,N_10872);
or U11305 (N_11305,N_10857,N_11165);
nand U11306 (N_11306,N_10888,N_11026);
nor U11307 (N_11307,N_11094,N_10816);
or U11308 (N_11308,N_10846,N_11101);
or U11309 (N_11309,N_11151,N_11157);
nand U11310 (N_11310,N_10942,N_10829);
and U11311 (N_11311,N_11055,N_11167);
and U11312 (N_11312,N_11049,N_10863);
and U11313 (N_11313,N_10878,N_10929);
nor U11314 (N_11314,N_10868,N_11057);
nor U11315 (N_11315,N_10944,N_10946);
or U11316 (N_11316,N_10813,N_11133);
xor U11317 (N_11317,N_11124,N_10996);
and U11318 (N_11318,N_11061,N_10890);
and U11319 (N_11319,N_10917,N_10838);
or U11320 (N_11320,N_11187,N_10828);
xnor U11321 (N_11321,N_11078,N_10833);
nand U11322 (N_11322,N_10862,N_11098);
nand U11323 (N_11323,N_11113,N_10916);
nand U11324 (N_11324,N_11076,N_10803);
xnor U11325 (N_11325,N_11052,N_10860);
nand U11326 (N_11326,N_10934,N_10818);
or U11327 (N_11327,N_11000,N_10807);
nand U11328 (N_11328,N_11023,N_11070);
nor U11329 (N_11329,N_10874,N_11119);
xnor U11330 (N_11330,N_11126,N_11091);
nor U11331 (N_11331,N_10805,N_10854);
nand U11332 (N_11332,N_11137,N_10981);
nor U11333 (N_11333,N_10969,N_11071);
nor U11334 (N_11334,N_10877,N_11132);
or U11335 (N_11335,N_11114,N_10895);
nor U11336 (N_11336,N_10806,N_11145);
and U11337 (N_11337,N_10935,N_10800);
nand U11338 (N_11338,N_11146,N_10802);
nor U11339 (N_11339,N_11086,N_11199);
or U11340 (N_11340,N_11120,N_11171);
or U11341 (N_11341,N_11079,N_10940);
or U11342 (N_11342,N_11188,N_11153);
nor U11343 (N_11343,N_10907,N_11111);
nand U11344 (N_11344,N_10968,N_10941);
or U11345 (N_11345,N_11030,N_10999);
or U11346 (N_11346,N_11180,N_11004);
and U11347 (N_11347,N_10851,N_11169);
nor U11348 (N_11348,N_11105,N_10994);
and U11349 (N_11349,N_10870,N_11095);
or U11350 (N_11350,N_10962,N_10947);
or U11351 (N_11351,N_10983,N_10879);
nand U11352 (N_11352,N_11022,N_10976);
nor U11353 (N_11353,N_11051,N_11096);
nor U11354 (N_11354,N_11149,N_10986);
nor U11355 (N_11355,N_10915,N_10837);
nor U11356 (N_11356,N_10840,N_11109);
xnor U11357 (N_11357,N_10998,N_11017);
and U11358 (N_11358,N_10979,N_10875);
and U11359 (N_11359,N_11115,N_11087);
nor U11360 (N_11360,N_10950,N_11058);
xor U11361 (N_11361,N_10919,N_10801);
and U11362 (N_11362,N_10836,N_10914);
xor U11363 (N_11363,N_11018,N_10937);
nor U11364 (N_11364,N_11154,N_11148);
nor U11365 (N_11365,N_10931,N_11177);
or U11366 (N_11366,N_11194,N_11195);
nor U11367 (N_11367,N_11046,N_11029);
nor U11368 (N_11368,N_10952,N_10910);
xor U11369 (N_11369,N_10864,N_11130);
nor U11370 (N_11370,N_10939,N_10978);
nor U11371 (N_11371,N_11054,N_11014);
and U11372 (N_11372,N_11069,N_10841);
or U11373 (N_11373,N_11181,N_10989);
or U11374 (N_11374,N_11122,N_11147);
nor U11375 (N_11375,N_11128,N_10821);
nand U11376 (N_11376,N_10893,N_11067);
xor U11377 (N_11377,N_11110,N_11144);
nand U11378 (N_11378,N_10970,N_10972);
or U11379 (N_11379,N_11168,N_10831);
and U11380 (N_11380,N_11197,N_10887);
nand U11381 (N_11381,N_11009,N_10959);
or U11382 (N_11382,N_11080,N_11085);
and U11383 (N_11383,N_11172,N_11121);
or U11384 (N_11384,N_10899,N_10928);
and U11385 (N_11385,N_11125,N_10932);
or U11386 (N_11386,N_11041,N_11118);
xnor U11387 (N_11387,N_10927,N_10918);
nand U11388 (N_11388,N_10943,N_10809);
nor U11389 (N_11389,N_11072,N_10884);
and U11390 (N_11390,N_11196,N_11112);
nand U11391 (N_11391,N_10824,N_10852);
nor U11392 (N_11392,N_11016,N_11179);
nor U11393 (N_11393,N_10957,N_10825);
nor U11394 (N_11394,N_11178,N_10906);
or U11395 (N_11395,N_10826,N_11193);
xor U11396 (N_11396,N_11163,N_11045);
nor U11397 (N_11397,N_11010,N_10897);
or U11398 (N_11398,N_10912,N_11015);
or U11399 (N_11399,N_11164,N_11191);
and U11400 (N_11400,N_10805,N_11006);
or U11401 (N_11401,N_11131,N_10951);
xnor U11402 (N_11402,N_10828,N_11036);
and U11403 (N_11403,N_10991,N_11102);
nand U11404 (N_11404,N_11017,N_11094);
and U11405 (N_11405,N_10867,N_10978);
xor U11406 (N_11406,N_11075,N_10995);
xnor U11407 (N_11407,N_10825,N_11142);
nor U11408 (N_11408,N_11132,N_11052);
or U11409 (N_11409,N_11186,N_10847);
or U11410 (N_11410,N_11131,N_11017);
nand U11411 (N_11411,N_11191,N_11172);
and U11412 (N_11412,N_10985,N_10865);
and U11413 (N_11413,N_10884,N_11032);
nand U11414 (N_11414,N_10840,N_10890);
nor U11415 (N_11415,N_10835,N_11142);
and U11416 (N_11416,N_10934,N_10994);
nor U11417 (N_11417,N_11123,N_10848);
or U11418 (N_11418,N_11140,N_10819);
xnor U11419 (N_11419,N_11036,N_11146);
or U11420 (N_11420,N_10893,N_10895);
nand U11421 (N_11421,N_11127,N_10970);
and U11422 (N_11422,N_10835,N_11193);
or U11423 (N_11423,N_11127,N_11038);
xor U11424 (N_11424,N_10924,N_10890);
nand U11425 (N_11425,N_10889,N_10888);
nor U11426 (N_11426,N_11138,N_10900);
or U11427 (N_11427,N_11195,N_11064);
and U11428 (N_11428,N_11197,N_11101);
xor U11429 (N_11429,N_11121,N_11100);
nand U11430 (N_11430,N_11014,N_11144);
or U11431 (N_11431,N_10833,N_10916);
or U11432 (N_11432,N_11122,N_10830);
and U11433 (N_11433,N_11127,N_10954);
nand U11434 (N_11434,N_11188,N_11103);
xor U11435 (N_11435,N_10939,N_10883);
and U11436 (N_11436,N_10914,N_11036);
nand U11437 (N_11437,N_11083,N_11146);
or U11438 (N_11438,N_11192,N_11188);
nor U11439 (N_11439,N_11020,N_11056);
nand U11440 (N_11440,N_10914,N_11199);
nor U11441 (N_11441,N_10985,N_11102);
nand U11442 (N_11442,N_10980,N_10944);
nand U11443 (N_11443,N_10861,N_11197);
xor U11444 (N_11444,N_10847,N_11093);
xor U11445 (N_11445,N_10994,N_11130);
and U11446 (N_11446,N_11114,N_10954);
nor U11447 (N_11447,N_11112,N_10926);
nand U11448 (N_11448,N_11035,N_10817);
xor U11449 (N_11449,N_10992,N_10829);
xnor U11450 (N_11450,N_10920,N_11096);
and U11451 (N_11451,N_10834,N_11163);
xnor U11452 (N_11452,N_10815,N_10902);
xor U11453 (N_11453,N_11081,N_11122);
or U11454 (N_11454,N_10999,N_11031);
and U11455 (N_11455,N_11048,N_10948);
nor U11456 (N_11456,N_11103,N_11041);
or U11457 (N_11457,N_11028,N_11091);
nor U11458 (N_11458,N_11089,N_10993);
nor U11459 (N_11459,N_10934,N_10868);
and U11460 (N_11460,N_11139,N_11015);
nor U11461 (N_11461,N_10871,N_11187);
and U11462 (N_11462,N_10826,N_11166);
or U11463 (N_11463,N_11158,N_10953);
xnor U11464 (N_11464,N_10865,N_11078);
and U11465 (N_11465,N_11054,N_11075);
nor U11466 (N_11466,N_11109,N_11049);
nor U11467 (N_11467,N_10856,N_10885);
nor U11468 (N_11468,N_10906,N_11008);
nand U11469 (N_11469,N_11083,N_10951);
or U11470 (N_11470,N_11099,N_10951);
xor U11471 (N_11471,N_10812,N_10823);
nor U11472 (N_11472,N_10998,N_10819);
nor U11473 (N_11473,N_10847,N_11169);
nor U11474 (N_11474,N_11099,N_11164);
and U11475 (N_11475,N_10840,N_11102);
nor U11476 (N_11476,N_11026,N_11004);
or U11477 (N_11477,N_11006,N_10818);
or U11478 (N_11478,N_10997,N_10934);
nand U11479 (N_11479,N_10823,N_10801);
xor U11480 (N_11480,N_11105,N_10980);
nand U11481 (N_11481,N_11045,N_11074);
xor U11482 (N_11482,N_11174,N_10870);
nand U11483 (N_11483,N_11066,N_10856);
or U11484 (N_11484,N_10919,N_11005);
nor U11485 (N_11485,N_11097,N_11122);
xor U11486 (N_11486,N_11073,N_10803);
nor U11487 (N_11487,N_10869,N_10804);
nand U11488 (N_11488,N_11194,N_10866);
nand U11489 (N_11489,N_11089,N_10821);
or U11490 (N_11490,N_11070,N_10924);
xor U11491 (N_11491,N_11000,N_11050);
or U11492 (N_11492,N_10960,N_10850);
nand U11493 (N_11493,N_10801,N_10908);
nand U11494 (N_11494,N_11141,N_10867);
xor U11495 (N_11495,N_10822,N_10859);
nor U11496 (N_11496,N_10925,N_10860);
xnor U11497 (N_11497,N_11008,N_11135);
nand U11498 (N_11498,N_11126,N_11172);
xor U11499 (N_11499,N_11168,N_11139);
or U11500 (N_11500,N_11083,N_11118);
xnor U11501 (N_11501,N_11085,N_11115);
nor U11502 (N_11502,N_11065,N_10995);
nor U11503 (N_11503,N_10835,N_11080);
xnor U11504 (N_11504,N_11169,N_10932);
and U11505 (N_11505,N_11184,N_10979);
or U11506 (N_11506,N_10857,N_10866);
nand U11507 (N_11507,N_10919,N_10882);
xnor U11508 (N_11508,N_10872,N_11195);
or U11509 (N_11509,N_10801,N_11039);
nand U11510 (N_11510,N_10879,N_11078);
and U11511 (N_11511,N_10829,N_11072);
and U11512 (N_11512,N_11023,N_11128);
or U11513 (N_11513,N_11129,N_10978);
nand U11514 (N_11514,N_10994,N_10868);
and U11515 (N_11515,N_11091,N_10832);
xor U11516 (N_11516,N_11188,N_11139);
and U11517 (N_11517,N_10919,N_11047);
xor U11518 (N_11518,N_11196,N_11043);
xor U11519 (N_11519,N_11015,N_11186);
nor U11520 (N_11520,N_11087,N_10875);
xor U11521 (N_11521,N_10866,N_11038);
nor U11522 (N_11522,N_10831,N_10985);
xor U11523 (N_11523,N_11090,N_10854);
xor U11524 (N_11524,N_10893,N_10921);
nand U11525 (N_11525,N_11066,N_11195);
nor U11526 (N_11526,N_11114,N_11188);
or U11527 (N_11527,N_10904,N_10801);
nor U11528 (N_11528,N_10897,N_11105);
or U11529 (N_11529,N_10978,N_11181);
nor U11530 (N_11530,N_11131,N_10858);
xnor U11531 (N_11531,N_11174,N_10916);
or U11532 (N_11532,N_10963,N_10989);
nor U11533 (N_11533,N_11178,N_11188);
xnor U11534 (N_11534,N_11122,N_11115);
or U11535 (N_11535,N_11048,N_11037);
xnor U11536 (N_11536,N_10863,N_10977);
nor U11537 (N_11537,N_11105,N_10850);
nor U11538 (N_11538,N_11169,N_11121);
and U11539 (N_11539,N_11136,N_10907);
xor U11540 (N_11540,N_10823,N_10817);
and U11541 (N_11541,N_11015,N_11014);
or U11542 (N_11542,N_10842,N_11064);
nor U11543 (N_11543,N_11022,N_10817);
xor U11544 (N_11544,N_11078,N_10911);
nand U11545 (N_11545,N_10944,N_11112);
xnor U11546 (N_11546,N_10844,N_10847);
xor U11547 (N_11547,N_11191,N_11045);
and U11548 (N_11548,N_11008,N_10911);
xnor U11549 (N_11549,N_11142,N_11036);
or U11550 (N_11550,N_10939,N_11178);
xor U11551 (N_11551,N_10924,N_10955);
or U11552 (N_11552,N_11106,N_11078);
xnor U11553 (N_11553,N_10973,N_11031);
nand U11554 (N_11554,N_11162,N_11066);
nor U11555 (N_11555,N_11009,N_11191);
xor U11556 (N_11556,N_10880,N_10951);
and U11557 (N_11557,N_11140,N_10876);
nor U11558 (N_11558,N_10905,N_11059);
xor U11559 (N_11559,N_11159,N_11122);
xnor U11560 (N_11560,N_11105,N_11075);
nor U11561 (N_11561,N_11182,N_11083);
or U11562 (N_11562,N_11114,N_11186);
or U11563 (N_11563,N_11049,N_11193);
and U11564 (N_11564,N_11046,N_10907);
nand U11565 (N_11565,N_10952,N_10967);
xnor U11566 (N_11566,N_11042,N_10918);
xor U11567 (N_11567,N_10815,N_11025);
or U11568 (N_11568,N_11070,N_10957);
xnor U11569 (N_11569,N_10895,N_11167);
and U11570 (N_11570,N_10815,N_10807);
xor U11571 (N_11571,N_11157,N_11083);
and U11572 (N_11572,N_10873,N_10962);
nor U11573 (N_11573,N_10982,N_10862);
nand U11574 (N_11574,N_11167,N_10871);
and U11575 (N_11575,N_11126,N_10892);
nor U11576 (N_11576,N_10893,N_10884);
nand U11577 (N_11577,N_11129,N_10922);
and U11578 (N_11578,N_10908,N_10885);
xor U11579 (N_11579,N_11141,N_11105);
nand U11580 (N_11580,N_10818,N_11016);
nand U11581 (N_11581,N_11121,N_11153);
or U11582 (N_11582,N_11163,N_11149);
and U11583 (N_11583,N_11088,N_10881);
and U11584 (N_11584,N_10993,N_11117);
nand U11585 (N_11585,N_11078,N_11162);
nand U11586 (N_11586,N_10897,N_10948);
or U11587 (N_11587,N_11112,N_11023);
and U11588 (N_11588,N_11155,N_11002);
and U11589 (N_11589,N_11138,N_11037);
nor U11590 (N_11590,N_10953,N_11085);
or U11591 (N_11591,N_10854,N_11143);
and U11592 (N_11592,N_11036,N_11045);
or U11593 (N_11593,N_11113,N_10841);
xnor U11594 (N_11594,N_10805,N_10901);
or U11595 (N_11595,N_10891,N_10934);
and U11596 (N_11596,N_11130,N_11054);
and U11597 (N_11597,N_11183,N_10899);
and U11598 (N_11598,N_11042,N_11050);
xnor U11599 (N_11599,N_10823,N_10855);
or U11600 (N_11600,N_11216,N_11315);
and U11601 (N_11601,N_11245,N_11511);
or U11602 (N_11602,N_11249,N_11594);
and U11603 (N_11603,N_11524,N_11481);
xor U11604 (N_11604,N_11548,N_11351);
and U11605 (N_11605,N_11332,N_11423);
xor U11606 (N_11606,N_11286,N_11321);
nor U11607 (N_11607,N_11488,N_11520);
nand U11608 (N_11608,N_11593,N_11257);
and U11609 (N_11609,N_11383,N_11455);
xnor U11610 (N_11610,N_11205,N_11405);
nor U11611 (N_11611,N_11562,N_11510);
nor U11612 (N_11612,N_11251,N_11290);
or U11613 (N_11613,N_11487,N_11209);
nor U11614 (N_11614,N_11428,N_11486);
or U11615 (N_11615,N_11381,N_11277);
xnor U11616 (N_11616,N_11443,N_11264);
nor U11617 (N_11617,N_11328,N_11576);
or U11618 (N_11618,N_11400,N_11538);
and U11619 (N_11619,N_11225,N_11206);
xor U11620 (N_11620,N_11402,N_11412);
nand U11621 (N_11621,N_11268,N_11541);
xnor U11622 (N_11622,N_11462,N_11410);
or U11623 (N_11623,N_11344,N_11472);
or U11624 (N_11624,N_11543,N_11378);
or U11625 (N_11625,N_11528,N_11440);
xor U11626 (N_11626,N_11363,N_11456);
xor U11627 (N_11627,N_11326,N_11222);
nand U11628 (N_11628,N_11558,N_11427);
or U11629 (N_11629,N_11388,N_11523);
nand U11630 (N_11630,N_11508,N_11208);
xor U11631 (N_11631,N_11358,N_11495);
and U11632 (N_11632,N_11275,N_11295);
or U11633 (N_11633,N_11228,N_11215);
nor U11634 (N_11634,N_11309,N_11273);
or U11635 (N_11635,N_11550,N_11557);
and U11636 (N_11636,N_11537,N_11409);
and U11637 (N_11637,N_11221,N_11573);
and U11638 (N_11638,N_11483,N_11577);
nor U11639 (N_11639,N_11255,N_11404);
and U11640 (N_11640,N_11392,N_11283);
nand U11641 (N_11641,N_11514,N_11376);
nand U11642 (N_11642,N_11564,N_11254);
or U11643 (N_11643,N_11329,N_11568);
xnor U11644 (N_11644,N_11287,N_11355);
xor U11645 (N_11645,N_11551,N_11248);
xnor U11646 (N_11646,N_11323,N_11201);
nor U11647 (N_11647,N_11203,N_11547);
xnor U11648 (N_11648,N_11438,N_11461);
nor U11649 (N_11649,N_11339,N_11253);
and U11650 (N_11650,N_11233,N_11210);
or U11651 (N_11651,N_11242,N_11469);
or U11652 (N_11652,N_11202,N_11213);
nand U11653 (N_11653,N_11407,N_11578);
xor U11654 (N_11654,N_11545,N_11308);
nand U11655 (N_11655,N_11281,N_11369);
nor U11656 (N_11656,N_11352,N_11333);
or U11657 (N_11657,N_11342,N_11529);
or U11658 (N_11658,N_11526,N_11360);
and U11659 (N_11659,N_11539,N_11503);
xnor U11660 (N_11660,N_11575,N_11552);
xnor U11661 (N_11661,N_11530,N_11554);
and U11662 (N_11662,N_11244,N_11570);
and U11663 (N_11663,N_11436,N_11294);
xor U11664 (N_11664,N_11331,N_11421);
or U11665 (N_11665,N_11289,N_11463);
or U11666 (N_11666,N_11274,N_11445);
nor U11667 (N_11667,N_11517,N_11343);
nand U11668 (N_11668,N_11297,N_11382);
nand U11669 (N_11669,N_11512,N_11347);
xnor U11670 (N_11670,N_11350,N_11411);
nand U11671 (N_11671,N_11466,N_11227);
xnor U11672 (N_11672,N_11306,N_11441);
xor U11673 (N_11673,N_11279,N_11263);
xnor U11674 (N_11674,N_11446,N_11460);
or U11675 (N_11675,N_11395,N_11403);
nand U11676 (N_11676,N_11569,N_11549);
or U11677 (N_11677,N_11498,N_11565);
xor U11678 (N_11678,N_11505,N_11373);
and U11679 (N_11679,N_11387,N_11319);
and U11680 (N_11680,N_11585,N_11223);
nand U11681 (N_11681,N_11497,N_11396);
nor U11682 (N_11682,N_11515,N_11327);
nor U11683 (N_11683,N_11596,N_11420);
or U11684 (N_11684,N_11507,N_11561);
and U11685 (N_11685,N_11540,N_11231);
nor U11686 (N_11686,N_11235,N_11482);
nor U11687 (N_11687,N_11470,N_11311);
nand U11688 (N_11688,N_11419,N_11371);
nand U11689 (N_11689,N_11285,N_11384);
nor U11690 (N_11690,N_11590,N_11491);
and U11691 (N_11691,N_11261,N_11240);
nand U11692 (N_11692,N_11340,N_11219);
nand U11693 (N_11693,N_11459,N_11348);
or U11694 (N_11694,N_11256,N_11313);
xnor U11695 (N_11695,N_11566,N_11485);
nand U11696 (N_11696,N_11424,N_11307);
nor U11697 (N_11697,N_11413,N_11303);
and U11698 (N_11698,N_11474,N_11574);
nor U11699 (N_11699,N_11418,N_11439);
and U11700 (N_11700,N_11316,N_11429);
or U11701 (N_11701,N_11494,N_11335);
nor U11702 (N_11702,N_11595,N_11238);
and U11703 (N_11703,N_11527,N_11572);
xor U11704 (N_11704,N_11252,N_11338);
nor U11705 (N_11705,N_11243,N_11581);
or U11706 (N_11706,N_11500,N_11533);
nand U11707 (N_11707,N_11467,N_11230);
or U11708 (N_11708,N_11431,N_11473);
nor U11709 (N_11709,N_11536,N_11324);
or U11710 (N_11710,N_11513,N_11598);
xor U11711 (N_11711,N_11531,N_11522);
and U11712 (N_11712,N_11372,N_11509);
and U11713 (N_11713,N_11296,N_11422);
nor U11714 (N_11714,N_11406,N_11506);
and U11715 (N_11715,N_11322,N_11563);
xnor U11716 (N_11716,N_11571,N_11379);
nor U11717 (N_11717,N_11229,N_11276);
nand U11718 (N_11718,N_11299,N_11386);
nand U11719 (N_11719,N_11265,N_11366);
nand U11720 (N_11720,N_11478,N_11361);
xnor U11721 (N_11721,N_11591,N_11259);
or U11722 (N_11722,N_11211,N_11239);
nand U11723 (N_11723,N_11451,N_11525);
xor U11724 (N_11724,N_11250,N_11452);
nand U11725 (N_11725,N_11367,N_11479);
nor U11726 (N_11726,N_11353,N_11375);
or U11727 (N_11727,N_11599,N_11320);
or U11728 (N_11728,N_11330,N_11458);
and U11729 (N_11729,N_11337,N_11317);
and U11730 (N_11730,N_11468,N_11288);
or U11731 (N_11731,N_11390,N_11586);
xnor U11732 (N_11732,N_11489,N_11368);
nand U11733 (N_11733,N_11302,N_11480);
nand U11734 (N_11734,N_11394,N_11555);
or U11735 (N_11735,N_11310,N_11496);
nor U11736 (N_11736,N_11582,N_11398);
nand U11737 (N_11737,N_11325,N_11224);
or U11738 (N_11738,N_11504,N_11393);
nand U11739 (N_11739,N_11501,N_11597);
or U11740 (N_11740,N_11204,N_11516);
and U11741 (N_11741,N_11280,N_11271);
nor U11742 (N_11742,N_11370,N_11544);
nor U11743 (N_11743,N_11262,N_11293);
xor U11744 (N_11744,N_11220,N_11484);
nand U11745 (N_11745,N_11282,N_11217);
and U11746 (N_11746,N_11534,N_11237);
xor U11747 (N_11747,N_11357,N_11354);
nor U11748 (N_11748,N_11414,N_11345);
nand U11749 (N_11749,N_11305,N_11397);
nor U11750 (N_11750,N_11212,N_11247);
or U11751 (N_11751,N_11492,N_11447);
or U11752 (N_11752,N_11437,N_11434);
nor U11753 (N_11753,N_11399,N_11475);
and U11754 (N_11754,N_11246,N_11365);
and U11755 (N_11755,N_11518,N_11448);
and U11756 (N_11756,N_11426,N_11385);
or U11757 (N_11757,N_11284,N_11587);
xnor U11758 (N_11758,N_11453,N_11493);
xnor U11759 (N_11759,N_11214,N_11477);
and U11760 (N_11760,N_11490,N_11234);
nand U11761 (N_11761,N_11270,N_11304);
nand U11762 (N_11762,N_11556,N_11389);
nor U11763 (N_11763,N_11521,N_11314);
nand U11764 (N_11764,N_11560,N_11291);
nand U11765 (N_11765,N_11380,N_11465);
xor U11766 (N_11766,N_11416,N_11583);
or U11767 (N_11767,N_11266,N_11300);
or U11768 (N_11768,N_11433,N_11359);
nand U11769 (N_11769,N_11218,N_11226);
nor U11770 (N_11770,N_11292,N_11236);
or U11771 (N_11771,N_11278,N_11318);
xnor U11772 (N_11772,N_11298,N_11542);
or U11773 (N_11773,N_11449,N_11499);
nor U11774 (N_11774,N_11312,N_11356);
xor U11775 (N_11775,N_11241,N_11374);
nor U11776 (N_11776,N_11430,N_11415);
nor U11777 (N_11777,N_11454,N_11559);
and U11778 (N_11778,N_11476,N_11364);
nand U11779 (N_11779,N_11435,N_11580);
xor U11780 (N_11780,N_11267,N_11584);
nand U11781 (N_11781,N_11532,N_11362);
or U11782 (N_11782,N_11553,N_11417);
or U11783 (N_11783,N_11260,N_11425);
xnor U11784 (N_11784,N_11502,N_11442);
or U11785 (N_11785,N_11450,N_11471);
nand U11786 (N_11786,N_11444,N_11567);
and U11787 (N_11787,N_11272,N_11336);
xor U11788 (N_11788,N_11579,N_11349);
nand U11789 (N_11789,N_11432,N_11269);
nor U11790 (N_11790,N_11232,N_11200);
nand U11791 (N_11791,N_11401,N_11408);
or U11792 (N_11792,N_11258,N_11464);
nand U11793 (N_11793,N_11546,N_11588);
or U11794 (N_11794,N_11589,N_11301);
or U11795 (N_11795,N_11334,N_11592);
nor U11796 (N_11796,N_11519,N_11346);
or U11797 (N_11797,N_11391,N_11341);
xnor U11798 (N_11798,N_11207,N_11457);
nand U11799 (N_11799,N_11535,N_11377);
nor U11800 (N_11800,N_11288,N_11278);
and U11801 (N_11801,N_11412,N_11523);
xnor U11802 (N_11802,N_11279,N_11546);
nor U11803 (N_11803,N_11458,N_11386);
and U11804 (N_11804,N_11491,N_11266);
xor U11805 (N_11805,N_11522,N_11552);
or U11806 (N_11806,N_11560,N_11483);
and U11807 (N_11807,N_11491,N_11563);
and U11808 (N_11808,N_11473,N_11589);
or U11809 (N_11809,N_11502,N_11445);
nand U11810 (N_11810,N_11432,N_11563);
xor U11811 (N_11811,N_11333,N_11435);
nand U11812 (N_11812,N_11475,N_11407);
xor U11813 (N_11813,N_11200,N_11252);
xor U11814 (N_11814,N_11245,N_11516);
or U11815 (N_11815,N_11552,N_11419);
or U11816 (N_11816,N_11577,N_11258);
nand U11817 (N_11817,N_11542,N_11551);
nand U11818 (N_11818,N_11289,N_11290);
nor U11819 (N_11819,N_11353,N_11200);
and U11820 (N_11820,N_11552,N_11232);
and U11821 (N_11821,N_11218,N_11478);
or U11822 (N_11822,N_11475,N_11372);
or U11823 (N_11823,N_11598,N_11425);
or U11824 (N_11824,N_11425,N_11561);
and U11825 (N_11825,N_11557,N_11460);
or U11826 (N_11826,N_11320,N_11391);
nor U11827 (N_11827,N_11355,N_11412);
nand U11828 (N_11828,N_11414,N_11529);
xnor U11829 (N_11829,N_11599,N_11237);
and U11830 (N_11830,N_11261,N_11527);
or U11831 (N_11831,N_11362,N_11446);
or U11832 (N_11832,N_11349,N_11413);
and U11833 (N_11833,N_11513,N_11462);
nand U11834 (N_11834,N_11375,N_11220);
nand U11835 (N_11835,N_11397,N_11595);
or U11836 (N_11836,N_11559,N_11297);
nor U11837 (N_11837,N_11481,N_11500);
xnor U11838 (N_11838,N_11482,N_11330);
nor U11839 (N_11839,N_11522,N_11241);
nand U11840 (N_11840,N_11204,N_11539);
and U11841 (N_11841,N_11509,N_11204);
nor U11842 (N_11842,N_11345,N_11227);
nor U11843 (N_11843,N_11563,N_11428);
nand U11844 (N_11844,N_11393,N_11577);
nand U11845 (N_11845,N_11241,N_11259);
nor U11846 (N_11846,N_11583,N_11484);
and U11847 (N_11847,N_11301,N_11310);
and U11848 (N_11848,N_11434,N_11514);
and U11849 (N_11849,N_11300,N_11466);
nor U11850 (N_11850,N_11398,N_11332);
and U11851 (N_11851,N_11305,N_11248);
or U11852 (N_11852,N_11213,N_11355);
xnor U11853 (N_11853,N_11280,N_11479);
or U11854 (N_11854,N_11209,N_11200);
nor U11855 (N_11855,N_11296,N_11598);
and U11856 (N_11856,N_11583,N_11207);
or U11857 (N_11857,N_11431,N_11322);
xor U11858 (N_11858,N_11270,N_11407);
and U11859 (N_11859,N_11546,N_11438);
or U11860 (N_11860,N_11308,N_11299);
and U11861 (N_11861,N_11250,N_11238);
nor U11862 (N_11862,N_11527,N_11289);
or U11863 (N_11863,N_11484,N_11390);
nor U11864 (N_11864,N_11593,N_11542);
xor U11865 (N_11865,N_11484,N_11346);
or U11866 (N_11866,N_11558,N_11313);
xnor U11867 (N_11867,N_11296,N_11242);
nor U11868 (N_11868,N_11421,N_11268);
and U11869 (N_11869,N_11593,N_11401);
nand U11870 (N_11870,N_11241,N_11322);
nand U11871 (N_11871,N_11569,N_11415);
nor U11872 (N_11872,N_11528,N_11574);
and U11873 (N_11873,N_11476,N_11316);
and U11874 (N_11874,N_11261,N_11571);
or U11875 (N_11875,N_11511,N_11371);
nand U11876 (N_11876,N_11337,N_11486);
or U11877 (N_11877,N_11528,N_11594);
xnor U11878 (N_11878,N_11563,N_11401);
and U11879 (N_11879,N_11390,N_11391);
xnor U11880 (N_11880,N_11366,N_11595);
nor U11881 (N_11881,N_11204,N_11482);
or U11882 (N_11882,N_11505,N_11271);
nand U11883 (N_11883,N_11298,N_11258);
and U11884 (N_11884,N_11382,N_11396);
xnor U11885 (N_11885,N_11485,N_11261);
and U11886 (N_11886,N_11294,N_11478);
nor U11887 (N_11887,N_11430,N_11448);
xnor U11888 (N_11888,N_11276,N_11559);
xor U11889 (N_11889,N_11522,N_11343);
nor U11890 (N_11890,N_11517,N_11406);
xnor U11891 (N_11891,N_11522,N_11350);
nor U11892 (N_11892,N_11283,N_11576);
nand U11893 (N_11893,N_11557,N_11234);
xor U11894 (N_11894,N_11538,N_11413);
or U11895 (N_11895,N_11464,N_11591);
xnor U11896 (N_11896,N_11532,N_11516);
nor U11897 (N_11897,N_11525,N_11536);
or U11898 (N_11898,N_11324,N_11425);
and U11899 (N_11899,N_11313,N_11266);
nand U11900 (N_11900,N_11450,N_11513);
nand U11901 (N_11901,N_11246,N_11256);
or U11902 (N_11902,N_11325,N_11335);
and U11903 (N_11903,N_11393,N_11557);
and U11904 (N_11904,N_11272,N_11352);
and U11905 (N_11905,N_11236,N_11403);
or U11906 (N_11906,N_11467,N_11415);
nor U11907 (N_11907,N_11582,N_11218);
xor U11908 (N_11908,N_11289,N_11405);
nor U11909 (N_11909,N_11449,N_11280);
xnor U11910 (N_11910,N_11515,N_11216);
nand U11911 (N_11911,N_11368,N_11541);
nor U11912 (N_11912,N_11348,N_11503);
or U11913 (N_11913,N_11303,N_11382);
xor U11914 (N_11914,N_11295,N_11591);
xnor U11915 (N_11915,N_11327,N_11574);
or U11916 (N_11916,N_11371,N_11339);
or U11917 (N_11917,N_11491,N_11596);
nor U11918 (N_11918,N_11474,N_11379);
and U11919 (N_11919,N_11377,N_11299);
nor U11920 (N_11920,N_11594,N_11320);
xor U11921 (N_11921,N_11562,N_11410);
nor U11922 (N_11922,N_11460,N_11455);
nor U11923 (N_11923,N_11356,N_11261);
and U11924 (N_11924,N_11436,N_11274);
nand U11925 (N_11925,N_11568,N_11431);
or U11926 (N_11926,N_11205,N_11246);
nand U11927 (N_11927,N_11597,N_11374);
and U11928 (N_11928,N_11437,N_11405);
and U11929 (N_11929,N_11369,N_11450);
nor U11930 (N_11930,N_11294,N_11489);
xor U11931 (N_11931,N_11357,N_11299);
nor U11932 (N_11932,N_11437,N_11490);
or U11933 (N_11933,N_11336,N_11329);
and U11934 (N_11934,N_11378,N_11325);
or U11935 (N_11935,N_11307,N_11537);
or U11936 (N_11936,N_11532,N_11570);
nor U11937 (N_11937,N_11595,N_11478);
nor U11938 (N_11938,N_11571,N_11206);
nand U11939 (N_11939,N_11304,N_11470);
nand U11940 (N_11940,N_11432,N_11422);
nor U11941 (N_11941,N_11238,N_11559);
nand U11942 (N_11942,N_11400,N_11506);
or U11943 (N_11943,N_11350,N_11396);
nor U11944 (N_11944,N_11455,N_11572);
and U11945 (N_11945,N_11208,N_11271);
xnor U11946 (N_11946,N_11581,N_11498);
xnor U11947 (N_11947,N_11372,N_11322);
xnor U11948 (N_11948,N_11315,N_11414);
nor U11949 (N_11949,N_11421,N_11248);
and U11950 (N_11950,N_11505,N_11502);
or U11951 (N_11951,N_11449,N_11396);
and U11952 (N_11952,N_11477,N_11490);
and U11953 (N_11953,N_11539,N_11310);
xor U11954 (N_11954,N_11221,N_11397);
or U11955 (N_11955,N_11206,N_11280);
xor U11956 (N_11956,N_11452,N_11469);
or U11957 (N_11957,N_11229,N_11509);
nor U11958 (N_11958,N_11382,N_11224);
and U11959 (N_11959,N_11371,N_11284);
xor U11960 (N_11960,N_11442,N_11532);
xnor U11961 (N_11961,N_11268,N_11293);
xnor U11962 (N_11962,N_11567,N_11255);
xnor U11963 (N_11963,N_11429,N_11270);
or U11964 (N_11964,N_11386,N_11551);
and U11965 (N_11965,N_11310,N_11238);
nand U11966 (N_11966,N_11230,N_11392);
and U11967 (N_11967,N_11224,N_11366);
and U11968 (N_11968,N_11509,N_11450);
or U11969 (N_11969,N_11483,N_11555);
nand U11970 (N_11970,N_11284,N_11257);
xor U11971 (N_11971,N_11396,N_11560);
and U11972 (N_11972,N_11364,N_11369);
or U11973 (N_11973,N_11423,N_11246);
nand U11974 (N_11974,N_11210,N_11205);
nand U11975 (N_11975,N_11338,N_11450);
nand U11976 (N_11976,N_11264,N_11576);
nand U11977 (N_11977,N_11347,N_11559);
xnor U11978 (N_11978,N_11485,N_11437);
and U11979 (N_11979,N_11382,N_11598);
nor U11980 (N_11980,N_11518,N_11354);
nand U11981 (N_11981,N_11237,N_11586);
or U11982 (N_11982,N_11467,N_11513);
xnor U11983 (N_11983,N_11271,N_11501);
nand U11984 (N_11984,N_11480,N_11495);
or U11985 (N_11985,N_11246,N_11472);
nor U11986 (N_11986,N_11359,N_11579);
and U11987 (N_11987,N_11499,N_11330);
nand U11988 (N_11988,N_11340,N_11237);
or U11989 (N_11989,N_11328,N_11284);
or U11990 (N_11990,N_11303,N_11264);
and U11991 (N_11991,N_11308,N_11382);
nor U11992 (N_11992,N_11530,N_11479);
and U11993 (N_11993,N_11570,N_11515);
and U11994 (N_11994,N_11320,N_11409);
nand U11995 (N_11995,N_11361,N_11488);
or U11996 (N_11996,N_11570,N_11555);
and U11997 (N_11997,N_11392,N_11483);
or U11998 (N_11998,N_11526,N_11444);
or U11999 (N_11999,N_11294,N_11350);
and U12000 (N_12000,N_11852,N_11975);
nand U12001 (N_12001,N_11986,N_11941);
xor U12002 (N_12002,N_11644,N_11711);
and U12003 (N_12003,N_11972,N_11656);
or U12004 (N_12004,N_11691,N_11912);
nor U12005 (N_12005,N_11672,N_11609);
xor U12006 (N_12006,N_11779,N_11903);
or U12007 (N_12007,N_11914,N_11991);
nand U12008 (N_12008,N_11771,N_11622);
nor U12009 (N_12009,N_11736,N_11824);
nand U12010 (N_12010,N_11806,N_11785);
or U12011 (N_12011,N_11643,N_11885);
and U12012 (N_12012,N_11620,N_11863);
nor U12013 (N_12013,N_11758,N_11678);
xnor U12014 (N_12014,N_11772,N_11807);
or U12015 (N_12015,N_11796,N_11786);
nand U12016 (N_12016,N_11649,N_11693);
and U12017 (N_12017,N_11831,N_11982);
nor U12018 (N_12018,N_11784,N_11640);
nor U12019 (N_12019,N_11613,N_11993);
or U12020 (N_12020,N_11989,N_11653);
and U12021 (N_12021,N_11834,N_11945);
and U12022 (N_12022,N_11988,N_11902);
and U12023 (N_12023,N_11837,N_11781);
or U12024 (N_12024,N_11857,N_11789);
xor U12025 (N_12025,N_11913,N_11616);
or U12026 (N_12026,N_11662,N_11985);
and U12027 (N_12027,N_11980,N_11900);
xor U12028 (N_12028,N_11718,N_11719);
nor U12029 (N_12029,N_11812,N_11872);
or U12030 (N_12030,N_11926,N_11753);
and U12031 (N_12031,N_11710,N_11652);
nor U12032 (N_12032,N_11998,N_11859);
xor U12033 (N_12033,N_11706,N_11875);
and U12034 (N_12034,N_11723,N_11610);
nor U12035 (N_12035,N_11897,N_11792);
nor U12036 (N_12036,N_11670,N_11651);
or U12037 (N_12037,N_11729,N_11970);
xor U12038 (N_12038,N_11948,N_11790);
nor U12039 (N_12039,N_11987,N_11674);
nand U12040 (N_12040,N_11821,N_11878);
nand U12041 (N_12041,N_11833,N_11876);
nor U12042 (N_12042,N_11759,N_11804);
and U12043 (N_12043,N_11898,N_11770);
nor U12044 (N_12044,N_11740,N_11665);
and U12045 (N_12045,N_11793,N_11720);
and U12046 (N_12046,N_11782,N_11922);
nand U12047 (N_12047,N_11637,N_11827);
nand U12048 (N_12048,N_11996,N_11743);
nor U12049 (N_12049,N_11754,N_11777);
or U12050 (N_12050,N_11932,N_11936);
or U12051 (N_12051,N_11992,N_11605);
or U12052 (N_12052,N_11825,N_11874);
nand U12053 (N_12053,N_11843,N_11883);
nor U12054 (N_12054,N_11939,N_11961);
xor U12055 (N_12055,N_11911,N_11990);
nor U12056 (N_12056,N_11684,N_11886);
xnor U12057 (N_12057,N_11994,N_11664);
and U12058 (N_12058,N_11632,N_11847);
nor U12059 (N_12059,N_11697,N_11947);
or U12060 (N_12060,N_11713,N_11960);
xnor U12061 (N_12061,N_11663,N_11956);
or U12062 (N_12062,N_11611,N_11716);
and U12063 (N_12063,N_11867,N_11924);
nor U12064 (N_12064,N_11881,N_11943);
and U12065 (N_12065,N_11692,N_11695);
or U12066 (N_12066,N_11908,N_11675);
xor U12067 (N_12067,N_11602,N_11788);
or U12068 (N_12068,N_11820,N_11735);
or U12069 (N_12069,N_11894,N_11764);
nor U12070 (N_12070,N_11889,N_11851);
and U12071 (N_12071,N_11959,N_11891);
nand U12072 (N_12072,N_11714,N_11767);
xnor U12073 (N_12073,N_11836,N_11938);
nand U12074 (N_12074,N_11808,N_11813);
xor U12075 (N_12075,N_11751,N_11978);
and U12076 (N_12076,N_11686,N_11606);
and U12077 (N_12077,N_11888,N_11928);
or U12078 (N_12078,N_11968,N_11787);
or U12079 (N_12079,N_11603,N_11687);
nor U12080 (N_12080,N_11638,N_11668);
nand U12081 (N_12081,N_11797,N_11919);
or U12082 (N_12082,N_11701,N_11944);
and U12083 (N_12083,N_11794,N_11957);
or U12084 (N_12084,N_11634,N_11722);
xnor U12085 (N_12085,N_11811,N_11800);
nor U12086 (N_12086,N_11830,N_11738);
and U12087 (N_12087,N_11906,N_11636);
or U12088 (N_12088,N_11870,N_11858);
and U12089 (N_12089,N_11783,N_11745);
and U12090 (N_12090,N_11817,N_11739);
and U12091 (N_12091,N_11696,N_11890);
or U12092 (N_12092,N_11750,N_11884);
nor U12093 (N_12093,N_11935,N_11899);
or U12094 (N_12094,N_11742,N_11731);
and U12095 (N_12095,N_11642,N_11918);
and U12096 (N_12096,N_11677,N_11955);
nand U12097 (N_12097,N_11965,N_11844);
nand U12098 (N_12098,N_11694,N_11845);
and U12099 (N_12099,N_11765,N_11712);
nor U12100 (N_12100,N_11882,N_11966);
xor U12101 (N_12101,N_11657,N_11953);
nand U12102 (N_12102,N_11964,N_11614);
nor U12103 (N_12103,N_11815,N_11828);
and U12104 (N_12104,N_11973,N_11930);
nand U12105 (N_12105,N_11608,N_11698);
nor U12106 (N_12106,N_11658,N_11755);
nand U12107 (N_12107,N_11703,N_11809);
or U12108 (N_12108,N_11839,N_11958);
and U12109 (N_12109,N_11627,N_11680);
or U12110 (N_12110,N_11976,N_11774);
nand U12111 (N_12111,N_11921,N_11682);
or U12112 (N_12112,N_11917,N_11814);
xnor U12113 (N_12113,N_11923,N_11866);
nor U12114 (N_12114,N_11717,N_11910);
xnor U12115 (N_12115,N_11660,N_11818);
nand U12116 (N_12116,N_11725,N_11934);
or U12117 (N_12117,N_11892,N_11734);
nand U12118 (N_12118,N_11756,N_11689);
nor U12119 (N_12119,N_11633,N_11728);
and U12120 (N_12120,N_11671,N_11877);
and U12121 (N_12121,N_11940,N_11679);
nand U12122 (N_12122,N_11915,N_11984);
and U12123 (N_12123,N_11775,N_11927);
nor U12124 (N_12124,N_11810,N_11648);
or U12125 (N_12125,N_11749,N_11974);
or U12126 (N_12126,N_11954,N_11816);
and U12127 (N_12127,N_11741,N_11952);
and U12128 (N_12128,N_11925,N_11893);
xnor U12129 (N_12129,N_11688,N_11766);
xor U12130 (N_12130,N_11748,N_11655);
xnor U12131 (N_12131,N_11916,N_11683);
nor U12132 (N_12132,N_11600,N_11624);
nand U12133 (N_12133,N_11829,N_11909);
and U12134 (N_12134,N_11744,N_11631);
and U12135 (N_12135,N_11879,N_11690);
nor U12136 (N_12136,N_11971,N_11715);
xor U12137 (N_12137,N_11981,N_11659);
or U12138 (N_12138,N_11746,N_11641);
or U12139 (N_12139,N_11907,N_11646);
and U12140 (N_12140,N_11773,N_11838);
nor U12141 (N_12141,N_11861,N_11681);
or U12142 (N_12142,N_11880,N_11760);
nand U12143 (N_12143,N_11769,N_11856);
and U12144 (N_12144,N_11799,N_11629);
or U12145 (N_12145,N_11645,N_11702);
nand U12146 (N_12146,N_11933,N_11607);
xnor U12147 (N_12147,N_11826,N_11650);
nand U12148 (N_12148,N_11798,N_11778);
and U12149 (N_12149,N_11623,N_11840);
nand U12150 (N_12150,N_11937,N_11647);
and U12151 (N_12151,N_11967,N_11950);
nand U12152 (N_12152,N_11865,N_11776);
nand U12153 (N_12153,N_11667,N_11639);
or U12154 (N_12154,N_11803,N_11848);
xor U12155 (N_12155,N_11707,N_11801);
xnor U12156 (N_12156,N_11855,N_11854);
nor U12157 (N_12157,N_11846,N_11604);
nand U12158 (N_12158,N_11995,N_11673);
nand U12159 (N_12159,N_11795,N_11850);
nand U12160 (N_12160,N_11724,N_11887);
xnor U12161 (N_12161,N_11628,N_11737);
nand U12162 (N_12162,N_11802,N_11705);
nand U12163 (N_12163,N_11615,N_11669);
xnor U12164 (N_12164,N_11904,N_11626);
xor U12165 (N_12165,N_11977,N_11979);
nand U12166 (N_12166,N_11685,N_11618);
nor U12167 (N_12167,N_11619,N_11832);
nor U12168 (N_12168,N_11661,N_11727);
nor U12169 (N_12169,N_11730,N_11666);
xnor U12170 (N_12170,N_11969,N_11871);
or U12171 (N_12171,N_11822,N_11997);
nand U12172 (N_12172,N_11849,N_11868);
nand U12173 (N_12173,N_11704,N_11732);
nor U12174 (N_12174,N_11612,N_11931);
xor U12175 (N_12175,N_11752,N_11835);
and U12176 (N_12176,N_11962,N_11920);
xor U12177 (N_12177,N_11700,N_11726);
nand U12178 (N_12178,N_11819,N_11761);
and U12179 (N_12179,N_11708,N_11617);
nand U12180 (N_12180,N_11896,N_11901);
nand U12181 (N_12181,N_11676,N_11805);
nand U12182 (N_12182,N_11630,N_11721);
or U12183 (N_12183,N_11601,N_11949);
xor U12184 (N_12184,N_11946,N_11942);
nand U12185 (N_12185,N_11762,N_11983);
nand U12186 (N_12186,N_11862,N_11873);
xor U12187 (N_12187,N_11905,N_11823);
xor U12188 (N_12188,N_11757,N_11963);
nor U12189 (N_12189,N_11654,N_11841);
or U12190 (N_12190,N_11864,N_11709);
xor U12191 (N_12191,N_11999,N_11699);
nor U12192 (N_12192,N_11733,N_11768);
and U12193 (N_12193,N_11860,N_11842);
nor U12194 (N_12194,N_11929,N_11747);
nor U12195 (N_12195,N_11869,N_11853);
nand U12196 (N_12196,N_11621,N_11625);
and U12197 (N_12197,N_11763,N_11895);
and U12198 (N_12198,N_11951,N_11791);
or U12199 (N_12199,N_11780,N_11635);
and U12200 (N_12200,N_11651,N_11776);
xor U12201 (N_12201,N_11691,N_11729);
and U12202 (N_12202,N_11747,N_11789);
nand U12203 (N_12203,N_11884,N_11622);
nor U12204 (N_12204,N_11753,N_11678);
nand U12205 (N_12205,N_11995,N_11703);
or U12206 (N_12206,N_11935,N_11951);
nand U12207 (N_12207,N_11845,N_11786);
xnor U12208 (N_12208,N_11603,N_11784);
nor U12209 (N_12209,N_11862,N_11644);
and U12210 (N_12210,N_11735,N_11908);
or U12211 (N_12211,N_11973,N_11843);
or U12212 (N_12212,N_11870,N_11696);
and U12213 (N_12213,N_11929,N_11836);
nand U12214 (N_12214,N_11691,N_11856);
nor U12215 (N_12215,N_11786,N_11826);
xor U12216 (N_12216,N_11926,N_11755);
and U12217 (N_12217,N_11660,N_11762);
xor U12218 (N_12218,N_11645,N_11740);
nor U12219 (N_12219,N_11641,N_11630);
nand U12220 (N_12220,N_11825,N_11762);
xor U12221 (N_12221,N_11687,N_11920);
nor U12222 (N_12222,N_11828,N_11630);
nand U12223 (N_12223,N_11606,N_11896);
and U12224 (N_12224,N_11666,N_11715);
or U12225 (N_12225,N_11686,N_11790);
nor U12226 (N_12226,N_11961,N_11691);
and U12227 (N_12227,N_11669,N_11892);
or U12228 (N_12228,N_11778,N_11659);
or U12229 (N_12229,N_11689,N_11671);
or U12230 (N_12230,N_11985,N_11689);
and U12231 (N_12231,N_11681,N_11860);
nor U12232 (N_12232,N_11970,N_11638);
or U12233 (N_12233,N_11615,N_11603);
nand U12234 (N_12234,N_11916,N_11690);
and U12235 (N_12235,N_11632,N_11618);
and U12236 (N_12236,N_11683,N_11840);
nor U12237 (N_12237,N_11932,N_11738);
or U12238 (N_12238,N_11621,N_11907);
nand U12239 (N_12239,N_11808,N_11715);
or U12240 (N_12240,N_11982,N_11663);
or U12241 (N_12241,N_11990,N_11895);
or U12242 (N_12242,N_11654,N_11739);
nand U12243 (N_12243,N_11938,N_11757);
nor U12244 (N_12244,N_11974,N_11686);
or U12245 (N_12245,N_11822,N_11962);
xor U12246 (N_12246,N_11984,N_11941);
nand U12247 (N_12247,N_11737,N_11798);
or U12248 (N_12248,N_11691,N_11843);
nor U12249 (N_12249,N_11826,N_11763);
nand U12250 (N_12250,N_11781,N_11698);
xor U12251 (N_12251,N_11909,N_11904);
nor U12252 (N_12252,N_11764,N_11653);
or U12253 (N_12253,N_11679,N_11846);
xor U12254 (N_12254,N_11623,N_11967);
and U12255 (N_12255,N_11847,N_11946);
nor U12256 (N_12256,N_11961,N_11942);
xnor U12257 (N_12257,N_11845,N_11789);
nor U12258 (N_12258,N_11944,N_11860);
xnor U12259 (N_12259,N_11940,N_11923);
or U12260 (N_12260,N_11714,N_11878);
or U12261 (N_12261,N_11939,N_11680);
or U12262 (N_12262,N_11962,N_11855);
nand U12263 (N_12263,N_11826,N_11893);
nand U12264 (N_12264,N_11704,N_11611);
and U12265 (N_12265,N_11635,N_11748);
xor U12266 (N_12266,N_11875,N_11999);
nand U12267 (N_12267,N_11694,N_11691);
nor U12268 (N_12268,N_11812,N_11902);
xor U12269 (N_12269,N_11671,N_11620);
or U12270 (N_12270,N_11674,N_11818);
nand U12271 (N_12271,N_11993,N_11982);
xnor U12272 (N_12272,N_11871,N_11688);
or U12273 (N_12273,N_11859,N_11796);
and U12274 (N_12274,N_11871,N_11747);
and U12275 (N_12275,N_11627,N_11879);
and U12276 (N_12276,N_11768,N_11623);
xnor U12277 (N_12277,N_11925,N_11675);
xnor U12278 (N_12278,N_11937,N_11674);
nor U12279 (N_12279,N_11771,N_11862);
and U12280 (N_12280,N_11624,N_11725);
nor U12281 (N_12281,N_11781,N_11622);
xnor U12282 (N_12282,N_11808,N_11706);
nand U12283 (N_12283,N_11718,N_11821);
nand U12284 (N_12284,N_11778,N_11764);
nand U12285 (N_12285,N_11674,N_11943);
nor U12286 (N_12286,N_11710,N_11910);
or U12287 (N_12287,N_11667,N_11786);
xor U12288 (N_12288,N_11819,N_11884);
and U12289 (N_12289,N_11666,N_11871);
nand U12290 (N_12290,N_11652,N_11864);
nor U12291 (N_12291,N_11648,N_11825);
and U12292 (N_12292,N_11947,N_11962);
nand U12293 (N_12293,N_11700,N_11904);
nand U12294 (N_12294,N_11719,N_11630);
nor U12295 (N_12295,N_11870,N_11712);
nand U12296 (N_12296,N_11917,N_11742);
and U12297 (N_12297,N_11706,N_11690);
nor U12298 (N_12298,N_11657,N_11915);
or U12299 (N_12299,N_11945,N_11883);
xnor U12300 (N_12300,N_11774,N_11884);
xor U12301 (N_12301,N_11989,N_11987);
xnor U12302 (N_12302,N_11674,N_11961);
nand U12303 (N_12303,N_11616,N_11626);
or U12304 (N_12304,N_11609,N_11715);
and U12305 (N_12305,N_11796,N_11983);
and U12306 (N_12306,N_11709,N_11676);
xor U12307 (N_12307,N_11607,N_11706);
nor U12308 (N_12308,N_11785,N_11990);
xnor U12309 (N_12309,N_11978,N_11973);
xor U12310 (N_12310,N_11601,N_11861);
nand U12311 (N_12311,N_11761,N_11736);
nor U12312 (N_12312,N_11918,N_11771);
or U12313 (N_12313,N_11929,N_11746);
nand U12314 (N_12314,N_11652,N_11781);
or U12315 (N_12315,N_11715,N_11683);
and U12316 (N_12316,N_11653,N_11929);
and U12317 (N_12317,N_11859,N_11745);
nand U12318 (N_12318,N_11768,N_11740);
nor U12319 (N_12319,N_11635,N_11987);
and U12320 (N_12320,N_11751,N_11699);
nor U12321 (N_12321,N_11633,N_11635);
nand U12322 (N_12322,N_11860,N_11779);
nor U12323 (N_12323,N_11814,N_11637);
nand U12324 (N_12324,N_11745,N_11655);
xnor U12325 (N_12325,N_11830,N_11618);
nand U12326 (N_12326,N_11642,N_11928);
nor U12327 (N_12327,N_11693,N_11959);
or U12328 (N_12328,N_11963,N_11830);
and U12329 (N_12329,N_11869,N_11630);
nand U12330 (N_12330,N_11740,N_11631);
nor U12331 (N_12331,N_11763,N_11874);
and U12332 (N_12332,N_11866,N_11728);
or U12333 (N_12333,N_11974,N_11603);
xor U12334 (N_12334,N_11657,N_11619);
or U12335 (N_12335,N_11809,N_11987);
or U12336 (N_12336,N_11720,N_11757);
xnor U12337 (N_12337,N_11778,N_11815);
xor U12338 (N_12338,N_11704,N_11877);
nor U12339 (N_12339,N_11696,N_11650);
xor U12340 (N_12340,N_11956,N_11764);
nor U12341 (N_12341,N_11646,N_11726);
xnor U12342 (N_12342,N_11879,N_11742);
or U12343 (N_12343,N_11869,N_11635);
nor U12344 (N_12344,N_11637,N_11618);
and U12345 (N_12345,N_11670,N_11721);
nor U12346 (N_12346,N_11937,N_11680);
xnor U12347 (N_12347,N_11816,N_11622);
or U12348 (N_12348,N_11781,N_11744);
or U12349 (N_12349,N_11888,N_11982);
nand U12350 (N_12350,N_11730,N_11781);
xnor U12351 (N_12351,N_11967,N_11848);
and U12352 (N_12352,N_11674,N_11670);
xnor U12353 (N_12353,N_11919,N_11986);
xnor U12354 (N_12354,N_11831,N_11732);
nand U12355 (N_12355,N_11888,N_11768);
or U12356 (N_12356,N_11760,N_11730);
and U12357 (N_12357,N_11786,N_11648);
or U12358 (N_12358,N_11834,N_11948);
xor U12359 (N_12359,N_11615,N_11878);
nand U12360 (N_12360,N_11974,N_11936);
nor U12361 (N_12361,N_11727,N_11765);
xnor U12362 (N_12362,N_11800,N_11662);
nor U12363 (N_12363,N_11636,N_11815);
xnor U12364 (N_12364,N_11858,N_11881);
xor U12365 (N_12365,N_11600,N_11933);
xnor U12366 (N_12366,N_11934,N_11957);
xnor U12367 (N_12367,N_11798,N_11955);
xor U12368 (N_12368,N_11668,N_11783);
and U12369 (N_12369,N_11800,N_11859);
nand U12370 (N_12370,N_11770,N_11779);
nor U12371 (N_12371,N_11944,N_11764);
xor U12372 (N_12372,N_11787,N_11839);
nand U12373 (N_12373,N_11833,N_11708);
or U12374 (N_12374,N_11672,N_11687);
nor U12375 (N_12375,N_11908,N_11893);
and U12376 (N_12376,N_11988,N_11931);
xnor U12377 (N_12377,N_11807,N_11606);
nand U12378 (N_12378,N_11903,N_11717);
xnor U12379 (N_12379,N_11912,N_11954);
and U12380 (N_12380,N_11958,N_11654);
nor U12381 (N_12381,N_11635,N_11876);
or U12382 (N_12382,N_11697,N_11737);
or U12383 (N_12383,N_11648,N_11991);
nor U12384 (N_12384,N_11841,N_11934);
nand U12385 (N_12385,N_11858,N_11836);
nor U12386 (N_12386,N_11725,N_11908);
nor U12387 (N_12387,N_11996,N_11951);
or U12388 (N_12388,N_11803,N_11743);
nand U12389 (N_12389,N_11643,N_11987);
xor U12390 (N_12390,N_11662,N_11795);
or U12391 (N_12391,N_11788,N_11820);
or U12392 (N_12392,N_11959,N_11892);
nor U12393 (N_12393,N_11611,N_11634);
nor U12394 (N_12394,N_11674,N_11779);
nand U12395 (N_12395,N_11977,N_11618);
nand U12396 (N_12396,N_11916,N_11966);
or U12397 (N_12397,N_11988,N_11986);
and U12398 (N_12398,N_11910,N_11689);
and U12399 (N_12399,N_11855,N_11824);
nand U12400 (N_12400,N_12210,N_12248);
or U12401 (N_12401,N_12020,N_12282);
and U12402 (N_12402,N_12025,N_12219);
or U12403 (N_12403,N_12368,N_12120);
and U12404 (N_12404,N_12389,N_12322);
and U12405 (N_12405,N_12174,N_12193);
or U12406 (N_12406,N_12233,N_12101);
nand U12407 (N_12407,N_12100,N_12222);
nand U12408 (N_12408,N_12060,N_12394);
nand U12409 (N_12409,N_12308,N_12034);
nor U12410 (N_12410,N_12142,N_12275);
or U12411 (N_12411,N_12170,N_12153);
nor U12412 (N_12412,N_12183,N_12220);
nor U12413 (N_12413,N_12125,N_12281);
nor U12414 (N_12414,N_12068,N_12397);
nor U12415 (N_12415,N_12190,N_12381);
nand U12416 (N_12416,N_12301,N_12070);
xnor U12417 (N_12417,N_12332,N_12307);
nand U12418 (N_12418,N_12265,N_12221);
or U12419 (N_12419,N_12270,N_12376);
nor U12420 (N_12420,N_12096,N_12379);
or U12421 (N_12421,N_12132,N_12319);
xor U12422 (N_12422,N_12127,N_12392);
or U12423 (N_12423,N_12296,N_12147);
nor U12424 (N_12424,N_12216,N_12202);
xor U12425 (N_12425,N_12110,N_12330);
nand U12426 (N_12426,N_12338,N_12178);
nand U12427 (N_12427,N_12244,N_12162);
or U12428 (N_12428,N_12357,N_12111);
and U12429 (N_12429,N_12294,N_12370);
nor U12430 (N_12430,N_12366,N_12138);
nor U12431 (N_12431,N_12093,N_12144);
or U12432 (N_12432,N_12195,N_12006);
or U12433 (N_12433,N_12327,N_12040);
or U12434 (N_12434,N_12230,N_12300);
nor U12435 (N_12435,N_12164,N_12215);
or U12436 (N_12436,N_12046,N_12361);
nor U12437 (N_12437,N_12390,N_12328);
and U12438 (N_12438,N_12158,N_12141);
nor U12439 (N_12439,N_12137,N_12066);
or U12440 (N_12440,N_12238,N_12228);
nor U12441 (N_12441,N_12155,N_12139);
or U12442 (N_12442,N_12283,N_12051);
nand U12443 (N_12443,N_12008,N_12041);
and U12444 (N_12444,N_12249,N_12026);
or U12445 (N_12445,N_12253,N_12395);
nor U12446 (N_12446,N_12117,N_12266);
nand U12447 (N_12447,N_12055,N_12004);
or U12448 (N_12448,N_12346,N_12204);
xor U12449 (N_12449,N_12354,N_12106);
nor U12450 (N_12450,N_12214,N_12022);
nor U12451 (N_12451,N_12149,N_12080);
and U12452 (N_12452,N_12028,N_12059);
nand U12453 (N_12453,N_12212,N_12385);
xor U12454 (N_12454,N_12045,N_12371);
and U12455 (N_12455,N_12269,N_12289);
nor U12456 (N_12456,N_12201,N_12262);
and U12457 (N_12457,N_12119,N_12373);
or U12458 (N_12458,N_12235,N_12049);
nor U12459 (N_12459,N_12131,N_12227);
nand U12460 (N_12460,N_12237,N_12350);
and U12461 (N_12461,N_12085,N_12200);
or U12462 (N_12462,N_12136,N_12116);
and U12463 (N_12463,N_12035,N_12165);
and U12464 (N_12464,N_12019,N_12166);
or U12465 (N_12465,N_12232,N_12287);
nor U12466 (N_12466,N_12240,N_12292);
and U12467 (N_12467,N_12115,N_12377);
nand U12468 (N_12468,N_12343,N_12391);
nand U12469 (N_12469,N_12172,N_12189);
nand U12470 (N_12470,N_12277,N_12134);
and U12471 (N_12471,N_12254,N_12077);
xor U12472 (N_12472,N_12358,N_12351);
nand U12473 (N_12473,N_12014,N_12316);
nor U12474 (N_12474,N_12314,N_12217);
nand U12475 (N_12475,N_12382,N_12191);
nor U12476 (N_12476,N_12205,N_12246);
nor U12477 (N_12477,N_12261,N_12364);
nand U12478 (N_12478,N_12029,N_12360);
xnor U12479 (N_12479,N_12298,N_12274);
nor U12480 (N_12480,N_12194,N_12126);
or U12481 (N_12481,N_12168,N_12239);
or U12482 (N_12482,N_12088,N_12092);
nand U12483 (N_12483,N_12304,N_12318);
and U12484 (N_12484,N_12245,N_12259);
xnor U12485 (N_12485,N_12387,N_12145);
xor U12486 (N_12486,N_12121,N_12039);
or U12487 (N_12487,N_12146,N_12310);
xnor U12488 (N_12488,N_12331,N_12355);
nand U12489 (N_12489,N_12352,N_12067);
or U12490 (N_12490,N_12181,N_12242);
and U12491 (N_12491,N_12344,N_12086);
nand U12492 (N_12492,N_12293,N_12148);
or U12493 (N_12493,N_12264,N_12347);
or U12494 (N_12494,N_12302,N_12323);
or U12495 (N_12495,N_12348,N_12184);
and U12496 (N_12496,N_12058,N_12023);
or U12497 (N_12497,N_12030,N_12072);
nand U12498 (N_12498,N_12396,N_12000);
or U12499 (N_12499,N_12208,N_12081);
and U12500 (N_12500,N_12130,N_12056);
or U12501 (N_12501,N_12231,N_12161);
and U12502 (N_12502,N_12295,N_12223);
and U12503 (N_12503,N_12384,N_12169);
or U12504 (N_12504,N_12209,N_12044);
nand U12505 (N_12505,N_12378,N_12114);
xnor U12506 (N_12506,N_12091,N_12353);
or U12507 (N_12507,N_12337,N_12124);
nand U12508 (N_12508,N_12156,N_12036);
and U12509 (N_12509,N_12150,N_12213);
nand U12510 (N_12510,N_12157,N_12263);
nor U12511 (N_12511,N_12197,N_12198);
and U12512 (N_12512,N_12179,N_12291);
and U12513 (N_12513,N_12069,N_12083);
and U12514 (N_12514,N_12324,N_12151);
nor U12515 (N_12515,N_12032,N_12065);
and U12516 (N_12516,N_12326,N_12186);
xnor U12517 (N_12517,N_12007,N_12226);
nor U12518 (N_12518,N_12313,N_12052);
nor U12519 (N_12519,N_12176,N_12342);
xnor U12520 (N_12520,N_12182,N_12105);
nor U12521 (N_12521,N_12011,N_12143);
and U12522 (N_12522,N_12001,N_12211);
or U12523 (N_12523,N_12053,N_12084);
nor U12524 (N_12524,N_12286,N_12188);
nor U12525 (N_12525,N_12251,N_12309);
or U12526 (N_12526,N_12071,N_12369);
nand U12527 (N_12527,N_12073,N_12280);
nor U12528 (N_12528,N_12002,N_12278);
nand U12529 (N_12529,N_12133,N_12118);
and U12530 (N_12530,N_12196,N_12393);
and U12531 (N_12531,N_12229,N_12128);
and U12532 (N_12532,N_12285,N_12163);
and U12533 (N_12533,N_12256,N_12271);
xor U12534 (N_12534,N_12374,N_12290);
or U12535 (N_12535,N_12013,N_12018);
or U12536 (N_12536,N_12003,N_12135);
xor U12537 (N_12537,N_12388,N_12383);
nand U12538 (N_12538,N_12255,N_12267);
and U12539 (N_12539,N_12123,N_12339);
xnor U12540 (N_12540,N_12129,N_12050);
or U12541 (N_12541,N_12345,N_12241);
nand U12542 (N_12542,N_12272,N_12021);
nor U12543 (N_12543,N_12187,N_12099);
xor U12544 (N_12544,N_12122,N_12033);
and U12545 (N_12545,N_12074,N_12037);
or U12546 (N_12546,N_12312,N_12103);
xnor U12547 (N_12547,N_12375,N_12024);
nand U12548 (N_12548,N_12365,N_12320);
xor U12549 (N_12549,N_12112,N_12082);
nor U12550 (N_12550,N_12064,N_12075);
xnor U12551 (N_12551,N_12311,N_12102);
nor U12552 (N_12552,N_12090,N_12257);
nor U12553 (N_12553,N_12224,N_12199);
nor U12554 (N_12554,N_12159,N_12284);
nand U12555 (N_12555,N_12340,N_12306);
and U12556 (N_12556,N_12333,N_12268);
and U12557 (N_12557,N_12325,N_12043);
and U12558 (N_12558,N_12288,N_12057);
and U12559 (N_12559,N_12017,N_12398);
nand U12560 (N_12560,N_12258,N_12010);
xnor U12561 (N_12561,N_12140,N_12154);
xnor U12562 (N_12562,N_12078,N_12107);
or U12563 (N_12563,N_12089,N_12372);
xor U12564 (N_12564,N_12336,N_12079);
or U12565 (N_12565,N_12273,N_12009);
and U12566 (N_12566,N_12367,N_12054);
xnor U12567 (N_12567,N_12362,N_12303);
and U12568 (N_12568,N_12276,N_12341);
or U12569 (N_12569,N_12097,N_12016);
and U12570 (N_12570,N_12063,N_12109);
xnor U12571 (N_12571,N_12012,N_12042);
xnor U12572 (N_12572,N_12218,N_12061);
xor U12573 (N_12573,N_12047,N_12203);
or U12574 (N_12574,N_12234,N_12152);
nor U12575 (N_12575,N_12048,N_12177);
nand U12576 (N_12576,N_12260,N_12250);
xnor U12577 (N_12577,N_12160,N_12236);
nand U12578 (N_12578,N_12321,N_12334);
xor U12579 (N_12579,N_12207,N_12087);
and U12580 (N_12580,N_12386,N_12297);
xor U12581 (N_12581,N_12363,N_12027);
nand U12582 (N_12582,N_12305,N_12185);
and U12583 (N_12583,N_12399,N_12031);
nand U12584 (N_12584,N_12095,N_12076);
nand U12585 (N_12585,N_12349,N_12247);
and U12586 (N_12586,N_12005,N_12113);
and U12587 (N_12587,N_12094,N_12225);
or U12588 (N_12588,N_12359,N_12173);
and U12589 (N_12589,N_12299,N_12167);
and U12590 (N_12590,N_12335,N_12279);
nor U12591 (N_12591,N_12015,N_12317);
nor U12592 (N_12592,N_12192,N_12171);
xnor U12593 (N_12593,N_12180,N_12252);
or U12594 (N_12594,N_12098,N_12380);
nand U12595 (N_12595,N_12038,N_12329);
nand U12596 (N_12596,N_12104,N_12062);
xor U12597 (N_12597,N_12356,N_12243);
xnor U12598 (N_12598,N_12108,N_12175);
and U12599 (N_12599,N_12315,N_12206);
xnor U12600 (N_12600,N_12211,N_12044);
and U12601 (N_12601,N_12173,N_12013);
xor U12602 (N_12602,N_12347,N_12268);
and U12603 (N_12603,N_12200,N_12282);
nor U12604 (N_12604,N_12049,N_12375);
xnor U12605 (N_12605,N_12262,N_12281);
nand U12606 (N_12606,N_12114,N_12150);
and U12607 (N_12607,N_12164,N_12111);
xnor U12608 (N_12608,N_12260,N_12353);
nor U12609 (N_12609,N_12257,N_12222);
nor U12610 (N_12610,N_12338,N_12301);
nand U12611 (N_12611,N_12119,N_12027);
nor U12612 (N_12612,N_12250,N_12263);
xor U12613 (N_12613,N_12324,N_12202);
nand U12614 (N_12614,N_12391,N_12056);
and U12615 (N_12615,N_12360,N_12092);
nand U12616 (N_12616,N_12073,N_12316);
nand U12617 (N_12617,N_12321,N_12319);
and U12618 (N_12618,N_12160,N_12264);
xnor U12619 (N_12619,N_12192,N_12135);
xor U12620 (N_12620,N_12085,N_12131);
nand U12621 (N_12621,N_12230,N_12399);
nand U12622 (N_12622,N_12115,N_12327);
nor U12623 (N_12623,N_12157,N_12383);
or U12624 (N_12624,N_12029,N_12332);
or U12625 (N_12625,N_12170,N_12368);
nor U12626 (N_12626,N_12024,N_12093);
nor U12627 (N_12627,N_12157,N_12363);
nor U12628 (N_12628,N_12022,N_12195);
xor U12629 (N_12629,N_12198,N_12366);
nor U12630 (N_12630,N_12163,N_12283);
or U12631 (N_12631,N_12081,N_12201);
nand U12632 (N_12632,N_12064,N_12145);
nand U12633 (N_12633,N_12092,N_12292);
nor U12634 (N_12634,N_12227,N_12335);
or U12635 (N_12635,N_12379,N_12083);
nor U12636 (N_12636,N_12394,N_12035);
nor U12637 (N_12637,N_12130,N_12307);
and U12638 (N_12638,N_12288,N_12077);
nor U12639 (N_12639,N_12348,N_12256);
xor U12640 (N_12640,N_12216,N_12288);
or U12641 (N_12641,N_12220,N_12025);
nor U12642 (N_12642,N_12032,N_12391);
nand U12643 (N_12643,N_12119,N_12242);
nor U12644 (N_12644,N_12064,N_12096);
and U12645 (N_12645,N_12096,N_12359);
xnor U12646 (N_12646,N_12051,N_12142);
xor U12647 (N_12647,N_12365,N_12025);
nor U12648 (N_12648,N_12145,N_12279);
nand U12649 (N_12649,N_12190,N_12204);
nor U12650 (N_12650,N_12318,N_12120);
nor U12651 (N_12651,N_12124,N_12092);
or U12652 (N_12652,N_12376,N_12186);
xnor U12653 (N_12653,N_12328,N_12304);
and U12654 (N_12654,N_12127,N_12399);
or U12655 (N_12655,N_12029,N_12295);
xor U12656 (N_12656,N_12364,N_12002);
xnor U12657 (N_12657,N_12095,N_12390);
nand U12658 (N_12658,N_12182,N_12257);
and U12659 (N_12659,N_12089,N_12240);
xor U12660 (N_12660,N_12083,N_12167);
and U12661 (N_12661,N_12387,N_12110);
xor U12662 (N_12662,N_12148,N_12207);
xor U12663 (N_12663,N_12343,N_12200);
nor U12664 (N_12664,N_12265,N_12006);
or U12665 (N_12665,N_12333,N_12388);
and U12666 (N_12666,N_12031,N_12338);
nand U12667 (N_12667,N_12326,N_12001);
nand U12668 (N_12668,N_12030,N_12177);
xor U12669 (N_12669,N_12229,N_12073);
nand U12670 (N_12670,N_12195,N_12391);
xor U12671 (N_12671,N_12156,N_12316);
or U12672 (N_12672,N_12113,N_12123);
xor U12673 (N_12673,N_12246,N_12377);
xor U12674 (N_12674,N_12028,N_12057);
nor U12675 (N_12675,N_12289,N_12394);
nor U12676 (N_12676,N_12184,N_12011);
or U12677 (N_12677,N_12157,N_12141);
nor U12678 (N_12678,N_12203,N_12397);
or U12679 (N_12679,N_12372,N_12196);
and U12680 (N_12680,N_12190,N_12319);
xor U12681 (N_12681,N_12338,N_12052);
and U12682 (N_12682,N_12329,N_12257);
or U12683 (N_12683,N_12317,N_12276);
nor U12684 (N_12684,N_12038,N_12337);
and U12685 (N_12685,N_12023,N_12175);
xnor U12686 (N_12686,N_12170,N_12116);
or U12687 (N_12687,N_12086,N_12314);
or U12688 (N_12688,N_12395,N_12061);
nor U12689 (N_12689,N_12247,N_12340);
xnor U12690 (N_12690,N_12222,N_12152);
xor U12691 (N_12691,N_12164,N_12042);
or U12692 (N_12692,N_12238,N_12251);
nand U12693 (N_12693,N_12163,N_12176);
nor U12694 (N_12694,N_12119,N_12264);
or U12695 (N_12695,N_12393,N_12231);
nand U12696 (N_12696,N_12010,N_12342);
xor U12697 (N_12697,N_12088,N_12244);
xor U12698 (N_12698,N_12014,N_12226);
nand U12699 (N_12699,N_12321,N_12375);
nand U12700 (N_12700,N_12029,N_12199);
and U12701 (N_12701,N_12081,N_12092);
or U12702 (N_12702,N_12101,N_12222);
nor U12703 (N_12703,N_12331,N_12096);
nor U12704 (N_12704,N_12100,N_12162);
xnor U12705 (N_12705,N_12220,N_12091);
nor U12706 (N_12706,N_12268,N_12209);
nor U12707 (N_12707,N_12093,N_12374);
nand U12708 (N_12708,N_12072,N_12280);
nor U12709 (N_12709,N_12067,N_12277);
xor U12710 (N_12710,N_12052,N_12020);
or U12711 (N_12711,N_12383,N_12289);
and U12712 (N_12712,N_12045,N_12345);
or U12713 (N_12713,N_12064,N_12362);
xor U12714 (N_12714,N_12170,N_12006);
or U12715 (N_12715,N_12227,N_12053);
or U12716 (N_12716,N_12201,N_12289);
xnor U12717 (N_12717,N_12139,N_12032);
nor U12718 (N_12718,N_12210,N_12397);
and U12719 (N_12719,N_12113,N_12051);
nor U12720 (N_12720,N_12283,N_12297);
nand U12721 (N_12721,N_12035,N_12218);
and U12722 (N_12722,N_12169,N_12142);
nand U12723 (N_12723,N_12102,N_12150);
nor U12724 (N_12724,N_12103,N_12045);
nor U12725 (N_12725,N_12014,N_12233);
xnor U12726 (N_12726,N_12093,N_12200);
and U12727 (N_12727,N_12326,N_12205);
xor U12728 (N_12728,N_12352,N_12197);
or U12729 (N_12729,N_12368,N_12107);
xor U12730 (N_12730,N_12001,N_12377);
and U12731 (N_12731,N_12371,N_12228);
nand U12732 (N_12732,N_12306,N_12059);
nand U12733 (N_12733,N_12167,N_12180);
and U12734 (N_12734,N_12256,N_12286);
nor U12735 (N_12735,N_12180,N_12099);
and U12736 (N_12736,N_12388,N_12246);
xnor U12737 (N_12737,N_12284,N_12038);
and U12738 (N_12738,N_12033,N_12017);
nand U12739 (N_12739,N_12143,N_12218);
xor U12740 (N_12740,N_12069,N_12252);
nor U12741 (N_12741,N_12205,N_12002);
nand U12742 (N_12742,N_12345,N_12087);
nor U12743 (N_12743,N_12035,N_12008);
or U12744 (N_12744,N_12239,N_12122);
nand U12745 (N_12745,N_12089,N_12079);
xnor U12746 (N_12746,N_12378,N_12246);
and U12747 (N_12747,N_12038,N_12275);
or U12748 (N_12748,N_12155,N_12173);
or U12749 (N_12749,N_12363,N_12117);
and U12750 (N_12750,N_12163,N_12133);
xor U12751 (N_12751,N_12161,N_12048);
or U12752 (N_12752,N_12060,N_12293);
and U12753 (N_12753,N_12010,N_12086);
nor U12754 (N_12754,N_12398,N_12358);
nor U12755 (N_12755,N_12380,N_12261);
and U12756 (N_12756,N_12317,N_12023);
and U12757 (N_12757,N_12020,N_12378);
xnor U12758 (N_12758,N_12337,N_12331);
nand U12759 (N_12759,N_12213,N_12211);
and U12760 (N_12760,N_12000,N_12316);
nor U12761 (N_12761,N_12012,N_12108);
xnor U12762 (N_12762,N_12157,N_12171);
or U12763 (N_12763,N_12015,N_12225);
nand U12764 (N_12764,N_12198,N_12180);
xor U12765 (N_12765,N_12259,N_12381);
nand U12766 (N_12766,N_12280,N_12170);
xor U12767 (N_12767,N_12083,N_12364);
xnor U12768 (N_12768,N_12233,N_12201);
and U12769 (N_12769,N_12208,N_12374);
nand U12770 (N_12770,N_12249,N_12125);
or U12771 (N_12771,N_12304,N_12362);
nor U12772 (N_12772,N_12288,N_12069);
nor U12773 (N_12773,N_12138,N_12273);
nand U12774 (N_12774,N_12240,N_12333);
xor U12775 (N_12775,N_12146,N_12308);
nor U12776 (N_12776,N_12185,N_12162);
nor U12777 (N_12777,N_12363,N_12304);
or U12778 (N_12778,N_12144,N_12264);
nor U12779 (N_12779,N_12140,N_12005);
nor U12780 (N_12780,N_12331,N_12387);
xnor U12781 (N_12781,N_12247,N_12170);
xnor U12782 (N_12782,N_12376,N_12185);
nand U12783 (N_12783,N_12366,N_12375);
xnor U12784 (N_12784,N_12183,N_12161);
nor U12785 (N_12785,N_12148,N_12119);
nand U12786 (N_12786,N_12361,N_12309);
nor U12787 (N_12787,N_12150,N_12155);
and U12788 (N_12788,N_12180,N_12126);
and U12789 (N_12789,N_12197,N_12025);
or U12790 (N_12790,N_12075,N_12225);
nor U12791 (N_12791,N_12003,N_12078);
nor U12792 (N_12792,N_12059,N_12234);
nand U12793 (N_12793,N_12044,N_12260);
xnor U12794 (N_12794,N_12296,N_12098);
nor U12795 (N_12795,N_12171,N_12149);
or U12796 (N_12796,N_12233,N_12319);
and U12797 (N_12797,N_12037,N_12095);
nor U12798 (N_12798,N_12375,N_12201);
nand U12799 (N_12799,N_12150,N_12305);
xor U12800 (N_12800,N_12667,N_12450);
or U12801 (N_12801,N_12702,N_12697);
nand U12802 (N_12802,N_12599,N_12563);
nor U12803 (N_12803,N_12505,N_12685);
nand U12804 (N_12804,N_12764,N_12578);
nor U12805 (N_12805,N_12757,N_12791);
nand U12806 (N_12806,N_12716,N_12596);
nand U12807 (N_12807,N_12725,N_12636);
xnor U12808 (N_12808,N_12419,N_12746);
or U12809 (N_12809,N_12477,N_12696);
or U12810 (N_12810,N_12500,N_12571);
xnor U12811 (N_12811,N_12625,N_12677);
and U12812 (N_12812,N_12695,N_12491);
or U12813 (N_12813,N_12640,N_12516);
nor U12814 (N_12814,N_12674,N_12462);
xor U12815 (N_12815,N_12736,N_12433);
or U12816 (N_12816,N_12569,N_12544);
or U12817 (N_12817,N_12490,N_12610);
and U12818 (N_12818,N_12690,N_12635);
or U12819 (N_12819,N_12469,N_12664);
xor U12820 (N_12820,N_12425,N_12644);
nand U12821 (N_12821,N_12788,N_12498);
and U12822 (N_12822,N_12503,N_12709);
nand U12823 (N_12823,N_12600,N_12799);
and U12824 (N_12824,N_12479,N_12735);
and U12825 (N_12825,N_12739,N_12564);
and U12826 (N_12826,N_12408,N_12603);
xnor U12827 (N_12827,N_12476,N_12464);
or U12828 (N_12828,N_12472,N_12779);
nor U12829 (N_12829,N_12793,N_12759);
xnor U12830 (N_12830,N_12639,N_12717);
or U12831 (N_12831,N_12649,N_12777);
nand U12832 (N_12832,N_12723,N_12642);
nor U12833 (N_12833,N_12634,N_12597);
xnor U12834 (N_12834,N_12551,N_12403);
nor U12835 (N_12835,N_12577,N_12765);
xnor U12836 (N_12836,N_12622,N_12688);
xnor U12837 (N_12837,N_12601,N_12492);
or U12838 (N_12838,N_12412,N_12556);
nor U12839 (N_12839,N_12481,N_12421);
and U12840 (N_12840,N_12595,N_12798);
nor U12841 (N_12841,N_12715,N_12430);
and U12842 (N_12842,N_12763,N_12797);
nor U12843 (N_12843,N_12771,N_12567);
xor U12844 (N_12844,N_12629,N_12658);
and U12845 (N_12845,N_12776,N_12570);
or U12846 (N_12846,N_12459,N_12553);
xnor U12847 (N_12847,N_12750,N_12444);
nand U12848 (N_12848,N_12770,N_12760);
nand U12849 (N_12849,N_12435,N_12478);
or U12850 (N_12850,N_12506,N_12766);
and U12851 (N_12851,N_12499,N_12573);
nand U12852 (N_12852,N_12698,N_12465);
nor U12853 (N_12853,N_12598,N_12730);
or U12854 (N_12854,N_12683,N_12404);
nand U12855 (N_12855,N_12582,N_12590);
or U12856 (N_12856,N_12449,N_12402);
nand U12857 (N_12857,N_12729,N_12761);
or U12858 (N_12858,N_12732,N_12415);
or U12859 (N_12859,N_12470,N_12747);
nand U12860 (N_12860,N_12485,N_12633);
nand U12861 (N_12861,N_12686,N_12645);
or U12862 (N_12862,N_12689,N_12781);
nor U12863 (N_12863,N_12726,N_12580);
nor U12864 (N_12864,N_12487,N_12699);
or U12865 (N_12865,N_12508,N_12756);
xnor U12866 (N_12866,N_12434,N_12515);
or U12867 (N_12867,N_12682,N_12539);
nand U12868 (N_12868,N_12653,N_12602);
nor U12869 (N_12869,N_12692,N_12720);
and U12870 (N_12870,N_12641,N_12537);
nor U12871 (N_12871,N_12769,N_12624);
and U12872 (N_12872,N_12438,N_12693);
nand U12873 (N_12873,N_12512,N_12703);
and U12874 (N_12874,N_12631,N_12458);
nor U12875 (N_12875,N_12733,N_12451);
or U12876 (N_12876,N_12795,N_12585);
nand U12877 (N_12877,N_12453,N_12687);
nor U12878 (N_12878,N_12426,N_12456);
or U12879 (N_12879,N_12773,N_12784);
nor U12880 (N_12880,N_12638,N_12718);
nor U12881 (N_12881,N_12783,N_12745);
xor U12882 (N_12882,N_12752,N_12486);
xor U12883 (N_12883,N_12668,N_12586);
nor U12884 (N_12884,N_12457,N_12427);
and U12885 (N_12885,N_12448,N_12753);
xor U12886 (N_12886,N_12460,N_12740);
or U12887 (N_12887,N_12681,N_12705);
xor U12888 (N_12888,N_12484,N_12751);
and U12889 (N_12889,N_12617,N_12611);
and U12890 (N_12890,N_12657,N_12443);
nand U12891 (N_12891,N_12418,N_12643);
nor U12892 (N_12892,N_12530,N_12620);
nand U12893 (N_12893,N_12767,N_12666);
or U12894 (N_12894,N_12519,N_12440);
and U12895 (N_12895,N_12768,N_12774);
nor U12896 (N_12896,N_12775,N_12615);
nor U12897 (N_12897,N_12663,N_12786);
or U12898 (N_12898,N_12475,N_12496);
nand U12899 (N_12899,N_12741,N_12561);
xnor U12900 (N_12900,N_12446,N_12670);
nor U12901 (N_12901,N_12521,N_12727);
nor U12902 (N_12902,N_12655,N_12436);
nor U12903 (N_12903,N_12424,N_12445);
xnor U12904 (N_12904,N_12704,N_12546);
xnor U12905 (N_12905,N_12742,N_12680);
xnor U12906 (N_12906,N_12559,N_12494);
nand U12907 (N_12907,N_12659,N_12731);
nand U12908 (N_12908,N_12785,N_12514);
and U12909 (N_12909,N_12708,N_12671);
xor U12910 (N_12910,N_12428,N_12592);
nand U12911 (N_12911,N_12637,N_12545);
nor U12912 (N_12912,N_12594,N_12787);
nand U12913 (N_12913,N_12557,N_12789);
and U12914 (N_12914,N_12468,N_12710);
xnor U12915 (N_12915,N_12628,N_12439);
nor U12916 (N_12916,N_12606,N_12432);
or U12917 (N_12917,N_12738,N_12414);
and U12918 (N_12918,N_12588,N_12630);
nand U12919 (N_12919,N_12714,N_12593);
nor U12920 (N_12920,N_12656,N_12591);
nand U12921 (N_12921,N_12608,N_12543);
xor U12922 (N_12922,N_12650,N_12507);
or U12923 (N_12923,N_12529,N_12581);
xor U12924 (N_12924,N_12648,N_12522);
and U12925 (N_12925,N_12417,N_12466);
or U12926 (N_12926,N_12724,N_12442);
nor U12927 (N_12927,N_12673,N_12541);
and U12928 (N_12928,N_12612,N_12712);
nand U12929 (N_12929,N_12605,N_12554);
and U12930 (N_12930,N_12755,N_12502);
xor U12931 (N_12931,N_12497,N_12647);
xnor U12932 (N_12932,N_12431,N_12662);
or U12933 (N_12933,N_12782,N_12744);
xnor U12934 (N_12934,N_12411,N_12675);
xnor U12935 (N_12935,N_12758,N_12510);
nand U12936 (N_12936,N_12558,N_12661);
xnor U12937 (N_12937,N_12748,N_12619);
xor U12938 (N_12938,N_12790,N_12616);
or U12939 (N_12939,N_12441,N_12565);
xor U12940 (N_12940,N_12583,N_12532);
nor U12941 (N_12941,N_12420,N_12413);
and U12942 (N_12942,N_12552,N_12627);
xnor U12943 (N_12943,N_12452,N_12493);
or U12944 (N_12944,N_12796,N_12646);
and U12945 (N_12945,N_12471,N_12547);
or U12946 (N_12946,N_12566,N_12778);
xor U12947 (N_12947,N_12579,N_12654);
nand U12948 (N_12948,N_12623,N_12400);
xnor U12949 (N_12949,N_12651,N_12694);
nand U12950 (N_12950,N_12762,N_12535);
and U12951 (N_12951,N_12713,N_12678);
or U12952 (N_12952,N_12527,N_12423);
and U12953 (N_12953,N_12405,N_12437);
nor U12954 (N_12954,N_12609,N_12706);
nand U12955 (N_12955,N_12589,N_12568);
xor U12956 (N_12956,N_12454,N_12792);
and U12957 (N_12957,N_12447,N_12429);
nor U12958 (N_12958,N_12401,N_12719);
xor U12959 (N_12959,N_12550,N_12734);
xnor U12960 (N_12960,N_12463,N_12542);
nand U12961 (N_12961,N_12632,N_12540);
xor U12962 (N_12962,N_12584,N_12409);
nand U12963 (N_12963,N_12495,N_12555);
and U12964 (N_12964,N_12517,N_12523);
nand U12965 (N_12965,N_12728,N_12772);
nor U12966 (N_12966,N_12669,N_12701);
and U12967 (N_12967,N_12575,N_12480);
xor U12968 (N_12968,N_12533,N_12618);
or U12969 (N_12969,N_12707,N_12672);
or U12970 (N_12970,N_12722,N_12406);
nand U12971 (N_12971,N_12474,N_12528);
or U12972 (N_12972,N_12660,N_12410);
xor U12973 (N_12973,N_12513,N_12572);
nor U12974 (N_12974,N_12562,N_12509);
xnor U12975 (N_12975,N_12538,N_12504);
and U12976 (N_12976,N_12422,N_12534);
and U12977 (N_12977,N_12501,N_12614);
xor U12978 (N_12978,N_12560,N_12576);
xor U12979 (N_12979,N_12473,N_12407);
and U12980 (N_12980,N_12461,N_12607);
nand U12981 (N_12981,N_12691,N_12754);
or U12982 (N_12982,N_12488,N_12679);
or U12983 (N_12983,N_12549,N_12520);
or U12984 (N_12984,N_12604,N_12737);
nor U12985 (N_12985,N_12743,N_12531);
xnor U12986 (N_12986,N_12511,N_12467);
and U12987 (N_12987,N_12455,N_12526);
nor U12988 (N_12988,N_12676,N_12536);
or U12989 (N_12989,N_12621,N_12524);
nand U12990 (N_12990,N_12711,N_12749);
or U12991 (N_12991,N_12518,N_12700);
or U12992 (N_12992,N_12794,N_12482);
nand U12993 (N_12993,N_12626,N_12416);
nand U12994 (N_12994,N_12780,N_12483);
and U12995 (N_12995,N_12548,N_12652);
nand U12996 (N_12996,N_12525,N_12489);
nor U12997 (N_12997,N_12587,N_12665);
or U12998 (N_12998,N_12721,N_12574);
or U12999 (N_12999,N_12684,N_12613);
and U13000 (N_13000,N_12462,N_12654);
nor U13001 (N_13001,N_12496,N_12778);
or U13002 (N_13002,N_12509,N_12664);
or U13003 (N_13003,N_12586,N_12494);
and U13004 (N_13004,N_12529,N_12561);
xor U13005 (N_13005,N_12770,N_12778);
nor U13006 (N_13006,N_12407,N_12641);
xor U13007 (N_13007,N_12506,N_12570);
nand U13008 (N_13008,N_12699,N_12519);
nor U13009 (N_13009,N_12680,N_12760);
and U13010 (N_13010,N_12665,N_12759);
and U13011 (N_13011,N_12784,N_12624);
and U13012 (N_13012,N_12484,N_12716);
xnor U13013 (N_13013,N_12623,N_12569);
xnor U13014 (N_13014,N_12788,N_12767);
xor U13015 (N_13015,N_12554,N_12665);
or U13016 (N_13016,N_12614,N_12660);
nand U13017 (N_13017,N_12438,N_12669);
nor U13018 (N_13018,N_12553,N_12676);
and U13019 (N_13019,N_12766,N_12615);
nor U13020 (N_13020,N_12713,N_12484);
xnor U13021 (N_13021,N_12664,N_12542);
nor U13022 (N_13022,N_12609,N_12683);
nor U13023 (N_13023,N_12797,N_12740);
and U13024 (N_13024,N_12446,N_12421);
and U13025 (N_13025,N_12764,N_12457);
nor U13026 (N_13026,N_12510,N_12567);
or U13027 (N_13027,N_12481,N_12473);
nor U13028 (N_13028,N_12621,N_12710);
xnor U13029 (N_13029,N_12712,N_12717);
nor U13030 (N_13030,N_12587,N_12727);
or U13031 (N_13031,N_12748,N_12731);
xor U13032 (N_13032,N_12451,N_12697);
and U13033 (N_13033,N_12551,N_12766);
nor U13034 (N_13034,N_12412,N_12499);
or U13035 (N_13035,N_12516,N_12538);
and U13036 (N_13036,N_12402,N_12505);
nor U13037 (N_13037,N_12659,N_12569);
and U13038 (N_13038,N_12770,N_12680);
nor U13039 (N_13039,N_12416,N_12749);
xnor U13040 (N_13040,N_12618,N_12768);
xor U13041 (N_13041,N_12742,N_12508);
and U13042 (N_13042,N_12704,N_12667);
or U13043 (N_13043,N_12580,N_12779);
nor U13044 (N_13044,N_12600,N_12442);
or U13045 (N_13045,N_12411,N_12694);
and U13046 (N_13046,N_12667,N_12657);
or U13047 (N_13047,N_12611,N_12690);
and U13048 (N_13048,N_12496,N_12792);
xor U13049 (N_13049,N_12417,N_12458);
or U13050 (N_13050,N_12743,N_12788);
nor U13051 (N_13051,N_12602,N_12744);
nor U13052 (N_13052,N_12724,N_12650);
xor U13053 (N_13053,N_12461,N_12706);
or U13054 (N_13054,N_12771,N_12630);
nor U13055 (N_13055,N_12723,N_12719);
and U13056 (N_13056,N_12785,N_12442);
or U13057 (N_13057,N_12586,N_12503);
or U13058 (N_13058,N_12741,N_12761);
nor U13059 (N_13059,N_12764,N_12427);
nor U13060 (N_13060,N_12717,N_12754);
nor U13061 (N_13061,N_12767,N_12750);
and U13062 (N_13062,N_12789,N_12569);
nand U13063 (N_13063,N_12516,N_12458);
and U13064 (N_13064,N_12679,N_12405);
nor U13065 (N_13065,N_12574,N_12401);
or U13066 (N_13066,N_12595,N_12755);
nor U13067 (N_13067,N_12561,N_12796);
or U13068 (N_13068,N_12758,N_12775);
or U13069 (N_13069,N_12543,N_12430);
or U13070 (N_13070,N_12624,N_12759);
nand U13071 (N_13071,N_12560,N_12704);
and U13072 (N_13072,N_12713,N_12477);
and U13073 (N_13073,N_12483,N_12543);
and U13074 (N_13074,N_12771,N_12439);
nand U13075 (N_13075,N_12620,N_12439);
and U13076 (N_13076,N_12556,N_12779);
and U13077 (N_13077,N_12685,N_12769);
or U13078 (N_13078,N_12674,N_12724);
xor U13079 (N_13079,N_12580,N_12550);
and U13080 (N_13080,N_12761,N_12411);
or U13081 (N_13081,N_12508,N_12424);
nor U13082 (N_13082,N_12436,N_12504);
and U13083 (N_13083,N_12734,N_12411);
or U13084 (N_13084,N_12681,N_12620);
xnor U13085 (N_13085,N_12436,N_12731);
nand U13086 (N_13086,N_12587,N_12481);
xnor U13087 (N_13087,N_12650,N_12412);
nor U13088 (N_13088,N_12430,N_12568);
nor U13089 (N_13089,N_12467,N_12686);
and U13090 (N_13090,N_12708,N_12575);
xor U13091 (N_13091,N_12551,N_12645);
xnor U13092 (N_13092,N_12440,N_12492);
xnor U13093 (N_13093,N_12478,N_12591);
or U13094 (N_13094,N_12538,N_12622);
xor U13095 (N_13095,N_12719,N_12500);
nor U13096 (N_13096,N_12786,N_12722);
or U13097 (N_13097,N_12563,N_12557);
nor U13098 (N_13098,N_12437,N_12760);
and U13099 (N_13099,N_12756,N_12635);
or U13100 (N_13100,N_12525,N_12540);
and U13101 (N_13101,N_12449,N_12710);
nand U13102 (N_13102,N_12441,N_12710);
xor U13103 (N_13103,N_12435,N_12776);
or U13104 (N_13104,N_12727,N_12480);
and U13105 (N_13105,N_12647,N_12487);
xnor U13106 (N_13106,N_12437,N_12415);
or U13107 (N_13107,N_12519,N_12550);
nor U13108 (N_13108,N_12731,N_12768);
nor U13109 (N_13109,N_12584,N_12678);
xor U13110 (N_13110,N_12518,N_12731);
nand U13111 (N_13111,N_12440,N_12443);
and U13112 (N_13112,N_12414,N_12742);
nor U13113 (N_13113,N_12602,N_12708);
nand U13114 (N_13114,N_12575,N_12584);
nand U13115 (N_13115,N_12686,N_12427);
or U13116 (N_13116,N_12789,N_12761);
xor U13117 (N_13117,N_12642,N_12499);
and U13118 (N_13118,N_12693,N_12793);
and U13119 (N_13119,N_12482,N_12434);
or U13120 (N_13120,N_12738,N_12629);
and U13121 (N_13121,N_12753,N_12565);
nor U13122 (N_13122,N_12455,N_12594);
and U13123 (N_13123,N_12664,N_12568);
nand U13124 (N_13124,N_12712,N_12460);
xor U13125 (N_13125,N_12779,N_12490);
nand U13126 (N_13126,N_12542,N_12722);
and U13127 (N_13127,N_12795,N_12577);
xnor U13128 (N_13128,N_12508,N_12530);
nor U13129 (N_13129,N_12472,N_12456);
xor U13130 (N_13130,N_12747,N_12477);
or U13131 (N_13131,N_12758,N_12449);
xor U13132 (N_13132,N_12536,N_12798);
and U13133 (N_13133,N_12499,N_12418);
or U13134 (N_13134,N_12532,N_12438);
xnor U13135 (N_13135,N_12432,N_12428);
xnor U13136 (N_13136,N_12543,N_12474);
nand U13137 (N_13137,N_12751,N_12709);
xor U13138 (N_13138,N_12582,N_12548);
or U13139 (N_13139,N_12410,N_12599);
or U13140 (N_13140,N_12603,N_12656);
nand U13141 (N_13141,N_12509,N_12446);
and U13142 (N_13142,N_12432,N_12457);
nand U13143 (N_13143,N_12778,N_12426);
or U13144 (N_13144,N_12646,N_12407);
or U13145 (N_13145,N_12445,N_12561);
xor U13146 (N_13146,N_12534,N_12649);
or U13147 (N_13147,N_12490,N_12680);
or U13148 (N_13148,N_12405,N_12404);
and U13149 (N_13149,N_12652,N_12471);
nand U13150 (N_13150,N_12435,N_12675);
nand U13151 (N_13151,N_12726,N_12687);
and U13152 (N_13152,N_12569,N_12663);
nand U13153 (N_13153,N_12604,N_12726);
nor U13154 (N_13154,N_12556,N_12780);
nand U13155 (N_13155,N_12457,N_12607);
and U13156 (N_13156,N_12515,N_12720);
or U13157 (N_13157,N_12787,N_12485);
nor U13158 (N_13158,N_12746,N_12522);
nand U13159 (N_13159,N_12431,N_12736);
and U13160 (N_13160,N_12785,N_12622);
xor U13161 (N_13161,N_12463,N_12722);
xnor U13162 (N_13162,N_12769,N_12676);
or U13163 (N_13163,N_12462,N_12487);
nor U13164 (N_13164,N_12717,N_12744);
or U13165 (N_13165,N_12545,N_12413);
nor U13166 (N_13166,N_12437,N_12554);
or U13167 (N_13167,N_12649,N_12767);
or U13168 (N_13168,N_12433,N_12473);
and U13169 (N_13169,N_12522,N_12482);
xor U13170 (N_13170,N_12429,N_12642);
nand U13171 (N_13171,N_12552,N_12515);
nor U13172 (N_13172,N_12565,N_12416);
or U13173 (N_13173,N_12408,N_12770);
or U13174 (N_13174,N_12600,N_12669);
or U13175 (N_13175,N_12502,N_12423);
nor U13176 (N_13176,N_12769,N_12564);
and U13177 (N_13177,N_12555,N_12704);
xnor U13178 (N_13178,N_12677,N_12531);
xor U13179 (N_13179,N_12706,N_12401);
or U13180 (N_13180,N_12472,N_12559);
xnor U13181 (N_13181,N_12796,N_12626);
and U13182 (N_13182,N_12542,N_12799);
nor U13183 (N_13183,N_12764,N_12652);
xor U13184 (N_13184,N_12423,N_12496);
nand U13185 (N_13185,N_12789,N_12540);
or U13186 (N_13186,N_12592,N_12597);
and U13187 (N_13187,N_12765,N_12750);
and U13188 (N_13188,N_12650,N_12633);
or U13189 (N_13189,N_12452,N_12614);
and U13190 (N_13190,N_12649,N_12791);
or U13191 (N_13191,N_12631,N_12401);
or U13192 (N_13192,N_12586,N_12442);
and U13193 (N_13193,N_12744,N_12682);
xnor U13194 (N_13194,N_12534,N_12413);
nand U13195 (N_13195,N_12604,N_12748);
nand U13196 (N_13196,N_12762,N_12542);
xnor U13197 (N_13197,N_12648,N_12510);
xor U13198 (N_13198,N_12764,N_12546);
nand U13199 (N_13199,N_12763,N_12703);
xor U13200 (N_13200,N_12806,N_12810);
nor U13201 (N_13201,N_12870,N_13033);
or U13202 (N_13202,N_12837,N_13061);
nand U13203 (N_13203,N_13087,N_13170);
xor U13204 (N_13204,N_13131,N_12890);
and U13205 (N_13205,N_13129,N_13139);
or U13206 (N_13206,N_12949,N_12801);
and U13207 (N_13207,N_13054,N_12873);
nand U13208 (N_13208,N_13042,N_12921);
nor U13209 (N_13209,N_13091,N_12906);
or U13210 (N_13210,N_12986,N_13010);
and U13211 (N_13211,N_13082,N_12958);
nand U13212 (N_13212,N_13050,N_13164);
xor U13213 (N_13213,N_13147,N_12970);
and U13214 (N_13214,N_12835,N_12966);
and U13215 (N_13215,N_12871,N_12972);
nor U13216 (N_13216,N_13132,N_13101);
or U13217 (N_13217,N_13074,N_12847);
nand U13218 (N_13218,N_13020,N_13017);
or U13219 (N_13219,N_12892,N_12868);
xor U13220 (N_13220,N_12975,N_13005);
xnor U13221 (N_13221,N_12998,N_12828);
xnor U13222 (N_13222,N_13071,N_13111);
or U13223 (N_13223,N_13048,N_13094);
or U13224 (N_13224,N_13148,N_13179);
nor U13225 (N_13225,N_12891,N_13055);
xnor U13226 (N_13226,N_13001,N_12991);
nand U13227 (N_13227,N_13143,N_13092);
and U13228 (N_13228,N_13014,N_13009);
and U13229 (N_13229,N_12914,N_12950);
nand U13230 (N_13230,N_13140,N_13159);
nand U13231 (N_13231,N_13052,N_13088);
xnor U13232 (N_13232,N_13122,N_12889);
xnor U13233 (N_13233,N_12814,N_12964);
and U13234 (N_13234,N_12925,N_13181);
nor U13235 (N_13235,N_12815,N_12827);
or U13236 (N_13236,N_13150,N_13135);
xnor U13237 (N_13237,N_13167,N_12875);
nor U13238 (N_13238,N_13166,N_13108);
nor U13239 (N_13239,N_13029,N_12984);
nor U13240 (N_13240,N_13188,N_13144);
nand U13241 (N_13241,N_13115,N_12956);
and U13242 (N_13242,N_12927,N_12955);
nand U13243 (N_13243,N_13025,N_13127);
or U13244 (N_13244,N_13060,N_13098);
and U13245 (N_13245,N_13165,N_12874);
or U13246 (N_13246,N_12907,N_12963);
nor U13247 (N_13247,N_12804,N_12823);
xor U13248 (N_13248,N_12940,N_13068);
and U13249 (N_13249,N_12866,N_12968);
and U13250 (N_13250,N_13110,N_12846);
nor U13251 (N_13251,N_13168,N_12820);
and U13252 (N_13252,N_13038,N_12812);
and U13253 (N_13253,N_12895,N_13109);
and U13254 (N_13254,N_13117,N_13039);
xnor U13255 (N_13255,N_13085,N_13134);
xor U13256 (N_13256,N_13174,N_12951);
and U13257 (N_13257,N_12863,N_12884);
and U13258 (N_13258,N_13193,N_12961);
nor U13259 (N_13259,N_12821,N_13194);
xor U13260 (N_13260,N_12886,N_13177);
and U13261 (N_13261,N_13057,N_12993);
nor U13262 (N_13262,N_12808,N_13128);
nand U13263 (N_13263,N_13104,N_13155);
and U13264 (N_13264,N_13173,N_13024);
or U13265 (N_13265,N_13044,N_12931);
nand U13266 (N_13266,N_13051,N_12905);
nor U13267 (N_13267,N_13083,N_12849);
or U13268 (N_13268,N_12899,N_12980);
or U13269 (N_13269,N_13078,N_12971);
nand U13270 (N_13270,N_12861,N_13099);
or U13271 (N_13271,N_13186,N_13130);
xor U13272 (N_13272,N_13192,N_13182);
nor U13273 (N_13273,N_13113,N_13016);
nand U13274 (N_13274,N_13124,N_12981);
nor U13275 (N_13275,N_12912,N_12826);
xnor U13276 (N_13276,N_12947,N_13069);
and U13277 (N_13277,N_12850,N_12976);
nor U13278 (N_13278,N_13156,N_12877);
and U13279 (N_13279,N_12953,N_12989);
and U13280 (N_13280,N_12973,N_12997);
xnor U13281 (N_13281,N_12946,N_12952);
and U13282 (N_13282,N_12830,N_13012);
xor U13283 (N_13283,N_13163,N_13106);
xor U13284 (N_13284,N_12864,N_12960);
xnor U13285 (N_13285,N_12908,N_13084);
nand U13286 (N_13286,N_12945,N_13080);
and U13287 (N_13287,N_12836,N_12813);
nor U13288 (N_13288,N_12865,N_12809);
and U13289 (N_13289,N_12932,N_13077);
nor U13290 (N_13290,N_13176,N_13089);
xor U13291 (N_13291,N_13013,N_12897);
or U13292 (N_13292,N_12974,N_12822);
xor U13293 (N_13293,N_12919,N_13197);
or U13294 (N_13294,N_12967,N_12918);
nor U13295 (N_13295,N_12954,N_13036);
or U13296 (N_13296,N_12957,N_13172);
nand U13297 (N_13297,N_13160,N_13119);
xor U13298 (N_13298,N_13035,N_12978);
xnor U13299 (N_13299,N_13162,N_12872);
xnor U13300 (N_13300,N_13000,N_13076);
and U13301 (N_13301,N_12941,N_12930);
nand U13302 (N_13302,N_13022,N_12934);
nand U13303 (N_13303,N_12883,N_13161);
xnor U13304 (N_13304,N_13026,N_13067);
or U13305 (N_13305,N_13096,N_12944);
and U13306 (N_13306,N_13027,N_13145);
nand U13307 (N_13307,N_13040,N_12840);
or U13308 (N_13308,N_13073,N_13105);
nor U13309 (N_13309,N_12922,N_12935);
or U13310 (N_13310,N_12857,N_12916);
or U13311 (N_13311,N_12988,N_12802);
nor U13312 (N_13312,N_13175,N_12985);
and U13313 (N_13313,N_12888,N_12881);
and U13314 (N_13314,N_12995,N_13072);
and U13315 (N_13315,N_12852,N_13102);
and U13316 (N_13316,N_13141,N_13075);
or U13317 (N_13317,N_12859,N_13146);
xnor U13318 (N_13318,N_13190,N_13100);
nor U13319 (N_13319,N_12844,N_12992);
nand U13320 (N_13320,N_13097,N_12856);
and U13321 (N_13321,N_13015,N_13004);
nor U13322 (N_13322,N_13183,N_13008);
xnor U13323 (N_13323,N_13199,N_13034);
nand U13324 (N_13324,N_13136,N_12851);
and U13325 (N_13325,N_13037,N_12896);
and U13326 (N_13326,N_12876,N_13196);
xnor U13327 (N_13327,N_12898,N_12869);
and U13328 (N_13328,N_12915,N_13121);
nor U13329 (N_13329,N_12816,N_13079);
or U13330 (N_13330,N_12885,N_12911);
and U13331 (N_13331,N_13154,N_13114);
or U13332 (N_13332,N_13142,N_13002);
and U13333 (N_13333,N_12839,N_13059);
xnor U13334 (N_13334,N_13032,N_12811);
xor U13335 (N_13335,N_13191,N_12878);
nor U13336 (N_13336,N_12800,N_13047);
nor U13337 (N_13337,N_12829,N_12803);
nand U13338 (N_13338,N_12969,N_12834);
xnor U13339 (N_13339,N_12903,N_12999);
or U13340 (N_13340,N_12841,N_12819);
nor U13341 (N_13341,N_13003,N_12933);
xor U13342 (N_13342,N_13066,N_12928);
nor U13343 (N_13343,N_13053,N_12858);
and U13344 (N_13344,N_13149,N_13064);
xor U13345 (N_13345,N_13151,N_13058);
nor U13346 (N_13346,N_12894,N_13063);
nand U13347 (N_13347,N_12936,N_13118);
nor U13348 (N_13348,N_13133,N_12893);
nor U13349 (N_13349,N_12962,N_12882);
xor U13350 (N_13350,N_13138,N_12862);
nand U13351 (N_13351,N_13011,N_12929);
and U13352 (N_13352,N_13116,N_12867);
nor U13353 (N_13353,N_12855,N_13049);
or U13354 (N_13354,N_13081,N_12920);
and U13355 (N_13355,N_13090,N_13045);
nor U13356 (N_13356,N_13107,N_13030);
nand U13357 (N_13357,N_13046,N_13178);
or U13358 (N_13358,N_12817,N_12818);
xnor U13359 (N_13359,N_13021,N_12979);
xor U13360 (N_13360,N_12832,N_12924);
nor U13361 (N_13361,N_12824,N_13043);
or U13362 (N_13362,N_13195,N_12994);
and U13363 (N_13363,N_12948,N_13019);
and U13364 (N_13364,N_13095,N_12848);
nor U13365 (N_13365,N_13171,N_13023);
and U13366 (N_13366,N_12942,N_13184);
xor U13367 (N_13367,N_12838,N_12880);
xnor U13368 (N_13368,N_13018,N_12825);
and U13369 (N_13369,N_13041,N_12860);
or U13370 (N_13370,N_12965,N_12990);
nand U13371 (N_13371,N_12996,N_12887);
nand U13372 (N_13372,N_12845,N_12926);
xor U13373 (N_13373,N_13185,N_12910);
or U13374 (N_13374,N_12879,N_12900);
or U13375 (N_13375,N_13158,N_12943);
nor U13376 (N_13376,N_12807,N_13086);
nand U13377 (N_13377,N_13006,N_12904);
nand U13378 (N_13378,N_13028,N_13070);
nand U13379 (N_13379,N_12831,N_12901);
nand U13380 (N_13380,N_12909,N_12805);
nand U13381 (N_13381,N_12987,N_12842);
nand U13382 (N_13382,N_13187,N_13056);
nand U13383 (N_13383,N_12923,N_13126);
nand U13384 (N_13384,N_13137,N_13157);
nor U13385 (N_13385,N_12854,N_13120);
and U13386 (N_13386,N_12853,N_13031);
nor U13387 (N_13387,N_13189,N_13065);
nor U13388 (N_13388,N_13198,N_12983);
xor U13389 (N_13389,N_13123,N_12939);
xor U13390 (N_13390,N_13152,N_13062);
xor U13391 (N_13391,N_13169,N_12917);
and U13392 (N_13392,N_12938,N_13093);
or U13393 (N_13393,N_13180,N_13125);
and U13394 (N_13394,N_12937,N_12902);
nor U13395 (N_13395,N_13112,N_12959);
nand U13396 (N_13396,N_12833,N_12843);
nand U13397 (N_13397,N_13007,N_12982);
or U13398 (N_13398,N_12913,N_12977);
nand U13399 (N_13399,N_13103,N_13153);
nand U13400 (N_13400,N_12960,N_13174);
nor U13401 (N_13401,N_13182,N_13091);
nor U13402 (N_13402,N_12956,N_13167);
xor U13403 (N_13403,N_13138,N_12896);
xnor U13404 (N_13404,N_13098,N_13108);
nor U13405 (N_13405,N_12960,N_12927);
nand U13406 (N_13406,N_12824,N_13001);
and U13407 (N_13407,N_13151,N_12876);
nand U13408 (N_13408,N_13057,N_13174);
and U13409 (N_13409,N_12967,N_12847);
xor U13410 (N_13410,N_13028,N_13043);
nor U13411 (N_13411,N_13096,N_12915);
nand U13412 (N_13412,N_13156,N_12808);
nor U13413 (N_13413,N_13025,N_12809);
and U13414 (N_13414,N_13112,N_12816);
or U13415 (N_13415,N_12974,N_12866);
and U13416 (N_13416,N_12901,N_13125);
nor U13417 (N_13417,N_13151,N_12841);
nand U13418 (N_13418,N_12821,N_12934);
or U13419 (N_13419,N_12965,N_13139);
or U13420 (N_13420,N_12914,N_12839);
and U13421 (N_13421,N_12918,N_12804);
nor U13422 (N_13422,N_12868,N_13168);
or U13423 (N_13423,N_12983,N_13044);
or U13424 (N_13424,N_12869,N_12884);
nor U13425 (N_13425,N_13141,N_12897);
nor U13426 (N_13426,N_13151,N_13159);
and U13427 (N_13427,N_13062,N_13002);
or U13428 (N_13428,N_13000,N_13120);
and U13429 (N_13429,N_12896,N_12957);
nand U13430 (N_13430,N_13025,N_13186);
and U13431 (N_13431,N_12880,N_13101);
or U13432 (N_13432,N_13079,N_12842);
nor U13433 (N_13433,N_13139,N_12876);
xor U13434 (N_13434,N_12940,N_13199);
nand U13435 (N_13435,N_13156,N_12962);
nor U13436 (N_13436,N_13033,N_13102);
or U13437 (N_13437,N_12932,N_13050);
or U13438 (N_13438,N_13134,N_12943);
and U13439 (N_13439,N_13116,N_13091);
nand U13440 (N_13440,N_12980,N_12839);
nand U13441 (N_13441,N_13067,N_13106);
or U13442 (N_13442,N_13109,N_12916);
nand U13443 (N_13443,N_13043,N_12805);
and U13444 (N_13444,N_13175,N_13153);
xnor U13445 (N_13445,N_12981,N_13144);
and U13446 (N_13446,N_13058,N_13137);
and U13447 (N_13447,N_13154,N_12920);
nand U13448 (N_13448,N_13116,N_12837);
nand U13449 (N_13449,N_13066,N_12911);
or U13450 (N_13450,N_13115,N_12866);
and U13451 (N_13451,N_12853,N_12927);
and U13452 (N_13452,N_12977,N_12988);
nor U13453 (N_13453,N_12940,N_13134);
nor U13454 (N_13454,N_12934,N_13113);
xor U13455 (N_13455,N_13195,N_13059);
xnor U13456 (N_13456,N_12869,N_13006);
nor U13457 (N_13457,N_13090,N_13191);
and U13458 (N_13458,N_12905,N_12916);
nor U13459 (N_13459,N_12931,N_13115);
nand U13460 (N_13460,N_12854,N_13075);
nand U13461 (N_13461,N_12924,N_12963);
nand U13462 (N_13462,N_13153,N_13187);
and U13463 (N_13463,N_12825,N_12966);
xnor U13464 (N_13464,N_13185,N_12959);
nor U13465 (N_13465,N_13163,N_12832);
or U13466 (N_13466,N_13060,N_13133);
nand U13467 (N_13467,N_12931,N_13060);
or U13468 (N_13468,N_12864,N_12915);
or U13469 (N_13469,N_12877,N_13197);
xor U13470 (N_13470,N_12957,N_12946);
nand U13471 (N_13471,N_12801,N_13081);
or U13472 (N_13472,N_12941,N_13132);
nand U13473 (N_13473,N_12889,N_13175);
and U13474 (N_13474,N_12859,N_12860);
xnor U13475 (N_13475,N_12850,N_13125);
and U13476 (N_13476,N_13069,N_12932);
nand U13477 (N_13477,N_13003,N_12870);
nand U13478 (N_13478,N_13140,N_13196);
xor U13479 (N_13479,N_13122,N_13132);
nor U13480 (N_13480,N_12981,N_13042);
or U13481 (N_13481,N_12920,N_13160);
nor U13482 (N_13482,N_13120,N_13109);
nand U13483 (N_13483,N_13066,N_13104);
nand U13484 (N_13484,N_13157,N_13164);
or U13485 (N_13485,N_13083,N_12856);
nand U13486 (N_13486,N_13146,N_12958);
nand U13487 (N_13487,N_13160,N_13163);
nor U13488 (N_13488,N_13182,N_12951);
nand U13489 (N_13489,N_13022,N_13077);
or U13490 (N_13490,N_12974,N_12803);
xor U13491 (N_13491,N_13157,N_12944);
and U13492 (N_13492,N_13185,N_12843);
or U13493 (N_13493,N_13132,N_13013);
nor U13494 (N_13494,N_12869,N_12814);
nand U13495 (N_13495,N_12858,N_13133);
xnor U13496 (N_13496,N_12938,N_12864);
and U13497 (N_13497,N_12988,N_12890);
xor U13498 (N_13498,N_12873,N_12911);
nand U13499 (N_13499,N_12930,N_12922);
or U13500 (N_13500,N_12837,N_12902);
xor U13501 (N_13501,N_13197,N_13073);
xor U13502 (N_13502,N_12871,N_13133);
and U13503 (N_13503,N_13173,N_13105);
and U13504 (N_13504,N_13001,N_13111);
nor U13505 (N_13505,N_13124,N_12828);
and U13506 (N_13506,N_13000,N_13134);
or U13507 (N_13507,N_12832,N_12958);
nand U13508 (N_13508,N_13183,N_12968);
or U13509 (N_13509,N_12856,N_13150);
nor U13510 (N_13510,N_12881,N_12876);
or U13511 (N_13511,N_13102,N_13084);
nor U13512 (N_13512,N_12987,N_13170);
or U13513 (N_13513,N_13040,N_12990);
nand U13514 (N_13514,N_12945,N_13138);
nand U13515 (N_13515,N_13070,N_12815);
nor U13516 (N_13516,N_13171,N_13091);
nor U13517 (N_13517,N_13091,N_12952);
nand U13518 (N_13518,N_12801,N_12825);
and U13519 (N_13519,N_13105,N_13124);
and U13520 (N_13520,N_12869,N_12961);
nor U13521 (N_13521,N_13159,N_12849);
and U13522 (N_13522,N_13075,N_13151);
or U13523 (N_13523,N_12957,N_13050);
nor U13524 (N_13524,N_13071,N_12987);
nor U13525 (N_13525,N_12810,N_12915);
or U13526 (N_13526,N_12945,N_12852);
nand U13527 (N_13527,N_12859,N_13095);
and U13528 (N_13528,N_13030,N_12992);
xor U13529 (N_13529,N_13119,N_13050);
or U13530 (N_13530,N_13072,N_12941);
nand U13531 (N_13531,N_13092,N_12939);
xnor U13532 (N_13532,N_12901,N_13129);
nor U13533 (N_13533,N_12892,N_12906);
nor U13534 (N_13534,N_12811,N_13060);
and U13535 (N_13535,N_13099,N_13059);
or U13536 (N_13536,N_13149,N_13122);
or U13537 (N_13537,N_13143,N_13170);
nand U13538 (N_13538,N_13001,N_13035);
nand U13539 (N_13539,N_13176,N_13141);
and U13540 (N_13540,N_13090,N_12919);
or U13541 (N_13541,N_13188,N_12962);
nor U13542 (N_13542,N_12870,N_13191);
nand U13543 (N_13543,N_13070,N_13005);
nand U13544 (N_13544,N_12823,N_12898);
or U13545 (N_13545,N_13189,N_13073);
or U13546 (N_13546,N_13177,N_13151);
and U13547 (N_13547,N_13031,N_12954);
xnor U13548 (N_13548,N_12946,N_13124);
and U13549 (N_13549,N_13087,N_12944);
xor U13550 (N_13550,N_12866,N_13192);
and U13551 (N_13551,N_13100,N_12844);
and U13552 (N_13552,N_12919,N_13194);
nand U13553 (N_13553,N_13138,N_13044);
nor U13554 (N_13554,N_12959,N_13037);
xnor U13555 (N_13555,N_12836,N_12932);
and U13556 (N_13556,N_13042,N_13192);
and U13557 (N_13557,N_13077,N_13070);
and U13558 (N_13558,N_12852,N_12977);
nor U13559 (N_13559,N_13067,N_12843);
or U13560 (N_13560,N_12955,N_13004);
nand U13561 (N_13561,N_12856,N_13005);
nor U13562 (N_13562,N_13143,N_12838);
and U13563 (N_13563,N_13097,N_12942);
and U13564 (N_13564,N_13167,N_12857);
nand U13565 (N_13565,N_12980,N_12809);
nand U13566 (N_13566,N_12829,N_12878);
or U13567 (N_13567,N_13083,N_12953);
or U13568 (N_13568,N_12923,N_12925);
nor U13569 (N_13569,N_12873,N_12979);
xnor U13570 (N_13570,N_12976,N_12860);
or U13571 (N_13571,N_13126,N_12924);
nor U13572 (N_13572,N_12863,N_13127);
nand U13573 (N_13573,N_12955,N_12988);
nor U13574 (N_13574,N_13146,N_12978);
xnor U13575 (N_13575,N_12824,N_12995);
nand U13576 (N_13576,N_13095,N_12837);
nand U13577 (N_13577,N_13054,N_13181);
or U13578 (N_13578,N_12865,N_13051);
and U13579 (N_13579,N_12989,N_13025);
xor U13580 (N_13580,N_12868,N_12956);
nand U13581 (N_13581,N_12892,N_13176);
nor U13582 (N_13582,N_13053,N_13026);
xor U13583 (N_13583,N_12965,N_12819);
or U13584 (N_13584,N_12960,N_13146);
or U13585 (N_13585,N_12861,N_13023);
nand U13586 (N_13586,N_12928,N_13141);
xor U13587 (N_13587,N_12951,N_13109);
nor U13588 (N_13588,N_12853,N_13040);
xor U13589 (N_13589,N_12858,N_12874);
xnor U13590 (N_13590,N_12964,N_13171);
nand U13591 (N_13591,N_13003,N_12925);
xnor U13592 (N_13592,N_13044,N_12940);
nor U13593 (N_13593,N_13156,N_13150);
nand U13594 (N_13594,N_12937,N_12847);
or U13595 (N_13595,N_12964,N_13156);
and U13596 (N_13596,N_13014,N_13029);
nand U13597 (N_13597,N_12872,N_12871);
and U13598 (N_13598,N_13036,N_12819);
xnor U13599 (N_13599,N_13176,N_13159);
nor U13600 (N_13600,N_13301,N_13352);
and U13601 (N_13601,N_13490,N_13277);
nand U13602 (N_13602,N_13365,N_13263);
and U13603 (N_13603,N_13373,N_13213);
and U13604 (N_13604,N_13564,N_13444);
nand U13605 (N_13605,N_13363,N_13331);
xor U13606 (N_13606,N_13510,N_13242);
or U13607 (N_13607,N_13558,N_13369);
or U13608 (N_13608,N_13281,N_13343);
xnor U13609 (N_13609,N_13514,N_13457);
nor U13610 (N_13610,N_13483,N_13315);
nand U13611 (N_13611,N_13561,N_13449);
or U13612 (N_13612,N_13416,N_13535);
or U13613 (N_13613,N_13505,N_13421);
and U13614 (N_13614,N_13295,N_13200);
and U13615 (N_13615,N_13446,N_13467);
or U13616 (N_13616,N_13225,N_13201);
xnor U13617 (N_13617,N_13428,N_13289);
xnor U13618 (N_13618,N_13323,N_13502);
xnor U13619 (N_13619,N_13526,N_13548);
nor U13620 (N_13620,N_13384,N_13485);
nand U13621 (N_13621,N_13357,N_13215);
xor U13622 (N_13622,N_13228,N_13403);
nand U13623 (N_13623,N_13298,N_13279);
nor U13624 (N_13624,N_13252,N_13344);
nand U13625 (N_13625,N_13224,N_13562);
nand U13626 (N_13626,N_13360,N_13304);
xnor U13627 (N_13627,N_13351,N_13453);
nor U13628 (N_13628,N_13227,N_13348);
nor U13629 (N_13629,N_13399,N_13524);
or U13630 (N_13630,N_13320,N_13405);
xnor U13631 (N_13631,N_13591,N_13381);
and U13632 (N_13632,N_13503,N_13541);
nor U13633 (N_13633,N_13547,N_13300);
nand U13634 (N_13634,N_13479,N_13390);
and U13635 (N_13635,N_13312,N_13582);
xor U13636 (N_13636,N_13486,N_13235);
nand U13637 (N_13637,N_13231,N_13572);
xnor U13638 (N_13638,N_13481,N_13529);
nor U13639 (N_13639,N_13487,N_13367);
nand U13640 (N_13640,N_13243,N_13368);
or U13641 (N_13641,N_13519,N_13478);
nand U13642 (N_13642,N_13245,N_13473);
nand U13643 (N_13643,N_13545,N_13511);
nand U13644 (N_13644,N_13212,N_13303);
and U13645 (N_13645,N_13556,N_13522);
or U13646 (N_13646,N_13376,N_13211);
nand U13647 (N_13647,N_13456,N_13570);
nor U13648 (N_13648,N_13273,N_13258);
and U13649 (N_13649,N_13538,N_13290);
or U13650 (N_13650,N_13282,N_13435);
or U13651 (N_13651,N_13397,N_13354);
xor U13652 (N_13652,N_13284,N_13317);
nand U13653 (N_13653,N_13527,N_13262);
nand U13654 (N_13654,N_13557,N_13434);
xor U13655 (N_13655,N_13571,N_13549);
nand U13656 (N_13656,N_13534,N_13313);
or U13657 (N_13657,N_13400,N_13432);
nand U13658 (N_13658,N_13402,N_13283);
nand U13659 (N_13659,N_13276,N_13546);
and U13660 (N_13660,N_13489,N_13297);
xor U13661 (N_13661,N_13240,N_13521);
xnor U13662 (N_13662,N_13496,N_13203);
nor U13663 (N_13663,N_13499,N_13458);
nand U13664 (N_13664,N_13349,N_13551);
xor U13665 (N_13665,N_13221,N_13379);
nor U13666 (N_13666,N_13305,N_13565);
or U13667 (N_13667,N_13568,N_13205);
nand U13668 (N_13668,N_13230,N_13214);
or U13669 (N_13669,N_13347,N_13267);
nor U13670 (N_13670,N_13468,N_13407);
xor U13671 (N_13671,N_13377,N_13335);
nor U13672 (N_13672,N_13555,N_13247);
xor U13673 (N_13673,N_13528,N_13234);
nand U13674 (N_13674,N_13455,N_13418);
nor U13675 (N_13675,N_13560,N_13540);
and U13676 (N_13676,N_13232,N_13274);
nor U13677 (N_13677,N_13294,N_13337);
and U13678 (N_13678,N_13575,N_13539);
nor U13679 (N_13679,N_13488,N_13382);
nand U13680 (N_13680,N_13583,N_13359);
or U13681 (N_13681,N_13553,N_13307);
or U13682 (N_13682,N_13208,N_13336);
or U13683 (N_13683,N_13469,N_13257);
and U13684 (N_13684,N_13353,N_13356);
and U13685 (N_13685,N_13306,N_13256);
and U13686 (N_13686,N_13477,N_13542);
xor U13687 (N_13687,N_13391,N_13471);
or U13688 (N_13688,N_13202,N_13419);
and U13689 (N_13689,N_13226,N_13255);
and U13690 (N_13690,N_13346,N_13248);
nor U13691 (N_13691,N_13508,N_13429);
and U13692 (N_13692,N_13392,N_13504);
and U13693 (N_13693,N_13311,N_13507);
nand U13694 (N_13694,N_13433,N_13414);
or U13695 (N_13695,N_13366,N_13345);
nor U13696 (N_13696,N_13475,N_13272);
and U13697 (N_13697,N_13461,N_13288);
or U13698 (N_13698,N_13448,N_13326);
xor U13699 (N_13699,N_13302,N_13334);
and U13700 (N_13700,N_13264,N_13525);
nor U13701 (N_13701,N_13394,N_13590);
xnor U13702 (N_13702,N_13574,N_13219);
xor U13703 (N_13703,N_13321,N_13222);
xnor U13704 (N_13704,N_13308,N_13374);
and U13705 (N_13705,N_13589,N_13513);
or U13706 (N_13706,N_13270,N_13427);
xnor U13707 (N_13707,N_13472,N_13309);
or U13708 (N_13708,N_13425,N_13569);
and U13709 (N_13709,N_13581,N_13285);
and U13710 (N_13710,N_13587,N_13410);
nor U13711 (N_13711,N_13512,N_13404);
nand U13712 (N_13712,N_13220,N_13380);
nand U13713 (N_13713,N_13566,N_13451);
or U13714 (N_13714,N_13338,N_13516);
or U13715 (N_13715,N_13375,N_13450);
xor U13716 (N_13716,N_13386,N_13577);
nand U13717 (N_13717,N_13246,N_13430);
or U13718 (N_13718,N_13415,N_13518);
or U13719 (N_13719,N_13398,N_13532);
and U13720 (N_13720,N_13426,N_13355);
and U13721 (N_13721,N_13217,N_13484);
nand U13722 (N_13722,N_13515,N_13466);
nor U13723 (N_13723,N_13586,N_13454);
and U13724 (N_13724,N_13436,N_13329);
or U13725 (N_13725,N_13445,N_13324);
nor U13726 (N_13726,N_13286,N_13580);
nor U13727 (N_13727,N_13544,N_13543);
or U13728 (N_13728,N_13494,N_13293);
xnor U13729 (N_13729,N_13480,N_13249);
xnor U13730 (N_13730,N_13576,N_13554);
nand U13731 (N_13731,N_13388,N_13501);
nor U13732 (N_13732,N_13424,N_13517);
nor U13733 (N_13733,N_13236,N_13319);
and U13734 (N_13734,N_13476,N_13462);
nand U13735 (N_13735,N_13218,N_13244);
nand U13736 (N_13736,N_13342,N_13563);
nand U13737 (N_13737,N_13389,N_13460);
and U13738 (N_13738,N_13442,N_13333);
xor U13739 (N_13739,N_13509,N_13210);
nand U13740 (N_13740,N_13420,N_13443);
nand U13741 (N_13741,N_13584,N_13408);
nor U13742 (N_13742,N_13266,N_13216);
or U13743 (N_13743,N_13598,N_13500);
or U13744 (N_13744,N_13441,N_13239);
or U13745 (N_13745,N_13371,N_13452);
and U13746 (N_13746,N_13260,N_13537);
and U13747 (N_13747,N_13250,N_13292);
xnor U13748 (N_13748,N_13209,N_13401);
nor U13749 (N_13749,N_13579,N_13271);
nand U13750 (N_13750,N_13422,N_13409);
or U13751 (N_13751,N_13387,N_13238);
nand U13752 (N_13752,N_13592,N_13383);
nand U13753 (N_13753,N_13330,N_13350);
nor U13754 (N_13754,N_13361,N_13464);
nand U13755 (N_13755,N_13296,N_13291);
or U13756 (N_13756,N_13229,N_13531);
or U13757 (N_13757,N_13411,N_13482);
or U13758 (N_13758,N_13378,N_13339);
xnor U13759 (N_13759,N_13423,N_13588);
xnor U13760 (N_13760,N_13437,N_13269);
nor U13761 (N_13761,N_13492,N_13204);
nor U13762 (N_13762,N_13497,N_13585);
nor U13763 (N_13763,N_13567,N_13395);
xor U13764 (N_13764,N_13506,N_13406);
nor U13765 (N_13765,N_13287,N_13393);
and U13766 (N_13766,N_13595,N_13596);
and U13767 (N_13767,N_13498,N_13578);
nand U13768 (N_13768,N_13533,N_13417);
or U13769 (N_13769,N_13268,N_13573);
xor U13770 (N_13770,N_13280,N_13241);
or U13771 (N_13771,N_13233,N_13207);
nand U13772 (N_13772,N_13318,N_13593);
nand U13773 (N_13773,N_13493,N_13328);
nor U13774 (N_13774,N_13316,N_13310);
nand U13775 (N_13775,N_13491,N_13474);
or U13776 (N_13776,N_13594,N_13530);
and U13777 (N_13777,N_13206,N_13520);
xor U13778 (N_13778,N_13523,N_13340);
xor U13779 (N_13779,N_13599,N_13332);
xnor U13780 (N_13780,N_13364,N_13440);
or U13781 (N_13781,N_13413,N_13495);
nand U13782 (N_13782,N_13223,N_13358);
or U13783 (N_13783,N_13261,N_13438);
and U13784 (N_13784,N_13459,N_13253);
nor U13785 (N_13785,N_13536,N_13259);
nand U13786 (N_13786,N_13559,N_13412);
nand U13787 (N_13787,N_13431,N_13275);
and U13788 (N_13788,N_13254,N_13597);
nand U13789 (N_13789,N_13327,N_13325);
xnor U13790 (N_13790,N_13552,N_13362);
nand U13791 (N_13791,N_13470,N_13251);
nor U13792 (N_13792,N_13237,N_13447);
nand U13793 (N_13793,N_13465,N_13278);
nor U13794 (N_13794,N_13299,N_13314);
nand U13795 (N_13795,N_13385,N_13439);
xnor U13796 (N_13796,N_13463,N_13341);
or U13797 (N_13797,N_13396,N_13372);
xor U13798 (N_13798,N_13265,N_13550);
nor U13799 (N_13799,N_13322,N_13370);
nand U13800 (N_13800,N_13423,N_13316);
xnor U13801 (N_13801,N_13409,N_13564);
and U13802 (N_13802,N_13390,N_13376);
xor U13803 (N_13803,N_13595,N_13266);
and U13804 (N_13804,N_13463,N_13484);
or U13805 (N_13805,N_13318,N_13208);
nor U13806 (N_13806,N_13458,N_13204);
or U13807 (N_13807,N_13273,N_13437);
and U13808 (N_13808,N_13552,N_13390);
nor U13809 (N_13809,N_13388,N_13506);
nand U13810 (N_13810,N_13211,N_13308);
nor U13811 (N_13811,N_13352,N_13304);
nand U13812 (N_13812,N_13438,N_13434);
nor U13813 (N_13813,N_13232,N_13592);
nor U13814 (N_13814,N_13494,N_13300);
xor U13815 (N_13815,N_13267,N_13566);
nor U13816 (N_13816,N_13588,N_13560);
or U13817 (N_13817,N_13481,N_13483);
nor U13818 (N_13818,N_13542,N_13520);
nand U13819 (N_13819,N_13575,N_13299);
and U13820 (N_13820,N_13449,N_13359);
nand U13821 (N_13821,N_13398,N_13478);
nor U13822 (N_13822,N_13267,N_13458);
nand U13823 (N_13823,N_13283,N_13555);
xnor U13824 (N_13824,N_13476,N_13381);
nor U13825 (N_13825,N_13430,N_13520);
nor U13826 (N_13826,N_13560,N_13462);
and U13827 (N_13827,N_13498,N_13271);
nor U13828 (N_13828,N_13531,N_13272);
and U13829 (N_13829,N_13526,N_13535);
nor U13830 (N_13830,N_13596,N_13526);
or U13831 (N_13831,N_13346,N_13391);
nand U13832 (N_13832,N_13353,N_13496);
nand U13833 (N_13833,N_13532,N_13240);
or U13834 (N_13834,N_13437,N_13511);
or U13835 (N_13835,N_13259,N_13422);
and U13836 (N_13836,N_13320,N_13264);
or U13837 (N_13837,N_13339,N_13371);
xnor U13838 (N_13838,N_13409,N_13513);
nand U13839 (N_13839,N_13284,N_13257);
xor U13840 (N_13840,N_13449,N_13553);
nor U13841 (N_13841,N_13433,N_13530);
xor U13842 (N_13842,N_13288,N_13573);
or U13843 (N_13843,N_13439,N_13445);
nor U13844 (N_13844,N_13467,N_13383);
or U13845 (N_13845,N_13209,N_13280);
or U13846 (N_13846,N_13516,N_13548);
nand U13847 (N_13847,N_13553,N_13218);
or U13848 (N_13848,N_13434,N_13282);
xnor U13849 (N_13849,N_13359,N_13263);
nand U13850 (N_13850,N_13383,N_13407);
and U13851 (N_13851,N_13331,N_13247);
nor U13852 (N_13852,N_13402,N_13307);
and U13853 (N_13853,N_13550,N_13411);
xor U13854 (N_13854,N_13377,N_13305);
or U13855 (N_13855,N_13500,N_13287);
nand U13856 (N_13856,N_13599,N_13510);
nand U13857 (N_13857,N_13576,N_13444);
or U13858 (N_13858,N_13313,N_13321);
nor U13859 (N_13859,N_13512,N_13427);
or U13860 (N_13860,N_13556,N_13364);
nor U13861 (N_13861,N_13558,N_13261);
and U13862 (N_13862,N_13550,N_13561);
and U13863 (N_13863,N_13373,N_13466);
or U13864 (N_13864,N_13386,N_13275);
or U13865 (N_13865,N_13354,N_13244);
nor U13866 (N_13866,N_13228,N_13304);
xor U13867 (N_13867,N_13354,N_13464);
nand U13868 (N_13868,N_13280,N_13363);
nor U13869 (N_13869,N_13422,N_13265);
or U13870 (N_13870,N_13204,N_13385);
nand U13871 (N_13871,N_13452,N_13416);
xnor U13872 (N_13872,N_13483,N_13593);
nand U13873 (N_13873,N_13456,N_13218);
nor U13874 (N_13874,N_13497,N_13520);
nand U13875 (N_13875,N_13212,N_13542);
or U13876 (N_13876,N_13492,N_13334);
xnor U13877 (N_13877,N_13271,N_13272);
or U13878 (N_13878,N_13543,N_13528);
and U13879 (N_13879,N_13267,N_13535);
and U13880 (N_13880,N_13401,N_13337);
xnor U13881 (N_13881,N_13331,N_13450);
and U13882 (N_13882,N_13537,N_13415);
xnor U13883 (N_13883,N_13361,N_13499);
or U13884 (N_13884,N_13430,N_13429);
nand U13885 (N_13885,N_13485,N_13241);
nor U13886 (N_13886,N_13537,N_13471);
nand U13887 (N_13887,N_13433,N_13430);
and U13888 (N_13888,N_13461,N_13593);
and U13889 (N_13889,N_13243,N_13511);
and U13890 (N_13890,N_13446,N_13255);
and U13891 (N_13891,N_13592,N_13251);
and U13892 (N_13892,N_13301,N_13223);
and U13893 (N_13893,N_13540,N_13397);
and U13894 (N_13894,N_13494,N_13219);
nand U13895 (N_13895,N_13342,N_13243);
and U13896 (N_13896,N_13211,N_13320);
or U13897 (N_13897,N_13247,N_13427);
xor U13898 (N_13898,N_13270,N_13483);
or U13899 (N_13899,N_13316,N_13517);
nand U13900 (N_13900,N_13408,N_13376);
nand U13901 (N_13901,N_13216,N_13309);
xor U13902 (N_13902,N_13423,N_13212);
xnor U13903 (N_13903,N_13341,N_13357);
xnor U13904 (N_13904,N_13288,N_13568);
xnor U13905 (N_13905,N_13222,N_13389);
and U13906 (N_13906,N_13452,N_13296);
nand U13907 (N_13907,N_13542,N_13463);
or U13908 (N_13908,N_13412,N_13439);
nand U13909 (N_13909,N_13533,N_13270);
and U13910 (N_13910,N_13421,N_13495);
nor U13911 (N_13911,N_13506,N_13579);
or U13912 (N_13912,N_13390,N_13357);
xnor U13913 (N_13913,N_13563,N_13214);
or U13914 (N_13914,N_13384,N_13253);
and U13915 (N_13915,N_13280,N_13457);
or U13916 (N_13916,N_13425,N_13353);
nand U13917 (N_13917,N_13474,N_13396);
and U13918 (N_13918,N_13288,N_13521);
xor U13919 (N_13919,N_13218,N_13344);
nand U13920 (N_13920,N_13461,N_13569);
xor U13921 (N_13921,N_13405,N_13305);
nor U13922 (N_13922,N_13367,N_13387);
nor U13923 (N_13923,N_13339,N_13247);
nor U13924 (N_13924,N_13456,N_13398);
or U13925 (N_13925,N_13310,N_13482);
and U13926 (N_13926,N_13409,N_13303);
xor U13927 (N_13927,N_13262,N_13489);
nand U13928 (N_13928,N_13335,N_13407);
or U13929 (N_13929,N_13362,N_13526);
nor U13930 (N_13930,N_13588,N_13531);
and U13931 (N_13931,N_13361,N_13444);
nor U13932 (N_13932,N_13342,N_13478);
and U13933 (N_13933,N_13406,N_13315);
xor U13934 (N_13934,N_13338,N_13245);
nand U13935 (N_13935,N_13565,N_13385);
xnor U13936 (N_13936,N_13546,N_13586);
and U13937 (N_13937,N_13433,N_13442);
xor U13938 (N_13938,N_13332,N_13382);
or U13939 (N_13939,N_13403,N_13377);
nor U13940 (N_13940,N_13237,N_13407);
or U13941 (N_13941,N_13571,N_13315);
nor U13942 (N_13942,N_13379,N_13471);
nand U13943 (N_13943,N_13299,N_13228);
or U13944 (N_13944,N_13230,N_13356);
xor U13945 (N_13945,N_13483,N_13252);
and U13946 (N_13946,N_13557,N_13382);
and U13947 (N_13947,N_13457,N_13237);
nand U13948 (N_13948,N_13486,N_13297);
or U13949 (N_13949,N_13283,N_13361);
nand U13950 (N_13950,N_13345,N_13362);
nor U13951 (N_13951,N_13326,N_13229);
or U13952 (N_13952,N_13311,N_13466);
and U13953 (N_13953,N_13281,N_13562);
nor U13954 (N_13954,N_13427,N_13447);
or U13955 (N_13955,N_13309,N_13283);
and U13956 (N_13956,N_13446,N_13511);
nor U13957 (N_13957,N_13383,N_13533);
nor U13958 (N_13958,N_13424,N_13569);
nand U13959 (N_13959,N_13231,N_13292);
nand U13960 (N_13960,N_13512,N_13467);
nand U13961 (N_13961,N_13365,N_13560);
nor U13962 (N_13962,N_13512,N_13595);
or U13963 (N_13963,N_13540,N_13519);
or U13964 (N_13964,N_13463,N_13436);
nor U13965 (N_13965,N_13368,N_13432);
or U13966 (N_13966,N_13576,N_13301);
xnor U13967 (N_13967,N_13402,N_13419);
and U13968 (N_13968,N_13486,N_13593);
nand U13969 (N_13969,N_13443,N_13590);
nand U13970 (N_13970,N_13575,N_13339);
xnor U13971 (N_13971,N_13345,N_13347);
xnor U13972 (N_13972,N_13264,N_13362);
xnor U13973 (N_13973,N_13484,N_13223);
nor U13974 (N_13974,N_13429,N_13520);
nand U13975 (N_13975,N_13413,N_13583);
xnor U13976 (N_13976,N_13212,N_13224);
nor U13977 (N_13977,N_13240,N_13540);
nor U13978 (N_13978,N_13419,N_13461);
or U13979 (N_13979,N_13298,N_13542);
xnor U13980 (N_13980,N_13429,N_13484);
nand U13981 (N_13981,N_13359,N_13355);
and U13982 (N_13982,N_13355,N_13222);
nand U13983 (N_13983,N_13246,N_13464);
and U13984 (N_13984,N_13561,N_13403);
nand U13985 (N_13985,N_13406,N_13261);
xnor U13986 (N_13986,N_13524,N_13359);
and U13987 (N_13987,N_13382,N_13575);
or U13988 (N_13988,N_13559,N_13581);
nand U13989 (N_13989,N_13293,N_13234);
nor U13990 (N_13990,N_13344,N_13469);
or U13991 (N_13991,N_13410,N_13532);
or U13992 (N_13992,N_13422,N_13464);
nor U13993 (N_13993,N_13256,N_13466);
or U13994 (N_13994,N_13420,N_13418);
or U13995 (N_13995,N_13566,N_13348);
and U13996 (N_13996,N_13454,N_13295);
and U13997 (N_13997,N_13342,N_13496);
nor U13998 (N_13998,N_13410,N_13362);
or U13999 (N_13999,N_13200,N_13310);
nor U14000 (N_14000,N_13879,N_13928);
nor U14001 (N_14001,N_13796,N_13764);
nor U14002 (N_14002,N_13685,N_13753);
or U14003 (N_14003,N_13695,N_13847);
and U14004 (N_14004,N_13667,N_13904);
or U14005 (N_14005,N_13974,N_13655);
and U14006 (N_14006,N_13773,N_13632);
nand U14007 (N_14007,N_13941,N_13801);
or U14008 (N_14008,N_13936,N_13938);
nor U14009 (N_14009,N_13827,N_13658);
xor U14010 (N_14010,N_13742,N_13991);
xnor U14011 (N_14011,N_13789,N_13835);
xor U14012 (N_14012,N_13724,N_13886);
or U14013 (N_14013,N_13869,N_13867);
nand U14014 (N_14014,N_13969,N_13907);
xnor U14015 (N_14015,N_13767,N_13730);
nand U14016 (N_14016,N_13778,N_13810);
nor U14017 (N_14017,N_13979,N_13825);
or U14018 (N_14018,N_13908,N_13903);
or U14019 (N_14019,N_13743,N_13761);
xor U14020 (N_14020,N_13814,N_13878);
and U14021 (N_14021,N_13917,N_13736);
nor U14022 (N_14022,N_13739,N_13618);
nand U14023 (N_14023,N_13838,N_13854);
nor U14024 (N_14024,N_13812,N_13627);
nor U14025 (N_14025,N_13906,N_13720);
and U14026 (N_14026,N_13981,N_13853);
or U14027 (N_14027,N_13890,N_13681);
nor U14028 (N_14028,N_13874,N_13826);
or U14029 (N_14029,N_13823,N_13640);
or U14030 (N_14030,N_13656,N_13709);
xnor U14031 (N_14031,N_13623,N_13843);
or U14032 (N_14032,N_13996,N_13792);
or U14033 (N_14033,N_13768,N_13841);
nor U14034 (N_14034,N_13716,N_13918);
nor U14035 (N_14035,N_13690,N_13740);
xnor U14036 (N_14036,N_13840,N_13619);
and U14037 (N_14037,N_13873,N_13708);
nor U14038 (N_14038,N_13975,N_13985);
and U14039 (N_14039,N_13613,N_13683);
or U14040 (N_14040,N_13808,N_13629);
nor U14041 (N_14041,N_13776,N_13661);
xor U14042 (N_14042,N_13729,N_13711);
and U14043 (N_14043,N_13758,N_13653);
nor U14044 (N_14044,N_13749,N_13967);
and U14045 (N_14045,N_13803,N_13948);
nor U14046 (N_14046,N_13602,N_13883);
nor U14047 (N_14047,N_13670,N_13726);
or U14048 (N_14048,N_13636,N_13615);
xnor U14049 (N_14049,N_13694,N_13651);
xnor U14050 (N_14050,N_13956,N_13944);
nand U14051 (N_14051,N_13872,N_13930);
or U14052 (N_14052,N_13710,N_13718);
or U14053 (N_14053,N_13631,N_13617);
nand U14054 (N_14054,N_13628,N_13824);
nor U14055 (N_14055,N_13947,N_13937);
nand U14056 (N_14056,N_13909,N_13750);
and U14057 (N_14057,N_13607,N_13786);
and U14058 (N_14058,N_13816,N_13897);
xor U14059 (N_14059,N_13833,N_13893);
and U14060 (N_14060,N_13983,N_13746);
and U14061 (N_14061,N_13677,N_13733);
nor U14062 (N_14062,N_13885,N_13963);
nor U14063 (N_14063,N_13832,N_13757);
and U14064 (N_14064,N_13714,N_13919);
or U14065 (N_14065,N_13772,N_13995);
nor U14066 (N_14066,N_13621,N_13706);
nand U14067 (N_14067,N_13807,N_13900);
and U14068 (N_14068,N_13822,N_13735);
and U14069 (N_14069,N_13756,N_13953);
nor U14070 (N_14070,N_13813,N_13682);
xor U14071 (N_14071,N_13675,N_13701);
nor U14072 (N_14072,N_13699,N_13696);
and U14073 (N_14073,N_13700,N_13986);
and U14074 (N_14074,N_13898,N_13999);
nand U14075 (N_14075,N_13732,N_13783);
nor U14076 (N_14076,N_13858,N_13647);
and U14077 (N_14077,N_13829,N_13678);
nor U14078 (N_14078,N_13751,N_13774);
nor U14079 (N_14079,N_13669,N_13952);
nand U14080 (N_14080,N_13663,N_13697);
xnor U14081 (N_14081,N_13760,N_13943);
xor U14082 (N_14082,N_13910,N_13857);
nand U14083 (N_14083,N_13950,N_13775);
xor U14084 (N_14084,N_13687,N_13608);
nand U14085 (N_14085,N_13781,N_13911);
xor U14086 (N_14086,N_13929,N_13924);
or U14087 (N_14087,N_13933,N_13649);
nor U14088 (N_14088,N_13762,N_13747);
nand U14089 (N_14089,N_13713,N_13992);
xnor U14090 (N_14090,N_13704,N_13755);
nor U14091 (N_14091,N_13959,N_13722);
xor U14092 (N_14092,N_13799,N_13795);
and U14093 (N_14093,N_13763,N_13748);
or U14094 (N_14094,N_13794,N_13844);
nand U14095 (N_14095,N_13921,N_13691);
or U14096 (N_14096,N_13728,N_13958);
and U14097 (N_14097,N_13915,N_13659);
or U14098 (N_14098,N_13849,N_13848);
nor U14099 (N_14099,N_13771,N_13644);
nor U14100 (N_14100,N_13845,N_13976);
and U14101 (N_14101,N_13856,N_13635);
xnor U14102 (N_14102,N_13988,N_13892);
or U14103 (N_14103,N_13606,N_13689);
nor U14104 (N_14104,N_13688,N_13891);
or U14105 (N_14105,N_13622,N_13980);
or U14106 (N_14106,N_13887,N_13620);
nor U14107 (N_14107,N_13693,N_13665);
or U14108 (N_14108,N_13966,N_13603);
nand U14109 (N_14109,N_13957,N_13940);
xnor U14110 (N_14110,N_13955,N_13942);
nor U14111 (N_14111,N_13637,N_13946);
or U14112 (N_14112,N_13782,N_13820);
or U14113 (N_14113,N_13962,N_13984);
or U14114 (N_14114,N_13671,N_13862);
and U14115 (N_14115,N_13790,N_13954);
and U14116 (N_14116,N_13638,N_13609);
nor U14117 (N_14117,N_13657,N_13881);
or U14118 (N_14118,N_13741,N_13960);
nand U14119 (N_14119,N_13723,N_13964);
nand U14120 (N_14120,N_13989,N_13643);
or U14121 (N_14121,N_13731,N_13779);
xnor U14122 (N_14122,N_13875,N_13806);
or U14123 (N_14123,N_13645,N_13923);
or U14124 (N_14124,N_13993,N_13777);
nand U14125 (N_14125,N_13828,N_13604);
nand U14126 (N_14126,N_13673,N_13650);
xor U14127 (N_14127,N_13895,N_13949);
or U14128 (N_14128,N_13641,N_13692);
nand U14129 (N_14129,N_13811,N_13821);
or U14130 (N_14130,N_13634,N_13601);
nor U14131 (N_14131,N_13754,N_13935);
and U14132 (N_14132,N_13668,N_13836);
xnor U14133 (N_14133,N_13932,N_13978);
and U14134 (N_14134,N_13680,N_13642);
nand U14135 (N_14135,N_13972,N_13994);
xnor U14136 (N_14136,N_13859,N_13846);
nand U14137 (N_14137,N_13961,N_13686);
or U14138 (N_14138,N_13759,N_13662);
nor U14139 (N_14139,N_13934,N_13765);
nor U14140 (N_14140,N_13676,N_13931);
nor U14141 (N_14141,N_13660,N_13672);
nand U14142 (N_14142,N_13654,N_13925);
and U14143 (N_14143,N_13815,N_13745);
xor U14144 (N_14144,N_13707,N_13600);
nand U14145 (N_14145,N_13702,N_13715);
or U14146 (N_14146,N_13861,N_13738);
xor U14147 (N_14147,N_13877,N_13834);
nor U14148 (N_14148,N_13717,N_13611);
xor U14149 (N_14149,N_13894,N_13725);
nor U14150 (N_14150,N_13666,N_13646);
nand U14151 (N_14151,N_13612,N_13837);
nor U14152 (N_14152,N_13805,N_13990);
xor U14153 (N_14153,N_13965,N_13852);
or U14154 (N_14154,N_13876,N_13850);
nand U14155 (N_14155,N_13605,N_13951);
nor U14156 (N_14156,N_13905,N_13970);
xnor U14157 (N_14157,N_13880,N_13842);
xor U14158 (N_14158,N_13896,N_13804);
or U14159 (N_14159,N_13851,N_13882);
nor U14160 (N_14160,N_13793,N_13684);
and U14161 (N_14161,N_13926,N_13787);
and U14162 (N_14162,N_13913,N_13912);
nand U14163 (N_14163,N_13791,N_13987);
or U14164 (N_14164,N_13639,N_13997);
xor U14165 (N_14165,N_13705,N_13674);
nand U14166 (N_14166,N_13625,N_13752);
and U14167 (N_14167,N_13802,N_13766);
xor U14168 (N_14168,N_13703,N_13614);
nand U14169 (N_14169,N_13977,N_13610);
or U14170 (N_14170,N_13945,N_13727);
nor U14171 (N_14171,N_13698,N_13920);
nand U14172 (N_14172,N_13721,N_13788);
or U14173 (N_14173,N_13809,N_13968);
and U14174 (N_14174,N_13616,N_13884);
nor U14175 (N_14175,N_13719,N_13899);
xnor U14176 (N_14176,N_13831,N_13902);
or U14177 (N_14177,N_13818,N_13648);
nor U14178 (N_14178,N_13652,N_13865);
and U14179 (N_14179,N_13939,N_13785);
xnor U14180 (N_14180,N_13914,N_13817);
and U14181 (N_14181,N_13630,N_13830);
or U14182 (N_14182,N_13770,N_13734);
or U14183 (N_14183,N_13922,N_13868);
nor U14184 (N_14184,N_13797,N_13819);
nor U14185 (N_14185,N_13866,N_13839);
or U14186 (N_14186,N_13780,N_13769);
and U14187 (N_14187,N_13664,N_13927);
xnor U14188 (N_14188,N_13737,N_13626);
or U14189 (N_14189,N_13870,N_13800);
and U14190 (N_14190,N_13784,N_13860);
xnor U14191 (N_14191,N_13855,N_13744);
and U14192 (N_14192,N_13982,N_13973);
and U14193 (N_14193,N_13798,N_13864);
xor U14194 (N_14194,N_13901,N_13633);
nand U14195 (N_14195,N_13871,N_13971);
nor U14196 (N_14196,N_13624,N_13712);
and U14197 (N_14197,N_13916,N_13863);
or U14198 (N_14198,N_13998,N_13679);
nand U14199 (N_14199,N_13889,N_13888);
nor U14200 (N_14200,N_13916,N_13690);
or U14201 (N_14201,N_13718,N_13659);
nand U14202 (N_14202,N_13967,N_13880);
and U14203 (N_14203,N_13891,N_13862);
nand U14204 (N_14204,N_13608,N_13712);
xnor U14205 (N_14205,N_13881,N_13717);
nand U14206 (N_14206,N_13745,N_13978);
or U14207 (N_14207,N_13745,N_13841);
nor U14208 (N_14208,N_13848,N_13992);
nand U14209 (N_14209,N_13854,N_13817);
and U14210 (N_14210,N_13873,N_13657);
nor U14211 (N_14211,N_13915,N_13808);
or U14212 (N_14212,N_13784,N_13693);
and U14213 (N_14213,N_13906,N_13841);
and U14214 (N_14214,N_13884,N_13716);
nor U14215 (N_14215,N_13750,N_13834);
nor U14216 (N_14216,N_13906,N_13898);
or U14217 (N_14217,N_13985,N_13613);
or U14218 (N_14218,N_13753,N_13769);
and U14219 (N_14219,N_13759,N_13969);
nor U14220 (N_14220,N_13867,N_13871);
nand U14221 (N_14221,N_13761,N_13847);
xnor U14222 (N_14222,N_13995,N_13979);
nand U14223 (N_14223,N_13980,N_13676);
nor U14224 (N_14224,N_13714,N_13613);
or U14225 (N_14225,N_13669,N_13977);
nand U14226 (N_14226,N_13640,N_13838);
nand U14227 (N_14227,N_13628,N_13987);
nand U14228 (N_14228,N_13712,N_13644);
or U14229 (N_14229,N_13795,N_13753);
or U14230 (N_14230,N_13614,N_13942);
xor U14231 (N_14231,N_13786,N_13853);
or U14232 (N_14232,N_13985,N_13677);
or U14233 (N_14233,N_13890,N_13702);
nand U14234 (N_14234,N_13810,N_13648);
or U14235 (N_14235,N_13995,N_13916);
and U14236 (N_14236,N_13657,N_13665);
and U14237 (N_14237,N_13985,N_13903);
or U14238 (N_14238,N_13871,N_13818);
and U14239 (N_14239,N_13604,N_13903);
or U14240 (N_14240,N_13855,N_13891);
and U14241 (N_14241,N_13833,N_13964);
or U14242 (N_14242,N_13809,N_13999);
nor U14243 (N_14243,N_13627,N_13992);
xor U14244 (N_14244,N_13953,N_13716);
and U14245 (N_14245,N_13618,N_13763);
xor U14246 (N_14246,N_13713,N_13820);
and U14247 (N_14247,N_13991,N_13936);
or U14248 (N_14248,N_13658,N_13770);
nor U14249 (N_14249,N_13797,N_13888);
or U14250 (N_14250,N_13741,N_13861);
or U14251 (N_14251,N_13637,N_13808);
or U14252 (N_14252,N_13904,N_13972);
and U14253 (N_14253,N_13917,N_13608);
xor U14254 (N_14254,N_13967,N_13930);
xor U14255 (N_14255,N_13841,N_13983);
or U14256 (N_14256,N_13600,N_13875);
nor U14257 (N_14257,N_13975,N_13644);
or U14258 (N_14258,N_13716,N_13771);
nand U14259 (N_14259,N_13828,N_13850);
xnor U14260 (N_14260,N_13869,N_13626);
nor U14261 (N_14261,N_13950,N_13747);
or U14262 (N_14262,N_13729,N_13951);
nand U14263 (N_14263,N_13863,N_13910);
and U14264 (N_14264,N_13880,N_13984);
nor U14265 (N_14265,N_13851,N_13652);
xor U14266 (N_14266,N_13949,N_13918);
nor U14267 (N_14267,N_13964,N_13620);
and U14268 (N_14268,N_13777,N_13683);
xor U14269 (N_14269,N_13964,N_13916);
xor U14270 (N_14270,N_13701,N_13654);
nand U14271 (N_14271,N_13815,N_13864);
xor U14272 (N_14272,N_13602,N_13807);
nand U14273 (N_14273,N_13619,N_13835);
xnor U14274 (N_14274,N_13810,N_13770);
or U14275 (N_14275,N_13631,N_13675);
xor U14276 (N_14276,N_13757,N_13639);
and U14277 (N_14277,N_13691,N_13724);
nor U14278 (N_14278,N_13733,N_13859);
xor U14279 (N_14279,N_13656,N_13811);
nand U14280 (N_14280,N_13894,N_13797);
nor U14281 (N_14281,N_13660,N_13663);
nand U14282 (N_14282,N_13980,N_13841);
xor U14283 (N_14283,N_13674,N_13871);
or U14284 (N_14284,N_13974,N_13953);
xnor U14285 (N_14285,N_13991,N_13790);
nand U14286 (N_14286,N_13960,N_13863);
or U14287 (N_14287,N_13742,N_13860);
or U14288 (N_14288,N_13703,N_13811);
nor U14289 (N_14289,N_13750,N_13951);
nor U14290 (N_14290,N_13735,N_13672);
nor U14291 (N_14291,N_13963,N_13938);
xnor U14292 (N_14292,N_13744,N_13705);
and U14293 (N_14293,N_13634,N_13937);
nand U14294 (N_14294,N_13805,N_13827);
and U14295 (N_14295,N_13924,N_13963);
xor U14296 (N_14296,N_13959,N_13827);
and U14297 (N_14297,N_13982,N_13672);
nand U14298 (N_14298,N_13728,N_13990);
xnor U14299 (N_14299,N_13753,N_13625);
and U14300 (N_14300,N_13883,N_13913);
nor U14301 (N_14301,N_13919,N_13901);
nand U14302 (N_14302,N_13665,N_13828);
nor U14303 (N_14303,N_13869,N_13755);
nand U14304 (N_14304,N_13993,N_13613);
nor U14305 (N_14305,N_13995,N_13721);
and U14306 (N_14306,N_13967,N_13836);
nor U14307 (N_14307,N_13668,N_13800);
and U14308 (N_14308,N_13733,N_13996);
nand U14309 (N_14309,N_13913,N_13999);
nand U14310 (N_14310,N_13796,N_13911);
or U14311 (N_14311,N_13946,N_13667);
nor U14312 (N_14312,N_13624,N_13989);
or U14313 (N_14313,N_13929,N_13832);
xnor U14314 (N_14314,N_13922,N_13802);
nor U14315 (N_14315,N_13864,N_13786);
nand U14316 (N_14316,N_13965,N_13799);
nand U14317 (N_14317,N_13847,N_13867);
nor U14318 (N_14318,N_13759,N_13624);
and U14319 (N_14319,N_13651,N_13873);
nand U14320 (N_14320,N_13655,N_13987);
xnor U14321 (N_14321,N_13747,N_13794);
nor U14322 (N_14322,N_13727,N_13817);
xor U14323 (N_14323,N_13661,N_13775);
xnor U14324 (N_14324,N_13965,N_13742);
nand U14325 (N_14325,N_13614,N_13699);
xnor U14326 (N_14326,N_13748,N_13918);
nor U14327 (N_14327,N_13841,N_13866);
xor U14328 (N_14328,N_13949,N_13615);
or U14329 (N_14329,N_13667,N_13820);
xnor U14330 (N_14330,N_13998,N_13637);
nand U14331 (N_14331,N_13627,N_13636);
xor U14332 (N_14332,N_13670,N_13839);
nand U14333 (N_14333,N_13815,N_13763);
nor U14334 (N_14334,N_13874,N_13773);
and U14335 (N_14335,N_13867,N_13854);
nor U14336 (N_14336,N_13864,N_13727);
nand U14337 (N_14337,N_13985,N_13826);
or U14338 (N_14338,N_13609,N_13613);
or U14339 (N_14339,N_13829,N_13710);
nor U14340 (N_14340,N_13642,N_13824);
nand U14341 (N_14341,N_13971,N_13710);
and U14342 (N_14342,N_13931,N_13897);
or U14343 (N_14343,N_13989,N_13913);
or U14344 (N_14344,N_13888,N_13957);
or U14345 (N_14345,N_13847,N_13698);
nor U14346 (N_14346,N_13798,N_13623);
xor U14347 (N_14347,N_13985,N_13766);
xor U14348 (N_14348,N_13857,N_13683);
and U14349 (N_14349,N_13683,N_13668);
or U14350 (N_14350,N_13907,N_13628);
or U14351 (N_14351,N_13682,N_13831);
or U14352 (N_14352,N_13911,N_13671);
or U14353 (N_14353,N_13944,N_13827);
or U14354 (N_14354,N_13654,N_13941);
nand U14355 (N_14355,N_13774,N_13837);
xnor U14356 (N_14356,N_13977,N_13702);
nand U14357 (N_14357,N_13720,N_13903);
nand U14358 (N_14358,N_13874,N_13649);
and U14359 (N_14359,N_13682,N_13641);
or U14360 (N_14360,N_13868,N_13786);
nor U14361 (N_14361,N_13697,N_13998);
or U14362 (N_14362,N_13789,N_13831);
nor U14363 (N_14363,N_13967,N_13900);
xor U14364 (N_14364,N_13808,N_13968);
or U14365 (N_14365,N_13976,N_13693);
or U14366 (N_14366,N_13795,N_13971);
nand U14367 (N_14367,N_13748,N_13646);
nor U14368 (N_14368,N_13757,N_13914);
xor U14369 (N_14369,N_13604,N_13857);
and U14370 (N_14370,N_13753,N_13881);
nor U14371 (N_14371,N_13989,N_13645);
xnor U14372 (N_14372,N_13865,N_13741);
nor U14373 (N_14373,N_13804,N_13679);
xor U14374 (N_14374,N_13621,N_13866);
nand U14375 (N_14375,N_13859,N_13887);
nand U14376 (N_14376,N_13978,N_13916);
and U14377 (N_14377,N_13838,N_13675);
nand U14378 (N_14378,N_13678,N_13671);
and U14379 (N_14379,N_13802,N_13970);
xor U14380 (N_14380,N_13940,N_13870);
nand U14381 (N_14381,N_13668,N_13745);
or U14382 (N_14382,N_13790,N_13963);
nor U14383 (N_14383,N_13815,N_13991);
xor U14384 (N_14384,N_13782,N_13700);
xnor U14385 (N_14385,N_13750,N_13747);
nand U14386 (N_14386,N_13983,N_13807);
or U14387 (N_14387,N_13999,N_13934);
nor U14388 (N_14388,N_13625,N_13864);
nor U14389 (N_14389,N_13814,N_13839);
nand U14390 (N_14390,N_13874,N_13669);
and U14391 (N_14391,N_13742,N_13975);
or U14392 (N_14392,N_13645,N_13734);
nand U14393 (N_14393,N_13650,N_13912);
nor U14394 (N_14394,N_13999,N_13942);
nand U14395 (N_14395,N_13769,N_13894);
nor U14396 (N_14396,N_13720,N_13959);
nand U14397 (N_14397,N_13708,N_13827);
nand U14398 (N_14398,N_13922,N_13783);
nor U14399 (N_14399,N_13795,N_13873);
nor U14400 (N_14400,N_14173,N_14305);
or U14401 (N_14401,N_14346,N_14073);
or U14402 (N_14402,N_14021,N_14083);
or U14403 (N_14403,N_14265,N_14300);
and U14404 (N_14404,N_14077,N_14000);
xor U14405 (N_14405,N_14210,N_14199);
or U14406 (N_14406,N_14274,N_14331);
nor U14407 (N_14407,N_14143,N_14110);
and U14408 (N_14408,N_14323,N_14111);
and U14409 (N_14409,N_14260,N_14091);
or U14410 (N_14410,N_14079,N_14024);
and U14411 (N_14411,N_14333,N_14357);
nor U14412 (N_14412,N_14159,N_14345);
or U14413 (N_14413,N_14095,N_14124);
or U14414 (N_14414,N_14360,N_14030);
xnor U14415 (N_14415,N_14202,N_14094);
nand U14416 (N_14416,N_14119,N_14087);
nand U14417 (N_14417,N_14043,N_14137);
nor U14418 (N_14418,N_14349,N_14239);
or U14419 (N_14419,N_14208,N_14232);
and U14420 (N_14420,N_14397,N_14211);
and U14421 (N_14421,N_14229,N_14179);
nand U14422 (N_14422,N_14389,N_14222);
or U14423 (N_14423,N_14193,N_14289);
nand U14424 (N_14424,N_14092,N_14186);
or U14425 (N_14425,N_14196,N_14154);
nand U14426 (N_14426,N_14285,N_14321);
nand U14427 (N_14427,N_14235,N_14054);
nand U14428 (N_14428,N_14145,N_14298);
and U14429 (N_14429,N_14053,N_14322);
xor U14430 (N_14430,N_14350,N_14135);
nor U14431 (N_14431,N_14234,N_14128);
nor U14432 (N_14432,N_14080,N_14306);
nor U14433 (N_14433,N_14342,N_14217);
and U14434 (N_14434,N_14004,N_14064);
nand U14435 (N_14435,N_14277,N_14050);
and U14436 (N_14436,N_14016,N_14393);
and U14437 (N_14437,N_14220,N_14212);
and U14438 (N_14438,N_14214,N_14266);
and U14439 (N_14439,N_14033,N_14329);
xnor U14440 (N_14440,N_14123,N_14007);
or U14441 (N_14441,N_14395,N_14187);
or U14442 (N_14442,N_14264,N_14125);
xor U14443 (N_14443,N_14276,N_14255);
nor U14444 (N_14444,N_14231,N_14078);
and U14445 (N_14445,N_14134,N_14197);
xor U14446 (N_14446,N_14215,N_14182);
or U14447 (N_14447,N_14028,N_14038);
nand U14448 (N_14448,N_14047,N_14074);
xnor U14449 (N_14449,N_14097,N_14251);
nor U14450 (N_14450,N_14181,N_14177);
or U14451 (N_14451,N_14262,N_14241);
xnor U14452 (N_14452,N_14219,N_14148);
nor U14453 (N_14453,N_14081,N_14103);
and U14454 (N_14454,N_14273,N_14390);
nand U14455 (N_14455,N_14367,N_14358);
nor U14456 (N_14456,N_14191,N_14108);
xnor U14457 (N_14457,N_14045,N_14051);
nor U14458 (N_14458,N_14006,N_14216);
nand U14459 (N_14459,N_14157,N_14308);
xnor U14460 (N_14460,N_14353,N_14138);
xor U14461 (N_14461,N_14250,N_14375);
xor U14462 (N_14462,N_14020,N_14259);
xor U14463 (N_14463,N_14242,N_14207);
and U14464 (N_14464,N_14105,N_14025);
xnor U14465 (N_14465,N_14213,N_14198);
xor U14466 (N_14466,N_14291,N_14171);
nand U14467 (N_14467,N_14385,N_14324);
nand U14468 (N_14468,N_14106,N_14023);
nor U14469 (N_14469,N_14090,N_14076);
xor U14470 (N_14470,N_14374,N_14351);
and U14471 (N_14471,N_14066,N_14046);
or U14472 (N_14472,N_14283,N_14263);
nor U14473 (N_14473,N_14354,N_14115);
xor U14474 (N_14474,N_14098,N_14101);
and U14475 (N_14475,N_14109,N_14335);
and U14476 (N_14476,N_14174,N_14227);
nor U14477 (N_14477,N_14003,N_14086);
nor U14478 (N_14478,N_14142,N_14280);
xnor U14479 (N_14479,N_14317,N_14188);
xor U14480 (N_14480,N_14194,N_14352);
or U14481 (N_14481,N_14133,N_14027);
xor U14482 (N_14482,N_14205,N_14200);
and U14483 (N_14483,N_14127,N_14293);
and U14484 (N_14484,N_14243,N_14132);
xnor U14485 (N_14485,N_14032,N_14309);
nor U14486 (N_14486,N_14096,N_14061);
or U14487 (N_14487,N_14052,N_14175);
and U14488 (N_14488,N_14294,N_14152);
nand U14489 (N_14489,N_14368,N_14141);
xnor U14490 (N_14490,N_14223,N_14019);
nor U14491 (N_14491,N_14249,N_14112);
nor U14492 (N_14492,N_14018,N_14378);
and U14493 (N_14493,N_14268,N_14359);
xnor U14494 (N_14494,N_14383,N_14151);
or U14495 (N_14495,N_14048,N_14224);
and U14496 (N_14496,N_14129,N_14203);
or U14497 (N_14497,N_14169,N_14258);
xnor U14498 (N_14498,N_14165,N_14313);
or U14499 (N_14499,N_14069,N_14085);
nor U14500 (N_14500,N_14218,N_14099);
and U14501 (N_14501,N_14271,N_14036);
and U14502 (N_14502,N_14136,N_14072);
or U14503 (N_14503,N_14278,N_14238);
or U14504 (N_14504,N_14387,N_14185);
and U14505 (N_14505,N_14270,N_14286);
nor U14506 (N_14506,N_14225,N_14284);
and U14507 (N_14507,N_14149,N_14183);
xnor U14508 (N_14508,N_14247,N_14155);
nand U14509 (N_14509,N_14176,N_14147);
nand U14510 (N_14510,N_14384,N_14049);
xnor U14511 (N_14511,N_14131,N_14337);
and U14512 (N_14512,N_14369,N_14319);
nor U14513 (N_14513,N_14257,N_14120);
nor U14514 (N_14514,N_14022,N_14339);
nand U14515 (N_14515,N_14236,N_14261);
nor U14516 (N_14516,N_14332,N_14288);
or U14517 (N_14517,N_14279,N_14292);
xnor U14518 (N_14518,N_14275,N_14068);
and U14519 (N_14519,N_14381,N_14035);
nor U14520 (N_14520,N_14282,N_14190);
and U14521 (N_14521,N_14362,N_14221);
xnor U14522 (N_14522,N_14060,N_14160);
and U14523 (N_14523,N_14348,N_14310);
nand U14524 (N_14524,N_14002,N_14399);
nor U14525 (N_14525,N_14082,N_14189);
nor U14526 (N_14526,N_14037,N_14156);
xor U14527 (N_14527,N_14245,N_14386);
or U14528 (N_14528,N_14314,N_14327);
or U14529 (N_14529,N_14014,N_14067);
nand U14530 (N_14530,N_14391,N_14167);
and U14531 (N_14531,N_14272,N_14040);
nand U14532 (N_14532,N_14341,N_14012);
and U14533 (N_14533,N_14244,N_14114);
or U14534 (N_14534,N_14304,N_14011);
and U14535 (N_14535,N_14372,N_14166);
nor U14536 (N_14536,N_14065,N_14376);
nand U14537 (N_14537,N_14059,N_14015);
or U14538 (N_14538,N_14008,N_14281);
and U14539 (N_14539,N_14315,N_14010);
or U14540 (N_14540,N_14195,N_14330);
nor U14541 (N_14541,N_14034,N_14139);
nor U14542 (N_14542,N_14340,N_14347);
nand U14543 (N_14543,N_14117,N_14233);
or U14544 (N_14544,N_14325,N_14089);
nand U14545 (N_14545,N_14240,N_14209);
or U14546 (N_14546,N_14102,N_14093);
or U14547 (N_14547,N_14248,N_14297);
nor U14548 (N_14548,N_14246,N_14084);
or U14549 (N_14549,N_14355,N_14170);
nor U14550 (N_14550,N_14204,N_14328);
nand U14551 (N_14551,N_14062,N_14026);
or U14552 (N_14552,N_14031,N_14017);
or U14553 (N_14553,N_14302,N_14338);
or U14554 (N_14554,N_14107,N_14075);
nor U14555 (N_14555,N_14256,N_14146);
xor U14556 (N_14556,N_14320,N_14013);
nor U14557 (N_14557,N_14254,N_14039);
and U14558 (N_14558,N_14334,N_14370);
xor U14559 (N_14559,N_14164,N_14162);
and U14560 (N_14560,N_14088,N_14377);
and U14561 (N_14561,N_14122,N_14230);
xnor U14562 (N_14562,N_14005,N_14373);
and U14563 (N_14563,N_14344,N_14253);
nor U14564 (N_14564,N_14366,N_14336);
xor U14565 (N_14565,N_14295,N_14252);
xnor U14566 (N_14566,N_14158,N_14057);
xnor U14567 (N_14567,N_14144,N_14121);
nand U14568 (N_14568,N_14290,N_14056);
nand U14569 (N_14569,N_14379,N_14226);
nor U14570 (N_14570,N_14178,N_14237);
nor U14571 (N_14571,N_14299,N_14041);
or U14572 (N_14572,N_14206,N_14058);
xnor U14573 (N_14573,N_14365,N_14269);
xnor U14574 (N_14574,N_14100,N_14398);
and U14575 (N_14575,N_14318,N_14163);
xnor U14576 (N_14576,N_14356,N_14361);
nor U14577 (N_14577,N_14396,N_14161);
or U14578 (N_14578,N_14392,N_14130);
nor U14579 (N_14579,N_14104,N_14388);
nand U14580 (N_14580,N_14150,N_14042);
xnor U14581 (N_14581,N_14070,N_14180);
and U14582 (N_14582,N_14380,N_14055);
and U14583 (N_14583,N_14316,N_14126);
nor U14584 (N_14584,N_14063,N_14168);
xor U14585 (N_14585,N_14296,N_14071);
nor U14586 (N_14586,N_14029,N_14364);
and U14587 (N_14587,N_14153,N_14192);
or U14588 (N_14588,N_14113,N_14140);
xnor U14589 (N_14589,N_14228,N_14044);
and U14590 (N_14590,N_14311,N_14307);
and U14591 (N_14591,N_14312,N_14301);
nor U14592 (N_14592,N_14303,N_14267);
nand U14593 (N_14593,N_14394,N_14116);
or U14594 (N_14594,N_14343,N_14118);
nand U14595 (N_14595,N_14001,N_14382);
and U14596 (N_14596,N_14184,N_14363);
nor U14597 (N_14597,N_14326,N_14287);
nand U14598 (N_14598,N_14009,N_14172);
xnor U14599 (N_14599,N_14371,N_14201);
nand U14600 (N_14600,N_14342,N_14220);
or U14601 (N_14601,N_14190,N_14301);
xnor U14602 (N_14602,N_14230,N_14150);
nand U14603 (N_14603,N_14166,N_14197);
nor U14604 (N_14604,N_14363,N_14046);
nor U14605 (N_14605,N_14081,N_14337);
or U14606 (N_14606,N_14222,N_14058);
nor U14607 (N_14607,N_14296,N_14153);
nor U14608 (N_14608,N_14032,N_14329);
and U14609 (N_14609,N_14224,N_14150);
nor U14610 (N_14610,N_14121,N_14385);
and U14611 (N_14611,N_14155,N_14006);
or U14612 (N_14612,N_14102,N_14110);
and U14613 (N_14613,N_14192,N_14201);
nand U14614 (N_14614,N_14044,N_14187);
nand U14615 (N_14615,N_14327,N_14239);
nor U14616 (N_14616,N_14336,N_14204);
and U14617 (N_14617,N_14083,N_14048);
nand U14618 (N_14618,N_14256,N_14116);
nor U14619 (N_14619,N_14307,N_14304);
or U14620 (N_14620,N_14206,N_14146);
or U14621 (N_14621,N_14240,N_14237);
xnor U14622 (N_14622,N_14348,N_14312);
and U14623 (N_14623,N_14096,N_14113);
or U14624 (N_14624,N_14106,N_14366);
xor U14625 (N_14625,N_14119,N_14239);
nand U14626 (N_14626,N_14123,N_14301);
xor U14627 (N_14627,N_14382,N_14123);
and U14628 (N_14628,N_14321,N_14001);
nor U14629 (N_14629,N_14339,N_14147);
nor U14630 (N_14630,N_14377,N_14293);
nor U14631 (N_14631,N_14021,N_14379);
and U14632 (N_14632,N_14151,N_14017);
xnor U14633 (N_14633,N_14389,N_14065);
nand U14634 (N_14634,N_14374,N_14143);
nor U14635 (N_14635,N_14331,N_14352);
or U14636 (N_14636,N_14283,N_14171);
nor U14637 (N_14637,N_14315,N_14061);
and U14638 (N_14638,N_14331,N_14198);
and U14639 (N_14639,N_14262,N_14377);
nand U14640 (N_14640,N_14246,N_14234);
xnor U14641 (N_14641,N_14258,N_14298);
xor U14642 (N_14642,N_14025,N_14198);
xor U14643 (N_14643,N_14239,N_14183);
or U14644 (N_14644,N_14129,N_14187);
or U14645 (N_14645,N_14169,N_14251);
xnor U14646 (N_14646,N_14012,N_14006);
nand U14647 (N_14647,N_14358,N_14228);
nor U14648 (N_14648,N_14375,N_14088);
nand U14649 (N_14649,N_14284,N_14167);
and U14650 (N_14650,N_14218,N_14359);
nor U14651 (N_14651,N_14166,N_14144);
nand U14652 (N_14652,N_14327,N_14283);
xor U14653 (N_14653,N_14008,N_14276);
xor U14654 (N_14654,N_14300,N_14237);
or U14655 (N_14655,N_14165,N_14251);
xor U14656 (N_14656,N_14189,N_14227);
nor U14657 (N_14657,N_14102,N_14127);
xor U14658 (N_14658,N_14077,N_14139);
nor U14659 (N_14659,N_14302,N_14153);
xnor U14660 (N_14660,N_14213,N_14287);
or U14661 (N_14661,N_14076,N_14061);
xor U14662 (N_14662,N_14343,N_14312);
xor U14663 (N_14663,N_14191,N_14186);
nand U14664 (N_14664,N_14002,N_14181);
and U14665 (N_14665,N_14109,N_14398);
and U14666 (N_14666,N_14342,N_14347);
and U14667 (N_14667,N_14274,N_14368);
nand U14668 (N_14668,N_14107,N_14364);
and U14669 (N_14669,N_14153,N_14228);
or U14670 (N_14670,N_14030,N_14229);
xnor U14671 (N_14671,N_14266,N_14324);
nand U14672 (N_14672,N_14173,N_14395);
and U14673 (N_14673,N_14040,N_14318);
nand U14674 (N_14674,N_14321,N_14044);
nand U14675 (N_14675,N_14047,N_14304);
or U14676 (N_14676,N_14068,N_14296);
nor U14677 (N_14677,N_14157,N_14298);
nand U14678 (N_14678,N_14134,N_14265);
and U14679 (N_14679,N_14173,N_14276);
nor U14680 (N_14680,N_14008,N_14372);
or U14681 (N_14681,N_14047,N_14184);
nor U14682 (N_14682,N_14095,N_14104);
nor U14683 (N_14683,N_14129,N_14375);
xnor U14684 (N_14684,N_14333,N_14396);
and U14685 (N_14685,N_14133,N_14237);
and U14686 (N_14686,N_14375,N_14107);
xor U14687 (N_14687,N_14178,N_14261);
xor U14688 (N_14688,N_14124,N_14148);
nor U14689 (N_14689,N_14128,N_14360);
nand U14690 (N_14690,N_14225,N_14158);
or U14691 (N_14691,N_14055,N_14114);
nor U14692 (N_14692,N_14265,N_14282);
xnor U14693 (N_14693,N_14154,N_14078);
nand U14694 (N_14694,N_14164,N_14222);
or U14695 (N_14695,N_14398,N_14337);
and U14696 (N_14696,N_14019,N_14078);
nor U14697 (N_14697,N_14100,N_14027);
nor U14698 (N_14698,N_14258,N_14237);
and U14699 (N_14699,N_14231,N_14009);
nand U14700 (N_14700,N_14333,N_14275);
or U14701 (N_14701,N_14320,N_14374);
nand U14702 (N_14702,N_14149,N_14186);
nor U14703 (N_14703,N_14136,N_14152);
nand U14704 (N_14704,N_14391,N_14227);
nand U14705 (N_14705,N_14288,N_14041);
xor U14706 (N_14706,N_14168,N_14125);
or U14707 (N_14707,N_14370,N_14247);
xnor U14708 (N_14708,N_14162,N_14080);
or U14709 (N_14709,N_14221,N_14182);
and U14710 (N_14710,N_14102,N_14099);
or U14711 (N_14711,N_14183,N_14271);
or U14712 (N_14712,N_14012,N_14071);
xnor U14713 (N_14713,N_14176,N_14222);
nand U14714 (N_14714,N_14217,N_14128);
and U14715 (N_14715,N_14379,N_14246);
or U14716 (N_14716,N_14114,N_14293);
xor U14717 (N_14717,N_14232,N_14300);
and U14718 (N_14718,N_14249,N_14002);
xnor U14719 (N_14719,N_14006,N_14231);
or U14720 (N_14720,N_14144,N_14058);
and U14721 (N_14721,N_14073,N_14107);
and U14722 (N_14722,N_14223,N_14119);
nor U14723 (N_14723,N_14076,N_14309);
nand U14724 (N_14724,N_14077,N_14003);
or U14725 (N_14725,N_14302,N_14267);
xor U14726 (N_14726,N_14202,N_14174);
nand U14727 (N_14727,N_14357,N_14241);
and U14728 (N_14728,N_14036,N_14269);
xnor U14729 (N_14729,N_14274,N_14298);
xor U14730 (N_14730,N_14208,N_14223);
or U14731 (N_14731,N_14263,N_14057);
nand U14732 (N_14732,N_14303,N_14004);
and U14733 (N_14733,N_14087,N_14076);
or U14734 (N_14734,N_14241,N_14028);
and U14735 (N_14735,N_14374,N_14296);
xor U14736 (N_14736,N_14148,N_14217);
xnor U14737 (N_14737,N_14231,N_14346);
and U14738 (N_14738,N_14306,N_14348);
or U14739 (N_14739,N_14238,N_14101);
and U14740 (N_14740,N_14307,N_14156);
nor U14741 (N_14741,N_14004,N_14197);
or U14742 (N_14742,N_14246,N_14007);
or U14743 (N_14743,N_14196,N_14179);
and U14744 (N_14744,N_14355,N_14393);
nor U14745 (N_14745,N_14352,N_14229);
or U14746 (N_14746,N_14047,N_14022);
and U14747 (N_14747,N_14266,N_14254);
and U14748 (N_14748,N_14316,N_14179);
nor U14749 (N_14749,N_14268,N_14357);
or U14750 (N_14750,N_14068,N_14021);
nor U14751 (N_14751,N_14340,N_14258);
nand U14752 (N_14752,N_14381,N_14265);
or U14753 (N_14753,N_14324,N_14274);
or U14754 (N_14754,N_14204,N_14348);
or U14755 (N_14755,N_14003,N_14187);
and U14756 (N_14756,N_14252,N_14064);
and U14757 (N_14757,N_14202,N_14097);
nand U14758 (N_14758,N_14086,N_14099);
xor U14759 (N_14759,N_14322,N_14371);
xor U14760 (N_14760,N_14091,N_14067);
nand U14761 (N_14761,N_14252,N_14309);
nand U14762 (N_14762,N_14178,N_14164);
and U14763 (N_14763,N_14101,N_14341);
and U14764 (N_14764,N_14331,N_14046);
nor U14765 (N_14765,N_14152,N_14322);
or U14766 (N_14766,N_14074,N_14084);
xnor U14767 (N_14767,N_14356,N_14261);
nor U14768 (N_14768,N_14001,N_14285);
and U14769 (N_14769,N_14060,N_14283);
xnor U14770 (N_14770,N_14088,N_14197);
and U14771 (N_14771,N_14395,N_14332);
and U14772 (N_14772,N_14043,N_14307);
or U14773 (N_14773,N_14241,N_14233);
and U14774 (N_14774,N_14282,N_14124);
and U14775 (N_14775,N_14101,N_14061);
and U14776 (N_14776,N_14012,N_14068);
nor U14777 (N_14777,N_14241,N_14378);
or U14778 (N_14778,N_14278,N_14313);
xnor U14779 (N_14779,N_14383,N_14048);
nor U14780 (N_14780,N_14263,N_14153);
xnor U14781 (N_14781,N_14135,N_14299);
nand U14782 (N_14782,N_14208,N_14310);
nand U14783 (N_14783,N_14286,N_14070);
xnor U14784 (N_14784,N_14050,N_14069);
and U14785 (N_14785,N_14376,N_14181);
and U14786 (N_14786,N_14321,N_14046);
xor U14787 (N_14787,N_14146,N_14208);
nor U14788 (N_14788,N_14085,N_14217);
or U14789 (N_14789,N_14188,N_14099);
or U14790 (N_14790,N_14176,N_14291);
and U14791 (N_14791,N_14103,N_14358);
nand U14792 (N_14792,N_14125,N_14048);
nor U14793 (N_14793,N_14099,N_14126);
nor U14794 (N_14794,N_14131,N_14019);
xnor U14795 (N_14795,N_14380,N_14300);
xor U14796 (N_14796,N_14226,N_14370);
nor U14797 (N_14797,N_14340,N_14285);
xnor U14798 (N_14798,N_14098,N_14294);
xnor U14799 (N_14799,N_14046,N_14308);
nand U14800 (N_14800,N_14512,N_14523);
nand U14801 (N_14801,N_14679,N_14508);
nand U14802 (N_14802,N_14715,N_14592);
and U14803 (N_14803,N_14431,N_14422);
nor U14804 (N_14804,N_14607,N_14582);
and U14805 (N_14805,N_14759,N_14664);
nand U14806 (N_14806,N_14553,N_14434);
or U14807 (N_14807,N_14792,N_14410);
and U14808 (N_14808,N_14625,N_14758);
and U14809 (N_14809,N_14565,N_14726);
nor U14810 (N_14810,N_14764,N_14620);
nand U14811 (N_14811,N_14490,N_14540);
or U14812 (N_14812,N_14420,N_14665);
and U14813 (N_14813,N_14405,N_14750);
nand U14814 (N_14814,N_14517,N_14707);
nand U14815 (N_14815,N_14690,N_14411);
or U14816 (N_14816,N_14534,N_14652);
xnor U14817 (N_14817,N_14748,N_14419);
nor U14818 (N_14818,N_14643,N_14735);
nor U14819 (N_14819,N_14404,N_14587);
nor U14820 (N_14820,N_14407,N_14791);
xnor U14821 (N_14821,N_14755,N_14595);
nor U14822 (N_14822,N_14589,N_14779);
or U14823 (N_14823,N_14599,N_14549);
and U14824 (N_14824,N_14501,N_14509);
or U14825 (N_14825,N_14653,N_14436);
xor U14826 (N_14826,N_14738,N_14452);
or U14827 (N_14827,N_14714,N_14711);
and U14828 (N_14828,N_14686,N_14684);
and U14829 (N_14829,N_14602,N_14533);
and U14830 (N_14830,N_14784,N_14539);
and U14831 (N_14831,N_14639,N_14729);
nor U14832 (N_14832,N_14586,N_14634);
xor U14833 (N_14833,N_14421,N_14633);
and U14834 (N_14834,N_14526,N_14521);
xor U14835 (N_14835,N_14756,N_14669);
nand U14836 (N_14836,N_14547,N_14524);
nand U14837 (N_14837,N_14573,N_14427);
nand U14838 (N_14838,N_14737,N_14594);
nor U14839 (N_14839,N_14515,N_14687);
or U14840 (N_14840,N_14782,N_14655);
nor U14841 (N_14841,N_14778,N_14767);
nand U14842 (N_14842,N_14498,N_14483);
nor U14843 (N_14843,N_14464,N_14462);
or U14844 (N_14844,N_14439,N_14603);
nor U14845 (N_14845,N_14775,N_14499);
or U14846 (N_14846,N_14604,N_14799);
nor U14847 (N_14847,N_14794,N_14771);
nor U14848 (N_14848,N_14641,N_14768);
and U14849 (N_14849,N_14471,N_14752);
nand U14850 (N_14850,N_14670,N_14456);
or U14851 (N_14851,N_14511,N_14660);
nand U14852 (N_14852,N_14504,N_14678);
or U14853 (N_14853,N_14642,N_14481);
nor U14854 (N_14854,N_14469,N_14635);
nor U14855 (N_14855,N_14701,N_14712);
or U14856 (N_14856,N_14721,N_14455);
nand U14857 (N_14857,N_14688,N_14785);
nor U14858 (N_14858,N_14566,N_14583);
or U14859 (N_14859,N_14488,N_14424);
nor U14860 (N_14860,N_14437,N_14507);
nand U14861 (N_14861,N_14662,N_14644);
nand U14862 (N_14862,N_14415,N_14522);
nor U14863 (N_14863,N_14659,N_14530);
nand U14864 (N_14864,N_14645,N_14581);
and U14865 (N_14865,N_14786,N_14449);
or U14866 (N_14866,N_14579,N_14555);
nand U14867 (N_14867,N_14485,N_14535);
nor U14868 (N_14868,N_14689,N_14740);
xnor U14869 (N_14869,N_14441,N_14454);
and U14870 (N_14870,N_14776,N_14495);
nand U14871 (N_14871,N_14596,N_14716);
and U14872 (N_14872,N_14629,N_14502);
and U14873 (N_14873,N_14546,N_14683);
xnor U14874 (N_14874,N_14733,N_14751);
or U14875 (N_14875,N_14700,N_14626);
nand U14876 (N_14876,N_14409,N_14691);
nor U14877 (N_14877,N_14706,N_14438);
nor U14878 (N_14878,N_14465,N_14487);
nor U14879 (N_14879,N_14703,N_14637);
nand U14880 (N_14880,N_14484,N_14468);
nor U14881 (N_14881,N_14693,N_14646);
nand U14882 (N_14882,N_14492,N_14731);
or U14883 (N_14883,N_14558,N_14567);
xor U14884 (N_14884,N_14519,N_14681);
and U14885 (N_14885,N_14463,N_14741);
xnor U14886 (N_14886,N_14542,N_14494);
and U14887 (N_14887,N_14467,N_14704);
xor U14888 (N_14888,N_14656,N_14457);
or U14889 (N_14889,N_14575,N_14561);
xor U14890 (N_14890,N_14450,N_14673);
nor U14891 (N_14891,N_14429,N_14552);
and U14892 (N_14892,N_14408,N_14401);
nor U14893 (N_14893,N_14772,N_14798);
nand U14894 (N_14894,N_14417,N_14598);
nand U14895 (N_14895,N_14541,N_14766);
or U14896 (N_14896,N_14649,N_14717);
nand U14897 (N_14897,N_14459,N_14537);
nor U14898 (N_14898,N_14577,N_14616);
nand U14899 (N_14899,N_14777,N_14479);
nand U14900 (N_14900,N_14482,N_14562);
or U14901 (N_14901,N_14632,N_14458);
nand U14902 (N_14902,N_14525,N_14654);
nor U14903 (N_14903,N_14722,N_14491);
or U14904 (N_14904,N_14710,N_14762);
or U14905 (N_14905,N_14430,N_14796);
nor U14906 (N_14906,N_14753,N_14739);
nand U14907 (N_14907,N_14795,N_14723);
nand U14908 (N_14908,N_14453,N_14569);
or U14909 (N_14909,N_14708,N_14412);
and U14910 (N_14910,N_14667,N_14601);
nand U14911 (N_14911,N_14568,N_14694);
and U14912 (N_14912,N_14647,N_14727);
nor U14913 (N_14913,N_14557,N_14418);
nor U14914 (N_14914,N_14531,N_14783);
nand U14915 (N_14915,N_14497,N_14496);
nor U14916 (N_14916,N_14680,N_14769);
xnor U14917 (N_14917,N_14675,N_14773);
and U14918 (N_14918,N_14651,N_14605);
nand U14919 (N_14919,N_14608,N_14702);
xnor U14920 (N_14920,N_14763,N_14527);
or U14921 (N_14921,N_14745,N_14445);
or U14922 (N_14922,N_14610,N_14513);
nand U14923 (N_14923,N_14663,N_14460);
or U14924 (N_14924,N_14584,N_14674);
nand U14925 (N_14925,N_14551,N_14671);
nand U14926 (N_14926,N_14480,N_14719);
and U14927 (N_14927,N_14624,N_14413);
xor U14928 (N_14928,N_14543,N_14698);
and U14929 (N_14929,N_14559,N_14746);
and U14930 (N_14930,N_14423,N_14477);
or U14931 (N_14931,N_14406,N_14563);
and U14932 (N_14932,N_14685,N_14600);
nor U14933 (N_14933,N_14630,N_14609);
nor U14934 (N_14934,N_14736,N_14442);
nor U14935 (N_14935,N_14742,N_14443);
xnor U14936 (N_14936,N_14780,N_14532);
nor U14937 (N_14937,N_14754,N_14590);
nand U14938 (N_14938,N_14572,N_14725);
and U14939 (N_14939,N_14612,N_14451);
or U14940 (N_14940,N_14520,N_14747);
nand U14941 (N_14941,N_14728,N_14470);
xnor U14942 (N_14942,N_14682,N_14514);
and U14943 (N_14943,N_14475,N_14614);
xor U14944 (N_14944,N_14506,N_14695);
nor U14945 (N_14945,N_14661,N_14743);
nand U14946 (N_14946,N_14621,N_14797);
nand U14947 (N_14947,N_14757,N_14518);
nand U14948 (N_14948,N_14571,N_14444);
or U14949 (N_14949,N_14461,N_14618);
nand U14950 (N_14950,N_14516,N_14774);
xnor U14951 (N_14951,N_14510,N_14446);
or U14952 (N_14952,N_14619,N_14744);
and U14953 (N_14953,N_14428,N_14615);
and U14954 (N_14954,N_14593,N_14529);
nand U14955 (N_14955,N_14472,N_14545);
nand U14956 (N_14956,N_14760,N_14554);
xnor U14957 (N_14957,N_14611,N_14734);
xnor U14958 (N_14958,N_14749,N_14440);
xnor U14959 (N_14959,N_14718,N_14597);
xor U14960 (N_14960,N_14433,N_14416);
and U14961 (N_14961,N_14585,N_14493);
and U14962 (N_14962,N_14466,N_14658);
nor U14963 (N_14963,N_14638,N_14447);
and U14964 (N_14964,N_14793,N_14548);
or U14965 (N_14965,N_14781,N_14709);
and U14966 (N_14966,N_14476,N_14697);
nand U14967 (N_14967,N_14400,N_14787);
nand U14968 (N_14968,N_14500,N_14668);
xor U14969 (N_14969,N_14425,N_14788);
xor U14970 (N_14970,N_14503,N_14576);
xor U14971 (N_14971,N_14414,N_14677);
nand U14972 (N_14972,N_14672,N_14617);
xor U14973 (N_14973,N_14505,N_14402);
nor U14974 (N_14974,N_14730,N_14574);
nand U14975 (N_14975,N_14627,N_14623);
nor U14976 (N_14976,N_14724,N_14696);
and U14977 (N_14977,N_14578,N_14650);
and U14978 (N_14978,N_14426,N_14648);
or U14979 (N_14979,N_14765,N_14556);
nor U14980 (N_14980,N_14606,N_14789);
xnor U14981 (N_14981,N_14790,N_14486);
nand U14982 (N_14982,N_14435,N_14636);
and U14983 (N_14983,N_14536,N_14538);
xor U14984 (N_14984,N_14570,N_14613);
nand U14985 (N_14985,N_14657,N_14403);
nand U14986 (N_14986,N_14474,N_14591);
nand U14987 (N_14987,N_14550,N_14676);
xnor U14988 (N_14988,N_14640,N_14580);
and U14989 (N_14989,N_14699,N_14713);
nand U14990 (N_14990,N_14732,N_14770);
nand U14991 (N_14991,N_14478,N_14588);
or U14992 (N_14992,N_14564,N_14528);
and U14993 (N_14993,N_14761,N_14720);
nor U14994 (N_14994,N_14560,N_14692);
and U14995 (N_14995,N_14544,N_14631);
nand U14996 (N_14996,N_14705,N_14628);
nand U14997 (N_14997,N_14489,N_14432);
nor U14998 (N_14998,N_14448,N_14666);
nand U14999 (N_14999,N_14622,N_14473);
nand U15000 (N_15000,N_14678,N_14515);
xnor U15001 (N_15001,N_14748,N_14706);
nand U15002 (N_15002,N_14608,N_14529);
and U15003 (N_15003,N_14535,N_14767);
nor U15004 (N_15004,N_14585,N_14693);
xor U15005 (N_15005,N_14508,N_14622);
xnor U15006 (N_15006,N_14631,N_14726);
nor U15007 (N_15007,N_14624,N_14565);
xnor U15008 (N_15008,N_14481,N_14767);
or U15009 (N_15009,N_14764,N_14674);
xor U15010 (N_15010,N_14674,N_14798);
and U15011 (N_15011,N_14433,N_14754);
nor U15012 (N_15012,N_14618,N_14566);
xor U15013 (N_15013,N_14619,N_14535);
nor U15014 (N_15014,N_14531,N_14472);
nand U15015 (N_15015,N_14537,N_14793);
or U15016 (N_15016,N_14547,N_14546);
nor U15017 (N_15017,N_14430,N_14655);
xor U15018 (N_15018,N_14632,N_14486);
or U15019 (N_15019,N_14733,N_14578);
or U15020 (N_15020,N_14751,N_14633);
or U15021 (N_15021,N_14572,N_14710);
or U15022 (N_15022,N_14690,N_14534);
nor U15023 (N_15023,N_14625,N_14766);
and U15024 (N_15024,N_14434,N_14789);
nand U15025 (N_15025,N_14646,N_14629);
nor U15026 (N_15026,N_14748,N_14538);
and U15027 (N_15027,N_14498,N_14725);
and U15028 (N_15028,N_14632,N_14710);
or U15029 (N_15029,N_14519,N_14564);
nor U15030 (N_15030,N_14423,N_14437);
nand U15031 (N_15031,N_14411,N_14474);
nand U15032 (N_15032,N_14415,N_14692);
xor U15033 (N_15033,N_14653,N_14750);
nand U15034 (N_15034,N_14581,N_14419);
or U15035 (N_15035,N_14649,N_14578);
nor U15036 (N_15036,N_14468,N_14665);
and U15037 (N_15037,N_14720,N_14515);
and U15038 (N_15038,N_14684,N_14796);
xnor U15039 (N_15039,N_14565,N_14409);
and U15040 (N_15040,N_14420,N_14730);
xnor U15041 (N_15041,N_14796,N_14622);
xor U15042 (N_15042,N_14484,N_14664);
nand U15043 (N_15043,N_14717,N_14460);
nor U15044 (N_15044,N_14746,N_14542);
nand U15045 (N_15045,N_14533,N_14692);
or U15046 (N_15046,N_14554,N_14697);
xor U15047 (N_15047,N_14410,N_14615);
xor U15048 (N_15048,N_14476,N_14515);
and U15049 (N_15049,N_14663,N_14560);
nor U15050 (N_15050,N_14530,N_14678);
nor U15051 (N_15051,N_14571,N_14684);
xor U15052 (N_15052,N_14711,N_14417);
nor U15053 (N_15053,N_14584,N_14697);
and U15054 (N_15054,N_14765,N_14404);
nand U15055 (N_15055,N_14592,N_14410);
xor U15056 (N_15056,N_14643,N_14540);
nand U15057 (N_15057,N_14632,N_14640);
or U15058 (N_15058,N_14763,N_14582);
nand U15059 (N_15059,N_14798,N_14459);
xnor U15060 (N_15060,N_14564,N_14706);
nand U15061 (N_15061,N_14746,N_14794);
xnor U15062 (N_15062,N_14435,N_14476);
xnor U15063 (N_15063,N_14567,N_14453);
nand U15064 (N_15064,N_14734,N_14542);
xnor U15065 (N_15065,N_14740,N_14482);
and U15066 (N_15066,N_14722,N_14493);
xnor U15067 (N_15067,N_14575,N_14461);
nor U15068 (N_15068,N_14699,N_14752);
or U15069 (N_15069,N_14435,N_14559);
and U15070 (N_15070,N_14554,N_14750);
nor U15071 (N_15071,N_14778,N_14553);
nand U15072 (N_15072,N_14475,N_14530);
nand U15073 (N_15073,N_14569,N_14644);
xnor U15074 (N_15074,N_14479,N_14715);
and U15075 (N_15075,N_14737,N_14787);
nor U15076 (N_15076,N_14489,N_14496);
nor U15077 (N_15077,N_14644,N_14435);
nand U15078 (N_15078,N_14421,N_14783);
and U15079 (N_15079,N_14550,N_14723);
xor U15080 (N_15080,N_14705,N_14408);
nor U15081 (N_15081,N_14450,N_14568);
or U15082 (N_15082,N_14732,N_14642);
nand U15083 (N_15083,N_14719,N_14773);
nand U15084 (N_15084,N_14725,N_14508);
or U15085 (N_15085,N_14693,N_14766);
nor U15086 (N_15086,N_14414,N_14505);
nand U15087 (N_15087,N_14428,N_14698);
nor U15088 (N_15088,N_14444,N_14740);
and U15089 (N_15089,N_14755,N_14584);
or U15090 (N_15090,N_14540,N_14458);
nand U15091 (N_15091,N_14779,N_14419);
nor U15092 (N_15092,N_14695,N_14650);
xor U15093 (N_15093,N_14535,N_14797);
and U15094 (N_15094,N_14455,N_14660);
and U15095 (N_15095,N_14709,N_14784);
or U15096 (N_15096,N_14759,N_14611);
nand U15097 (N_15097,N_14531,N_14510);
nand U15098 (N_15098,N_14678,N_14469);
nand U15099 (N_15099,N_14573,N_14662);
nand U15100 (N_15100,N_14709,N_14559);
and U15101 (N_15101,N_14416,N_14543);
xor U15102 (N_15102,N_14644,N_14458);
nand U15103 (N_15103,N_14542,N_14794);
nor U15104 (N_15104,N_14415,N_14514);
nand U15105 (N_15105,N_14742,N_14619);
and U15106 (N_15106,N_14609,N_14688);
or U15107 (N_15107,N_14756,N_14626);
and U15108 (N_15108,N_14502,N_14729);
nor U15109 (N_15109,N_14736,N_14712);
nor U15110 (N_15110,N_14423,N_14764);
nand U15111 (N_15111,N_14421,N_14740);
xor U15112 (N_15112,N_14472,N_14678);
nand U15113 (N_15113,N_14616,N_14723);
or U15114 (N_15114,N_14567,N_14637);
and U15115 (N_15115,N_14636,N_14586);
or U15116 (N_15116,N_14417,N_14443);
or U15117 (N_15117,N_14588,N_14657);
xor U15118 (N_15118,N_14734,N_14606);
or U15119 (N_15119,N_14679,N_14542);
nor U15120 (N_15120,N_14548,N_14720);
xor U15121 (N_15121,N_14583,N_14706);
nand U15122 (N_15122,N_14550,N_14677);
and U15123 (N_15123,N_14410,N_14465);
and U15124 (N_15124,N_14578,N_14745);
nand U15125 (N_15125,N_14417,N_14702);
nor U15126 (N_15126,N_14455,N_14448);
xor U15127 (N_15127,N_14602,N_14676);
and U15128 (N_15128,N_14500,N_14659);
and U15129 (N_15129,N_14454,N_14511);
or U15130 (N_15130,N_14561,N_14797);
or U15131 (N_15131,N_14560,N_14496);
nand U15132 (N_15132,N_14707,N_14418);
xnor U15133 (N_15133,N_14436,N_14430);
and U15134 (N_15134,N_14412,N_14555);
and U15135 (N_15135,N_14649,N_14494);
or U15136 (N_15136,N_14434,N_14456);
or U15137 (N_15137,N_14535,N_14638);
nor U15138 (N_15138,N_14417,N_14538);
and U15139 (N_15139,N_14539,N_14599);
or U15140 (N_15140,N_14515,N_14599);
and U15141 (N_15141,N_14479,N_14562);
and U15142 (N_15142,N_14543,N_14708);
or U15143 (N_15143,N_14668,N_14612);
nand U15144 (N_15144,N_14491,N_14437);
nor U15145 (N_15145,N_14465,N_14697);
or U15146 (N_15146,N_14677,N_14467);
nor U15147 (N_15147,N_14694,N_14656);
nand U15148 (N_15148,N_14576,N_14679);
or U15149 (N_15149,N_14506,N_14525);
xor U15150 (N_15150,N_14675,N_14515);
or U15151 (N_15151,N_14476,N_14443);
nand U15152 (N_15152,N_14433,N_14758);
and U15153 (N_15153,N_14603,N_14733);
nand U15154 (N_15154,N_14466,N_14696);
xnor U15155 (N_15155,N_14563,N_14656);
or U15156 (N_15156,N_14548,N_14746);
xnor U15157 (N_15157,N_14710,N_14790);
or U15158 (N_15158,N_14432,N_14614);
nor U15159 (N_15159,N_14648,N_14568);
xnor U15160 (N_15160,N_14749,N_14792);
and U15161 (N_15161,N_14789,N_14722);
and U15162 (N_15162,N_14789,N_14642);
or U15163 (N_15163,N_14715,N_14621);
nor U15164 (N_15164,N_14479,N_14417);
xor U15165 (N_15165,N_14729,N_14758);
nand U15166 (N_15166,N_14785,N_14603);
or U15167 (N_15167,N_14775,N_14412);
nand U15168 (N_15168,N_14562,N_14539);
nand U15169 (N_15169,N_14465,N_14781);
or U15170 (N_15170,N_14637,N_14701);
nor U15171 (N_15171,N_14716,N_14410);
nand U15172 (N_15172,N_14515,N_14484);
or U15173 (N_15173,N_14619,N_14453);
xor U15174 (N_15174,N_14591,N_14502);
and U15175 (N_15175,N_14761,N_14608);
or U15176 (N_15176,N_14700,N_14734);
or U15177 (N_15177,N_14532,N_14521);
nand U15178 (N_15178,N_14626,N_14400);
nor U15179 (N_15179,N_14502,N_14688);
xor U15180 (N_15180,N_14749,N_14430);
nand U15181 (N_15181,N_14640,N_14788);
nor U15182 (N_15182,N_14787,N_14770);
or U15183 (N_15183,N_14680,N_14759);
xor U15184 (N_15184,N_14621,N_14522);
xnor U15185 (N_15185,N_14614,N_14612);
nor U15186 (N_15186,N_14543,N_14483);
nor U15187 (N_15187,N_14435,N_14768);
or U15188 (N_15188,N_14640,N_14755);
nand U15189 (N_15189,N_14419,N_14792);
xor U15190 (N_15190,N_14623,N_14597);
or U15191 (N_15191,N_14479,N_14706);
nor U15192 (N_15192,N_14596,N_14557);
xor U15193 (N_15193,N_14740,N_14672);
xnor U15194 (N_15194,N_14588,N_14790);
xnor U15195 (N_15195,N_14672,N_14548);
nand U15196 (N_15196,N_14640,N_14445);
nor U15197 (N_15197,N_14415,N_14664);
and U15198 (N_15198,N_14740,N_14695);
nor U15199 (N_15199,N_14688,N_14525);
and U15200 (N_15200,N_15147,N_14928);
nor U15201 (N_15201,N_15109,N_14853);
nand U15202 (N_15202,N_14916,N_14860);
nand U15203 (N_15203,N_15118,N_14809);
nor U15204 (N_15204,N_15151,N_15000);
and U15205 (N_15205,N_14927,N_14847);
nand U15206 (N_15206,N_14863,N_15120);
nor U15207 (N_15207,N_14816,N_15005);
or U15208 (N_15208,N_15158,N_15076);
xor U15209 (N_15209,N_15077,N_15171);
xor U15210 (N_15210,N_14901,N_14957);
nor U15211 (N_15211,N_15061,N_14970);
or U15212 (N_15212,N_14905,N_15153);
nor U15213 (N_15213,N_14993,N_14880);
xor U15214 (N_15214,N_15152,N_15090);
nand U15215 (N_15215,N_15006,N_15156);
xor U15216 (N_15216,N_14969,N_15154);
nor U15217 (N_15217,N_14845,N_15085);
nand U15218 (N_15218,N_14828,N_14836);
xnor U15219 (N_15219,N_14861,N_14887);
nand U15220 (N_15220,N_15102,N_15064);
nand U15221 (N_15221,N_15081,N_15115);
xor U15222 (N_15222,N_15044,N_15092);
and U15223 (N_15223,N_14884,N_15124);
nor U15224 (N_15224,N_14923,N_15049);
nand U15225 (N_15225,N_14823,N_14800);
and U15226 (N_15226,N_15123,N_15140);
and U15227 (N_15227,N_14839,N_15180);
nand U15228 (N_15228,N_15088,N_15071);
nand U15229 (N_15229,N_15160,N_15028);
or U15230 (N_15230,N_15125,N_14891);
xnor U15231 (N_15231,N_14911,N_15117);
or U15232 (N_15232,N_15083,N_14908);
and U15233 (N_15233,N_15106,N_15057);
and U15234 (N_15234,N_14972,N_14895);
and U15235 (N_15235,N_14904,N_14801);
and U15236 (N_15236,N_15013,N_15136);
nor U15237 (N_15237,N_14940,N_14837);
nand U15238 (N_15238,N_15165,N_14941);
nor U15239 (N_15239,N_15078,N_15075);
nor U15240 (N_15240,N_14854,N_14840);
nand U15241 (N_15241,N_15003,N_15034);
and U15242 (N_15242,N_15048,N_14919);
and U15243 (N_15243,N_15027,N_14843);
nor U15244 (N_15244,N_14900,N_15186);
nand U15245 (N_15245,N_14890,N_15073);
xor U15246 (N_15246,N_15195,N_14902);
and U15247 (N_15247,N_14859,N_15111);
or U15248 (N_15248,N_15063,N_14952);
xor U15249 (N_15249,N_14811,N_14846);
and U15250 (N_15250,N_14945,N_14917);
and U15251 (N_15251,N_15119,N_15146);
and U15252 (N_15252,N_14804,N_14925);
and U15253 (N_15253,N_15187,N_15086);
or U15254 (N_15254,N_15197,N_14985);
nand U15255 (N_15255,N_14942,N_14921);
or U15256 (N_15256,N_14949,N_15060);
nand U15257 (N_15257,N_15132,N_14934);
and U15258 (N_15258,N_14812,N_15101);
and U15259 (N_15259,N_14947,N_15131);
nor U15260 (N_15260,N_15030,N_14879);
or U15261 (N_15261,N_15108,N_15052);
xor U15262 (N_15262,N_14991,N_14935);
nand U15263 (N_15263,N_15189,N_15020);
nand U15264 (N_15264,N_14933,N_15056);
or U15265 (N_15265,N_15084,N_14877);
or U15266 (N_15266,N_14903,N_15142);
nand U15267 (N_15267,N_14838,N_15135);
xnor U15268 (N_15268,N_15033,N_14960);
nand U15269 (N_15269,N_15193,N_14842);
xor U15270 (N_15270,N_15041,N_14876);
xor U15271 (N_15271,N_14959,N_15127);
or U15272 (N_15272,N_15051,N_15178);
or U15273 (N_15273,N_14924,N_15031);
or U15274 (N_15274,N_15017,N_14990);
nor U15275 (N_15275,N_14892,N_14871);
and U15276 (N_15276,N_15148,N_14978);
nor U15277 (N_15277,N_14951,N_14995);
and U15278 (N_15278,N_15008,N_14963);
xor U15279 (N_15279,N_15173,N_14815);
or U15280 (N_15280,N_14936,N_14943);
and U15281 (N_15281,N_14896,N_15054);
xor U15282 (N_15282,N_15068,N_15045);
or U15283 (N_15283,N_14849,N_14906);
nor U15284 (N_15284,N_14899,N_14888);
xor U15285 (N_15285,N_14869,N_15177);
nand U15286 (N_15286,N_15163,N_14817);
and U15287 (N_15287,N_14964,N_15058);
and U15288 (N_15288,N_15129,N_14973);
or U15289 (N_15289,N_15059,N_15175);
and U15290 (N_15290,N_14954,N_14992);
nand U15291 (N_15291,N_15097,N_15122);
or U15292 (N_15292,N_14999,N_14855);
nand U15293 (N_15293,N_15066,N_15168);
or U15294 (N_15294,N_15065,N_14979);
nor U15295 (N_15295,N_14950,N_14810);
nand U15296 (N_15296,N_14866,N_15026);
xor U15297 (N_15297,N_15004,N_14805);
nand U15298 (N_15298,N_14883,N_15198);
nor U15299 (N_15299,N_14918,N_14989);
xor U15300 (N_15300,N_14841,N_14803);
nand U15301 (N_15301,N_14835,N_14833);
nor U15302 (N_15302,N_14894,N_14832);
nor U15303 (N_15303,N_15087,N_14850);
nand U15304 (N_15304,N_14873,N_15167);
nand U15305 (N_15305,N_14889,N_15018);
and U15306 (N_15306,N_15093,N_15121);
or U15307 (N_15307,N_14965,N_15022);
xnor U15308 (N_15308,N_14994,N_15103);
nor U15309 (N_15309,N_15082,N_15188);
nor U15310 (N_15310,N_15007,N_14829);
nand U15311 (N_15311,N_14820,N_15032);
nand U15312 (N_15312,N_14914,N_14856);
xor U15313 (N_15313,N_14920,N_14819);
nand U15314 (N_15314,N_15183,N_15062);
nand U15315 (N_15315,N_15010,N_15029);
xor U15316 (N_15316,N_14808,N_14814);
xnor U15317 (N_15317,N_14864,N_14834);
or U15318 (N_15318,N_15134,N_14885);
nor U15319 (N_15319,N_15199,N_15116);
xnor U15320 (N_15320,N_14912,N_14851);
nand U15321 (N_15321,N_14930,N_15036);
xor U15322 (N_15322,N_15172,N_14848);
and U15323 (N_15323,N_14898,N_15162);
nor U15324 (N_15324,N_15100,N_15046);
xnor U15325 (N_15325,N_15190,N_14875);
nand U15326 (N_15326,N_15094,N_15144);
nand U15327 (N_15327,N_14881,N_14862);
nand U15328 (N_15328,N_14858,N_14961);
nor U15329 (N_15329,N_15196,N_15164);
or U15330 (N_15330,N_14946,N_15169);
or U15331 (N_15331,N_14984,N_15037);
or U15332 (N_15332,N_15176,N_14955);
nand U15333 (N_15333,N_14938,N_15128);
or U15334 (N_15334,N_15130,N_14986);
xnor U15335 (N_15335,N_14806,N_14824);
and U15336 (N_15336,N_14909,N_15112);
nand U15337 (N_15337,N_14910,N_14987);
or U15338 (N_15338,N_14802,N_15149);
or U15339 (N_15339,N_14958,N_15099);
xnor U15340 (N_15340,N_15110,N_14974);
xnor U15341 (N_15341,N_15021,N_15079);
or U15342 (N_15342,N_15023,N_15067);
or U15343 (N_15343,N_14893,N_14981);
nor U15344 (N_15344,N_15042,N_15184);
xnor U15345 (N_15345,N_14998,N_15011);
or U15346 (N_15346,N_15069,N_15192);
or U15347 (N_15347,N_15001,N_15040);
nor U15348 (N_15348,N_15080,N_15145);
and U15349 (N_15349,N_15053,N_15074);
xnor U15350 (N_15350,N_15091,N_15166);
nor U15351 (N_15351,N_15096,N_15181);
nor U15352 (N_15352,N_14865,N_15114);
nor U15353 (N_15353,N_14966,N_15015);
nand U15354 (N_15354,N_14913,N_15194);
or U15355 (N_15355,N_14874,N_15072);
and U15356 (N_15356,N_14983,N_15055);
and U15357 (N_15357,N_14915,N_15002);
nor U15358 (N_15358,N_15105,N_14830);
or U15359 (N_15359,N_14818,N_14929);
nor U15360 (N_15360,N_14976,N_15043);
or U15361 (N_15361,N_14997,N_14852);
nor U15362 (N_15362,N_14827,N_15038);
nor U15363 (N_15363,N_15024,N_15174);
xnor U15364 (N_15364,N_15179,N_15143);
and U15365 (N_15365,N_14878,N_14980);
or U15366 (N_15366,N_15009,N_15141);
or U15367 (N_15367,N_14813,N_14996);
nand U15368 (N_15368,N_15012,N_15113);
xor U15369 (N_15369,N_14968,N_14962);
or U15370 (N_15370,N_15025,N_14821);
xnor U15371 (N_15371,N_14988,N_14932);
xor U15372 (N_15372,N_15159,N_15089);
xor U15373 (N_15373,N_14926,N_14870);
nand U15374 (N_15374,N_15170,N_14886);
nand U15375 (N_15375,N_14971,N_14977);
and U15376 (N_15376,N_14822,N_14937);
xnor U15377 (N_15377,N_14857,N_14967);
nand U15378 (N_15378,N_14897,N_15107);
xnor U15379 (N_15379,N_15137,N_15016);
xnor U15380 (N_15380,N_14872,N_15185);
xor U15381 (N_15381,N_14868,N_15035);
nor U15382 (N_15382,N_15182,N_14931);
xnor U15383 (N_15383,N_14953,N_14956);
nor U15384 (N_15384,N_15191,N_15039);
xnor U15385 (N_15385,N_14939,N_14948);
xnor U15386 (N_15386,N_14907,N_15155);
nor U15387 (N_15387,N_15095,N_14867);
nand U15388 (N_15388,N_15070,N_15047);
or U15389 (N_15389,N_14825,N_15126);
and U15390 (N_15390,N_15133,N_14975);
nand U15391 (N_15391,N_15098,N_15157);
nand U15392 (N_15392,N_14922,N_14826);
or U15393 (N_15393,N_15138,N_15139);
or U15394 (N_15394,N_15161,N_15019);
nand U15395 (N_15395,N_15104,N_14944);
xor U15396 (N_15396,N_14807,N_15150);
nor U15397 (N_15397,N_14844,N_14982);
or U15398 (N_15398,N_15050,N_15014);
nand U15399 (N_15399,N_14831,N_14882);
nor U15400 (N_15400,N_14958,N_15123);
nor U15401 (N_15401,N_14915,N_14945);
nor U15402 (N_15402,N_14913,N_15163);
or U15403 (N_15403,N_14934,N_14830);
nor U15404 (N_15404,N_14952,N_15199);
or U15405 (N_15405,N_15119,N_15060);
or U15406 (N_15406,N_15150,N_14924);
nand U15407 (N_15407,N_14893,N_15027);
or U15408 (N_15408,N_15083,N_15106);
xnor U15409 (N_15409,N_14944,N_15008);
or U15410 (N_15410,N_15114,N_15192);
nor U15411 (N_15411,N_14999,N_15193);
nand U15412 (N_15412,N_15084,N_15142);
xnor U15413 (N_15413,N_14945,N_14981);
nor U15414 (N_15414,N_14894,N_14912);
nor U15415 (N_15415,N_15071,N_15180);
and U15416 (N_15416,N_15040,N_15138);
xor U15417 (N_15417,N_14851,N_15031);
nand U15418 (N_15418,N_15179,N_15005);
or U15419 (N_15419,N_14820,N_14880);
nand U15420 (N_15420,N_14848,N_14993);
or U15421 (N_15421,N_14866,N_14870);
xor U15422 (N_15422,N_15088,N_15093);
nand U15423 (N_15423,N_14940,N_15105);
or U15424 (N_15424,N_15085,N_15139);
and U15425 (N_15425,N_15142,N_14874);
and U15426 (N_15426,N_15052,N_15184);
and U15427 (N_15427,N_14851,N_14841);
xnor U15428 (N_15428,N_15195,N_15077);
xor U15429 (N_15429,N_14956,N_15022);
nand U15430 (N_15430,N_15021,N_15071);
nand U15431 (N_15431,N_14820,N_14953);
xnor U15432 (N_15432,N_14882,N_14918);
nand U15433 (N_15433,N_15111,N_14891);
and U15434 (N_15434,N_14980,N_15107);
and U15435 (N_15435,N_15007,N_15162);
nand U15436 (N_15436,N_14931,N_14837);
and U15437 (N_15437,N_15119,N_15109);
or U15438 (N_15438,N_15059,N_15156);
nor U15439 (N_15439,N_15116,N_14936);
or U15440 (N_15440,N_14995,N_15184);
or U15441 (N_15441,N_15004,N_15194);
nor U15442 (N_15442,N_14976,N_14889);
nand U15443 (N_15443,N_15170,N_14809);
xor U15444 (N_15444,N_14938,N_14926);
and U15445 (N_15445,N_14901,N_15182);
nand U15446 (N_15446,N_15119,N_15198);
or U15447 (N_15447,N_14882,N_15002);
xnor U15448 (N_15448,N_14866,N_15041);
and U15449 (N_15449,N_14834,N_15007);
and U15450 (N_15450,N_14997,N_15152);
nor U15451 (N_15451,N_15166,N_15113);
or U15452 (N_15452,N_15197,N_15183);
nor U15453 (N_15453,N_15167,N_14839);
and U15454 (N_15454,N_14922,N_15185);
or U15455 (N_15455,N_15001,N_15120);
or U15456 (N_15456,N_14800,N_15146);
xor U15457 (N_15457,N_15047,N_15058);
and U15458 (N_15458,N_14960,N_15007);
xnor U15459 (N_15459,N_14950,N_14971);
nor U15460 (N_15460,N_15005,N_15093);
and U15461 (N_15461,N_14853,N_15188);
nor U15462 (N_15462,N_14957,N_14845);
and U15463 (N_15463,N_15186,N_14993);
or U15464 (N_15464,N_15192,N_15106);
and U15465 (N_15465,N_14986,N_14850);
nor U15466 (N_15466,N_15171,N_15186);
nor U15467 (N_15467,N_14869,N_15099);
nor U15468 (N_15468,N_14982,N_15052);
xor U15469 (N_15469,N_14945,N_14804);
nand U15470 (N_15470,N_15034,N_14857);
nand U15471 (N_15471,N_15099,N_15199);
and U15472 (N_15472,N_14953,N_14852);
xor U15473 (N_15473,N_14858,N_14944);
xnor U15474 (N_15474,N_14898,N_14810);
xor U15475 (N_15475,N_14847,N_15048);
or U15476 (N_15476,N_15095,N_15094);
and U15477 (N_15477,N_14944,N_15132);
and U15478 (N_15478,N_15054,N_14831);
nand U15479 (N_15479,N_15092,N_15167);
nor U15480 (N_15480,N_14881,N_15066);
or U15481 (N_15481,N_15126,N_14916);
or U15482 (N_15482,N_14942,N_15030);
xor U15483 (N_15483,N_14923,N_15016);
xor U15484 (N_15484,N_14906,N_14872);
nand U15485 (N_15485,N_15041,N_14961);
and U15486 (N_15486,N_15031,N_15024);
nand U15487 (N_15487,N_15173,N_15067);
nand U15488 (N_15488,N_14989,N_14991);
and U15489 (N_15489,N_15158,N_14836);
or U15490 (N_15490,N_14926,N_15014);
nor U15491 (N_15491,N_15002,N_14834);
nand U15492 (N_15492,N_14937,N_15052);
nand U15493 (N_15493,N_15013,N_15107);
nor U15494 (N_15494,N_15167,N_15082);
nor U15495 (N_15495,N_14808,N_15090);
or U15496 (N_15496,N_15028,N_14854);
nand U15497 (N_15497,N_15068,N_15195);
nand U15498 (N_15498,N_14968,N_14933);
and U15499 (N_15499,N_14952,N_14979);
or U15500 (N_15500,N_15033,N_15023);
or U15501 (N_15501,N_14883,N_15111);
and U15502 (N_15502,N_14977,N_15154);
or U15503 (N_15503,N_15099,N_15187);
or U15504 (N_15504,N_14943,N_15005);
or U15505 (N_15505,N_14803,N_15196);
nor U15506 (N_15506,N_15125,N_14902);
and U15507 (N_15507,N_15170,N_14807);
or U15508 (N_15508,N_14825,N_15170);
nand U15509 (N_15509,N_14869,N_15064);
or U15510 (N_15510,N_14901,N_14837);
and U15511 (N_15511,N_15089,N_15010);
or U15512 (N_15512,N_14955,N_15189);
xnor U15513 (N_15513,N_15055,N_14973);
nand U15514 (N_15514,N_15072,N_14984);
and U15515 (N_15515,N_15036,N_15050);
nand U15516 (N_15516,N_15125,N_15191);
nor U15517 (N_15517,N_14824,N_14877);
or U15518 (N_15518,N_15144,N_15014);
nand U15519 (N_15519,N_15072,N_15172);
xor U15520 (N_15520,N_15159,N_14815);
or U15521 (N_15521,N_15039,N_14971);
nor U15522 (N_15522,N_15123,N_15197);
nor U15523 (N_15523,N_15139,N_15029);
or U15524 (N_15524,N_15166,N_14983);
nand U15525 (N_15525,N_14861,N_15092);
or U15526 (N_15526,N_15025,N_15167);
nor U15527 (N_15527,N_15044,N_14851);
xnor U15528 (N_15528,N_15064,N_14978);
nand U15529 (N_15529,N_15138,N_15184);
nor U15530 (N_15530,N_14860,N_14982);
xor U15531 (N_15531,N_15075,N_14970);
nor U15532 (N_15532,N_15026,N_15151);
nor U15533 (N_15533,N_15111,N_14949);
nor U15534 (N_15534,N_14839,N_14830);
xor U15535 (N_15535,N_15073,N_14905);
xor U15536 (N_15536,N_15176,N_14930);
xor U15537 (N_15537,N_15032,N_15161);
or U15538 (N_15538,N_15038,N_15060);
xor U15539 (N_15539,N_14915,N_14921);
and U15540 (N_15540,N_14935,N_15063);
xnor U15541 (N_15541,N_14898,N_15007);
and U15542 (N_15542,N_14825,N_15193);
or U15543 (N_15543,N_15015,N_14989);
nand U15544 (N_15544,N_14884,N_14910);
nor U15545 (N_15545,N_15112,N_15180);
or U15546 (N_15546,N_15055,N_15128);
or U15547 (N_15547,N_14940,N_15075);
xnor U15548 (N_15548,N_14927,N_15064);
and U15549 (N_15549,N_14909,N_15142);
nor U15550 (N_15550,N_14809,N_14813);
xor U15551 (N_15551,N_15102,N_14938);
nand U15552 (N_15552,N_15123,N_15168);
and U15553 (N_15553,N_14852,N_15138);
xnor U15554 (N_15554,N_14923,N_14855);
nand U15555 (N_15555,N_14859,N_14889);
and U15556 (N_15556,N_14808,N_14892);
nor U15557 (N_15557,N_14837,N_15019);
xor U15558 (N_15558,N_14907,N_15138);
xnor U15559 (N_15559,N_14817,N_14812);
or U15560 (N_15560,N_15102,N_15068);
nand U15561 (N_15561,N_14984,N_15054);
nor U15562 (N_15562,N_15181,N_14915);
xnor U15563 (N_15563,N_15012,N_15089);
nand U15564 (N_15564,N_15066,N_15073);
nor U15565 (N_15565,N_15096,N_14898);
and U15566 (N_15566,N_15058,N_15032);
and U15567 (N_15567,N_14810,N_14897);
nand U15568 (N_15568,N_15005,N_14868);
xor U15569 (N_15569,N_15160,N_15199);
xnor U15570 (N_15570,N_14956,N_15107);
or U15571 (N_15571,N_15142,N_15141);
and U15572 (N_15572,N_14979,N_15176);
and U15573 (N_15573,N_14837,N_15116);
and U15574 (N_15574,N_14905,N_14937);
and U15575 (N_15575,N_15187,N_15051);
or U15576 (N_15576,N_14863,N_14801);
and U15577 (N_15577,N_14833,N_15023);
nand U15578 (N_15578,N_15143,N_15050);
or U15579 (N_15579,N_14913,N_14998);
nand U15580 (N_15580,N_14903,N_14918);
nand U15581 (N_15581,N_15169,N_15160);
xor U15582 (N_15582,N_15038,N_15126);
or U15583 (N_15583,N_15082,N_14917);
nand U15584 (N_15584,N_15060,N_15160);
nand U15585 (N_15585,N_14982,N_14872);
or U15586 (N_15586,N_15126,N_15184);
or U15587 (N_15587,N_15052,N_15002);
nand U15588 (N_15588,N_14908,N_14989);
and U15589 (N_15589,N_15020,N_15118);
nor U15590 (N_15590,N_15113,N_14932);
or U15591 (N_15591,N_15003,N_14980);
and U15592 (N_15592,N_14874,N_14834);
or U15593 (N_15593,N_15188,N_14959);
nand U15594 (N_15594,N_14915,N_14876);
nand U15595 (N_15595,N_14937,N_15104);
or U15596 (N_15596,N_15071,N_14974);
xnor U15597 (N_15597,N_14874,N_14828);
and U15598 (N_15598,N_14855,N_15089);
xor U15599 (N_15599,N_15071,N_15182);
and U15600 (N_15600,N_15517,N_15450);
nor U15601 (N_15601,N_15424,N_15374);
and U15602 (N_15602,N_15500,N_15285);
and U15603 (N_15603,N_15435,N_15428);
xnor U15604 (N_15604,N_15440,N_15378);
and U15605 (N_15605,N_15337,N_15361);
and U15606 (N_15606,N_15544,N_15298);
nor U15607 (N_15607,N_15347,N_15321);
or U15608 (N_15608,N_15372,N_15259);
and U15609 (N_15609,N_15338,N_15322);
nand U15610 (N_15610,N_15496,N_15559);
or U15611 (N_15611,N_15569,N_15340);
and U15612 (N_15612,N_15379,N_15385);
and U15613 (N_15613,N_15245,N_15525);
xnor U15614 (N_15614,N_15498,N_15466);
xor U15615 (N_15615,N_15309,N_15279);
or U15616 (N_15616,N_15409,N_15214);
or U15617 (N_15617,N_15402,N_15530);
nor U15618 (N_15618,N_15578,N_15494);
xor U15619 (N_15619,N_15389,N_15513);
and U15620 (N_15620,N_15594,N_15277);
nand U15621 (N_15621,N_15456,N_15420);
nor U15622 (N_15622,N_15505,N_15463);
nand U15623 (N_15623,N_15327,N_15455);
xnor U15624 (N_15624,N_15438,N_15218);
nand U15625 (N_15625,N_15224,N_15432);
nor U15626 (N_15626,N_15572,N_15430);
xnor U15627 (N_15627,N_15223,N_15464);
nor U15628 (N_15628,N_15394,N_15370);
or U15629 (N_15629,N_15215,N_15256);
or U15630 (N_15630,N_15492,N_15357);
nor U15631 (N_15631,N_15558,N_15523);
and U15632 (N_15632,N_15547,N_15244);
nand U15633 (N_15633,N_15242,N_15565);
or U15634 (N_15634,N_15273,N_15299);
nor U15635 (N_15635,N_15446,N_15490);
nor U15636 (N_15636,N_15254,N_15520);
nor U15637 (N_15637,N_15581,N_15468);
and U15638 (N_15638,N_15236,N_15552);
nand U15639 (N_15639,N_15509,N_15445);
or U15640 (N_15640,N_15238,N_15323);
and U15641 (N_15641,N_15307,N_15425);
nor U15642 (N_15642,N_15577,N_15566);
nand U15643 (N_15643,N_15380,N_15333);
or U15644 (N_15644,N_15518,N_15336);
nor U15645 (N_15645,N_15411,N_15568);
xnor U15646 (N_15646,N_15251,N_15452);
or U15647 (N_15647,N_15349,N_15553);
and U15648 (N_15648,N_15548,N_15493);
nand U15649 (N_15649,N_15228,N_15339);
nand U15650 (N_15650,N_15431,N_15437);
and U15651 (N_15651,N_15417,N_15589);
nand U15652 (N_15652,N_15232,N_15293);
nor U15653 (N_15653,N_15311,N_15272);
xnor U15654 (N_15654,N_15316,N_15229);
nand U15655 (N_15655,N_15376,N_15392);
or U15656 (N_15656,N_15555,N_15308);
and U15657 (N_15657,N_15222,N_15270);
nor U15658 (N_15658,N_15382,N_15262);
nand U15659 (N_15659,N_15250,N_15599);
nand U15660 (N_15660,N_15528,N_15536);
and U15661 (N_15661,N_15551,N_15433);
xor U15662 (N_15662,N_15516,N_15355);
nor U15663 (N_15663,N_15332,N_15358);
or U15664 (N_15664,N_15596,N_15470);
or U15665 (N_15665,N_15534,N_15451);
nor U15666 (N_15666,N_15227,N_15287);
nand U15667 (N_15667,N_15454,N_15314);
nand U15668 (N_15668,N_15571,N_15297);
nand U15669 (N_15669,N_15502,N_15434);
nor U15670 (N_15670,N_15258,N_15248);
nand U15671 (N_15671,N_15597,N_15207);
or U15672 (N_15672,N_15478,N_15306);
and U15673 (N_15673,N_15280,N_15461);
or U15674 (N_15674,N_15598,N_15482);
nor U15675 (N_15675,N_15587,N_15289);
and U15676 (N_15676,N_15532,N_15331);
xor U15677 (N_15677,N_15557,N_15217);
and U15678 (N_15678,N_15317,N_15545);
xnor U15679 (N_15679,N_15512,N_15211);
and U15680 (N_15680,N_15449,N_15441);
and U15681 (N_15681,N_15419,N_15584);
nand U15682 (N_15682,N_15260,N_15550);
or U15683 (N_15683,N_15295,N_15243);
or U15684 (N_15684,N_15474,N_15312);
or U15685 (N_15685,N_15585,N_15554);
xnor U15686 (N_15686,N_15443,N_15324);
xnor U15687 (N_15687,N_15413,N_15447);
nor U15688 (N_15688,N_15514,N_15271);
nor U15689 (N_15689,N_15234,N_15510);
and U15690 (N_15690,N_15592,N_15479);
or U15691 (N_15691,N_15202,N_15398);
nand U15692 (N_15692,N_15416,N_15286);
xor U15693 (N_15693,N_15252,N_15210);
nor U15694 (N_15694,N_15407,N_15546);
and U15695 (N_15695,N_15484,N_15368);
or U15696 (N_15696,N_15560,N_15294);
nand U15697 (N_15697,N_15562,N_15576);
xor U15698 (N_15698,N_15381,N_15415);
nor U15699 (N_15699,N_15330,N_15564);
nand U15700 (N_15700,N_15353,N_15561);
xor U15701 (N_15701,N_15458,N_15233);
or U15702 (N_15702,N_15595,N_15208);
xnor U15703 (N_15703,N_15268,N_15395);
and U15704 (N_15704,N_15475,N_15400);
and U15705 (N_15705,N_15320,N_15212);
nor U15706 (N_15706,N_15405,N_15412);
or U15707 (N_15707,N_15503,N_15539);
or U15708 (N_15708,N_15575,N_15276);
nor U15709 (N_15709,N_15329,N_15573);
or U15710 (N_15710,N_15570,N_15206);
nor U15711 (N_15711,N_15226,N_15342);
xor U15712 (N_15712,N_15352,N_15418);
nand U15713 (N_15713,N_15404,N_15302);
nor U15714 (N_15714,N_15473,N_15315);
nand U15715 (N_15715,N_15469,N_15367);
nand U15716 (N_15716,N_15531,N_15497);
and U15717 (N_15717,N_15288,N_15300);
or U15718 (N_15718,N_15350,N_15346);
and U15719 (N_15719,N_15593,N_15292);
and U15720 (N_15720,N_15393,N_15267);
nand U15721 (N_15721,N_15465,N_15290);
nand U15722 (N_15722,N_15291,N_15511);
xnor U15723 (N_15723,N_15220,N_15221);
nand U15724 (N_15724,N_15282,N_15537);
nor U15725 (N_15725,N_15556,N_15239);
or U15726 (N_15726,N_15506,N_15472);
nand U15727 (N_15727,N_15356,N_15535);
or U15728 (N_15728,N_15335,N_15540);
and U15729 (N_15729,N_15401,N_15310);
nand U15730 (N_15730,N_15489,N_15457);
or U15731 (N_15731,N_15403,N_15387);
xor U15732 (N_15732,N_15410,N_15591);
or U15733 (N_15733,N_15348,N_15487);
or U15734 (N_15734,N_15231,N_15278);
nor U15735 (N_15735,N_15524,N_15423);
nor U15736 (N_15736,N_15235,N_15319);
xnor U15737 (N_15737,N_15541,N_15240);
and U15738 (N_15738,N_15481,N_15371);
nand U15739 (N_15739,N_15363,N_15366);
nand U15740 (N_15740,N_15249,N_15359);
xnor U15741 (N_15741,N_15313,N_15390);
xnor U15742 (N_15742,N_15507,N_15460);
and U15743 (N_15743,N_15542,N_15275);
xor U15744 (N_15744,N_15426,N_15201);
xor U15745 (N_15745,N_15480,N_15486);
or U15746 (N_15746,N_15519,N_15203);
nand U15747 (N_15747,N_15422,N_15365);
xor U15748 (N_15748,N_15444,N_15508);
nor U15749 (N_15749,N_15301,N_15515);
or U15750 (N_15750,N_15406,N_15200);
or U15751 (N_15751,N_15476,N_15219);
nor U15752 (N_15752,N_15427,N_15283);
nand U15753 (N_15753,N_15216,N_15266);
xor U15754 (N_15754,N_15533,N_15281);
nand U15755 (N_15755,N_15471,N_15388);
nor U15756 (N_15756,N_15391,N_15448);
xnor U15757 (N_15757,N_15326,N_15501);
and U15758 (N_15758,N_15334,N_15442);
nor U15759 (N_15759,N_15549,N_15429);
nand U15760 (N_15760,N_15225,N_15343);
or U15761 (N_15761,N_15205,N_15375);
and U15762 (N_15762,N_15521,N_15527);
nor U15763 (N_15763,N_15213,N_15209);
nand U15764 (N_15764,N_15241,N_15383);
nor U15765 (N_15765,N_15318,N_15408);
nor U15766 (N_15766,N_15284,N_15328);
nand U15767 (N_15767,N_15499,N_15529);
nand U15768 (N_15768,N_15567,N_15459);
nor U15769 (N_15769,N_15462,N_15261);
nand U15770 (N_15770,N_15483,N_15488);
and U15771 (N_15771,N_15491,N_15485);
nand U15772 (N_15772,N_15263,N_15477);
nand U15773 (N_15773,N_15305,N_15543);
nor U15774 (N_15774,N_15247,N_15351);
nor U15775 (N_15775,N_15384,N_15586);
nor U15776 (N_15776,N_15354,N_15257);
and U15777 (N_15777,N_15396,N_15304);
xor U15778 (N_15778,N_15526,N_15421);
xnor U15779 (N_15779,N_15522,N_15360);
and U15780 (N_15780,N_15504,N_15582);
nand U15781 (N_15781,N_15345,N_15495);
nor U15782 (N_15782,N_15397,N_15377);
xnor U15783 (N_15783,N_15467,N_15230);
or U15784 (N_15784,N_15255,N_15344);
nand U15785 (N_15785,N_15265,N_15590);
or U15786 (N_15786,N_15274,N_15341);
nand U15787 (N_15787,N_15269,N_15303);
nand U15788 (N_15788,N_15453,N_15369);
nand U15789 (N_15789,N_15580,N_15414);
or U15790 (N_15790,N_15364,N_15325);
and U15791 (N_15791,N_15373,N_15264);
and U15792 (N_15792,N_15253,N_15237);
or U15793 (N_15793,N_15439,N_15579);
and U15794 (N_15794,N_15574,N_15204);
and U15795 (N_15795,N_15362,N_15386);
nor U15796 (N_15796,N_15583,N_15246);
or U15797 (N_15797,N_15563,N_15436);
and U15798 (N_15798,N_15399,N_15538);
xor U15799 (N_15799,N_15296,N_15588);
and U15800 (N_15800,N_15231,N_15591);
nor U15801 (N_15801,N_15327,N_15482);
nand U15802 (N_15802,N_15259,N_15532);
or U15803 (N_15803,N_15500,N_15582);
xor U15804 (N_15804,N_15268,N_15382);
or U15805 (N_15805,N_15410,N_15536);
xnor U15806 (N_15806,N_15332,N_15427);
nand U15807 (N_15807,N_15206,N_15290);
and U15808 (N_15808,N_15335,N_15591);
xor U15809 (N_15809,N_15323,N_15504);
nor U15810 (N_15810,N_15430,N_15294);
and U15811 (N_15811,N_15513,N_15271);
or U15812 (N_15812,N_15305,N_15431);
and U15813 (N_15813,N_15504,N_15575);
or U15814 (N_15814,N_15307,N_15320);
nand U15815 (N_15815,N_15572,N_15235);
or U15816 (N_15816,N_15216,N_15210);
and U15817 (N_15817,N_15462,N_15571);
nand U15818 (N_15818,N_15320,N_15405);
or U15819 (N_15819,N_15220,N_15262);
or U15820 (N_15820,N_15392,N_15599);
and U15821 (N_15821,N_15591,N_15419);
nor U15822 (N_15822,N_15295,N_15264);
or U15823 (N_15823,N_15222,N_15319);
nor U15824 (N_15824,N_15381,N_15582);
nand U15825 (N_15825,N_15464,N_15441);
nor U15826 (N_15826,N_15308,N_15420);
xor U15827 (N_15827,N_15520,N_15259);
nand U15828 (N_15828,N_15563,N_15231);
nand U15829 (N_15829,N_15509,N_15587);
nor U15830 (N_15830,N_15484,N_15294);
or U15831 (N_15831,N_15380,N_15233);
xnor U15832 (N_15832,N_15205,N_15248);
or U15833 (N_15833,N_15354,N_15304);
or U15834 (N_15834,N_15287,N_15339);
and U15835 (N_15835,N_15485,N_15320);
or U15836 (N_15836,N_15444,N_15252);
nor U15837 (N_15837,N_15341,N_15384);
xor U15838 (N_15838,N_15293,N_15532);
nand U15839 (N_15839,N_15404,N_15402);
nand U15840 (N_15840,N_15272,N_15336);
nor U15841 (N_15841,N_15570,N_15404);
or U15842 (N_15842,N_15468,N_15307);
and U15843 (N_15843,N_15531,N_15230);
xnor U15844 (N_15844,N_15322,N_15507);
and U15845 (N_15845,N_15549,N_15339);
or U15846 (N_15846,N_15328,N_15403);
and U15847 (N_15847,N_15471,N_15317);
and U15848 (N_15848,N_15291,N_15371);
nand U15849 (N_15849,N_15550,N_15272);
xor U15850 (N_15850,N_15272,N_15457);
nor U15851 (N_15851,N_15449,N_15322);
or U15852 (N_15852,N_15520,N_15212);
xnor U15853 (N_15853,N_15584,N_15329);
xor U15854 (N_15854,N_15343,N_15448);
nor U15855 (N_15855,N_15295,N_15307);
and U15856 (N_15856,N_15228,N_15594);
and U15857 (N_15857,N_15225,N_15223);
or U15858 (N_15858,N_15372,N_15439);
nor U15859 (N_15859,N_15491,N_15519);
and U15860 (N_15860,N_15445,N_15221);
xor U15861 (N_15861,N_15331,N_15586);
and U15862 (N_15862,N_15426,N_15578);
and U15863 (N_15863,N_15582,N_15458);
xnor U15864 (N_15864,N_15396,N_15320);
and U15865 (N_15865,N_15297,N_15213);
or U15866 (N_15866,N_15573,N_15325);
nand U15867 (N_15867,N_15243,N_15384);
or U15868 (N_15868,N_15376,N_15497);
and U15869 (N_15869,N_15366,N_15391);
xnor U15870 (N_15870,N_15359,N_15363);
and U15871 (N_15871,N_15282,N_15247);
or U15872 (N_15872,N_15303,N_15449);
nor U15873 (N_15873,N_15412,N_15372);
xnor U15874 (N_15874,N_15454,N_15224);
nor U15875 (N_15875,N_15416,N_15264);
nand U15876 (N_15876,N_15598,N_15512);
nand U15877 (N_15877,N_15326,N_15431);
xnor U15878 (N_15878,N_15455,N_15374);
and U15879 (N_15879,N_15515,N_15289);
or U15880 (N_15880,N_15407,N_15401);
nor U15881 (N_15881,N_15514,N_15350);
or U15882 (N_15882,N_15282,N_15383);
xor U15883 (N_15883,N_15244,N_15206);
nor U15884 (N_15884,N_15494,N_15308);
nor U15885 (N_15885,N_15555,N_15507);
or U15886 (N_15886,N_15446,N_15371);
xor U15887 (N_15887,N_15518,N_15207);
xnor U15888 (N_15888,N_15459,N_15587);
nand U15889 (N_15889,N_15474,N_15276);
xnor U15890 (N_15890,N_15548,N_15497);
nand U15891 (N_15891,N_15345,N_15217);
and U15892 (N_15892,N_15490,N_15562);
xnor U15893 (N_15893,N_15476,N_15572);
nand U15894 (N_15894,N_15559,N_15490);
nor U15895 (N_15895,N_15224,N_15310);
nor U15896 (N_15896,N_15563,N_15355);
nand U15897 (N_15897,N_15499,N_15429);
or U15898 (N_15898,N_15347,N_15260);
and U15899 (N_15899,N_15200,N_15377);
xor U15900 (N_15900,N_15557,N_15222);
or U15901 (N_15901,N_15452,N_15206);
or U15902 (N_15902,N_15323,N_15236);
nand U15903 (N_15903,N_15587,N_15214);
nand U15904 (N_15904,N_15286,N_15499);
nor U15905 (N_15905,N_15550,N_15252);
and U15906 (N_15906,N_15521,N_15454);
and U15907 (N_15907,N_15555,N_15380);
and U15908 (N_15908,N_15318,N_15392);
nand U15909 (N_15909,N_15521,N_15213);
or U15910 (N_15910,N_15454,N_15409);
nor U15911 (N_15911,N_15324,N_15304);
nand U15912 (N_15912,N_15525,N_15388);
xor U15913 (N_15913,N_15517,N_15488);
nand U15914 (N_15914,N_15525,N_15483);
and U15915 (N_15915,N_15598,N_15416);
nand U15916 (N_15916,N_15497,N_15360);
and U15917 (N_15917,N_15263,N_15440);
nor U15918 (N_15918,N_15457,N_15226);
nand U15919 (N_15919,N_15424,N_15299);
nor U15920 (N_15920,N_15230,N_15248);
and U15921 (N_15921,N_15598,N_15524);
xor U15922 (N_15922,N_15490,N_15394);
xor U15923 (N_15923,N_15230,N_15558);
and U15924 (N_15924,N_15264,N_15298);
xor U15925 (N_15925,N_15377,N_15356);
and U15926 (N_15926,N_15523,N_15336);
nor U15927 (N_15927,N_15337,N_15557);
and U15928 (N_15928,N_15219,N_15508);
nand U15929 (N_15929,N_15505,N_15340);
and U15930 (N_15930,N_15514,N_15531);
nand U15931 (N_15931,N_15345,N_15285);
nor U15932 (N_15932,N_15537,N_15295);
xor U15933 (N_15933,N_15399,N_15447);
nor U15934 (N_15934,N_15520,N_15444);
and U15935 (N_15935,N_15224,N_15477);
xnor U15936 (N_15936,N_15526,N_15359);
xor U15937 (N_15937,N_15276,N_15234);
nand U15938 (N_15938,N_15487,N_15422);
nor U15939 (N_15939,N_15333,N_15286);
xor U15940 (N_15940,N_15464,N_15336);
xor U15941 (N_15941,N_15562,N_15311);
nor U15942 (N_15942,N_15424,N_15312);
nor U15943 (N_15943,N_15480,N_15381);
or U15944 (N_15944,N_15402,N_15293);
nand U15945 (N_15945,N_15333,N_15573);
xor U15946 (N_15946,N_15384,N_15486);
xnor U15947 (N_15947,N_15589,N_15301);
or U15948 (N_15948,N_15270,N_15283);
and U15949 (N_15949,N_15391,N_15514);
nor U15950 (N_15950,N_15488,N_15571);
and U15951 (N_15951,N_15217,N_15598);
or U15952 (N_15952,N_15212,N_15273);
or U15953 (N_15953,N_15250,N_15446);
xor U15954 (N_15954,N_15237,N_15272);
nor U15955 (N_15955,N_15396,N_15272);
and U15956 (N_15956,N_15535,N_15436);
or U15957 (N_15957,N_15395,N_15217);
or U15958 (N_15958,N_15364,N_15545);
or U15959 (N_15959,N_15301,N_15478);
xor U15960 (N_15960,N_15410,N_15237);
nand U15961 (N_15961,N_15209,N_15237);
nand U15962 (N_15962,N_15213,N_15330);
nand U15963 (N_15963,N_15490,N_15516);
nor U15964 (N_15964,N_15559,N_15488);
nor U15965 (N_15965,N_15570,N_15507);
xnor U15966 (N_15966,N_15422,N_15240);
and U15967 (N_15967,N_15358,N_15263);
nand U15968 (N_15968,N_15442,N_15333);
xor U15969 (N_15969,N_15236,N_15569);
xor U15970 (N_15970,N_15573,N_15521);
xor U15971 (N_15971,N_15520,N_15450);
and U15972 (N_15972,N_15220,N_15538);
nand U15973 (N_15973,N_15487,N_15489);
or U15974 (N_15974,N_15293,N_15367);
nor U15975 (N_15975,N_15467,N_15519);
or U15976 (N_15976,N_15221,N_15473);
xor U15977 (N_15977,N_15234,N_15384);
and U15978 (N_15978,N_15524,N_15463);
nor U15979 (N_15979,N_15502,N_15571);
and U15980 (N_15980,N_15386,N_15493);
nand U15981 (N_15981,N_15442,N_15235);
or U15982 (N_15982,N_15446,N_15476);
nor U15983 (N_15983,N_15303,N_15206);
nand U15984 (N_15984,N_15503,N_15294);
and U15985 (N_15985,N_15298,N_15251);
nand U15986 (N_15986,N_15471,N_15352);
nand U15987 (N_15987,N_15519,N_15316);
or U15988 (N_15988,N_15281,N_15333);
xnor U15989 (N_15989,N_15472,N_15218);
nand U15990 (N_15990,N_15497,N_15266);
nand U15991 (N_15991,N_15473,N_15325);
and U15992 (N_15992,N_15407,N_15371);
nand U15993 (N_15993,N_15469,N_15412);
or U15994 (N_15994,N_15223,N_15210);
and U15995 (N_15995,N_15230,N_15240);
xor U15996 (N_15996,N_15509,N_15201);
or U15997 (N_15997,N_15326,N_15569);
xnor U15998 (N_15998,N_15452,N_15366);
or U15999 (N_15999,N_15588,N_15265);
xnor U16000 (N_16000,N_15611,N_15963);
or U16001 (N_16001,N_15897,N_15754);
nor U16002 (N_16002,N_15889,N_15741);
nand U16003 (N_16003,N_15772,N_15994);
nand U16004 (N_16004,N_15868,N_15895);
nor U16005 (N_16005,N_15990,N_15801);
nand U16006 (N_16006,N_15985,N_15669);
nor U16007 (N_16007,N_15945,N_15892);
nand U16008 (N_16008,N_15885,N_15818);
xor U16009 (N_16009,N_15796,N_15872);
and U16010 (N_16010,N_15789,N_15643);
nor U16011 (N_16011,N_15968,N_15664);
xor U16012 (N_16012,N_15859,N_15776);
and U16013 (N_16013,N_15824,N_15704);
or U16014 (N_16014,N_15902,N_15983);
nand U16015 (N_16015,N_15609,N_15615);
xor U16016 (N_16016,N_15732,N_15831);
xor U16017 (N_16017,N_15974,N_15866);
nand U16018 (N_16018,N_15761,N_15667);
xor U16019 (N_16019,N_15689,N_15840);
xor U16020 (N_16020,N_15815,N_15802);
or U16021 (N_16021,N_15708,N_15660);
and U16022 (N_16022,N_15809,N_15903);
or U16023 (N_16023,N_15896,N_15767);
nor U16024 (N_16024,N_15672,N_15680);
nor U16025 (N_16025,N_15798,N_15898);
nand U16026 (N_16026,N_15799,N_15830);
or U16027 (N_16027,N_15700,N_15663);
nor U16028 (N_16028,N_15722,N_15899);
and U16029 (N_16029,N_15774,N_15964);
and U16030 (N_16030,N_15607,N_15999);
nand U16031 (N_16031,N_15793,N_15883);
or U16032 (N_16032,N_15944,N_15942);
xnor U16033 (N_16033,N_15987,N_15684);
or U16034 (N_16034,N_15676,N_15752);
xor U16035 (N_16035,N_15804,N_15756);
and U16036 (N_16036,N_15919,N_15931);
and U16037 (N_16037,N_15744,N_15881);
or U16038 (N_16038,N_15878,N_15936);
nor U16039 (N_16039,N_15694,N_15659);
and U16040 (N_16040,N_15842,N_15650);
nand U16041 (N_16041,N_15876,N_15869);
nand U16042 (N_16042,N_15748,N_15602);
or U16043 (N_16043,N_15871,N_15965);
or U16044 (N_16044,N_15787,N_15707);
xor U16045 (N_16045,N_15907,N_15850);
xor U16046 (N_16046,N_15706,N_15717);
or U16047 (N_16047,N_15806,N_15836);
nand U16048 (N_16048,N_15906,N_15636);
and U16049 (N_16049,N_15856,N_15913);
xnor U16050 (N_16050,N_15647,N_15739);
and U16051 (N_16051,N_15870,N_15735);
nor U16052 (N_16052,N_15781,N_15803);
xor U16053 (N_16053,N_15668,N_15657);
nand U16054 (N_16054,N_15746,N_15697);
nand U16055 (N_16055,N_15751,N_15675);
nor U16056 (N_16056,N_15758,N_15665);
and U16057 (N_16057,N_15834,N_15832);
xnor U16058 (N_16058,N_15601,N_15846);
or U16059 (N_16059,N_15749,N_15841);
and U16060 (N_16060,N_15605,N_15630);
or U16061 (N_16061,N_15938,N_15645);
or U16062 (N_16062,N_15710,N_15703);
xor U16063 (N_16063,N_15890,N_15957);
or U16064 (N_16064,N_15996,N_15687);
or U16065 (N_16065,N_15825,N_15918);
nand U16066 (N_16066,N_15606,N_15783);
or U16067 (N_16067,N_15966,N_15702);
nand U16068 (N_16068,N_15853,N_15959);
xor U16069 (N_16069,N_15695,N_15674);
and U16070 (N_16070,N_15691,N_15972);
nor U16071 (N_16071,N_15613,N_15600);
nor U16072 (N_16072,N_15975,N_15768);
and U16073 (N_16073,N_15709,N_15845);
nor U16074 (N_16074,N_15688,N_15893);
nor U16075 (N_16075,N_15730,N_15860);
and U16076 (N_16076,N_15971,N_15731);
nand U16077 (N_16077,N_15843,N_15617);
or U16078 (N_16078,N_15901,N_15880);
or U16079 (N_16079,N_15848,N_15620);
and U16080 (N_16080,N_15948,N_15622);
nand U16081 (N_16081,N_15631,N_15810);
or U16082 (N_16082,N_15637,N_15629);
nor U16083 (N_16083,N_15929,N_15666);
or U16084 (N_16084,N_15656,N_15719);
nand U16085 (N_16085,N_15970,N_15978);
and U16086 (N_16086,N_15894,N_15862);
and U16087 (N_16087,N_15692,N_15921);
and U16088 (N_16088,N_15822,N_15679);
nor U16089 (N_16089,N_15808,N_15632);
and U16090 (N_16090,N_15791,N_15775);
nand U16091 (N_16091,N_15750,N_15884);
xnor U16092 (N_16092,N_15992,N_15891);
nand U16093 (N_16093,N_15956,N_15967);
xor U16094 (N_16094,N_15727,N_15973);
nand U16095 (N_16095,N_15733,N_15648);
nor U16096 (N_16096,N_15952,N_15927);
nand U16097 (N_16097,N_15770,N_15920);
nand U16098 (N_16098,N_15673,N_15816);
nand U16099 (N_16099,N_15784,N_15628);
or U16100 (N_16100,N_15950,N_15723);
and U16101 (N_16101,N_15819,N_15888);
xnor U16102 (N_16102,N_15875,N_15640);
xor U16103 (N_16103,N_15928,N_15886);
nor U16104 (N_16104,N_15934,N_15635);
and U16105 (N_16105,N_15685,N_15951);
and U16106 (N_16106,N_15827,N_15740);
xnor U16107 (N_16107,N_15788,N_15734);
nor U16108 (N_16108,N_15813,N_15955);
nand U16109 (N_16109,N_15619,N_15867);
and U16110 (N_16110,N_15771,N_15724);
nor U16111 (N_16111,N_15726,N_15721);
and U16112 (N_16112,N_15759,N_15686);
or U16113 (N_16113,N_15716,N_15743);
xnor U16114 (N_16114,N_15654,N_15812);
and U16115 (N_16115,N_15949,N_15807);
nor U16116 (N_16116,N_15641,N_15737);
and U16117 (N_16117,N_15713,N_15954);
xor U16118 (N_16118,N_15696,N_15782);
xnor U16119 (N_16119,N_15800,N_15984);
xor U16120 (N_16120,N_15797,N_15701);
or U16121 (N_16121,N_15915,N_15714);
or U16122 (N_16122,N_15779,N_15905);
and U16123 (N_16123,N_15773,N_15851);
or U16124 (N_16124,N_15821,N_15625);
or U16125 (N_16125,N_15720,N_15947);
nand U16126 (N_16126,N_15616,N_15823);
nor U16127 (N_16127,N_15833,N_15979);
nand U16128 (N_16128,N_15982,N_15926);
nand U16129 (N_16129,N_15661,N_15908);
nand U16130 (N_16130,N_15718,N_15887);
xnor U16131 (N_16131,N_15785,N_15769);
nor U16132 (N_16132,N_15849,N_15933);
or U16133 (N_16133,N_15838,N_15627);
nor U16134 (N_16134,N_15814,N_15711);
or U16135 (N_16135,N_15626,N_15837);
xnor U16136 (N_16136,N_15760,N_15925);
nand U16137 (N_16137,N_15861,N_15763);
nand U16138 (N_16138,N_15924,N_15678);
or U16139 (N_16139,N_15828,N_15604);
nor U16140 (N_16140,N_15780,N_15829);
xor U16141 (N_16141,N_15738,N_15712);
or U16142 (N_16142,N_15835,N_15614);
xor U16143 (N_16143,N_15922,N_15864);
or U16144 (N_16144,N_15805,N_15705);
nor U16145 (N_16145,N_15728,N_15683);
nor U16146 (N_16146,N_15960,N_15603);
and U16147 (N_16147,N_15981,N_15725);
or U16148 (N_16148,N_15930,N_15795);
or U16149 (N_16149,N_15764,N_15991);
xnor U16150 (N_16150,N_15790,N_15755);
or U16151 (N_16151,N_15976,N_15698);
nor U16152 (N_16152,N_15917,N_15638);
nor U16153 (N_16153,N_15995,N_15873);
nor U16154 (N_16154,N_15877,N_15715);
and U16155 (N_16155,N_15916,N_15634);
xnor U16156 (N_16156,N_15882,N_15935);
and U16157 (N_16157,N_15826,N_15874);
and U16158 (N_16158,N_15757,N_15847);
nor U16159 (N_16159,N_15729,N_15753);
nand U16160 (N_16160,N_15969,N_15977);
xnor U16161 (N_16161,N_15699,N_15946);
and U16162 (N_16162,N_15910,N_15633);
nor U16163 (N_16163,N_15858,N_15612);
nor U16164 (N_16164,N_15655,N_15653);
and U16165 (N_16165,N_15621,N_15777);
or U16166 (N_16166,N_15794,N_15693);
or U16167 (N_16167,N_15765,N_15855);
or U16168 (N_16168,N_15610,N_15644);
nor U16169 (N_16169,N_15961,N_15998);
nor U16170 (N_16170,N_15623,N_15747);
or U16171 (N_16171,N_15778,N_15912);
nor U16172 (N_16172,N_15677,N_15865);
nand U16173 (N_16173,N_15904,N_15742);
and U16174 (N_16174,N_15937,N_15940);
nor U16175 (N_16175,N_15989,N_15844);
xnor U16176 (N_16176,N_15980,N_15652);
xnor U16177 (N_16177,N_15671,N_15988);
nand U16178 (N_16178,N_15879,N_15854);
nand U16179 (N_16179,N_15943,N_15939);
nand U16180 (N_16180,N_15690,N_15900);
or U16181 (N_16181,N_15820,N_15993);
xnor U16182 (N_16182,N_15941,N_15932);
or U16183 (N_16183,N_15651,N_15909);
nor U16184 (N_16184,N_15839,N_15857);
or U16185 (N_16185,N_15642,N_15852);
or U16186 (N_16186,N_15786,N_15745);
nand U16187 (N_16187,N_15962,N_15624);
nor U16188 (N_16188,N_15682,N_15670);
xor U16189 (N_16189,N_15817,N_15911);
or U16190 (N_16190,N_15762,N_15662);
or U16191 (N_16191,N_15986,N_15766);
or U16192 (N_16192,N_15639,N_15811);
nor U16193 (N_16193,N_15658,N_15914);
nor U16194 (N_16194,N_15608,N_15646);
nor U16195 (N_16195,N_15958,N_15792);
xnor U16196 (N_16196,N_15681,N_15923);
nand U16197 (N_16197,N_15618,N_15649);
xor U16198 (N_16198,N_15953,N_15997);
nor U16199 (N_16199,N_15863,N_15736);
nand U16200 (N_16200,N_15746,N_15614);
and U16201 (N_16201,N_15622,N_15814);
nor U16202 (N_16202,N_15612,N_15762);
and U16203 (N_16203,N_15902,N_15853);
nand U16204 (N_16204,N_15976,N_15973);
or U16205 (N_16205,N_15717,N_15922);
nand U16206 (N_16206,N_15944,N_15681);
xor U16207 (N_16207,N_15872,N_15759);
and U16208 (N_16208,N_15771,N_15694);
or U16209 (N_16209,N_15965,N_15685);
nor U16210 (N_16210,N_15905,N_15626);
or U16211 (N_16211,N_15984,N_15839);
or U16212 (N_16212,N_15789,N_15735);
and U16213 (N_16213,N_15963,N_15736);
nand U16214 (N_16214,N_15605,N_15612);
nor U16215 (N_16215,N_15791,N_15908);
nand U16216 (N_16216,N_15625,N_15644);
nor U16217 (N_16217,N_15775,N_15967);
and U16218 (N_16218,N_15792,N_15787);
nand U16219 (N_16219,N_15632,N_15716);
xnor U16220 (N_16220,N_15888,N_15657);
or U16221 (N_16221,N_15836,N_15685);
xor U16222 (N_16222,N_15807,N_15939);
nand U16223 (N_16223,N_15646,N_15925);
nand U16224 (N_16224,N_15644,N_15971);
nand U16225 (N_16225,N_15700,N_15796);
and U16226 (N_16226,N_15730,N_15750);
nor U16227 (N_16227,N_15616,N_15865);
or U16228 (N_16228,N_15798,N_15794);
nand U16229 (N_16229,N_15852,N_15799);
nor U16230 (N_16230,N_15862,N_15891);
or U16231 (N_16231,N_15828,N_15831);
nor U16232 (N_16232,N_15808,N_15631);
xor U16233 (N_16233,N_15773,N_15714);
nor U16234 (N_16234,N_15889,N_15734);
or U16235 (N_16235,N_15830,N_15973);
nor U16236 (N_16236,N_15889,N_15748);
and U16237 (N_16237,N_15663,N_15907);
and U16238 (N_16238,N_15672,N_15988);
and U16239 (N_16239,N_15881,N_15971);
or U16240 (N_16240,N_15632,N_15835);
and U16241 (N_16241,N_15732,N_15692);
or U16242 (N_16242,N_15898,N_15701);
xor U16243 (N_16243,N_15626,N_15716);
and U16244 (N_16244,N_15997,N_15752);
and U16245 (N_16245,N_15629,N_15720);
or U16246 (N_16246,N_15824,N_15637);
xnor U16247 (N_16247,N_15812,N_15865);
and U16248 (N_16248,N_15776,N_15980);
and U16249 (N_16249,N_15620,N_15688);
xor U16250 (N_16250,N_15812,N_15783);
xor U16251 (N_16251,N_15938,N_15719);
and U16252 (N_16252,N_15914,N_15768);
nor U16253 (N_16253,N_15811,N_15766);
xnor U16254 (N_16254,N_15904,N_15773);
or U16255 (N_16255,N_15663,N_15927);
and U16256 (N_16256,N_15947,N_15690);
nor U16257 (N_16257,N_15619,N_15825);
nor U16258 (N_16258,N_15644,N_15735);
and U16259 (N_16259,N_15905,N_15851);
or U16260 (N_16260,N_15698,N_15762);
and U16261 (N_16261,N_15831,N_15731);
xor U16262 (N_16262,N_15698,N_15729);
nand U16263 (N_16263,N_15897,N_15735);
nor U16264 (N_16264,N_15632,N_15670);
or U16265 (N_16265,N_15829,N_15686);
nand U16266 (N_16266,N_15764,N_15976);
nand U16267 (N_16267,N_15770,N_15962);
xnor U16268 (N_16268,N_15785,N_15731);
nor U16269 (N_16269,N_15882,N_15629);
xor U16270 (N_16270,N_15758,N_15824);
nand U16271 (N_16271,N_15674,N_15721);
and U16272 (N_16272,N_15844,N_15616);
nor U16273 (N_16273,N_15920,N_15656);
xnor U16274 (N_16274,N_15637,N_15967);
nor U16275 (N_16275,N_15859,N_15697);
nand U16276 (N_16276,N_15636,N_15984);
and U16277 (N_16277,N_15625,N_15882);
xor U16278 (N_16278,N_15617,N_15866);
xor U16279 (N_16279,N_15785,N_15660);
nand U16280 (N_16280,N_15773,N_15685);
or U16281 (N_16281,N_15917,N_15992);
or U16282 (N_16282,N_15964,N_15615);
nand U16283 (N_16283,N_15785,N_15927);
nor U16284 (N_16284,N_15777,N_15843);
and U16285 (N_16285,N_15727,N_15626);
and U16286 (N_16286,N_15832,N_15850);
or U16287 (N_16287,N_15679,N_15841);
nand U16288 (N_16288,N_15781,N_15782);
nand U16289 (N_16289,N_15636,N_15678);
or U16290 (N_16290,N_15689,N_15956);
nor U16291 (N_16291,N_15631,N_15990);
nor U16292 (N_16292,N_15846,N_15829);
nand U16293 (N_16293,N_15959,N_15752);
xor U16294 (N_16294,N_15923,N_15754);
nand U16295 (N_16295,N_15651,N_15657);
and U16296 (N_16296,N_15664,N_15750);
or U16297 (N_16297,N_15993,N_15844);
or U16298 (N_16298,N_15783,N_15907);
nand U16299 (N_16299,N_15742,N_15709);
xnor U16300 (N_16300,N_15977,N_15790);
and U16301 (N_16301,N_15978,N_15926);
and U16302 (N_16302,N_15869,N_15905);
and U16303 (N_16303,N_15795,N_15863);
or U16304 (N_16304,N_15916,N_15984);
and U16305 (N_16305,N_15813,N_15720);
xnor U16306 (N_16306,N_15842,N_15947);
xor U16307 (N_16307,N_15929,N_15716);
or U16308 (N_16308,N_15898,N_15635);
and U16309 (N_16309,N_15950,N_15647);
nand U16310 (N_16310,N_15882,N_15926);
xor U16311 (N_16311,N_15722,N_15692);
nand U16312 (N_16312,N_15909,N_15662);
or U16313 (N_16313,N_15865,N_15666);
or U16314 (N_16314,N_15657,N_15904);
nor U16315 (N_16315,N_15783,N_15940);
xor U16316 (N_16316,N_15813,N_15788);
nor U16317 (N_16317,N_15680,N_15789);
nor U16318 (N_16318,N_15793,N_15613);
nor U16319 (N_16319,N_15948,N_15989);
and U16320 (N_16320,N_15890,N_15906);
and U16321 (N_16321,N_15756,N_15734);
or U16322 (N_16322,N_15777,N_15756);
and U16323 (N_16323,N_15612,N_15911);
or U16324 (N_16324,N_15964,N_15781);
and U16325 (N_16325,N_15697,N_15640);
nand U16326 (N_16326,N_15766,N_15974);
or U16327 (N_16327,N_15919,N_15854);
nand U16328 (N_16328,N_15923,N_15793);
or U16329 (N_16329,N_15788,N_15714);
or U16330 (N_16330,N_15960,N_15671);
or U16331 (N_16331,N_15870,N_15671);
and U16332 (N_16332,N_15847,N_15625);
nor U16333 (N_16333,N_15848,N_15646);
nor U16334 (N_16334,N_15637,N_15908);
xor U16335 (N_16335,N_15900,N_15763);
nor U16336 (N_16336,N_15607,N_15817);
and U16337 (N_16337,N_15734,N_15785);
xnor U16338 (N_16338,N_15821,N_15994);
nor U16339 (N_16339,N_15701,N_15941);
or U16340 (N_16340,N_15991,N_15933);
xnor U16341 (N_16341,N_15682,N_15664);
and U16342 (N_16342,N_15709,N_15963);
or U16343 (N_16343,N_15843,N_15678);
xor U16344 (N_16344,N_15928,N_15676);
nor U16345 (N_16345,N_15947,N_15983);
or U16346 (N_16346,N_15920,N_15826);
xnor U16347 (N_16347,N_15739,N_15877);
nand U16348 (N_16348,N_15746,N_15747);
or U16349 (N_16349,N_15881,N_15638);
nand U16350 (N_16350,N_15864,N_15614);
nor U16351 (N_16351,N_15661,N_15699);
xor U16352 (N_16352,N_15908,N_15846);
nor U16353 (N_16353,N_15895,N_15645);
nor U16354 (N_16354,N_15768,N_15747);
nand U16355 (N_16355,N_15824,N_15840);
or U16356 (N_16356,N_15659,N_15851);
and U16357 (N_16357,N_15847,N_15766);
nand U16358 (N_16358,N_15842,N_15620);
nand U16359 (N_16359,N_15808,N_15918);
nand U16360 (N_16360,N_15877,N_15909);
nor U16361 (N_16361,N_15642,N_15657);
nor U16362 (N_16362,N_15665,N_15945);
nor U16363 (N_16363,N_15671,N_15766);
and U16364 (N_16364,N_15829,N_15852);
nand U16365 (N_16365,N_15830,N_15907);
nand U16366 (N_16366,N_15646,N_15834);
or U16367 (N_16367,N_15625,N_15693);
and U16368 (N_16368,N_15656,N_15714);
nand U16369 (N_16369,N_15835,N_15815);
or U16370 (N_16370,N_15686,N_15665);
xnor U16371 (N_16371,N_15933,N_15853);
nand U16372 (N_16372,N_15988,N_15667);
xor U16373 (N_16373,N_15624,N_15692);
xnor U16374 (N_16374,N_15783,N_15808);
nor U16375 (N_16375,N_15665,N_15873);
nand U16376 (N_16376,N_15986,N_15755);
xnor U16377 (N_16377,N_15852,N_15762);
nand U16378 (N_16378,N_15668,N_15953);
nand U16379 (N_16379,N_15832,N_15848);
and U16380 (N_16380,N_15776,N_15616);
nand U16381 (N_16381,N_15763,N_15913);
or U16382 (N_16382,N_15768,N_15994);
and U16383 (N_16383,N_15658,N_15758);
and U16384 (N_16384,N_15664,N_15644);
or U16385 (N_16385,N_15734,N_15945);
nand U16386 (N_16386,N_15715,N_15781);
xnor U16387 (N_16387,N_15978,N_15707);
nand U16388 (N_16388,N_15913,N_15852);
xor U16389 (N_16389,N_15657,N_15971);
and U16390 (N_16390,N_15918,N_15747);
or U16391 (N_16391,N_15905,N_15855);
xnor U16392 (N_16392,N_15881,N_15647);
nor U16393 (N_16393,N_15969,N_15673);
nand U16394 (N_16394,N_15866,N_15732);
nor U16395 (N_16395,N_15798,N_15669);
or U16396 (N_16396,N_15905,N_15748);
xnor U16397 (N_16397,N_15802,N_15927);
and U16398 (N_16398,N_15953,N_15931);
nand U16399 (N_16399,N_15739,N_15771);
and U16400 (N_16400,N_16391,N_16096);
nor U16401 (N_16401,N_16145,N_16061);
nand U16402 (N_16402,N_16095,N_16223);
or U16403 (N_16403,N_16029,N_16250);
nor U16404 (N_16404,N_16293,N_16330);
or U16405 (N_16405,N_16378,N_16278);
xor U16406 (N_16406,N_16085,N_16317);
or U16407 (N_16407,N_16141,N_16217);
and U16408 (N_16408,N_16148,N_16060);
and U16409 (N_16409,N_16197,N_16111);
nand U16410 (N_16410,N_16078,N_16183);
or U16411 (N_16411,N_16295,N_16094);
or U16412 (N_16412,N_16261,N_16017);
nor U16413 (N_16413,N_16064,N_16069);
or U16414 (N_16414,N_16336,N_16304);
nand U16415 (N_16415,N_16359,N_16132);
nor U16416 (N_16416,N_16354,N_16025);
nand U16417 (N_16417,N_16097,N_16311);
and U16418 (N_16418,N_16142,N_16288);
and U16419 (N_16419,N_16159,N_16030);
and U16420 (N_16420,N_16086,N_16074);
xnor U16421 (N_16421,N_16027,N_16325);
or U16422 (N_16422,N_16289,N_16101);
nand U16423 (N_16423,N_16053,N_16249);
or U16424 (N_16424,N_16081,N_16001);
nand U16425 (N_16425,N_16372,N_16076);
or U16426 (N_16426,N_16343,N_16012);
and U16427 (N_16427,N_16389,N_16260);
nor U16428 (N_16428,N_16328,N_16283);
and U16429 (N_16429,N_16088,N_16107);
nor U16430 (N_16430,N_16298,N_16157);
nand U16431 (N_16431,N_16005,N_16356);
or U16432 (N_16432,N_16167,N_16349);
nand U16433 (N_16433,N_16015,N_16386);
or U16434 (N_16434,N_16114,N_16385);
nand U16435 (N_16435,N_16266,N_16133);
and U16436 (N_16436,N_16307,N_16160);
nand U16437 (N_16437,N_16302,N_16301);
or U16438 (N_16438,N_16251,N_16264);
nand U16439 (N_16439,N_16263,N_16327);
xnor U16440 (N_16440,N_16171,N_16051);
or U16441 (N_16441,N_16320,N_16040);
nand U16442 (N_16442,N_16208,N_16033);
and U16443 (N_16443,N_16065,N_16286);
nand U16444 (N_16444,N_16109,N_16257);
nor U16445 (N_16445,N_16398,N_16357);
and U16446 (N_16446,N_16241,N_16070);
or U16447 (N_16447,N_16315,N_16043);
or U16448 (N_16448,N_16122,N_16276);
and U16449 (N_16449,N_16265,N_16262);
nand U16450 (N_16450,N_16049,N_16098);
nor U16451 (N_16451,N_16310,N_16351);
or U16452 (N_16452,N_16185,N_16082);
nor U16453 (N_16453,N_16077,N_16207);
and U16454 (N_16454,N_16150,N_16104);
xor U16455 (N_16455,N_16396,N_16180);
nor U16456 (N_16456,N_16300,N_16013);
and U16457 (N_16457,N_16034,N_16370);
xnor U16458 (N_16458,N_16243,N_16100);
nand U16459 (N_16459,N_16192,N_16238);
nor U16460 (N_16460,N_16369,N_16007);
nand U16461 (N_16461,N_16387,N_16376);
and U16462 (N_16462,N_16189,N_16239);
and U16463 (N_16463,N_16232,N_16340);
and U16464 (N_16464,N_16269,N_16038);
and U16465 (N_16465,N_16139,N_16121);
or U16466 (N_16466,N_16216,N_16173);
nand U16467 (N_16467,N_16113,N_16028);
nand U16468 (N_16468,N_16196,N_16259);
xnor U16469 (N_16469,N_16136,N_16014);
and U16470 (N_16470,N_16321,N_16165);
xor U16471 (N_16471,N_16072,N_16155);
and U16472 (N_16472,N_16003,N_16089);
xnor U16473 (N_16473,N_16240,N_16031);
or U16474 (N_16474,N_16147,N_16346);
xor U16475 (N_16475,N_16390,N_16123);
and U16476 (N_16476,N_16274,N_16258);
nand U16477 (N_16477,N_16292,N_16270);
or U16478 (N_16478,N_16297,N_16119);
nor U16479 (N_16479,N_16339,N_16368);
nand U16480 (N_16480,N_16345,N_16394);
nand U16481 (N_16481,N_16050,N_16073);
and U16482 (N_16482,N_16191,N_16329);
xnor U16483 (N_16483,N_16229,N_16154);
or U16484 (N_16484,N_16395,N_16365);
nor U16485 (N_16485,N_16242,N_16044);
nand U16486 (N_16486,N_16209,N_16153);
nor U16487 (N_16487,N_16335,N_16367);
nand U16488 (N_16488,N_16084,N_16203);
and U16489 (N_16489,N_16056,N_16117);
nand U16490 (N_16490,N_16275,N_16202);
nor U16491 (N_16491,N_16152,N_16120);
nand U16492 (N_16492,N_16041,N_16322);
and U16493 (N_16493,N_16268,N_16093);
xor U16494 (N_16494,N_16380,N_16331);
xnor U16495 (N_16495,N_16057,N_16226);
nor U16496 (N_16496,N_16308,N_16182);
nor U16497 (N_16497,N_16219,N_16112);
nor U16498 (N_16498,N_16256,N_16245);
xnor U16499 (N_16499,N_16174,N_16316);
nor U16500 (N_16500,N_16127,N_16023);
xnor U16501 (N_16501,N_16246,N_16285);
nand U16502 (N_16502,N_16392,N_16248);
and U16503 (N_16503,N_16233,N_16348);
and U16504 (N_16504,N_16211,N_16035);
xnor U16505 (N_16505,N_16149,N_16252);
nor U16506 (N_16506,N_16143,N_16080);
nor U16507 (N_16507,N_16254,N_16324);
nor U16508 (N_16508,N_16313,N_16342);
nand U16509 (N_16509,N_16210,N_16366);
or U16510 (N_16510,N_16178,N_16135);
and U16511 (N_16511,N_16032,N_16287);
and U16512 (N_16512,N_16186,N_16099);
nor U16513 (N_16513,N_16362,N_16230);
xnor U16514 (N_16514,N_16164,N_16021);
nand U16515 (N_16515,N_16039,N_16375);
nor U16516 (N_16516,N_16272,N_16071);
nand U16517 (N_16517,N_16079,N_16175);
and U16518 (N_16518,N_16338,N_16019);
or U16519 (N_16519,N_16234,N_16237);
or U16520 (N_16520,N_16036,N_16194);
and U16521 (N_16521,N_16103,N_16090);
xor U16522 (N_16522,N_16170,N_16009);
xor U16523 (N_16523,N_16002,N_16004);
nand U16524 (N_16524,N_16000,N_16224);
nand U16525 (N_16525,N_16062,N_16187);
or U16526 (N_16526,N_16228,N_16280);
and U16527 (N_16527,N_16220,N_16008);
nand U16528 (N_16528,N_16309,N_16253);
nor U16529 (N_16529,N_16225,N_16190);
nor U16530 (N_16530,N_16358,N_16018);
or U16531 (N_16531,N_16299,N_16231);
and U16532 (N_16532,N_16255,N_16212);
xor U16533 (N_16533,N_16350,N_16334);
nor U16534 (N_16534,N_16199,N_16054);
and U16535 (N_16535,N_16277,N_16124);
xnor U16536 (N_16536,N_16290,N_16052);
and U16537 (N_16537,N_16010,N_16393);
or U16538 (N_16538,N_16016,N_16129);
and U16539 (N_16539,N_16116,N_16046);
and U16540 (N_16540,N_16227,N_16205);
xor U16541 (N_16541,N_16172,N_16323);
xor U16542 (N_16542,N_16303,N_16218);
nor U16543 (N_16543,N_16193,N_16213);
xor U16544 (N_16544,N_16091,N_16244);
nor U16545 (N_16545,N_16115,N_16195);
nand U16546 (N_16546,N_16382,N_16279);
and U16547 (N_16547,N_16326,N_16271);
or U16548 (N_16548,N_16130,N_16314);
nor U16549 (N_16549,N_16222,N_16045);
nand U16550 (N_16550,N_16221,N_16024);
or U16551 (N_16551,N_16318,N_16355);
or U16552 (N_16552,N_16118,N_16305);
or U16553 (N_16553,N_16188,N_16134);
xor U16554 (N_16554,N_16083,N_16011);
or U16555 (N_16555,N_16361,N_16381);
xor U16556 (N_16556,N_16063,N_16176);
and U16557 (N_16557,N_16377,N_16281);
nand U16558 (N_16558,N_16105,N_16181);
xor U16559 (N_16559,N_16306,N_16158);
or U16560 (N_16560,N_16151,N_16291);
xnor U16561 (N_16561,N_16022,N_16179);
xnor U16562 (N_16562,N_16200,N_16384);
and U16563 (N_16563,N_16102,N_16282);
xnor U16564 (N_16564,N_16144,N_16296);
nor U16565 (N_16565,N_16047,N_16273);
nand U16566 (N_16566,N_16379,N_16201);
and U16567 (N_16567,N_16374,N_16371);
xnor U16568 (N_16568,N_16198,N_16138);
xnor U16569 (N_16569,N_16332,N_16075);
nand U16570 (N_16570,N_16110,N_16177);
nand U16571 (N_16571,N_16204,N_16140);
nand U16572 (N_16572,N_16068,N_16399);
and U16573 (N_16573,N_16347,N_16363);
nand U16574 (N_16574,N_16388,N_16284);
nand U16575 (N_16575,N_16206,N_16126);
and U16576 (N_16576,N_16184,N_16236);
xnor U16577 (N_16577,N_16026,N_16383);
or U16578 (N_16578,N_16214,N_16048);
nor U16579 (N_16579,N_16364,N_16235);
nor U16580 (N_16580,N_16169,N_16337);
nor U16581 (N_16581,N_16067,N_16163);
nor U16582 (N_16582,N_16058,N_16333);
xnor U16583 (N_16583,N_16215,N_16042);
and U16584 (N_16584,N_16020,N_16106);
and U16585 (N_16585,N_16294,N_16344);
or U16586 (N_16586,N_16373,N_16267);
or U16587 (N_16587,N_16352,N_16006);
nor U16588 (N_16588,N_16166,N_16360);
nor U16589 (N_16589,N_16156,N_16125);
and U16590 (N_16590,N_16092,N_16353);
and U16591 (N_16591,N_16037,N_16087);
xor U16592 (N_16592,N_16397,N_16137);
nor U16593 (N_16593,N_16108,N_16312);
xnor U16594 (N_16594,N_16146,N_16247);
nor U16595 (N_16595,N_16168,N_16162);
and U16596 (N_16596,N_16066,N_16055);
xnor U16597 (N_16597,N_16128,N_16161);
nor U16598 (N_16598,N_16341,N_16131);
nor U16599 (N_16599,N_16319,N_16059);
or U16600 (N_16600,N_16326,N_16071);
and U16601 (N_16601,N_16373,N_16279);
xor U16602 (N_16602,N_16326,N_16315);
xnor U16603 (N_16603,N_16370,N_16248);
nor U16604 (N_16604,N_16054,N_16310);
xnor U16605 (N_16605,N_16193,N_16330);
and U16606 (N_16606,N_16049,N_16181);
nand U16607 (N_16607,N_16106,N_16292);
and U16608 (N_16608,N_16387,N_16386);
xnor U16609 (N_16609,N_16379,N_16364);
and U16610 (N_16610,N_16086,N_16264);
nand U16611 (N_16611,N_16058,N_16343);
xor U16612 (N_16612,N_16070,N_16292);
xnor U16613 (N_16613,N_16067,N_16244);
and U16614 (N_16614,N_16231,N_16328);
nand U16615 (N_16615,N_16165,N_16352);
or U16616 (N_16616,N_16161,N_16120);
xor U16617 (N_16617,N_16249,N_16380);
nor U16618 (N_16618,N_16212,N_16357);
nor U16619 (N_16619,N_16060,N_16278);
xnor U16620 (N_16620,N_16112,N_16232);
xnor U16621 (N_16621,N_16131,N_16325);
xor U16622 (N_16622,N_16263,N_16158);
and U16623 (N_16623,N_16178,N_16234);
or U16624 (N_16624,N_16099,N_16152);
or U16625 (N_16625,N_16018,N_16163);
and U16626 (N_16626,N_16157,N_16192);
nor U16627 (N_16627,N_16286,N_16290);
xnor U16628 (N_16628,N_16029,N_16142);
nor U16629 (N_16629,N_16351,N_16289);
nor U16630 (N_16630,N_16081,N_16353);
and U16631 (N_16631,N_16058,N_16254);
or U16632 (N_16632,N_16003,N_16391);
nor U16633 (N_16633,N_16173,N_16128);
xnor U16634 (N_16634,N_16294,N_16123);
or U16635 (N_16635,N_16087,N_16277);
and U16636 (N_16636,N_16072,N_16075);
and U16637 (N_16637,N_16292,N_16122);
and U16638 (N_16638,N_16064,N_16349);
nand U16639 (N_16639,N_16181,N_16250);
nor U16640 (N_16640,N_16290,N_16345);
nor U16641 (N_16641,N_16144,N_16353);
and U16642 (N_16642,N_16089,N_16365);
xnor U16643 (N_16643,N_16241,N_16289);
and U16644 (N_16644,N_16188,N_16233);
nor U16645 (N_16645,N_16120,N_16150);
or U16646 (N_16646,N_16058,N_16050);
xnor U16647 (N_16647,N_16048,N_16372);
nand U16648 (N_16648,N_16283,N_16288);
xor U16649 (N_16649,N_16050,N_16002);
xnor U16650 (N_16650,N_16291,N_16196);
nor U16651 (N_16651,N_16294,N_16032);
and U16652 (N_16652,N_16073,N_16065);
xor U16653 (N_16653,N_16087,N_16269);
xnor U16654 (N_16654,N_16199,N_16125);
and U16655 (N_16655,N_16274,N_16186);
nand U16656 (N_16656,N_16304,N_16175);
nand U16657 (N_16657,N_16129,N_16125);
nor U16658 (N_16658,N_16001,N_16029);
xor U16659 (N_16659,N_16344,N_16365);
nor U16660 (N_16660,N_16375,N_16234);
nand U16661 (N_16661,N_16055,N_16354);
or U16662 (N_16662,N_16344,N_16041);
nor U16663 (N_16663,N_16315,N_16200);
xnor U16664 (N_16664,N_16057,N_16341);
nor U16665 (N_16665,N_16186,N_16258);
or U16666 (N_16666,N_16361,N_16355);
nor U16667 (N_16667,N_16016,N_16288);
nor U16668 (N_16668,N_16054,N_16168);
and U16669 (N_16669,N_16015,N_16276);
nand U16670 (N_16670,N_16298,N_16022);
nand U16671 (N_16671,N_16055,N_16314);
and U16672 (N_16672,N_16232,N_16386);
or U16673 (N_16673,N_16033,N_16023);
nand U16674 (N_16674,N_16020,N_16350);
and U16675 (N_16675,N_16109,N_16188);
nand U16676 (N_16676,N_16023,N_16389);
and U16677 (N_16677,N_16096,N_16041);
and U16678 (N_16678,N_16213,N_16019);
and U16679 (N_16679,N_16358,N_16319);
and U16680 (N_16680,N_16390,N_16037);
xor U16681 (N_16681,N_16217,N_16238);
or U16682 (N_16682,N_16303,N_16070);
nor U16683 (N_16683,N_16359,N_16157);
nor U16684 (N_16684,N_16307,N_16102);
or U16685 (N_16685,N_16180,N_16051);
and U16686 (N_16686,N_16183,N_16367);
xnor U16687 (N_16687,N_16055,N_16316);
nand U16688 (N_16688,N_16331,N_16072);
or U16689 (N_16689,N_16005,N_16207);
xor U16690 (N_16690,N_16208,N_16097);
nand U16691 (N_16691,N_16308,N_16213);
and U16692 (N_16692,N_16375,N_16047);
nor U16693 (N_16693,N_16025,N_16377);
nor U16694 (N_16694,N_16348,N_16341);
xnor U16695 (N_16695,N_16141,N_16176);
and U16696 (N_16696,N_16272,N_16372);
nand U16697 (N_16697,N_16256,N_16020);
and U16698 (N_16698,N_16076,N_16094);
nor U16699 (N_16699,N_16036,N_16065);
nand U16700 (N_16700,N_16288,N_16073);
nand U16701 (N_16701,N_16348,N_16358);
nor U16702 (N_16702,N_16094,N_16234);
and U16703 (N_16703,N_16119,N_16290);
and U16704 (N_16704,N_16302,N_16239);
xor U16705 (N_16705,N_16234,N_16192);
and U16706 (N_16706,N_16243,N_16015);
xor U16707 (N_16707,N_16399,N_16388);
nand U16708 (N_16708,N_16362,N_16223);
nor U16709 (N_16709,N_16040,N_16210);
nor U16710 (N_16710,N_16103,N_16387);
or U16711 (N_16711,N_16322,N_16131);
or U16712 (N_16712,N_16055,N_16154);
nor U16713 (N_16713,N_16201,N_16057);
nand U16714 (N_16714,N_16369,N_16203);
and U16715 (N_16715,N_16397,N_16105);
xnor U16716 (N_16716,N_16113,N_16030);
xor U16717 (N_16717,N_16310,N_16302);
nor U16718 (N_16718,N_16258,N_16088);
or U16719 (N_16719,N_16120,N_16128);
nand U16720 (N_16720,N_16269,N_16213);
nor U16721 (N_16721,N_16319,N_16148);
and U16722 (N_16722,N_16372,N_16119);
nor U16723 (N_16723,N_16087,N_16263);
nor U16724 (N_16724,N_16006,N_16365);
xor U16725 (N_16725,N_16064,N_16366);
and U16726 (N_16726,N_16088,N_16195);
nand U16727 (N_16727,N_16268,N_16296);
and U16728 (N_16728,N_16189,N_16234);
nand U16729 (N_16729,N_16044,N_16311);
and U16730 (N_16730,N_16308,N_16176);
xnor U16731 (N_16731,N_16198,N_16158);
and U16732 (N_16732,N_16362,N_16192);
nor U16733 (N_16733,N_16346,N_16396);
and U16734 (N_16734,N_16237,N_16223);
nand U16735 (N_16735,N_16040,N_16041);
xor U16736 (N_16736,N_16000,N_16132);
or U16737 (N_16737,N_16008,N_16056);
xnor U16738 (N_16738,N_16007,N_16254);
nand U16739 (N_16739,N_16024,N_16364);
or U16740 (N_16740,N_16205,N_16212);
nand U16741 (N_16741,N_16325,N_16066);
nor U16742 (N_16742,N_16262,N_16185);
nor U16743 (N_16743,N_16377,N_16296);
or U16744 (N_16744,N_16107,N_16312);
nor U16745 (N_16745,N_16284,N_16145);
xor U16746 (N_16746,N_16146,N_16321);
nand U16747 (N_16747,N_16192,N_16115);
or U16748 (N_16748,N_16265,N_16161);
xor U16749 (N_16749,N_16040,N_16171);
or U16750 (N_16750,N_16383,N_16106);
xnor U16751 (N_16751,N_16171,N_16362);
xnor U16752 (N_16752,N_16002,N_16383);
nor U16753 (N_16753,N_16293,N_16191);
or U16754 (N_16754,N_16094,N_16042);
nand U16755 (N_16755,N_16184,N_16364);
nand U16756 (N_16756,N_16288,N_16352);
or U16757 (N_16757,N_16226,N_16061);
xnor U16758 (N_16758,N_16067,N_16193);
nand U16759 (N_16759,N_16148,N_16137);
nand U16760 (N_16760,N_16216,N_16388);
nand U16761 (N_16761,N_16130,N_16297);
nand U16762 (N_16762,N_16277,N_16154);
or U16763 (N_16763,N_16273,N_16049);
or U16764 (N_16764,N_16078,N_16116);
nor U16765 (N_16765,N_16291,N_16337);
xnor U16766 (N_16766,N_16257,N_16281);
nor U16767 (N_16767,N_16168,N_16182);
xor U16768 (N_16768,N_16283,N_16313);
nor U16769 (N_16769,N_16022,N_16359);
xor U16770 (N_16770,N_16007,N_16049);
and U16771 (N_16771,N_16219,N_16154);
nor U16772 (N_16772,N_16171,N_16367);
nor U16773 (N_16773,N_16176,N_16305);
nand U16774 (N_16774,N_16061,N_16312);
or U16775 (N_16775,N_16033,N_16121);
or U16776 (N_16776,N_16162,N_16192);
nand U16777 (N_16777,N_16022,N_16391);
xnor U16778 (N_16778,N_16382,N_16070);
xnor U16779 (N_16779,N_16391,N_16358);
and U16780 (N_16780,N_16216,N_16314);
nand U16781 (N_16781,N_16165,N_16343);
nand U16782 (N_16782,N_16294,N_16312);
xor U16783 (N_16783,N_16318,N_16033);
and U16784 (N_16784,N_16007,N_16041);
xnor U16785 (N_16785,N_16368,N_16190);
or U16786 (N_16786,N_16079,N_16355);
nor U16787 (N_16787,N_16105,N_16338);
nor U16788 (N_16788,N_16266,N_16094);
or U16789 (N_16789,N_16042,N_16393);
nand U16790 (N_16790,N_16034,N_16317);
and U16791 (N_16791,N_16208,N_16217);
or U16792 (N_16792,N_16022,N_16390);
nand U16793 (N_16793,N_16221,N_16256);
nand U16794 (N_16794,N_16029,N_16192);
and U16795 (N_16795,N_16162,N_16150);
and U16796 (N_16796,N_16300,N_16284);
nor U16797 (N_16797,N_16302,N_16238);
nand U16798 (N_16798,N_16139,N_16277);
nand U16799 (N_16799,N_16170,N_16215);
or U16800 (N_16800,N_16663,N_16793);
nor U16801 (N_16801,N_16408,N_16625);
or U16802 (N_16802,N_16491,N_16533);
and U16803 (N_16803,N_16529,N_16690);
xor U16804 (N_16804,N_16583,N_16574);
nor U16805 (N_16805,N_16613,N_16682);
xor U16806 (N_16806,N_16758,N_16775);
and U16807 (N_16807,N_16748,N_16471);
nor U16808 (N_16808,N_16428,N_16716);
nor U16809 (N_16809,N_16412,N_16524);
or U16810 (N_16810,N_16627,N_16603);
nand U16811 (N_16811,N_16484,N_16451);
xnor U16812 (N_16812,N_16470,N_16591);
xor U16813 (N_16813,N_16735,N_16441);
nand U16814 (N_16814,N_16632,N_16606);
nor U16815 (N_16815,N_16526,N_16521);
nor U16816 (N_16816,N_16499,N_16414);
nor U16817 (N_16817,N_16440,N_16416);
and U16818 (N_16818,N_16502,N_16545);
or U16819 (N_16819,N_16458,N_16723);
xnor U16820 (N_16820,N_16647,N_16679);
nand U16821 (N_16821,N_16559,N_16599);
nand U16822 (N_16822,N_16695,N_16651);
or U16823 (N_16823,N_16799,N_16421);
nand U16824 (N_16824,N_16742,N_16552);
nor U16825 (N_16825,N_16563,N_16797);
nor U16826 (N_16826,N_16721,N_16641);
xor U16827 (N_16827,N_16774,N_16555);
and U16828 (N_16828,N_16717,N_16537);
xnor U16829 (N_16829,N_16406,N_16427);
nand U16830 (N_16830,N_16478,N_16417);
xor U16831 (N_16831,N_16634,N_16560);
nand U16832 (N_16832,N_16546,N_16612);
nor U16833 (N_16833,N_16454,N_16405);
and U16834 (N_16834,N_16622,N_16637);
nor U16835 (N_16835,N_16575,N_16595);
and U16836 (N_16836,N_16419,N_16649);
nand U16837 (N_16837,N_16553,N_16557);
nand U16838 (N_16838,N_16724,N_16746);
nor U16839 (N_16839,N_16718,N_16788);
and U16840 (N_16840,N_16768,N_16794);
or U16841 (N_16841,N_16745,N_16402);
nor U16842 (N_16842,N_16645,N_16755);
or U16843 (N_16843,N_16683,N_16636);
nor U16844 (N_16844,N_16468,N_16436);
and U16845 (N_16845,N_16761,N_16496);
nand U16846 (N_16846,N_16701,N_16586);
xnor U16847 (N_16847,N_16530,N_16507);
and U16848 (N_16848,N_16517,N_16602);
and U16849 (N_16849,N_16539,N_16593);
and U16850 (N_16850,N_16617,N_16462);
xnor U16851 (N_16851,N_16475,N_16660);
xnor U16852 (N_16852,N_16477,N_16518);
or U16853 (N_16853,N_16608,N_16767);
and U16854 (N_16854,N_16509,N_16676);
nand U16855 (N_16855,N_16624,N_16561);
nor U16856 (N_16856,N_16536,N_16661);
xnor U16857 (N_16857,N_16747,N_16469);
or U16858 (N_16858,N_16777,N_16413);
or U16859 (N_16859,N_16776,N_16750);
nand U16860 (N_16860,N_16486,N_16512);
nor U16861 (N_16861,N_16596,N_16658);
xor U16862 (N_16862,N_16435,N_16404);
xnor U16863 (N_16863,N_16752,N_16714);
xor U16864 (N_16864,N_16688,N_16453);
xnor U16865 (N_16865,N_16494,N_16571);
and U16866 (N_16866,N_16704,N_16433);
xnor U16867 (N_16867,N_16578,N_16744);
and U16868 (N_16868,N_16719,N_16525);
or U16869 (N_16869,N_16639,N_16738);
nand U16870 (N_16870,N_16673,N_16543);
nand U16871 (N_16871,N_16439,N_16771);
and U16872 (N_16872,N_16640,N_16769);
nor U16873 (N_16873,N_16527,N_16707);
nor U16874 (N_16874,N_16488,N_16444);
nor U16875 (N_16875,N_16548,N_16653);
xnor U16876 (N_16876,N_16646,N_16756);
nor U16877 (N_16877,N_16443,N_16549);
nand U16878 (N_16878,N_16766,N_16731);
or U16879 (N_16879,N_16664,N_16694);
or U16880 (N_16880,N_16540,N_16538);
nand U16881 (N_16881,N_16696,N_16792);
or U16882 (N_16882,N_16759,N_16722);
and U16883 (N_16883,N_16523,N_16445);
nand U16884 (N_16884,N_16505,N_16698);
nand U16885 (N_16885,N_16515,N_16550);
xor U16886 (N_16886,N_16728,N_16420);
nand U16887 (N_16887,N_16620,N_16449);
or U16888 (N_16888,N_16423,N_16784);
nor U16889 (N_16889,N_16732,N_16588);
nor U16890 (N_16890,N_16567,N_16630);
nor U16891 (N_16891,N_16418,N_16584);
nor U16892 (N_16892,N_16592,N_16710);
nor U16893 (N_16893,N_16554,N_16765);
and U16894 (N_16894,N_16654,N_16411);
and U16895 (N_16895,N_16778,N_16562);
nand U16896 (N_16896,N_16659,N_16466);
nand U16897 (N_16897,N_16482,N_16670);
or U16898 (N_16898,N_16697,N_16626);
or U16899 (N_16899,N_16648,N_16763);
nor U16900 (N_16900,N_16481,N_16501);
or U16901 (N_16901,N_16712,N_16594);
and U16902 (N_16902,N_16590,N_16459);
nand U16903 (N_16903,N_16531,N_16506);
and U16904 (N_16904,N_16407,N_16479);
xnor U16905 (N_16905,N_16424,N_16666);
xnor U16906 (N_16906,N_16770,N_16460);
nand U16907 (N_16907,N_16609,N_16432);
xnor U16908 (N_16908,N_16483,N_16504);
or U16909 (N_16909,N_16587,N_16671);
or U16910 (N_16910,N_16558,N_16655);
nor U16911 (N_16911,N_16422,N_16700);
and U16912 (N_16912,N_16450,N_16564);
xnor U16913 (N_16913,N_16503,N_16669);
nand U16914 (N_16914,N_16410,N_16403);
or U16915 (N_16915,N_16455,N_16572);
or U16916 (N_16916,N_16534,N_16431);
or U16917 (N_16917,N_16643,N_16691);
nand U16918 (N_16918,N_16452,N_16544);
xor U16919 (N_16919,N_16760,N_16490);
nand U16920 (N_16920,N_16522,N_16787);
xor U16921 (N_16921,N_16581,N_16513);
and U16922 (N_16922,N_16429,N_16535);
or U16923 (N_16923,N_16693,N_16614);
nand U16924 (N_16924,N_16657,N_16785);
and U16925 (N_16925,N_16610,N_16569);
nand U16926 (N_16926,N_16448,N_16615);
nand U16927 (N_16927,N_16628,N_16665);
nand U16928 (N_16928,N_16400,N_16743);
xor U16929 (N_16929,N_16631,N_16464);
nand U16930 (N_16930,N_16598,N_16607);
or U16931 (N_16931,N_16685,N_16437);
and U16932 (N_16932,N_16623,N_16740);
nand U16933 (N_16933,N_16430,N_16489);
nand U16934 (N_16934,N_16605,N_16795);
and U16935 (N_16935,N_16751,N_16689);
nor U16936 (N_16936,N_16789,N_16667);
and U16937 (N_16937,N_16638,N_16635);
xor U16938 (N_16938,N_16725,N_16674);
xor U16939 (N_16939,N_16729,N_16668);
xor U16940 (N_16940,N_16467,N_16465);
and U16941 (N_16941,N_16681,N_16772);
nand U16942 (N_16942,N_16741,N_16753);
or U16943 (N_16943,N_16642,N_16487);
xnor U16944 (N_16944,N_16713,N_16532);
nand U16945 (N_16945,N_16456,N_16576);
or U16946 (N_16946,N_16699,N_16680);
or U16947 (N_16947,N_16798,N_16409);
xnor U16948 (N_16948,N_16662,N_16565);
nor U16949 (N_16949,N_16715,N_16425);
and U16950 (N_16950,N_16650,N_16510);
nand U16951 (N_16951,N_16675,N_16446);
and U16952 (N_16952,N_16498,N_16730);
nor U16953 (N_16953,N_16426,N_16500);
xor U16954 (N_16954,N_16519,N_16621);
xor U16955 (N_16955,N_16783,N_16790);
xnor U16956 (N_16956,N_16597,N_16677);
and U16957 (N_16957,N_16585,N_16629);
xnor U16958 (N_16958,N_16791,N_16434);
nand U16959 (N_16959,N_16709,N_16779);
or U16960 (N_16960,N_16516,N_16566);
and U16961 (N_16961,N_16438,N_16705);
xnor U16962 (N_16962,N_16692,N_16514);
nand U16963 (N_16963,N_16582,N_16589);
nand U16964 (N_16964,N_16401,N_16568);
xnor U16965 (N_16965,N_16508,N_16447);
or U16966 (N_16966,N_16736,N_16547);
or U16967 (N_16967,N_16472,N_16442);
xnor U16968 (N_16968,N_16618,N_16457);
and U16969 (N_16969,N_16684,N_16633);
xnor U16970 (N_16970,N_16644,N_16737);
nand U16971 (N_16971,N_16619,N_16687);
and U16972 (N_16972,N_16739,N_16786);
xnor U16973 (N_16973,N_16485,N_16601);
and U16974 (N_16974,N_16656,N_16473);
and U16975 (N_16975,N_16757,N_16497);
xnor U16976 (N_16976,N_16493,N_16480);
or U16977 (N_16977,N_16541,N_16528);
xnor U16978 (N_16978,N_16796,N_16773);
and U16979 (N_16979,N_16542,N_16780);
xnor U16980 (N_16980,N_16754,N_16711);
nor U16981 (N_16981,N_16476,N_16703);
or U16982 (N_16982,N_16611,N_16726);
and U16983 (N_16983,N_16580,N_16733);
and U16984 (N_16984,N_16495,N_16463);
nand U16985 (N_16985,N_16415,N_16762);
and U16986 (N_16986,N_16686,N_16556);
nor U16987 (N_16987,N_16492,N_16672);
and U16988 (N_16988,N_16570,N_16461);
and U16989 (N_16989,N_16474,N_16782);
nand U16990 (N_16990,N_16781,N_16604);
nand U16991 (N_16991,N_16600,N_16579);
and U16992 (N_16992,N_16652,N_16727);
xor U16993 (N_16993,N_16749,N_16734);
nor U16994 (N_16994,N_16678,N_16708);
nand U16995 (N_16995,N_16551,N_16520);
or U16996 (N_16996,N_16577,N_16573);
nand U16997 (N_16997,N_16511,N_16706);
or U16998 (N_16998,N_16616,N_16702);
nor U16999 (N_16999,N_16720,N_16764);
or U17000 (N_17000,N_16480,N_16638);
nand U17001 (N_17001,N_16708,N_16469);
xnor U17002 (N_17002,N_16552,N_16555);
and U17003 (N_17003,N_16547,N_16532);
nand U17004 (N_17004,N_16596,N_16547);
and U17005 (N_17005,N_16446,N_16670);
or U17006 (N_17006,N_16449,N_16645);
and U17007 (N_17007,N_16642,N_16631);
and U17008 (N_17008,N_16608,N_16454);
or U17009 (N_17009,N_16733,N_16637);
or U17010 (N_17010,N_16620,N_16415);
nand U17011 (N_17011,N_16467,N_16785);
xor U17012 (N_17012,N_16410,N_16655);
or U17013 (N_17013,N_16496,N_16455);
nor U17014 (N_17014,N_16728,N_16626);
and U17015 (N_17015,N_16583,N_16785);
nand U17016 (N_17016,N_16730,N_16500);
xor U17017 (N_17017,N_16592,N_16451);
nor U17018 (N_17018,N_16788,N_16424);
nor U17019 (N_17019,N_16770,N_16781);
xnor U17020 (N_17020,N_16439,N_16401);
or U17021 (N_17021,N_16690,N_16512);
nor U17022 (N_17022,N_16589,N_16686);
and U17023 (N_17023,N_16780,N_16531);
xor U17024 (N_17024,N_16493,N_16437);
and U17025 (N_17025,N_16609,N_16611);
or U17026 (N_17026,N_16445,N_16538);
nor U17027 (N_17027,N_16515,N_16607);
or U17028 (N_17028,N_16467,N_16586);
and U17029 (N_17029,N_16762,N_16600);
nand U17030 (N_17030,N_16650,N_16526);
or U17031 (N_17031,N_16599,N_16647);
nor U17032 (N_17032,N_16697,N_16619);
or U17033 (N_17033,N_16759,N_16411);
nand U17034 (N_17034,N_16493,N_16542);
and U17035 (N_17035,N_16672,N_16779);
and U17036 (N_17036,N_16746,N_16562);
nand U17037 (N_17037,N_16659,N_16414);
and U17038 (N_17038,N_16764,N_16760);
nor U17039 (N_17039,N_16707,N_16461);
or U17040 (N_17040,N_16431,N_16784);
nand U17041 (N_17041,N_16544,N_16482);
and U17042 (N_17042,N_16578,N_16724);
xnor U17043 (N_17043,N_16768,N_16481);
and U17044 (N_17044,N_16615,N_16536);
nor U17045 (N_17045,N_16410,N_16483);
nor U17046 (N_17046,N_16486,N_16550);
xor U17047 (N_17047,N_16436,N_16603);
and U17048 (N_17048,N_16512,N_16531);
or U17049 (N_17049,N_16401,N_16532);
or U17050 (N_17050,N_16691,N_16699);
or U17051 (N_17051,N_16695,N_16432);
nor U17052 (N_17052,N_16448,N_16680);
nor U17053 (N_17053,N_16520,N_16438);
and U17054 (N_17054,N_16514,N_16501);
or U17055 (N_17055,N_16453,N_16441);
and U17056 (N_17056,N_16620,N_16569);
xnor U17057 (N_17057,N_16677,N_16433);
and U17058 (N_17058,N_16599,N_16777);
or U17059 (N_17059,N_16410,N_16643);
or U17060 (N_17060,N_16693,N_16483);
or U17061 (N_17061,N_16608,N_16776);
nand U17062 (N_17062,N_16722,N_16590);
nor U17063 (N_17063,N_16798,N_16460);
or U17064 (N_17064,N_16636,N_16428);
nor U17065 (N_17065,N_16438,N_16681);
nand U17066 (N_17066,N_16466,N_16536);
or U17067 (N_17067,N_16447,N_16787);
and U17068 (N_17068,N_16787,N_16746);
nand U17069 (N_17069,N_16594,N_16506);
xnor U17070 (N_17070,N_16556,N_16786);
nand U17071 (N_17071,N_16648,N_16685);
nor U17072 (N_17072,N_16703,N_16707);
or U17073 (N_17073,N_16671,N_16505);
nor U17074 (N_17074,N_16611,N_16705);
nor U17075 (N_17075,N_16756,N_16678);
or U17076 (N_17076,N_16400,N_16697);
or U17077 (N_17077,N_16475,N_16544);
xnor U17078 (N_17078,N_16643,N_16580);
nor U17079 (N_17079,N_16709,N_16449);
nand U17080 (N_17080,N_16495,N_16791);
or U17081 (N_17081,N_16555,N_16726);
nor U17082 (N_17082,N_16456,N_16585);
nand U17083 (N_17083,N_16461,N_16786);
or U17084 (N_17084,N_16610,N_16589);
xnor U17085 (N_17085,N_16529,N_16620);
nor U17086 (N_17086,N_16568,N_16627);
xnor U17087 (N_17087,N_16431,N_16795);
or U17088 (N_17088,N_16743,N_16651);
nand U17089 (N_17089,N_16569,N_16648);
xnor U17090 (N_17090,N_16701,N_16786);
nor U17091 (N_17091,N_16630,N_16459);
or U17092 (N_17092,N_16449,N_16678);
or U17093 (N_17093,N_16443,N_16795);
and U17094 (N_17094,N_16663,N_16693);
and U17095 (N_17095,N_16759,N_16610);
xnor U17096 (N_17096,N_16478,N_16562);
and U17097 (N_17097,N_16746,N_16456);
and U17098 (N_17098,N_16720,N_16510);
nand U17099 (N_17099,N_16562,N_16615);
or U17100 (N_17100,N_16535,N_16423);
or U17101 (N_17101,N_16655,N_16670);
xor U17102 (N_17102,N_16480,N_16647);
xor U17103 (N_17103,N_16524,N_16508);
and U17104 (N_17104,N_16793,N_16474);
xor U17105 (N_17105,N_16607,N_16548);
xor U17106 (N_17106,N_16630,N_16696);
xnor U17107 (N_17107,N_16405,N_16464);
xnor U17108 (N_17108,N_16412,N_16738);
nor U17109 (N_17109,N_16762,N_16700);
xnor U17110 (N_17110,N_16766,N_16424);
xnor U17111 (N_17111,N_16645,N_16611);
nor U17112 (N_17112,N_16784,N_16603);
nand U17113 (N_17113,N_16583,N_16673);
xor U17114 (N_17114,N_16549,N_16649);
or U17115 (N_17115,N_16777,N_16744);
xor U17116 (N_17116,N_16493,N_16643);
xnor U17117 (N_17117,N_16442,N_16445);
and U17118 (N_17118,N_16401,N_16640);
nor U17119 (N_17119,N_16728,N_16665);
xor U17120 (N_17120,N_16754,N_16649);
or U17121 (N_17121,N_16504,N_16578);
or U17122 (N_17122,N_16707,N_16423);
nand U17123 (N_17123,N_16489,N_16687);
xor U17124 (N_17124,N_16582,N_16753);
nand U17125 (N_17125,N_16663,N_16741);
nand U17126 (N_17126,N_16780,N_16485);
and U17127 (N_17127,N_16699,N_16660);
and U17128 (N_17128,N_16520,N_16482);
nand U17129 (N_17129,N_16623,N_16556);
or U17130 (N_17130,N_16708,N_16716);
nand U17131 (N_17131,N_16658,N_16544);
and U17132 (N_17132,N_16482,N_16466);
nand U17133 (N_17133,N_16402,N_16648);
nand U17134 (N_17134,N_16702,N_16754);
and U17135 (N_17135,N_16599,N_16584);
nor U17136 (N_17136,N_16547,N_16659);
or U17137 (N_17137,N_16740,N_16667);
nor U17138 (N_17138,N_16682,N_16596);
xor U17139 (N_17139,N_16472,N_16626);
nand U17140 (N_17140,N_16798,N_16640);
nor U17141 (N_17141,N_16418,N_16523);
nand U17142 (N_17142,N_16776,N_16515);
xor U17143 (N_17143,N_16496,N_16532);
or U17144 (N_17144,N_16610,N_16408);
nor U17145 (N_17145,N_16509,N_16623);
nor U17146 (N_17146,N_16558,N_16704);
nand U17147 (N_17147,N_16703,N_16455);
nor U17148 (N_17148,N_16662,N_16514);
nor U17149 (N_17149,N_16533,N_16772);
nand U17150 (N_17150,N_16767,N_16582);
xnor U17151 (N_17151,N_16415,N_16470);
xor U17152 (N_17152,N_16699,N_16799);
xnor U17153 (N_17153,N_16574,N_16665);
xor U17154 (N_17154,N_16527,N_16717);
xnor U17155 (N_17155,N_16429,N_16580);
nor U17156 (N_17156,N_16539,N_16403);
xnor U17157 (N_17157,N_16609,N_16406);
or U17158 (N_17158,N_16627,N_16601);
nor U17159 (N_17159,N_16632,N_16556);
nor U17160 (N_17160,N_16404,N_16512);
or U17161 (N_17161,N_16686,N_16408);
xor U17162 (N_17162,N_16732,N_16444);
xor U17163 (N_17163,N_16570,N_16660);
xnor U17164 (N_17164,N_16766,N_16503);
nor U17165 (N_17165,N_16672,N_16576);
or U17166 (N_17166,N_16502,N_16588);
nor U17167 (N_17167,N_16497,N_16571);
and U17168 (N_17168,N_16430,N_16761);
nand U17169 (N_17169,N_16689,N_16472);
or U17170 (N_17170,N_16762,N_16742);
and U17171 (N_17171,N_16477,N_16416);
xor U17172 (N_17172,N_16560,N_16515);
nand U17173 (N_17173,N_16404,N_16424);
and U17174 (N_17174,N_16701,N_16789);
nor U17175 (N_17175,N_16418,N_16702);
xor U17176 (N_17176,N_16600,N_16606);
nand U17177 (N_17177,N_16740,N_16508);
and U17178 (N_17178,N_16601,N_16751);
and U17179 (N_17179,N_16560,N_16617);
xor U17180 (N_17180,N_16729,N_16612);
xor U17181 (N_17181,N_16472,N_16755);
and U17182 (N_17182,N_16400,N_16709);
xor U17183 (N_17183,N_16445,N_16491);
and U17184 (N_17184,N_16666,N_16653);
or U17185 (N_17185,N_16698,N_16799);
or U17186 (N_17186,N_16430,N_16741);
nor U17187 (N_17187,N_16506,N_16486);
nand U17188 (N_17188,N_16608,N_16691);
nand U17189 (N_17189,N_16472,N_16650);
nor U17190 (N_17190,N_16607,N_16618);
xnor U17191 (N_17191,N_16747,N_16766);
xor U17192 (N_17192,N_16466,N_16653);
nor U17193 (N_17193,N_16570,N_16704);
xnor U17194 (N_17194,N_16661,N_16671);
nor U17195 (N_17195,N_16668,N_16741);
nor U17196 (N_17196,N_16552,N_16743);
or U17197 (N_17197,N_16576,N_16405);
nand U17198 (N_17198,N_16755,N_16736);
or U17199 (N_17199,N_16402,N_16431);
or U17200 (N_17200,N_16901,N_16882);
and U17201 (N_17201,N_17119,N_16812);
nand U17202 (N_17202,N_16919,N_16878);
or U17203 (N_17203,N_17049,N_17128);
or U17204 (N_17204,N_16840,N_17120);
xnor U17205 (N_17205,N_16941,N_16921);
or U17206 (N_17206,N_16881,N_17004);
and U17207 (N_17207,N_16996,N_17000);
xnor U17208 (N_17208,N_16802,N_16999);
nand U17209 (N_17209,N_17032,N_16864);
xnor U17210 (N_17210,N_17159,N_17152);
xnor U17211 (N_17211,N_16819,N_17001);
xor U17212 (N_17212,N_17192,N_17015);
or U17213 (N_17213,N_16994,N_16857);
xor U17214 (N_17214,N_16816,N_16839);
nor U17215 (N_17215,N_16833,N_16905);
xnor U17216 (N_17216,N_16981,N_17053);
and U17217 (N_17217,N_17117,N_16866);
nor U17218 (N_17218,N_17023,N_17027);
nand U17219 (N_17219,N_17174,N_17002);
xor U17220 (N_17220,N_17167,N_16873);
nand U17221 (N_17221,N_17103,N_17022);
or U17222 (N_17222,N_17112,N_16897);
nand U17223 (N_17223,N_17131,N_16960);
or U17224 (N_17224,N_16966,N_17104);
and U17225 (N_17225,N_16975,N_16877);
xnor U17226 (N_17226,N_17020,N_17029);
or U17227 (N_17227,N_17074,N_16929);
nand U17228 (N_17228,N_17101,N_17130);
xnor U17229 (N_17229,N_16829,N_16846);
nand U17230 (N_17230,N_17005,N_16931);
and U17231 (N_17231,N_16800,N_17180);
xor U17232 (N_17232,N_17081,N_17045);
xnor U17233 (N_17233,N_17150,N_16952);
or U17234 (N_17234,N_16945,N_16969);
xnor U17235 (N_17235,N_17105,N_16880);
nand U17236 (N_17236,N_16944,N_16888);
xor U17237 (N_17237,N_16847,N_16814);
nor U17238 (N_17238,N_17118,N_16834);
and U17239 (N_17239,N_16976,N_17108);
nand U17240 (N_17240,N_16923,N_17144);
and U17241 (N_17241,N_17151,N_16946);
nand U17242 (N_17242,N_16957,N_17037);
and U17243 (N_17243,N_17197,N_17087);
nor U17244 (N_17244,N_17088,N_16920);
or U17245 (N_17245,N_16815,N_16998);
nor U17246 (N_17246,N_16886,N_17082);
nor U17247 (N_17247,N_16980,N_17134);
nand U17248 (N_17248,N_17086,N_17161);
or U17249 (N_17249,N_16841,N_16933);
nand U17250 (N_17250,N_17066,N_16821);
xor U17251 (N_17251,N_17048,N_17011);
nand U17252 (N_17252,N_16871,N_17107);
or U17253 (N_17253,N_17021,N_16965);
nor U17254 (N_17254,N_16836,N_16979);
nor U17255 (N_17255,N_16989,N_16934);
xor U17256 (N_17256,N_16926,N_16948);
nand U17257 (N_17257,N_16907,N_16982);
or U17258 (N_17258,N_16854,N_17041);
nand U17259 (N_17259,N_16902,N_16959);
or U17260 (N_17260,N_17162,N_17019);
nand U17261 (N_17261,N_16826,N_17196);
or U17262 (N_17262,N_16937,N_17052);
and U17263 (N_17263,N_17025,N_17127);
xor U17264 (N_17264,N_16867,N_16911);
or U17265 (N_17265,N_17132,N_17098);
nor U17266 (N_17266,N_16968,N_17110);
nand U17267 (N_17267,N_16848,N_17016);
or U17268 (N_17268,N_16887,N_17126);
or U17269 (N_17269,N_16987,N_17044);
nand U17270 (N_17270,N_17036,N_16884);
or U17271 (N_17271,N_17047,N_17010);
nand U17272 (N_17272,N_17040,N_16862);
or U17273 (N_17273,N_17146,N_17125);
nor U17274 (N_17274,N_17035,N_17133);
xor U17275 (N_17275,N_16828,N_16870);
nor U17276 (N_17276,N_17075,N_17172);
and U17277 (N_17277,N_16983,N_17184);
xor U17278 (N_17278,N_16851,N_16947);
or U17279 (N_17279,N_17168,N_16874);
xor U17280 (N_17280,N_17073,N_17008);
and U17281 (N_17281,N_16868,N_16804);
nand U17282 (N_17282,N_17195,N_17080);
xnor U17283 (N_17283,N_17154,N_17064);
and U17284 (N_17284,N_16974,N_17137);
and U17285 (N_17285,N_16938,N_16883);
nand U17286 (N_17286,N_17177,N_16973);
nor U17287 (N_17287,N_16942,N_16962);
nand U17288 (N_17288,N_16894,N_16986);
and U17289 (N_17289,N_17089,N_17099);
xnor U17290 (N_17290,N_17114,N_17153);
xor U17291 (N_17291,N_17149,N_17057);
or U17292 (N_17292,N_16809,N_17078);
and U17293 (N_17293,N_17123,N_17182);
nor U17294 (N_17294,N_16838,N_16845);
nor U17295 (N_17295,N_16978,N_17141);
nor U17296 (N_17296,N_17175,N_16956);
nand U17297 (N_17297,N_16849,N_17111);
xnor U17298 (N_17298,N_17046,N_17030);
and U17299 (N_17299,N_17007,N_17033);
nor U17300 (N_17300,N_16817,N_17042);
nand U17301 (N_17301,N_17116,N_16990);
nor U17302 (N_17302,N_17124,N_16936);
nand U17303 (N_17303,N_16955,N_17090);
nand U17304 (N_17304,N_16916,N_17173);
or U17305 (N_17305,N_17155,N_17163);
and U17306 (N_17306,N_17062,N_17018);
and U17307 (N_17307,N_17138,N_17060);
and U17308 (N_17308,N_16820,N_16925);
and U17309 (N_17309,N_16991,N_17135);
or U17310 (N_17310,N_16806,N_16900);
nand U17311 (N_17311,N_17079,N_16885);
nand U17312 (N_17312,N_16895,N_16927);
nor U17313 (N_17313,N_16801,N_16964);
nor U17314 (N_17314,N_16899,N_17013);
nand U17315 (N_17315,N_16837,N_16805);
or U17316 (N_17316,N_17147,N_17024);
nand U17317 (N_17317,N_16813,N_16958);
xnor U17318 (N_17318,N_16872,N_17058);
and U17319 (N_17319,N_16928,N_16924);
nor U17320 (N_17320,N_17003,N_17059);
or U17321 (N_17321,N_16997,N_17109);
or U17322 (N_17322,N_16825,N_16904);
xnor U17323 (N_17323,N_16930,N_17193);
xnor U17324 (N_17324,N_16909,N_16984);
xor U17325 (N_17325,N_16935,N_17158);
xor U17326 (N_17326,N_17092,N_17014);
or U17327 (N_17327,N_17102,N_16988);
xor U17328 (N_17328,N_16843,N_16860);
nand U17329 (N_17329,N_16865,N_17054);
or U17330 (N_17330,N_16912,N_17106);
or U17331 (N_17331,N_17160,N_17050);
nand U17332 (N_17332,N_16852,N_16939);
nor U17333 (N_17333,N_17148,N_17113);
xor U17334 (N_17334,N_17100,N_17121);
xor U17335 (N_17335,N_16835,N_17039);
and U17336 (N_17336,N_16971,N_16844);
or U17337 (N_17337,N_17095,N_17143);
and U17338 (N_17338,N_16914,N_16967);
xor U17339 (N_17339,N_16808,N_17028);
nor U17340 (N_17340,N_16915,N_17009);
nand U17341 (N_17341,N_17188,N_16879);
and U17342 (N_17342,N_16993,N_17077);
or U17343 (N_17343,N_16977,N_17140);
and U17344 (N_17344,N_17051,N_17094);
or U17345 (N_17345,N_17115,N_16869);
nor U17346 (N_17346,N_16832,N_17038);
and U17347 (N_17347,N_16861,N_16893);
and U17348 (N_17348,N_17069,N_16954);
or U17349 (N_17349,N_17181,N_17191);
xor U17350 (N_17350,N_16811,N_17026);
xor U17351 (N_17351,N_16824,N_17198);
xor U17352 (N_17352,N_17006,N_16961);
xnor U17353 (N_17353,N_17186,N_17171);
nand U17354 (N_17354,N_17043,N_17190);
and U17355 (N_17355,N_17071,N_16892);
nand U17356 (N_17356,N_17085,N_16823);
and U17357 (N_17357,N_16890,N_17194);
nor U17358 (N_17358,N_17169,N_16972);
xor U17359 (N_17359,N_17083,N_16855);
xor U17360 (N_17360,N_16951,N_16949);
nand U17361 (N_17361,N_17179,N_17068);
and U17362 (N_17362,N_16827,N_16917);
nor U17363 (N_17363,N_16932,N_17076);
nor U17364 (N_17364,N_17084,N_17165);
or U17365 (N_17365,N_17170,N_17129);
and U17366 (N_17366,N_17185,N_16830);
nand U17367 (N_17367,N_17136,N_16918);
xnor U17368 (N_17368,N_16995,N_16842);
or U17369 (N_17369,N_17176,N_16803);
xnor U17370 (N_17370,N_17166,N_16953);
xor U17371 (N_17371,N_17145,N_16853);
or U17372 (N_17372,N_16850,N_16992);
or U17373 (N_17373,N_17070,N_16859);
or U17374 (N_17374,N_17012,N_16910);
and U17375 (N_17375,N_16985,N_17164);
and U17376 (N_17376,N_17056,N_17063);
or U17377 (N_17377,N_17055,N_16810);
and U17378 (N_17378,N_17187,N_17017);
nor U17379 (N_17379,N_16858,N_17097);
or U17380 (N_17380,N_16903,N_16922);
or U17381 (N_17381,N_17093,N_16856);
or U17382 (N_17382,N_16889,N_16898);
nand U17383 (N_17383,N_17156,N_16818);
or U17384 (N_17384,N_17072,N_16950);
nand U17385 (N_17385,N_17091,N_17122);
or U17386 (N_17386,N_17061,N_17065);
nand U17387 (N_17387,N_16940,N_17199);
or U17388 (N_17388,N_16908,N_16822);
and U17389 (N_17389,N_16963,N_16970);
or U17390 (N_17390,N_16896,N_16876);
nor U17391 (N_17391,N_17183,N_16913);
nand U17392 (N_17392,N_17031,N_16807);
and U17393 (N_17393,N_17142,N_17157);
and U17394 (N_17394,N_17189,N_17178);
nand U17395 (N_17395,N_16891,N_17096);
xor U17396 (N_17396,N_17139,N_16875);
and U17397 (N_17397,N_16943,N_16863);
nor U17398 (N_17398,N_16831,N_17034);
and U17399 (N_17399,N_17067,N_16906);
and U17400 (N_17400,N_16890,N_17115);
and U17401 (N_17401,N_16802,N_17068);
nor U17402 (N_17402,N_16885,N_16812);
nor U17403 (N_17403,N_17147,N_17150);
nor U17404 (N_17404,N_16824,N_17034);
nor U17405 (N_17405,N_17109,N_17183);
or U17406 (N_17406,N_16912,N_16965);
nand U17407 (N_17407,N_16800,N_17142);
xor U17408 (N_17408,N_17012,N_17091);
xnor U17409 (N_17409,N_17010,N_17016);
and U17410 (N_17410,N_16932,N_17146);
nor U17411 (N_17411,N_16900,N_16864);
nand U17412 (N_17412,N_17164,N_16806);
nand U17413 (N_17413,N_17052,N_16801);
and U17414 (N_17414,N_17137,N_16891);
xnor U17415 (N_17415,N_17127,N_16848);
nor U17416 (N_17416,N_16818,N_17172);
and U17417 (N_17417,N_16802,N_16915);
nand U17418 (N_17418,N_16802,N_16994);
and U17419 (N_17419,N_17155,N_16805);
or U17420 (N_17420,N_17025,N_16877);
nor U17421 (N_17421,N_16800,N_16960);
and U17422 (N_17422,N_16810,N_17092);
or U17423 (N_17423,N_16949,N_16966);
nand U17424 (N_17424,N_17151,N_16865);
or U17425 (N_17425,N_17081,N_16922);
nor U17426 (N_17426,N_16871,N_17084);
and U17427 (N_17427,N_16842,N_17051);
xor U17428 (N_17428,N_17046,N_17124);
nor U17429 (N_17429,N_16846,N_17127);
nor U17430 (N_17430,N_17117,N_17196);
nand U17431 (N_17431,N_17007,N_16933);
or U17432 (N_17432,N_16992,N_17103);
nand U17433 (N_17433,N_16875,N_16870);
and U17434 (N_17434,N_17166,N_17044);
nand U17435 (N_17435,N_16886,N_17114);
or U17436 (N_17436,N_16961,N_17013);
or U17437 (N_17437,N_16936,N_17047);
or U17438 (N_17438,N_16869,N_16874);
and U17439 (N_17439,N_17096,N_17030);
nor U17440 (N_17440,N_17060,N_17150);
xor U17441 (N_17441,N_16967,N_17091);
xor U17442 (N_17442,N_16935,N_17111);
xor U17443 (N_17443,N_17150,N_16811);
or U17444 (N_17444,N_16968,N_17012);
and U17445 (N_17445,N_17062,N_16932);
and U17446 (N_17446,N_16915,N_16998);
xor U17447 (N_17447,N_16807,N_17020);
nor U17448 (N_17448,N_16952,N_16838);
or U17449 (N_17449,N_16807,N_17166);
and U17450 (N_17450,N_17177,N_17139);
and U17451 (N_17451,N_16978,N_16832);
nand U17452 (N_17452,N_16974,N_16985);
or U17453 (N_17453,N_17116,N_17056);
or U17454 (N_17454,N_17132,N_17008);
and U17455 (N_17455,N_16932,N_17016);
nor U17456 (N_17456,N_16953,N_17193);
xnor U17457 (N_17457,N_16888,N_16909);
and U17458 (N_17458,N_17011,N_16851);
and U17459 (N_17459,N_16827,N_16967);
xor U17460 (N_17460,N_17123,N_17184);
nand U17461 (N_17461,N_16818,N_17106);
xnor U17462 (N_17462,N_16926,N_17068);
nand U17463 (N_17463,N_17140,N_17059);
or U17464 (N_17464,N_17081,N_16895);
nor U17465 (N_17465,N_16856,N_17024);
and U17466 (N_17466,N_17058,N_17011);
and U17467 (N_17467,N_17000,N_16821);
and U17468 (N_17468,N_17015,N_17017);
and U17469 (N_17469,N_16966,N_16807);
and U17470 (N_17470,N_17076,N_17167);
and U17471 (N_17471,N_16894,N_16871);
and U17472 (N_17472,N_17100,N_16995);
and U17473 (N_17473,N_17125,N_16907);
nor U17474 (N_17474,N_16913,N_16828);
or U17475 (N_17475,N_16892,N_17035);
or U17476 (N_17476,N_16896,N_17018);
nand U17477 (N_17477,N_16903,N_17194);
or U17478 (N_17478,N_16921,N_17057);
xor U17479 (N_17479,N_17101,N_17078);
or U17480 (N_17480,N_17015,N_17048);
nor U17481 (N_17481,N_17179,N_16935);
xor U17482 (N_17482,N_16815,N_16857);
or U17483 (N_17483,N_16895,N_16940);
or U17484 (N_17484,N_16843,N_17154);
or U17485 (N_17485,N_16891,N_16926);
nor U17486 (N_17486,N_17163,N_16894);
nand U17487 (N_17487,N_17107,N_16996);
nand U17488 (N_17488,N_17118,N_16938);
nor U17489 (N_17489,N_16978,N_17106);
nand U17490 (N_17490,N_17056,N_16862);
nand U17491 (N_17491,N_17153,N_17018);
or U17492 (N_17492,N_17192,N_17164);
nor U17493 (N_17493,N_17007,N_16981);
xor U17494 (N_17494,N_17127,N_16862);
and U17495 (N_17495,N_16889,N_17030);
or U17496 (N_17496,N_17071,N_17143);
and U17497 (N_17497,N_17089,N_17162);
xnor U17498 (N_17498,N_16867,N_16919);
or U17499 (N_17499,N_17125,N_16879);
and U17500 (N_17500,N_17069,N_16859);
and U17501 (N_17501,N_17119,N_16826);
nor U17502 (N_17502,N_16946,N_16878);
xnor U17503 (N_17503,N_16811,N_16803);
nand U17504 (N_17504,N_16857,N_16942);
nor U17505 (N_17505,N_17137,N_17104);
nand U17506 (N_17506,N_17032,N_16884);
xnor U17507 (N_17507,N_17177,N_17058);
and U17508 (N_17508,N_17059,N_16835);
nand U17509 (N_17509,N_17029,N_17143);
or U17510 (N_17510,N_17167,N_17016);
xor U17511 (N_17511,N_17085,N_17151);
nand U17512 (N_17512,N_16931,N_17020);
or U17513 (N_17513,N_17035,N_16804);
and U17514 (N_17514,N_16895,N_16811);
and U17515 (N_17515,N_16986,N_17043);
and U17516 (N_17516,N_16918,N_16957);
xnor U17517 (N_17517,N_16891,N_17190);
and U17518 (N_17518,N_17102,N_17105);
xnor U17519 (N_17519,N_17108,N_17095);
nand U17520 (N_17520,N_17108,N_17005);
xor U17521 (N_17521,N_16921,N_16969);
or U17522 (N_17522,N_16932,N_16931);
nand U17523 (N_17523,N_16814,N_17054);
nor U17524 (N_17524,N_16942,N_17086);
and U17525 (N_17525,N_17110,N_17013);
xor U17526 (N_17526,N_17126,N_16880);
and U17527 (N_17527,N_17140,N_16965);
nor U17528 (N_17528,N_16993,N_17160);
and U17529 (N_17529,N_17067,N_16943);
or U17530 (N_17530,N_17193,N_17104);
xor U17531 (N_17531,N_17077,N_16944);
nand U17532 (N_17532,N_17061,N_16922);
nand U17533 (N_17533,N_17176,N_17062);
or U17534 (N_17534,N_17165,N_16973);
nor U17535 (N_17535,N_16914,N_17102);
and U17536 (N_17536,N_16848,N_16923);
or U17537 (N_17537,N_16908,N_17180);
xor U17538 (N_17538,N_16889,N_17187);
nor U17539 (N_17539,N_16864,N_16997);
and U17540 (N_17540,N_16943,N_17087);
or U17541 (N_17541,N_16951,N_17057);
xnor U17542 (N_17542,N_17062,N_17071);
and U17543 (N_17543,N_17063,N_17030);
nand U17544 (N_17544,N_16835,N_17174);
and U17545 (N_17545,N_16887,N_16874);
nor U17546 (N_17546,N_17055,N_17037);
nand U17547 (N_17547,N_16888,N_16864);
nand U17548 (N_17548,N_16953,N_16852);
nand U17549 (N_17549,N_16958,N_17137);
nand U17550 (N_17550,N_17042,N_16828);
xnor U17551 (N_17551,N_17172,N_17166);
xor U17552 (N_17552,N_16904,N_16863);
nor U17553 (N_17553,N_16951,N_17189);
and U17554 (N_17554,N_16976,N_17198);
xnor U17555 (N_17555,N_16995,N_17057);
and U17556 (N_17556,N_16953,N_16805);
nor U17557 (N_17557,N_16917,N_16967);
and U17558 (N_17558,N_17039,N_17156);
or U17559 (N_17559,N_16808,N_16800);
xor U17560 (N_17560,N_16917,N_17166);
nand U17561 (N_17561,N_16888,N_17020);
nand U17562 (N_17562,N_16856,N_17101);
and U17563 (N_17563,N_17083,N_16944);
xor U17564 (N_17564,N_16883,N_16814);
or U17565 (N_17565,N_16839,N_17032);
or U17566 (N_17566,N_17022,N_16974);
or U17567 (N_17567,N_17139,N_16947);
nor U17568 (N_17568,N_16897,N_17138);
nand U17569 (N_17569,N_17192,N_17196);
nand U17570 (N_17570,N_16928,N_16875);
xnor U17571 (N_17571,N_16950,N_16952);
nor U17572 (N_17572,N_16867,N_17122);
nand U17573 (N_17573,N_16987,N_16890);
or U17574 (N_17574,N_16839,N_17092);
or U17575 (N_17575,N_17193,N_16803);
nor U17576 (N_17576,N_17158,N_17128);
nand U17577 (N_17577,N_16970,N_17195);
and U17578 (N_17578,N_16882,N_17002);
or U17579 (N_17579,N_17178,N_17055);
nor U17580 (N_17580,N_17001,N_16833);
nand U17581 (N_17581,N_17016,N_17198);
nand U17582 (N_17582,N_17154,N_16943);
or U17583 (N_17583,N_16951,N_17065);
or U17584 (N_17584,N_16820,N_16860);
or U17585 (N_17585,N_16906,N_17111);
and U17586 (N_17586,N_17076,N_17125);
nand U17587 (N_17587,N_17158,N_16903);
nand U17588 (N_17588,N_17077,N_16825);
xor U17589 (N_17589,N_17110,N_17194);
xnor U17590 (N_17590,N_16995,N_16944);
xor U17591 (N_17591,N_17031,N_17095);
xnor U17592 (N_17592,N_16978,N_16862);
nor U17593 (N_17593,N_16849,N_16933);
nor U17594 (N_17594,N_16913,N_16992);
or U17595 (N_17595,N_16809,N_16847);
nor U17596 (N_17596,N_17051,N_16907);
xnor U17597 (N_17597,N_16934,N_16939);
xnor U17598 (N_17598,N_17106,N_17140);
and U17599 (N_17599,N_16885,N_16934);
nand U17600 (N_17600,N_17256,N_17591);
nor U17601 (N_17601,N_17290,N_17219);
or U17602 (N_17602,N_17294,N_17531);
nor U17603 (N_17603,N_17434,N_17554);
nor U17604 (N_17604,N_17509,N_17351);
nor U17605 (N_17605,N_17289,N_17540);
nand U17606 (N_17606,N_17454,N_17566);
nand U17607 (N_17607,N_17203,N_17246);
xnor U17608 (N_17608,N_17589,N_17374);
and U17609 (N_17609,N_17369,N_17239);
or U17610 (N_17610,N_17574,N_17423);
or U17611 (N_17611,N_17295,N_17393);
xor U17612 (N_17612,N_17223,N_17302);
or U17613 (N_17613,N_17511,N_17598);
nor U17614 (N_17614,N_17495,N_17237);
xor U17615 (N_17615,N_17534,N_17499);
and U17616 (N_17616,N_17587,N_17414);
nor U17617 (N_17617,N_17451,N_17270);
nor U17618 (N_17618,N_17240,N_17292);
nand U17619 (N_17619,N_17552,N_17225);
xor U17620 (N_17620,N_17400,N_17426);
or U17621 (N_17621,N_17593,N_17530);
nand U17622 (N_17622,N_17396,N_17323);
or U17623 (N_17623,N_17267,N_17420);
nor U17624 (N_17624,N_17250,N_17583);
nor U17625 (N_17625,N_17458,N_17529);
nor U17626 (N_17626,N_17522,N_17367);
and U17627 (N_17627,N_17291,N_17427);
nor U17628 (N_17628,N_17460,N_17537);
nand U17629 (N_17629,N_17413,N_17504);
and U17630 (N_17630,N_17425,N_17263);
or U17631 (N_17631,N_17354,N_17325);
nand U17632 (N_17632,N_17415,N_17462);
xor U17633 (N_17633,N_17528,N_17467);
xor U17634 (N_17634,N_17503,N_17404);
nand U17635 (N_17635,N_17496,N_17355);
and U17636 (N_17636,N_17334,N_17359);
nor U17637 (N_17637,N_17444,N_17274);
nand U17638 (N_17638,N_17500,N_17306);
and U17639 (N_17639,N_17200,N_17364);
nand U17640 (N_17640,N_17436,N_17582);
and U17641 (N_17641,N_17391,N_17505);
xnor U17642 (N_17642,N_17271,N_17486);
nand U17643 (N_17643,N_17258,N_17304);
xnor U17644 (N_17644,N_17555,N_17429);
and U17645 (N_17645,N_17453,N_17517);
or U17646 (N_17646,N_17314,N_17287);
nor U17647 (N_17647,N_17281,N_17218);
or U17648 (N_17648,N_17553,N_17432);
xnor U17649 (N_17649,N_17483,N_17241);
xnor U17650 (N_17650,N_17443,N_17470);
nor U17651 (N_17651,N_17473,N_17547);
or U17652 (N_17652,N_17560,N_17515);
and U17653 (N_17653,N_17206,N_17526);
nor U17654 (N_17654,N_17348,N_17224);
xnor U17655 (N_17655,N_17254,N_17447);
or U17656 (N_17656,N_17232,N_17253);
xor U17657 (N_17657,N_17559,N_17578);
nor U17658 (N_17658,N_17358,N_17356);
xnor U17659 (N_17659,N_17216,N_17539);
nor U17660 (N_17660,N_17576,N_17410);
and U17661 (N_17661,N_17328,N_17373);
xnor U17662 (N_17662,N_17561,N_17536);
xor U17663 (N_17663,N_17312,N_17448);
nor U17664 (N_17664,N_17442,N_17320);
or U17665 (N_17665,N_17450,N_17366);
and U17666 (N_17666,N_17471,N_17251);
xnor U17667 (N_17667,N_17247,N_17384);
or U17668 (N_17668,N_17405,N_17335);
nor U17669 (N_17669,N_17278,N_17370);
xnor U17670 (N_17670,N_17379,N_17494);
nand U17671 (N_17671,N_17466,N_17599);
and U17672 (N_17672,N_17376,N_17333);
and U17673 (N_17673,N_17513,N_17437);
nand U17674 (N_17674,N_17244,N_17277);
and U17675 (N_17675,N_17497,N_17301);
nand U17676 (N_17676,N_17449,N_17362);
or U17677 (N_17677,N_17523,N_17319);
nor U17678 (N_17678,N_17435,N_17548);
nand U17679 (N_17679,N_17461,N_17406);
xor U17680 (N_17680,N_17516,N_17363);
xnor U17681 (N_17681,N_17493,N_17543);
nand U17682 (N_17682,N_17243,N_17378);
nand U17683 (N_17683,N_17299,N_17303);
and U17684 (N_17684,N_17257,N_17440);
nand U17685 (N_17685,N_17468,N_17490);
nor U17686 (N_17686,N_17395,N_17550);
or U17687 (N_17687,N_17212,N_17472);
nand U17688 (N_17688,N_17527,N_17389);
and U17689 (N_17689,N_17214,N_17399);
or U17690 (N_17690,N_17455,N_17307);
xor U17691 (N_17691,N_17422,N_17383);
and U17692 (N_17692,N_17365,N_17562);
or U17693 (N_17693,N_17315,N_17568);
nand U17694 (N_17694,N_17545,N_17236);
or U17695 (N_17695,N_17242,N_17204);
and U17696 (N_17696,N_17482,N_17342);
nand U17697 (N_17697,N_17533,N_17469);
and U17698 (N_17698,N_17514,N_17345);
xor U17699 (N_17699,N_17344,N_17538);
nand U17700 (N_17700,N_17549,N_17403);
and U17701 (N_17701,N_17313,N_17228);
nor U17702 (N_17702,N_17544,N_17512);
or U17703 (N_17703,N_17387,N_17476);
and U17704 (N_17704,N_17201,N_17329);
nor U17705 (N_17705,N_17507,N_17408);
nand U17706 (N_17706,N_17282,N_17248);
or U17707 (N_17707,N_17430,N_17491);
nor U17708 (N_17708,N_17385,N_17532);
nor U17709 (N_17709,N_17226,N_17592);
or U17710 (N_17710,N_17388,N_17317);
and U17711 (N_17711,N_17519,N_17298);
or U17712 (N_17712,N_17322,N_17336);
or U17713 (N_17713,N_17398,N_17424);
and U17714 (N_17714,N_17478,N_17594);
and U17715 (N_17715,N_17488,N_17577);
or U17716 (N_17716,N_17372,N_17474);
nand U17717 (N_17717,N_17445,N_17564);
nand U17718 (N_17718,N_17418,N_17205);
and U17719 (N_17719,N_17262,N_17390);
xnor U17720 (N_17720,N_17520,N_17268);
nor U17721 (N_17721,N_17350,N_17202);
or U17722 (N_17722,N_17284,N_17318);
nor U17723 (N_17723,N_17394,N_17338);
nor U17724 (N_17724,N_17211,N_17381);
nand U17725 (N_17725,N_17215,N_17433);
nor U17726 (N_17726,N_17386,N_17286);
and U17727 (N_17727,N_17492,N_17407);
and U17728 (N_17728,N_17441,N_17402);
and U17729 (N_17729,N_17464,N_17227);
or U17730 (N_17730,N_17296,N_17457);
xor U17731 (N_17731,N_17276,N_17337);
nand U17732 (N_17732,N_17480,N_17249);
nand U17733 (N_17733,N_17580,N_17331);
nand U17734 (N_17734,N_17309,N_17446);
and U17735 (N_17735,N_17475,N_17573);
and U17736 (N_17736,N_17349,N_17222);
nand U17737 (N_17737,N_17273,N_17220);
nor U17738 (N_17738,N_17259,N_17481);
nand U17739 (N_17739,N_17221,N_17459);
and U17740 (N_17740,N_17238,N_17285);
nor U17741 (N_17741,N_17368,N_17330);
or U17742 (N_17742,N_17579,N_17308);
and U17743 (N_17743,N_17570,N_17524);
nor U17744 (N_17744,N_17347,N_17272);
xor U17745 (N_17745,N_17421,N_17264);
and U17746 (N_17746,N_17510,N_17485);
xnor U17747 (N_17747,N_17326,N_17557);
or U17748 (N_17748,N_17518,N_17556);
xor U17749 (N_17749,N_17585,N_17230);
nand U17750 (N_17750,N_17300,N_17452);
nand U17751 (N_17751,N_17586,N_17305);
and U17752 (N_17752,N_17275,N_17332);
xnor U17753 (N_17753,N_17558,N_17575);
nand U17754 (N_17754,N_17502,N_17357);
and U17755 (N_17755,N_17584,N_17563);
nor U17756 (N_17756,N_17261,N_17489);
nand U17757 (N_17757,N_17525,N_17417);
or U17758 (N_17758,N_17377,N_17311);
nand U17759 (N_17759,N_17506,N_17297);
nand U17760 (N_17760,N_17361,N_17590);
and U17761 (N_17761,N_17283,N_17572);
nand U17762 (N_17762,N_17213,N_17465);
and U17763 (N_17763,N_17431,N_17463);
and U17764 (N_17764,N_17498,N_17569);
xor U17765 (N_17765,N_17419,N_17375);
or U17766 (N_17766,N_17346,N_17234);
nand U17767 (N_17767,N_17245,N_17380);
and U17768 (N_17768,N_17265,N_17508);
nand U17769 (N_17769,N_17551,N_17401);
or U17770 (N_17770,N_17280,N_17229);
nand U17771 (N_17771,N_17542,N_17210);
xnor U17772 (N_17772,N_17321,N_17231);
or U17773 (N_17773,N_17416,N_17327);
and U17774 (N_17774,N_17581,N_17324);
nand U17775 (N_17775,N_17535,N_17343);
or U17776 (N_17776,N_17288,N_17521);
xnor U17777 (N_17777,N_17255,N_17487);
nor U17778 (N_17778,N_17207,N_17341);
nand U17779 (N_17779,N_17597,N_17546);
nand U17780 (N_17780,N_17411,N_17352);
and U17781 (N_17781,N_17392,N_17208);
nor U17782 (N_17782,N_17233,N_17428);
nand U17783 (N_17783,N_17260,N_17567);
xnor U17784 (N_17784,N_17595,N_17266);
or U17785 (N_17785,N_17479,N_17217);
or U17786 (N_17786,N_17439,N_17269);
xnor U17787 (N_17787,N_17501,N_17382);
and U17788 (N_17788,N_17571,N_17293);
nand U17789 (N_17789,N_17360,N_17371);
nand U17790 (N_17790,N_17310,N_17565);
xor U17791 (N_17791,N_17438,N_17209);
xor U17792 (N_17792,N_17339,N_17541);
or U17793 (N_17793,N_17340,N_17484);
nor U17794 (N_17794,N_17353,N_17477);
or U17795 (N_17795,N_17235,N_17412);
nor U17796 (N_17796,N_17456,N_17409);
or U17797 (N_17797,N_17588,N_17252);
nand U17798 (N_17798,N_17397,N_17316);
and U17799 (N_17799,N_17279,N_17596);
xor U17800 (N_17800,N_17485,N_17570);
nor U17801 (N_17801,N_17595,N_17480);
nor U17802 (N_17802,N_17571,N_17389);
nor U17803 (N_17803,N_17492,N_17574);
and U17804 (N_17804,N_17344,N_17290);
nand U17805 (N_17805,N_17317,N_17236);
and U17806 (N_17806,N_17241,N_17388);
or U17807 (N_17807,N_17510,N_17596);
nand U17808 (N_17808,N_17289,N_17282);
and U17809 (N_17809,N_17259,N_17313);
or U17810 (N_17810,N_17494,N_17339);
or U17811 (N_17811,N_17370,N_17239);
nor U17812 (N_17812,N_17223,N_17586);
nand U17813 (N_17813,N_17259,N_17325);
or U17814 (N_17814,N_17404,N_17521);
and U17815 (N_17815,N_17313,N_17343);
nand U17816 (N_17816,N_17583,N_17220);
and U17817 (N_17817,N_17303,N_17501);
xnor U17818 (N_17818,N_17244,N_17437);
or U17819 (N_17819,N_17408,N_17544);
nor U17820 (N_17820,N_17461,N_17479);
or U17821 (N_17821,N_17269,N_17351);
or U17822 (N_17822,N_17249,N_17383);
and U17823 (N_17823,N_17324,N_17571);
nand U17824 (N_17824,N_17457,N_17432);
and U17825 (N_17825,N_17597,N_17579);
nand U17826 (N_17826,N_17567,N_17544);
nand U17827 (N_17827,N_17405,N_17535);
nand U17828 (N_17828,N_17392,N_17234);
nor U17829 (N_17829,N_17244,N_17283);
xnor U17830 (N_17830,N_17360,N_17573);
nor U17831 (N_17831,N_17236,N_17544);
nand U17832 (N_17832,N_17272,N_17491);
or U17833 (N_17833,N_17370,N_17593);
or U17834 (N_17834,N_17326,N_17384);
or U17835 (N_17835,N_17258,N_17331);
nor U17836 (N_17836,N_17321,N_17360);
nor U17837 (N_17837,N_17378,N_17468);
xor U17838 (N_17838,N_17432,N_17236);
nand U17839 (N_17839,N_17341,N_17251);
nand U17840 (N_17840,N_17267,N_17402);
nor U17841 (N_17841,N_17595,N_17352);
and U17842 (N_17842,N_17261,N_17344);
or U17843 (N_17843,N_17565,N_17575);
xor U17844 (N_17844,N_17428,N_17442);
and U17845 (N_17845,N_17520,N_17396);
nor U17846 (N_17846,N_17386,N_17551);
nor U17847 (N_17847,N_17425,N_17389);
or U17848 (N_17848,N_17502,N_17367);
and U17849 (N_17849,N_17293,N_17462);
nor U17850 (N_17850,N_17509,N_17264);
nand U17851 (N_17851,N_17449,N_17288);
or U17852 (N_17852,N_17571,N_17427);
xnor U17853 (N_17853,N_17450,N_17321);
or U17854 (N_17854,N_17483,N_17509);
nand U17855 (N_17855,N_17393,N_17458);
nand U17856 (N_17856,N_17326,N_17286);
nor U17857 (N_17857,N_17317,N_17543);
nor U17858 (N_17858,N_17387,N_17440);
nor U17859 (N_17859,N_17416,N_17550);
nand U17860 (N_17860,N_17283,N_17473);
nand U17861 (N_17861,N_17493,N_17596);
nor U17862 (N_17862,N_17303,N_17272);
xnor U17863 (N_17863,N_17345,N_17593);
xnor U17864 (N_17864,N_17441,N_17373);
or U17865 (N_17865,N_17415,N_17499);
or U17866 (N_17866,N_17423,N_17243);
xor U17867 (N_17867,N_17400,N_17587);
nand U17868 (N_17868,N_17516,N_17496);
nor U17869 (N_17869,N_17497,N_17228);
or U17870 (N_17870,N_17280,N_17231);
or U17871 (N_17871,N_17575,N_17274);
and U17872 (N_17872,N_17263,N_17249);
xor U17873 (N_17873,N_17512,N_17315);
or U17874 (N_17874,N_17519,N_17408);
and U17875 (N_17875,N_17389,N_17594);
nand U17876 (N_17876,N_17464,N_17482);
and U17877 (N_17877,N_17384,N_17275);
nand U17878 (N_17878,N_17365,N_17278);
xnor U17879 (N_17879,N_17469,N_17437);
and U17880 (N_17880,N_17303,N_17311);
nand U17881 (N_17881,N_17498,N_17225);
nor U17882 (N_17882,N_17469,N_17347);
and U17883 (N_17883,N_17474,N_17392);
or U17884 (N_17884,N_17278,N_17416);
xnor U17885 (N_17885,N_17559,N_17218);
xnor U17886 (N_17886,N_17580,N_17492);
nand U17887 (N_17887,N_17335,N_17414);
xnor U17888 (N_17888,N_17223,N_17348);
xor U17889 (N_17889,N_17245,N_17238);
xor U17890 (N_17890,N_17512,N_17479);
or U17891 (N_17891,N_17598,N_17351);
xor U17892 (N_17892,N_17325,N_17473);
xnor U17893 (N_17893,N_17329,N_17231);
nor U17894 (N_17894,N_17544,N_17311);
nand U17895 (N_17895,N_17220,N_17441);
xor U17896 (N_17896,N_17594,N_17579);
xor U17897 (N_17897,N_17264,N_17534);
xor U17898 (N_17898,N_17530,N_17265);
nand U17899 (N_17899,N_17422,N_17453);
or U17900 (N_17900,N_17462,N_17315);
or U17901 (N_17901,N_17589,N_17503);
or U17902 (N_17902,N_17513,N_17419);
or U17903 (N_17903,N_17274,N_17558);
or U17904 (N_17904,N_17230,N_17416);
and U17905 (N_17905,N_17264,N_17401);
xnor U17906 (N_17906,N_17399,N_17462);
or U17907 (N_17907,N_17598,N_17487);
and U17908 (N_17908,N_17563,N_17484);
or U17909 (N_17909,N_17491,N_17271);
nand U17910 (N_17910,N_17401,N_17580);
or U17911 (N_17911,N_17499,N_17253);
or U17912 (N_17912,N_17238,N_17205);
nand U17913 (N_17913,N_17479,N_17420);
nor U17914 (N_17914,N_17353,N_17397);
xor U17915 (N_17915,N_17543,N_17290);
xor U17916 (N_17916,N_17297,N_17466);
or U17917 (N_17917,N_17562,N_17443);
and U17918 (N_17918,N_17299,N_17373);
nand U17919 (N_17919,N_17328,N_17208);
nand U17920 (N_17920,N_17475,N_17343);
and U17921 (N_17921,N_17216,N_17268);
nor U17922 (N_17922,N_17570,N_17513);
xor U17923 (N_17923,N_17328,N_17496);
nand U17924 (N_17924,N_17213,N_17395);
xnor U17925 (N_17925,N_17487,N_17217);
nor U17926 (N_17926,N_17417,N_17434);
xor U17927 (N_17927,N_17201,N_17474);
or U17928 (N_17928,N_17296,N_17290);
nor U17929 (N_17929,N_17438,N_17300);
xor U17930 (N_17930,N_17519,N_17365);
nor U17931 (N_17931,N_17412,N_17534);
xnor U17932 (N_17932,N_17219,N_17229);
and U17933 (N_17933,N_17291,N_17361);
nor U17934 (N_17934,N_17443,N_17251);
xor U17935 (N_17935,N_17546,N_17521);
and U17936 (N_17936,N_17474,N_17357);
xor U17937 (N_17937,N_17463,N_17309);
nor U17938 (N_17938,N_17366,N_17498);
and U17939 (N_17939,N_17566,N_17471);
or U17940 (N_17940,N_17217,N_17275);
nand U17941 (N_17941,N_17220,N_17232);
and U17942 (N_17942,N_17227,N_17267);
nor U17943 (N_17943,N_17571,N_17267);
nor U17944 (N_17944,N_17439,N_17223);
xor U17945 (N_17945,N_17376,N_17415);
xor U17946 (N_17946,N_17506,N_17451);
nor U17947 (N_17947,N_17286,N_17299);
and U17948 (N_17948,N_17463,N_17376);
nor U17949 (N_17949,N_17211,N_17377);
and U17950 (N_17950,N_17441,N_17333);
and U17951 (N_17951,N_17447,N_17544);
or U17952 (N_17952,N_17560,N_17531);
nor U17953 (N_17953,N_17241,N_17282);
nor U17954 (N_17954,N_17316,N_17478);
nand U17955 (N_17955,N_17216,N_17487);
and U17956 (N_17956,N_17345,N_17238);
nand U17957 (N_17957,N_17575,N_17403);
nand U17958 (N_17958,N_17364,N_17323);
xor U17959 (N_17959,N_17302,N_17517);
nor U17960 (N_17960,N_17417,N_17408);
or U17961 (N_17961,N_17261,N_17230);
nor U17962 (N_17962,N_17532,N_17361);
nor U17963 (N_17963,N_17204,N_17209);
and U17964 (N_17964,N_17485,N_17384);
and U17965 (N_17965,N_17336,N_17253);
and U17966 (N_17966,N_17525,N_17365);
nor U17967 (N_17967,N_17328,N_17560);
xnor U17968 (N_17968,N_17431,N_17222);
nor U17969 (N_17969,N_17493,N_17569);
or U17970 (N_17970,N_17400,N_17367);
nor U17971 (N_17971,N_17525,N_17313);
or U17972 (N_17972,N_17475,N_17504);
or U17973 (N_17973,N_17245,N_17345);
nand U17974 (N_17974,N_17296,N_17348);
nand U17975 (N_17975,N_17466,N_17493);
nor U17976 (N_17976,N_17372,N_17329);
or U17977 (N_17977,N_17447,N_17245);
nor U17978 (N_17978,N_17499,N_17421);
nor U17979 (N_17979,N_17486,N_17230);
and U17980 (N_17980,N_17428,N_17586);
xor U17981 (N_17981,N_17413,N_17242);
and U17982 (N_17982,N_17303,N_17308);
or U17983 (N_17983,N_17530,N_17263);
nor U17984 (N_17984,N_17322,N_17447);
nor U17985 (N_17985,N_17346,N_17456);
and U17986 (N_17986,N_17319,N_17232);
nor U17987 (N_17987,N_17427,N_17483);
nand U17988 (N_17988,N_17518,N_17485);
xnor U17989 (N_17989,N_17453,N_17423);
nor U17990 (N_17990,N_17561,N_17206);
xnor U17991 (N_17991,N_17257,N_17314);
or U17992 (N_17992,N_17400,N_17340);
xor U17993 (N_17993,N_17355,N_17523);
and U17994 (N_17994,N_17271,N_17571);
nor U17995 (N_17995,N_17385,N_17361);
and U17996 (N_17996,N_17345,N_17509);
nor U17997 (N_17997,N_17249,N_17418);
and U17998 (N_17998,N_17291,N_17317);
xor U17999 (N_17999,N_17297,N_17560);
or U18000 (N_18000,N_17773,N_17696);
or U18001 (N_18001,N_17792,N_17655);
xnor U18002 (N_18002,N_17746,N_17737);
or U18003 (N_18003,N_17879,N_17791);
or U18004 (N_18004,N_17892,N_17883);
and U18005 (N_18005,N_17612,N_17925);
and U18006 (N_18006,N_17998,N_17714);
nor U18007 (N_18007,N_17888,N_17710);
xor U18008 (N_18008,N_17635,N_17797);
or U18009 (N_18009,N_17867,N_17893);
nand U18010 (N_18010,N_17795,N_17928);
and U18011 (N_18011,N_17638,N_17755);
or U18012 (N_18012,N_17924,N_17858);
nor U18013 (N_18013,N_17882,N_17663);
nand U18014 (N_18014,N_17674,N_17688);
nor U18015 (N_18015,N_17918,N_17835);
nand U18016 (N_18016,N_17813,N_17631);
or U18017 (N_18017,N_17640,N_17701);
nand U18018 (N_18018,N_17622,N_17680);
nor U18019 (N_18019,N_17643,N_17722);
nor U18020 (N_18020,N_17985,N_17717);
nand U18021 (N_18021,N_17652,N_17770);
nand U18022 (N_18022,N_17861,N_17926);
nand U18023 (N_18023,N_17846,N_17890);
and U18024 (N_18024,N_17708,N_17604);
xor U18025 (N_18025,N_17979,N_17899);
and U18026 (N_18026,N_17641,N_17745);
xor U18027 (N_18027,N_17806,N_17881);
xor U18028 (N_18028,N_17917,N_17695);
or U18029 (N_18029,N_17699,N_17627);
or U18030 (N_18030,N_17620,N_17712);
nand U18031 (N_18031,N_17771,N_17684);
nand U18032 (N_18032,N_17700,N_17816);
or U18033 (N_18033,N_17617,N_17765);
and U18034 (N_18034,N_17954,N_17841);
and U18035 (N_18035,N_17783,N_17930);
and U18036 (N_18036,N_17965,N_17839);
and U18037 (N_18037,N_17693,N_17973);
nor U18038 (N_18038,N_17984,N_17694);
or U18039 (N_18039,N_17931,N_17720);
xor U18040 (N_18040,N_17955,N_17726);
nand U18041 (N_18041,N_17686,N_17647);
and U18042 (N_18042,N_17891,N_17724);
nor U18043 (N_18043,N_17733,N_17801);
and U18044 (N_18044,N_17919,N_17789);
nand U18045 (N_18045,N_17732,N_17877);
or U18046 (N_18046,N_17796,N_17634);
nand U18047 (N_18047,N_17653,N_17731);
nand U18048 (N_18048,N_17817,N_17629);
nand U18049 (N_18049,N_17943,N_17845);
xnor U18050 (N_18050,N_17980,N_17650);
and U18051 (N_18051,N_17703,N_17802);
and U18052 (N_18052,N_17921,N_17705);
or U18053 (N_18053,N_17804,N_17934);
xor U18054 (N_18054,N_17615,N_17902);
nor U18055 (N_18055,N_17681,N_17654);
and U18056 (N_18056,N_17739,N_17898);
nor U18057 (N_18057,N_17675,N_17644);
nor U18058 (N_18058,N_17763,N_17992);
xor U18059 (N_18059,N_17608,N_17672);
xnor U18060 (N_18060,N_17905,N_17847);
xor U18061 (N_18061,N_17676,N_17865);
or U18062 (N_18062,N_17605,N_17639);
xor U18063 (N_18063,N_17912,N_17851);
and U18064 (N_18064,N_17633,N_17936);
xor U18065 (N_18065,N_17719,N_17809);
nor U18066 (N_18066,N_17750,N_17761);
nor U18067 (N_18067,N_17751,N_17968);
nand U18068 (N_18068,N_17698,N_17785);
or U18069 (N_18069,N_17683,N_17793);
and U18070 (N_18070,N_17673,N_17900);
xnor U18071 (N_18071,N_17786,N_17738);
xnor U18072 (N_18072,N_17614,N_17961);
nor U18073 (N_18073,N_17628,N_17857);
and U18074 (N_18074,N_17685,N_17971);
nor U18075 (N_18075,N_17916,N_17906);
xnor U18076 (N_18076,N_17651,N_17624);
and U18077 (N_18077,N_17963,N_17774);
nand U18078 (N_18078,N_17836,N_17807);
or U18079 (N_18079,N_17725,N_17621);
and U18080 (N_18080,N_17664,N_17929);
xnor U18081 (N_18081,N_17875,N_17866);
or U18082 (N_18082,N_17977,N_17779);
and U18083 (N_18083,N_17938,N_17728);
nor U18084 (N_18084,N_17660,N_17601);
nand U18085 (N_18085,N_17996,N_17993);
or U18086 (N_18086,N_17721,N_17994);
nor U18087 (N_18087,N_17788,N_17910);
or U18088 (N_18088,N_17850,N_17610);
xnor U18089 (N_18089,N_17966,N_17758);
xnor U18090 (N_18090,N_17715,N_17764);
nor U18091 (N_18091,N_17646,N_17702);
and U18092 (N_18092,N_17872,N_17814);
and U18093 (N_18093,N_17856,N_17939);
nor U18094 (N_18094,N_17904,N_17999);
nor U18095 (N_18095,N_17842,N_17616);
nand U18096 (N_18096,N_17838,N_17947);
nand U18097 (N_18097,N_17941,N_17778);
nand U18098 (N_18098,N_17927,N_17658);
or U18099 (N_18099,N_17920,N_17844);
and U18100 (N_18100,N_17747,N_17602);
nor U18101 (N_18101,N_17944,N_17989);
nor U18102 (N_18102,N_17670,N_17782);
xnor U18103 (N_18103,N_17908,N_17618);
nor U18104 (N_18104,N_17887,N_17830);
xnor U18105 (N_18105,N_17871,N_17709);
and U18106 (N_18106,N_17937,N_17742);
and U18107 (N_18107,N_17625,N_17642);
or U18108 (N_18108,N_17603,N_17697);
xnor U18109 (N_18109,N_17976,N_17752);
xor U18110 (N_18110,N_17945,N_17860);
xor U18111 (N_18111,N_17957,N_17983);
nand U18112 (N_18112,N_17909,N_17704);
xnor U18113 (N_18113,N_17897,N_17824);
nor U18114 (N_18114,N_17645,N_17870);
or U18115 (N_18115,N_17808,N_17707);
and U18116 (N_18116,N_17942,N_17772);
or U18117 (N_18117,N_17950,N_17744);
xor U18118 (N_18118,N_17854,N_17648);
nand U18119 (N_18119,N_17711,N_17986);
or U18120 (N_18120,N_17864,N_17834);
xnor U18121 (N_18121,N_17754,N_17922);
nor U18122 (N_18122,N_17606,N_17767);
xor U18123 (N_18123,N_17915,N_17964);
nor U18124 (N_18124,N_17874,N_17776);
or U18125 (N_18125,N_17810,N_17768);
nor U18126 (N_18126,N_17753,N_17727);
nand U18127 (N_18127,N_17649,N_17815);
nor U18128 (N_18128,N_17960,N_17769);
xor U18129 (N_18129,N_17749,N_17923);
and U18130 (N_18130,N_17690,N_17896);
nand U18131 (N_18131,N_17800,N_17607);
and U18132 (N_18132,N_17730,N_17671);
nand U18133 (N_18133,N_17829,N_17679);
nand U18134 (N_18134,N_17886,N_17831);
and U18135 (N_18135,N_17743,N_17869);
and U18136 (N_18136,N_17991,N_17656);
or U18137 (N_18137,N_17689,N_17790);
nand U18138 (N_18138,N_17862,N_17828);
and U18139 (N_18139,N_17995,N_17981);
nor U18140 (N_18140,N_17805,N_17687);
or U18141 (N_18141,N_17799,N_17833);
nor U18142 (N_18142,N_17682,N_17784);
and U18143 (N_18143,N_17885,N_17997);
nor U18144 (N_18144,N_17880,N_17818);
or U18145 (N_18145,N_17820,N_17734);
xor U18146 (N_18146,N_17781,N_17803);
nand U18147 (N_18147,N_17970,N_17812);
and U18148 (N_18148,N_17853,N_17969);
or U18149 (N_18149,N_17975,N_17787);
and U18150 (N_18150,N_17873,N_17777);
and U18151 (N_18151,N_17962,N_17878);
and U18152 (N_18152,N_17903,N_17843);
nor U18153 (N_18153,N_17766,N_17825);
or U18154 (N_18154,N_17868,N_17982);
and U18155 (N_18155,N_17756,N_17822);
xor U18156 (N_18156,N_17668,N_17667);
and U18157 (N_18157,N_17678,N_17626);
or U18158 (N_18158,N_17665,N_17819);
or U18159 (N_18159,N_17827,N_17987);
xnor U18160 (N_18160,N_17884,N_17619);
xnor U18161 (N_18161,N_17748,N_17952);
nor U18162 (N_18162,N_17848,N_17630);
and U18163 (N_18163,N_17811,N_17632);
and U18164 (N_18164,N_17859,N_17636);
or U18165 (N_18165,N_17613,N_17911);
nand U18166 (N_18166,N_17823,N_17716);
or U18167 (N_18167,N_17895,N_17953);
nand U18168 (N_18168,N_17935,N_17736);
and U18169 (N_18169,N_17959,N_17889);
nand U18170 (N_18170,N_17757,N_17609);
nand U18171 (N_18171,N_17623,N_17978);
nor U18172 (N_18172,N_17913,N_17932);
or U18173 (N_18173,N_17760,N_17659);
nand U18174 (N_18174,N_17949,N_17972);
nor U18175 (N_18175,N_17762,N_17677);
nand U18176 (N_18176,N_17914,N_17691);
nand U18177 (N_18177,N_17826,N_17863);
or U18178 (N_18178,N_17948,N_17735);
and U18179 (N_18179,N_17907,N_17821);
nand U18180 (N_18180,N_17706,N_17974);
or U18181 (N_18181,N_17600,N_17990);
nand U18182 (N_18182,N_17780,N_17666);
nand U18183 (N_18183,N_17958,N_17832);
nor U18184 (N_18184,N_17852,N_17840);
or U18185 (N_18185,N_17894,N_17775);
or U18186 (N_18186,N_17901,N_17798);
nand U18187 (N_18187,N_17723,N_17713);
nor U18188 (N_18188,N_17956,N_17692);
or U18189 (N_18189,N_17988,N_17951);
or U18190 (N_18190,N_17855,N_17662);
xor U18191 (N_18191,N_17661,N_17837);
or U18192 (N_18192,N_17611,N_17718);
nand U18193 (N_18193,N_17849,N_17657);
xnor U18194 (N_18194,N_17876,N_17741);
nand U18195 (N_18195,N_17794,N_17729);
and U18196 (N_18196,N_17967,N_17637);
nand U18197 (N_18197,N_17940,N_17759);
xnor U18198 (N_18198,N_17933,N_17740);
or U18199 (N_18199,N_17669,N_17946);
nor U18200 (N_18200,N_17638,N_17993);
xor U18201 (N_18201,N_17990,N_17778);
nand U18202 (N_18202,N_17739,N_17907);
and U18203 (N_18203,N_17650,N_17623);
xor U18204 (N_18204,N_17950,N_17868);
and U18205 (N_18205,N_17970,N_17826);
or U18206 (N_18206,N_17915,N_17803);
nand U18207 (N_18207,N_17862,N_17848);
and U18208 (N_18208,N_17909,N_17661);
or U18209 (N_18209,N_17952,N_17971);
nor U18210 (N_18210,N_17875,N_17910);
and U18211 (N_18211,N_17786,N_17979);
nor U18212 (N_18212,N_17944,N_17614);
or U18213 (N_18213,N_17713,N_17970);
nor U18214 (N_18214,N_17821,N_17850);
nand U18215 (N_18215,N_17840,N_17985);
xor U18216 (N_18216,N_17910,N_17690);
nand U18217 (N_18217,N_17887,N_17988);
and U18218 (N_18218,N_17855,N_17876);
nand U18219 (N_18219,N_17709,N_17695);
or U18220 (N_18220,N_17715,N_17722);
and U18221 (N_18221,N_17904,N_17762);
xor U18222 (N_18222,N_17856,N_17843);
nor U18223 (N_18223,N_17827,N_17995);
nor U18224 (N_18224,N_17815,N_17822);
nand U18225 (N_18225,N_17655,N_17802);
xnor U18226 (N_18226,N_17880,N_17643);
nand U18227 (N_18227,N_17946,N_17890);
nand U18228 (N_18228,N_17625,N_17681);
xor U18229 (N_18229,N_17617,N_17703);
nor U18230 (N_18230,N_17959,N_17697);
and U18231 (N_18231,N_17750,N_17818);
nand U18232 (N_18232,N_17664,N_17993);
nand U18233 (N_18233,N_17862,N_17633);
xnor U18234 (N_18234,N_17836,N_17718);
nor U18235 (N_18235,N_17861,N_17975);
nand U18236 (N_18236,N_17670,N_17883);
xnor U18237 (N_18237,N_17815,N_17609);
nand U18238 (N_18238,N_17842,N_17693);
nor U18239 (N_18239,N_17976,N_17784);
xor U18240 (N_18240,N_17683,N_17636);
nor U18241 (N_18241,N_17744,N_17945);
xnor U18242 (N_18242,N_17893,N_17757);
xnor U18243 (N_18243,N_17834,N_17667);
and U18244 (N_18244,N_17820,N_17796);
or U18245 (N_18245,N_17626,N_17879);
nand U18246 (N_18246,N_17993,N_17734);
and U18247 (N_18247,N_17937,N_17796);
nor U18248 (N_18248,N_17840,N_17832);
and U18249 (N_18249,N_17897,N_17694);
nor U18250 (N_18250,N_17929,N_17730);
nor U18251 (N_18251,N_17957,N_17863);
and U18252 (N_18252,N_17608,N_17652);
xor U18253 (N_18253,N_17785,N_17739);
xor U18254 (N_18254,N_17987,N_17662);
nor U18255 (N_18255,N_17612,N_17752);
nand U18256 (N_18256,N_17963,N_17750);
xor U18257 (N_18257,N_17852,N_17682);
xor U18258 (N_18258,N_17667,N_17618);
nand U18259 (N_18259,N_17672,N_17787);
nor U18260 (N_18260,N_17913,N_17886);
and U18261 (N_18261,N_17993,N_17933);
or U18262 (N_18262,N_17910,N_17752);
nor U18263 (N_18263,N_17932,N_17821);
xnor U18264 (N_18264,N_17873,N_17805);
nor U18265 (N_18265,N_17957,N_17664);
or U18266 (N_18266,N_17676,N_17867);
or U18267 (N_18267,N_17977,N_17609);
and U18268 (N_18268,N_17758,N_17971);
xor U18269 (N_18269,N_17623,N_17851);
nand U18270 (N_18270,N_17726,N_17933);
and U18271 (N_18271,N_17792,N_17754);
nand U18272 (N_18272,N_17718,N_17827);
or U18273 (N_18273,N_17986,N_17840);
nor U18274 (N_18274,N_17885,N_17801);
nand U18275 (N_18275,N_17941,N_17885);
or U18276 (N_18276,N_17870,N_17638);
or U18277 (N_18277,N_17643,N_17666);
xor U18278 (N_18278,N_17736,N_17929);
nand U18279 (N_18279,N_17906,N_17974);
nand U18280 (N_18280,N_17814,N_17956);
or U18281 (N_18281,N_17651,N_17988);
or U18282 (N_18282,N_17778,N_17620);
nand U18283 (N_18283,N_17857,N_17681);
xnor U18284 (N_18284,N_17730,N_17871);
nand U18285 (N_18285,N_17665,N_17811);
or U18286 (N_18286,N_17642,N_17902);
xnor U18287 (N_18287,N_17644,N_17897);
nand U18288 (N_18288,N_17611,N_17978);
nor U18289 (N_18289,N_17719,N_17606);
nand U18290 (N_18290,N_17702,N_17674);
nor U18291 (N_18291,N_17691,N_17820);
nand U18292 (N_18292,N_17880,N_17928);
nor U18293 (N_18293,N_17994,N_17814);
nand U18294 (N_18294,N_17760,N_17720);
nand U18295 (N_18295,N_17993,N_17875);
xor U18296 (N_18296,N_17622,N_17951);
nor U18297 (N_18297,N_17904,N_17612);
nor U18298 (N_18298,N_17910,N_17930);
or U18299 (N_18299,N_17871,N_17913);
xor U18300 (N_18300,N_17805,N_17809);
and U18301 (N_18301,N_17701,N_17744);
and U18302 (N_18302,N_17949,N_17996);
or U18303 (N_18303,N_17842,N_17972);
nand U18304 (N_18304,N_17801,N_17997);
or U18305 (N_18305,N_17779,N_17642);
xnor U18306 (N_18306,N_17811,N_17881);
or U18307 (N_18307,N_17613,N_17802);
and U18308 (N_18308,N_17921,N_17937);
and U18309 (N_18309,N_17983,N_17668);
or U18310 (N_18310,N_17663,N_17657);
and U18311 (N_18311,N_17649,N_17624);
or U18312 (N_18312,N_17913,N_17777);
nand U18313 (N_18313,N_17616,N_17861);
nor U18314 (N_18314,N_17747,N_17787);
or U18315 (N_18315,N_17622,N_17718);
nand U18316 (N_18316,N_17971,N_17873);
and U18317 (N_18317,N_17801,N_17836);
xnor U18318 (N_18318,N_17861,N_17726);
and U18319 (N_18319,N_17900,N_17928);
and U18320 (N_18320,N_17776,N_17662);
nand U18321 (N_18321,N_17761,N_17762);
or U18322 (N_18322,N_17801,N_17720);
xor U18323 (N_18323,N_17914,N_17892);
nor U18324 (N_18324,N_17739,N_17765);
and U18325 (N_18325,N_17647,N_17707);
or U18326 (N_18326,N_17723,N_17616);
or U18327 (N_18327,N_17652,N_17627);
or U18328 (N_18328,N_17871,N_17906);
or U18329 (N_18329,N_17857,N_17912);
and U18330 (N_18330,N_17924,N_17662);
xor U18331 (N_18331,N_17960,N_17924);
xnor U18332 (N_18332,N_17804,N_17671);
or U18333 (N_18333,N_17845,N_17703);
xnor U18334 (N_18334,N_17806,N_17836);
nand U18335 (N_18335,N_17618,N_17648);
or U18336 (N_18336,N_17762,N_17874);
or U18337 (N_18337,N_17872,N_17621);
xnor U18338 (N_18338,N_17924,N_17995);
or U18339 (N_18339,N_17629,N_17902);
nand U18340 (N_18340,N_17943,N_17756);
and U18341 (N_18341,N_17998,N_17815);
nand U18342 (N_18342,N_17978,N_17691);
nor U18343 (N_18343,N_17897,N_17804);
and U18344 (N_18344,N_17886,N_17998);
or U18345 (N_18345,N_17710,N_17937);
or U18346 (N_18346,N_17649,N_17930);
nor U18347 (N_18347,N_17805,N_17715);
xnor U18348 (N_18348,N_17749,N_17652);
and U18349 (N_18349,N_17925,N_17680);
nor U18350 (N_18350,N_17796,N_17888);
or U18351 (N_18351,N_17972,N_17731);
and U18352 (N_18352,N_17608,N_17977);
nor U18353 (N_18353,N_17981,N_17922);
nor U18354 (N_18354,N_17911,N_17742);
nand U18355 (N_18355,N_17667,N_17603);
or U18356 (N_18356,N_17766,N_17837);
nand U18357 (N_18357,N_17810,N_17825);
nor U18358 (N_18358,N_17758,N_17781);
or U18359 (N_18359,N_17825,N_17984);
nand U18360 (N_18360,N_17770,N_17960);
or U18361 (N_18361,N_17760,N_17966);
xor U18362 (N_18362,N_17752,N_17679);
or U18363 (N_18363,N_17933,N_17999);
nor U18364 (N_18364,N_17974,N_17653);
or U18365 (N_18365,N_17795,N_17672);
nor U18366 (N_18366,N_17916,N_17713);
or U18367 (N_18367,N_17839,N_17638);
and U18368 (N_18368,N_17824,N_17859);
nand U18369 (N_18369,N_17972,N_17600);
nand U18370 (N_18370,N_17750,N_17882);
and U18371 (N_18371,N_17883,N_17764);
and U18372 (N_18372,N_17848,N_17960);
or U18373 (N_18373,N_17765,N_17728);
or U18374 (N_18374,N_17728,N_17986);
and U18375 (N_18375,N_17961,N_17819);
nor U18376 (N_18376,N_17760,N_17992);
xor U18377 (N_18377,N_17663,N_17926);
nand U18378 (N_18378,N_17612,N_17930);
and U18379 (N_18379,N_17659,N_17815);
or U18380 (N_18380,N_17998,N_17897);
nor U18381 (N_18381,N_17837,N_17870);
nand U18382 (N_18382,N_17718,N_17962);
xor U18383 (N_18383,N_17672,N_17819);
nand U18384 (N_18384,N_17993,N_17683);
nand U18385 (N_18385,N_17921,N_17760);
or U18386 (N_18386,N_17769,N_17975);
nor U18387 (N_18387,N_17654,N_17751);
nor U18388 (N_18388,N_17857,N_17876);
nand U18389 (N_18389,N_17897,N_17816);
nor U18390 (N_18390,N_17661,N_17610);
nand U18391 (N_18391,N_17862,N_17781);
and U18392 (N_18392,N_17913,N_17943);
nand U18393 (N_18393,N_17762,N_17983);
xnor U18394 (N_18394,N_17746,N_17975);
or U18395 (N_18395,N_17672,N_17984);
or U18396 (N_18396,N_17849,N_17733);
nor U18397 (N_18397,N_17976,N_17768);
or U18398 (N_18398,N_17910,N_17787);
nand U18399 (N_18399,N_17838,N_17756);
and U18400 (N_18400,N_18166,N_18082);
nor U18401 (N_18401,N_18185,N_18372);
nand U18402 (N_18402,N_18022,N_18306);
or U18403 (N_18403,N_18282,N_18289);
nor U18404 (N_18404,N_18340,N_18333);
xor U18405 (N_18405,N_18154,N_18172);
nor U18406 (N_18406,N_18115,N_18277);
and U18407 (N_18407,N_18267,N_18347);
and U18408 (N_18408,N_18018,N_18205);
and U18409 (N_18409,N_18396,N_18009);
nand U18410 (N_18410,N_18157,N_18011);
or U18411 (N_18411,N_18091,N_18352);
and U18412 (N_18412,N_18094,N_18376);
xor U18413 (N_18413,N_18032,N_18005);
nand U18414 (N_18414,N_18109,N_18153);
or U18415 (N_18415,N_18084,N_18040);
xnor U18416 (N_18416,N_18268,N_18211);
and U18417 (N_18417,N_18142,N_18042);
xnor U18418 (N_18418,N_18139,N_18353);
nor U18419 (N_18419,N_18390,N_18100);
or U18420 (N_18420,N_18138,N_18290);
or U18421 (N_18421,N_18370,N_18252);
xor U18422 (N_18422,N_18328,N_18055);
xnor U18423 (N_18423,N_18046,N_18304);
nor U18424 (N_18424,N_18341,N_18335);
nor U18425 (N_18425,N_18300,N_18285);
xor U18426 (N_18426,N_18116,N_18024);
nor U18427 (N_18427,N_18065,N_18044);
nor U18428 (N_18428,N_18284,N_18035);
nand U18429 (N_18429,N_18201,N_18127);
nor U18430 (N_18430,N_18010,N_18229);
or U18431 (N_18431,N_18113,N_18363);
or U18432 (N_18432,N_18008,N_18243);
or U18433 (N_18433,N_18398,N_18129);
xnor U18434 (N_18434,N_18192,N_18253);
or U18435 (N_18435,N_18150,N_18235);
or U18436 (N_18436,N_18274,N_18021);
nand U18437 (N_18437,N_18312,N_18118);
or U18438 (N_18438,N_18336,N_18356);
and U18439 (N_18439,N_18343,N_18198);
nor U18440 (N_18440,N_18119,N_18206);
nor U18441 (N_18441,N_18251,N_18240);
nor U18442 (N_18442,N_18393,N_18384);
nor U18443 (N_18443,N_18278,N_18088);
nor U18444 (N_18444,N_18069,N_18310);
nor U18445 (N_18445,N_18231,N_18379);
nor U18446 (N_18446,N_18388,N_18123);
nand U18447 (N_18447,N_18230,N_18258);
xor U18448 (N_18448,N_18080,N_18216);
nor U18449 (N_18449,N_18074,N_18107);
and U18450 (N_18450,N_18193,N_18015);
or U18451 (N_18451,N_18199,N_18238);
xor U18452 (N_18452,N_18339,N_18190);
nand U18453 (N_18453,N_18215,N_18232);
nor U18454 (N_18454,N_18257,N_18359);
nor U18455 (N_18455,N_18381,N_18355);
nor U18456 (N_18456,N_18093,N_18124);
or U18457 (N_18457,N_18038,N_18125);
xnor U18458 (N_18458,N_18334,N_18034);
or U18459 (N_18459,N_18027,N_18162);
nor U18460 (N_18460,N_18176,N_18320);
nand U18461 (N_18461,N_18283,N_18006);
xnor U18462 (N_18462,N_18095,N_18313);
nor U18463 (N_18463,N_18323,N_18121);
and U18464 (N_18464,N_18383,N_18303);
nor U18465 (N_18465,N_18371,N_18259);
nand U18466 (N_18466,N_18148,N_18007);
and U18467 (N_18467,N_18332,N_18321);
and U18468 (N_18468,N_18087,N_18030);
nor U18469 (N_18469,N_18067,N_18322);
and U18470 (N_18470,N_18077,N_18296);
and U18471 (N_18471,N_18203,N_18064);
nor U18472 (N_18472,N_18308,N_18264);
xor U18473 (N_18473,N_18063,N_18291);
nand U18474 (N_18474,N_18218,N_18365);
nor U18475 (N_18475,N_18319,N_18213);
xnor U18476 (N_18476,N_18221,N_18210);
xnor U18477 (N_18477,N_18337,N_18292);
xnor U18478 (N_18478,N_18047,N_18098);
xnor U18479 (N_18479,N_18207,N_18019);
nand U18480 (N_18480,N_18182,N_18177);
nand U18481 (N_18481,N_18362,N_18137);
nor U18482 (N_18482,N_18023,N_18307);
nor U18483 (N_18483,N_18373,N_18146);
nor U18484 (N_18484,N_18220,N_18163);
nor U18485 (N_18485,N_18317,N_18208);
nand U18486 (N_18486,N_18255,N_18126);
nand U18487 (N_18487,N_18299,N_18070);
nor U18488 (N_18488,N_18263,N_18085);
or U18489 (N_18489,N_18271,N_18043);
or U18490 (N_18490,N_18059,N_18342);
nor U18491 (N_18491,N_18066,N_18288);
xor U18492 (N_18492,N_18227,N_18103);
and U18493 (N_18493,N_18228,N_18256);
xnor U18494 (N_18494,N_18349,N_18394);
or U18495 (N_18495,N_18078,N_18195);
nor U18496 (N_18496,N_18265,N_18245);
or U18497 (N_18497,N_18302,N_18244);
and U18498 (N_18498,N_18212,N_18375);
nor U18499 (N_18499,N_18097,N_18382);
nor U18500 (N_18500,N_18366,N_18387);
xor U18501 (N_18501,N_18287,N_18017);
nor U18502 (N_18502,N_18294,N_18311);
nor U18503 (N_18503,N_18392,N_18073);
nand U18504 (N_18504,N_18112,N_18060);
nor U18505 (N_18505,N_18187,N_18135);
xor U18506 (N_18506,N_18039,N_18189);
and U18507 (N_18507,N_18036,N_18068);
xor U18508 (N_18508,N_18037,N_18051);
nand U18509 (N_18509,N_18086,N_18298);
or U18510 (N_18510,N_18001,N_18314);
or U18511 (N_18511,N_18378,N_18071);
xor U18512 (N_18512,N_18133,N_18262);
or U18513 (N_18513,N_18083,N_18297);
nand U18514 (N_18514,N_18248,N_18062);
nor U18515 (N_18515,N_18367,N_18161);
nor U18516 (N_18516,N_18101,N_18058);
nand U18517 (N_18517,N_18013,N_18266);
nand U18518 (N_18518,N_18076,N_18305);
xnor U18519 (N_18519,N_18000,N_18186);
nand U18520 (N_18520,N_18075,N_18241);
xnor U18521 (N_18521,N_18270,N_18226);
nor U18522 (N_18522,N_18134,N_18145);
and U18523 (N_18523,N_18102,N_18397);
nor U18524 (N_18524,N_18130,N_18079);
and U18525 (N_18525,N_18175,N_18316);
and U18526 (N_18526,N_18194,N_18260);
nand U18527 (N_18527,N_18279,N_18159);
xor U18528 (N_18528,N_18269,N_18250);
nand U18529 (N_18529,N_18170,N_18164);
nand U18530 (N_18530,N_18049,N_18181);
or U18531 (N_18531,N_18196,N_18089);
and U18532 (N_18532,N_18108,N_18167);
and U18533 (N_18533,N_18016,N_18180);
or U18534 (N_18534,N_18217,N_18204);
and U18535 (N_18535,N_18151,N_18272);
nand U18536 (N_18536,N_18143,N_18057);
nand U18537 (N_18537,N_18053,N_18160);
xor U18538 (N_18538,N_18106,N_18152);
nor U18539 (N_18539,N_18357,N_18338);
nand U18540 (N_18540,N_18351,N_18179);
or U18541 (N_18541,N_18155,N_18399);
and U18542 (N_18542,N_18045,N_18056);
or U18543 (N_18543,N_18004,N_18234);
xor U18544 (N_18544,N_18276,N_18233);
nand U18545 (N_18545,N_18033,N_18090);
and U18546 (N_18546,N_18389,N_18149);
nor U18547 (N_18547,N_18326,N_18131);
xnor U18548 (N_18548,N_18325,N_18295);
or U18549 (N_18549,N_18041,N_18012);
or U18550 (N_18550,N_18318,N_18224);
xnor U18551 (N_18551,N_18377,N_18242);
nand U18552 (N_18552,N_18246,N_18183);
xor U18553 (N_18553,N_18197,N_18368);
nor U18554 (N_18554,N_18141,N_18081);
nand U18555 (N_18555,N_18280,N_18354);
nor U18556 (N_18556,N_18165,N_18391);
or U18557 (N_18557,N_18050,N_18140);
or U18558 (N_18558,N_18344,N_18031);
xor U18559 (N_18559,N_18222,N_18360);
and U18560 (N_18560,N_18395,N_18169);
xor U18561 (N_18561,N_18324,N_18315);
and U18562 (N_18562,N_18117,N_18003);
xnor U18563 (N_18563,N_18184,N_18136);
and U18564 (N_18564,N_18358,N_18329);
nand U18565 (N_18565,N_18330,N_18114);
nor U18566 (N_18566,N_18249,N_18099);
nor U18567 (N_18567,N_18369,N_18188);
and U18568 (N_18568,N_18293,N_18092);
xnor U18569 (N_18569,N_18219,N_18209);
nor U18570 (N_18570,N_18029,N_18380);
xor U18571 (N_18571,N_18301,N_18054);
and U18572 (N_18572,N_18239,N_18025);
nand U18573 (N_18573,N_18026,N_18147);
xor U18574 (N_18574,N_18104,N_18122);
nand U18575 (N_18575,N_18200,N_18132);
nand U18576 (N_18576,N_18111,N_18156);
nor U18577 (N_18577,N_18158,N_18128);
xnor U18578 (N_18578,N_18275,N_18171);
or U18579 (N_18579,N_18002,N_18237);
or U18580 (N_18580,N_18173,N_18168);
nand U18581 (N_18581,N_18028,N_18374);
or U18582 (N_18582,N_18236,N_18309);
or U18583 (N_18583,N_18223,N_18214);
and U18584 (N_18584,N_18385,N_18364);
and U18585 (N_18585,N_18061,N_18191);
nor U18586 (N_18586,N_18072,N_18020);
xnor U18587 (N_18587,N_18254,N_18386);
and U18588 (N_18588,N_18225,N_18202);
nand U18589 (N_18589,N_18174,N_18273);
or U18590 (N_18590,N_18247,N_18110);
xnor U18591 (N_18591,N_18052,N_18331);
nand U18592 (N_18592,N_18281,N_18361);
or U18593 (N_18593,N_18327,N_18120);
nand U18594 (N_18594,N_18014,N_18144);
xnor U18595 (N_18595,N_18105,N_18346);
nand U18596 (N_18596,N_18345,N_18096);
or U18597 (N_18597,N_18350,N_18286);
and U18598 (N_18598,N_18261,N_18178);
xnor U18599 (N_18599,N_18348,N_18048);
and U18600 (N_18600,N_18389,N_18068);
nor U18601 (N_18601,N_18073,N_18060);
and U18602 (N_18602,N_18255,N_18253);
and U18603 (N_18603,N_18310,N_18381);
nand U18604 (N_18604,N_18233,N_18137);
or U18605 (N_18605,N_18053,N_18345);
nor U18606 (N_18606,N_18007,N_18233);
or U18607 (N_18607,N_18396,N_18258);
xor U18608 (N_18608,N_18188,N_18259);
nor U18609 (N_18609,N_18134,N_18278);
and U18610 (N_18610,N_18001,N_18220);
nand U18611 (N_18611,N_18020,N_18016);
and U18612 (N_18612,N_18232,N_18140);
or U18613 (N_18613,N_18256,N_18310);
xor U18614 (N_18614,N_18372,N_18358);
xor U18615 (N_18615,N_18361,N_18042);
or U18616 (N_18616,N_18224,N_18043);
nor U18617 (N_18617,N_18194,N_18151);
nand U18618 (N_18618,N_18152,N_18295);
nor U18619 (N_18619,N_18185,N_18271);
nand U18620 (N_18620,N_18171,N_18220);
and U18621 (N_18621,N_18326,N_18348);
nand U18622 (N_18622,N_18382,N_18211);
nand U18623 (N_18623,N_18398,N_18286);
xor U18624 (N_18624,N_18358,N_18198);
or U18625 (N_18625,N_18192,N_18342);
or U18626 (N_18626,N_18140,N_18338);
or U18627 (N_18627,N_18279,N_18140);
nor U18628 (N_18628,N_18299,N_18322);
nor U18629 (N_18629,N_18367,N_18181);
and U18630 (N_18630,N_18051,N_18073);
nor U18631 (N_18631,N_18034,N_18071);
nor U18632 (N_18632,N_18152,N_18101);
nand U18633 (N_18633,N_18388,N_18031);
nor U18634 (N_18634,N_18349,N_18157);
nor U18635 (N_18635,N_18202,N_18192);
nand U18636 (N_18636,N_18017,N_18166);
and U18637 (N_18637,N_18079,N_18280);
xnor U18638 (N_18638,N_18330,N_18015);
or U18639 (N_18639,N_18034,N_18219);
nand U18640 (N_18640,N_18352,N_18330);
nand U18641 (N_18641,N_18011,N_18012);
or U18642 (N_18642,N_18351,N_18106);
and U18643 (N_18643,N_18129,N_18302);
or U18644 (N_18644,N_18236,N_18182);
and U18645 (N_18645,N_18187,N_18363);
xnor U18646 (N_18646,N_18353,N_18282);
or U18647 (N_18647,N_18146,N_18067);
and U18648 (N_18648,N_18302,N_18333);
nand U18649 (N_18649,N_18279,N_18275);
or U18650 (N_18650,N_18387,N_18076);
or U18651 (N_18651,N_18310,N_18042);
nand U18652 (N_18652,N_18279,N_18163);
xnor U18653 (N_18653,N_18135,N_18207);
nor U18654 (N_18654,N_18164,N_18304);
or U18655 (N_18655,N_18242,N_18222);
or U18656 (N_18656,N_18189,N_18355);
nand U18657 (N_18657,N_18076,N_18087);
xor U18658 (N_18658,N_18113,N_18352);
nor U18659 (N_18659,N_18364,N_18145);
or U18660 (N_18660,N_18313,N_18363);
nand U18661 (N_18661,N_18384,N_18158);
nor U18662 (N_18662,N_18154,N_18106);
and U18663 (N_18663,N_18355,N_18343);
or U18664 (N_18664,N_18353,N_18336);
nor U18665 (N_18665,N_18336,N_18015);
or U18666 (N_18666,N_18289,N_18077);
and U18667 (N_18667,N_18353,N_18200);
and U18668 (N_18668,N_18065,N_18346);
or U18669 (N_18669,N_18072,N_18157);
or U18670 (N_18670,N_18291,N_18239);
and U18671 (N_18671,N_18144,N_18269);
and U18672 (N_18672,N_18115,N_18086);
nand U18673 (N_18673,N_18291,N_18358);
nor U18674 (N_18674,N_18347,N_18353);
nor U18675 (N_18675,N_18185,N_18058);
xor U18676 (N_18676,N_18211,N_18397);
nor U18677 (N_18677,N_18227,N_18137);
and U18678 (N_18678,N_18101,N_18040);
nand U18679 (N_18679,N_18142,N_18058);
nand U18680 (N_18680,N_18004,N_18030);
nor U18681 (N_18681,N_18116,N_18331);
xnor U18682 (N_18682,N_18059,N_18379);
nor U18683 (N_18683,N_18355,N_18216);
xor U18684 (N_18684,N_18133,N_18006);
and U18685 (N_18685,N_18149,N_18038);
nand U18686 (N_18686,N_18242,N_18071);
or U18687 (N_18687,N_18114,N_18286);
xor U18688 (N_18688,N_18220,N_18232);
or U18689 (N_18689,N_18083,N_18292);
or U18690 (N_18690,N_18276,N_18361);
nor U18691 (N_18691,N_18164,N_18038);
or U18692 (N_18692,N_18263,N_18320);
xnor U18693 (N_18693,N_18335,N_18047);
nor U18694 (N_18694,N_18244,N_18164);
nand U18695 (N_18695,N_18112,N_18137);
or U18696 (N_18696,N_18391,N_18340);
or U18697 (N_18697,N_18383,N_18353);
and U18698 (N_18698,N_18362,N_18337);
nor U18699 (N_18699,N_18159,N_18019);
xor U18700 (N_18700,N_18347,N_18286);
nor U18701 (N_18701,N_18178,N_18061);
xor U18702 (N_18702,N_18254,N_18109);
nand U18703 (N_18703,N_18347,N_18349);
nand U18704 (N_18704,N_18321,N_18006);
or U18705 (N_18705,N_18087,N_18101);
and U18706 (N_18706,N_18253,N_18206);
xor U18707 (N_18707,N_18327,N_18344);
nand U18708 (N_18708,N_18382,N_18316);
xor U18709 (N_18709,N_18234,N_18028);
nor U18710 (N_18710,N_18181,N_18237);
xor U18711 (N_18711,N_18279,N_18065);
nand U18712 (N_18712,N_18345,N_18291);
or U18713 (N_18713,N_18351,N_18329);
xnor U18714 (N_18714,N_18354,N_18384);
xnor U18715 (N_18715,N_18388,N_18276);
or U18716 (N_18716,N_18257,N_18260);
or U18717 (N_18717,N_18270,N_18173);
or U18718 (N_18718,N_18208,N_18332);
and U18719 (N_18719,N_18250,N_18335);
nor U18720 (N_18720,N_18069,N_18223);
nor U18721 (N_18721,N_18398,N_18003);
xnor U18722 (N_18722,N_18051,N_18341);
or U18723 (N_18723,N_18316,N_18317);
nor U18724 (N_18724,N_18308,N_18112);
and U18725 (N_18725,N_18001,N_18054);
and U18726 (N_18726,N_18104,N_18008);
nor U18727 (N_18727,N_18211,N_18321);
nor U18728 (N_18728,N_18146,N_18217);
nor U18729 (N_18729,N_18154,N_18320);
nor U18730 (N_18730,N_18305,N_18125);
nor U18731 (N_18731,N_18248,N_18317);
and U18732 (N_18732,N_18353,N_18382);
and U18733 (N_18733,N_18085,N_18150);
nor U18734 (N_18734,N_18207,N_18233);
xor U18735 (N_18735,N_18238,N_18239);
or U18736 (N_18736,N_18042,N_18163);
or U18737 (N_18737,N_18201,N_18037);
or U18738 (N_18738,N_18148,N_18253);
nor U18739 (N_18739,N_18265,N_18262);
and U18740 (N_18740,N_18218,N_18123);
nor U18741 (N_18741,N_18304,N_18141);
or U18742 (N_18742,N_18321,N_18220);
nand U18743 (N_18743,N_18181,N_18379);
nor U18744 (N_18744,N_18203,N_18220);
and U18745 (N_18745,N_18342,N_18171);
xor U18746 (N_18746,N_18173,N_18361);
and U18747 (N_18747,N_18055,N_18107);
or U18748 (N_18748,N_18201,N_18307);
or U18749 (N_18749,N_18271,N_18136);
xnor U18750 (N_18750,N_18276,N_18087);
or U18751 (N_18751,N_18011,N_18168);
or U18752 (N_18752,N_18315,N_18206);
nand U18753 (N_18753,N_18313,N_18242);
and U18754 (N_18754,N_18133,N_18223);
xnor U18755 (N_18755,N_18385,N_18136);
and U18756 (N_18756,N_18097,N_18172);
nand U18757 (N_18757,N_18341,N_18176);
xnor U18758 (N_18758,N_18383,N_18064);
nand U18759 (N_18759,N_18199,N_18118);
or U18760 (N_18760,N_18293,N_18244);
nand U18761 (N_18761,N_18366,N_18024);
xor U18762 (N_18762,N_18183,N_18032);
xor U18763 (N_18763,N_18028,N_18379);
nand U18764 (N_18764,N_18009,N_18322);
nor U18765 (N_18765,N_18170,N_18244);
xor U18766 (N_18766,N_18347,N_18295);
xor U18767 (N_18767,N_18349,N_18060);
xnor U18768 (N_18768,N_18021,N_18194);
nor U18769 (N_18769,N_18162,N_18251);
nand U18770 (N_18770,N_18392,N_18164);
or U18771 (N_18771,N_18220,N_18055);
and U18772 (N_18772,N_18021,N_18358);
or U18773 (N_18773,N_18263,N_18252);
nand U18774 (N_18774,N_18249,N_18133);
and U18775 (N_18775,N_18067,N_18098);
xnor U18776 (N_18776,N_18060,N_18220);
and U18777 (N_18777,N_18009,N_18330);
nand U18778 (N_18778,N_18366,N_18338);
nand U18779 (N_18779,N_18183,N_18363);
and U18780 (N_18780,N_18124,N_18306);
nand U18781 (N_18781,N_18101,N_18235);
and U18782 (N_18782,N_18287,N_18359);
xnor U18783 (N_18783,N_18172,N_18030);
nor U18784 (N_18784,N_18067,N_18090);
and U18785 (N_18785,N_18336,N_18066);
xnor U18786 (N_18786,N_18253,N_18210);
nor U18787 (N_18787,N_18224,N_18056);
xor U18788 (N_18788,N_18383,N_18200);
nor U18789 (N_18789,N_18018,N_18160);
or U18790 (N_18790,N_18186,N_18323);
and U18791 (N_18791,N_18326,N_18278);
or U18792 (N_18792,N_18159,N_18238);
or U18793 (N_18793,N_18159,N_18141);
or U18794 (N_18794,N_18061,N_18132);
xor U18795 (N_18795,N_18034,N_18067);
nand U18796 (N_18796,N_18339,N_18292);
or U18797 (N_18797,N_18181,N_18052);
or U18798 (N_18798,N_18328,N_18053);
nand U18799 (N_18799,N_18063,N_18253);
and U18800 (N_18800,N_18726,N_18584);
and U18801 (N_18801,N_18784,N_18592);
or U18802 (N_18802,N_18744,N_18568);
xor U18803 (N_18803,N_18670,N_18580);
xnor U18804 (N_18804,N_18732,N_18415);
nor U18805 (N_18805,N_18721,N_18658);
nand U18806 (N_18806,N_18677,N_18542);
or U18807 (N_18807,N_18579,N_18432);
xnor U18808 (N_18808,N_18761,N_18451);
nor U18809 (N_18809,N_18668,N_18434);
and U18810 (N_18810,N_18619,N_18782);
nor U18811 (N_18811,N_18679,N_18735);
and U18812 (N_18812,N_18541,N_18591);
xor U18813 (N_18813,N_18609,N_18763);
and U18814 (N_18814,N_18714,N_18509);
nor U18815 (N_18815,N_18689,N_18643);
or U18816 (N_18816,N_18758,N_18773);
nor U18817 (N_18817,N_18479,N_18687);
and U18818 (N_18818,N_18659,N_18532);
nor U18819 (N_18819,N_18661,N_18565);
nand U18820 (N_18820,N_18752,N_18406);
or U18821 (N_18821,N_18620,N_18740);
nand U18822 (N_18822,N_18555,N_18738);
or U18823 (N_18823,N_18711,N_18443);
and U18824 (N_18824,N_18540,N_18460);
xor U18825 (N_18825,N_18422,N_18666);
nor U18826 (N_18826,N_18582,N_18446);
or U18827 (N_18827,N_18767,N_18690);
or U18828 (N_18828,N_18458,N_18583);
nor U18829 (N_18829,N_18790,N_18543);
nand U18830 (N_18830,N_18742,N_18627);
xnor U18831 (N_18831,N_18611,N_18483);
or U18832 (N_18832,N_18786,N_18548);
nand U18833 (N_18833,N_18599,N_18707);
and U18834 (N_18834,N_18577,N_18510);
and U18835 (N_18835,N_18400,N_18547);
nor U18836 (N_18836,N_18696,N_18553);
xnor U18837 (N_18837,N_18589,N_18678);
nand U18838 (N_18838,N_18745,N_18566);
or U18839 (N_18839,N_18657,N_18475);
nand U18840 (N_18840,N_18642,N_18667);
and U18841 (N_18841,N_18676,N_18675);
nand U18842 (N_18842,N_18777,N_18533);
nor U18843 (N_18843,N_18724,N_18424);
nand U18844 (N_18844,N_18612,N_18426);
nand U18845 (N_18845,N_18720,N_18640);
and U18846 (N_18846,N_18454,N_18606);
nor U18847 (N_18847,N_18603,N_18794);
xnor U18848 (N_18848,N_18420,N_18428);
xor U18849 (N_18849,N_18755,N_18710);
nor U18850 (N_18850,N_18470,N_18605);
nor U18851 (N_18851,N_18438,N_18537);
xor U18852 (N_18852,N_18671,N_18455);
nor U18853 (N_18853,N_18445,N_18713);
or U18854 (N_18854,N_18636,N_18594);
nor U18855 (N_18855,N_18536,N_18481);
xnor U18856 (N_18856,N_18504,N_18461);
and U18857 (N_18857,N_18703,N_18762);
and U18858 (N_18858,N_18550,N_18493);
nand U18859 (N_18859,N_18515,N_18650);
nor U18860 (N_18860,N_18476,N_18512);
nor U18861 (N_18861,N_18549,N_18608);
or U18862 (N_18862,N_18474,N_18746);
xor U18863 (N_18863,N_18754,N_18465);
nor U18864 (N_18864,N_18647,N_18495);
or U18865 (N_18865,N_18558,N_18625);
nor U18866 (N_18866,N_18665,N_18792);
and U18867 (N_18867,N_18712,N_18523);
and U18868 (N_18868,N_18616,N_18576);
and U18869 (N_18869,N_18598,N_18624);
and U18870 (N_18870,N_18440,N_18688);
and U18871 (N_18871,N_18575,N_18638);
xor U18872 (N_18872,N_18596,N_18748);
and U18873 (N_18873,N_18405,N_18613);
nand U18874 (N_18874,N_18663,N_18653);
nand U18875 (N_18875,N_18702,N_18453);
or U18876 (N_18876,N_18519,N_18718);
or U18877 (N_18877,N_18545,N_18501);
or U18878 (N_18878,N_18567,N_18681);
or U18879 (N_18879,N_18435,N_18494);
or U18880 (N_18880,N_18750,N_18514);
or U18881 (N_18881,N_18564,N_18680);
and U18882 (N_18882,N_18631,N_18645);
nor U18883 (N_18883,N_18441,N_18634);
nand U18884 (N_18884,N_18705,N_18448);
and U18885 (N_18885,N_18499,N_18516);
nor U18886 (N_18886,N_18795,N_18462);
xor U18887 (N_18887,N_18587,N_18772);
or U18888 (N_18888,N_18464,N_18478);
nor U18889 (N_18889,N_18528,N_18684);
or U18890 (N_18890,N_18651,N_18730);
xor U18891 (N_18891,N_18734,N_18507);
nor U18892 (N_18892,N_18496,N_18753);
nor U18893 (N_18893,N_18569,N_18601);
nand U18894 (N_18894,N_18637,N_18517);
nand U18895 (N_18895,N_18610,N_18433);
nand U18896 (N_18896,N_18563,N_18708);
xor U18897 (N_18897,N_18437,N_18429);
xnor U18898 (N_18898,N_18595,N_18488);
and U18899 (N_18899,N_18655,N_18442);
nor U18900 (N_18900,N_18449,N_18685);
xnor U18901 (N_18901,N_18602,N_18469);
or U18902 (N_18902,N_18467,N_18617);
xor U18903 (N_18903,N_18492,N_18572);
and U18904 (N_18904,N_18502,N_18779);
nand U18905 (N_18905,N_18737,N_18739);
xnor U18906 (N_18906,N_18692,N_18444);
xor U18907 (N_18907,N_18717,N_18704);
and U18908 (N_18908,N_18403,N_18747);
and U18909 (N_18909,N_18497,N_18412);
nor U18910 (N_18910,N_18673,N_18546);
nor U18911 (N_18911,N_18471,N_18503);
or U18912 (N_18912,N_18628,N_18559);
xnor U18913 (N_18913,N_18622,N_18505);
nor U18914 (N_18914,N_18725,N_18418);
xnor U18915 (N_18915,N_18425,N_18538);
and U18916 (N_18916,N_18727,N_18522);
and U18917 (N_18917,N_18551,N_18588);
xor U18918 (N_18918,N_18459,N_18452);
nand U18919 (N_18919,N_18401,N_18656);
and U18920 (N_18920,N_18529,N_18796);
or U18921 (N_18921,N_18633,N_18527);
nand U18922 (N_18922,N_18506,N_18785);
nor U18923 (N_18923,N_18783,N_18694);
nor U18924 (N_18924,N_18757,N_18485);
nand U18925 (N_18925,N_18780,N_18581);
nor U18926 (N_18926,N_18654,N_18427);
or U18927 (N_18927,N_18423,N_18788);
nor U18928 (N_18928,N_18408,N_18430);
xnor U18929 (N_18929,N_18554,N_18770);
nand U18930 (N_18930,N_18562,N_18604);
or U18931 (N_18931,N_18662,N_18719);
or U18932 (N_18932,N_18741,N_18614);
and U18933 (N_18933,N_18781,N_18669);
and U18934 (N_18934,N_18706,N_18729);
nor U18935 (N_18935,N_18701,N_18530);
nand U18936 (N_18936,N_18477,N_18644);
and U18937 (N_18937,N_18556,N_18695);
xor U18938 (N_18938,N_18693,N_18728);
xor U18939 (N_18939,N_18574,N_18799);
or U18940 (N_18940,N_18743,N_18402);
and U18941 (N_18941,N_18570,N_18674);
nand U18942 (N_18942,N_18463,N_18797);
nand U18943 (N_18943,N_18411,N_18491);
and U18944 (N_18944,N_18544,N_18766);
and U18945 (N_18945,N_18760,N_18646);
nand U18946 (N_18946,N_18586,N_18749);
or U18947 (N_18947,N_18552,N_18736);
or U18948 (N_18948,N_18447,N_18699);
nand U18949 (N_18949,N_18722,N_18539);
xor U18950 (N_18950,N_18487,N_18416);
nand U18951 (N_18951,N_18793,N_18791);
or U18952 (N_18952,N_18578,N_18571);
or U18953 (N_18953,N_18421,N_18526);
or U18954 (N_18954,N_18561,N_18649);
and U18955 (N_18955,N_18404,N_18431);
or U18956 (N_18956,N_18626,N_18630);
or U18957 (N_18957,N_18511,N_18798);
nand U18958 (N_18958,N_18641,N_18716);
or U18959 (N_18959,N_18607,N_18660);
and U18960 (N_18960,N_18490,N_18531);
xnor U18961 (N_18961,N_18414,N_18664);
nor U18962 (N_18962,N_18618,N_18407);
nand U18963 (N_18963,N_18520,N_18486);
or U18964 (N_18964,N_18776,N_18417);
or U18965 (N_18965,N_18573,N_18751);
or U18966 (N_18966,N_18733,N_18629);
and U18967 (N_18967,N_18723,N_18764);
or U18968 (N_18968,N_18632,N_18436);
or U18969 (N_18969,N_18700,N_18525);
nor U18970 (N_18970,N_18450,N_18648);
and U18971 (N_18971,N_18731,N_18652);
or U18972 (N_18972,N_18489,N_18557);
and U18973 (N_18973,N_18789,N_18419);
or U18974 (N_18974,N_18778,N_18535);
xnor U18975 (N_18975,N_18410,N_18682);
xnor U18976 (N_18976,N_18639,N_18524);
nand U18977 (N_18977,N_18683,N_18756);
nor U18978 (N_18978,N_18590,N_18484);
nor U18979 (N_18979,N_18771,N_18508);
nand U18980 (N_18980,N_18709,N_18472);
nor U18981 (N_18981,N_18621,N_18769);
nor U18982 (N_18982,N_18765,N_18686);
nor U18983 (N_18983,N_18456,N_18597);
and U18984 (N_18984,N_18691,N_18473);
nand U18985 (N_18985,N_18498,N_18534);
or U18986 (N_18986,N_18715,N_18560);
nor U18987 (N_18987,N_18768,N_18635);
xnor U18988 (N_18988,N_18521,N_18513);
and U18989 (N_18989,N_18593,N_18518);
or U18990 (N_18990,N_18759,N_18774);
nand U18991 (N_18991,N_18468,N_18457);
or U18992 (N_18992,N_18413,N_18697);
nand U18993 (N_18993,N_18480,N_18672);
nor U18994 (N_18994,N_18500,N_18482);
and U18995 (N_18995,N_18585,N_18409);
nor U18996 (N_18996,N_18787,N_18466);
nand U18997 (N_18997,N_18439,N_18775);
nand U18998 (N_18998,N_18600,N_18623);
xor U18999 (N_18999,N_18698,N_18615);
or U19000 (N_19000,N_18666,N_18483);
or U19001 (N_19001,N_18759,N_18620);
nand U19002 (N_19002,N_18459,N_18468);
xnor U19003 (N_19003,N_18660,N_18699);
nor U19004 (N_19004,N_18797,N_18675);
and U19005 (N_19005,N_18487,N_18402);
nor U19006 (N_19006,N_18770,N_18526);
nand U19007 (N_19007,N_18682,N_18721);
and U19008 (N_19008,N_18795,N_18487);
xnor U19009 (N_19009,N_18489,N_18754);
or U19010 (N_19010,N_18445,N_18411);
nor U19011 (N_19011,N_18509,N_18540);
nor U19012 (N_19012,N_18465,N_18691);
or U19013 (N_19013,N_18478,N_18511);
nand U19014 (N_19014,N_18791,N_18407);
or U19015 (N_19015,N_18796,N_18589);
nand U19016 (N_19016,N_18732,N_18458);
or U19017 (N_19017,N_18546,N_18716);
xor U19018 (N_19018,N_18575,N_18407);
or U19019 (N_19019,N_18739,N_18407);
xnor U19020 (N_19020,N_18444,N_18670);
xor U19021 (N_19021,N_18534,N_18615);
and U19022 (N_19022,N_18474,N_18603);
nand U19023 (N_19023,N_18441,N_18425);
nand U19024 (N_19024,N_18554,N_18602);
nor U19025 (N_19025,N_18451,N_18418);
nand U19026 (N_19026,N_18645,N_18606);
nand U19027 (N_19027,N_18728,N_18437);
nor U19028 (N_19028,N_18555,N_18778);
xor U19029 (N_19029,N_18732,N_18717);
nand U19030 (N_19030,N_18466,N_18749);
and U19031 (N_19031,N_18775,N_18688);
and U19032 (N_19032,N_18738,N_18609);
nand U19033 (N_19033,N_18454,N_18433);
xnor U19034 (N_19034,N_18679,N_18463);
xnor U19035 (N_19035,N_18701,N_18590);
and U19036 (N_19036,N_18544,N_18535);
or U19037 (N_19037,N_18746,N_18464);
nand U19038 (N_19038,N_18508,N_18590);
or U19039 (N_19039,N_18492,N_18743);
nand U19040 (N_19040,N_18719,N_18417);
and U19041 (N_19041,N_18693,N_18442);
xor U19042 (N_19042,N_18484,N_18630);
and U19043 (N_19043,N_18414,N_18666);
or U19044 (N_19044,N_18408,N_18697);
nor U19045 (N_19045,N_18655,N_18798);
or U19046 (N_19046,N_18489,N_18527);
or U19047 (N_19047,N_18483,N_18491);
or U19048 (N_19048,N_18585,N_18416);
nand U19049 (N_19049,N_18767,N_18748);
nand U19050 (N_19050,N_18748,N_18677);
nor U19051 (N_19051,N_18796,N_18430);
xor U19052 (N_19052,N_18414,N_18615);
xor U19053 (N_19053,N_18690,N_18669);
nor U19054 (N_19054,N_18764,N_18672);
xnor U19055 (N_19055,N_18493,N_18599);
nand U19056 (N_19056,N_18588,N_18484);
or U19057 (N_19057,N_18761,N_18746);
nand U19058 (N_19058,N_18547,N_18534);
or U19059 (N_19059,N_18661,N_18634);
xnor U19060 (N_19060,N_18437,N_18745);
nor U19061 (N_19061,N_18709,N_18467);
and U19062 (N_19062,N_18607,N_18400);
nor U19063 (N_19063,N_18471,N_18501);
or U19064 (N_19064,N_18712,N_18522);
nor U19065 (N_19065,N_18769,N_18417);
nor U19066 (N_19066,N_18773,N_18605);
or U19067 (N_19067,N_18652,N_18560);
xnor U19068 (N_19068,N_18484,N_18768);
and U19069 (N_19069,N_18663,N_18765);
and U19070 (N_19070,N_18671,N_18767);
nand U19071 (N_19071,N_18524,N_18648);
nand U19072 (N_19072,N_18586,N_18462);
and U19073 (N_19073,N_18427,N_18725);
nand U19074 (N_19074,N_18626,N_18612);
nand U19075 (N_19075,N_18477,N_18466);
nand U19076 (N_19076,N_18687,N_18777);
xor U19077 (N_19077,N_18571,N_18416);
nand U19078 (N_19078,N_18432,N_18789);
nor U19079 (N_19079,N_18429,N_18640);
and U19080 (N_19080,N_18418,N_18509);
xnor U19081 (N_19081,N_18681,N_18620);
nor U19082 (N_19082,N_18703,N_18783);
and U19083 (N_19083,N_18769,N_18464);
or U19084 (N_19084,N_18778,N_18464);
nor U19085 (N_19085,N_18638,N_18643);
or U19086 (N_19086,N_18442,N_18494);
xnor U19087 (N_19087,N_18754,N_18747);
and U19088 (N_19088,N_18554,N_18433);
nand U19089 (N_19089,N_18660,N_18784);
or U19090 (N_19090,N_18732,N_18663);
and U19091 (N_19091,N_18691,N_18439);
xnor U19092 (N_19092,N_18650,N_18753);
nand U19093 (N_19093,N_18459,N_18438);
and U19094 (N_19094,N_18733,N_18676);
nor U19095 (N_19095,N_18745,N_18747);
or U19096 (N_19096,N_18643,N_18611);
or U19097 (N_19097,N_18578,N_18659);
xnor U19098 (N_19098,N_18757,N_18631);
and U19099 (N_19099,N_18411,N_18798);
or U19100 (N_19100,N_18748,N_18438);
xor U19101 (N_19101,N_18441,N_18655);
nand U19102 (N_19102,N_18598,N_18462);
or U19103 (N_19103,N_18479,N_18525);
and U19104 (N_19104,N_18701,N_18547);
or U19105 (N_19105,N_18772,N_18663);
and U19106 (N_19106,N_18590,N_18538);
xor U19107 (N_19107,N_18797,N_18468);
and U19108 (N_19108,N_18410,N_18685);
xnor U19109 (N_19109,N_18566,N_18795);
and U19110 (N_19110,N_18724,N_18774);
xnor U19111 (N_19111,N_18571,N_18679);
nand U19112 (N_19112,N_18558,N_18786);
xnor U19113 (N_19113,N_18718,N_18483);
nand U19114 (N_19114,N_18637,N_18444);
xnor U19115 (N_19115,N_18684,N_18511);
nand U19116 (N_19116,N_18665,N_18776);
xor U19117 (N_19117,N_18709,N_18587);
nand U19118 (N_19118,N_18602,N_18646);
nand U19119 (N_19119,N_18436,N_18715);
xor U19120 (N_19120,N_18714,N_18541);
and U19121 (N_19121,N_18725,N_18645);
or U19122 (N_19122,N_18723,N_18647);
nor U19123 (N_19123,N_18780,N_18564);
nor U19124 (N_19124,N_18665,N_18434);
or U19125 (N_19125,N_18449,N_18751);
and U19126 (N_19126,N_18418,N_18549);
nand U19127 (N_19127,N_18428,N_18532);
nor U19128 (N_19128,N_18418,N_18642);
and U19129 (N_19129,N_18780,N_18592);
and U19130 (N_19130,N_18424,N_18766);
nor U19131 (N_19131,N_18471,N_18707);
xnor U19132 (N_19132,N_18766,N_18551);
nand U19133 (N_19133,N_18539,N_18729);
or U19134 (N_19134,N_18447,N_18458);
and U19135 (N_19135,N_18490,N_18516);
or U19136 (N_19136,N_18784,N_18698);
xnor U19137 (N_19137,N_18727,N_18789);
xnor U19138 (N_19138,N_18409,N_18442);
xnor U19139 (N_19139,N_18759,N_18797);
nand U19140 (N_19140,N_18701,N_18768);
xor U19141 (N_19141,N_18756,N_18703);
xnor U19142 (N_19142,N_18486,N_18419);
xor U19143 (N_19143,N_18666,N_18442);
xnor U19144 (N_19144,N_18560,N_18577);
xor U19145 (N_19145,N_18734,N_18790);
and U19146 (N_19146,N_18451,N_18720);
xor U19147 (N_19147,N_18616,N_18665);
nand U19148 (N_19148,N_18505,N_18428);
nor U19149 (N_19149,N_18540,N_18514);
nor U19150 (N_19150,N_18552,N_18570);
xor U19151 (N_19151,N_18418,N_18721);
or U19152 (N_19152,N_18418,N_18416);
or U19153 (N_19153,N_18525,N_18449);
or U19154 (N_19154,N_18600,N_18678);
nor U19155 (N_19155,N_18560,N_18616);
nor U19156 (N_19156,N_18607,N_18575);
nor U19157 (N_19157,N_18570,N_18516);
nor U19158 (N_19158,N_18493,N_18404);
nand U19159 (N_19159,N_18424,N_18638);
nand U19160 (N_19160,N_18461,N_18667);
nand U19161 (N_19161,N_18554,N_18774);
and U19162 (N_19162,N_18561,N_18526);
nand U19163 (N_19163,N_18620,N_18499);
xor U19164 (N_19164,N_18635,N_18563);
xor U19165 (N_19165,N_18778,N_18716);
xor U19166 (N_19166,N_18571,N_18701);
nand U19167 (N_19167,N_18759,N_18549);
and U19168 (N_19168,N_18553,N_18699);
nand U19169 (N_19169,N_18709,N_18689);
or U19170 (N_19170,N_18663,N_18551);
nand U19171 (N_19171,N_18491,N_18496);
or U19172 (N_19172,N_18485,N_18750);
xor U19173 (N_19173,N_18581,N_18404);
nor U19174 (N_19174,N_18545,N_18626);
xor U19175 (N_19175,N_18663,N_18403);
xnor U19176 (N_19176,N_18435,N_18731);
and U19177 (N_19177,N_18450,N_18765);
and U19178 (N_19178,N_18493,N_18772);
and U19179 (N_19179,N_18405,N_18633);
nor U19180 (N_19180,N_18538,N_18629);
nor U19181 (N_19181,N_18647,N_18584);
nand U19182 (N_19182,N_18566,N_18450);
and U19183 (N_19183,N_18647,N_18709);
or U19184 (N_19184,N_18594,N_18568);
nor U19185 (N_19185,N_18515,N_18511);
xnor U19186 (N_19186,N_18798,N_18733);
nor U19187 (N_19187,N_18602,N_18566);
nand U19188 (N_19188,N_18765,N_18746);
nor U19189 (N_19189,N_18438,N_18647);
nor U19190 (N_19190,N_18595,N_18638);
nor U19191 (N_19191,N_18469,N_18440);
nor U19192 (N_19192,N_18552,N_18612);
nor U19193 (N_19193,N_18585,N_18754);
and U19194 (N_19194,N_18661,N_18450);
nand U19195 (N_19195,N_18570,N_18456);
nor U19196 (N_19196,N_18709,N_18726);
xnor U19197 (N_19197,N_18411,N_18737);
nand U19198 (N_19198,N_18480,N_18579);
xor U19199 (N_19199,N_18655,N_18731);
and U19200 (N_19200,N_19129,N_19100);
nor U19201 (N_19201,N_18833,N_18825);
nand U19202 (N_19202,N_19119,N_18859);
or U19203 (N_19203,N_19011,N_19038);
nor U19204 (N_19204,N_18900,N_18856);
nand U19205 (N_19205,N_19024,N_18801);
xor U19206 (N_19206,N_19001,N_19145);
xnor U19207 (N_19207,N_19182,N_18849);
or U19208 (N_19208,N_19142,N_19097);
xnor U19209 (N_19209,N_19177,N_18938);
or U19210 (N_19210,N_19081,N_18803);
xor U19211 (N_19211,N_18926,N_19149);
nor U19212 (N_19212,N_18884,N_19108);
nor U19213 (N_19213,N_19076,N_19186);
and U19214 (N_19214,N_19103,N_18818);
nor U19215 (N_19215,N_18934,N_19066);
nor U19216 (N_19216,N_19137,N_18930);
xnor U19217 (N_19217,N_19075,N_19049);
xor U19218 (N_19218,N_18872,N_18921);
and U19219 (N_19219,N_18890,N_19150);
nor U19220 (N_19220,N_19164,N_18946);
xor U19221 (N_19221,N_19092,N_19087);
nand U19222 (N_19222,N_18901,N_19102);
nor U19223 (N_19223,N_18980,N_19190);
xnor U19224 (N_19224,N_18911,N_19062);
and U19225 (N_19225,N_18875,N_18916);
xnor U19226 (N_19226,N_19130,N_18808);
xor U19227 (N_19227,N_18919,N_19163);
nand U19228 (N_19228,N_18909,N_19157);
nor U19229 (N_19229,N_18958,N_18999);
nand U19230 (N_19230,N_19135,N_19156);
nand U19231 (N_19231,N_19016,N_19029);
nor U19232 (N_19232,N_18943,N_19060);
nand U19233 (N_19233,N_19197,N_18972);
and U19234 (N_19234,N_19140,N_19065);
xnor U19235 (N_19235,N_19046,N_19041);
or U19236 (N_19236,N_19008,N_18983);
nor U19237 (N_19237,N_19078,N_19159);
nor U19238 (N_19238,N_19055,N_19032);
xnor U19239 (N_19239,N_19193,N_18874);
nor U19240 (N_19240,N_19125,N_19005);
xor U19241 (N_19241,N_18932,N_19187);
or U19242 (N_19242,N_19117,N_19199);
nand U19243 (N_19243,N_19014,N_19086);
nand U19244 (N_19244,N_18809,N_19059);
and U19245 (N_19245,N_18893,N_18853);
nor U19246 (N_19246,N_18997,N_18965);
and U19247 (N_19247,N_18877,N_19120);
nand U19248 (N_19248,N_19124,N_18894);
and U19249 (N_19249,N_18827,N_18941);
nand U19250 (N_19250,N_19183,N_19138);
and U19251 (N_19251,N_19002,N_18804);
or U19252 (N_19252,N_18981,N_19000);
nand U19253 (N_19253,N_19180,N_19147);
nand U19254 (N_19254,N_18954,N_19198);
and U19255 (N_19255,N_18903,N_19143);
or U19256 (N_19256,N_18918,N_19171);
xnor U19257 (N_19257,N_19044,N_18881);
nor U19258 (N_19258,N_19185,N_19162);
and U19259 (N_19259,N_18913,N_18993);
or U19260 (N_19260,N_19084,N_19184);
and U19261 (N_19261,N_19074,N_18865);
and U19262 (N_19262,N_19173,N_19152);
nand U19263 (N_19263,N_19175,N_18952);
or U19264 (N_19264,N_19111,N_18840);
xor U19265 (N_19265,N_18824,N_18889);
nand U19266 (N_19266,N_19045,N_18984);
or U19267 (N_19267,N_18908,N_19015);
or U19268 (N_19268,N_18848,N_19189);
nor U19269 (N_19269,N_18988,N_19088);
or U19270 (N_19270,N_19082,N_19007);
nand U19271 (N_19271,N_18979,N_18845);
xor U19272 (N_19272,N_19118,N_18977);
xnor U19273 (N_19273,N_19027,N_18936);
xor U19274 (N_19274,N_18867,N_18844);
nand U19275 (N_19275,N_19099,N_18857);
nor U19276 (N_19276,N_18986,N_19192);
and U19277 (N_19277,N_18923,N_18895);
nor U19278 (N_19278,N_18960,N_19020);
and U19279 (N_19279,N_19121,N_19047);
nand U19280 (N_19280,N_19158,N_18974);
and U19281 (N_19281,N_18951,N_18950);
xor U19282 (N_19282,N_18937,N_19035);
xnor U19283 (N_19283,N_18998,N_19096);
nand U19284 (N_19284,N_18886,N_19191);
nand U19285 (N_19285,N_19188,N_18800);
nor U19286 (N_19286,N_18870,N_18817);
nand U19287 (N_19287,N_18805,N_18969);
or U19288 (N_19288,N_18996,N_18878);
and U19289 (N_19289,N_18846,N_18994);
nand U19290 (N_19290,N_18975,N_19141);
nor U19291 (N_19291,N_18802,N_19028);
nor U19292 (N_19292,N_19160,N_19018);
and U19293 (N_19293,N_19128,N_19181);
xor U19294 (N_19294,N_18892,N_19053);
nor U19295 (N_19295,N_18907,N_19110);
xor U19296 (N_19296,N_19168,N_18822);
or U19297 (N_19297,N_18957,N_19042);
nor U19298 (N_19298,N_19022,N_19132);
nand U19299 (N_19299,N_19107,N_19133);
or U19300 (N_19300,N_19048,N_18953);
nor U19301 (N_19301,N_18873,N_18855);
nand U19302 (N_19302,N_19079,N_19095);
xor U19303 (N_19303,N_19073,N_18862);
nand U19304 (N_19304,N_19179,N_18968);
and U19305 (N_19305,N_18929,N_18842);
nand U19306 (N_19306,N_18815,N_18905);
and U19307 (N_19307,N_19051,N_19104);
nor U19308 (N_19308,N_18869,N_18902);
or U19309 (N_19309,N_19021,N_18864);
nand U19310 (N_19310,N_18876,N_18990);
or U19311 (N_19311,N_18962,N_19054);
nand U19312 (N_19312,N_18854,N_18832);
xor U19313 (N_19313,N_18863,N_18806);
nor U19314 (N_19314,N_18971,N_19167);
nand U19315 (N_19315,N_18959,N_18834);
xnor U19316 (N_19316,N_19040,N_19064);
and U19317 (N_19317,N_18879,N_18924);
nor U19318 (N_19318,N_18917,N_19112);
nand U19319 (N_19319,N_19089,N_19052);
nand U19320 (N_19320,N_18920,N_19113);
nor U19321 (N_19321,N_18826,N_18807);
nand U19322 (N_19322,N_18871,N_19127);
and U19323 (N_19323,N_18987,N_18899);
xnor U19324 (N_19324,N_18811,N_18847);
xnor U19325 (N_19325,N_19116,N_19067);
and U19326 (N_19326,N_19036,N_19169);
and U19327 (N_19327,N_19172,N_19126);
nor U19328 (N_19328,N_19037,N_19004);
and U19329 (N_19329,N_18830,N_19056);
or U19330 (N_19330,N_19148,N_18922);
or U19331 (N_19331,N_18897,N_19165);
xor U19332 (N_19332,N_18939,N_19039);
xnor U19333 (N_19333,N_19151,N_18944);
xor U19334 (N_19334,N_18963,N_19161);
nor U19335 (N_19335,N_19083,N_18810);
nor U19336 (N_19336,N_19069,N_19043);
nand U19337 (N_19337,N_19134,N_19122);
nand U19338 (N_19338,N_19063,N_19033);
nor U19339 (N_19339,N_18821,N_19114);
and U19340 (N_19340,N_19106,N_18989);
nor U19341 (N_19341,N_19166,N_18882);
or U19342 (N_19342,N_18843,N_19072);
nor U19343 (N_19343,N_18914,N_19153);
nor U19344 (N_19344,N_18940,N_18888);
and U19345 (N_19345,N_18942,N_19023);
nor U19346 (N_19346,N_19058,N_18956);
nand U19347 (N_19347,N_19123,N_19061);
nor U19348 (N_19348,N_18906,N_18967);
or U19349 (N_19349,N_19006,N_18896);
xnor U19350 (N_19350,N_19105,N_18931);
xor U19351 (N_19351,N_18819,N_19090);
nand U19352 (N_19352,N_18992,N_18860);
or U19353 (N_19353,N_18891,N_18836);
nand U19354 (N_19354,N_19136,N_19091);
or U19355 (N_19355,N_19085,N_19070);
xnor U19356 (N_19356,N_18816,N_18928);
and U19357 (N_19357,N_19154,N_18828);
nor U19358 (N_19358,N_18955,N_19115);
nand U19359 (N_19359,N_18831,N_18883);
nor U19360 (N_19360,N_19196,N_18978);
or U19361 (N_19361,N_18904,N_18841);
xnor U19362 (N_19362,N_19109,N_18880);
nand U19363 (N_19363,N_18966,N_18982);
and U19364 (N_19364,N_18945,N_19025);
nor U19365 (N_19365,N_18868,N_18898);
nor U19366 (N_19366,N_19195,N_19017);
or U19367 (N_19367,N_18839,N_19194);
or U19368 (N_19368,N_18925,N_18820);
nor U19369 (N_19369,N_19093,N_19139);
nor U19370 (N_19370,N_18915,N_19131);
or U19371 (N_19371,N_18973,N_19050);
or U19372 (N_19372,N_18838,N_19098);
xnor U19373 (N_19373,N_19026,N_18829);
xnor U19374 (N_19374,N_19034,N_19170);
nor U19375 (N_19375,N_19010,N_18850);
nand U19376 (N_19376,N_19068,N_18948);
nor U19377 (N_19377,N_19012,N_19174);
nor U19378 (N_19378,N_18964,N_19071);
nand U19379 (N_19379,N_19019,N_18976);
and U19380 (N_19380,N_18837,N_18995);
xnor U19381 (N_19381,N_19101,N_19003);
nand U19382 (N_19382,N_18912,N_19077);
or U19383 (N_19383,N_18887,N_19146);
and U19384 (N_19384,N_19030,N_19057);
xnor U19385 (N_19385,N_19094,N_18823);
xor U19386 (N_19386,N_18991,N_18927);
or U19387 (N_19387,N_18866,N_19155);
and U19388 (N_19388,N_18852,N_18935);
xnor U19389 (N_19389,N_18985,N_19013);
xnor U19390 (N_19390,N_19080,N_18961);
nand U19391 (N_19391,N_18933,N_18814);
xnor U19392 (N_19392,N_19178,N_18812);
nor U19393 (N_19393,N_19009,N_18851);
nand U19394 (N_19394,N_18949,N_18835);
nand U19395 (N_19395,N_18861,N_18885);
nand U19396 (N_19396,N_18947,N_19031);
xor U19397 (N_19397,N_18970,N_19176);
nand U19398 (N_19398,N_18910,N_19144);
xnor U19399 (N_19399,N_18858,N_18813);
nor U19400 (N_19400,N_19043,N_18871);
or U19401 (N_19401,N_18943,N_18923);
nor U19402 (N_19402,N_18929,N_19026);
or U19403 (N_19403,N_19092,N_19099);
nand U19404 (N_19404,N_18849,N_19032);
nand U19405 (N_19405,N_19049,N_18956);
and U19406 (N_19406,N_19112,N_18800);
and U19407 (N_19407,N_18947,N_18957);
xnor U19408 (N_19408,N_19111,N_19152);
nor U19409 (N_19409,N_19036,N_18833);
nor U19410 (N_19410,N_18981,N_19014);
nand U19411 (N_19411,N_19026,N_19149);
or U19412 (N_19412,N_19088,N_18956);
nor U19413 (N_19413,N_18901,N_19197);
nor U19414 (N_19414,N_18883,N_18870);
or U19415 (N_19415,N_18902,N_19100);
or U19416 (N_19416,N_18803,N_18969);
xnor U19417 (N_19417,N_19089,N_19118);
nand U19418 (N_19418,N_18890,N_18842);
nor U19419 (N_19419,N_18998,N_18844);
or U19420 (N_19420,N_19170,N_19091);
xnor U19421 (N_19421,N_19137,N_19024);
nand U19422 (N_19422,N_18952,N_18967);
nor U19423 (N_19423,N_18886,N_18974);
nor U19424 (N_19424,N_19061,N_18957);
nor U19425 (N_19425,N_19168,N_18873);
or U19426 (N_19426,N_18841,N_19155);
nand U19427 (N_19427,N_19044,N_19164);
nand U19428 (N_19428,N_18940,N_19182);
xor U19429 (N_19429,N_19060,N_19058);
xnor U19430 (N_19430,N_19080,N_19005);
or U19431 (N_19431,N_18888,N_19098);
or U19432 (N_19432,N_19160,N_19046);
nor U19433 (N_19433,N_18812,N_19175);
xnor U19434 (N_19434,N_18808,N_18816);
xor U19435 (N_19435,N_18832,N_18836);
or U19436 (N_19436,N_18881,N_19061);
or U19437 (N_19437,N_19116,N_18978);
nor U19438 (N_19438,N_18800,N_18938);
xor U19439 (N_19439,N_18824,N_18965);
and U19440 (N_19440,N_18863,N_19102);
nor U19441 (N_19441,N_19129,N_19170);
xnor U19442 (N_19442,N_19105,N_18979);
xnor U19443 (N_19443,N_18898,N_18929);
nand U19444 (N_19444,N_19096,N_18961);
or U19445 (N_19445,N_18945,N_19196);
xnor U19446 (N_19446,N_19119,N_18940);
nor U19447 (N_19447,N_19008,N_18969);
and U19448 (N_19448,N_19178,N_19163);
and U19449 (N_19449,N_19030,N_19051);
nand U19450 (N_19450,N_19187,N_18977);
and U19451 (N_19451,N_19184,N_19038);
nor U19452 (N_19452,N_18866,N_18892);
nor U19453 (N_19453,N_19196,N_19002);
xor U19454 (N_19454,N_19122,N_19165);
nand U19455 (N_19455,N_19146,N_18998);
nand U19456 (N_19456,N_18875,N_19096);
xnor U19457 (N_19457,N_19083,N_19082);
or U19458 (N_19458,N_19166,N_18932);
nor U19459 (N_19459,N_19181,N_18872);
and U19460 (N_19460,N_19000,N_18996);
or U19461 (N_19461,N_18855,N_19017);
xnor U19462 (N_19462,N_18988,N_18868);
xor U19463 (N_19463,N_19028,N_19180);
and U19464 (N_19464,N_19165,N_19057);
xor U19465 (N_19465,N_18831,N_19005);
nor U19466 (N_19466,N_18898,N_19110);
nor U19467 (N_19467,N_19165,N_19102);
nand U19468 (N_19468,N_18872,N_19089);
nor U19469 (N_19469,N_19080,N_19131);
and U19470 (N_19470,N_19143,N_19176);
nor U19471 (N_19471,N_19170,N_19090);
or U19472 (N_19472,N_18810,N_18950);
nand U19473 (N_19473,N_19075,N_18812);
xor U19474 (N_19474,N_19037,N_18808);
xor U19475 (N_19475,N_19152,N_19138);
and U19476 (N_19476,N_18961,N_19057);
or U19477 (N_19477,N_18962,N_19138);
nand U19478 (N_19478,N_18881,N_19045);
nand U19479 (N_19479,N_18889,N_18968);
and U19480 (N_19480,N_19184,N_18997);
xor U19481 (N_19481,N_19120,N_19021);
nor U19482 (N_19482,N_18895,N_18988);
nor U19483 (N_19483,N_18801,N_18814);
xor U19484 (N_19484,N_18867,N_18935);
or U19485 (N_19485,N_19010,N_19082);
nand U19486 (N_19486,N_19168,N_19184);
xor U19487 (N_19487,N_19050,N_18912);
and U19488 (N_19488,N_18877,N_18976);
nand U19489 (N_19489,N_18842,N_18852);
nand U19490 (N_19490,N_19039,N_19064);
nand U19491 (N_19491,N_18992,N_19007);
or U19492 (N_19492,N_19178,N_18920);
nor U19493 (N_19493,N_19109,N_18838);
xnor U19494 (N_19494,N_19123,N_19159);
or U19495 (N_19495,N_18848,N_19102);
nand U19496 (N_19496,N_19060,N_19096);
nor U19497 (N_19497,N_19121,N_18922);
nand U19498 (N_19498,N_18957,N_18968);
nand U19499 (N_19499,N_18981,N_19122);
and U19500 (N_19500,N_19177,N_18819);
or U19501 (N_19501,N_19160,N_19118);
or U19502 (N_19502,N_18839,N_18942);
nand U19503 (N_19503,N_18892,N_19016);
nor U19504 (N_19504,N_18977,N_18846);
xor U19505 (N_19505,N_18943,N_19010);
nor U19506 (N_19506,N_19190,N_19149);
xnor U19507 (N_19507,N_18876,N_18853);
nand U19508 (N_19508,N_19049,N_19079);
xnor U19509 (N_19509,N_19059,N_18954);
nand U19510 (N_19510,N_19049,N_19174);
nand U19511 (N_19511,N_19137,N_19009);
nand U19512 (N_19512,N_19042,N_19089);
nor U19513 (N_19513,N_19127,N_18876);
nor U19514 (N_19514,N_19154,N_19168);
nand U19515 (N_19515,N_19184,N_18841);
nand U19516 (N_19516,N_19081,N_18962);
xnor U19517 (N_19517,N_18913,N_19191);
and U19518 (N_19518,N_18918,N_19003);
and U19519 (N_19519,N_19115,N_19024);
xnor U19520 (N_19520,N_19021,N_19003);
or U19521 (N_19521,N_19188,N_18939);
nand U19522 (N_19522,N_19176,N_19045);
nor U19523 (N_19523,N_18880,N_18972);
nor U19524 (N_19524,N_18901,N_19022);
xor U19525 (N_19525,N_18833,N_19110);
nand U19526 (N_19526,N_18851,N_18972);
and U19527 (N_19527,N_18828,N_19132);
nand U19528 (N_19528,N_18952,N_18964);
or U19529 (N_19529,N_19072,N_19105);
xor U19530 (N_19530,N_18808,N_18971);
nand U19531 (N_19531,N_18871,N_18925);
or U19532 (N_19532,N_18878,N_18875);
nand U19533 (N_19533,N_18994,N_19157);
nand U19534 (N_19534,N_18824,N_19187);
or U19535 (N_19535,N_18901,N_19065);
nand U19536 (N_19536,N_18945,N_18961);
nand U19537 (N_19537,N_19154,N_18911);
xnor U19538 (N_19538,N_18901,N_19036);
nand U19539 (N_19539,N_19181,N_19071);
or U19540 (N_19540,N_18860,N_18893);
and U19541 (N_19541,N_19190,N_18992);
or U19542 (N_19542,N_19162,N_19150);
or U19543 (N_19543,N_19049,N_18891);
nand U19544 (N_19544,N_18918,N_18851);
nand U19545 (N_19545,N_18934,N_18939);
xnor U19546 (N_19546,N_18935,N_18846);
or U19547 (N_19547,N_19053,N_18952);
xor U19548 (N_19548,N_19146,N_18925);
nor U19549 (N_19549,N_18814,N_19155);
or U19550 (N_19550,N_18920,N_18999);
xnor U19551 (N_19551,N_18856,N_19129);
nor U19552 (N_19552,N_18976,N_19015);
or U19553 (N_19553,N_19143,N_18926);
nor U19554 (N_19554,N_19026,N_18800);
nor U19555 (N_19555,N_18929,N_19151);
xor U19556 (N_19556,N_18839,N_19032);
xor U19557 (N_19557,N_18878,N_18867);
xor U19558 (N_19558,N_18897,N_19009);
nand U19559 (N_19559,N_18804,N_19119);
nor U19560 (N_19560,N_18963,N_18988);
and U19561 (N_19561,N_19158,N_18969);
nor U19562 (N_19562,N_19174,N_19120);
or U19563 (N_19563,N_18803,N_18819);
nand U19564 (N_19564,N_18925,N_18934);
nand U19565 (N_19565,N_18860,N_18864);
nand U19566 (N_19566,N_18853,N_18831);
and U19567 (N_19567,N_19100,N_19121);
nor U19568 (N_19568,N_18887,N_18820);
xnor U19569 (N_19569,N_18992,N_19048);
or U19570 (N_19570,N_19009,N_18926);
or U19571 (N_19571,N_19019,N_18857);
nor U19572 (N_19572,N_18824,N_19031);
nand U19573 (N_19573,N_19134,N_18958);
nand U19574 (N_19574,N_18834,N_19154);
nor U19575 (N_19575,N_18983,N_19142);
nand U19576 (N_19576,N_18863,N_18991);
or U19577 (N_19577,N_18946,N_19139);
nand U19578 (N_19578,N_18932,N_18896);
nand U19579 (N_19579,N_18827,N_19060);
and U19580 (N_19580,N_19023,N_18908);
and U19581 (N_19581,N_19199,N_18931);
nor U19582 (N_19582,N_19041,N_18872);
and U19583 (N_19583,N_18919,N_19117);
nand U19584 (N_19584,N_19166,N_19030);
or U19585 (N_19585,N_18936,N_19059);
and U19586 (N_19586,N_18899,N_19111);
and U19587 (N_19587,N_19088,N_18952);
and U19588 (N_19588,N_18938,N_19158);
nor U19589 (N_19589,N_18932,N_19067);
and U19590 (N_19590,N_18882,N_19198);
nand U19591 (N_19591,N_19015,N_18920);
nor U19592 (N_19592,N_18833,N_19102);
nor U19593 (N_19593,N_18883,N_18996);
xnor U19594 (N_19594,N_18920,N_18811);
xor U19595 (N_19595,N_18870,N_19040);
xor U19596 (N_19596,N_18997,N_19158);
or U19597 (N_19597,N_19057,N_19033);
or U19598 (N_19598,N_19131,N_18971);
and U19599 (N_19599,N_18884,N_18858);
or U19600 (N_19600,N_19569,N_19485);
nor U19601 (N_19601,N_19375,N_19216);
or U19602 (N_19602,N_19499,N_19361);
or U19603 (N_19603,N_19405,N_19565);
or U19604 (N_19604,N_19319,N_19278);
xor U19605 (N_19605,N_19433,N_19283);
or U19606 (N_19606,N_19312,N_19544);
nor U19607 (N_19607,N_19504,N_19310);
xnor U19608 (N_19608,N_19464,N_19462);
or U19609 (N_19609,N_19291,N_19223);
or U19610 (N_19610,N_19584,N_19437);
and U19611 (N_19611,N_19248,N_19335);
or U19612 (N_19612,N_19376,N_19436);
nand U19613 (N_19613,N_19556,N_19257);
nand U19614 (N_19614,N_19358,N_19261);
xor U19615 (N_19615,N_19457,N_19355);
nor U19616 (N_19616,N_19325,N_19262);
xor U19617 (N_19617,N_19545,N_19541);
nand U19618 (N_19618,N_19547,N_19435);
or U19619 (N_19619,N_19419,N_19525);
xnor U19620 (N_19620,N_19285,N_19532);
nand U19621 (N_19621,N_19593,N_19254);
or U19622 (N_19622,N_19482,N_19542);
nor U19623 (N_19623,N_19264,N_19299);
nand U19624 (N_19624,N_19377,N_19490);
nand U19625 (N_19625,N_19586,N_19200);
xor U19626 (N_19626,N_19587,N_19311);
or U19627 (N_19627,N_19566,N_19467);
nand U19628 (N_19628,N_19395,N_19445);
or U19629 (N_19629,N_19233,N_19511);
or U19630 (N_19630,N_19336,N_19468);
xor U19631 (N_19631,N_19480,N_19305);
xor U19632 (N_19632,N_19318,N_19364);
and U19633 (N_19633,N_19580,N_19362);
nand U19634 (N_19634,N_19380,N_19323);
xnor U19635 (N_19635,N_19409,N_19360);
and U19636 (N_19636,N_19507,N_19366);
nand U19637 (N_19637,N_19267,N_19501);
or U19638 (N_19638,N_19564,N_19347);
or U19639 (N_19639,N_19350,N_19241);
or U19640 (N_19640,N_19455,N_19222);
and U19641 (N_19641,N_19440,N_19372);
nor U19642 (N_19642,N_19270,N_19280);
xor U19643 (N_19643,N_19448,N_19263);
xor U19644 (N_19644,N_19210,N_19272);
or U19645 (N_19645,N_19406,N_19220);
xor U19646 (N_19646,N_19474,N_19416);
and U19647 (N_19647,N_19374,N_19450);
nor U19648 (N_19648,N_19337,N_19338);
and U19649 (N_19649,N_19522,N_19402);
nand U19650 (N_19650,N_19573,N_19424);
and U19651 (N_19651,N_19378,N_19316);
and U19652 (N_19652,N_19592,N_19255);
nor U19653 (N_19653,N_19492,N_19413);
and U19654 (N_19654,N_19290,N_19397);
nand U19655 (N_19655,N_19428,N_19206);
and U19656 (N_19656,N_19354,N_19313);
xnor U19657 (N_19657,N_19329,N_19326);
nor U19658 (N_19658,N_19208,N_19357);
or U19659 (N_19659,N_19275,N_19543);
or U19660 (N_19660,N_19389,N_19509);
xor U19661 (N_19661,N_19379,N_19598);
nand U19662 (N_19662,N_19595,N_19321);
and U19663 (N_19663,N_19351,N_19236);
xnor U19664 (N_19664,N_19562,N_19471);
xnor U19665 (N_19665,N_19552,N_19476);
xnor U19666 (N_19666,N_19568,N_19469);
or U19667 (N_19667,N_19317,N_19218);
xor U19668 (N_19668,N_19415,N_19591);
nand U19669 (N_19669,N_19286,N_19540);
nand U19670 (N_19670,N_19453,N_19237);
or U19671 (N_19671,N_19258,N_19201);
xor U19672 (N_19672,N_19211,N_19282);
xor U19673 (N_19673,N_19488,N_19230);
nand U19674 (N_19674,N_19596,N_19517);
or U19675 (N_19675,N_19212,N_19537);
and U19676 (N_19676,N_19266,N_19349);
xor U19677 (N_19677,N_19417,N_19470);
nand U19678 (N_19678,N_19473,N_19503);
or U19679 (N_19679,N_19268,N_19340);
xnor U19680 (N_19680,N_19363,N_19202);
nand U19681 (N_19681,N_19577,N_19232);
nand U19682 (N_19682,N_19253,N_19365);
and U19683 (N_19683,N_19369,N_19554);
nor U19684 (N_19684,N_19472,N_19400);
and U19685 (N_19685,N_19359,N_19439);
xnor U19686 (N_19686,N_19444,N_19486);
or U19687 (N_19687,N_19234,N_19520);
nor U19688 (N_19688,N_19570,N_19306);
nor U19689 (N_19689,N_19422,N_19259);
nor U19690 (N_19690,N_19500,N_19578);
xnor U19691 (N_19691,N_19381,N_19432);
xnor U19692 (N_19692,N_19459,N_19203);
nor U19693 (N_19693,N_19442,N_19226);
or U19694 (N_19694,N_19209,N_19399);
xnor U19695 (N_19695,N_19309,N_19583);
nor U19696 (N_19696,N_19224,N_19551);
nand U19697 (N_19697,N_19315,N_19599);
nor U19698 (N_19698,N_19597,N_19493);
xor U19699 (N_19699,N_19506,N_19465);
or U19700 (N_19700,N_19484,N_19523);
or U19701 (N_19701,N_19454,N_19301);
and U19702 (N_19702,N_19452,N_19243);
nor U19703 (N_19703,N_19303,N_19367);
nand U19704 (N_19704,N_19308,N_19461);
and U19705 (N_19705,N_19414,N_19271);
nor U19706 (N_19706,N_19341,N_19496);
nand U19707 (N_19707,N_19348,N_19478);
nand U19708 (N_19708,N_19518,N_19277);
xnor U19709 (N_19709,N_19487,N_19328);
xnor U19710 (N_19710,N_19494,N_19368);
and U19711 (N_19711,N_19585,N_19385);
nor U19712 (N_19712,N_19383,N_19590);
xnor U19713 (N_19713,N_19346,N_19456);
xnor U19714 (N_19714,N_19269,N_19449);
nand U19715 (N_19715,N_19524,N_19549);
or U19716 (N_19716,N_19535,N_19249);
or U19717 (N_19717,N_19332,N_19398);
or U19718 (N_19718,N_19307,N_19373);
and U19719 (N_19719,N_19557,N_19244);
and U19720 (N_19720,N_19434,N_19247);
nor U19721 (N_19721,N_19214,N_19466);
or U19722 (N_19722,N_19333,N_19294);
nor U19723 (N_19723,N_19371,N_19529);
nor U19724 (N_19724,N_19561,N_19527);
xor U19725 (N_19725,N_19219,N_19477);
or U19726 (N_19726,N_19563,N_19281);
nor U19727 (N_19727,N_19392,N_19429);
or U19728 (N_19728,N_19594,N_19297);
nor U19729 (N_19729,N_19582,N_19207);
or U19730 (N_19730,N_19238,N_19370);
nor U19731 (N_19731,N_19411,N_19327);
nand U19732 (N_19732,N_19251,N_19344);
xor U19733 (N_19733,N_19443,N_19403);
or U19734 (N_19734,N_19553,N_19495);
or U19735 (N_19735,N_19235,N_19412);
and U19736 (N_19736,N_19431,N_19546);
or U19737 (N_19737,N_19225,N_19528);
nor U19738 (N_19738,N_19571,N_19572);
and U19739 (N_19739,N_19284,N_19228);
xnor U19740 (N_19740,N_19205,N_19458);
nand U19741 (N_19741,N_19288,N_19300);
nor U19742 (N_19742,N_19555,N_19322);
nor U19743 (N_19743,N_19246,N_19276);
nand U19744 (N_19744,N_19293,N_19356);
xor U19745 (N_19745,N_19343,N_19531);
or U19746 (N_19746,N_19292,N_19215);
and U19747 (N_19747,N_19404,N_19491);
or U19748 (N_19748,N_19274,N_19388);
nor U19749 (N_19749,N_19229,N_19260);
or U19750 (N_19750,N_19289,N_19589);
nor U19751 (N_19751,N_19353,N_19302);
nand U19752 (N_19752,N_19221,N_19314);
or U19753 (N_19753,N_19386,N_19418);
and U19754 (N_19754,N_19483,N_19217);
xor U19755 (N_19755,N_19408,N_19256);
nand U19756 (N_19756,N_19463,N_19514);
or U19757 (N_19757,N_19387,N_19295);
xor U19758 (N_19758,N_19421,N_19451);
nor U19759 (N_19759,N_19550,N_19530);
nor U19760 (N_19760,N_19460,N_19245);
nor U19761 (N_19761,N_19426,N_19420);
and U19762 (N_19762,N_19512,N_19342);
xor U19763 (N_19763,N_19441,N_19489);
and U19764 (N_19764,N_19273,N_19324);
or U19765 (N_19765,N_19382,N_19533);
nor U19766 (N_19766,N_19250,N_19446);
nand U19767 (N_19767,N_19502,N_19567);
or U19768 (N_19768,N_19581,N_19239);
nand U19769 (N_19769,N_19558,N_19475);
xnor U19770 (N_19770,N_19265,N_19352);
xnor U19771 (N_19771,N_19391,N_19515);
and U19772 (N_19772,N_19213,N_19410);
and U19773 (N_19773,N_19345,N_19481);
nor U19774 (N_19774,N_19560,N_19479);
xor U19775 (N_19775,N_19394,N_19227);
and U19776 (N_19776,N_19279,N_19296);
and U19777 (N_19777,N_19498,N_19339);
nor U19778 (N_19778,N_19430,N_19510);
and U19779 (N_19779,N_19384,N_19576);
xor U19780 (N_19780,N_19539,N_19559);
nor U19781 (N_19781,N_19538,N_19536);
nor U19782 (N_19782,N_19401,N_19390);
xnor U19783 (N_19783,N_19588,N_19513);
nand U19784 (N_19784,N_19526,N_19505);
xnor U19785 (N_19785,N_19548,N_19579);
or U19786 (N_19786,N_19497,N_19574);
nor U19787 (N_19787,N_19304,N_19334);
nand U19788 (N_19788,N_19425,N_19330);
and U19789 (N_19789,N_19521,N_19423);
nand U19790 (N_19790,N_19331,N_19231);
nor U19791 (N_19791,N_19407,N_19438);
nor U19792 (N_19792,N_19204,N_19508);
and U19793 (N_19793,N_19298,N_19287);
or U19794 (N_19794,N_19320,N_19242);
or U19795 (N_19795,N_19447,N_19396);
nor U19796 (N_19796,N_19252,N_19516);
xor U19797 (N_19797,N_19393,N_19240);
and U19798 (N_19798,N_19575,N_19534);
nor U19799 (N_19799,N_19427,N_19519);
nand U19800 (N_19800,N_19232,N_19568);
and U19801 (N_19801,N_19434,N_19362);
or U19802 (N_19802,N_19314,N_19473);
xnor U19803 (N_19803,N_19337,N_19325);
nor U19804 (N_19804,N_19223,N_19467);
or U19805 (N_19805,N_19493,N_19338);
xor U19806 (N_19806,N_19444,N_19305);
nand U19807 (N_19807,N_19363,N_19315);
or U19808 (N_19808,N_19388,N_19363);
nand U19809 (N_19809,N_19409,N_19456);
xor U19810 (N_19810,N_19548,N_19438);
nand U19811 (N_19811,N_19435,N_19478);
and U19812 (N_19812,N_19535,N_19557);
nand U19813 (N_19813,N_19310,N_19306);
and U19814 (N_19814,N_19389,N_19342);
and U19815 (N_19815,N_19270,N_19498);
nand U19816 (N_19816,N_19326,N_19304);
nand U19817 (N_19817,N_19329,N_19495);
and U19818 (N_19818,N_19588,N_19512);
nor U19819 (N_19819,N_19294,N_19532);
and U19820 (N_19820,N_19246,N_19573);
nor U19821 (N_19821,N_19247,N_19572);
nand U19822 (N_19822,N_19312,N_19384);
xnor U19823 (N_19823,N_19524,N_19327);
or U19824 (N_19824,N_19219,N_19321);
or U19825 (N_19825,N_19494,N_19227);
nand U19826 (N_19826,N_19304,N_19216);
xnor U19827 (N_19827,N_19302,N_19347);
or U19828 (N_19828,N_19595,N_19499);
or U19829 (N_19829,N_19559,N_19466);
nor U19830 (N_19830,N_19402,N_19501);
and U19831 (N_19831,N_19293,N_19469);
nor U19832 (N_19832,N_19311,N_19213);
nor U19833 (N_19833,N_19418,N_19540);
or U19834 (N_19834,N_19319,N_19366);
xor U19835 (N_19835,N_19468,N_19271);
nor U19836 (N_19836,N_19339,N_19250);
xor U19837 (N_19837,N_19477,N_19444);
and U19838 (N_19838,N_19371,N_19264);
and U19839 (N_19839,N_19310,N_19545);
and U19840 (N_19840,N_19543,N_19464);
nand U19841 (N_19841,N_19297,N_19320);
nor U19842 (N_19842,N_19496,N_19538);
nand U19843 (N_19843,N_19470,N_19551);
or U19844 (N_19844,N_19200,N_19297);
nand U19845 (N_19845,N_19549,N_19485);
xnor U19846 (N_19846,N_19245,N_19445);
and U19847 (N_19847,N_19546,N_19434);
and U19848 (N_19848,N_19264,N_19495);
xnor U19849 (N_19849,N_19510,N_19495);
nor U19850 (N_19850,N_19452,N_19268);
nor U19851 (N_19851,N_19383,N_19341);
nor U19852 (N_19852,N_19415,N_19549);
or U19853 (N_19853,N_19567,N_19260);
nand U19854 (N_19854,N_19298,N_19456);
nand U19855 (N_19855,N_19314,N_19255);
or U19856 (N_19856,N_19210,N_19257);
xor U19857 (N_19857,N_19424,N_19437);
nand U19858 (N_19858,N_19344,N_19320);
nand U19859 (N_19859,N_19324,N_19477);
nand U19860 (N_19860,N_19322,N_19567);
nor U19861 (N_19861,N_19258,N_19257);
and U19862 (N_19862,N_19544,N_19434);
nor U19863 (N_19863,N_19563,N_19321);
nor U19864 (N_19864,N_19219,N_19452);
nor U19865 (N_19865,N_19341,N_19320);
nand U19866 (N_19866,N_19440,N_19201);
or U19867 (N_19867,N_19292,N_19284);
and U19868 (N_19868,N_19507,N_19465);
nor U19869 (N_19869,N_19406,N_19525);
nor U19870 (N_19870,N_19219,N_19274);
and U19871 (N_19871,N_19463,N_19352);
or U19872 (N_19872,N_19231,N_19471);
and U19873 (N_19873,N_19498,N_19458);
and U19874 (N_19874,N_19334,N_19413);
and U19875 (N_19875,N_19537,N_19563);
and U19876 (N_19876,N_19404,N_19493);
and U19877 (N_19877,N_19323,N_19202);
nand U19878 (N_19878,N_19367,N_19272);
xnor U19879 (N_19879,N_19336,N_19266);
nand U19880 (N_19880,N_19368,N_19203);
xnor U19881 (N_19881,N_19577,N_19204);
xor U19882 (N_19882,N_19490,N_19504);
nor U19883 (N_19883,N_19220,N_19367);
and U19884 (N_19884,N_19545,N_19579);
nand U19885 (N_19885,N_19371,N_19378);
nand U19886 (N_19886,N_19258,N_19207);
nand U19887 (N_19887,N_19520,N_19544);
xnor U19888 (N_19888,N_19259,N_19380);
or U19889 (N_19889,N_19552,N_19285);
and U19890 (N_19890,N_19315,N_19393);
nand U19891 (N_19891,N_19531,N_19347);
or U19892 (N_19892,N_19576,N_19586);
xnor U19893 (N_19893,N_19427,N_19565);
and U19894 (N_19894,N_19259,N_19208);
xnor U19895 (N_19895,N_19276,N_19473);
or U19896 (N_19896,N_19399,N_19234);
nor U19897 (N_19897,N_19263,N_19417);
xor U19898 (N_19898,N_19529,N_19271);
and U19899 (N_19899,N_19392,N_19536);
nand U19900 (N_19900,N_19560,N_19285);
nor U19901 (N_19901,N_19580,N_19208);
nand U19902 (N_19902,N_19464,N_19595);
and U19903 (N_19903,N_19271,N_19476);
xnor U19904 (N_19904,N_19524,N_19418);
nor U19905 (N_19905,N_19552,N_19514);
nand U19906 (N_19906,N_19258,N_19327);
and U19907 (N_19907,N_19587,N_19244);
or U19908 (N_19908,N_19403,N_19204);
or U19909 (N_19909,N_19274,N_19257);
nand U19910 (N_19910,N_19585,N_19398);
and U19911 (N_19911,N_19304,N_19537);
nor U19912 (N_19912,N_19492,N_19393);
xor U19913 (N_19913,N_19322,N_19269);
or U19914 (N_19914,N_19393,N_19417);
or U19915 (N_19915,N_19520,N_19511);
nor U19916 (N_19916,N_19271,N_19433);
or U19917 (N_19917,N_19533,N_19428);
or U19918 (N_19918,N_19582,N_19224);
and U19919 (N_19919,N_19512,N_19365);
or U19920 (N_19920,N_19278,N_19363);
and U19921 (N_19921,N_19308,N_19468);
nand U19922 (N_19922,N_19563,N_19278);
nor U19923 (N_19923,N_19447,N_19262);
nand U19924 (N_19924,N_19362,N_19530);
nor U19925 (N_19925,N_19429,N_19472);
nor U19926 (N_19926,N_19300,N_19489);
and U19927 (N_19927,N_19381,N_19565);
nor U19928 (N_19928,N_19362,N_19592);
or U19929 (N_19929,N_19462,N_19389);
or U19930 (N_19930,N_19223,N_19428);
xnor U19931 (N_19931,N_19561,N_19394);
nand U19932 (N_19932,N_19387,N_19584);
and U19933 (N_19933,N_19338,N_19457);
or U19934 (N_19934,N_19520,N_19236);
xor U19935 (N_19935,N_19591,N_19368);
nor U19936 (N_19936,N_19527,N_19409);
nand U19937 (N_19937,N_19243,N_19516);
or U19938 (N_19938,N_19545,N_19352);
xor U19939 (N_19939,N_19285,N_19238);
or U19940 (N_19940,N_19293,N_19538);
or U19941 (N_19941,N_19441,N_19342);
nand U19942 (N_19942,N_19402,N_19380);
xor U19943 (N_19943,N_19536,N_19207);
xnor U19944 (N_19944,N_19343,N_19597);
nand U19945 (N_19945,N_19360,N_19585);
and U19946 (N_19946,N_19300,N_19533);
and U19947 (N_19947,N_19390,N_19393);
and U19948 (N_19948,N_19459,N_19579);
nor U19949 (N_19949,N_19491,N_19486);
and U19950 (N_19950,N_19342,N_19530);
xor U19951 (N_19951,N_19488,N_19311);
or U19952 (N_19952,N_19563,N_19453);
and U19953 (N_19953,N_19318,N_19533);
and U19954 (N_19954,N_19240,N_19271);
or U19955 (N_19955,N_19363,N_19231);
or U19956 (N_19956,N_19532,N_19379);
nor U19957 (N_19957,N_19414,N_19200);
nand U19958 (N_19958,N_19421,N_19328);
nand U19959 (N_19959,N_19260,N_19458);
nand U19960 (N_19960,N_19515,N_19386);
or U19961 (N_19961,N_19226,N_19380);
xor U19962 (N_19962,N_19374,N_19552);
xor U19963 (N_19963,N_19403,N_19354);
and U19964 (N_19964,N_19474,N_19221);
xor U19965 (N_19965,N_19512,N_19231);
nor U19966 (N_19966,N_19201,N_19527);
nor U19967 (N_19967,N_19338,N_19221);
xor U19968 (N_19968,N_19577,N_19326);
nor U19969 (N_19969,N_19483,N_19544);
xnor U19970 (N_19970,N_19509,N_19458);
and U19971 (N_19971,N_19312,N_19411);
or U19972 (N_19972,N_19220,N_19576);
or U19973 (N_19973,N_19553,N_19396);
nand U19974 (N_19974,N_19443,N_19311);
nor U19975 (N_19975,N_19353,N_19439);
or U19976 (N_19976,N_19340,N_19332);
and U19977 (N_19977,N_19429,N_19335);
nand U19978 (N_19978,N_19551,N_19396);
and U19979 (N_19979,N_19442,N_19285);
or U19980 (N_19980,N_19557,N_19382);
or U19981 (N_19981,N_19320,N_19296);
or U19982 (N_19982,N_19459,N_19244);
nor U19983 (N_19983,N_19204,N_19465);
nor U19984 (N_19984,N_19238,N_19585);
xnor U19985 (N_19985,N_19314,N_19457);
xor U19986 (N_19986,N_19352,N_19377);
nor U19987 (N_19987,N_19464,N_19353);
nor U19988 (N_19988,N_19314,N_19480);
xnor U19989 (N_19989,N_19593,N_19292);
and U19990 (N_19990,N_19310,N_19383);
nand U19991 (N_19991,N_19480,N_19291);
nand U19992 (N_19992,N_19310,N_19349);
nor U19993 (N_19993,N_19410,N_19500);
and U19994 (N_19994,N_19357,N_19462);
nand U19995 (N_19995,N_19422,N_19421);
nor U19996 (N_19996,N_19488,N_19300);
nand U19997 (N_19997,N_19511,N_19210);
xor U19998 (N_19998,N_19580,N_19235);
nor U19999 (N_19999,N_19453,N_19536);
nand UO_0 (O_0,N_19870,N_19773);
nor UO_1 (O_1,N_19968,N_19992);
nor UO_2 (O_2,N_19643,N_19669);
nor UO_3 (O_3,N_19935,N_19829);
xor UO_4 (O_4,N_19993,N_19614);
nand UO_5 (O_5,N_19649,N_19952);
nand UO_6 (O_6,N_19705,N_19794);
xnor UO_7 (O_7,N_19792,N_19891);
or UO_8 (O_8,N_19977,N_19732);
nor UO_9 (O_9,N_19662,N_19898);
or UO_10 (O_10,N_19695,N_19927);
and UO_11 (O_11,N_19889,N_19668);
xor UO_12 (O_12,N_19802,N_19838);
and UO_13 (O_13,N_19890,N_19625);
and UO_14 (O_14,N_19951,N_19698);
nor UO_15 (O_15,N_19921,N_19896);
and UO_16 (O_16,N_19736,N_19756);
nand UO_17 (O_17,N_19758,N_19973);
nand UO_18 (O_18,N_19863,N_19928);
and UO_19 (O_19,N_19711,N_19623);
nand UO_20 (O_20,N_19855,N_19607);
nand UO_21 (O_21,N_19663,N_19634);
or UO_22 (O_22,N_19729,N_19801);
nor UO_23 (O_23,N_19965,N_19842);
xor UO_24 (O_24,N_19957,N_19866);
and UO_25 (O_25,N_19845,N_19856);
xnor UO_26 (O_26,N_19949,N_19804);
and UO_27 (O_27,N_19962,N_19657);
or UO_28 (O_28,N_19997,N_19721);
nor UO_29 (O_29,N_19956,N_19703);
or UO_30 (O_30,N_19672,N_19602);
nor UO_31 (O_31,N_19946,N_19708);
or UO_32 (O_32,N_19616,N_19642);
xnor UO_33 (O_33,N_19766,N_19816);
xor UO_34 (O_34,N_19661,N_19976);
and UO_35 (O_35,N_19803,N_19610);
nor UO_36 (O_36,N_19772,N_19782);
xor UO_37 (O_37,N_19947,N_19955);
nor UO_38 (O_38,N_19631,N_19608);
and UO_39 (O_39,N_19847,N_19624);
or UO_40 (O_40,N_19980,N_19822);
xnor UO_41 (O_41,N_19694,N_19735);
xor UO_42 (O_42,N_19938,N_19991);
xor UO_43 (O_43,N_19906,N_19770);
nand UO_44 (O_44,N_19984,N_19680);
nand UO_45 (O_45,N_19741,N_19988);
and UO_46 (O_46,N_19742,N_19818);
xnor UO_47 (O_47,N_19718,N_19783);
nand UO_48 (O_48,N_19733,N_19633);
nand UO_49 (O_49,N_19959,N_19644);
or UO_50 (O_50,N_19895,N_19660);
or UO_51 (O_51,N_19873,N_19755);
xnor UO_52 (O_52,N_19740,N_19950);
nor UO_53 (O_53,N_19894,N_19702);
nor UO_54 (O_54,N_19797,N_19665);
nand UO_55 (O_55,N_19728,N_19875);
nor UO_56 (O_56,N_19969,N_19826);
or UO_57 (O_57,N_19958,N_19903);
xor UO_58 (O_58,N_19776,N_19834);
or UO_59 (O_59,N_19931,N_19656);
xor UO_60 (O_60,N_19620,N_19611);
or UO_61 (O_61,N_19989,N_19995);
nand UO_62 (O_62,N_19765,N_19990);
nor UO_63 (O_63,N_19884,N_19681);
or UO_64 (O_64,N_19692,N_19983);
xor UO_65 (O_65,N_19730,N_19747);
xnor UO_66 (O_66,N_19823,N_19697);
nor UO_67 (O_67,N_19916,N_19864);
and UO_68 (O_68,N_19859,N_19601);
and UO_69 (O_69,N_19954,N_19813);
xor UO_70 (O_70,N_19979,N_19638);
nor UO_71 (O_71,N_19945,N_19833);
nand UO_72 (O_72,N_19707,N_19897);
xor UO_73 (O_73,N_19805,N_19650);
or UO_74 (O_74,N_19912,N_19727);
and UO_75 (O_75,N_19861,N_19904);
and UO_76 (O_76,N_19796,N_19798);
nand UO_77 (O_77,N_19971,N_19930);
or UO_78 (O_78,N_19932,N_19846);
xor UO_79 (O_79,N_19820,N_19723);
xor UO_80 (O_80,N_19769,N_19664);
xor UO_81 (O_81,N_19716,N_19911);
and UO_82 (O_82,N_19639,N_19793);
xnor UO_83 (O_83,N_19637,N_19720);
nor UO_84 (O_84,N_19835,N_19636);
and UO_85 (O_85,N_19937,N_19821);
and UO_86 (O_86,N_19871,N_19754);
and UO_87 (O_87,N_19900,N_19651);
and UO_88 (O_88,N_19817,N_19853);
xnor UO_89 (O_89,N_19600,N_19612);
and UO_90 (O_90,N_19693,N_19632);
nor UO_91 (O_91,N_19771,N_19676);
nand UO_92 (O_92,N_19691,N_19974);
nand UO_93 (O_93,N_19605,N_19868);
or UO_94 (O_94,N_19815,N_19924);
or UO_95 (O_95,N_19909,N_19628);
nor UO_96 (O_96,N_19749,N_19824);
and UO_97 (O_97,N_19779,N_19748);
nor UO_98 (O_98,N_19750,N_19603);
and UO_99 (O_99,N_19677,N_19719);
xor UO_100 (O_100,N_19923,N_19926);
or UO_101 (O_101,N_19934,N_19841);
nor UO_102 (O_102,N_19806,N_19999);
and UO_103 (O_103,N_19918,N_19996);
xor UO_104 (O_104,N_19655,N_19867);
and UO_105 (O_105,N_19674,N_19761);
xor UO_106 (O_106,N_19737,N_19808);
or UO_107 (O_107,N_19629,N_19762);
or UO_108 (O_108,N_19621,N_19961);
nand UO_109 (O_109,N_19940,N_19706);
nor UO_110 (O_110,N_19799,N_19763);
or UO_111 (O_111,N_19878,N_19830);
and UO_112 (O_112,N_19836,N_19819);
nor UO_113 (O_113,N_19837,N_19757);
nand UO_114 (O_114,N_19978,N_19854);
xnor UO_115 (O_115,N_19832,N_19807);
or UO_116 (O_116,N_19948,N_19809);
and UO_117 (O_117,N_19986,N_19872);
xor UO_118 (O_118,N_19684,N_19893);
or UO_119 (O_119,N_19925,N_19919);
and UO_120 (O_120,N_19953,N_19615);
and UO_121 (O_121,N_19690,N_19787);
xor UO_122 (O_122,N_19877,N_19645);
nor UO_123 (O_123,N_19627,N_19673);
and UO_124 (O_124,N_19767,N_19778);
xor UO_125 (O_125,N_19812,N_19667);
nor UO_126 (O_126,N_19910,N_19701);
or UO_127 (O_127,N_19654,N_19800);
or UO_128 (O_128,N_19860,N_19679);
nand UO_129 (O_129,N_19851,N_19666);
nand UO_130 (O_130,N_19780,N_19678);
and UO_131 (O_131,N_19715,N_19905);
xor UO_132 (O_132,N_19791,N_19972);
xor UO_133 (O_133,N_19790,N_19975);
nand UO_134 (O_134,N_19685,N_19942);
nand UO_135 (O_135,N_19887,N_19775);
and UO_136 (O_136,N_19722,N_19709);
xnor UO_137 (O_137,N_19985,N_19970);
nor UO_138 (O_138,N_19994,N_19683);
nor UO_139 (O_139,N_19609,N_19652);
or UO_140 (O_140,N_19981,N_19936);
xor UO_141 (O_141,N_19865,N_19883);
or UO_142 (O_142,N_19622,N_19713);
nor UO_143 (O_143,N_19699,N_19939);
or UO_144 (O_144,N_19659,N_19941);
or UO_145 (O_145,N_19876,N_19751);
or UO_146 (O_146,N_19635,N_19647);
nand UO_147 (O_147,N_19901,N_19917);
and UO_148 (O_148,N_19786,N_19682);
nand UO_149 (O_149,N_19908,N_19619);
xnor UO_150 (O_150,N_19784,N_19670);
xnor UO_151 (O_151,N_19831,N_19888);
or UO_152 (O_152,N_19671,N_19885);
nand UO_153 (O_153,N_19907,N_19882);
nor UO_154 (O_154,N_19966,N_19617);
nand UO_155 (O_155,N_19746,N_19745);
xnor UO_156 (O_156,N_19811,N_19827);
or UO_157 (O_157,N_19613,N_19753);
nand UO_158 (O_158,N_19777,N_19828);
nand UO_159 (O_159,N_19892,N_19963);
xor UO_160 (O_160,N_19734,N_19920);
xnor UO_161 (O_161,N_19686,N_19998);
xor UO_162 (O_162,N_19849,N_19858);
nand UO_163 (O_163,N_19653,N_19739);
or UO_164 (O_164,N_19738,N_19850);
and UO_165 (O_165,N_19899,N_19774);
nor UO_166 (O_166,N_19922,N_19840);
or UO_167 (O_167,N_19726,N_19879);
xnor UO_168 (O_168,N_19768,N_19844);
xor UO_169 (O_169,N_19626,N_19886);
nor UO_170 (O_170,N_19915,N_19743);
and UO_171 (O_171,N_19982,N_19714);
nand UO_172 (O_172,N_19874,N_19752);
nor UO_173 (O_173,N_19960,N_19789);
nor UO_174 (O_174,N_19913,N_19675);
or UO_175 (O_175,N_19687,N_19881);
and UO_176 (O_176,N_19933,N_19658);
xor UO_177 (O_177,N_19943,N_19869);
nor UO_178 (O_178,N_19967,N_19839);
nor UO_179 (O_179,N_19862,N_19880);
or UO_180 (O_180,N_19795,N_19606);
and UO_181 (O_181,N_19764,N_19987);
or UO_182 (O_182,N_19785,N_19810);
nor UO_183 (O_183,N_19843,N_19704);
xnor UO_184 (O_184,N_19760,N_19618);
and UO_185 (O_185,N_19964,N_19781);
and UO_186 (O_186,N_19725,N_19852);
or UO_187 (O_187,N_19825,N_19929);
or UO_188 (O_188,N_19914,N_19944);
or UO_189 (O_189,N_19688,N_19641);
nand UO_190 (O_190,N_19648,N_19700);
and UO_191 (O_191,N_19731,N_19788);
nand UO_192 (O_192,N_19696,N_19848);
nor UO_193 (O_193,N_19630,N_19744);
nand UO_194 (O_194,N_19902,N_19604);
nor UO_195 (O_195,N_19710,N_19857);
xnor UO_196 (O_196,N_19724,N_19646);
xor UO_197 (O_197,N_19759,N_19689);
xor UO_198 (O_198,N_19712,N_19717);
nand UO_199 (O_199,N_19640,N_19814);
xnor UO_200 (O_200,N_19687,N_19662);
and UO_201 (O_201,N_19975,N_19718);
or UO_202 (O_202,N_19972,N_19787);
xnor UO_203 (O_203,N_19919,N_19716);
nand UO_204 (O_204,N_19917,N_19859);
xnor UO_205 (O_205,N_19989,N_19771);
nor UO_206 (O_206,N_19663,N_19826);
nand UO_207 (O_207,N_19703,N_19943);
nor UO_208 (O_208,N_19805,N_19796);
nor UO_209 (O_209,N_19819,N_19913);
nor UO_210 (O_210,N_19910,N_19851);
nand UO_211 (O_211,N_19655,N_19888);
or UO_212 (O_212,N_19792,N_19776);
nor UO_213 (O_213,N_19779,N_19799);
nand UO_214 (O_214,N_19638,N_19879);
xor UO_215 (O_215,N_19937,N_19997);
xnor UO_216 (O_216,N_19872,N_19968);
and UO_217 (O_217,N_19614,N_19627);
and UO_218 (O_218,N_19796,N_19969);
xnor UO_219 (O_219,N_19906,N_19746);
or UO_220 (O_220,N_19726,N_19841);
or UO_221 (O_221,N_19775,N_19717);
xnor UO_222 (O_222,N_19702,N_19613);
nand UO_223 (O_223,N_19930,N_19859);
nor UO_224 (O_224,N_19667,N_19927);
nor UO_225 (O_225,N_19839,N_19796);
nor UO_226 (O_226,N_19836,N_19954);
or UO_227 (O_227,N_19684,N_19870);
xor UO_228 (O_228,N_19617,N_19647);
nand UO_229 (O_229,N_19725,N_19884);
nor UO_230 (O_230,N_19957,N_19671);
and UO_231 (O_231,N_19833,N_19979);
xnor UO_232 (O_232,N_19992,N_19977);
nand UO_233 (O_233,N_19962,N_19801);
nor UO_234 (O_234,N_19901,N_19696);
xor UO_235 (O_235,N_19843,N_19901);
xor UO_236 (O_236,N_19952,N_19626);
and UO_237 (O_237,N_19922,N_19647);
nor UO_238 (O_238,N_19805,N_19797);
nand UO_239 (O_239,N_19927,N_19632);
nand UO_240 (O_240,N_19637,N_19712);
nor UO_241 (O_241,N_19735,N_19670);
or UO_242 (O_242,N_19933,N_19748);
nand UO_243 (O_243,N_19927,N_19745);
nor UO_244 (O_244,N_19714,N_19725);
nand UO_245 (O_245,N_19863,N_19788);
or UO_246 (O_246,N_19707,N_19984);
xor UO_247 (O_247,N_19608,N_19746);
nor UO_248 (O_248,N_19750,N_19810);
or UO_249 (O_249,N_19805,N_19800);
or UO_250 (O_250,N_19854,N_19891);
nor UO_251 (O_251,N_19760,N_19792);
nand UO_252 (O_252,N_19813,N_19774);
nor UO_253 (O_253,N_19608,N_19909);
nand UO_254 (O_254,N_19757,N_19889);
or UO_255 (O_255,N_19699,N_19824);
or UO_256 (O_256,N_19662,N_19618);
and UO_257 (O_257,N_19755,N_19804);
and UO_258 (O_258,N_19905,N_19831);
nor UO_259 (O_259,N_19779,N_19981);
nor UO_260 (O_260,N_19933,N_19795);
xor UO_261 (O_261,N_19808,N_19626);
xor UO_262 (O_262,N_19959,N_19683);
nor UO_263 (O_263,N_19617,N_19771);
or UO_264 (O_264,N_19765,N_19780);
xor UO_265 (O_265,N_19705,N_19734);
nand UO_266 (O_266,N_19672,N_19915);
nand UO_267 (O_267,N_19781,N_19601);
xor UO_268 (O_268,N_19743,N_19922);
nand UO_269 (O_269,N_19763,N_19942);
and UO_270 (O_270,N_19666,N_19872);
nor UO_271 (O_271,N_19705,N_19933);
xnor UO_272 (O_272,N_19638,N_19929);
nor UO_273 (O_273,N_19958,N_19647);
xnor UO_274 (O_274,N_19950,N_19631);
nor UO_275 (O_275,N_19734,N_19818);
nand UO_276 (O_276,N_19804,N_19900);
or UO_277 (O_277,N_19725,N_19795);
nand UO_278 (O_278,N_19721,N_19753);
and UO_279 (O_279,N_19974,N_19673);
xnor UO_280 (O_280,N_19738,N_19704);
nand UO_281 (O_281,N_19603,N_19951);
or UO_282 (O_282,N_19957,N_19863);
or UO_283 (O_283,N_19812,N_19840);
and UO_284 (O_284,N_19880,N_19947);
and UO_285 (O_285,N_19612,N_19900);
xnor UO_286 (O_286,N_19740,N_19812);
xnor UO_287 (O_287,N_19612,N_19717);
and UO_288 (O_288,N_19791,N_19883);
xnor UO_289 (O_289,N_19696,N_19843);
xnor UO_290 (O_290,N_19918,N_19620);
nand UO_291 (O_291,N_19942,N_19705);
and UO_292 (O_292,N_19813,N_19790);
or UO_293 (O_293,N_19846,N_19696);
xnor UO_294 (O_294,N_19850,N_19960);
and UO_295 (O_295,N_19683,N_19740);
and UO_296 (O_296,N_19814,N_19638);
nand UO_297 (O_297,N_19898,N_19721);
nand UO_298 (O_298,N_19866,N_19655);
nand UO_299 (O_299,N_19693,N_19704);
or UO_300 (O_300,N_19651,N_19672);
and UO_301 (O_301,N_19807,N_19686);
and UO_302 (O_302,N_19907,N_19784);
nand UO_303 (O_303,N_19837,N_19925);
or UO_304 (O_304,N_19897,N_19957);
nand UO_305 (O_305,N_19766,N_19946);
xnor UO_306 (O_306,N_19620,N_19663);
xor UO_307 (O_307,N_19791,N_19750);
and UO_308 (O_308,N_19748,N_19863);
and UO_309 (O_309,N_19804,N_19606);
nand UO_310 (O_310,N_19628,N_19637);
and UO_311 (O_311,N_19626,N_19844);
and UO_312 (O_312,N_19960,N_19910);
and UO_313 (O_313,N_19924,N_19778);
or UO_314 (O_314,N_19829,N_19629);
nor UO_315 (O_315,N_19796,N_19736);
or UO_316 (O_316,N_19877,N_19902);
nand UO_317 (O_317,N_19894,N_19736);
or UO_318 (O_318,N_19969,N_19611);
nor UO_319 (O_319,N_19951,N_19810);
xor UO_320 (O_320,N_19621,N_19763);
xnor UO_321 (O_321,N_19857,N_19921);
nor UO_322 (O_322,N_19938,N_19808);
nor UO_323 (O_323,N_19706,N_19979);
nand UO_324 (O_324,N_19693,N_19714);
nor UO_325 (O_325,N_19945,N_19697);
or UO_326 (O_326,N_19639,N_19733);
nor UO_327 (O_327,N_19868,N_19973);
nand UO_328 (O_328,N_19916,N_19678);
nor UO_329 (O_329,N_19793,N_19614);
xnor UO_330 (O_330,N_19943,N_19755);
or UO_331 (O_331,N_19825,N_19839);
nor UO_332 (O_332,N_19922,N_19891);
and UO_333 (O_333,N_19722,N_19784);
or UO_334 (O_334,N_19997,N_19963);
xor UO_335 (O_335,N_19969,N_19651);
and UO_336 (O_336,N_19970,N_19753);
xnor UO_337 (O_337,N_19661,N_19759);
nand UO_338 (O_338,N_19644,N_19736);
nand UO_339 (O_339,N_19643,N_19670);
xor UO_340 (O_340,N_19610,N_19661);
nand UO_341 (O_341,N_19735,N_19719);
or UO_342 (O_342,N_19730,N_19837);
xor UO_343 (O_343,N_19808,N_19796);
nor UO_344 (O_344,N_19632,N_19675);
and UO_345 (O_345,N_19741,N_19777);
and UO_346 (O_346,N_19860,N_19782);
or UO_347 (O_347,N_19673,N_19943);
xnor UO_348 (O_348,N_19845,N_19915);
or UO_349 (O_349,N_19627,N_19636);
nand UO_350 (O_350,N_19606,N_19999);
and UO_351 (O_351,N_19805,N_19831);
and UO_352 (O_352,N_19697,N_19668);
nand UO_353 (O_353,N_19986,N_19845);
or UO_354 (O_354,N_19990,N_19658);
nor UO_355 (O_355,N_19618,N_19792);
nor UO_356 (O_356,N_19866,N_19687);
nand UO_357 (O_357,N_19650,N_19905);
xnor UO_358 (O_358,N_19997,N_19662);
nand UO_359 (O_359,N_19718,N_19981);
and UO_360 (O_360,N_19691,N_19728);
nand UO_361 (O_361,N_19986,N_19942);
xnor UO_362 (O_362,N_19870,N_19825);
or UO_363 (O_363,N_19606,N_19650);
xnor UO_364 (O_364,N_19808,N_19636);
nor UO_365 (O_365,N_19937,N_19674);
xor UO_366 (O_366,N_19717,N_19974);
xnor UO_367 (O_367,N_19851,N_19703);
nor UO_368 (O_368,N_19842,N_19679);
or UO_369 (O_369,N_19760,N_19901);
nor UO_370 (O_370,N_19782,N_19804);
nand UO_371 (O_371,N_19811,N_19937);
or UO_372 (O_372,N_19758,N_19855);
xor UO_373 (O_373,N_19850,N_19955);
nor UO_374 (O_374,N_19803,N_19983);
nand UO_375 (O_375,N_19740,N_19761);
nand UO_376 (O_376,N_19911,N_19893);
and UO_377 (O_377,N_19918,N_19981);
or UO_378 (O_378,N_19980,N_19949);
nor UO_379 (O_379,N_19831,N_19750);
and UO_380 (O_380,N_19956,N_19783);
nor UO_381 (O_381,N_19904,N_19797);
nor UO_382 (O_382,N_19783,N_19666);
nand UO_383 (O_383,N_19739,N_19967);
or UO_384 (O_384,N_19725,N_19846);
and UO_385 (O_385,N_19693,N_19853);
or UO_386 (O_386,N_19839,N_19621);
and UO_387 (O_387,N_19766,N_19685);
nand UO_388 (O_388,N_19843,N_19963);
xnor UO_389 (O_389,N_19834,N_19736);
nand UO_390 (O_390,N_19922,N_19889);
xor UO_391 (O_391,N_19675,N_19829);
nor UO_392 (O_392,N_19653,N_19658);
nor UO_393 (O_393,N_19639,N_19743);
or UO_394 (O_394,N_19611,N_19980);
xnor UO_395 (O_395,N_19645,N_19701);
nor UO_396 (O_396,N_19786,N_19915);
xnor UO_397 (O_397,N_19722,N_19990);
xnor UO_398 (O_398,N_19879,N_19632);
nor UO_399 (O_399,N_19700,N_19938);
or UO_400 (O_400,N_19819,N_19944);
and UO_401 (O_401,N_19603,N_19691);
nand UO_402 (O_402,N_19960,N_19662);
xnor UO_403 (O_403,N_19900,N_19828);
nand UO_404 (O_404,N_19854,N_19604);
xnor UO_405 (O_405,N_19749,N_19661);
and UO_406 (O_406,N_19604,N_19823);
xor UO_407 (O_407,N_19951,N_19780);
xor UO_408 (O_408,N_19779,N_19934);
xnor UO_409 (O_409,N_19694,N_19773);
or UO_410 (O_410,N_19609,N_19663);
nor UO_411 (O_411,N_19613,N_19697);
xnor UO_412 (O_412,N_19724,N_19819);
xor UO_413 (O_413,N_19614,N_19763);
nand UO_414 (O_414,N_19878,N_19730);
or UO_415 (O_415,N_19736,N_19799);
xnor UO_416 (O_416,N_19647,N_19747);
nand UO_417 (O_417,N_19953,N_19921);
nand UO_418 (O_418,N_19946,N_19868);
nor UO_419 (O_419,N_19952,N_19652);
nor UO_420 (O_420,N_19897,N_19799);
and UO_421 (O_421,N_19677,N_19781);
or UO_422 (O_422,N_19629,N_19684);
nand UO_423 (O_423,N_19672,N_19834);
nor UO_424 (O_424,N_19643,N_19608);
nor UO_425 (O_425,N_19895,N_19646);
xor UO_426 (O_426,N_19785,N_19725);
nand UO_427 (O_427,N_19683,N_19794);
or UO_428 (O_428,N_19635,N_19653);
nor UO_429 (O_429,N_19705,N_19721);
and UO_430 (O_430,N_19801,N_19889);
and UO_431 (O_431,N_19873,N_19845);
nor UO_432 (O_432,N_19828,N_19730);
nand UO_433 (O_433,N_19925,N_19932);
and UO_434 (O_434,N_19868,N_19979);
or UO_435 (O_435,N_19719,N_19800);
or UO_436 (O_436,N_19793,N_19846);
nand UO_437 (O_437,N_19881,N_19608);
or UO_438 (O_438,N_19650,N_19980);
nor UO_439 (O_439,N_19643,N_19610);
xor UO_440 (O_440,N_19608,N_19841);
xor UO_441 (O_441,N_19697,N_19851);
or UO_442 (O_442,N_19846,N_19710);
and UO_443 (O_443,N_19850,N_19987);
nand UO_444 (O_444,N_19728,N_19924);
nor UO_445 (O_445,N_19793,N_19987);
nand UO_446 (O_446,N_19851,N_19890);
xor UO_447 (O_447,N_19661,N_19758);
nand UO_448 (O_448,N_19720,N_19802);
nand UO_449 (O_449,N_19681,N_19733);
nor UO_450 (O_450,N_19977,N_19987);
xor UO_451 (O_451,N_19757,N_19641);
nand UO_452 (O_452,N_19691,N_19997);
nand UO_453 (O_453,N_19623,N_19869);
and UO_454 (O_454,N_19931,N_19689);
nor UO_455 (O_455,N_19754,N_19669);
xnor UO_456 (O_456,N_19996,N_19630);
and UO_457 (O_457,N_19980,N_19812);
or UO_458 (O_458,N_19983,N_19678);
nor UO_459 (O_459,N_19737,N_19886);
nand UO_460 (O_460,N_19826,N_19643);
and UO_461 (O_461,N_19882,N_19872);
nand UO_462 (O_462,N_19785,N_19710);
nor UO_463 (O_463,N_19809,N_19926);
nand UO_464 (O_464,N_19940,N_19908);
nand UO_465 (O_465,N_19750,N_19844);
or UO_466 (O_466,N_19867,N_19920);
and UO_467 (O_467,N_19824,N_19646);
xnor UO_468 (O_468,N_19658,N_19778);
xnor UO_469 (O_469,N_19678,N_19959);
xnor UO_470 (O_470,N_19752,N_19643);
xor UO_471 (O_471,N_19698,N_19791);
or UO_472 (O_472,N_19979,N_19916);
and UO_473 (O_473,N_19683,N_19923);
nand UO_474 (O_474,N_19703,N_19844);
and UO_475 (O_475,N_19949,N_19896);
xnor UO_476 (O_476,N_19976,N_19642);
nand UO_477 (O_477,N_19859,N_19947);
nor UO_478 (O_478,N_19611,N_19801);
nand UO_479 (O_479,N_19697,N_19891);
and UO_480 (O_480,N_19935,N_19605);
nor UO_481 (O_481,N_19673,N_19863);
xor UO_482 (O_482,N_19988,N_19804);
nor UO_483 (O_483,N_19795,N_19923);
nor UO_484 (O_484,N_19924,N_19990);
nand UO_485 (O_485,N_19692,N_19694);
xnor UO_486 (O_486,N_19832,N_19709);
or UO_487 (O_487,N_19685,N_19988);
xnor UO_488 (O_488,N_19989,N_19752);
and UO_489 (O_489,N_19907,N_19975);
or UO_490 (O_490,N_19891,N_19943);
nand UO_491 (O_491,N_19605,N_19815);
or UO_492 (O_492,N_19721,N_19847);
and UO_493 (O_493,N_19863,N_19937);
nand UO_494 (O_494,N_19781,N_19610);
and UO_495 (O_495,N_19949,N_19976);
xnor UO_496 (O_496,N_19600,N_19922);
nand UO_497 (O_497,N_19645,N_19930);
or UO_498 (O_498,N_19618,N_19653);
xor UO_499 (O_499,N_19984,N_19946);
and UO_500 (O_500,N_19659,N_19632);
nor UO_501 (O_501,N_19792,N_19674);
nand UO_502 (O_502,N_19749,N_19696);
or UO_503 (O_503,N_19866,N_19705);
or UO_504 (O_504,N_19764,N_19753);
xor UO_505 (O_505,N_19918,N_19682);
xor UO_506 (O_506,N_19769,N_19823);
nor UO_507 (O_507,N_19965,N_19939);
or UO_508 (O_508,N_19833,N_19795);
and UO_509 (O_509,N_19731,N_19609);
or UO_510 (O_510,N_19969,N_19778);
nand UO_511 (O_511,N_19651,N_19974);
and UO_512 (O_512,N_19663,N_19725);
nand UO_513 (O_513,N_19744,N_19940);
or UO_514 (O_514,N_19936,N_19719);
xnor UO_515 (O_515,N_19698,N_19815);
or UO_516 (O_516,N_19771,N_19804);
nor UO_517 (O_517,N_19824,N_19683);
or UO_518 (O_518,N_19870,N_19977);
and UO_519 (O_519,N_19748,N_19685);
or UO_520 (O_520,N_19952,N_19971);
or UO_521 (O_521,N_19633,N_19827);
nand UO_522 (O_522,N_19746,N_19984);
nand UO_523 (O_523,N_19845,N_19601);
and UO_524 (O_524,N_19744,N_19656);
or UO_525 (O_525,N_19867,N_19709);
or UO_526 (O_526,N_19826,N_19717);
nor UO_527 (O_527,N_19878,N_19660);
nor UO_528 (O_528,N_19762,N_19865);
or UO_529 (O_529,N_19928,N_19776);
nor UO_530 (O_530,N_19656,N_19638);
nand UO_531 (O_531,N_19947,N_19633);
nand UO_532 (O_532,N_19763,N_19832);
nor UO_533 (O_533,N_19939,N_19737);
xnor UO_534 (O_534,N_19761,N_19616);
nand UO_535 (O_535,N_19619,N_19886);
and UO_536 (O_536,N_19987,N_19729);
nand UO_537 (O_537,N_19605,N_19806);
and UO_538 (O_538,N_19944,N_19907);
nand UO_539 (O_539,N_19610,N_19985);
or UO_540 (O_540,N_19764,N_19959);
nand UO_541 (O_541,N_19850,N_19647);
nor UO_542 (O_542,N_19782,N_19684);
nand UO_543 (O_543,N_19870,N_19809);
and UO_544 (O_544,N_19751,N_19918);
or UO_545 (O_545,N_19600,N_19831);
nor UO_546 (O_546,N_19688,N_19729);
nand UO_547 (O_547,N_19975,N_19794);
and UO_548 (O_548,N_19944,N_19748);
nor UO_549 (O_549,N_19801,N_19957);
xor UO_550 (O_550,N_19620,N_19669);
xor UO_551 (O_551,N_19912,N_19802);
xnor UO_552 (O_552,N_19626,N_19981);
or UO_553 (O_553,N_19655,N_19765);
or UO_554 (O_554,N_19610,N_19680);
or UO_555 (O_555,N_19759,N_19669);
xnor UO_556 (O_556,N_19857,N_19640);
xnor UO_557 (O_557,N_19866,N_19886);
xor UO_558 (O_558,N_19946,N_19925);
nand UO_559 (O_559,N_19634,N_19972);
or UO_560 (O_560,N_19618,N_19774);
nand UO_561 (O_561,N_19809,N_19700);
nor UO_562 (O_562,N_19616,N_19954);
or UO_563 (O_563,N_19852,N_19613);
or UO_564 (O_564,N_19653,N_19813);
xnor UO_565 (O_565,N_19991,N_19704);
xor UO_566 (O_566,N_19754,N_19987);
nand UO_567 (O_567,N_19928,N_19896);
and UO_568 (O_568,N_19839,N_19716);
nor UO_569 (O_569,N_19903,N_19997);
nor UO_570 (O_570,N_19758,N_19603);
and UO_571 (O_571,N_19765,N_19841);
xnor UO_572 (O_572,N_19888,N_19950);
and UO_573 (O_573,N_19813,N_19807);
nor UO_574 (O_574,N_19692,N_19800);
xnor UO_575 (O_575,N_19674,N_19809);
xor UO_576 (O_576,N_19987,N_19769);
or UO_577 (O_577,N_19796,N_19774);
nand UO_578 (O_578,N_19704,N_19686);
nor UO_579 (O_579,N_19920,N_19931);
nand UO_580 (O_580,N_19706,N_19696);
nor UO_581 (O_581,N_19969,N_19923);
nor UO_582 (O_582,N_19947,N_19973);
or UO_583 (O_583,N_19894,N_19815);
or UO_584 (O_584,N_19675,N_19792);
nor UO_585 (O_585,N_19667,N_19886);
and UO_586 (O_586,N_19707,N_19776);
or UO_587 (O_587,N_19616,N_19763);
nand UO_588 (O_588,N_19951,N_19884);
or UO_589 (O_589,N_19931,N_19769);
nor UO_590 (O_590,N_19986,N_19920);
nand UO_591 (O_591,N_19751,N_19851);
xor UO_592 (O_592,N_19930,N_19861);
nor UO_593 (O_593,N_19992,N_19852);
nor UO_594 (O_594,N_19690,N_19850);
xor UO_595 (O_595,N_19700,N_19939);
or UO_596 (O_596,N_19944,N_19611);
nand UO_597 (O_597,N_19657,N_19701);
and UO_598 (O_598,N_19738,N_19625);
nand UO_599 (O_599,N_19812,N_19852);
or UO_600 (O_600,N_19734,N_19805);
or UO_601 (O_601,N_19742,N_19898);
and UO_602 (O_602,N_19752,N_19814);
or UO_603 (O_603,N_19798,N_19621);
and UO_604 (O_604,N_19956,N_19916);
xnor UO_605 (O_605,N_19993,N_19930);
nor UO_606 (O_606,N_19669,N_19931);
and UO_607 (O_607,N_19850,N_19641);
nand UO_608 (O_608,N_19900,N_19768);
and UO_609 (O_609,N_19934,N_19603);
and UO_610 (O_610,N_19690,N_19614);
or UO_611 (O_611,N_19810,N_19729);
nor UO_612 (O_612,N_19787,N_19790);
nor UO_613 (O_613,N_19956,N_19899);
xnor UO_614 (O_614,N_19704,N_19730);
xor UO_615 (O_615,N_19780,N_19617);
xnor UO_616 (O_616,N_19675,N_19771);
xor UO_617 (O_617,N_19884,N_19825);
or UO_618 (O_618,N_19813,N_19862);
xor UO_619 (O_619,N_19986,N_19814);
nor UO_620 (O_620,N_19720,N_19926);
and UO_621 (O_621,N_19624,N_19716);
or UO_622 (O_622,N_19721,N_19955);
nor UO_623 (O_623,N_19826,N_19789);
or UO_624 (O_624,N_19754,N_19736);
nor UO_625 (O_625,N_19773,N_19857);
nand UO_626 (O_626,N_19780,N_19860);
and UO_627 (O_627,N_19829,N_19812);
and UO_628 (O_628,N_19803,N_19910);
nor UO_629 (O_629,N_19603,N_19717);
and UO_630 (O_630,N_19806,N_19884);
or UO_631 (O_631,N_19775,N_19900);
nand UO_632 (O_632,N_19917,N_19774);
and UO_633 (O_633,N_19623,N_19816);
and UO_634 (O_634,N_19610,N_19866);
or UO_635 (O_635,N_19769,N_19833);
nand UO_636 (O_636,N_19662,N_19971);
nand UO_637 (O_637,N_19900,N_19922);
xnor UO_638 (O_638,N_19884,N_19812);
nand UO_639 (O_639,N_19879,N_19647);
or UO_640 (O_640,N_19867,N_19955);
and UO_641 (O_641,N_19743,N_19676);
and UO_642 (O_642,N_19698,N_19654);
nand UO_643 (O_643,N_19787,N_19873);
nor UO_644 (O_644,N_19798,N_19844);
or UO_645 (O_645,N_19829,N_19759);
and UO_646 (O_646,N_19814,N_19629);
or UO_647 (O_647,N_19762,N_19754);
nand UO_648 (O_648,N_19747,N_19684);
or UO_649 (O_649,N_19708,N_19645);
xnor UO_650 (O_650,N_19798,N_19738);
xor UO_651 (O_651,N_19962,N_19964);
nor UO_652 (O_652,N_19991,N_19826);
nor UO_653 (O_653,N_19855,N_19643);
and UO_654 (O_654,N_19710,N_19782);
and UO_655 (O_655,N_19633,N_19641);
xor UO_656 (O_656,N_19926,N_19635);
nand UO_657 (O_657,N_19693,N_19794);
and UO_658 (O_658,N_19979,N_19710);
and UO_659 (O_659,N_19869,N_19769);
and UO_660 (O_660,N_19688,N_19911);
xnor UO_661 (O_661,N_19737,N_19976);
or UO_662 (O_662,N_19665,N_19653);
xnor UO_663 (O_663,N_19891,N_19702);
xor UO_664 (O_664,N_19652,N_19662);
or UO_665 (O_665,N_19692,N_19998);
nand UO_666 (O_666,N_19889,N_19869);
nor UO_667 (O_667,N_19899,N_19941);
xnor UO_668 (O_668,N_19828,N_19685);
xnor UO_669 (O_669,N_19626,N_19689);
or UO_670 (O_670,N_19873,N_19770);
xor UO_671 (O_671,N_19987,N_19637);
and UO_672 (O_672,N_19696,N_19932);
xnor UO_673 (O_673,N_19851,N_19780);
xor UO_674 (O_674,N_19885,N_19812);
or UO_675 (O_675,N_19612,N_19839);
or UO_676 (O_676,N_19744,N_19616);
nand UO_677 (O_677,N_19739,N_19877);
nor UO_678 (O_678,N_19745,N_19733);
or UO_679 (O_679,N_19674,N_19636);
or UO_680 (O_680,N_19722,N_19968);
nor UO_681 (O_681,N_19722,N_19662);
nor UO_682 (O_682,N_19928,N_19840);
nand UO_683 (O_683,N_19844,N_19939);
nor UO_684 (O_684,N_19652,N_19963);
nor UO_685 (O_685,N_19657,N_19699);
and UO_686 (O_686,N_19737,N_19626);
or UO_687 (O_687,N_19635,N_19722);
and UO_688 (O_688,N_19601,N_19875);
xnor UO_689 (O_689,N_19911,N_19779);
nand UO_690 (O_690,N_19986,N_19723);
xor UO_691 (O_691,N_19927,N_19681);
xor UO_692 (O_692,N_19961,N_19987);
and UO_693 (O_693,N_19814,N_19891);
xnor UO_694 (O_694,N_19798,N_19755);
or UO_695 (O_695,N_19906,N_19684);
nand UO_696 (O_696,N_19905,N_19787);
nand UO_697 (O_697,N_19926,N_19704);
xnor UO_698 (O_698,N_19696,N_19720);
or UO_699 (O_699,N_19675,N_19827);
nand UO_700 (O_700,N_19830,N_19626);
and UO_701 (O_701,N_19650,N_19972);
xor UO_702 (O_702,N_19797,N_19763);
nand UO_703 (O_703,N_19651,N_19770);
or UO_704 (O_704,N_19834,N_19862);
or UO_705 (O_705,N_19927,N_19707);
nand UO_706 (O_706,N_19787,N_19799);
nand UO_707 (O_707,N_19857,N_19917);
and UO_708 (O_708,N_19916,N_19959);
nand UO_709 (O_709,N_19700,N_19663);
nor UO_710 (O_710,N_19695,N_19672);
xor UO_711 (O_711,N_19882,N_19694);
xor UO_712 (O_712,N_19769,N_19858);
nor UO_713 (O_713,N_19736,N_19712);
xnor UO_714 (O_714,N_19675,N_19751);
nand UO_715 (O_715,N_19750,N_19687);
nand UO_716 (O_716,N_19626,N_19602);
xnor UO_717 (O_717,N_19744,N_19705);
or UO_718 (O_718,N_19928,N_19893);
xnor UO_719 (O_719,N_19972,N_19883);
xor UO_720 (O_720,N_19974,N_19626);
and UO_721 (O_721,N_19900,N_19762);
nor UO_722 (O_722,N_19862,N_19629);
nand UO_723 (O_723,N_19740,N_19691);
nor UO_724 (O_724,N_19939,N_19635);
or UO_725 (O_725,N_19962,N_19709);
nor UO_726 (O_726,N_19840,N_19893);
xnor UO_727 (O_727,N_19815,N_19921);
nand UO_728 (O_728,N_19828,N_19747);
nand UO_729 (O_729,N_19760,N_19790);
or UO_730 (O_730,N_19651,N_19800);
nor UO_731 (O_731,N_19786,N_19858);
xnor UO_732 (O_732,N_19910,N_19829);
and UO_733 (O_733,N_19617,N_19831);
and UO_734 (O_734,N_19807,N_19860);
xnor UO_735 (O_735,N_19660,N_19901);
and UO_736 (O_736,N_19637,N_19870);
nor UO_737 (O_737,N_19655,N_19801);
and UO_738 (O_738,N_19790,N_19618);
and UO_739 (O_739,N_19861,N_19806);
and UO_740 (O_740,N_19906,N_19651);
xnor UO_741 (O_741,N_19924,N_19903);
nor UO_742 (O_742,N_19919,N_19751);
or UO_743 (O_743,N_19605,N_19905);
xnor UO_744 (O_744,N_19895,N_19899);
xor UO_745 (O_745,N_19786,N_19978);
nand UO_746 (O_746,N_19635,N_19620);
or UO_747 (O_747,N_19677,N_19790);
nor UO_748 (O_748,N_19946,N_19664);
xnor UO_749 (O_749,N_19753,N_19922);
nor UO_750 (O_750,N_19787,N_19865);
nand UO_751 (O_751,N_19965,N_19607);
and UO_752 (O_752,N_19853,N_19991);
xnor UO_753 (O_753,N_19683,N_19768);
nor UO_754 (O_754,N_19707,N_19623);
nor UO_755 (O_755,N_19902,N_19735);
or UO_756 (O_756,N_19822,N_19897);
and UO_757 (O_757,N_19831,N_19649);
xnor UO_758 (O_758,N_19800,N_19867);
xnor UO_759 (O_759,N_19744,N_19975);
and UO_760 (O_760,N_19886,N_19947);
and UO_761 (O_761,N_19963,N_19666);
and UO_762 (O_762,N_19921,N_19880);
and UO_763 (O_763,N_19839,N_19922);
nand UO_764 (O_764,N_19949,N_19629);
nor UO_765 (O_765,N_19737,N_19958);
nor UO_766 (O_766,N_19778,N_19922);
xor UO_767 (O_767,N_19888,N_19842);
xnor UO_768 (O_768,N_19906,N_19814);
nor UO_769 (O_769,N_19645,N_19840);
nand UO_770 (O_770,N_19851,N_19738);
and UO_771 (O_771,N_19949,N_19639);
nor UO_772 (O_772,N_19610,N_19819);
xnor UO_773 (O_773,N_19632,N_19803);
nor UO_774 (O_774,N_19982,N_19884);
xor UO_775 (O_775,N_19790,N_19682);
or UO_776 (O_776,N_19892,N_19902);
nand UO_777 (O_777,N_19803,N_19853);
xor UO_778 (O_778,N_19972,N_19961);
and UO_779 (O_779,N_19785,N_19697);
and UO_780 (O_780,N_19756,N_19732);
nor UO_781 (O_781,N_19615,N_19819);
and UO_782 (O_782,N_19930,N_19932);
xor UO_783 (O_783,N_19825,N_19819);
xor UO_784 (O_784,N_19672,N_19752);
nor UO_785 (O_785,N_19726,N_19675);
nand UO_786 (O_786,N_19785,N_19958);
nor UO_787 (O_787,N_19857,N_19652);
nand UO_788 (O_788,N_19927,N_19916);
xnor UO_789 (O_789,N_19631,N_19639);
nand UO_790 (O_790,N_19641,N_19630);
xor UO_791 (O_791,N_19797,N_19949);
or UO_792 (O_792,N_19649,N_19852);
or UO_793 (O_793,N_19688,N_19935);
nor UO_794 (O_794,N_19747,N_19822);
or UO_795 (O_795,N_19807,N_19920);
nor UO_796 (O_796,N_19749,N_19673);
and UO_797 (O_797,N_19707,N_19712);
nor UO_798 (O_798,N_19906,N_19745);
nor UO_799 (O_799,N_19661,N_19942);
nand UO_800 (O_800,N_19754,N_19986);
nor UO_801 (O_801,N_19789,N_19707);
or UO_802 (O_802,N_19910,N_19807);
nor UO_803 (O_803,N_19852,N_19645);
nor UO_804 (O_804,N_19931,N_19604);
or UO_805 (O_805,N_19862,N_19918);
or UO_806 (O_806,N_19633,N_19798);
or UO_807 (O_807,N_19889,N_19719);
nand UO_808 (O_808,N_19929,N_19630);
nand UO_809 (O_809,N_19739,N_19809);
and UO_810 (O_810,N_19786,N_19658);
nand UO_811 (O_811,N_19955,N_19601);
and UO_812 (O_812,N_19816,N_19957);
nand UO_813 (O_813,N_19916,N_19934);
xor UO_814 (O_814,N_19890,N_19995);
nor UO_815 (O_815,N_19608,N_19777);
and UO_816 (O_816,N_19958,N_19940);
nand UO_817 (O_817,N_19773,N_19844);
nor UO_818 (O_818,N_19750,N_19839);
and UO_819 (O_819,N_19736,N_19933);
nand UO_820 (O_820,N_19762,N_19931);
and UO_821 (O_821,N_19633,N_19796);
or UO_822 (O_822,N_19615,N_19625);
and UO_823 (O_823,N_19998,N_19741);
and UO_824 (O_824,N_19861,N_19984);
nand UO_825 (O_825,N_19614,N_19835);
or UO_826 (O_826,N_19626,N_19960);
or UO_827 (O_827,N_19858,N_19812);
xnor UO_828 (O_828,N_19759,N_19980);
or UO_829 (O_829,N_19661,N_19820);
and UO_830 (O_830,N_19980,N_19757);
xnor UO_831 (O_831,N_19650,N_19925);
xor UO_832 (O_832,N_19866,N_19980);
and UO_833 (O_833,N_19869,N_19964);
nand UO_834 (O_834,N_19999,N_19706);
and UO_835 (O_835,N_19860,N_19805);
xnor UO_836 (O_836,N_19829,N_19907);
or UO_837 (O_837,N_19722,N_19658);
or UO_838 (O_838,N_19778,N_19789);
nand UO_839 (O_839,N_19663,N_19828);
nand UO_840 (O_840,N_19626,N_19761);
or UO_841 (O_841,N_19841,N_19818);
or UO_842 (O_842,N_19731,N_19818);
xor UO_843 (O_843,N_19623,N_19946);
or UO_844 (O_844,N_19936,N_19679);
or UO_845 (O_845,N_19747,N_19768);
or UO_846 (O_846,N_19966,N_19651);
xor UO_847 (O_847,N_19677,N_19730);
xor UO_848 (O_848,N_19732,N_19817);
or UO_849 (O_849,N_19731,N_19803);
nand UO_850 (O_850,N_19859,N_19740);
or UO_851 (O_851,N_19730,N_19973);
and UO_852 (O_852,N_19881,N_19610);
nand UO_853 (O_853,N_19880,N_19750);
nor UO_854 (O_854,N_19863,N_19650);
or UO_855 (O_855,N_19846,N_19629);
nor UO_856 (O_856,N_19698,N_19656);
or UO_857 (O_857,N_19815,N_19944);
or UO_858 (O_858,N_19896,N_19789);
nand UO_859 (O_859,N_19768,N_19931);
nand UO_860 (O_860,N_19682,N_19989);
or UO_861 (O_861,N_19863,N_19678);
nand UO_862 (O_862,N_19988,N_19908);
nor UO_863 (O_863,N_19686,N_19629);
or UO_864 (O_864,N_19997,N_19700);
nand UO_865 (O_865,N_19880,N_19870);
and UO_866 (O_866,N_19751,N_19857);
and UO_867 (O_867,N_19619,N_19763);
nand UO_868 (O_868,N_19612,N_19639);
nand UO_869 (O_869,N_19930,N_19946);
nor UO_870 (O_870,N_19611,N_19762);
nor UO_871 (O_871,N_19821,N_19682);
and UO_872 (O_872,N_19653,N_19887);
or UO_873 (O_873,N_19900,N_19737);
nand UO_874 (O_874,N_19680,N_19943);
nor UO_875 (O_875,N_19722,N_19624);
or UO_876 (O_876,N_19752,N_19923);
or UO_877 (O_877,N_19873,N_19874);
and UO_878 (O_878,N_19601,N_19896);
nand UO_879 (O_879,N_19974,N_19851);
nand UO_880 (O_880,N_19843,N_19909);
or UO_881 (O_881,N_19802,N_19608);
nand UO_882 (O_882,N_19767,N_19834);
and UO_883 (O_883,N_19927,N_19726);
or UO_884 (O_884,N_19638,N_19807);
and UO_885 (O_885,N_19922,N_19843);
nand UO_886 (O_886,N_19650,N_19865);
or UO_887 (O_887,N_19900,N_19821);
and UO_888 (O_888,N_19974,N_19655);
nand UO_889 (O_889,N_19669,N_19823);
nor UO_890 (O_890,N_19784,N_19772);
nor UO_891 (O_891,N_19714,N_19874);
and UO_892 (O_892,N_19831,N_19809);
or UO_893 (O_893,N_19756,N_19882);
xnor UO_894 (O_894,N_19882,N_19639);
xor UO_895 (O_895,N_19814,N_19818);
xnor UO_896 (O_896,N_19822,N_19715);
and UO_897 (O_897,N_19980,N_19993);
nor UO_898 (O_898,N_19778,N_19927);
nor UO_899 (O_899,N_19961,N_19705);
nand UO_900 (O_900,N_19854,N_19842);
xnor UO_901 (O_901,N_19660,N_19617);
nor UO_902 (O_902,N_19886,N_19996);
or UO_903 (O_903,N_19663,N_19925);
nand UO_904 (O_904,N_19891,N_19992);
and UO_905 (O_905,N_19669,N_19767);
and UO_906 (O_906,N_19931,N_19603);
and UO_907 (O_907,N_19744,N_19637);
xor UO_908 (O_908,N_19973,N_19894);
or UO_909 (O_909,N_19897,N_19803);
nor UO_910 (O_910,N_19881,N_19948);
nor UO_911 (O_911,N_19921,N_19787);
nor UO_912 (O_912,N_19852,N_19977);
or UO_913 (O_913,N_19935,N_19714);
or UO_914 (O_914,N_19725,N_19966);
or UO_915 (O_915,N_19945,N_19947);
nand UO_916 (O_916,N_19930,N_19666);
xor UO_917 (O_917,N_19885,N_19667);
and UO_918 (O_918,N_19990,N_19956);
or UO_919 (O_919,N_19841,N_19879);
and UO_920 (O_920,N_19857,N_19793);
or UO_921 (O_921,N_19938,N_19852);
nor UO_922 (O_922,N_19882,N_19716);
nand UO_923 (O_923,N_19854,N_19998);
or UO_924 (O_924,N_19727,N_19979);
and UO_925 (O_925,N_19620,N_19884);
xor UO_926 (O_926,N_19970,N_19612);
nand UO_927 (O_927,N_19844,N_19868);
nand UO_928 (O_928,N_19737,N_19856);
or UO_929 (O_929,N_19747,N_19829);
and UO_930 (O_930,N_19798,N_19602);
and UO_931 (O_931,N_19835,N_19604);
nand UO_932 (O_932,N_19602,N_19847);
nand UO_933 (O_933,N_19823,N_19630);
xor UO_934 (O_934,N_19722,N_19619);
and UO_935 (O_935,N_19979,N_19757);
nand UO_936 (O_936,N_19928,N_19962);
or UO_937 (O_937,N_19745,N_19879);
nor UO_938 (O_938,N_19840,N_19716);
or UO_939 (O_939,N_19812,N_19665);
nor UO_940 (O_940,N_19729,N_19765);
or UO_941 (O_941,N_19690,N_19780);
nand UO_942 (O_942,N_19680,N_19966);
and UO_943 (O_943,N_19916,N_19682);
nand UO_944 (O_944,N_19691,N_19929);
xor UO_945 (O_945,N_19758,N_19914);
or UO_946 (O_946,N_19665,N_19916);
and UO_947 (O_947,N_19920,N_19835);
nor UO_948 (O_948,N_19602,N_19994);
and UO_949 (O_949,N_19705,N_19708);
and UO_950 (O_950,N_19705,N_19697);
or UO_951 (O_951,N_19929,N_19727);
nand UO_952 (O_952,N_19959,N_19934);
xor UO_953 (O_953,N_19989,N_19773);
or UO_954 (O_954,N_19800,N_19764);
nor UO_955 (O_955,N_19983,N_19683);
nor UO_956 (O_956,N_19912,N_19901);
nand UO_957 (O_957,N_19714,N_19814);
nand UO_958 (O_958,N_19806,N_19857);
nor UO_959 (O_959,N_19932,N_19670);
or UO_960 (O_960,N_19600,N_19841);
nand UO_961 (O_961,N_19811,N_19690);
xor UO_962 (O_962,N_19990,N_19846);
and UO_963 (O_963,N_19806,N_19988);
nand UO_964 (O_964,N_19756,N_19978);
and UO_965 (O_965,N_19916,N_19656);
xnor UO_966 (O_966,N_19667,N_19745);
xor UO_967 (O_967,N_19672,N_19928);
nand UO_968 (O_968,N_19820,N_19892);
nand UO_969 (O_969,N_19873,N_19980);
and UO_970 (O_970,N_19684,N_19633);
xnor UO_971 (O_971,N_19848,N_19837);
or UO_972 (O_972,N_19845,N_19687);
nor UO_973 (O_973,N_19902,N_19659);
or UO_974 (O_974,N_19680,N_19981);
or UO_975 (O_975,N_19656,N_19631);
nand UO_976 (O_976,N_19930,N_19683);
and UO_977 (O_977,N_19922,N_19780);
or UO_978 (O_978,N_19790,N_19649);
or UO_979 (O_979,N_19610,N_19928);
nor UO_980 (O_980,N_19982,N_19866);
nor UO_981 (O_981,N_19860,N_19666);
nand UO_982 (O_982,N_19706,N_19876);
and UO_983 (O_983,N_19913,N_19879);
nor UO_984 (O_984,N_19994,N_19858);
and UO_985 (O_985,N_19762,N_19659);
or UO_986 (O_986,N_19625,N_19783);
nor UO_987 (O_987,N_19953,N_19728);
and UO_988 (O_988,N_19672,N_19760);
nor UO_989 (O_989,N_19659,N_19638);
and UO_990 (O_990,N_19968,N_19868);
xor UO_991 (O_991,N_19784,N_19912);
xor UO_992 (O_992,N_19907,N_19992);
nand UO_993 (O_993,N_19850,N_19653);
or UO_994 (O_994,N_19605,N_19698);
xor UO_995 (O_995,N_19945,N_19741);
nand UO_996 (O_996,N_19954,N_19997);
or UO_997 (O_997,N_19894,N_19705);
xor UO_998 (O_998,N_19856,N_19922);
nand UO_999 (O_999,N_19986,N_19668);
and UO_1000 (O_1000,N_19641,N_19769);
and UO_1001 (O_1001,N_19852,N_19921);
or UO_1002 (O_1002,N_19979,N_19849);
and UO_1003 (O_1003,N_19900,N_19832);
nand UO_1004 (O_1004,N_19735,N_19825);
nor UO_1005 (O_1005,N_19619,N_19608);
nor UO_1006 (O_1006,N_19675,N_19889);
or UO_1007 (O_1007,N_19702,N_19615);
or UO_1008 (O_1008,N_19858,N_19863);
nand UO_1009 (O_1009,N_19693,N_19862);
and UO_1010 (O_1010,N_19822,N_19975);
nor UO_1011 (O_1011,N_19965,N_19673);
nor UO_1012 (O_1012,N_19863,N_19710);
nand UO_1013 (O_1013,N_19657,N_19947);
nor UO_1014 (O_1014,N_19727,N_19925);
or UO_1015 (O_1015,N_19931,N_19810);
and UO_1016 (O_1016,N_19861,N_19652);
nand UO_1017 (O_1017,N_19885,N_19659);
nand UO_1018 (O_1018,N_19806,N_19891);
xor UO_1019 (O_1019,N_19852,N_19984);
and UO_1020 (O_1020,N_19622,N_19634);
xor UO_1021 (O_1021,N_19815,N_19793);
nand UO_1022 (O_1022,N_19700,N_19951);
or UO_1023 (O_1023,N_19974,N_19778);
or UO_1024 (O_1024,N_19743,N_19875);
or UO_1025 (O_1025,N_19814,N_19843);
nor UO_1026 (O_1026,N_19790,N_19858);
nand UO_1027 (O_1027,N_19919,N_19620);
nand UO_1028 (O_1028,N_19744,N_19612);
or UO_1029 (O_1029,N_19726,N_19691);
and UO_1030 (O_1030,N_19935,N_19812);
nor UO_1031 (O_1031,N_19798,N_19646);
nor UO_1032 (O_1032,N_19893,N_19853);
or UO_1033 (O_1033,N_19925,N_19601);
nor UO_1034 (O_1034,N_19629,N_19935);
or UO_1035 (O_1035,N_19741,N_19687);
nand UO_1036 (O_1036,N_19921,N_19699);
or UO_1037 (O_1037,N_19791,N_19881);
nand UO_1038 (O_1038,N_19988,N_19840);
nand UO_1039 (O_1039,N_19631,N_19752);
xor UO_1040 (O_1040,N_19678,N_19882);
xor UO_1041 (O_1041,N_19633,N_19958);
xor UO_1042 (O_1042,N_19906,N_19819);
xor UO_1043 (O_1043,N_19711,N_19708);
and UO_1044 (O_1044,N_19928,N_19809);
xnor UO_1045 (O_1045,N_19723,N_19634);
nand UO_1046 (O_1046,N_19899,N_19640);
nor UO_1047 (O_1047,N_19775,N_19665);
nor UO_1048 (O_1048,N_19959,N_19618);
or UO_1049 (O_1049,N_19813,N_19849);
nand UO_1050 (O_1050,N_19710,N_19754);
nand UO_1051 (O_1051,N_19901,N_19887);
nor UO_1052 (O_1052,N_19688,N_19770);
and UO_1053 (O_1053,N_19666,N_19723);
and UO_1054 (O_1054,N_19870,N_19603);
and UO_1055 (O_1055,N_19911,N_19821);
nand UO_1056 (O_1056,N_19763,N_19687);
nor UO_1057 (O_1057,N_19913,N_19801);
and UO_1058 (O_1058,N_19772,N_19834);
xnor UO_1059 (O_1059,N_19906,N_19720);
or UO_1060 (O_1060,N_19851,N_19665);
nor UO_1061 (O_1061,N_19991,N_19838);
or UO_1062 (O_1062,N_19857,N_19927);
xor UO_1063 (O_1063,N_19899,N_19601);
xnor UO_1064 (O_1064,N_19649,N_19686);
nand UO_1065 (O_1065,N_19808,N_19880);
nand UO_1066 (O_1066,N_19695,N_19684);
nand UO_1067 (O_1067,N_19906,N_19849);
nand UO_1068 (O_1068,N_19616,N_19623);
nor UO_1069 (O_1069,N_19616,N_19628);
nand UO_1070 (O_1070,N_19960,N_19721);
or UO_1071 (O_1071,N_19883,N_19700);
and UO_1072 (O_1072,N_19856,N_19976);
xnor UO_1073 (O_1073,N_19627,N_19676);
nand UO_1074 (O_1074,N_19688,N_19984);
or UO_1075 (O_1075,N_19691,N_19715);
or UO_1076 (O_1076,N_19849,N_19916);
or UO_1077 (O_1077,N_19989,N_19645);
nand UO_1078 (O_1078,N_19865,N_19661);
or UO_1079 (O_1079,N_19791,N_19757);
nand UO_1080 (O_1080,N_19956,N_19604);
xor UO_1081 (O_1081,N_19919,N_19889);
nand UO_1082 (O_1082,N_19887,N_19722);
or UO_1083 (O_1083,N_19606,N_19941);
nor UO_1084 (O_1084,N_19941,N_19969);
xnor UO_1085 (O_1085,N_19912,N_19896);
xnor UO_1086 (O_1086,N_19765,N_19985);
xnor UO_1087 (O_1087,N_19894,N_19813);
xor UO_1088 (O_1088,N_19759,N_19644);
nand UO_1089 (O_1089,N_19626,N_19957);
nor UO_1090 (O_1090,N_19628,N_19708);
and UO_1091 (O_1091,N_19973,N_19970);
nand UO_1092 (O_1092,N_19928,N_19816);
nand UO_1093 (O_1093,N_19846,N_19637);
nand UO_1094 (O_1094,N_19698,N_19981);
and UO_1095 (O_1095,N_19965,N_19891);
nand UO_1096 (O_1096,N_19716,N_19792);
and UO_1097 (O_1097,N_19736,N_19724);
or UO_1098 (O_1098,N_19994,N_19610);
or UO_1099 (O_1099,N_19879,N_19882);
and UO_1100 (O_1100,N_19894,N_19988);
or UO_1101 (O_1101,N_19900,N_19813);
nor UO_1102 (O_1102,N_19749,N_19890);
xor UO_1103 (O_1103,N_19797,N_19643);
nor UO_1104 (O_1104,N_19697,N_19615);
nand UO_1105 (O_1105,N_19772,N_19777);
nor UO_1106 (O_1106,N_19673,N_19975);
nand UO_1107 (O_1107,N_19674,N_19712);
nor UO_1108 (O_1108,N_19747,N_19898);
xor UO_1109 (O_1109,N_19852,N_19882);
or UO_1110 (O_1110,N_19949,N_19666);
nand UO_1111 (O_1111,N_19806,N_19827);
or UO_1112 (O_1112,N_19752,N_19886);
and UO_1113 (O_1113,N_19901,N_19704);
xor UO_1114 (O_1114,N_19966,N_19658);
nor UO_1115 (O_1115,N_19899,N_19938);
and UO_1116 (O_1116,N_19828,N_19671);
nand UO_1117 (O_1117,N_19957,N_19690);
xor UO_1118 (O_1118,N_19829,N_19801);
xor UO_1119 (O_1119,N_19710,N_19783);
nand UO_1120 (O_1120,N_19737,N_19877);
and UO_1121 (O_1121,N_19630,N_19836);
xor UO_1122 (O_1122,N_19879,N_19914);
and UO_1123 (O_1123,N_19972,N_19758);
or UO_1124 (O_1124,N_19613,N_19969);
nor UO_1125 (O_1125,N_19940,N_19613);
nor UO_1126 (O_1126,N_19939,N_19865);
xnor UO_1127 (O_1127,N_19920,N_19811);
and UO_1128 (O_1128,N_19819,N_19647);
xnor UO_1129 (O_1129,N_19966,N_19751);
xor UO_1130 (O_1130,N_19882,N_19751);
and UO_1131 (O_1131,N_19685,N_19606);
or UO_1132 (O_1132,N_19784,N_19657);
nor UO_1133 (O_1133,N_19699,N_19933);
nand UO_1134 (O_1134,N_19614,N_19667);
or UO_1135 (O_1135,N_19713,N_19760);
or UO_1136 (O_1136,N_19768,N_19788);
xnor UO_1137 (O_1137,N_19772,N_19750);
or UO_1138 (O_1138,N_19827,N_19857);
and UO_1139 (O_1139,N_19631,N_19919);
or UO_1140 (O_1140,N_19917,N_19946);
nor UO_1141 (O_1141,N_19987,N_19812);
nor UO_1142 (O_1142,N_19904,N_19852);
nand UO_1143 (O_1143,N_19738,N_19990);
xor UO_1144 (O_1144,N_19630,N_19715);
or UO_1145 (O_1145,N_19605,N_19651);
xor UO_1146 (O_1146,N_19661,N_19853);
xnor UO_1147 (O_1147,N_19715,N_19679);
nand UO_1148 (O_1148,N_19612,N_19869);
nor UO_1149 (O_1149,N_19994,N_19983);
nor UO_1150 (O_1150,N_19758,N_19685);
xnor UO_1151 (O_1151,N_19832,N_19670);
nor UO_1152 (O_1152,N_19879,N_19822);
nor UO_1153 (O_1153,N_19744,N_19968);
xnor UO_1154 (O_1154,N_19603,N_19805);
and UO_1155 (O_1155,N_19817,N_19798);
xnor UO_1156 (O_1156,N_19781,N_19873);
xnor UO_1157 (O_1157,N_19687,N_19684);
xor UO_1158 (O_1158,N_19891,N_19691);
and UO_1159 (O_1159,N_19673,N_19967);
and UO_1160 (O_1160,N_19918,N_19771);
nor UO_1161 (O_1161,N_19828,N_19817);
and UO_1162 (O_1162,N_19844,N_19680);
xor UO_1163 (O_1163,N_19803,N_19614);
nor UO_1164 (O_1164,N_19657,N_19615);
nor UO_1165 (O_1165,N_19821,N_19865);
or UO_1166 (O_1166,N_19617,N_19775);
or UO_1167 (O_1167,N_19726,N_19624);
nor UO_1168 (O_1168,N_19915,N_19670);
nand UO_1169 (O_1169,N_19832,N_19691);
nand UO_1170 (O_1170,N_19843,N_19753);
or UO_1171 (O_1171,N_19694,N_19739);
and UO_1172 (O_1172,N_19876,N_19822);
nor UO_1173 (O_1173,N_19738,N_19870);
nand UO_1174 (O_1174,N_19874,N_19927);
or UO_1175 (O_1175,N_19887,N_19689);
and UO_1176 (O_1176,N_19820,N_19767);
nor UO_1177 (O_1177,N_19784,N_19801);
nor UO_1178 (O_1178,N_19669,N_19717);
xnor UO_1179 (O_1179,N_19618,N_19743);
xor UO_1180 (O_1180,N_19701,N_19951);
nor UO_1181 (O_1181,N_19775,N_19686);
xor UO_1182 (O_1182,N_19688,N_19902);
nor UO_1183 (O_1183,N_19623,N_19820);
nor UO_1184 (O_1184,N_19624,N_19712);
nor UO_1185 (O_1185,N_19802,N_19978);
nor UO_1186 (O_1186,N_19880,N_19925);
nand UO_1187 (O_1187,N_19881,N_19727);
and UO_1188 (O_1188,N_19695,N_19957);
nand UO_1189 (O_1189,N_19879,N_19693);
nor UO_1190 (O_1190,N_19661,N_19926);
nor UO_1191 (O_1191,N_19988,N_19855);
nor UO_1192 (O_1192,N_19892,N_19628);
nor UO_1193 (O_1193,N_19914,N_19862);
xnor UO_1194 (O_1194,N_19740,N_19737);
nand UO_1195 (O_1195,N_19621,N_19998);
nor UO_1196 (O_1196,N_19995,N_19605);
or UO_1197 (O_1197,N_19779,N_19689);
or UO_1198 (O_1198,N_19889,N_19627);
nand UO_1199 (O_1199,N_19966,N_19891);
nor UO_1200 (O_1200,N_19663,N_19741);
nand UO_1201 (O_1201,N_19718,N_19927);
nor UO_1202 (O_1202,N_19748,N_19963);
or UO_1203 (O_1203,N_19672,N_19655);
and UO_1204 (O_1204,N_19874,N_19839);
or UO_1205 (O_1205,N_19694,N_19706);
nand UO_1206 (O_1206,N_19705,N_19994);
xor UO_1207 (O_1207,N_19957,N_19987);
nand UO_1208 (O_1208,N_19988,N_19881);
and UO_1209 (O_1209,N_19791,N_19703);
and UO_1210 (O_1210,N_19888,N_19807);
and UO_1211 (O_1211,N_19606,N_19916);
nand UO_1212 (O_1212,N_19731,N_19815);
xnor UO_1213 (O_1213,N_19613,N_19982);
nor UO_1214 (O_1214,N_19935,N_19656);
nand UO_1215 (O_1215,N_19664,N_19907);
or UO_1216 (O_1216,N_19945,N_19932);
xor UO_1217 (O_1217,N_19616,N_19860);
nand UO_1218 (O_1218,N_19821,N_19973);
xor UO_1219 (O_1219,N_19893,N_19913);
xnor UO_1220 (O_1220,N_19676,N_19873);
nand UO_1221 (O_1221,N_19603,N_19986);
xor UO_1222 (O_1222,N_19917,N_19619);
nor UO_1223 (O_1223,N_19988,N_19828);
or UO_1224 (O_1224,N_19818,N_19993);
or UO_1225 (O_1225,N_19815,N_19956);
xnor UO_1226 (O_1226,N_19754,N_19897);
xor UO_1227 (O_1227,N_19768,N_19790);
nor UO_1228 (O_1228,N_19780,N_19670);
nor UO_1229 (O_1229,N_19815,N_19764);
nand UO_1230 (O_1230,N_19689,N_19660);
xnor UO_1231 (O_1231,N_19960,N_19972);
nor UO_1232 (O_1232,N_19630,N_19815);
nor UO_1233 (O_1233,N_19920,N_19945);
nand UO_1234 (O_1234,N_19622,N_19878);
nor UO_1235 (O_1235,N_19847,N_19931);
nor UO_1236 (O_1236,N_19636,N_19697);
nand UO_1237 (O_1237,N_19694,N_19902);
and UO_1238 (O_1238,N_19815,N_19741);
or UO_1239 (O_1239,N_19780,N_19901);
and UO_1240 (O_1240,N_19859,N_19769);
nor UO_1241 (O_1241,N_19811,N_19736);
nand UO_1242 (O_1242,N_19798,N_19937);
nor UO_1243 (O_1243,N_19900,N_19779);
and UO_1244 (O_1244,N_19643,N_19791);
xor UO_1245 (O_1245,N_19767,N_19962);
xor UO_1246 (O_1246,N_19645,N_19664);
nor UO_1247 (O_1247,N_19740,N_19958);
and UO_1248 (O_1248,N_19895,N_19908);
nor UO_1249 (O_1249,N_19918,N_19756);
nor UO_1250 (O_1250,N_19946,N_19618);
or UO_1251 (O_1251,N_19860,N_19620);
or UO_1252 (O_1252,N_19645,N_19979);
and UO_1253 (O_1253,N_19874,N_19850);
nand UO_1254 (O_1254,N_19804,N_19916);
nand UO_1255 (O_1255,N_19675,N_19997);
nor UO_1256 (O_1256,N_19827,N_19750);
xor UO_1257 (O_1257,N_19799,N_19852);
or UO_1258 (O_1258,N_19691,N_19967);
xnor UO_1259 (O_1259,N_19729,N_19691);
nor UO_1260 (O_1260,N_19704,N_19985);
and UO_1261 (O_1261,N_19906,N_19823);
xnor UO_1262 (O_1262,N_19965,N_19688);
nand UO_1263 (O_1263,N_19819,N_19758);
nor UO_1264 (O_1264,N_19910,N_19964);
nor UO_1265 (O_1265,N_19664,N_19982);
xor UO_1266 (O_1266,N_19954,N_19839);
or UO_1267 (O_1267,N_19768,N_19886);
and UO_1268 (O_1268,N_19652,N_19969);
nand UO_1269 (O_1269,N_19928,N_19867);
or UO_1270 (O_1270,N_19797,N_19937);
and UO_1271 (O_1271,N_19839,N_19781);
xor UO_1272 (O_1272,N_19852,N_19640);
or UO_1273 (O_1273,N_19997,N_19698);
nor UO_1274 (O_1274,N_19756,N_19764);
and UO_1275 (O_1275,N_19792,N_19619);
nand UO_1276 (O_1276,N_19700,N_19956);
nor UO_1277 (O_1277,N_19886,N_19877);
nand UO_1278 (O_1278,N_19734,N_19674);
or UO_1279 (O_1279,N_19903,N_19918);
or UO_1280 (O_1280,N_19762,N_19652);
nor UO_1281 (O_1281,N_19697,N_19991);
and UO_1282 (O_1282,N_19956,N_19952);
nor UO_1283 (O_1283,N_19878,N_19864);
nand UO_1284 (O_1284,N_19951,N_19974);
and UO_1285 (O_1285,N_19819,N_19895);
xor UO_1286 (O_1286,N_19844,N_19823);
nor UO_1287 (O_1287,N_19719,N_19618);
or UO_1288 (O_1288,N_19907,N_19604);
and UO_1289 (O_1289,N_19960,N_19927);
or UO_1290 (O_1290,N_19664,N_19900);
nor UO_1291 (O_1291,N_19941,N_19743);
xor UO_1292 (O_1292,N_19708,N_19799);
nor UO_1293 (O_1293,N_19907,N_19766);
or UO_1294 (O_1294,N_19852,N_19630);
or UO_1295 (O_1295,N_19600,N_19633);
or UO_1296 (O_1296,N_19825,N_19978);
xor UO_1297 (O_1297,N_19848,N_19916);
or UO_1298 (O_1298,N_19666,N_19609);
nand UO_1299 (O_1299,N_19859,N_19985);
xnor UO_1300 (O_1300,N_19917,N_19759);
nor UO_1301 (O_1301,N_19896,N_19825);
nor UO_1302 (O_1302,N_19720,N_19694);
or UO_1303 (O_1303,N_19938,N_19634);
and UO_1304 (O_1304,N_19980,N_19687);
nor UO_1305 (O_1305,N_19633,N_19859);
or UO_1306 (O_1306,N_19805,N_19794);
xor UO_1307 (O_1307,N_19813,N_19686);
xnor UO_1308 (O_1308,N_19695,N_19852);
and UO_1309 (O_1309,N_19681,N_19987);
nand UO_1310 (O_1310,N_19619,N_19609);
and UO_1311 (O_1311,N_19820,N_19707);
or UO_1312 (O_1312,N_19627,N_19810);
nand UO_1313 (O_1313,N_19805,N_19604);
or UO_1314 (O_1314,N_19622,N_19887);
nand UO_1315 (O_1315,N_19659,N_19927);
nor UO_1316 (O_1316,N_19874,N_19957);
nand UO_1317 (O_1317,N_19889,N_19838);
nor UO_1318 (O_1318,N_19798,N_19943);
nor UO_1319 (O_1319,N_19718,N_19811);
or UO_1320 (O_1320,N_19801,N_19675);
or UO_1321 (O_1321,N_19663,N_19682);
xnor UO_1322 (O_1322,N_19621,N_19824);
and UO_1323 (O_1323,N_19663,N_19618);
nand UO_1324 (O_1324,N_19837,N_19844);
nand UO_1325 (O_1325,N_19881,N_19903);
and UO_1326 (O_1326,N_19895,N_19913);
or UO_1327 (O_1327,N_19946,N_19709);
nand UO_1328 (O_1328,N_19969,N_19917);
or UO_1329 (O_1329,N_19917,N_19750);
and UO_1330 (O_1330,N_19794,N_19915);
or UO_1331 (O_1331,N_19839,N_19618);
nor UO_1332 (O_1332,N_19647,N_19827);
or UO_1333 (O_1333,N_19629,N_19988);
nand UO_1334 (O_1334,N_19601,N_19784);
nor UO_1335 (O_1335,N_19971,N_19990);
xnor UO_1336 (O_1336,N_19861,N_19844);
nand UO_1337 (O_1337,N_19734,N_19851);
and UO_1338 (O_1338,N_19913,N_19990);
nand UO_1339 (O_1339,N_19716,N_19741);
nor UO_1340 (O_1340,N_19618,N_19985);
and UO_1341 (O_1341,N_19811,N_19976);
or UO_1342 (O_1342,N_19943,N_19900);
or UO_1343 (O_1343,N_19834,N_19611);
and UO_1344 (O_1344,N_19747,N_19795);
or UO_1345 (O_1345,N_19930,N_19651);
nor UO_1346 (O_1346,N_19865,N_19743);
xor UO_1347 (O_1347,N_19660,N_19813);
and UO_1348 (O_1348,N_19812,N_19699);
xnor UO_1349 (O_1349,N_19959,N_19986);
or UO_1350 (O_1350,N_19730,N_19685);
nand UO_1351 (O_1351,N_19979,N_19826);
and UO_1352 (O_1352,N_19771,N_19693);
nor UO_1353 (O_1353,N_19657,N_19880);
or UO_1354 (O_1354,N_19786,N_19668);
nand UO_1355 (O_1355,N_19681,N_19787);
nand UO_1356 (O_1356,N_19752,N_19760);
nor UO_1357 (O_1357,N_19944,N_19970);
xnor UO_1358 (O_1358,N_19728,N_19954);
nand UO_1359 (O_1359,N_19663,N_19817);
or UO_1360 (O_1360,N_19662,N_19760);
xor UO_1361 (O_1361,N_19745,N_19750);
or UO_1362 (O_1362,N_19631,N_19679);
and UO_1363 (O_1363,N_19893,N_19869);
nand UO_1364 (O_1364,N_19843,N_19800);
xnor UO_1365 (O_1365,N_19669,N_19900);
nor UO_1366 (O_1366,N_19764,N_19782);
xnor UO_1367 (O_1367,N_19647,N_19770);
xnor UO_1368 (O_1368,N_19684,N_19842);
xor UO_1369 (O_1369,N_19804,N_19961);
nor UO_1370 (O_1370,N_19892,N_19782);
nand UO_1371 (O_1371,N_19682,N_19667);
nand UO_1372 (O_1372,N_19782,N_19904);
nand UO_1373 (O_1373,N_19788,N_19675);
nor UO_1374 (O_1374,N_19949,N_19889);
nand UO_1375 (O_1375,N_19737,N_19946);
or UO_1376 (O_1376,N_19747,N_19740);
or UO_1377 (O_1377,N_19615,N_19711);
nor UO_1378 (O_1378,N_19729,N_19911);
xnor UO_1379 (O_1379,N_19920,N_19855);
xnor UO_1380 (O_1380,N_19719,N_19797);
xnor UO_1381 (O_1381,N_19997,N_19899);
and UO_1382 (O_1382,N_19906,N_19696);
nor UO_1383 (O_1383,N_19674,N_19908);
xor UO_1384 (O_1384,N_19857,N_19951);
nor UO_1385 (O_1385,N_19709,N_19650);
and UO_1386 (O_1386,N_19626,N_19966);
nand UO_1387 (O_1387,N_19774,N_19700);
and UO_1388 (O_1388,N_19827,N_19826);
xnor UO_1389 (O_1389,N_19607,N_19746);
nand UO_1390 (O_1390,N_19916,N_19758);
xnor UO_1391 (O_1391,N_19726,N_19967);
and UO_1392 (O_1392,N_19863,N_19786);
or UO_1393 (O_1393,N_19820,N_19876);
xor UO_1394 (O_1394,N_19742,N_19899);
nor UO_1395 (O_1395,N_19887,N_19951);
nor UO_1396 (O_1396,N_19613,N_19728);
xor UO_1397 (O_1397,N_19981,N_19611);
or UO_1398 (O_1398,N_19951,N_19890);
xnor UO_1399 (O_1399,N_19759,N_19855);
nor UO_1400 (O_1400,N_19619,N_19955);
nand UO_1401 (O_1401,N_19916,N_19810);
nand UO_1402 (O_1402,N_19876,N_19812);
nor UO_1403 (O_1403,N_19745,N_19786);
xor UO_1404 (O_1404,N_19601,N_19901);
nor UO_1405 (O_1405,N_19655,N_19644);
or UO_1406 (O_1406,N_19685,N_19795);
nand UO_1407 (O_1407,N_19741,N_19854);
or UO_1408 (O_1408,N_19832,N_19895);
or UO_1409 (O_1409,N_19646,N_19677);
or UO_1410 (O_1410,N_19936,N_19788);
nor UO_1411 (O_1411,N_19713,N_19722);
nand UO_1412 (O_1412,N_19673,N_19739);
and UO_1413 (O_1413,N_19671,N_19845);
nor UO_1414 (O_1414,N_19742,N_19666);
or UO_1415 (O_1415,N_19856,N_19750);
or UO_1416 (O_1416,N_19643,N_19945);
nand UO_1417 (O_1417,N_19727,N_19662);
nand UO_1418 (O_1418,N_19750,N_19819);
nor UO_1419 (O_1419,N_19969,N_19933);
and UO_1420 (O_1420,N_19821,N_19725);
xor UO_1421 (O_1421,N_19773,N_19668);
nand UO_1422 (O_1422,N_19904,N_19752);
and UO_1423 (O_1423,N_19929,N_19814);
and UO_1424 (O_1424,N_19699,N_19955);
nor UO_1425 (O_1425,N_19776,N_19976);
nor UO_1426 (O_1426,N_19868,N_19783);
nor UO_1427 (O_1427,N_19783,N_19627);
or UO_1428 (O_1428,N_19795,N_19691);
or UO_1429 (O_1429,N_19760,N_19737);
and UO_1430 (O_1430,N_19761,N_19684);
xnor UO_1431 (O_1431,N_19938,N_19620);
nor UO_1432 (O_1432,N_19604,N_19633);
or UO_1433 (O_1433,N_19616,N_19920);
nand UO_1434 (O_1434,N_19898,N_19906);
nand UO_1435 (O_1435,N_19806,N_19745);
or UO_1436 (O_1436,N_19858,N_19627);
and UO_1437 (O_1437,N_19683,N_19671);
xnor UO_1438 (O_1438,N_19792,N_19748);
xor UO_1439 (O_1439,N_19965,N_19663);
xnor UO_1440 (O_1440,N_19803,N_19760);
nand UO_1441 (O_1441,N_19658,N_19931);
nor UO_1442 (O_1442,N_19887,N_19928);
and UO_1443 (O_1443,N_19890,N_19652);
nand UO_1444 (O_1444,N_19756,N_19600);
and UO_1445 (O_1445,N_19659,N_19858);
xnor UO_1446 (O_1446,N_19981,N_19817);
nand UO_1447 (O_1447,N_19849,N_19682);
xnor UO_1448 (O_1448,N_19791,N_19607);
xnor UO_1449 (O_1449,N_19953,N_19758);
or UO_1450 (O_1450,N_19994,N_19791);
nor UO_1451 (O_1451,N_19895,N_19692);
and UO_1452 (O_1452,N_19656,N_19742);
and UO_1453 (O_1453,N_19616,N_19630);
nand UO_1454 (O_1454,N_19935,N_19789);
nand UO_1455 (O_1455,N_19924,N_19829);
xnor UO_1456 (O_1456,N_19640,N_19603);
or UO_1457 (O_1457,N_19663,N_19771);
nor UO_1458 (O_1458,N_19778,N_19627);
and UO_1459 (O_1459,N_19854,N_19689);
nor UO_1460 (O_1460,N_19875,N_19814);
or UO_1461 (O_1461,N_19686,N_19810);
xor UO_1462 (O_1462,N_19686,N_19856);
or UO_1463 (O_1463,N_19669,N_19736);
nand UO_1464 (O_1464,N_19855,N_19762);
nand UO_1465 (O_1465,N_19789,N_19793);
nand UO_1466 (O_1466,N_19696,N_19639);
xnor UO_1467 (O_1467,N_19805,N_19938);
xor UO_1468 (O_1468,N_19690,N_19809);
or UO_1469 (O_1469,N_19932,N_19838);
xor UO_1470 (O_1470,N_19713,N_19679);
xor UO_1471 (O_1471,N_19837,N_19712);
and UO_1472 (O_1472,N_19943,N_19810);
xnor UO_1473 (O_1473,N_19673,N_19800);
and UO_1474 (O_1474,N_19873,N_19754);
nor UO_1475 (O_1475,N_19816,N_19880);
nor UO_1476 (O_1476,N_19925,N_19859);
or UO_1477 (O_1477,N_19688,N_19659);
xor UO_1478 (O_1478,N_19839,N_19884);
or UO_1479 (O_1479,N_19714,N_19679);
xor UO_1480 (O_1480,N_19770,N_19897);
xnor UO_1481 (O_1481,N_19902,N_19721);
nand UO_1482 (O_1482,N_19998,N_19646);
and UO_1483 (O_1483,N_19851,N_19684);
nand UO_1484 (O_1484,N_19617,N_19953);
xnor UO_1485 (O_1485,N_19738,N_19800);
and UO_1486 (O_1486,N_19924,N_19810);
nand UO_1487 (O_1487,N_19774,N_19601);
nand UO_1488 (O_1488,N_19688,N_19784);
or UO_1489 (O_1489,N_19785,N_19849);
nor UO_1490 (O_1490,N_19835,N_19643);
or UO_1491 (O_1491,N_19676,N_19837);
nand UO_1492 (O_1492,N_19758,N_19826);
xnor UO_1493 (O_1493,N_19856,N_19860);
xor UO_1494 (O_1494,N_19683,N_19857);
nand UO_1495 (O_1495,N_19647,N_19847);
or UO_1496 (O_1496,N_19721,N_19613);
and UO_1497 (O_1497,N_19691,N_19895);
and UO_1498 (O_1498,N_19875,N_19651);
and UO_1499 (O_1499,N_19910,N_19815);
xnor UO_1500 (O_1500,N_19928,N_19669);
xnor UO_1501 (O_1501,N_19610,N_19991);
xor UO_1502 (O_1502,N_19789,N_19958);
and UO_1503 (O_1503,N_19653,N_19821);
xor UO_1504 (O_1504,N_19705,N_19875);
xor UO_1505 (O_1505,N_19738,N_19728);
xnor UO_1506 (O_1506,N_19782,N_19679);
nand UO_1507 (O_1507,N_19684,N_19682);
nand UO_1508 (O_1508,N_19703,N_19906);
nand UO_1509 (O_1509,N_19856,N_19813);
nor UO_1510 (O_1510,N_19663,N_19782);
and UO_1511 (O_1511,N_19967,N_19893);
nand UO_1512 (O_1512,N_19893,N_19933);
nand UO_1513 (O_1513,N_19715,N_19758);
xor UO_1514 (O_1514,N_19998,N_19788);
xor UO_1515 (O_1515,N_19641,N_19929);
or UO_1516 (O_1516,N_19716,N_19873);
nor UO_1517 (O_1517,N_19965,N_19893);
or UO_1518 (O_1518,N_19819,N_19752);
and UO_1519 (O_1519,N_19742,N_19945);
xnor UO_1520 (O_1520,N_19993,N_19905);
xor UO_1521 (O_1521,N_19621,N_19958);
or UO_1522 (O_1522,N_19957,N_19840);
nor UO_1523 (O_1523,N_19706,N_19660);
or UO_1524 (O_1524,N_19920,N_19856);
or UO_1525 (O_1525,N_19828,N_19673);
and UO_1526 (O_1526,N_19767,N_19734);
and UO_1527 (O_1527,N_19789,N_19973);
or UO_1528 (O_1528,N_19988,N_19913);
and UO_1529 (O_1529,N_19911,N_19701);
nand UO_1530 (O_1530,N_19947,N_19771);
or UO_1531 (O_1531,N_19897,N_19891);
nor UO_1532 (O_1532,N_19712,N_19913);
and UO_1533 (O_1533,N_19872,N_19905);
or UO_1534 (O_1534,N_19856,N_19772);
nor UO_1535 (O_1535,N_19722,N_19670);
nor UO_1536 (O_1536,N_19692,N_19822);
or UO_1537 (O_1537,N_19604,N_19946);
nand UO_1538 (O_1538,N_19838,N_19640);
nor UO_1539 (O_1539,N_19877,N_19870);
or UO_1540 (O_1540,N_19949,N_19691);
nand UO_1541 (O_1541,N_19837,N_19897);
or UO_1542 (O_1542,N_19765,N_19908);
xnor UO_1543 (O_1543,N_19952,N_19878);
nand UO_1544 (O_1544,N_19971,N_19947);
and UO_1545 (O_1545,N_19662,N_19826);
xnor UO_1546 (O_1546,N_19915,N_19758);
and UO_1547 (O_1547,N_19644,N_19946);
xor UO_1548 (O_1548,N_19984,N_19610);
or UO_1549 (O_1549,N_19967,N_19957);
nand UO_1550 (O_1550,N_19699,N_19703);
or UO_1551 (O_1551,N_19990,N_19962);
nor UO_1552 (O_1552,N_19879,N_19760);
and UO_1553 (O_1553,N_19845,N_19705);
and UO_1554 (O_1554,N_19886,N_19984);
and UO_1555 (O_1555,N_19915,N_19671);
xor UO_1556 (O_1556,N_19787,N_19952);
nor UO_1557 (O_1557,N_19736,N_19892);
or UO_1558 (O_1558,N_19832,N_19835);
xnor UO_1559 (O_1559,N_19965,N_19953);
and UO_1560 (O_1560,N_19623,N_19663);
or UO_1561 (O_1561,N_19948,N_19947);
nand UO_1562 (O_1562,N_19912,N_19996);
or UO_1563 (O_1563,N_19754,N_19961);
and UO_1564 (O_1564,N_19971,N_19827);
or UO_1565 (O_1565,N_19682,N_19828);
nand UO_1566 (O_1566,N_19936,N_19800);
xor UO_1567 (O_1567,N_19675,N_19691);
xor UO_1568 (O_1568,N_19871,N_19734);
and UO_1569 (O_1569,N_19834,N_19858);
or UO_1570 (O_1570,N_19917,N_19734);
nor UO_1571 (O_1571,N_19611,N_19691);
nand UO_1572 (O_1572,N_19829,N_19953);
and UO_1573 (O_1573,N_19622,N_19631);
xor UO_1574 (O_1574,N_19885,N_19804);
nand UO_1575 (O_1575,N_19666,N_19832);
nand UO_1576 (O_1576,N_19951,N_19628);
nor UO_1577 (O_1577,N_19815,N_19646);
nor UO_1578 (O_1578,N_19618,N_19851);
xnor UO_1579 (O_1579,N_19909,N_19638);
xnor UO_1580 (O_1580,N_19716,N_19929);
nor UO_1581 (O_1581,N_19772,N_19721);
nor UO_1582 (O_1582,N_19742,N_19704);
nand UO_1583 (O_1583,N_19732,N_19954);
or UO_1584 (O_1584,N_19850,N_19603);
nor UO_1585 (O_1585,N_19819,N_19896);
or UO_1586 (O_1586,N_19680,N_19638);
nand UO_1587 (O_1587,N_19843,N_19606);
xnor UO_1588 (O_1588,N_19854,N_19945);
xor UO_1589 (O_1589,N_19637,N_19738);
xor UO_1590 (O_1590,N_19625,N_19637);
or UO_1591 (O_1591,N_19913,N_19723);
or UO_1592 (O_1592,N_19996,N_19899);
or UO_1593 (O_1593,N_19993,N_19799);
nor UO_1594 (O_1594,N_19834,N_19969);
nand UO_1595 (O_1595,N_19895,N_19664);
nor UO_1596 (O_1596,N_19985,N_19752);
nand UO_1597 (O_1597,N_19929,N_19640);
nor UO_1598 (O_1598,N_19769,N_19955);
nor UO_1599 (O_1599,N_19650,N_19808);
or UO_1600 (O_1600,N_19832,N_19811);
nor UO_1601 (O_1601,N_19835,N_19659);
nor UO_1602 (O_1602,N_19932,N_19611);
xnor UO_1603 (O_1603,N_19641,N_19790);
or UO_1604 (O_1604,N_19618,N_19634);
nand UO_1605 (O_1605,N_19631,N_19699);
nor UO_1606 (O_1606,N_19915,N_19718);
nor UO_1607 (O_1607,N_19723,N_19990);
nor UO_1608 (O_1608,N_19633,N_19784);
or UO_1609 (O_1609,N_19857,N_19988);
nand UO_1610 (O_1610,N_19725,N_19803);
xnor UO_1611 (O_1611,N_19993,N_19678);
or UO_1612 (O_1612,N_19624,N_19928);
nor UO_1613 (O_1613,N_19903,N_19611);
nand UO_1614 (O_1614,N_19753,N_19645);
or UO_1615 (O_1615,N_19768,N_19823);
and UO_1616 (O_1616,N_19724,N_19858);
nand UO_1617 (O_1617,N_19930,N_19647);
nor UO_1618 (O_1618,N_19921,N_19705);
nand UO_1619 (O_1619,N_19750,N_19611);
xor UO_1620 (O_1620,N_19672,N_19917);
and UO_1621 (O_1621,N_19656,N_19824);
xor UO_1622 (O_1622,N_19798,N_19839);
nand UO_1623 (O_1623,N_19765,N_19929);
nor UO_1624 (O_1624,N_19946,N_19962);
nor UO_1625 (O_1625,N_19746,N_19881);
nand UO_1626 (O_1626,N_19823,N_19759);
nand UO_1627 (O_1627,N_19812,N_19922);
nand UO_1628 (O_1628,N_19887,N_19707);
or UO_1629 (O_1629,N_19626,N_19736);
xnor UO_1630 (O_1630,N_19832,N_19702);
nand UO_1631 (O_1631,N_19741,N_19623);
nand UO_1632 (O_1632,N_19977,N_19940);
nand UO_1633 (O_1633,N_19631,N_19968);
and UO_1634 (O_1634,N_19824,N_19993);
nor UO_1635 (O_1635,N_19859,N_19764);
and UO_1636 (O_1636,N_19748,N_19831);
and UO_1637 (O_1637,N_19677,N_19886);
xor UO_1638 (O_1638,N_19655,N_19796);
or UO_1639 (O_1639,N_19877,N_19648);
or UO_1640 (O_1640,N_19855,N_19652);
nand UO_1641 (O_1641,N_19643,N_19786);
xnor UO_1642 (O_1642,N_19808,N_19862);
nand UO_1643 (O_1643,N_19886,N_19632);
nand UO_1644 (O_1644,N_19852,N_19660);
and UO_1645 (O_1645,N_19935,N_19701);
xnor UO_1646 (O_1646,N_19682,N_19941);
and UO_1647 (O_1647,N_19875,N_19619);
xor UO_1648 (O_1648,N_19778,N_19706);
and UO_1649 (O_1649,N_19862,N_19719);
and UO_1650 (O_1650,N_19831,N_19995);
or UO_1651 (O_1651,N_19760,N_19799);
and UO_1652 (O_1652,N_19721,N_19604);
nor UO_1653 (O_1653,N_19999,N_19949);
nor UO_1654 (O_1654,N_19652,N_19837);
nor UO_1655 (O_1655,N_19986,N_19811);
and UO_1656 (O_1656,N_19815,N_19655);
nand UO_1657 (O_1657,N_19989,N_19711);
xor UO_1658 (O_1658,N_19735,N_19833);
nor UO_1659 (O_1659,N_19992,N_19634);
nand UO_1660 (O_1660,N_19610,N_19893);
or UO_1661 (O_1661,N_19664,N_19958);
and UO_1662 (O_1662,N_19728,N_19851);
or UO_1663 (O_1663,N_19773,N_19665);
nand UO_1664 (O_1664,N_19766,N_19854);
xnor UO_1665 (O_1665,N_19785,N_19703);
nand UO_1666 (O_1666,N_19935,N_19770);
nand UO_1667 (O_1667,N_19772,N_19875);
or UO_1668 (O_1668,N_19694,N_19832);
xor UO_1669 (O_1669,N_19791,N_19807);
or UO_1670 (O_1670,N_19965,N_19840);
xor UO_1671 (O_1671,N_19871,N_19653);
xor UO_1672 (O_1672,N_19935,N_19614);
nor UO_1673 (O_1673,N_19643,N_19827);
nor UO_1674 (O_1674,N_19841,N_19681);
nand UO_1675 (O_1675,N_19863,N_19636);
nand UO_1676 (O_1676,N_19730,N_19880);
nor UO_1677 (O_1677,N_19802,N_19663);
nand UO_1678 (O_1678,N_19663,N_19938);
xor UO_1679 (O_1679,N_19639,N_19685);
nand UO_1680 (O_1680,N_19949,N_19823);
nor UO_1681 (O_1681,N_19702,N_19676);
xor UO_1682 (O_1682,N_19650,N_19959);
nor UO_1683 (O_1683,N_19732,N_19869);
nor UO_1684 (O_1684,N_19760,N_19917);
nand UO_1685 (O_1685,N_19712,N_19693);
nand UO_1686 (O_1686,N_19961,N_19716);
nand UO_1687 (O_1687,N_19959,N_19948);
xnor UO_1688 (O_1688,N_19868,N_19743);
and UO_1689 (O_1689,N_19623,N_19991);
and UO_1690 (O_1690,N_19828,N_19605);
nand UO_1691 (O_1691,N_19904,N_19786);
nor UO_1692 (O_1692,N_19886,N_19645);
and UO_1693 (O_1693,N_19924,N_19841);
nand UO_1694 (O_1694,N_19628,N_19692);
and UO_1695 (O_1695,N_19617,N_19726);
or UO_1696 (O_1696,N_19655,N_19603);
xor UO_1697 (O_1697,N_19614,N_19823);
xor UO_1698 (O_1698,N_19694,N_19958);
nand UO_1699 (O_1699,N_19938,N_19738);
nand UO_1700 (O_1700,N_19742,N_19793);
xor UO_1701 (O_1701,N_19613,N_19605);
and UO_1702 (O_1702,N_19725,N_19759);
or UO_1703 (O_1703,N_19951,N_19627);
xnor UO_1704 (O_1704,N_19645,N_19641);
nor UO_1705 (O_1705,N_19727,N_19986);
xor UO_1706 (O_1706,N_19875,N_19642);
and UO_1707 (O_1707,N_19701,N_19783);
nand UO_1708 (O_1708,N_19820,N_19852);
xor UO_1709 (O_1709,N_19971,N_19755);
and UO_1710 (O_1710,N_19859,N_19876);
or UO_1711 (O_1711,N_19752,N_19909);
and UO_1712 (O_1712,N_19983,N_19696);
xnor UO_1713 (O_1713,N_19829,N_19952);
xor UO_1714 (O_1714,N_19882,N_19698);
nor UO_1715 (O_1715,N_19654,N_19711);
and UO_1716 (O_1716,N_19941,N_19747);
or UO_1717 (O_1717,N_19946,N_19816);
and UO_1718 (O_1718,N_19997,N_19822);
and UO_1719 (O_1719,N_19716,N_19865);
and UO_1720 (O_1720,N_19810,N_19869);
nand UO_1721 (O_1721,N_19986,N_19770);
xor UO_1722 (O_1722,N_19980,N_19778);
or UO_1723 (O_1723,N_19797,N_19813);
or UO_1724 (O_1724,N_19644,N_19939);
and UO_1725 (O_1725,N_19692,N_19681);
nor UO_1726 (O_1726,N_19693,N_19807);
xor UO_1727 (O_1727,N_19680,N_19864);
and UO_1728 (O_1728,N_19804,N_19693);
nand UO_1729 (O_1729,N_19870,N_19971);
nor UO_1730 (O_1730,N_19672,N_19737);
or UO_1731 (O_1731,N_19856,N_19809);
nor UO_1732 (O_1732,N_19859,N_19668);
and UO_1733 (O_1733,N_19735,N_19660);
or UO_1734 (O_1734,N_19942,N_19871);
and UO_1735 (O_1735,N_19869,N_19703);
xor UO_1736 (O_1736,N_19713,N_19821);
nand UO_1737 (O_1737,N_19752,N_19735);
nand UO_1738 (O_1738,N_19720,N_19656);
nor UO_1739 (O_1739,N_19603,N_19668);
nor UO_1740 (O_1740,N_19700,N_19981);
xor UO_1741 (O_1741,N_19724,N_19618);
nor UO_1742 (O_1742,N_19980,N_19672);
nand UO_1743 (O_1743,N_19820,N_19873);
or UO_1744 (O_1744,N_19609,N_19856);
nand UO_1745 (O_1745,N_19776,N_19997);
and UO_1746 (O_1746,N_19797,N_19768);
xnor UO_1747 (O_1747,N_19953,N_19625);
or UO_1748 (O_1748,N_19887,N_19606);
and UO_1749 (O_1749,N_19717,N_19697);
nand UO_1750 (O_1750,N_19868,N_19752);
nor UO_1751 (O_1751,N_19871,N_19789);
nor UO_1752 (O_1752,N_19615,N_19613);
nand UO_1753 (O_1753,N_19638,N_19653);
or UO_1754 (O_1754,N_19844,N_19859);
xnor UO_1755 (O_1755,N_19752,N_19711);
and UO_1756 (O_1756,N_19773,N_19715);
and UO_1757 (O_1757,N_19609,N_19878);
and UO_1758 (O_1758,N_19820,N_19821);
or UO_1759 (O_1759,N_19718,N_19780);
nand UO_1760 (O_1760,N_19794,N_19723);
or UO_1761 (O_1761,N_19621,N_19815);
nand UO_1762 (O_1762,N_19811,N_19877);
and UO_1763 (O_1763,N_19779,N_19654);
xnor UO_1764 (O_1764,N_19988,N_19936);
and UO_1765 (O_1765,N_19875,N_19961);
nand UO_1766 (O_1766,N_19644,N_19887);
xnor UO_1767 (O_1767,N_19983,N_19927);
nand UO_1768 (O_1768,N_19948,N_19603);
or UO_1769 (O_1769,N_19795,N_19642);
and UO_1770 (O_1770,N_19717,N_19743);
nand UO_1771 (O_1771,N_19676,N_19830);
xnor UO_1772 (O_1772,N_19763,N_19970);
nor UO_1773 (O_1773,N_19855,N_19706);
nand UO_1774 (O_1774,N_19903,N_19899);
nand UO_1775 (O_1775,N_19907,N_19801);
xnor UO_1776 (O_1776,N_19608,N_19769);
xnor UO_1777 (O_1777,N_19708,N_19832);
or UO_1778 (O_1778,N_19725,N_19707);
or UO_1779 (O_1779,N_19834,N_19692);
nor UO_1780 (O_1780,N_19778,N_19983);
and UO_1781 (O_1781,N_19904,N_19698);
nor UO_1782 (O_1782,N_19873,N_19788);
and UO_1783 (O_1783,N_19669,N_19990);
nand UO_1784 (O_1784,N_19931,N_19905);
nand UO_1785 (O_1785,N_19795,N_19924);
nand UO_1786 (O_1786,N_19934,N_19984);
xnor UO_1787 (O_1787,N_19675,N_19670);
or UO_1788 (O_1788,N_19929,N_19902);
nand UO_1789 (O_1789,N_19707,N_19930);
nor UO_1790 (O_1790,N_19880,N_19946);
xnor UO_1791 (O_1791,N_19982,N_19870);
nand UO_1792 (O_1792,N_19629,N_19803);
nor UO_1793 (O_1793,N_19938,N_19659);
nand UO_1794 (O_1794,N_19848,N_19743);
xnor UO_1795 (O_1795,N_19727,N_19621);
nor UO_1796 (O_1796,N_19774,N_19647);
and UO_1797 (O_1797,N_19951,N_19782);
xnor UO_1798 (O_1798,N_19905,N_19928);
xor UO_1799 (O_1799,N_19875,N_19774);
nor UO_1800 (O_1800,N_19785,N_19998);
nand UO_1801 (O_1801,N_19677,N_19711);
xor UO_1802 (O_1802,N_19757,N_19957);
and UO_1803 (O_1803,N_19938,N_19820);
or UO_1804 (O_1804,N_19615,N_19792);
nor UO_1805 (O_1805,N_19951,N_19892);
or UO_1806 (O_1806,N_19799,N_19616);
nand UO_1807 (O_1807,N_19698,N_19845);
xor UO_1808 (O_1808,N_19702,N_19864);
or UO_1809 (O_1809,N_19933,N_19710);
xor UO_1810 (O_1810,N_19710,N_19818);
or UO_1811 (O_1811,N_19946,N_19724);
nand UO_1812 (O_1812,N_19755,N_19927);
xnor UO_1813 (O_1813,N_19886,N_19698);
nand UO_1814 (O_1814,N_19773,N_19830);
nand UO_1815 (O_1815,N_19636,N_19716);
xnor UO_1816 (O_1816,N_19877,N_19952);
nor UO_1817 (O_1817,N_19809,N_19611);
nand UO_1818 (O_1818,N_19762,N_19816);
xnor UO_1819 (O_1819,N_19762,N_19896);
nor UO_1820 (O_1820,N_19744,N_19941);
nor UO_1821 (O_1821,N_19998,N_19867);
nand UO_1822 (O_1822,N_19633,N_19661);
nand UO_1823 (O_1823,N_19667,N_19788);
nand UO_1824 (O_1824,N_19842,N_19833);
nand UO_1825 (O_1825,N_19816,N_19737);
and UO_1826 (O_1826,N_19605,N_19702);
xnor UO_1827 (O_1827,N_19933,N_19846);
xnor UO_1828 (O_1828,N_19684,N_19781);
or UO_1829 (O_1829,N_19716,N_19733);
nand UO_1830 (O_1830,N_19640,N_19710);
nor UO_1831 (O_1831,N_19699,N_19910);
nand UO_1832 (O_1832,N_19889,N_19641);
nand UO_1833 (O_1833,N_19906,N_19687);
and UO_1834 (O_1834,N_19634,N_19831);
nor UO_1835 (O_1835,N_19885,N_19709);
nand UO_1836 (O_1836,N_19653,N_19827);
or UO_1837 (O_1837,N_19662,N_19764);
nand UO_1838 (O_1838,N_19919,N_19880);
nand UO_1839 (O_1839,N_19816,N_19616);
and UO_1840 (O_1840,N_19896,N_19696);
xnor UO_1841 (O_1841,N_19748,N_19660);
nand UO_1842 (O_1842,N_19656,N_19835);
or UO_1843 (O_1843,N_19652,N_19741);
nand UO_1844 (O_1844,N_19805,N_19861);
or UO_1845 (O_1845,N_19680,N_19965);
nor UO_1846 (O_1846,N_19957,N_19980);
or UO_1847 (O_1847,N_19722,N_19648);
xor UO_1848 (O_1848,N_19758,N_19909);
nor UO_1849 (O_1849,N_19724,N_19790);
or UO_1850 (O_1850,N_19724,N_19942);
and UO_1851 (O_1851,N_19793,N_19921);
or UO_1852 (O_1852,N_19795,N_19905);
or UO_1853 (O_1853,N_19843,N_19951);
nand UO_1854 (O_1854,N_19952,N_19702);
nand UO_1855 (O_1855,N_19752,N_19812);
nand UO_1856 (O_1856,N_19923,N_19911);
nor UO_1857 (O_1857,N_19962,N_19670);
and UO_1858 (O_1858,N_19660,N_19907);
xnor UO_1859 (O_1859,N_19942,N_19931);
xor UO_1860 (O_1860,N_19604,N_19870);
xnor UO_1861 (O_1861,N_19636,N_19737);
and UO_1862 (O_1862,N_19902,N_19778);
or UO_1863 (O_1863,N_19938,N_19928);
nor UO_1864 (O_1864,N_19642,N_19633);
nor UO_1865 (O_1865,N_19620,N_19665);
xnor UO_1866 (O_1866,N_19866,N_19914);
and UO_1867 (O_1867,N_19689,N_19841);
nand UO_1868 (O_1868,N_19617,N_19714);
nand UO_1869 (O_1869,N_19775,N_19967);
or UO_1870 (O_1870,N_19734,N_19966);
or UO_1871 (O_1871,N_19610,N_19926);
xnor UO_1872 (O_1872,N_19855,N_19716);
nor UO_1873 (O_1873,N_19824,N_19662);
nor UO_1874 (O_1874,N_19742,N_19777);
or UO_1875 (O_1875,N_19867,N_19884);
or UO_1876 (O_1876,N_19850,N_19607);
or UO_1877 (O_1877,N_19866,N_19834);
or UO_1878 (O_1878,N_19710,N_19665);
xor UO_1879 (O_1879,N_19878,N_19840);
or UO_1880 (O_1880,N_19687,N_19690);
nor UO_1881 (O_1881,N_19700,N_19712);
nand UO_1882 (O_1882,N_19641,N_19908);
nor UO_1883 (O_1883,N_19634,N_19795);
or UO_1884 (O_1884,N_19990,N_19681);
and UO_1885 (O_1885,N_19967,N_19715);
and UO_1886 (O_1886,N_19619,N_19757);
or UO_1887 (O_1887,N_19635,N_19792);
xor UO_1888 (O_1888,N_19845,N_19895);
nor UO_1889 (O_1889,N_19815,N_19697);
xnor UO_1890 (O_1890,N_19918,N_19649);
xnor UO_1891 (O_1891,N_19945,N_19830);
or UO_1892 (O_1892,N_19867,N_19786);
nor UO_1893 (O_1893,N_19861,N_19780);
or UO_1894 (O_1894,N_19656,N_19621);
xor UO_1895 (O_1895,N_19642,N_19622);
nor UO_1896 (O_1896,N_19844,N_19808);
nor UO_1897 (O_1897,N_19833,N_19611);
xnor UO_1898 (O_1898,N_19929,N_19633);
and UO_1899 (O_1899,N_19698,N_19809);
xor UO_1900 (O_1900,N_19910,N_19707);
or UO_1901 (O_1901,N_19660,N_19841);
xnor UO_1902 (O_1902,N_19651,N_19933);
and UO_1903 (O_1903,N_19736,N_19838);
nand UO_1904 (O_1904,N_19614,N_19799);
nor UO_1905 (O_1905,N_19858,N_19672);
nand UO_1906 (O_1906,N_19972,N_19990);
nand UO_1907 (O_1907,N_19814,N_19698);
or UO_1908 (O_1908,N_19894,N_19942);
nand UO_1909 (O_1909,N_19909,N_19768);
and UO_1910 (O_1910,N_19913,N_19692);
or UO_1911 (O_1911,N_19835,N_19890);
xnor UO_1912 (O_1912,N_19752,N_19720);
or UO_1913 (O_1913,N_19994,N_19901);
nor UO_1914 (O_1914,N_19679,N_19706);
and UO_1915 (O_1915,N_19713,N_19851);
and UO_1916 (O_1916,N_19769,N_19952);
and UO_1917 (O_1917,N_19849,N_19829);
or UO_1918 (O_1918,N_19946,N_19671);
nand UO_1919 (O_1919,N_19756,N_19747);
or UO_1920 (O_1920,N_19945,N_19918);
nor UO_1921 (O_1921,N_19944,N_19677);
nand UO_1922 (O_1922,N_19602,N_19888);
nand UO_1923 (O_1923,N_19715,N_19867);
or UO_1924 (O_1924,N_19848,N_19894);
nand UO_1925 (O_1925,N_19740,N_19937);
nand UO_1926 (O_1926,N_19860,N_19788);
nand UO_1927 (O_1927,N_19828,N_19910);
or UO_1928 (O_1928,N_19616,N_19957);
nand UO_1929 (O_1929,N_19867,N_19910);
nand UO_1930 (O_1930,N_19828,N_19957);
nor UO_1931 (O_1931,N_19883,N_19713);
xor UO_1932 (O_1932,N_19809,N_19722);
nor UO_1933 (O_1933,N_19783,N_19937);
nor UO_1934 (O_1934,N_19871,N_19963);
xor UO_1935 (O_1935,N_19901,N_19716);
and UO_1936 (O_1936,N_19819,N_19970);
or UO_1937 (O_1937,N_19985,N_19986);
xor UO_1938 (O_1938,N_19823,N_19625);
nand UO_1939 (O_1939,N_19687,N_19908);
and UO_1940 (O_1940,N_19835,N_19885);
nand UO_1941 (O_1941,N_19680,N_19739);
and UO_1942 (O_1942,N_19808,N_19828);
xor UO_1943 (O_1943,N_19635,N_19769);
xnor UO_1944 (O_1944,N_19756,N_19844);
xnor UO_1945 (O_1945,N_19676,N_19715);
nor UO_1946 (O_1946,N_19700,N_19666);
or UO_1947 (O_1947,N_19687,N_19656);
xor UO_1948 (O_1948,N_19860,N_19726);
or UO_1949 (O_1949,N_19641,N_19668);
nor UO_1950 (O_1950,N_19927,N_19827);
xor UO_1951 (O_1951,N_19889,N_19937);
nand UO_1952 (O_1952,N_19984,N_19953);
nand UO_1953 (O_1953,N_19949,N_19985);
xor UO_1954 (O_1954,N_19986,N_19734);
nor UO_1955 (O_1955,N_19817,N_19662);
nand UO_1956 (O_1956,N_19646,N_19617);
xor UO_1957 (O_1957,N_19699,N_19869);
and UO_1958 (O_1958,N_19826,N_19940);
nor UO_1959 (O_1959,N_19697,N_19972);
nor UO_1960 (O_1960,N_19810,N_19991);
nand UO_1961 (O_1961,N_19749,N_19981);
nor UO_1962 (O_1962,N_19665,N_19855);
xor UO_1963 (O_1963,N_19655,N_19701);
or UO_1964 (O_1964,N_19830,N_19911);
or UO_1965 (O_1965,N_19760,N_19969);
nand UO_1966 (O_1966,N_19703,N_19819);
nand UO_1967 (O_1967,N_19875,N_19693);
and UO_1968 (O_1968,N_19990,N_19651);
nand UO_1969 (O_1969,N_19783,N_19672);
nor UO_1970 (O_1970,N_19765,N_19934);
and UO_1971 (O_1971,N_19621,N_19855);
and UO_1972 (O_1972,N_19951,N_19967);
xnor UO_1973 (O_1973,N_19886,N_19843);
or UO_1974 (O_1974,N_19983,N_19620);
nor UO_1975 (O_1975,N_19623,N_19861);
or UO_1976 (O_1976,N_19863,N_19737);
nor UO_1977 (O_1977,N_19658,N_19902);
and UO_1978 (O_1978,N_19834,N_19874);
nand UO_1979 (O_1979,N_19669,N_19890);
nand UO_1980 (O_1980,N_19873,N_19776);
xnor UO_1981 (O_1981,N_19985,N_19698);
nand UO_1982 (O_1982,N_19737,N_19632);
or UO_1983 (O_1983,N_19955,N_19923);
and UO_1984 (O_1984,N_19982,N_19703);
xor UO_1985 (O_1985,N_19687,N_19953);
xor UO_1986 (O_1986,N_19877,N_19895);
nor UO_1987 (O_1987,N_19868,N_19911);
nor UO_1988 (O_1988,N_19951,N_19793);
nand UO_1989 (O_1989,N_19944,N_19866);
or UO_1990 (O_1990,N_19923,N_19706);
nor UO_1991 (O_1991,N_19669,N_19861);
nand UO_1992 (O_1992,N_19753,N_19784);
and UO_1993 (O_1993,N_19723,N_19752);
or UO_1994 (O_1994,N_19720,N_19855);
nand UO_1995 (O_1995,N_19700,N_19852);
nor UO_1996 (O_1996,N_19740,N_19720);
and UO_1997 (O_1997,N_19803,N_19640);
or UO_1998 (O_1998,N_19613,N_19825);
nor UO_1999 (O_1999,N_19754,N_19821);
and UO_2000 (O_2000,N_19757,N_19848);
nor UO_2001 (O_2001,N_19968,N_19689);
nor UO_2002 (O_2002,N_19721,N_19647);
and UO_2003 (O_2003,N_19916,N_19954);
and UO_2004 (O_2004,N_19673,N_19883);
nand UO_2005 (O_2005,N_19636,N_19893);
or UO_2006 (O_2006,N_19645,N_19826);
nand UO_2007 (O_2007,N_19663,N_19851);
xnor UO_2008 (O_2008,N_19674,N_19909);
or UO_2009 (O_2009,N_19675,N_19850);
xnor UO_2010 (O_2010,N_19641,N_19795);
xor UO_2011 (O_2011,N_19981,N_19603);
xor UO_2012 (O_2012,N_19924,N_19931);
xor UO_2013 (O_2013,N_19800,N_19789);
nor UO_2014 (O_2014,N_19768,N_19760);
and UO_2015 (O_2015,N_19695,N_19915);
nor UO_2016 (O_2016,N_19965,N_19748);
or UO_2017 (O_2017,N_19859,N_19747);
xnor UO_2018 (O_2018,N_19656,N_19979);
xnor UO_2019 (O_2019,N_19809,N_19821);
nand UO_2020 (O_2020,N_19950,N_19712);
nor UO_2021 (O_2021,N_19704,N_19603);
nor UO_2022 (O_2022,N_19808,N_19744);
nand UO_2023 (O_2023,N_19633,N_19687);
nor UO_2024 (O_2024,N_19625,N_19694);
or UO_2025 (O_2025,N_19758,N_19648);
nor UO_2026 (O_2026,N_19847,N_19680);
xor UO_2027 (O_2027,N_19622,N_19823);
and UO_2028 (O_2028,N_19707,N_19906);
or UO_2029 (O_2029,N_19962,N_19634);
and UO_2030 (O_2030,N_19706,N_19958);
xor UO_2031 (O_2031,N_19729,N_19967);
and UO_2032 (O_2032,N_19981,N_19873);
and UO_2033 (O_2033,N_19659,N_19819);
nor UO_2034 (O_2034,N_19633,N_19847);
and UO_2035 (O_2035,N_19944,N_19932);
and UO_2036 (O_2036,N_19651,N_19880);
or UO_2037 (O_2037,N_19847,N_19771);
nor UO_2038 (O_2038,N_19679,N_19830);
xor UO_2039 (O_2039,N_19783,N_19770);
xnor UO_2040 (O_2040,N_19870,N_19778);
xnor UO_2041 (O_2041,N_19809,N_19990);
xor UO_2042 (O_2042,N_19632,N_19708);
nor UO_2043 (O_2043,N_19945,N_19717);
nand UO_2044 (O_2044,N_19865,N_19901);
or UO_2045 (O_2045,N_19933,N_19678);
xnor UO_2046 (O_2046,N_19971,N_19770);
nand UO_2047 (O_2047,N_19639,N_19768);
and UO_2048 (O_2048,N_19784,N_19741);
nand UO_2049 (O_2049,N_19731,N_19635);
or UO_2050 (O_2050,N_19606,N_19734);
and UO_2051 (O_2051,N_19647,N_19642);
xor UO_2052 (O_2052,N_19737,N_19867);
nor UO_2053 (O_2053,N_19990,N_19674);
nor UO_2054 (O_2054,N_19756,N_19977);
nand UO_2055 (O_2055,N_19663,N_19945);
nand UO_2056 (O_2056,N_19684,N_19707);
or UO_2057 (O_2057,N_19851,N_19808);
or UO_2058 (O_2058,N_19938,N_19922);
and UO_2059 (O_2059,N_19950,N_19628);
and UO_2060 (O_2060,N_19725,N_19734);
xor UO_2061 (O_2061,N_19833,N_19633);
and UO_2062 (O_2062,N_19688,N_19840);
nand UO_2063 (O_2063,N_19926,N_19767);
or UO_2064 (O_2064,N_19809,N_19955);
and UO_2065 (O_2065,N_19862,N_19695);
and UO_2066 (O_2066,N_19744,N_19817);
xor UO_2067 (O_2067,N_19625,N_19764);
nor UO_2068 (O_2068,N_19667,N_19704);
xor UO_2069 (O_2069,N_19833,N_19636);
nor UO_2070 (O_2070,N_19751,N_19867);
and UO_2071 (O_2071,N_19722,N_19996);
or UO_2072 (O_2072,N_19775,N_19654);
nand UO_2073 (O_2073,N_19713,N_19819);
xor UO_2074 (O_2074,N_19750,N_19860);
and UO_2075 (O_2075,N_19735,N_19820);
and UO_2076 (O_2076,N_19769,N_19918);
and UO_2077 (O_2077,N_19855,N_19907);
nand UO_2078 (O_2078,N_19828,N_19688);
and UO_2079 (O_2079,N_19665,N_19663);
xnor UO_2080 (O_2080,N_19733,N_19802);
or UO_2081 (O_2081,N_19837,N_19858);
xor UO_2082 (O_2082,N_19873,N_19734);
or UO_2083 (O_2083,N_19784,N_19749);
nand UO_2084 (O_2084,N_19801,N_19728);
xnor UO_2085 (O_2085,N_19753,N_19615);
xnor UO_2086 (O_2086,N_19807,N_19929);
xnor UO_2087 (O_2087,N_19634,N_19837);
and UO_2088 (O_2088,N_19938,N_19801);
xnor UO_2089 (O_2089,N_19800,N_19790);
xor UO_2090 (O_2090,N_19781,N_19940);
nor UO_2091 (O_2091,N_19865,N_19775);
nor UO_2092 (O_2092,N_19637,N_19814);
or UO_2093 (O_2093,N_19964,N_19799);
nor UO_2094 (O_2094,N_19827,N_19977);
or UO_2095 (O_2095,N_19849,N_19903);
nand UO_2096 (O_2096,N_19869,N_19849);
and UO_2097 (O_2097,N_19662,N_19629);
nand UO_2098 (O_2098,N_19618,N_19602);
nor UO_2099 (O_2099,N_19975,N_19845);
nand UO_2100 (O_2100,N_19707,N_19895);
xnor UO_2101 (O_2101,N_19621,N_19894);
nand UO_2102 (O_2102,N_19698,N_19894);
nand UO_2103 (O_2103,N_19950,N_19731);
nor UO_2104 (O_2104,N_19924,N_19944);
nand UO_2105 (O_2105,N_19736,N_19623);
or UO_2106 (O_2106,N_19902,N_19810);
nor UO_2107 (O_2107,N_19989,N_19873);
xor UO_2108 (O_2108,N_19876,N_19978);
nand UO_2109 (O_2109,N_19998,N_19617);
nand UO_2110 (O_2110,N_19602,N_19816);
or UO_2111 (O_2111,N_19999,N_19608);
and UO_2112 (O_2112,N_19721,N_19886);
xnor UO_2113 (O_2113,N_19847,N_19786);
nand UO_2114 (O_2114,N_19729,N_19713);
xnor UO_2115 (O_2115,N_19993,N_19738);
nor UO_2116 (O_2116,N_19780,N_19822);
nor UO_2117 (O_2117,N_19640,N_19658);
nand UO_2118 (O_2118,N_19909,N_19634);
and UO_2119 (O_2119,N_19820,N_19688);
and UO_2120 (O_2120,N_19931,N_19791);
and UO_2121 (O_2121,N_19787,N_19924);
nor UO_2122 (O_2122,N_19756,N_19704);
and UO_2123 (O_2123,N_19614,N_19972);
or UO_2124 (O_2124,N_19841,N_19656);
nor UO_2125 (O_2125,N_19894,N_19689);
nand UO_2126 (O_2126,N_19749,N_19637);
xor UO_2127 (O_2127,N_19956,N_19667);
or UO_2128 (O_2128,N_19819,N_19948);
or UO_2129 (O_2129,N_19605,N_19845);
xnor UO_2130 (O_2130,N_19800,N_19732);
nor UO_2131 (O_2131,N_19834,N_19710);
or UO_2132 (O_2132,N_19869,N_19809);
nand UO_2133 (O_2133,N_19756,N_19963);
nor UO_2134 (O_2134,N_19737,N_19929);
nor UO_2135 (O_2135,N_19624,N_19858);
xor UO_2136 (O_2136,N_19722,N_19644);
xnor UO_2137 (O_2137,N_19748,N_19799);
or UO_2138 (O_2138,N_19817,N_19988);
or UO_2139 (O_2139,N_19770,N_19985);
nand UO_2140 (O_2140,N_19677,N_19648);
and UO_2141 (O_2141,N_19853,N_19725);
nor UO_2142 (O_2142,N_19822,N_19700);
nor UO_2143 (O_2143,N_19999,N_19622);
and UO_2144 (O_2144,N_19716,N_19847);
and UO_2145 (O_2145,N_19766,N_19773);
xnor UO_2146 (O_2146,N_19865,N_19684);
and UO_2147 (O_2147,N_19642,N_19807);
xor UO_2148 (O_2148,N_19605,N_19997);
xor UO_2149 (O_2149,N_19938,N_19607);
or UO_2150 (O_2150,N_19641,N_19853);
xor UO_2151 (O_2151,N_19770,N_19649);
nor UO_2152 (O_2152,N_19634,N_19818);
xor UO_2153 (O_2153,N_19600,N_19943);
xnor UO_2154 (O_2154,N_19963,N_19991);
nand UO_2155 (O_2155,N_19671,N_19664);
nor UO_2156 (O_2156,N_19623,N_19828);
nand UO_2157 (O_2157,N_19927,N_19640);
nor UO_2158 (O_2158,N_19609,N_19897);
or UO_2159 (O_2159,N_19812,N_19793);
and UO_2160 (O_2160,N_19723,N_19831);
or UO_2161 (O_2161,N_19855,N_19678);
nor UO_2162 (O_2162,N_19897,N_19640);
nor UO_2163 (O_2163,N_19726,N_19954);
nand UO_2164 (O_2164,N_19617,N_19924);
or UO_2165 (O_2165,N_19782,N_19776);
or UO_2166 (O_2166,N_19780,N_19654);
nand UO_2167 (O_2167,N_19665,N_19947);
and UO_2168 (O_2168,N_19699,N_19681);
xor UO_2169 (O_2169,N_19914,N_19753);
nor UO_2170 (O_2170,N_19608,N_19990);
and UO_2171 (O_2171,N_19631,N_19844);
and UO_2172 (O_2172,N_19900,N_19935);
nand UO_2173 (O_2173,N_19639,N_19626);
or UO_2174 (O_2174,N_19823,N_19793);
or UO_2175 (O_2175,N_19600,N_19727);
and UO_2176 (O_2176,N_19949,N_19979);
and UO_2177 (O_2177,N_19796,N_19930);
xnor UO_2178 (O_2178,N_19883,N_19704);
or UO_2179 (O_2179,N_19603,N_19677);
xor UO_2180 (O_2180,N_19831,N_19868);
nand UO_2181 (O_2181,N_19889,N_19995);
nor UO_2182 (O_2182,N_19900,N_19635);
nor UO_2183 (O_2183,N_19600,N_19990);
xor UO_2184 (O_2184,N_19915,N_19750);
xor UO_2185 (O_2185,N_19793,N_19962);
xor UO_2186 (O_2186,N_19614,N_19713);
nand UO_2187 (O_2187,N_19723,N_19663);
and UO_2188 (O_2188,N_19735,N_19662);
nand UO_2189 (O_2189,N_19838,N_19651);
and UO_2190 (O_2190,N_19723,N_19851);
nand UO_2191 (O_2191,N_19750,N_19967);
nor UO_2192 (O_2192,N_19609,N_19708);
nor UO_2193 (O_2193,N_19788,N_19958);
nor UO_2194 (O_2194,N_19627,N_19935);
and UO_2195 (O_2195,N_19625,N_19963);
and UO_2196 (O_2196,N_19851,N_19782);
or UO_2197 (O_2197,N_19641,N_19956);
xnor UO_2198 (O_2198,N_19931,N_19781);
nor UO_2199 (O_2199,N_19962,N_19884);
or UO_2200 (O_2200,N_19872,N_19848);
xor UO_2201 (O_2201,N_19936,N_19798);
or UO_2202 (O_2202,N_19810,N_19690);
or UO_2203 (O_2203,N_19942,N_19619);
or UO_2204 (O_2204,N_19684,N_19683);
nor UO_2205 (O_2205,N_19673,N_19667);
or UO_2206 (O_2206,N_19739,N_19996);
nand UO_2207 (O_2207,N_19892,N_19929);
and UO_2208 (O_2208,N_19613,N_19878);
nand UO_2209 (O_2209,N_19770,N_19847);
nor UO_2210 (O_2210,N_19618,N_19603);
nor UO_2211 (O_2211,N_19840,N_19821);
and UO_2212 (O_2212,N_19690,N_19709);
nor UO_2213 (O_2213,N_19992,N_19816);
xor UO_2214 (O_2214,N_19930,N_19878);
nor UO_2215 (O_2215,N_19796,N_19861);
and UO_2216 (O_2216,N_19889,N_19808);
nand UO_2217 (O_2217,N_19715,N_19695);
xnor UO_2218 (O_2218,N_19951,N_19637);
xnor UO_2219 (O_2219,N_19852,N_19994);
or UO_2220 (O_2220,N_19825,N_19874);
and UO_2221 (O_2221,N_19736,N_19868);
and UO_2222 (O_2222,N_19636,N_19901);
xor UO_2223 (O_2223,N_19685,N_19796);
xnor UO_2224 (O_2224,N_19833,N_19901);
xnor UO_2225 (O_2225,N_19625,N_19603);
nor UO_2226 (O_2226,N_19914,N_19874);
nand UO_2227 (O_2227,N_19964,N_19898);
nor UO_2228 (O_2228,N_19882,N_19606);
and UO_2229 (O_2229,N_19723,N_19873);
xor UO_2230 (O_2230,N_19875,N_19936);
nand UO_2231 (O_2231,N_19912,N_19838);
nand UO_2232 (O_2232,N_19769,N_19878);
nor UO_2233 (O_2233,N_19928,N_19954);
or UO_2234 (O_2234,N_19893,N_19829);
nor UO_2235 (O_2235,N_19852,N_19782);
nor UO_2236 (O_2236,N_19637,N_19626);
nand UO_2237 (O_2237,N_19780,N_19658);
and UO_2238 (O_2238,N_19849,N_19920);
nor UO_2239 (O_2239,N_19974,N_19743);
nor UO_2240 (O_2240,N_19925,N_19603);
nor UO_2241 (O_2241,N_19914,N_19858);
and UO_2242 (O_2242,N_19732,N_19853);
nand UO_2243 (O_2243,N_19905,N_19609);
and UO_2244 (O_2244,N_19602,N_19720);
nor UO_2245 (O_2245,N_19651,N_19846);
nand UO_2246 (O_2246,N_19710,N_19731);
nor UO_2247 (O_2247,N_19611,N_19978);
xnor UO_2248 (O_2248,N_19915,N_19676);
or UO_2249 (O_2249,N_19923,N_19680);
or UO_2250 (O_2250,N_19921,N_19831);
nand UO_2251 (O_2251,N_19708,N_19801);
and UO_2252 (O_2252,N_19894,N_19997);
nand UO_2253 (O_2253,N_19984,N_19700);
and UO_2254 (O_2254,N_19784,N_19649);
nand UO_2255 (O_2255,N_19674,N_19776);
or UO_2256 (O_2256,N_19742,N_19724);
or UO_2257 (O_2257,N_19971,N_19610);
xor UO_2258 (O_2258,N_19940,N_19854);
and UO_2259 (O_2259,N_19992,N_19835);
nor UO_2260 (O_2260,N_19762,N_19743);
or UO_2261 (O_2261,N_19717,N_19625);
nor UO_2262 (O_2262,N_19794,N_19699);
nor UO_2263 (O_2263,N_19741,N_19603);
xor UO_2264 (O_2264,N_19927,N_19975);
nor UO_2265 (O_2265,N_19770,N_19903);
xor UO_2266 (O_2266,N_19603,N_19743);
or UO_2267 (O_2267,N_19790,N_19982);
nand UO_2268 (O_2268,N_19942,N_19662);
nor UO_2269 (O_2269,N_19990,N_19713);
nor UO_2270 (O_2270,N_19861,N_19759);
nand UO_2271 (O_2271,N_19665,N_19666);
nand UO_2272 (O_2272,N_19936,N_19953);
nand UO_2273 (O_2273,N_19601,N_19847);
nand UO_2274 (O_2274,N_19793,N_19899);
nand UO_2275 (O_2275,N_19887,N_19896);
nor UO_2276 (O_2276,N_19627,N_19779);
nor UO_2277 (O_2277,N_19622,N_19852);
nand UO_2278 (O_2278,N_19881,N_19955);
xor UO_2279 (O_2279,N_19607,N_19954);
nor UO_2280 (O_2280,N_19859,N_19873);
nor UO_2281 (O_2281,N_19933,N_19914);
nor UO_2282 (O_2282,N_19845,N_19677);
and UO_2283 (O_2283,N_19685,N_19934);
or UO_2284 (O_2284,N_19760,N_19773);
nor UO_2285 (O_2285,N_19640,N_19965);
nand UO_2286 (O_2286,N_19917,N_19956);
and UO_2287 (O_2287,N_19813,N_19634);
xor UO_2288 (O_2288,N_19718,N_19832);
and UO_2289 (O_2289,N_19844,N_19742);
xor UO_2290 (O_2290,N_19824,N_19830);
or UO_2291 (O_2291,N_19628,N_19799);
and UO_2292 (O_2292,N_19696,N_19731);
xor UO_2293 (O_2293,N_19953,N_19683);
nand UO_2294 (O_2294,N_19698,N_19667);
and UO_2295 (O_2295,N_19882,N_19685);
xnor UO_2296 (O_2296,N_19746,N_19912);
or UO_2297 (O_2297,N_19754,N_19892);
or UO_2298 (O_2298,N_19614,N_19626);
nor UO_2299 (O_2299,N_19825,N_19920);
and UO_2300 (O_2300,N_19733,N_19933);
nand UO_2301 (O_2301,N_19662,N_19866);
xor UO_2302 (O_2302,N_19784,N_19669);
xor UO_2303 (O_2303,N_19622,N_19664);
nand UO_2304 (O_2304,N_19948,N_19977);
xor UO_2305 (O_2305,N_19617,N_19815);
xor UO_2306 (O_2306,N_19904,N_19812);
nor UO_2307 (O_2307,N_19783,N_19847);
nor UO_2308 (O_2308,N_19872,N_19801);
and UO_2309 (O_2309,N_19756,N_19976);
xnor UO_2310 (O_2310,N_19914,N_19679);
xnor UO_2311 (O_2311,N_19630,N_19618);
nor UO_2312 (O_2312,N_19874,N_19806);
nor UO_2313 (O_2313,N_19897,N_19929);
nor UO_2314 (O_2314,N_19910,N_19965);
xor UO_2315 (O_2315,N_19650,N_19968);
and UO_2316 (O_2316,N_19712,N_19826);
and UO_2317 (O_2317,N_19697,N_19671);
or UO_2318 (O_2318,N_19996,N_19717);
and UO_2319 (O_2319,N_19686,N_19679);
or UO_2320 (O_2320,N_19989,N_19949);
and UO_2321 (O_2321,N_19874,N_19773);
or UO_2322 (O_2322,N_19786,N_19642);
xor UO_2323 (O_2323,N_19681,N_19943);
xor UO_2324 (O_2324,N_19895,N_19645);
and UO_2325 (O_2325,N_19713,N_19899);
or UO_2326 (O_2326,N_19870,N_19793);
and UO_2327 (O_2327,N_19781,N_19649);
nand UO_2328 (O_2328,N_19676,N_19626);
nand UO_2329 (O_2329,N_19780,N_19828);
and UO_2330 (O_2330,N_19698,N_19800);
and UO_2331 (O_2331,N_19868,N_19984);
xnor UO_2332 (O_2332,N_19839,N_19720);
or UO_2333 (O_2333,N_19635,N_19846);
xor UO_2334 (O_2334,N_19785,N_19783);
nor UO_2335 (O_2335,N_19849,N_19666);
or UO_2336 (O_2336,N_19641,N_19683);
and UO_2337 (O_2337,N_19638,N_19988);
nand UO_2338 (O_2338,N_19824,N_19654);
nand UO_2339 (O_2339,N_19944,N_19994);
or UO_2340 (O_2340,N_19693,N_19868);
nand UO_2341 (O_2341,N_19928,N_19803);
nor UO_2342 (O_2342,N_19885,N_19700);
xnor UO_2343 (O_2343,N_19970,N_19629);
nand UO_2344 (O_2344,N_19795,N_19621);
or UO_2345 (O_2345,N_19906,N_19910);
nor UO_2346 (O_2346,N_19904,N_19817);
nand UO_2347 (O_2347,N_19945,N_19811);
and UO_2348 (O_2348,N_19839,N_19693);
and UO_2349 (O_2349,N_19909,N_19971);
or UO_2350 (O_2350,N_19727,N_19990);
and UO_2351 (O_2351,N_19949,N_19865);
or UO_2352 (O_2352,N_19817,N_19606);
xnor UO_2353 (O_2353,N_19648,N_19951);
and UO_2354 (O_2354,N_19695,N_19896);
nor UO_2355 (O_2355,N_19845,N_19912);
and UO_2356 (O_2356,N_19643,N_19897);
nor UO_2357 (O_2357,N_19987,N_19629);
xnor UO_2358 (O_2358,N_19768,N_19864);
nor UO_2359 (O_2359,N_19773,N_19755);
nand UO_2360 (O_2360,N_19861,N_19731);
nand UO_2361 (O_2361,N_19664,N_19653);
and UO_2362 (O_2362,N_19772,N_19930);
xor UO_2363 (O_2363,N_19715,N_19765);
xnor UO_2364 (O_2364,N_19938,N_19866);
nand UO_2365 (O_2365,N_19827,N_19619);
nand UO_2366 (O_2366,N_19822,N_19718);
nand UO_2367 (O_2367,N_19976,N_19958);
xnor UO_2368 (O_2368,N_19838,N_19873);
or UO_2369 (O_2369,N_19925,N_19682);
xnor UO_2370 (O_2370,N_19957,N_19736);
nor UO_2371 (O_2371,N_19777,N_19754);
or UO_2372 (O_2372,N_19882,N_19966);
nand UO_2373 (O_2373,N_19955,N_19984);
and UO_2374 (O_2374,N_19827,N_19761);
xnor UO_2375 (O_2375,N_19953,N_19968);
xnor UO_2376 (O_2376,N_19639,N_19622);
nor UO_2377 (O_2377,N_19645,N_19963);
nor UO_2378 (O_2378,N_19944,N_19923);
xnor UO_2379 (O_2379,N_19806,N_19904);
xor UO_2380 (O_2380,N_19968,N_19998);
nand UO_2381 (O_2381,N_19705,N_19804);
or UO_2382 (O_2382,N_19763,N_19622);
or UO_2383 (O_2383,N_19888,N_19809);
or UO_2384 (O_2384,N_19629,N_19671);
and UO_2385 (O_2385,N_19924,N_19791);
nand UO_2386 (O_2386,N_19770,N_19797);
xnor UO_2387 (O_2387,N_19912,N_19847);
and UO_2388 (O_2388,N_19785,N_19772);
and UO_2389 (O_2389,N_19929,N_19977);
nor UO_2390 (O_2390,N_19945,N_19967);
nor UO_2391 (O_2391,N_19708,N_19745);
and UO_2392 (O_2392,N_19885,N_19696);
or UO_2393 (O_2393,N_19690,N_19768);
or UO_2394 (O_2394,N_19969,N_19980);
nand UO_2395 (O_2395,N_19811,N_19867);
nand UO_2396 (O_2396,N_19912,N_19665);
or UO_2397 (O_2397,N_19667,N_19913);
nor UO_2398 (O_2398,N_19667,N_19922);
or UO_2399 (O_2399,N_19648,N_19942);
or UO_2400 (O_2400,N_19894,N_19864);
or UO_2401 (O_2401,N_19797,N_19809);
and UO_2402 (O_2402,N_19875,N_19776);
xnor UO_2403 (O_2403,N_19863,N_19744);
nand UO_2404 (O_2404,N_19798,N_19896);
or UO_2405 (O_2405,N_19996,N_19802);
nand UO_2406 (O_2406,N_19689,N_19862);
or UO_2407 (O_2407,N_19838,N_19682);
xnor UO_2408 (O_2408,N_19874,N_19680);
nor UO_2409 (O_2409,N_19774,N_19892);
or UO_2410 (O_2410,N_19830,N_19666);
nand UO_2411 (O_2411,N_19668,N_19874);
xor UO_2412 (O_2412,N_19705,N_19696);
nor UO_2413 (O_2413,N_19710,N_19618);
and UO_2414 (O_2414,N_19668,N_19742);
nand UO_2415 (O_2415,N_19746,N_19718);
xor UO_2416 (O_2416,N_19609,N_19858);
nor UO_2417 (O_2417,N_19930,N_19692);
nor UO_2418 (O_2418,N_19638,N_19654);
nand UO_2419 (O_2419,N_19869,N_19915);
and UO_2420 (O_2420,N_19675,N_19688);
or UO_2421 (O_2421,N_19738,N_19721);
nand UO_2422 (O_2422,N_19915,N_19937);
nand UO_2423 (O_2423,N_19695,N_19955);
nor UO_2424 (O_2424,N_19623,N_19763);
nand UO_2425 (O_2425,N_19957,N_19798);
nand UO_2426 (O_2426,N_19748,N_19607);
and UO_2427 (O_2427,N_19676,N_19805);
nor UO_2428 (O_2428,N_19712,N_19842);
or UO_2429 (O_2429,N_19679,N_19604);
nor UO_2430 (O_2430,N_19737,N_19969);
xor UO_2431 (O_2431,N_19743,N_19653);
and UO_2432 (O_2432,N_19823,N_19662);
nor UO_2433 (O_2433,N_19828,N_19635);
nor UO_2434 (O_2434,N_19806,N_19759);
and UO_2435 (O_2435,N_19656,N_19875);
nor UO_2436 (O_2436,N_19648,N_19680);
and UO_2437 (O_2437,N_19977,N_19774);
nor UO_2438 (O_2438,N_19675,N_19852);
or UO_2439 (O_2439,N_19600,N_19889);
xnor UO_2440 (O_2440,N_19623,N_19973);
or UO_2441 (O_2441,N_19785,N_19899);
xnor UO_2442 (O_2442,N_19867,N_19621);
or UO_2443 (O_2443,N_19643,N_19665);
or UO_2444 (O_2444,N_19674,N_19723);
nor UO_2445 (O_2445,N_19747,N_19927);
nor UO_2446 (O_2446,N_19625,N_19828);
and UO_2447 (O_2447,N_19744,N_19964);
nor UO_2448 (O_2448,N_19639,N_19930);
nor UO_2449 (O_2449,N_19919,N_19865);
and UO_2450 (O_2450,N_19947,N_19974);
nand UO_2451 (O_2451,N_19808,N_19623);
xnor UO_2452 (O_2452,N_19814,N_19749);
xnor UO_2453 (O_2453,N_19777,N_19954);
and UO_2454 (O_2454,N_19753,N_19918);
xor UO_2455 (O_2455,N_19807,N_19665);
and UO_2456 (O_2456,N_19772,N_19633);
nor UO_2457 (O_2457,N_19863,N_19792);
nor UO_2458 (O_2458,N_19877,N_19677);
nand UO_2459 (O_2459,N_19861,N_19723);
and UO_2460 (O_2460,N_19842,N_19709);
nand UO_2461 (O_2461,N_19664,N_19608);
xor UO_2462 (O_2462,N_19996,N_19982);
and UO_2463 (O_2463,N_19776,N_19809);
nand UO_2464 (O_2464,N_19951,N_19841);
nor UO_2465 (O_2465,N_19904,N_19962);
nand UO_2466 (O_2466,N_19912,N_19871);
nor UO_2467 (O_2467,N_19781,N_19848);
or UO_2468 (O_2468,N_19672,N_19851);
or UO_2469 (O_2469,N_19873,N_19712);
xnor UO_2470 (O_2470,N_19946,N_19952);
nor UO_2471 (O_2471,N_19900,N_19729);
or UO_2472 (O_2472,N_19960,N_19769);
or UO_2473 (O_2473,N_19793,N_19685);
xor UO_2474 (O_2474,N_19762,N_19712);
nor UO_2475 (O_2475,N_19925,N_19951);
xnor UO_2476 (O_2476,N_19990,N_19873);
xnor UO_2477 (O_2477,N_19616,N_19876);
nand UO_2478 (O_2478,N_19965,N_19759);
xnor UO_2479 (O_2479,N_19767,N_19733);
and UO_2480 (O_2480,N_19635,N_19849);
xnor UO_2481 (O_2481,N_19768,N_19828);
nor UO_2482 (O_2482,N_19995,N_19988);
and UO_2483 (O_2483,N_19916,N_19601);
nor UO_2484 (O_2484,N_19659,N_19852);
and UO_2485 (O_2485,N_19746,N_19950);
or UO_2486 (O_2486,N_19959,N_19890);
or UO_2487 (O_2487,N_19629,N_19923);
xor UO_2488 (O_2488,N_19671,N_19905);
nor UO_2489 (O_2489,N_19959,N_19738);
and UO_2490 (O_2490,N_19724,N_19932);
nor UO_2491 (O_2491,N_19905,N_19824);
or UO_2492 (O_2492,N_19602,N_19903);
nand UO_2493 (O_2493,N_19737,N_19728);
and UO_2494 (O_2494,N_19799,N_19689);
or UO_2495 (O_2495,N_19726,N_19745);
or UO_2496 (O_2496,N_19960,N_19869);
xor UO_2497 (O_2497,N_19819,N_19626);
xor UO_2498 (O_2498,N_19896,N_19616);
nand UO_2499 (O_2499,N_19697,N_19898);
endmodule