module basic_2000_20000_2500_40_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1749,In_1163);
and U1 (N_1,In_1784,In_1484);
and U2 (N_2,In_610,In_932);
or U3 (N_3,In_1182,In_1577);
nor U4 (N_4,In_1499,In_1454);
nand U5 (N_5,In_1666,In_1194);
nor U6 (N_6,In_1426,In_1311);
nand U7 (N_7,In_1564,In_721);
nand U8 (N_8,In_1628,In_785);
or U9 (N_9,In_465,In_977);
and U10 (N_10,In_1330,In_965);
or U11 (N_11,In_1133,In_438);
nor U12 (N_12,In_1579,In_1334);
and U13 (N_13,In_582,In_990);
nand U14 (N_14,In_1364,In_1957);
xnor U15 (N_15,In_65,In_1595);
and U16 (N_16,In_1070,In_1800);
and U17 (N_17,In_1025,In_650);
nor U18 (N_18,In_949,In_1064);
or U19 (N_19,In_1604,In_889);
nand U20 (N_20,In_98,In_1820);
and U21 (N_21,In_894,In_353);
nand U22 (N_22,In_912,In_529);
nor U23 (N_23,In_466,In_779);
or U24 (N_24,In_809,In_420);
nor U25 (N_25,In_16,In_584);
and U26 (N_26,In_1411,In_941);
nor U27 (N_27,In_1925,In_1891);
and U28 (N_28,In_1262,In_846);
nor U29 (N_29,In_100,In_1022);
nand U30 (N_30,In_1162,In_1729);
nor U31 (N_31,In_693,In_1218);
or U32 (N_32,In_1637,In_775);
nor U33 (N_33,In_250,In_1200);
and U34 (N_34,In_504,In_601);
nand U35 (N_35,In_1605,In_503);
and U36 (N_36,In_1992,In_166);
nand U37 (N_37,In_1489,In_814);
nand U38 (N_38,In_1075,In_1221);
and U39 (N_39,In_352,In_848);
nand U40 (N_40,In_477,In_1977);
nor U41 (N_41,In_1352,In_1219);
nand U42 (N_42,In_994,In_1861);
nand U43 (N_43,In_706,In_1537);
and U44 (N_44,In_663,In_1929);
nor U45 (N_45,In_1155,In_1389);
nor U46 (N_46,In_1363,In_1517);
nand U47 (N_47,In_1348,In_1129);
or U48 (N_48,In_478,In_1545);
and U49 (N_49,In_1771,In_845);
xnor U50 (N_50,In_1934,In_1035);
nand U51 (N_51,In_1094,In_1947);
nand U52 (N_52,In_1650,In_951);
or U53 (N_53,In_871,In_1309);
or U54 (N_54,In_430,In_1447);
nor U55 (N_55,In_1049,In_1435);
nand U56 (N_56,In_1146,In_690);
nor U57 (N_57,In_1469,In_411);
and U58 (N_58,In_859,In_1900);
nor U59 (N_59,In_1067,In_718);
nor U60 (N_60,In_1935,In_699);
or U61 (N_61,In_605,In_403);
and U62 (N_62,In_426,In_696);
or U63 (N_63,In_1692,In_920);
nor U64 (N_64,In_1370,In_955);
nor U65 (N_65,In_767,In_164);
or U66 (N_66,In_1151,In_1763);
nor U67 (N_67,In_761,In_590);
and U68 (N_68,In_54,In_792);
nor U69 (N_69,In_919,In_1716);
and U70 (N_70,In_270,In_414);
nor U71 (N_71,In_437,In_1697);
and U72 (N_72,In_905,In_1889);
and U73 (N_73,In_1799,In_868);
nand U74 (N_74,In_844,In_838);
and U75 (N_75,In_433,In_799);
nor U76 (N_76,In_1552,In_874);
nand U77 (N_77,In_1117,In_408);
nand U78 (N_78,In_1758,In_1639);
nor U79 (N_79,In_1388,In_1588);
and U80 (N_80,In_483,In_1058);
nor U81 (N_81,In_1096,In_370);
or U82 (N_82,In_688,In_1984);
nor U83 (N_83,In_825,In_355);
and U84 (N_84,In_1590,In_899);
nand U85 (N_85,In_25,In_1908);
nor U86 (N_86,In_1148,In_1169);
or U87 (N_87,In_1598,In_640);
or U88 (N_88,In_1089,In_497);
nor U89 (N_89,In_542,In_307);
and U90 (N_90,In_971,In_765);
and U91 (N_91,In_762,In_985);
or U92 (N_92,In_101,In_1476);
nor U93 (N_93,In_1337,In_537);
nor U94 (N_94,In_881,In_1733);
and U95 (N_95,In_1013,In_1027);
nor U96 (N_96,In_1135,In_514);
or U97 (N_97,In_1264,In_1177);
or U98 (N_98,In_1037,In_243);
and U99 (N_99,In_872,In_1278);
or U100 (N_100,In_434,In_999);
nor U101 (N_101,In_1483,In_1786);
nand U102 (N_102,In_256,In_1712);
and U103 (N_103,In_976,In_428);
and U104 (N_104,In_1358,In_831);
nand U105 (N_105,In_1020,In_1596);
nand U106 (N_106,In_1134,In_1314);
and U107 (N_107,In_509,In_10);
or U108 (N_108,In_863,In_310);
nor U109 (N_109,In_1396,In_1005);
nor U110 (N_110,In_153,In_656);
nand U111 (N_111,In_1792,In_1016);
nand U112 (N_112,In_984,In_926);
or U113 (N_113,In_302,In_593);
nand U114 (N_114,In_987,In_1848);
and U115 (N_115,In_273,In_530);
and U116 (N_116,In_178,In_1072);
and U117 (N_117,In_1030,In_959);
nor U118 (N_118,In_1913,In_522);
or U119 (N_119,In_1896,In_416);
and U120 (N_120,In_350,In_1805);
and U121 (N_121,In_42,In_1018);
nand U122 (N_122,In_413,In_1098);
and U123 (N_123,In_1582,In_1863);
nand U124 (N_124,In_1850,In_1972);
nand U125 (N_125,In_1529,In_388);
nor U126 (N_126,In_67,In_1317);
or U127 (N_127,In_940,In_210);
xor U128 (N_128,In_1230,In_820);
nor U129 (N_129,In_764,In_760);
nand U130 (N_130,In_1462,In_40);
nor U131 (N_131,In_1463,In_1190);
or U132 (N_132,In_673,In_704);
nand U133 (N_133,In_85,In_960);
and U134 (N_134,In_1014,In_1899);
and U135 (N_135,In_563,In_1015);
and U136 (N_136,In_1099,In_644);
or U137 (N_137,In_957,In_1256);
nor U138 (N_138,In_1980,In_1157);
or U139 (N_139,In_910,In_463);
or U140 (N_140,In_1362,In_1371);
or U141 (N_141,In_1885,In_27);
nand U142 (N_142,In_251,In_1486);
or U143 (N_143,In_546,In_1390);
nand U144 (N_144,In_583,In_950);
or U145 (N_145,In_1292,In_832);
and U146 (N_146,In_1316,In_1467);
nand U147 (N_147,In_1635,In_261);
nand U148 (N_148,In_1558,In_1167);
nor U149 (N_149,In_655,In_268);
and U150 (N_150,In_769,In_404);
nand U151 (N_151,In_1281,In_1449);
nor U152 (N_152,In_389,In_1696);
or U153 (N_153,In_212,In_415);
nand U154 (N_154,In_1715,In_1803);
or U155 (N_155,In_1132,In_55);
and U156 (N_156,In_1857,In_954);
and U157 (N_157,In_1826,In_685);
or U158 (N_158,In_1207,In_1275);
and U159 (N_159,In_1926,In_1420);
or U160 (N_160,In_1719,In_1834);
nor U161 (N_161,In_649,In_1455);
or U162 (N_162,In_579,In_1199);
and U163 (N_163,In_345,In_69);
xor U164 (N_164,In_968,In_1241);
nor U165 (N_165,In_1421,In_402);
nor U166 (N_166,In_1153,In_739);
and U167 (N_167,In_109,In_1277);
nor U168 (N_168,In_710,In_1830);
nor U169 (N_169,In_1229,In_385);
nor U170 (N_170,In_1217,In_664);
or U171 (N_171,In_1888,In_1575);
and U172 (N_172,In_1503,In_519);
nand U173 (N_173,In_1626,In_1141);
nor U174 (N_174,In_259,In_1315);
or U175 (N_175,In_982,In_1559);
and U176 (N_176,In_807,In_226);
or U177 (N_177,In_666,In_1299);
or U178 (N_178,In_836,In_786);
or U179 (N_179,In_1136,In_347);
or U180 (N_180,In_177,In_66);
xnor U181 (N_181,In_933,In_1516);
nor U182 (N_182,In_60,In_216);
or U183 (N_183,In_925,In_384);
nor U184 (N_184,In_707,In_30);
and U185 (N_185,In_120,In_168);
nor U186 (N_186,In_1429,In_469);
nand U187 (N_187,In_1076,In_1448);
nand U188 (N_188,In_665,In_195);
nand U189 (N_189,In_1198,In_1078);
and U190 (N_190,In_674,In_1988);
nand U191 (N_191,In_571,In_1875);
and U192 (N_192,In_1122,In_283);
and U193 (N_193,In_200,In_1297);
or U194 (N_194,In_459,In_1368);
nand U195 (N_195,In_37,In_1050);
and U196 (N_196,In_708,In_1270);
nand U197 (N_197,In_1104,In_1498);
nand U198 (N_198,In_123,In_1986);
nor U199 (N_199,In_1663,In_1224);
or U200 (N_200,In_1865,In_12);
and U201 (N_201,In_850,In_1474);
and U202 (N_202,In_801,In_561);
nand U203 (N_203,In_417,In_1779);
nand U204 (N_204,In_1982,In_1051);
nand U205 (N_205,In_205,In_962);
nor U206 (N_206,In_643,In_154);
or U207 (N_207,In_218,In_804);
and U208 (N_208,In_810,In_1118);
and U209 (N_209,In_716,In_147);
nor U210 (N_210,In_732,In_197);
and U211 (N_211,In_486,In_111);
nand U212 (N_212,In_52,In_1731);
or U213 (N_213,In_1497,In_1251);
nand U214 (N_214,In_1748,In_1287);
or U215 (N_215,In_262,In_1647);
and U216 (N_216,In_1240,In_827);
nand U217 (N_217,In_654,In_400);
and U218 (N_218,In_1761,In_1744);
or U219 (N_219,In_1773,In_1730);
nor U220 (N_220,In_365,In_1664);
nand U221 (N_221,In_81,In_183);
and U222 (N_222,In_1958,In_170);
or U223 (N_223,In_596,In_1538);
nor U224 (N_224,In_375,In_1487);
nor U225 (N_225,In_1906,In_1107);
nor U226 (N_226,In_121,In_1062);
nand U227 (N_227,In_516,In_677);
nor U228 (N_228,In_1404,In_1086);
nor U229 (N_229,In_224,In_288);
nand U230 (N_230,In_1031,In_877);
and U231 (N_231,In_659,In_1446);
nor U232 (N_232,In_612,In_1048);
nor U233 (N_233,In_199,In_125);
and U234 (N_234,In_1717,In_684);
nand U235 (N_235,In_1927,In_1243);
and U236 (N_236,In_1933,In_713);
nand U237 (N_237,In_771,In_1427);
or U238 (N_238,In_711,In_1032);
or U239 (N_239,In_326,In_980);
and U240 (N_240,In_1678,In_983);
and U241 (N_241,In_75,In_759);
nand U242 (N_242,In_429,In_1154);
nand U243 (N_243,In_264,In_1751);
nand U244 (N_244,In_1422,In_1453);
nor U245 (N_245,In_1145,In_505);
and U246 (N_246,In_146,In_1424);
or U247 (N_247,In_1366,In_1535);
nand U248 (N_248,In_233,In_189);
nor U249 (N_249,In_1556,In_358);
or U250 (N_250,In_1894,In_485);
nand U251 (N_251,In_703,In_1480);
nand U252 (N_252,In_875,In_180);
and U253 (N_253,In_1962,In_369);
nor U254 (N_254,In_914,In_1284);
nand U255 (N_255,In_1402,In_939);
and U256 (N_256,In_1393,In_1441);
nor U257 (N_257,In_196,In_1641);
nor U258 (N_258,In_5,In_23);
or U259 (N_259,In_1653,In_336);
nor U260 (N_260,In_1568,In_45);
or U261 (N_261,In_493,In_34);
or U262 (N_262,In_869,In_322);
or U263 (N_263,In_247,In_858);
or U264 (N_264,In_1365,In_886);
nand U265 (N_265,In_637,In_298);
nor U266 (N_266,In_958,In_21);
nand U267 (N_267,In_1788,In_1767);
and U268 (N_268,In_61,In_1079);
or U269 (N_269,In_679,In_1581);
nand U270 (N_270,In_97,In_1534);
nor U271 (N_271,In_179,In_311);
or U272 (N_272,In_1391,In_126);
nand U273 (N_273,In_1354,In_1116);
xor U274 (N_274,In_1423,In_1795);
nor U275 (N_275,In_1995,In_312);
or U276 (N_276,In_1335,In_462);
or U277 (N_277,In_1540,In_1776);
nor U278 (N_278,In_723,In_712);
and U279 (N_279,In_1502,In_453);
and U280 (N_280,In_1431,In_140);
nand U281 (N_281,In_174,In_1196);
or U282 (N_282,In_1548,In_47);
nor U283 (N_283,In_1917,In_1591);
nor U284 (N_284,In_1520,In_412);
or U285 (N_285,In_172,In_290);
and U286 (N_286,In_570,In_1488);
and U287 (N_287,In_1331,In_159);
or U288 (N_288,In_1379,In_856);
and U289 (N_289,In_1818,In_938);
nor U290 (N_290,In_110,In_623);
nor U291 (N_291,In_1130,In_619);
and U292 (N_292,In_293,In_1144);
nand U293 (N_293,In_754,In_309);
nand U294 (N_294,In_1987,In_1879);
nand U295 (N_295,In_777,In_1526);
nand U296 (N_296,In_709,In_1533);
nor U297 (N_297,In_722,In_254);
and U298 (N_298,In_525,In_791);
nand U299 (N_299,In_1959,In_48);
or U300 (N_300,In_1797,In_1225);
or U301 (N_301,In_1768,In_1044);
nor U302 (N_302,In_324,In_876);
and U303 (N_303,In_953,In_1718);
nand U304 (N_304,In_1655,In_1438);
and U305 (N_305,In_692,In_1103);
nand U306 (N_306,In_1747,In_1216);
and U307 (N_307,In_1127,In_94);
nor U308 (N_308,In_552,In_734);
or U309 (N_309,In_1415,In_1560);
nor U310 (N_310,In_1739,In_630);
nor U311 (N_311,In_440,In_323);
and U312 (N_312,In_1745,In_538);
nor U313 (N_313,In_1759,In_686);
nor U314 (N_314,In_1521,In_1807);
nand U315 (N_315,In_1827,In_1753);
nor U316 (N_316,In_622,In_227);
and U317 (N_317,In_1823,In_1530);
or U318 (N_318,In_670,In_1868);
nand U319 (N_319,In_1912,In_510);
and U320 (N_320,In_209,In_1515);
or U321 (N_321,In_1464,In_1675);
nand U322 (N_322,In_1720,In_92);
or U323 (N_323,In_62,In_272);
and U324 (N_324,In_857,In_1321);
or U325 (N_325,In_986,In_1047);
or U326 (N_326,In_1110,In_1835);
nand U327 (N_327,In_946,In_22);
nor U328 (N_328,In_1054,In_329);
and U329 (N_329,In_1689,In_447);
nor U330 (N_330,In_432,In_1065);
or U331 (N_331,In_1869,In_468);
or U332 (N_332,In_824,In_318);
nand U333 (N_333,In_1833,In_1244);
and U334 (N_334,In_1838,In_1512);
or U335 (N_335,In_1849,In_1059);
nand U336 (N_336,In_1142,In_366);
and U337 (N_337,In_1380,In_1247);
nor U338 (N_338,In_1858,In_738);
or U339 (N_339,In_354,In_278);
and U340 (N_340,In_1140,In_474);
and U341 (N_341,In_800,In_1041);
and U342 (N_342,In_1332,In_569);
nor U343 (N_343,In_849,In_996);
and U344 (N_344,In_1223,In_207);
and U345 (N_345,In_1757,In_305);
or U346 (N_346,In_240,In_1623);
and U347 (N_347,In_443,In_833);
nor U348 (N_348,In_589,In_888);
nor U349 (N_349,In_851,In_1175);
or U350 (N_350,In_181,In_1152);
nand U351 (N_351,In_332,In_471);
nand U352 (N_352,In_1306,In_625);
and U353 (N_353,In_578,In_1310);
and U354 (N_354,In_488,In_1397);
nor U355 (N_355,In_1011,In_1288);
nand U356 (N_356,In_176,In_338);
nor U357 (N_357,In_1694,In_1349);
or U358 (N_358,In_1578,In_1019);
nand U359 (N_359,In_84,In_751);
nand U360 (N_360,In_1852,In_57);
nand U361 (N_361,In_1741,In_74);
and U362 (N_362,In_119,In_794);
nor U363 (N_363,In_1114,In_591);
or U364 (N_364,In_1304,In_1042);
and U365 (N_365,In_639,In_333);
nand U366 (N_366,In_134,In_1966);
nand U367 (N_367,In_1828,In_1704);
and U368 (N_368,In_1250,In_1787);
nor U369 (N_369,In_523,In_1341);
or U370 (N_370,In_544,In_1322);
nand U371 (N_371,In_361,In_1570);
or U372 (N_372,In_1989,In_1994);
nor U373 (N_373,In_339,In_1921);
nor U374 (N_374,In_1562,In_1644);
and U375 (N_375,In_1482,In_1810);
or U376 (N_376,In_1408,In_1023);
nand U377 (N_377,In_768,In_1174);
nor U378 (N_378,In_328,In_1102);
and U379 (N_379,In_911,In_1105);
and U380 (N_380,In_78,In_1300);
or U381 (N_381,In_1001,In_1907);
and U382 (N_382,In_1479,In_943);
or U383 (N_383,In_517,In_76);
xor U384 (N_384,In_1381,In_1632);
nor U385 (N_385,In_379,In_892);
nor U386 (N_386,In_864,In_1645);
nor U387 (N_387,In_1737,In_1202);
nand U388 (N_388,In_878,In_648);
nor U389 (N_389,In_286,In_918);
and U390 (N_390,In_834,In_1892);
or U391 (N_391,In_252,In_1943);
xnor U392 (N_392,In_1312,In_1772);
nand U393 (N_393,In_201,In_1629);
nor U394 (N_394,In_280,In_694);
and U395 (N_395,In_1410,In_551);
nand U396 (N_396,In_1770,In_1355);
and U397 (N_397,In_560,In_816);
or U398 (N_398,In_1361,In_1181);
and U399 (N_399,In_150,In_1923);
nand U400 (N_400,In_1793,In_1407);
or U401 (N_401,In_1043,In_1074);
or U402 (N_402,In_1339,In_1948);
and U403 (N_403,In_1658,In_808);
and U404 (N_404,In_1657,In_1481);
and U405 (N_405,In_1791,In_163);
nor U406 (N_406,In_72,In_1961);
nor U407 (N_407,In_492,In_325);
nor U408 (N_408,In_766,In_746);
nor U409 (N_409,In_1842,In_817);
nand U410 (N_410,In_620,In_129);
or U411 (N_411,In_1289,In_452);
and U412 (N_412,In_1350,In_161);
and U413 (N_413,In_217,In_904);
or U414 (N_414,In_1950,In_744);
nor U415 (N_415,In_803,In_1513);
nand U416 (N_416,In_1192,In_607);
or U417 (N_417,In_865,In_444);
nand U418 (N_418,In_952,In_1670);
nand U419 (N_419,In_50,In_1967);
or U420 (N_420,In_380,In_464);
and U421 (N_421,In_1708,In_127);
or U422 (N_422,In_839,In_1413);
or U423 (N_423,In_1711,In_854);
nor U424 (N_424,In_1640,In_1783);
or U425 (N_425,In_1097,In_1066);
nand U426 (N_426,In_1659,In_13);
nor U427 (N_427,In_235,In_145);
and U428 (N_428,In_114,In_974);
or U429 (N_429,In_211,In_1880);
and U430 (N_430,In_399,In_1269);
nor U431 (N_431,In_229,In_539);
and U432 (N_432,In_557,In_1295);
nor U433 (N_433,In_1924,In_635);
nor U434 (N_434,In_564,In_24);
nor U435 (N_435,In_879,In_1607);
nor U436 (N_436,In_1845,In_1686);
nand U437 (N_437,In_1755,In_1425);
nor U438 (N_438,In_1606,In_1746);
or U439 (N_439,In_1274,In_99);
nor U440 (N_440,In_646,In_1384);
or U441 (N_441,In_1974,In_1395);
or U442 (N_442,In_44,In_454);
or U443 (N_443,In_1963,In_1280);
and U444 (N_444,In_508,In_873);
nand U445 (N_445,In_1915,In_371);
and U446 (N_446,In_1851,In_1553);
xnor U447 (N_447,In_276,In_482);
and U448 (N_448,In_963,In_981);
nor U449 (N_449,In_1024,In_1814);
nand U450 (N_450,In_1461,In_698);
or U451 (N_451,In_435,In_1170);
nand U452 (N_452,In_774,In_822);
nand U453 (N_453,In_1360,In_1197);
or U454 (N_454,In_1353,In_691);
nor U455 (N_455,In_1672,In_1752);
nor U456 (N_456,In_966,In_930);
and U457 (N_457,In_1012,In_258);
nand U458 (N_458,In_1500,In_1674);
nand U459 (N_459,In_687,In_733);
nor U460 (N_460,In_1485,In_1608);
and U461 (N_461,In_819,In_260);
nand U462 (N_462,In_1890,In_151);
or U463 (N_463,In_1101,In_1205);
and U464 (N_464,In_317,In_1416);
or U465 (N_465,In_1296,In_342);
nand U466 (N_466,In_1855,In_1511);
and U467 (N_467,In_796,In_364);
nor U468 (N_468,In_853,In_1611);
and U469 (N_469,In_1137,In_63);
and U470 (N_470,In_1831,In_1258);
nor U471 (N_471,In_89,In_1893);
and U472 (N_472,In_80,In_135);
nand U473 (N_473,In_728,In_1166);
nand U474 (N_474,In_1220,In_909);
nor U475 (N_475,In_675,In_992);
nor U476 (N_476,In_1189,In_495);
nand U477 (N_477,In_396,In_1457);
nand U478 (N_478,In_1774,In_1226);
nor U479 (N_479,In_1093,In_1245);
and U480 (N_480,In_487,In_1620);
or U481 (N_481,In_68,In_1061);
nor U482 (N_482,In_138,In_841);
or U483 (N_483,In_1572,In_1291);
nand U484 (N_484,In_296,In_1555);
and U485 (N_485,In_829,In_1508);
and U486 (N_486,In_1298,In_167);
nor U487 (N_487,In_373,In_993);
nor U488 (N_488,In_449,In_1904);
nand U489 (N_489,In_214,In_1777);
nor U490 (N_490,In_1206,In_1239);
nand U491 (N_491,In_747,In_191);
nand U492 (N_492,In_594,In_1853);
nor U493 (N_493,In_58,In_1294);
or U494 (N_494,In_852,In_1878);
and U495 (N_495,In_297,In_1584);
and U496 (N_496,In_1460,In_1496);
nand U497 (N_497,In_1883,In_658);
nor U498 (N_498,In_128,In_294);
or U499 (N_499,In_1528,In_245);
or U500 (N_500,In_1928,N_211);
or U501 (N_501,In_1478,In_903);
nor U502 (N_502,In_1970,N_177);
nor U503 (N_503,In_1340,In_1680);
or U504 (N_504,In_567,N_118);
and U505 (N_505,In_705,In_1053);
nand U506 (N_506,In_1532,N_362);
nand U507 (N_507,In_1087,In_1633);
nor U508 (N_508,N_38,In_1039);
nand U509 (N_509,In_609,N_329);
or U510 (N_510,In_559,N_461);
or U511 (N_511,N_430,In_395);
or U512 (N_512,In_1060,In_653);
and U513 (N_513,N_376,In_587);
nor U514 (N_514,In_271,In_660);
and U515 (N_515,In_1418,In_1045);
and U516 (N_516,In_1616,In_1125);
and U517 (N_517,In_376,In_363);
or U518 (N_518,In_1318,N_335);
or U519 (N_519,In_882,In_173);
or U520 (N_520,In_165,N_364);
and U521 (N_521,In_964,N_139);
nand U522 (N_522,N_276,In_652);
or U523 (N_523,In_840,N_97);
or U524 (N_524,N_46,In_1610);
and U525 (N_525,In_742,In_533);
nand U526 (N_526,In_945,In_1592);
nor U527 (N_527,In_575,In_202);
nor U528 (N_528,N_57,In_1385);
or U529 (N_529,In_418,In_753);
and U530 (N_530,In_1652,In_287);
and U531 (N_531,N_209,In_467);
or U532 (N_532,N_389,In_662);
and U533 (N_533,N_263,In_1522);
or U534 (N_534,In_1910,N_166);
and U535 (N_535,In_1527,In_618);
and U536 (N_536,N_226,N_313);
and U537 (N_537,In_26,In_228);
and U538 (N_538,In_1939,In_1510);
nand U539 (N_539,N_333,In_292);
and U540 (N_540,N_18,N_233);
nor U541 (N_541,N_179,In_1124);
or U542 (N_542,In_1756,N_230);
or U543 (N_543,In_1983,In_1029);
or U544 (N_544,In_1369,N_398);
and U545 (N_545,N_149,In_6);
and U546 (N_546,In_1108,In_1952);
or U547 (N_547,N_167,In_772);
or U548 (N_548,In_1,In_1956);
nand U549 (N_549,In_931,In_18);
and U550 (N_550,In_924,In_1622);
or U551 (N_551,In_1518,N_271);
or U552 (N_552,In_967,In_1618);
nand U553 (N_553,In_611,In_634);
or U554 (N_554,N_251,In_1812);
nand U555 (N_555,N_62,In_1405);
nor U556 (N_556,N_221,N_168);
nand U557 (N_557,N_184,N_21);
nor U558 (N_558,In_548,In_1524);
and U559 (N_559,In_1235,In_90);
nor U560 (N_560,N_463,N_66);
or U561 (N_561,In_883,In_599);
and U562 (N_562,N_208,N_172);
or U563 (N_563,In_1073,N_93);
and U564 (N_564,In_1392,In_1257);
or U565 (N_565,In_344,In_1614);
and U566 (N_566,In_855,N_387);
or U567 (N_567,In_1343,In_531);
nand U568 (N_568,In_1228,N_444);
nor U569 (N_569,In_798,In_900);
nor U570 (N_570,In_203,N_484);
nand U571 (N_571,In_1874,In_1801);
nor U572 (N_572,N_156,In_835);
or U573 (N_573,In_1612,In_53);
xor U574 (N_574,In_249,N_296);
nor U575 (N_575,N_289,In_187);
nor U576 (N_576,In_1844,In_1769);
and U577 (N_577,In_104,In_93);
nand U578 (N_578,In_1550,In_921);
nor U579 (N_579,In_720,N_386);
nand U580 (N_580,N_29,In_614);
and U581 (N_581,In_1063,N_352);
or U582 (N_582,N_310,N_187);
and U583 (N_583,In_1846,In_223);
and U584 (N_584,N_191,In_1525);
nor U585 (N_585,N_228,N_426);
nand U586 (N_586,In_1433,N_185);
and U587 (N_587,N_348,In_1176);
nor U588 (N_588,In_436,In_1147);
nor U589 (N_589,In_301,N_303);
nand U590 (N_590,In_1473,In_313);
and U591 (N_591,In_185,N_35);
nand U592 (N_592,N_419,N_110);
or U593 (N_593,N_402,In_1386);
nand U594 (N_594,In_1293,In_729);
nor U595 (N_595,In_935,In_1960);
and U596 (N_596,In_1914,In_441);
nand U597 (N_597,In_96,In_162);
or U598 (N_598,N_286,In_1740);
and U599 (N_599,In_1685,In_885);
nand U600 (N_600,In_1290,N_8);
or U601 (N_601,N_493,In_1036);
nand U602 (N_602,In_944,In_1208);
nand U603 (N_603,In_1714,In_554);
nor U604 (N_604,In_1877,N_240);
or U605 (N_605,In_1750,In_337);
or U606 (N_606,In_248,In_295);
or U607 (N_607,In_1662,In_1843);
or U608 (N_608,N_297,N_64);
or U609 (N_609,N_272,In_1897);
or U610 (N_610,In_1651,In_1266);
nand U611 (N_611,In_107,N_258);
or U612 (N_612,N_195,N_411);
nor U613 (N_613,N_197,In_386);
nand U614 (N_614,In_1862,In_645);
and U615 (N_615,In_1253,N_366);
nand U616 (N_616,In_499,N_302);
nor U617 (N_617,N_314,In_602);
nand U618 (N_618,In_1702,In_489);
and U619 (N_619,In_749,In_736);
nand U620 (N_620,N_481,In_577);
and U621 (N_621,In_520,N_359);
nand U622 (N_622,N_395,N_182);
nor U623 (N_623,N_44,In_927);
or U624 (N_624,In_1683,In_368);
or U625 (N_625,In_1286,N_227);
or U626 (N_626,In_263,In_1249);
nand U627 (N_627,N_356,In_39);
or U628 (N_628,In_242,In_1519);
and U629 (N_629,In_1412,N_455);
nand U630 (N_630,In_88,In_1656);
nor U631 (N_631,In_35,In_1399);
and U632 (N_632,In_232,In_535);
nand U633 (N_633,In_473,In_1706);
nor U634 (N_634,In_1809,In_215);
or U635 (N_635,In_1542,N_305);
nand U636 (N_636,N_238,In_802);
and U637 (N_637,In_281,N_229);
nand U638 (N_638,N_332,In_528);
or U639 (N_639,In_241,In_1285);
or U640 (N_640,In_1100,N_341);
nor U641 (N_641,In_756,N_246);
and U642 (N_642,N_100,N_384);
nand U643 (N_643,In_1593,N_262);
nor U644 (N_644,In_431,In_422);
or U645 (N_645,N_418,In_545);
xor U646 (N_646,In_647,In_11);
and U647 (N_647,N_406,In_1585);
nor U648 (N_648,In_923,In_512);
nand U649 (N_649,In_41,N_33);
nand U650 (N_650,In_1255,N_299);
and U651 (N_651,In_1403,N_54);
nand U652 (N_652,N_171,N_214);
or U653 (N_653,N_365,In_1973);
and U654 (N_654,In_1673,In_31);
and U655 (N_655,In_1942,In_1836);
nor U656 (N_656,N_193,In_755);
and U657 (N_657,N_235,In_1840);
and U658 (N_658,In_661,N_123);
nand U659 (N_659,N_317,In_1186);
and U660 (N_660,N_290,In_613);
and U661 (N_661,N_279,In_540);
nor U662 (N_662,N_468,In_1008);
nand U663 (N_663,In_142,In_1667);
nor U664 (N_664,In_550,N_42);
or U665 (N_665,In_1459,N_466);
or U666 (N_666,In_1778,N_43);
and U667 (N_667,N_351,In_1684);
nand U668 (N_668,In_847,In_870);
or U669 (N_669,N_327,In_277);
or U670 (N_670,N_83,In_1038);
nand U671 (N_671,N_392,In_1794);
or U672 (N_672,In_221,N_321);
nand U673 (N_673,In_390,In_942);
and U674 (N_674,In_770,N_451);
and U675 (N_675,In_143,In_702);
and U676 (N_676,N_27,In_175);
nor U677 (N_677,N_436,In_424);
nand U678 (N_678,N_127,In_1985);
nor U679 (N_679,In_1374,N_134);
or U680 (N_680,In_451,N_422);
and U681 (N_681,In_616,N_486);
nor U682 (N_682,N_124,N_316);
nand U683 (N_683,In_319,In_1382);
nand U684 (N_684,In_1886,N_180);
or U685 (N_685,In_1876,In_568);
and U686 (N_686,In_1922,In_105);
and U687 (N_687,In_157,N_108);
nor U688 (N_688,In_239,In_1785);
nor U689 (N_689,N_116,In_1938);
nor U690 (N_690,N_89,In_526);
nand U691 (N_691,In_1507,N_76);
and U692 (N_692,In_382,In_1839);
or U693 (N_693,In_657,In_978);
nor U694 (N_694,In_1726,N_433);
and U695 (N_695,N_45,N_391);
or U696 (N_696,N_261,In_1601);
and U697 (N_697,N_70,In_1346);
nor U698 (N_698,N_388,In_419);
nor U699 (N_699,In_308,In_275);
nand U700 (N_700,N_155,In_86);
nor U701 (N_701,In_182,In_576);
or U702 (N_702,In_51,In_511);
nand U703 (N_703,In_502,N_370);
and U704 (N_704,In_1267,In_122);
and U705 (N_705,N_479,In_1302);
nor U706 (N_706,In_837,In_1808);
nand U707 (N_707,In_676,N_142);
nor U708 (N_708,In_193,N_339);
and U709 (N_709,In_124,In_1009);
or U710 (N_710,N_408,In_1617);
and U711 (N_711,In_401,In_1969);
nor U712 (N_712,In_4,In_1789);
nor U713 (N_713,N_274,In_830);
and U714 (N_714,N_125,In_1856);
nor U715 (N_715,N_5,In_7);
and U716 (N_716,N_53,N_255);
and U717 (N_717,In_1955,N_98);
nand U718 (N_718,In_1319,In_1871);
nor U719 (N_719,N_417,In_1895);
and U720 (N_720,In_1326,In_341);
nand U721 (N_721,In_1760,In_1728);
and U722 (N_722,N_450,N_128);
xnor U723 (N_723,In_1901,N_37);
or U724 (N_724,In_82,In_669);
or U725 (N_725,N_114,N_80);
nand U726 (N_726,In_719,In_1214);
nor U727 (N_727,In_1627,In_184);
nor U728 (N_728,In_1941,In_1599);
nor U729 (N_729,In_351,In_566);
nand U730 (N_730,In_773,N_148);
nor U731 (N_731,In_1121,N_39);
xnor U732 (N_732,N_17,In_71);
nor U733 (N_733,In_600,N_181);
or U734 (N_734,In_1069,N_371);
nand U735 (N_735,In_667,N_41);
or U736 (N_736,In_1383,N_318);
or U737 (N_737,N_361,N_264);
and U738 (N_738,In_956,N_278);
or U739 (N_739,In_1010,N_212);
or U740 (N_740,In_1347,In_1991);
and U741 (N_741,N_87,In_274);
and U742 (N_742,In_700,In_1695);
nor U743 (N_743,N_69,In_1642);
and U744 (N_744,In_1320,In_636);
nand U745 (N_745,In_1993,In_1547);
nor U746 (N_746,N_122,In_1514);
or U747 (N_747,In_884,N_320);
nor U748 (N_748,In_748,N_96);
and U749 (N_749,N_399,N_11);
nand U750 (N_750,In_1734,In_1238);
and U751 (N_751,In_1359,In_997);
nor U752 (N_752,N_9,N_56);
nor U753 (N_753,In_998,In_752);
nor U754 (N_754,In_1283,In_1998);
nor U755 (N_755,In_204,N_369);
nor U756 (N_756,In_378,In_1603);
nand U757 (N_757,In_265,In_1325);
xnor U758 (N_758,N_103,In_1710);
and U759 (N_759,In_314,N_225);
nor U760 (N_760,In_137,N_470);
nor U761 (N_761,In_778,In_1766);
nand U762 (N_762,In_797,N_298);
and U763 (N_763,N_315,In_304);
nor U764 (N_764,In_108,In_334);
and U765 (N_765,In_893,In_574);
nor U766 (N_766,In_1077,In_1236);
nand U767 (N_767,In_668,N_248);
nor U768 (N_768,In_1246,N_253);
nand U769 (N_769,In_190,N_311);
or U770 (N_770,N_244,In_1345);
or U771 (N_771,N_173,In_1092);
nor U772 (N_772,N_322,N_480);
nand U773 (N_773,In_1273,In_1705);
and U774 (N_774,In_763,In_787);
nand U775 (N_775,In_1456,In_117);
nand U776 (N_776,In_1439,In_860);
nand U777 (N_777,N_48,In_890);
nor U778 (N_778,In_1468,In_357);
nor U779 (N_779,In_405,In_206);
and U780 (N_780,In_472,In_572);
nor U781 (N_781,In_367,N_407);
and U782 (N_782,N_377,N_325);
nand U783 (N_783,N_219,N_355);
xor U784 (N_784,In_1301,In_547);
and U785 (N_785,In_320,N_107);
xor U786 (N_786,In_1040,In_1796);
and U787 (N_787,In_1090,In_1713);
nand U788 (N_788,N_55,N_88);
nand U789 (N_789,N_165,N_354);
or U790 (N_790,In_1829,In_532);
nor U791 (N_791,In_491,In_356);
or U792 (N_792,In_383,In_158);
and U793 (N_793,In_1732,In_1679);
nor U794 (N_794,In_284,In_1549);
or U795 (N_795,In_812,N_75);
nor U796 (N_796,In_234,In_149);
or U797 (N_797,In_1775,In_255);
nand U798 (N_798,N_133,In_682);
xor U799 (N_799,In_898,N_259);
and U800 (N_800,N_342,In_442);
and U801 (N_801,N_222,In_112);
and U802 (N_802,In_1551,In_1884);
and U803 (N_803,N_154,N_36);
nor U804 (N_804,In_1434,In_1115);
or U805 (N_805,N_192,N_79);
nand U806 (N_806,N_82,In_1028);
and U807 (N_807,N_363,N_266);
or U808 (N_808,In_1372,In_651);
or U809 (N_809,In_20,In_1944);
nor U810 (N_810,In_562,In_597);
nor U811 (N_811,In_1495,N_283);
xor U812 (N_812,In_15,In_592);
nand U813 (N_813,In_1798,N_454);
and U814 (N_814,N_346,In_1721);
and U815 (N_815,N_414,In_188);
nor U816 (N_816,In_1209,In_222);
or U817 (N_817,In_811,In_1400);
and U818 (N_818,In_1139,In_1722);
nand U819 (N_819,N_23,In_1313);
and U820 (N_820,In_257,In_1213);
and U821 (N_821,In_1375,In_1417);
nand U822 (N_822,N_291,N_74);
nand U823 (N_823,N_220,In_335);
or U824 (N_824,N_441,N_427);
or U825 (N_825,In_1440,In_750);
or U826 (N_826,In_1997,N_92);
xor U827 (N_827,In_103,N_292);
and U828 (N_828,In_783,N_51);
or U829 (N_829,In_1817,N_4);
or U830 (N_830,N_52,In_169);
and U831 (N_831,In_1164,In_327);
and U832 (N_832,In_500,In_1261);
nor U833 (N_833,In_758,In_343);
and U834 (N_834,In_1180,In_1187);
nor U835 (N_835,In_1376,In_726);
nand U836 (N_836,In_741,In_1837);
xnor U837 (N_837,In_1887,In_237);
and U838 (N_838,N_488,In_1701);
or U839 (N_839,N_94,In_289);
and U840 (N_840,In_2,N_428);
and U841 (N_841,In_1477,N_336);
nand U842 (N_842,In_1723,N_343);
nor U843 (N_843,In_1567,In_1665);
nor U844 (N_844,In_1574,N_404);
or U845 (N_845,N_378,In_1565);
or U846 (N_846,In_1272,N_216);
and U847 (N_847,N_494,In_1693);
nand U848 (N_848,In_1212,In_410);
nor U849 (N_849,N_326,In_1242);
and U850 (N_850,In_1327,In_1007);
and U851 (N_851,In_790,N_338);
nor U852 (N_852,N_19,In_1866);
or U853 (N_853,In_1159,In_1017);
nor U854 (N_854,In_1265,In_19);
and U855 (N_855,In_1654,In_1873);
and U856 (N_856,In_1859,In_1539);
and U857 (N_857,In_225,N_353);
nor U858 (N_858,In_806,In_156);
and U859 (N_859,In_1764,In_781);
and U860 (N_860,N_456,In_1832);
and U861 (N_861,In_14,In_1172);
or U862 (N_862,N_105,In_553);
nor U863 (N_863,In_632,N_163);
and U864 (N_864,In_1902,In_937);
or U865 (N_865,In_1687,N_50);
nor U866 (N_866,In_1493,In_116);
and U867 (N_867,In_244,In_501);
nor U868 (N_868,In_236,In_282);
nand U869 (N_869,In_972,N_217);
or U870 (N_870,N_476,In_1765);
or U871 (N_871,N_337,In_1700);
nand U872 (N_872,In_717,In_1046);
and U873 (N_873,In_36,N_449);
and U874 (N_874,In_1954,N_6);
nor U875 (N_875,In_77,In_1357);
and U876 (N_876,N_424,N_143);
nor U877 (N_877,In_1782,In_1536);
and U878 (N_878,In_1636,N_199);
or U879 (N_879,N_295,N_3);
and U880 (N_880,In_1119,In_1002);
or U881 (N_881,N_475,In_1905);
nand U882 (N_882,In_907,In_866);
and U883 (N_883,In_291,N_7);
nor U884 (N_884,In_118,In_1597);
nand U885 (N_885,In_1113,In_1882);
or U886 (N_886,In_1080,N_0);
and U887 (N_887,N_260,In_446);
nor U888 (N_888,In_1123,In_1609);
or U889 (N_889,In_1490,In_303);
nor U890 (N_890,In_1143,N_194);
nor U891 (N_891,N_151,In_543);
nor U892 (N_892,In_697,In_1543);
and U893 (N_893,In_928,In_59);
or U894 (N_894,In_1649,In_633);
nor U895 (N_895,In_1949,In_346);
or U896 (N_896,In_1813,N_270);
nor U897 (N_897,In_1648,In_678);
or U898 (N_898,In_1978,In_595);
nand U899 (N_899,In_1619,In_340);
and U900 (N_900,In_672,N_446);
nor U901 (N_901,In_1630,N_497);
or U902 (N_902,In_1589,In_795);
nor U903 (N_903,In_1237,In_1822);
nand U904 (N_904,N_495,In_615);
nor U905 (N_905,In_1401,N_301);
or U906 (N_906,In_934,N_437);
or U907 (N_907,In_861,In_475);
nand U908 (N_908,In_299,In_1587);
and U909 (N_909,In_624,In_524);
or U910 (N_910,In_715,In_1178);
nand U911 (N_911,In_476,In_479);
nand U912 (N_912,N_249,In_1055);
or U913 (N_913,N_256,N_429);
nand U914 (N_914,In_541,In_598);
or U915 (N_915,In_1328,In_1308);
nand U916 (N_916,In_1971,In_1248);
nand U917 (N_917,In_460,In_1802);
nor U918 (N_918,N_65,In_1323);
or U919 (N_919,In_208,N_385);
nor U920 (N_920,In_1387,In_1436);
nand U921 (N_921,N_294,In_973);
xor U922 (N_922,In_782,In_113);
or U923 (N_923,N_90,In_397);
or U924 (N_924,In_1344,In_776);
nand U925 (N_925,In_1168,N_442);
nand U926 (N_926,In_780,In_316);
nor U927 (N_927,N_170,In_891);
nand U928 (N_928,N_323,In_1471);
nor U929 (N_929,In_1688,In_1682);
or U930 (N_930,In_490,In_1305);
nor U931 (N_931,In_507,In_409);
nor U932 (N_932,In_991,In_1909);
or U933 (N_933,In_1450,N_120);
nor U934 (N_934,N_443,In_1409);
and U935 (N_935,N_492,N_25);
nand U936 (N_936,N_91,In_1563);
nor U937 (N_937,N_59,In_33);
or U938 (N_938,In_1600,In_1573);
nor U939 (N_939,N_206,In_1088);
nand U940 (N_940,In_349,N_203);
and U941 (N_941,N_241,N_400);
and U942 (N_942,In_269,In_549);
nor U943 (N_943,N_113,In_1561);
nand U944 (N_944,In_1624,In_1081);
or U945 (N_945,In_427,In_246);
and U946 (N_946,In_1979,In_391);
nand U947 (N_947,N_28,In_701);
and U948 (N_948,In_1106,In_518);
and U949 (N_949,In_456,In_1259);
xor U950 (N_950,N_401,In_230);
nand U951 (N_951,In_91,N_257);
nor U952 (N_952,In_1437,In_603);
nand U953 (N_953,In_1068,In_527);
nor U954 (N_954,In_29,In_73);
nor U955 (N_955,N_447,In_1095);
and U956 (N_956,N_132,In_1338);
and U957 (N_957,In_1506,N_73);
nand U958 (N_958,In_1373,In_1149);
or U959 (N_959,In_1804,In_1034);
or U960 (N_960,In_1638,N_358);
and U961 (N_961,In_1819,In_266);
and U962 (N_962,N_111,N_381);
nand U963 (N_963,N_237,In_1580);
and U964 (N_964,N_77,In_1201);
nand U965 (N_965,N_405,N_138);
nor U966 (N_966,In_1351,In_1211);
nor U967 (N_967,In_1445,N_334);
xor U968 (N_968,In_1492,N_1);
or U969 (N_969,In_1505,N_13);
or U970 (N_970,In_484,N_347);
and U971 (N_971,N_324,N_198);
and U972 (N_972,In_638,In_481);
nor U973 (N_973,N_478,In_1193);
nand U974 (N_974,In_49,In_1583);
or U975 (N_975,N_499,N_491);
nand U976 (N_976,N_129,N_16);
and U977 (N_977,In_580,N_117);
or U978 (N_978,In_393,N_269);
nor U979 (N_979,In_1919,N_421);
nand U980 (N_980,In_695,N_445);
or U981 (N_981,In_1470,N_141);
nand U982 (N_982,N_410,In_805);
and U983 (N_983,In_1727,N_174);
nand U984 (N_984,In_948,N_425);
and U985 (N_985,N_458,In_1691);
nor U986 (N_986,N_130,In_823);
nor U987 (N_987,N_496,In_913);
and U988 (N_988,In_1523,N_288);
and U989 (N_989,N_498,N_15);
nor U990 (N_990,N_137,N_68);
nor U991 (N_991,In_1676,N_146);
nor U992 (N_992,In_1699,In_961);
or U993 (N_993,In_1936,N_413);
nor U994 (N_994,In_1419,In_586);
nor U995 (N_995,N_350,In_1033);
or U996 (N_996,In_1307,In_606);
nand U997 (N_997,In_1613,N_368);
nand U998 (N_998,In_1004,N_306);
or U999 (N_999,N_345,In_455);
and U1000 (N_1000,N_994,N_541);
nand U1001 (N_1001,N_714,In_887);
and U1002 (N_1002,In_1222,N_593);
nand U1003 (N_1003,In_392,N_724);
nor U1004 (N_1004,In_381,N_189);
nor U1005 (N_1005,N_833,In_642);
and U1006 (N_1006,In_285,N_894);
nand U1007 (N_1007,N_504,N_594);
nor U1008 (N_1008,N_692,N_511);
nor U1009 (N_1009,In_714,N_659);
nand U1010 (N_1010,In_1000,In_498);
or U1011 (N_1011,In_360,N_853);
or U1012 (N_1012,N_610,N_112);
or U1013 (N_1013,N_554,N_438);
and U1014 (N_1014,N_243,N_390);
or U1015 (N_1015,N_462,In_1191);
nor U1016 (N_1016,N_285,In_867);
and U1017 (N_1017,N_556,N_612);
and U1018 (N_1018,N_690,N_686);
nand U1019 (N_1019,N_749,N_810);
nand U1020 (N_1020,N_106,In_916);
and U1021 (N_1021,N_795,In_1150);
and U1022 (N_1022,In_213,N_995);
or U1023 (N_1023,N_975,N_627);
or U1024 (N_1024,In_689,In_1491);
nand U1025 (N_1025,In_534,N_720);
nand U1026 (N_1026,N_540,In_1160);
or U1027 (N_1027,N_921,N_768);
or U1028 (N_1028,In_445,N_697);
or U1029 (N_1029,In_1084,N_619);
nor U1030 (N_1030,In_1981,N_675);
nand U1031 (N_1031,N_14,N_489);
nor U1032 (N_1032,N_762,In_1743);
nand U1033 (N_1033,N_763,N_704);
nand U1034 (N_1034,In_901,N_160);
nand U1035 (N_1035,N_277,N_534);
or U1036 (N_1036,N_988,N_634);
nand U1037 (N_1037,In_1171,N_755);
nor U1038 (N_1038,N_867,In_1932);
or U1039 (N_1039,N_706,In_377);
or U1040 (N_1040,N_819,N_699);
nand U1041 (N_1041,N_662,N_245);
nor U1042 (N_1042,N_874,In_1762);
or U1043 (N_1043,N_903,N_696);
nand U1044 (N_1044,N_157,N_655);
nand U1045 (N_1045,In_1378,N_787);
nand U1046 (N_1046,N_863,In_194);
or U1047 (N_1047,In_131,N_764);
nand U1048 (N_1048,In_1571,In_1188);
nor U1049 (N_1049,In_826,N_917);
nor U1050 (N_1050,N_613,In_450);
and U1051 (N_1051,N_420,In_1999);
nor U1052 (N_1052,N_962,N_772);
nor U1053 (N_1053,N_681,N_983);
nand U1054 (N_1054,In_1472,N_207);
nand U1055 (N_1055,N_252,N_58);
nand U1056 (N_1056,In_731,N_563);
and U1057 (N_1057,In_0,In_279);
nor U1058 (N_1058,N_667,In_979);
and U1059 (N_1059,N_929,N_570);
nor U1060 (N_1060,N_20,In_219);
or U1061 (N_1061,N_809,In_132);
and U1062 (N_1062,N_601,In_1725);
nand U1063 (N_1063,In_1398,N_818);
and U1064 (N_1064,N_785,In_1681);
or U1065 (N_1065,N_175,In_1203);
nor U1066 (N_1066,N_218,In_83);
nand U1067 (N_1067,In_1990,N_561);
and U1068 (N_1068,N_708,N_394);
nand U1069 (N_1069,In_588,N_828);
nand U1070 (N_1070,In_1052,N_713);
or U1071 (N_1071,In_1085,In_555);
and U1072 (N_1072,In_267,N_615);
and U1073 (N_1073,In_1367,In_406);
and U1074 (N_1074,N_946,N_799);
nand U1075 (N_1075,In_573,N_911);
nor U1076 (N_1076,In_1964,In_1195);
or U1077 (N_1077,N_604,N_607);
xnor U1078 (N_1078,N_707,N_415);
nand U1079 (N_1079,N_529,N_866);
nor U1080 (N_1080,N_614,N_982);
nand U1081 (N_1081,N_596,N_473);
or U1082 (N_1082,N_553,N_934);
nor U1083 (N_1083,In_1509,In_735);
and U1084 (N_1084,N_144,N_161);
nand U1085 (N_1085,N_611,N_367);
and U1086 (N_1086,N_736,N_521);
or U1087 (N_1087,N_744,N_701);
or U1088 (N_1088,In_1021,N_247);
nand U1089 (N_1089,In_1825,N_660);
or U1090 (N_1090,In_1996,In_818);
nor U1091 (N_1091,N_448,N_293);
nor U1092 (N_1092,N_663,In_1254);
and U1093 (N_1093,N_849,N_176);
nand U1094 (N_1094,In_1501,N_517);
nand U1095 (N_1095,N_357,In_1975);
nor U1096 (N_1096,N_726,N_633);
and U1097 (N_1097,N_985,N_152);
nor U1098 (N_1098,N_769,N_746);
nand U1099 (N_1099,N_865,N_992);
nor U1100 (N_1100,N_330,N_582);
or U1101 (N_1101,N_885,In_1576);
and U1102 (N_1102,N_782,In_1356);
nand U1103 (N_1103,N_586,N_647);
nor U1104 (N_1104,N_501,In_1931);
nand U1105 (N_1105,N_213,N_200);
and U1106 (N_1106,N_568,N_850);
nand U1107 (N_1107,N_268,N_609);
and U1108 (N_1108,N_431,In_975);
and U1109 (N_1109,N_86,N_731);
nor U1110 (N_1110,N_694,N_215);
nor U1111 (N_1111,N_914,N_464);
or U1112 (N_1112,N_505,In_457);
or U1113 (N_1113,In_1634,In_136);
or U1114 (N_1114,In_38,N_642);
nor U1115 (N_1115,N_580,N_904);
xor U1116 (N_1116,N_34,N_453);
or U1117 (N_1117,N_432,In_46);
or U1118 (N_1118,N_957,In_740);
nor U1119 (N_1119,N_602,In_1210);
nand U1120 (N_1120,In_32,N_862);
nand U1121 (N_1121,In_439,N_526);
and U1122 (N_1122,N_925,In_1279);
or U1123 (N_1123,N_753,N_820);
nor U1124 (N_1124,N_516,In_1442);
and U1125 (N_1125,N_656,N_490);
nor U1126 (N_1126,N_703,N_300);
and U1127 (N_1127,N_668,In_1475);
nor U1128 (N_1128,In_1282,N_472);
nor U1129 (N_1129,N_331,In_198);
nand U1130 (N_1130,N_523,N_485);
or U1131 (N_1131,In_922,N_966);
nand U1132 (N_1132,In_1444,In_880);
nor U1133 (N_1133,N_913,In_813);
nor U1134 (N_1134,N_508,N_588);
nor U1135 (N_1135,N_883,N_629);
nor U1136 (N_1136,N_571,In_585);
or U1137 (N_1137,N_765,In_1126);
and U1138 (N_1138,N_936,N_700);
nor U1139 (N_1139,In_902,In_458);
or U1140 (N_1140,In_1690,N_807);
nor U1141 (N_1141,N_728,N_698);
or U1142 (N_1142,N_932,N_986);
and U1143 (N_1143,N_635,N_81);
and U1144 (N_1144,N_282,N_49);
or U1145 (N_1145,N_528,N_319);
or U1146 (N_1146,N_826,N_680);
or U1147 (N_1147,N_971,In_1452);
or U1148 (N_1148,N_560,N_628);
and U1149 (N_1149,N_899,N_636);
and U1150 (N_1150,In_1263,In_915);
or U1151 (N_1151,N_671,In_506);
or U1152 (N_1152,N_375,N_757);
and U1153 (N_1153,In_862,N_630);
or U1154 (N_1154,In_788,N_789);
nand U1155 (N_1155,In_1602,In_513);
nor U1156 (N_1156,N_716,N_895);
nand U1157 (N_1157,N_581,N_920);
nand U1158 (N_1158,N_823,In_1303);
and U1159 (N_1159,N_836,N_889);
nand U1160 (N_1160,N_831,In_680);
xor U1161 (N_1161,N_374,N_578);
nor U1162 (N_1162,N_931,In_1621);
and U1163 (N_1163,N_881,N_952);
nand U1164 (N_1164,N_597,N_340);
nand U1165 (N_1165,In_1231,N_705);
and U1166 (N_1166,In_1707,N_10);
nor U1167 (N_1167,N_978,N_649);
nand U1168 (N_1168,N_915,In_743);
nor U1169 (N_1169,N_891,N_482);
nand U1170 (N_1170,In_1668,In_1466);
or U1171 (N_1171,N_811,N_848);
or U1172 (N_1172,N_880,N_31);
nand U1173 (N_1173,N_543,N_725);
nand U1174 (N_1174,N_435,In_1860);
nand U1175 (N_1175,In_629,N_743);
nor U1176 (N_1176,In_1677,In_56);
or U1177 (N_1177,N_732,N_178);
and U1178 (N_1178,N_632,N_572);
or U1179 (N_1179,In_3,N_555);
nor U1180 (N_1180,N_61,In_1268);
or U1181 (N_1181,N_188,N_839);
nor U1182 (N_1182,N_758,N_774);
and U1183 (N_1183,N_382,In_106);
and U1184 (N_1184,N_841,N_109);
nand U1185 (N_1185,N_205,N_679);
or U1186 (N_1186,N_201,In_398);
nor U1187 (N_1187,N_905,In_1083);
and U1188 (N_1188,In_133,N_723);
and U1189 (N_1189,N_439,N_864);
nor U1190 (N_1190,N_509,N_530);
and U1191 (N_1191,In_1930,N_734);
or U1192 (N_1192,N_40,In_1671);
nand U1193 (N_1193,N_416,In_1260);
nor U1194 (N_1194,In_641,N_842);
nor U1195 (N_1195,N_549,N_779);
nand U1196 (N_1196,In_1179,N_372);
or U1197 (N_1197,In_480,N_676);
nand U1198 (N_1198,N_965,In_1951);
nor U1199 (N_1199,N_652,N_532);
nor U1200 (N_1200,In_1494,N_741);
and U1201 (N_1201,N_875,N_608);
and U1202 (N_1202,N_474,N_797);
nand U1203 (N_1203,N_162,In_1394);
nand U1204 (N_1204,In_1546,N_791);
and U1205 (N_1205,N_231,In_1204);
or U1206 (N_1206,In_628,N_585);
or U1207 (N_1207,N_858,N_623);
and U1208 (N_1208,In_1158,In_1569);
nand U1209 (N_1209,N_670,In_95);
and U1210 (N_1210,N_890,In_995);
and U1211 (N_1211,N_718,In_1465);
nand U1212 (N_1212,N_527,In_186);
or U1213 (N_1213,N_645,In_1735);
or U1214 (N_1214,N_773,N_832);
nor U1215 (N_1215,N_661,In_1324);
and U1216 (N_1216,N_837,N_948);
and U1217 (N_1217,N_403,N_600);
nor U1218 (N_1218,In_617,N_603);
or U1219 (N_1219,In_929,In_461);
and U1220 (N_1220,In_1815,N_775);
nor U1221 (N_1221,N_906,N_868);
nor U1222 (N_1222,N_916,In_1112);
or U1223 (N_1223,N_963,In_1811);
nor U1224 (N_1224,N_794,N_510);
or U1225 (N_1225,N_236,N_186);
nand U1226 (N_1226,N_544,N_760);
or U1227 (N_1227,N_712,In_1111);
nor U1228 (N_1228,N_164,N_945);
and U1229 (N_1229,N_522,N_525);
or U1230 (N_1230,N_941,N_595);
nor U1231 (N_1231,N_829,N_469);
or U1232 (N_1232,N_577,N_202);
and U1233 (N_1233,N_800,In_1841);
nand U1234 (N_1234,N_900,N_434);
nand U1235 (N_1235,In_789,N_545);
or U1236 (N_1236,In_330,N_976);
and U1237 (N_1237,In_372,In_17);
or U1238 (N_1238,N_396,N_727);
nand U1239 (N_1239,N_467,N_922);
nor U1240 (N_1240,N_273,In_1428);
or U1241 (N_1241,N_751,N_869);
or U1242 (N_1242,In_1131,N_267);
nor U1243 (N_1243,In_1138,N_938);
and U1244 (N_1244,N_308,N_781);
and U1245 (N_1245,N_150,N_591);
nor U1246 (N_1246,N_616,N_617);
or U1247 (N_1247,In_1660,In_730);
and U1248 (N_1248,In_407,In_969);
and U1249 (N_1249,N_977,In_608);
or U1250 (N_1250,N_967,N_951);
nand U1251 (N_1251,N_897,In_1184);
or U1252 (N_1252,In_1738,In_1165);
nand U1253 (N_1253,N_695,N_575);
and U1254 (N_1254,N_590,N_275);
nand U1255 (N_1255,In_793,N_131);
nand U1256 (N_1256,N_520,N_816);
and U1257 (N_1257,N_598,N_304);
or U1258 (N_1258,N_964,N_730);
or U1259 (N_1259,N_955,N_830);
or U1260 (N_1260,In_496,N_557);
or U1261 (N_1261,N_584,N_902);
nor U1262 (N_1262,N_959,In_1082);
or U1263 (N_1263,In_1120,In_448);
xnor U1264 (N_1264,In_43,N_981);
nand U1265 (N_1265,N_968,N_815);
nand U1266 (N_1266,N_583,N_60);
nand U1267 (N_1267,N_870,N_566);
nor U1268 (N_1268,N_592,N_878);
and U1269 (N_1269,N_856,N_30);
nor U1270 (N_1270,N_879,In_1342);
and U1271 (N_1271,N_898,N_834);
or U1272 (N_1272,In_1903,In_821);
or U1273 (N_1273,N_806,In_1541);
or U1274 (N_1274,In_626,In_1227);
nor U1275 (N_1275,In_1790,N_658);
nand U1276 (N_1276,N_737,In_1091);
and U1277 (N_1277,N_78,In_231);
nor U1278 (N_1278,N_907,N_638);
xnor U1279 (N_1279,In_1336,N_969);
nor U1280 (N_1280,In_1276,In_917);
or U1281 (N_1281,In_1432,In_1183);
nand U1282 (N_1282,In_970,N_970);
nor U1283 (N_1283,N_190,In_1816);
or U1284 (N_1284,N_119,In_362);
and U1285 (N_1285,N_961,N_84);
nor U1286 (N_1286,N_812,N_767);
or U1287 (N_1287,N_783,N_722);
nor U1288 (N_1288,N_158,In_1173);
nor U1289 (N_1289,In_238,N_232);
nor U1290 (N_1290,In_536,In_1451);
and U1291 (N_1291,In_828,In_102);
nand U1292 (N_1292,N_852,N_747);
and U1293 (N_1293,In_1945,In_300);
or U1294 (N_1294,N_855,In_87);
or U1295 (N_1295,N_719,N_672);
or U1296 (N_1296,N_935,In_1271);
nor U1297 (N_1297,N_711,In_745);
nand U1298 (N_1298,N_620,In_115);
xnor U1299 (N_1299,N_973,N_792);
nor U1300 (N_1300,In_1918,N_825);
or U1301 (N_1301,N_559,In_989);
or U1302 (N_1302,In_1594,N_383);
and U1303 (N_1303,N_857,In_148);
nand U1304 (N_1304,N_888,N_683);
nand U1305 (N_1305,In_724,In_348);
or U1306 (N_1306,In_1443,N_547);
nor U1307 (N_1307,N_85,In_1646);
xnor U1308 (N_1308,In_515,In_843);
nand U1309 (N_1309,N_689,N_551);
nor U1310 (N_1310,N_665,N_284);
nand U1311 (N_1311,In_1742,N_693);
nor U1312 (N_1312,N_631,N_412);
or U1313 (N_1313,N_440,In_565);
nand U1314 (N_1314,N_802,In_1056);
or U1315 (N_1315,N_621,In_1911);
nor U1316 (N_1316,N_960,N_459);
xor U1317 (N_1317,N_104,In_1233);
nor U1318 (N_1318,In_1557,N_984);
nand U1319 (N_1319,In_1458,N_729);
nand U1320 (N_1320,In_1615,N_745);
and U1321 (N_1321,N_803,In_725);
nand U1322 (N_1322,N_506,In_1864);
or U1323 (N_1323,N_835,N_989);
nand U1324 (N_1324,N_861,N_854);
or U1325 (N_1325,N_987,N_804);
and U1326 (N_1326,N_717,In_757);
nand U1327 (N_1327,In_1128,N_709);
nor U1328 (N_1328,N_483,N_309);
nor U1329 (N_1329,In_1780,N_756);
and U1330 (N_1330,N_998,N_847);
nor U1331 (N_1331,N_640,N_536);
nand U1332 (N_1332,N_924,N_673);
nor U1333 (N_1333,N_908,N_979);
or U1334 (N_1334,In_70,N_877);
or U1335 (N_1335,N_750,In_1071);
and U1336 (N_1336,In_1625,In_1781);
or U1337 (N_1337,In_79,N_953);
nand U1338 (N_1338,In_681,N_234);
and U1339 (N_1339,N_605,N_822);
nor U1340 (N_1340,In_1333,N_574);
nand U1341 (N_1341,In_727,N_754);
nand U1342 (N_1342,N_778,N_126);
nor U1343 (N_1343,N_788,N_533);
and U1344 (N_1344,In_315,In_1854);
xnor U1345 (N_1345,N_909,In_1937);
nand U1346 (N_1346,In_423,N_524);
and U1347 (N_1347,In_1544,In_1847);
and U1348 (N_1348,N_884,N_827);
or U1349 (N_1349,In_1406,N_379);
nor U1350 (N_1350,N_145,N_606);
or U1351 (N_1351,N_738,N_876);
or U1352 (N_1352,N_882,N_579);
or U1353 (N_1353,N_24,In_815);
nand U1354 (N_1354,N_954,N_140);
nand U1355 (N_1355,N_63,N_928);
nor U1356 (N_1356,N_587,In_1161);
or U1357 (N_1357,N_204,N_859);
nand U1358 (N_1358,In_160,N_813);
and U1359 (N_1359,In_331,In_1703);
or U1360 (N_1360,In_842,N_912);
and U1361 (N_1361,N_846,In_1531);
or U1362 (N_1362,In_425,N_512);
and U1363 (N_1363,N_242,N_513);
or U1364 (N_1364,N_265,N_102);
or U1365 (N_1365,N_72,N_618);
and U1366 (N_1366,N_487,N_798);
or U1367 (N_1367,N_886,In_1430);
and U1368 (N_1368,In_1898,N_22);
or U1369 (N_1369,N_759,N_691);
nor U1370 (N_1370,N_801,N_653);
nand U1371 (N_1371,In_139,N_589);
and U1372 (N_1372,N_739,N_183);
or U1373 (N_1373,N_624,In_1736);
nand U1374 (N_1374,N_950,N_344);
nand U1375 (N_1375,In_9,N_666);
nand U1376 (N_1376,N_871,N_682);
and U1377 (N_1377,N_927,N_958);
and U1378 (N_1378,In_220,In_1872);
and U1379 (N_1379,N_573,In_394);
and U1380 (N_1380,N_12,N_26);
or U1381 (N_1381,In_1806,In_387);
nor U1382 (N_1382,N_397,In_1586);
nor U1383 (N_1383,N_838,In_784);
nor U1384 (N_1384,N_393,N_771);
nor U1385 (N_1385,N_71,N_793);
nor U1386 (N_1386,N_742,N_558);
or U1387 (N_1387,N_542,N_651);
nand U1388 (N_1388,N_307,N_644);
or U1389 (N_1389,In_737,In_470);
or U1390 (N_1390,In_631,In_1156);
nand U1391 (N_1391,N_786,In_155);
nand U1392 (N_1392,In_1643,N_991);
or U1393 (N_1393,In_683,In_359);
or U1394 (N_1394,N_639,N_817);
nor U1395 (N_1395,N_919,In_521);
and U1396 (N_1396,In_1870,N_923);
nand U1397 (N_1397,N_896,N_677);
nand U1398 (N_1398,In_1754,N_685);
nand U1399 (N_1399,N_507,N_159);
nor U1400 (N_1400,In_144,N_502);
nor U1401 (N_1401,N_669,In_1026);
nor U1402 (N_1402,N_990,In_1940);
nor U1403 (N_1403,In_1824,In_558);
nor U1404 (N_1404,In_141,In_896);
nor U1405 (N_1405,In_1881,In_421);
or U1406 (N_1406,In_581,N_567);
or U1407 (N_1407,In_947,In_936);
or U1408 (N_1408,N_873,N_674);
nand U1409 (N_1409,N_457,N_784);
or U1410 (N_1410,N_790,In_1232);
and U1411 (N_1411,N_153,N_777);
nand U1412 (N_1412,N_872,N_648);
and U1413 (N_1413,N_576,N_538);
or U1414 (N_1414,N_360,N_646);
nor U1415 (N_1415,N_552,N_423);
and U1416 (N_1416,In_1234,In_1377);
and U1417 (N_1417,N_254,N_892);
and U1418 (N_1418,N_721,In_1006);
nor U1419 (N_1419,N_996,In_1976);
nand U1420 (N_1420,N_860,N_2);
and U1421 (N_1421,N_287,N_688);
nor U1422 (N_1422,In_621,N_471);
xnor U1423 (N_1423,In_1003,In_1504);
and U1424 (N_1424,N_599,N_328);
nor U1425 (N_1425,N_539,N_956);
and U1426 (N_1426,N_548,In_1669);
or U1427 (N_1427,N_752,N_625);
nand U1428 (N_1428,N_546,In_306);
nand U1429 (N_1429,N_531,N_47);
nand U1430 (N_1430,N_503,N_814);
or U1431 (N_1431,In_28,In_988);
nand U1432 (N_1432,N_239,N_780);
and U1433 (N_1433,N_569,In_1916);
and U1434 (N_1434,In_671,N_196);
nand U1435 (N_1435,N_943,N_115);
and U1436 (N_1436,N_135,N_942);
xor U1437 (N_1437,N_710,In_1968);
nor U1438 (N_1438,N_678,N_409);
nand U1439 (N_1439,N_514,N_147);
or U1440 (N_1440,In_1709,N_477);
nor U1441 (N_1441,N_937,N_840);
nor U1442 (N_1442,In_1867,In_1057);
or U1443 (N_1443,N_933,N_626);
nand U1444 (N_1444,N_949,N_939);
nor U1445 (N_1445,In_627,N_210);
or U1446 (N_1446,N_452,N_944);
nand U1447 (N_1447,N_515,N_845);
nand U1448 (N_1448,N_761,N_67);
or U1449 (N_1449,N_650,N_887);
nor U1450 (N_1450,N_733,In_1953);
nor U1451 (N_1451,N_562,N_980);
xor U1452 (N_1452,N_281,In_895);
nand U1453 (N_1453,In_1661,N_550);
and U1454 (N_1454,N_844,N_664);
nand U1455 (N_1455,In_556,In_1109);
nor U1456 (N_1456,N_280,N_715);
or U1457 (N_1457,N_918,N_796);
or U1458 (N_1458,N_740,In_1329);
nand U1459 (N_1459,N_657,N_641);
nor U1460 (N_1460,N_926,N_940);
and U1461 (N_1461,N_518,N_843);
nor U1462 (N_1462,In_1698,N_999);
and U1463 (N_1463,In_152,N_349);
or U1464 (N_1464,N_851,N_974);
and U1465 (N_1465,N_748,N_312);
nor U1466 (N_1466,In_1631,N_824);
and U1467 (N_1467,In_604,N_564);
nand U1468 (N_1468,N_460,In_897);
nor U1469 (N_1469,In_253,In_8);
or U1470 (N_1470,In_908,In_1414);
nor U1471 (N_1471,N_972,N_622);
nor U1472 (N_1472,N_684,N_519);
nor U1473 (N_1473,In_374,In_1252);
nand U1474 (N_1474,N_910,In_494);
and U1475 (N_1475,In_1185,N_99);
and U1476 (N_1476,In_1821,N_224);
nor U1477 (N_1477,In_192,N_32);
nor U1478 (N_1478,N_805,In_1566);
and U1479 (N_1479,N_654,N_169);
nor U1480 (N_1480,In_321,N_535);
xnor U1481 (N_1481,N_930,N_465);
nor U1482 (N_1482,N_687,N_735);
and U1483 (N_1483,N_373,N_947);
and U1484 (N_1484,N_901,N_95);
and U1485 (N_1485,N_101,N_808);
nor U1486 (N_1486,N_500,In_1554);
nor U1487 (N_1487,In_1965,N_893);
nor U1488 (N_1488,N_380,N_537);
and U1489 (N_1489,In_1724,N_643);
nand U1490 (N_1490,N_136,In_906);
and U1491 (N_1491,In_1946,N_702);
nor U1492 (N_1492,In_64,N_565);
nor U1493 (N_1493,N_121,In_1215);
nand U1494 (N_1494,N_997,In_1920);
nand U1495 (N_1495,N_776,N_250);
and U1496 (N_1496,N_770,In_171);
nor U1497 (N_1497,N_637,N_993);
nor U1498 (N_1498,N_223,N_821);
nand U1499 (N_1499,In_130,N_766);
nand U1500 (N_1500,N_1436,N_1138);
and U1501 (N_1501,N_1231,N_1479);
nor U1502 (N_1502,N_1449,N_1053);
or U1503 (N_1503,N_1492,N_1294);
nand U1504 (N_1504,N_1391,N_1260);
nand U1505 (N_1505,N_1451,N_1413);
nand U1506 (N_1506,N_1111,N_1181);
nor U1507 (N_1507,N_1196,N_1408);
and U1508 (N_1508,N_1169,N_1210);
nand U1509 (N_1509,N_1163,N_1175);
or U1510 (N_1510,N_1070,N_1208);
or U1511 (N_1511,N_1377,N_1179);
and U1512 (N_1512,N_1452,N_1368);
or U1513 (N_1513,N_1085,N_1024);
and U1514 (N_1514,N_1469,N_1109);
nor U1515 (N_1515,N_1438,N_1284);
nand U1516 (N_1516,N_1228,N_1456);
nand U1517 (N_1517,N_1427,N_1470);
nor U1518 (N_1518,N_1097,N_1343);
nor U1519 (N_1519,N_1001,N_1203);
nand U1520 (N_1520,N_1201,N_1441);
nor U1521 (N_1521,N_1014,N_1009);
and U1522 (N_1522,N_1158,N_1033);
nor U1523 (N_1523,N_1172,N_1326);
or U1524 (N_1524,N_1266,N_1322);
nand U1525 (N_1525,N_1274,N_1037);
nand U1526 (N_1526,N_1405,N_1161);
and U1527 (N_1527,N_1299,N_1047);
and U1528 (N_1528,N_1307,N_1333);
nand U1529 (N_1529,N_1240,N_1280);
nor U1530 (N_1530,N_1151,N_1335);
or U1531 (N_1531,N_1485,N_1336);
nand U1532 (N_1532,N_1011,N_1200);
or U1533 (N_1533,N_1372,N_1384);
and U1534 (N_1534,N_1184,N_1481);
or U1535 (N_1535,N_1004,N_1232);
or U1536 (N_1536,N_1360,N_1348);
and U1537 (N_1537,N_1282,N_1153);
and U1538 (N_1538,N_1244,N_1426);
nor U1539 (N_1539,N_1304,N_1386);
and U1540 (N_1540,N_1027,N_1084);
or U1541 (N_1541,N_1021,N_1393);
nand U1542 (N_1542,N_1023,N_1300);
or U1543 (N_1543,N_1136,N_1221);
and U1544 (N_1544,N_1341,N_1418);
and U1545 (N_1545,N_1134,N_1132);
and U1546 (N_1546,N_1432,N_1054);
and U1547 (N_1547,N_1370,N_1487);
nand U1548 (N_1548,N_1482,N_1057);
or U1549 (N_1549,N_1433,N_1465);
nand U1550 (N_1550,N_1440,N_1050);
and U1551 (N_1551,N_1499,N_1474);
or U1552 (N_1552,N_1303,N_1058);
nor U1553 (N_1553,N_1291,N_1059);
or U1554 (N_1554,N_1013,N_1356);
and U1555 (N_1555,N_1270,N_1403);
nor U1556 (N_1556,N_1218,N_1083);
and U1557 (N_1557,N_1020,N_1064);
and U1558 (N_1558,N_1030,N_1026);
nor U1559 (N_1559,N_1332,N_1293);
nand U1560 (N_1560,N_1347,N_1416);
nand U1561 (N_1561,N_1353,N_1351);
nand U1562 (N_1562,N_1005,N_1486);
or U1563 (N_1563,N_1042,N_1071);
nand U1564 (N_1564,N_1325,N_1252);
and U1565 (N_1565,N_1073,N_1204);
nor U1566 (N_1566,N_1334,N_1242);
and U1567 (N_1567,N_1245,N_1087);
nor U1568 (N_1568,N_1223,N_1066);
and U1569 (N_1569,N_1226,N_1437);
nand U1570 (N_1570,N_1146,N_1301);
nor U1571 (N_1571,N_1421,N_1285);
or U1572 (N_1572,N_1396,N_1114);
and U1573 (N_1573,N_1034,N_1116);
or U1574 (N_1574,N_1106,N_1435);
nand U1575 (N_1575,N_1189,N_1081);
nand U1576 (N_1576,N_1044,N_1170);
nor U1577 (N_1577,N_1458,N_1061);
nor U1578 (N_1578,N_1447,N_1233);
or U1579 (N_1579,N_1191,N_1174);
nor U1580 (N_1580,N_1075,N_1092);
nand U1581 (N_1581,N_1103,N_1065);
or U1582 (N_1582,N_1466,N_1067);
nor U1583 (N_1583,N_1471,N_1430);
or U1584 (N_1584,N_1467,N_1096);
or U1585 (N_1585,N_1168,N_1248);
and U1586 (N_1586,N_1329,N_1354);
or U1587 (N_1587,N_1213,N_1055);
and U1588 (N_1588,N_1150,N_1239);
or U1589 (N_1589,N_1025,N_1137);
or U1590 (N_1590,N_1445,N_1464);
nor U1591 (N_1591,N_1258,N_1115);
or U1592 (N_1592,N_1344,N_1394);
and U1593 (N_1593,N_1273,N_1323);
and U1594 (N_1594,N_1331,N_1399);
and U1595 (N_1595,N_1383,N_1375);
nand U1596 (N_1596,N_1045,N_1450);
or U1597 (N_1597,N_1147,N_1080);
or U1598 (N_1598,N_1359,N_1094);
nor U1599 (N_1599,N_1446,N_1357);
nor U1600 (N_1600,N_1246,N_1063);
or U1601 (N_1601,N_1389,N_1443);
or U1602 (N_1602,N_1180,N_1488);
nand U1603 (N_1603,N_1475,N_1490);
and U1604 (N_1604,N_1090,N_1062);
or U1605 (N_1605,N_1288,N_1306);
or U1606 (N_1606,N_1156,N_1207);
or U1607 (N_1607,N_1091,N_1038);
and U1608 (N_1608,N_1035,N_1483);
and U1609 (N_1609,N_1298,N_1216);
or U1610 (N_1610,N_1363,N_1039);
and U1611 (N_1611,N_1310,N_1448);
nor U1612 (N_1612,N_1126,N_1374);
or U1613 (N_1613,N_1002,N_1143);
and U1614 (N_1614,N_1197,N_1472);
xnor U1615 (N_1615,N_1496,N_1439);
or U1616 (N_1616,N_1355,N_1086);
nor U1617 (N_1617,N_1032,N_1415);
or U1618 (N_1618,N_1366,N_1192);
or U1619 (N_1619,N_1017,N_1202);
and U1620 (N_1620,N_1468,N_1337);
or U1621 (N_1621,N_1262,N_1398);
and U1622 (N_1622,N_1183,N_1302);
nand U1623 (N_1623,N_1295,N_1498);
or U1624 (N_1624,N_1431,N_1493);
or U1625 (N_1625,N_1473,N_1477);
or U1626 (N_1626,N_1238,N_1434);
and U1627 (N_1627,N_1041,N_1100);
and U1628 (N_1628,N_1049,N_1319);
nand U1629 (N_1629,N_1243,N_1124);
or U1630 (N_1630,N_1236,N_1235);
nor U1631 (N_1631,N_1271,N_1406);
nor U1632 (N_1632,N_1123,N_1480);
or U1633 (N_1633,N_1186,N_1358);
or U1634 (N_1634,N_1107,N_1060);
or U1635 (N_1635,N_1118,N_1423);
nor U1636 (N_1636,N_1308,N_1278);
and U1637 (N_1637,N_1251,N_1379);
nor U1638 (N_1638,N_1089,N_1407);
nor U1639 (N_1639,N_1157,N_1364);
and U1640 (N_1640,N_1108,N_1410);
or U1641 (N_1641,N_1387,N_1217);
and U1642 (N_1642,N_1140,N_1209);
or U1643 (N_1643,N_1112,N_1402);
and U1644 (N_1644,N_1076,N_1442);
nor U1645 (N_1645,N_1162,N_1489);
or U1646 (N_1646,N_1129,N_1234);
or U1647 (N_1647,N_1411,N_1088);
nor U1648 (N_1648,N_1267,N_1018);
or U1649 (N_1649,N_1424,N_1257);
nand U1650 (N_1650,N_1247,N_1139);
nor U1651 (N_1651,N_1255,N_1012);
and U1652 (N_1652,N_1036,N_1376);
and U1653 (N_1653,N_1164,N_1417);
or U1654 (N_1654,N_1269,N_1225);
nand U1655 (N_1655,N_1367,N_1149);
nand U1656 (N_1656,N_1212,N_1029);
or U1657 (N_1657,N_1105,N_1457);
nand U1658 (N_1658,N_1342,N_1313);
and U1659 (N_1659,N_1078,N_1484);
nand U1660 (N_1660,N_1382,N_1371);
nand U1661 (N_1661,N_1215,N_1093);
nor U1662 (N_1662,N_1194,N_1127);
nor U1663 (N_1663,N_1429,N_1072);
or U1664 (N_1664,N_1077,N_1206);
or U1665 (N_1665,N_1462,N_1121);
or U1666 (N_1666,N_1340,N_1350);
or U1667 (N_1667,N_1287,N_1224);
or U1668 (N_1668,N_1193,N_1292);
nor U1669 (N_1669,N_1128,N_1229);
and U1670 (N_1670,N_1199,N_1476);
nand U1671 (N_1671,N_1178,N_1003);
or U1672 (N_1672,N_1276,N_1000);
and U1673 (N_1673,N_1414,N_1491);
nand U1674 (N_1674,N_1283,N_1290);
nand U1675 (N_1675,N_1316,N_1380);
or U1676 (N_1676,N_1214,N_1385);
or U1677 (N_1677,N_1122,N_1007);
or U1678 (N_1678,N_1422,N_1110);
nand U1679 (N_1679,N_1141,N_1237);
nor U1680 (N_1680,N_1079,N_1040);
and U1681 (N_1681,N_1052,N_1051);
nand U1682 (N_1682,N_1056,N_1272);
or U1683 (N_1683,N_1119,N_1265);
nor U1684 (N_1684,N_1152,N_1173);
and U1685 (N_1685,N_1145,N_1428);
and U1686 (N_1686,N_1275,N_1185);
nor U1687 (N_1687,N_1125,N_1074);
nand U1688 (N_1688,N_1098,N_1155);
or U1689 (N_1689,N_1043,N_1095);
and U1690 (N_1690,N_1268,N_1130);
nand U1691 (N_1691,N_1345,N_1305);
nand U1692 (N_1692,N_1362,N_1425);
and U1693 (N_1693,N_1286,N_1453);
nor U1694 (N_1694,N_1068,N_1241);
nor U1695 (N_1695,N_1346,N_1311);
and U1696 (N_1696,N_1222,N_1019);
nand U1697 (N_1697,N_1378,N_1006);
and U1698 (N_1698,N_1412,N_1395);
or U1699 (N_1699,N_1135,N_1198);
and U1700 (N_1700,N_1016,N_1008);
nand U1701 (N_1701,N_1176,N_1230);
or U1702 (N_1702,N_1166,N_1069);
xor U1703 (N_1703,N_1381,N_1419);
nor U1704 (N_1704,N_1361,N_1205);
nand U1705 (N_1705,N_1082,N_1390);
nor U1706 (N_1706,N_1314,N_1478);
or U1707 (N_1707,N_1142,N_1369);
or U1708 (N_1708,N_1324,N_1165);
or U1709 (N_1709,N_1289,N_1373);
nand U1710 (N_1710,N_1159,N_1349);
nor U1711 (N_1711,N_1400,N_1022);
and U1712 (N_1712,N_1171,N_1296);
nand U1713 (N_1713,N_1250,N_1028);
nand U1714 (N_1714,N_1015,N_1120);
or U1715 (N_1715,N_1167,N_1277);
nand U1716 (N_1716,N_1392,N_1317);
nand U1717 (N_1717,N_1494,N_1048);
nor U1718 (N_1718,N_1321,N_1031);
nand U1719 (N_1719,N_1160,N_1104);
nor U1720 (N_1720,N_1144,N_1388);
and U1721 (N_1721,N_1154,N_1297);
and U1722 (N_1722,N_1312,N_1454);
nand U1723 (N_1723,N_1279,N_1188);
or U1724 (N_1724,N_1328,N_1460);
nor U1725 (N_1725,N_1249,N_1117);
and U1726 (N_1726,N_1113,N_1404);
xnor U1727 (N_1727,N_1339,N_1261);
or U1728 (N_1728,N_1309,N_1338);
or U1729 (N_1729,N_1259,N_1330);
and U1730 (N_1730,N_1263,N_1131);
nand U1731 (N_1731,N_1461,N_1102);
nand U1732 (N_1732,N_1497,N_1211);
nor U1733 (N_1733,N_1133,N_1409);
or U1734 (N_1734,N_1352,N_1010);
nand U1735 (N_1735,N_1318,N_1420);
and U1736 (N_1736,N_1397,N_1365);
or U1737 (N_1737,N_1459,N_1148);
or U1738 (N_1738,N_1253,N_1101);
nand U1739 (N_1739,N_1182,N_1190);
and U1740 (N_1740,N_1099,N_1254);
and U1741 (N_1741,N_1327,N_1220);
nand U1742 (N_1742,N_1187,N_1455);
nor U1743 (N_1743,N_1401,N_1495);
and U1744 (N_1744,N_1264,N_1320);
and U1745 (N_1745,N_1227,N_1046);
nand U1746 (N_1746,N_1219,N_1444);
and U1747 (N_1747,N_1281,N_1177);
nand U1748 (N_1748,N_1315,N_1195);
nand U1749 (N_1749,N_1256,N_1463);
or U1750 (N_1750,N_1202,N_1008);
and U1751 (N_1751,N_1480,N_1205);
nand U1752 (N_1752,N_1144,N_1061);
nand U1753 (N_1753,N_1156,N_1103);
nor U1754 (N_1754,N_1257,N_1328);
nor U1755 (N_1755,N_1359,N_1223);
or U1756 (N_1756,N_1044,N_1202);
nand U1757 (N_1757,N_1208,N_1293);
nor U1758 (N_1758,N_1230,N_1309);
xor U1759 (N_1759,N_1122,N_1496);
nand U1760 (N_1760,N_1133,N_1032);
and U1761 (N_1761,N_1053,N_1105);
or U1762 (N_1762,N_1052,N_1466);
nand U1763 (N_1763,N_1098,N_1254);
or U1764 (N_1764,N_1489,N_1089);
or U1765 (N_1765,N_1399,N_1199);
and U1766 (N_1766,N_1416,N_1359);
and U1767 (N_1767,N_1221,N_1339);
nand U1768 (N_1768,N_1481,N_1240);
nand U1769 (N_1769,N_1449,N_1130);
nand U1770 (N_1770,N_1368,N_1052);
and U1771 (N_1771,N_1208,N_1034);
nand U1772 (N_1772,N_1273,N_1188);
or U1773 (N_1773,N_1042,N_1357);
and U1774 (N_1774,N_1318,N_1212);
nor U1775 (N_1775,N_1298,N_1247);
and U1776 (N_1776,N_1278,N_1434);
nor U1777 (N_1777,N_1239,N_1105);
and U1778 (N_1778,N_1475,N_1183);
or U1779 (N_1779,N_1488,N_1235);
nor U1780 (N_1780,N_1483,N_1428);
nand U1781 (N_1781,N_1159,N_1219);
nand U1782 (N_1782,N_1145,N_1391);
nor U1783 (N_1783,N_1011,N_1429);
nor U1784 (N_1784,N_1116,N_1017);
nor U1785 (N_1785,N_1010,N_1278);
nor U1786 (N_1786,N_1245,N_1111);
or U1787 (N_1787,N_1456,N_1116);
and U1788 (N_1788,N_1294,N_1378);
nand U1789 (N_1789,N_1414,N_1144);
nand U1790 (N_1790,N_1233,N_1237);
xnor U1791 (N_1791,N_1026,N_1101);
nor U1792 (N_1792,N_1181,N_1435);
nand U1793 (N_1793,N_1487,N_1165);
and U1794 (N_1794,N_1031,N_1372);
nor U1795 (N_1795,N_1401,N_1088);
nand U1796 (N_1796,N_1079,N_1461);
nand U1797 (N_1797,N_1429,N_1325);
and U1798 (N_1798,N_1301,N_1479);
or U1799 (N_1799,N_1156,N_1248);
nor U1800 (N_1800,N_1460,N_1395);
and U1801 (N_1801,N_1096,N_1074);
and U1802 (N_1802,N_1481,N_1489);
or U1803 (N_1803,N_1230,N_1020);
or U1804 (N_1804,N_1056,N_1097);
nor U1805 (N_1805,N_1381,N_1384);
or U1806 (N_1806,N_1060,N_1467);
or U1807 (N_1807,N_1101,N_1209);
nor U1808 (N_1808,N_1152,N_1243);
nor U1809 (N_1809,N_1288,N_1469);
nand U1810 (N_1810,N_1079,N_1130);
and U1811 (N_1811,N_1428,N_1076);
nor U1812 (N_1812,N_1030,N_1290);
and U1813 (N_1813,N_1241,N_1418);
and U1814 (N_1814,N_1172,N_1167);
and U1815 (N_1815,N_1217,N_1160);
nand U1816 (N_1816,N_1337,N_1135);
and U1817 (N_1817,N_1060,N_1339);
or U1818 (N_1818,N_1042,N_1269);
or U1819 (N_1819,N_1456,N_1076);
or U1820 (N_1820,N_1344,N_1107);
nor U1821 (N_1821,N_1291,N_1281);
and U1822 (N_1822,N_1143,N_1011);
nor U1823 (N_1823,N_1141,N_1369);
nand U1824 (N_1824,N_1319,N_1490);
nor U1825 (N_1825,N_1134,N_1211);
nor U1826 (N_1826,N_1018,N_1020);
nand U1827 (N_1827,N_1270,N_1005);
nor U1828 (N_1828,N_1118,N_1401);
and U1829 (N_1829,N_1071,N_1462);
nor U1830 (N_1830,N_1321,N_1477);
and U1831 (N_1831,N_1360,N_1376);
nor U1832 (N_1832,N_1064,N_1238);
nand U1833 (N_1833,N_1337,N_1282);
nand U1834 (N_1834,N_1176,N_1291);
nand U1835 (N_1835,N_1146,N_1398);
nor U1836 (N_1836,N_1123,N_1297);
or U1837 (N_1837,N_1465,N_1299);
and U1838 (N_1838,N_1408,N_1418);
nor U1839 (N_1839,N_1156,N_1470);
nor U1840 (N_1840,N_1320,N_1273);
or U1841 (N_1841,N_1229,N_1467);
or U1842 (N_1842,N_1022,N_1446);
and U1843 (N_1843,N_1156,N_1380);
and U1844 (N_1844,N_1002,N_1236);
nand U1845 (N_1845,N_1344,N_1333);
and U1846 (N_1846,N_1306,N_1009);
or U1847 (N_1847,N_1023,N_1380);
or U1848 (N_1848,N_1221,N_1114);
nand U1849 (N_1849,N_1109,N_1191);
and U1850 (N_1850,N_1389,N_1129);
and U1851 (N_1851,N_1166,N_1351);
or U1852 (N_1852,N_1360,N_1230);
and U1853 (N_1853,N_1055,N_1414);
nand U1854 (N_1854,N_1265,N_1474);
nor U1855 (N_1855,N_1171,N_1223);
or U1856 (N_1856,N_1074,N_1126);
or U1857 (N_1857,N_1215,N_1227);
and U1858 (N_1858,N_1469,N_1272);
nand U1859 (N_1859,N_1166,N_1189);
nor U1860 (N_1860,N_1226,N_1320);
and U1861 (N_1861,N_1375,N_1129);
nand U1862 (N_1862,N_1155,N_1146);
nand U1863 (N_1863,N_1226,N_1401);
and U1864 (N_1864,N_1322,N_1068);
or U1865 (N_1865,N_1035,N_1045);
and U1866 (N_1866,N_1484,N_1003);
nor U1867 (N_1867,N_1445,N_1187);
or U1868 (N_1868,N_1462,N_1460);
or U1869 (N_1869,N_1189,N_1232);
and U1870 (N_1870,N_1153,N_1353);
and U1871 (N_1871,N_1211,N_1201);
or U1872 (N_1872,N_1391,N_1085);
and U1873 (N_1873,N_1177,N_1494);
nand U1874 (N_1874,N_1140,N_1418);
or U1875 (N_1875,N_1152,N_1220);
nor U1876 (N_1876,N_1040,N_1421);
and U1877 (N_1877,N_1008,N_1087);
nor U1878 (N_1878,N_1025,N_1427);
nor U1879 (N_1879,N_1289,N_1108);
nor U1880 (N_1880,N_1048,N_1440);
nor U1881 (N_1881,N_1378,N_1298);
nand U1882 (N_1882,N_1131,N_1496);
or U1883 (N_1883,N_1298,N_1166);
nand U1884 (N_1884,N_1431,N_1448);
or U1885 (N_1885,N_1325,N_1490);
nand U1886 (N_1886,N_1495,N_1166);
and U1887 (N_1887,N_1245,N_1198);
and U1888 (N_1888,N_1448,N_1265);
nand U1889 (N_1889,N_1355,N_1177);
nor U1890 (N_1890,N_1189,N_1172);
or U1891 (N_1891,N_1390,N_1289);
and U1892 (N_1892,N_1141,N_1445);
nor U1893 (N_1893,N_1174,N_1480);
nand U1894 (N_1894,N_1494,N_1120);
and U1895 (N_1895,N_1296,N_1014);
and U1896 (N_1896,N_1331,N_1222);
nor U1897 (N_1897,N_1060,N_1211);
nand U1898 (N_1898,N_1303,N_1011);
nor U1899 (N_1899,N_1264,N_1334);
and U1900 (N_1900,N_1002,N_1426);
and U1901 (N_1901,N_1007,N_1493);
and U1902 (N_1902,N_1406,N_1478);
nand U1903 (N_1903,N_1499,N_1452);
or U1904 (N_1904,N_1062,N_1497);
and U1905 (N_1905,N_1048,N_1424);
or U1906 (N_1906,N_1435,N_1214);
or U1907 (N_1907,N_1333,N_1216);
nand U1908 (N_1908,N_1252,N_1432);
and U1909 (N_1909,N_1427,N_1435);
and U1910 (N_1910,N_1344,N_1095);
nor U1911 (N_1911,N_1392,N_1094);
nand U1912 (N_1912,N_1421,N_1490);
or U1913 (N_1913,N_1414,N_1061);
nor U1914 (N_1914,N_1242,N_1015);
nor U1915 (N_1915,N_1290,N_1396);
or U1916 (N_1916,N_1334,N_1141);
or U1917 (N_1917,N_1499,N_1425);
nand U1918 (N_1918,N_1041,N_1231);
and U1919 (N_1919,N_1262,N_1348);
and U1920 (N_1920,N_1221,N_1389);
nand U1921 (N_1921,N_1374,N_1473);
nor U1922 (N_1922,N_1056,N_1226);
and U1923 (N_1923,N_1102,N_1286);
nor U1924 (N_1924,N_1435,N_1466);
nor U1925 (N_1925,N_1062,N_1318);
nand U1926 (N_1926,N_1241,N_1096);
nor U1927 (N_1927,N_1045,N_1466);
and U1928 (N_1928,N_1444,N_1342);
and U1929 (N_1929,N_1291,N_1283);
nand U1930 (N_1930,N_1409,N_1225);
nor U1931 (N_1931,N_1431,N_1460);
and U1932 (N_1932,N_1474,N_1087);
or U1933 (N_1933,N_1321,N_1169);
and U1934 (N_1934,N_1079,N_1486);
nand U1935 (N_1935,N_1171,N_1327);
nor U1936 (N_1936,N_1166,N_1429);
and U1937 (N_1937,N_1445,N_1076);
nor U1938 (N_1938,N_1275,N_1068);
nor U1939 (N_1939,N_1326,N_1103);
nand U1940 (N_1940,N_1216,N_1379);
or U1941 (N_1941,N_1182,N_1083);
or U1942 (N_1942,N_1171,N_1118);
and U1943 (N_1943,N_1277,N_1129);
or U1944 (N_1944,N_1120,N_1345);
nor U1945 (N_1945,N_1152,N_1286);
nand U1946 (N_1946,N_1186,N_1356);
nand U1947 (N_1947,N_1229,N_1028);
or U1948 (N_1948,N_1275,N_1137);
nor U1949 (N_1949,N_1278,N_1217);
or U1950 (N_1950,N_1184,N_1231);
nand U1951 (N_1951,N_1036,N_1347);
nor U1952 (N_1952,N_1097,N_1425);
nand U1953 (N_1953,N_1414,N_1252);
nand U1954 (N_1954,N_1453,N_1421);
nand U1955 (N_1955,N_1294,N_1367);
or U1956 (N_1956,N_1322,N_1109);
nand U1957 (N_1957,N_1035,N_1146);
and U1958 (N_1958,N_1115,N_1218);
nand U1959 (N_1959,N_1324,N_1482);
and U1960 (N_1960,N_1469,N_1365);
and U1961 (N_1961,N_1123,N_1340);
nand U1962 (N_1962,N_1110,N_1464);
and U1963 (N_1963,N_1389,N_1424);
nor U1964 (N_1964,N_1336,N_1393);
nand U1965 (N_1965,N_1207,N_1075);
nand U1966 (N_1966,N_1188,N_1378);
or U1967 (N_1967,N_1199,N_1447);
nor U1968 (N_1968,N_1032,N_1421);
nand U1969 (N_1969,N_1152,N_1427);
or U1970 (N_1970,N_1129,N_1173);
and U1971 (N_1971,N_1439,N_1434);
or U1972 (N_1972,N_1051,N_1201);
xor U1973 (N_1973,N_1037,N_1244);
nor U1974 (N_1974,N_1175,N_1241);
nor U1975 (N_1975,N_1492,N_1048);
nand U1976 (N_1976,N_1395,N_1279);
or U1977 (N_1977,N_1256,N_1041);
nand U1978 (N_1978,N_1037,N_1366);
nand U1979 (N_1979,N_1305,N_1211);
or U1980 (N_1980,N_1110,N_1202);
or U1981 (N_1981,N_1183,N_1000);
nand U1982 (N_1982,N_1147,N_1402);
and U1983 (N_1983,N_1400,N_1275);
or U1984 (N_1984,N_1168,N_1415);
nor U1985 (N_1985,N_1294,N_1472);
and U1986 (N_1986,N_1425,N_1435);
nand U1987 (N_1987,N_1279,N_1251);
and U1988 (N_1988,N_1149,N_1304);
or U1989 (N_1989,N_1206,N_1088);
nand U1990 (N_1990,N_1339,N_1420);
nor U1991 (N_1991,N_1324,N_1313);
nand U1992 (N_1992,N_1286,N_1123);
nand U1993 (N_1993,N_1124,N_1010);
nand U1994 (N_1994,N_1382,N_1196);
nand U1995 (N_1995,N_1102,N_1444);
or U1996 (N_1996,N_1106,N_1279);
nand U1997 (N_1997,N_1302,N_1499);
or U1998 (N_1998,N_1241,N_1426);
nor U1999 (N_1999,N_1133,N_1062);
nand U2000 (N_2000,N_1823,N_1820);
or U2001 (N_2001,N_1922,N_1819);
nand U2002 (N_2002,N_1904,N_1560);
and U2003 (N_2003,N_1759,N_1865);
and U2004 (N_2004,N_1968,N_1509);
nand U2005 (N_2005,N_1825,N_1885);
or U2006 (N_2006,N_1866,N_1650);
nand U2007 (N_2007,N_1649,N_1886);
nand U2008 (N_2008,N_1745,N_1986);
and U2009 (N_2009,N_1673,N_1752);
xnor U2010 (N_2010,N_1540,N_1903);
nor U2011 (N_2011,N_1973,N_1785);
and U2012 (N_2012,N_1623,N_1985);
nand U2013 (N_2013,N_1925,N_1889);
nor U2014 (N_2014,N_1854,N_1639);
and U2015 (N_2015,N_1891,N_1770);
or U2016 (N_2016,N_1954,N_1796);
nand U2017 (N_2017,N_1773,N_1593);
nand U2018 (N_2018,N_1665,N_1652);
nor U2019 (N_2019,N_1972,N_1746);
and U2020 (N_2020,N_1726,N_1520);
nand U2021 (N_2021,N_1531,N_1856);
nand U2022 (N_2022,N_1761,N_1533);
or U2023 (N_2023,N_1813,N_1918);
nand U2024 (N_2024,N_1681,N_1599);
and U2025 (N_2025,N_1682,N_1571);
nor U2026 (N_2026,N_1879,N_1655);
nor U2027 (N_2027,N_1651,N_1568);
or U2028 (N_2028,N_1948,N_1936);
or U2029 (N_2029,N_1843,N_1713);
nand U2030 (N_2030,N_1826,N_1640);
nor U2031 (N_2031,N_1578,N_1670);
and U2032 (N_2032,N_1778,N_1711);
nand U2033 (N_2033,N_1787,N_1645);
nor U2034 (N_2034,N_1878,N_1803);
and U2035 (N_2035,N_1589,N_1753);
nand U2036 (N_2036,N_1699,N_1888);
nand U2037 (N_2037,N_1953,N_1700);
nor U2038 (N_2038,N_1622,N_1905);
or U2039 (N_2039,N_1775,N_1992);
and U2040 (N_2040,N_1980,N_1989);
and U2041 (N_2041,N_1933,N_1798);
nand U2042 (N_2042,N_1527,N_1931);
and U2043 (N_2043,N_1841,N_1714);
xnor U2044 (N_2044,N_1698,N_1551);
or U2045 (N_2045,N_1988,N_1683);
and U2046 (N_2046,N_1707,N_1610);
and U2047 (N_2047,N_1940,N_1957);
nand U2048 (N_2048,N_1967,N_1774);
nor U2049 (N_2049,N_1704,N_1853);
and U2050 (N_2050,N_1884,N_1515);
nor U2051 (N_2051,N_1762,N_1519);
or U2052 (N_2052,N_1919,N_1597);
or U2053 (N_2053,N_1653,N_1934);
nand U2054 (N_2054,N_1847,N_1680);
or U2055 (N_2055,N_1620,N_1857);
and U2056 (N_2056,N_1812,N_1791);
nor U2057 (N_2057,N_1742,N_1976);
or U2058 (N_2058,N_1894,N_1522);
or U2059 (N_2059,N_1712,N_1732);
nand U2060 (N_2060,N_1757,N_1617);
or U2061 (N_2061,N_1626,N_1930);
and U2062 (N_2062,N_1910,N_1737);
or U2063 (N_2063,N_1873,N_1671);
nand U2064 (N_2064,N_1760,N_1830);
nand U2065 (N_2065,N_1600,N_1944);
nand U2066 (N_2066,N_1952,N_1928);
nor U2067 (N_2067,N_1780,N_1536);
or U2068 (N_2068,N_1902,N_1720);
or U2069 (N_2069,N_1662,N_1908);
xor U2070 (N_2070,N_1874,N_1521);
nand U2071 (N_2071,N_1828,N_1595);
and U2072 (N_2072,N_1999,N_1664);
and U2073 (N_2073,N_1821,N_1864);
nor U2074 (N_2074,N_1559,N_1604);
nor U2075 (N_2075,N_1781,N_1518);
nor U2076 (N_2076,N_1523,N_1790);
nor U2077 (N_2077,N_1541,N_1660);
nand U2078 (N_2078,N_1558,N_1900);
nand U2079 (N_2079,N_1958,N_1895);
or U2080 (N_2080,N_1942,N_1689);
or U2081 (N_2081,N_1946,N_1935);
nand U2082 (N_2082,N_1990,N_1921);
and U2083 (N_2083,N_1920,N_1917);
or U2084 (N_2084,N_1658,N_1555);
nor U2085 (N_2085,N_1634,N_1835);
nand U2086 (N_2086,N_1701,N_1625);
nor U2087 (N_2087,N_1890,N_1754);
nor U2088 (N_2088,N_1697,N_1818);
or U2089 (N_2089,N_1811,N_1612);
nor U2090 (N_2090,N_1624,N_1995);
nor U2091 (N_2091,N_1945,N_1566);
nor U2092 (N_2092,N_1586,N_1709);
and U2093 (N_2093,N_1557,N_1896);
nand U2094 (N_2094,N_1556,N_1603);
nor U2095 (N_2095,N_1686,N_1733);
and U2096 (N_2096,N_1982,N_1800);
nor U2097 (N_2097,N_1744,N_1859);
nor U2098 (N_2098,N_1638,N_1837);
nor U2099 (N_2099,N_1977,N_1739);
and U2100 (N_2100,N_1949,N_1609);
or U2101 (N_2101,N_1667,N_1749);
nand U2102 (N_2102,N_1814,N_1892);
and U2103 (N_2103,N_1743,N_1633);
nor U2104 (N_2104,N_1817,N_1602);
nand U2105 (N_2105,N_1850,N_1983);
and U2106 (N_2106,N_1950,N_1998);
and U2107 (N_2107,N_1569,N_1528);
nor U2108 (N_2108,N_1844,N_1550);
nor U2109 (N_2109,N_1758,N_1897);
and U2110 (N_2110,N_1926,N_1806);
nor U2111 (N_2111,N_1996,N_1719);
nor U2112 (N_2112,N_1659,N_1590);
nand U2113 (N_2113,N_1849,N_1974);
or U2114 (N_2114,N_1584,N_1899);
or U2115 (N_2115,N_1598,N_1690);
and U2116 (N_2116,N_1628,N_1635);
nor U2117 (N_2117,N_1516,N_1510);
and U2118 (N_2118,N_1875,N_1549);
and U2119 (N_2119,N_1769,N_1619);
nand U2120 (N_2120,N_1504,N_1526);
or U2121 (N_2121,N_1675,N_1514);
and U2122 (N_2122,N_1862,N_1901);
or U2123 (N_2123,N_1962,N_1688);
and U2124 (N_2124,N_1573,N_1554);
nor U2125 (N_2125,N_1668,N_1631);
nor U2126 (N_2126,N_1721,N_1836);
or U2127 (N_2127,N_1637,N_1929);
nand U2128 (N_2128,N_1538,N_1927);
nor U2129 (N_2129,N_1672,N_1611);
and U2130 (N_2130,N_1613,N_1924);
or U2131 (N_2131,N_1574,N_1723);
nor U2132 (N_2132,N_1706,N_1718);
nor U2133 (N_2133,N_1851,N_1801);
nand U2134 (N_2134,N_1525,N_1687);
or U2135 (N_2135,N_1630,N_1883);
or U2136 (N_2136,N_1674,N_1881);
nor U2137 (N_2137,N_1583,N_1702);
or U2138 (N_2138,N_1961,N_1722);
nand U2139 (N_2139,N_1923,N_1766);
nor U2140 (N_2140,N_1632,N_1804);
xor U2141 (N_2141,N_1975,N_1941);
or U2142 (N_2142,N_1575,N_1756);
nand U2143 (N_2143,N_1717,N_1772);
or U2144 (N_2144,N_1861,N_1715);
nand U2145 (N_2145,N_1647,N_1693);
or U2146 (N_2146,N_1994,N_1963);
xor U2147 (N_2147,N_1822,N_1959);
or U2148 (N_2148,N_1565,N_1751);
and U2149 (N_2149,N_1694,N_1740);
nor U2150 (N_2150,N_1727,N_1765);
and U2151 (N_2151,N_1676,N_1588);
or U2152 (N_2152,N_1816,N_1502);
and U2153 (N_2153,N_1615,N_1829);
and U2154 (N_2154,N_1955,N_1691);
nor U2155 (N_2155,N_1730,N_1616);
nand U2156 (N_2156,N_1552,N_1838);
and U2157 (N_2157,N_1511,N_1777);
or U2158 (N_2158,N_1545,N_1606);
nand U2159 (N_2159,N_1741,N_1997);
nor U2160 (N_2160,N_1731,N_1679);
or U2161 (N_2161,N_1534,N_1563);
or U2162 (N_2162,N_1543,N_1582);
nand U2163 (N_2163,N_1776,N_1779);
and U2164 (N_2164,N_1795,N_1669);
or U2165 (N_2165,N_1585,N_1734);
nand U2166 (N_2166,N_1710,N_1579);
nor U2167 (N_2167,N_1939,N_1783);
nor U2168 (N_2168,N_1692,N_1839);
or U2169 (N_2169,N_1914,N_1789);
and U2170 (N_2170,N_1943,N_1601);
nand U2171 (N_2171,N_1627,N_1716);
nand U2172 (N_2172,N_1663,N_1629);
and U2173 (N_2173,N_1771,N_1876);
nand U2174 (N_2174,N_1792,N_1842);
nor U2175 (N_2175,N_1951,N_1735);
xor U2176 (N_2176,N_1547,N_1564);
nand U2177 (N_2177,N_1797,N_1648);
and U2178 (N_2178,N_1909,N_1845);
nor U2179 (N_2179,N_1546,N_1561);
and U2180 (N_2180,N_1869,N_1971);
or U2181 (N_2181,N_1696,N_1807);
and U2182 (N_2182,N_1840,N_1913);
or U2183 (N_2183,N_1855,N_1508);
nor U2184 (N_2184,N_1788,N_1863);
and U2185 (N_2185,N_1832,N_1979);
and U2186 (N_2186,N_1501,N_1764);
nand U2187 (N_2187,N_1646,N_1993);
nand U2188 (N_2188,N_1542,N_1657);
or U2189 (N_2189,N_1506,N_1906);
and U2190 (N_2190,N_1517,N_1572);
nand U2191 (N_2191,N_1824,N_1587);
and U2192 (N_2192,N_1870,N_1618);
and U2193 (N_2193,N_1786,N_1535);
nor U2194 (N_2194,N_1581,N_1656);
nor U2195 (N_2195,N_1747,N_1591);
or U2196 (N_2196,N_1978,N_1887);
nand U2197 (N_2197,N_1708,N_1768);
and U2198 (N_2198,N_1724,N_1570);
and U2199 (N_2199,N_1763,N_1767);
nor U2200 (N_2200,N_1907,N_1605);
or U2201 (N_2201,N_1608,N_1852);
nand U2202 (N_2202,N_1915,N_1539);
and U2203 (N_2203,N_1809,N_1831);
or U2204 (N_2204,N_1893,N_1641);
nand U2205 (N_2205,N_1614,N_1607);
and U2206 (N_2206,N_1642,N_1937);
nor U2207 (N_2207,N_1562,N_1815);
or U2208 (N_2208,N_1932,N_1738);
and U2209 (N_2209,N_1553,N_1970);
or U2210 (N_2210,N_1576,N_1882);
nand U2211 (N_2211,N_1782,N_1621);
nand U2212 (N_2212,N_1793,N_1529);
nand U2213 (N_2213,N_1805,N_1799);
nand U2214 (N_2214,N_1705,N_1567);
and U2215 (N_2215,N_1938,N_1725);
nand U2216 (N_2216,N_1871,N_1860);
or U2217 (N_2217,N_1872,N_1748);
nand U2218 (N_2218,N_1846,N_1678);
nor U2219 (N_2219,N_1984,N_1729);
or U2220 (N_2220,N_1636,N_1784);
and U2221 (N_2221,N_1685,N_1524);
nor U2222 (N_2222,N_1794,N_1969);
and U2223 (N_2223,N_1810,N_1512);
and U2224 (N_2224,N_1808,N_1750);
nor U2225 (N_2225,N_1964,N_1966);
or U2226 (N_2226,N_1544,N_1507);
nand U2227 (N_2227,N_1848,N_1703);
nor U2228 (N_2228,N_1965,N_1513);
nor U2229 (N_2229,N_1987,N_1643);
nor U2230 (N_2230,N_1802,N_1596);
nand U2231 (N_2231,N_1503,N_1644);
or U2232 (N_2232,N_1500,N_1592);
nor U2233 (N_2233,N_1594,N_1898);
nand U2234 (N_2234,N_1505,N_1728);
nor U2235 (N_2235,N_1833,N_1695);
nor U2236 (N_2236,N_1960,N_1912);
nor U2237 (N_2237,N_1661,N_1911);
or U2238 (N_2238,N_1991,N_1755);
or U2239 (N_2239,N_1532,N_1880);
nor U2240 (N_2240,N_1981,N_1677);
nor U2241 (N_2241,N_1530,N_1867);
and U2242 (N_2242,N_1947,N_1666);
nor U2243 (N_2243,N_1858,N_1868);
nand U2244 (N_2244,N_1827,N_1580);
and U2245 (N_2245,N_1834,N_1736);
nor U2246 (N_2246,N_1916,N_1684);
nor U2247 (N_2247,N_1654,N_1548);
and U2248 (N_2248,N_1956,N_1537);
nand U2249 (N_2249,N_1577,N_1877);
nor U2250 (N_2250,N_1782,N_1775);
nor U2251 (N_2251,N_1993,N_1847);
nand U2252 (N_2252,N_1880,N_1663);
nor U2253 (N_2253,N_1946,N_1688);
or U2254 (N_2254,N_1894,N_1574);
nor U2255 (N_2255,N_1795,N_1638);
or U2256 (N_2256,N_1723,N_1581);
and U2257 (N_2257,N_1893,N_1923);
and U2258 (N_2258,N_1709,N_1890);
or U2259 (N_2259,N_1757,N_1872);
nor U2260 (N_2260,N_1943,N_1537);
or U2261 (N_2261,N_1609,N_1698);
xor U2262 (N_2262,N_1867,N_1678);
or U2263 (N_2263,N_1767,N_1799);
nor U2264 (N_2264,N_1657,N_1611);
or U2265 (N_2265,N_1702,N_1869);
nor U2266 (N_2266,N_1738,N_1612);
nand U2267 (N_2267,N_1764,N_1549);
and U2268 (N_2268,N_1546,N_1629);
nor U2269 (N_2269,N_1802,N_1853);
nand U2270 (N_2270,N_1796,N_1802);
and U2271 (N_2271,N_1832,N_1563);
nor U2272 (N_2272,N_1942,N_1996);
nand U2273 (N_2273,N_1536,N_1933);
nand U2274 (N_2274,N_1784,N_1660);
nand U2275 (N_2275,N_1547,N_1520);
nor U2276 (N_2276,N_1993,N_1578);
and U2277 (N_2277,N_1577,N_1740);
and U2278 (N_2278,N_1570,N_1878);
nand U2279 (N_2279,N_1779,N_1636);
or U2280 (N_2280,N_1662,N_1576);
or U2281 (N_2281,N_1570,N_1587);
nor U2282 (N_2282,N_1931,N_1818);
nor U2283 (N_2283,N_1839,N_1667);
nor U2284 (N_2284,N_1728,N_1787);
nand U2285 (N_2285,N_1512,N_1720);
nor U2286 (N_2286,N_1802,N_1911);
nor U2287 (N_2287,N_1644,N_1550);
xnor U2288 (N_2288,N_1699,N_1823);
or U2289 (N_2289,N_1823,N_1738);
and U2290 (N_2290,N_1964,N_1890);
and U2291 (N_2291,N_1786,N_1544);
nor U2292 (N_2292,N_1510,N_1739);
and U2293 (N_2293,N_1580,N_1607);
and U2294 (N_2294,N_1910,N_1635);
or U2295 (N_2295,N_1848,N_1828);
nor U2296 (N_2296,N_1857,N_1839);
xnor U2297 (N_2297,N_1588,N_1977);
or U2298 (N_2298,N_1927,N_1884);
or U2299 (N_2299,N_1965,N_1992);
and U2300 (N_2300,N_1539,N_1788);
and U2301 (N_2301,N_1906,N_1867);
nand U2302 (N_2302,N_1607,N_1501);
nand U2303 (N_2303,N_1668,N_1698);
nand U2304 (N_2304,N_1736,N_1550);
or U2305 (N_2305,N_1824,N_1787);
nand U2306 (N_2306,N_1602,N_1760);
nor U2307 (N_2307,N_1969,N_1789);
nor U2308 (N_2308,N_1552,N_1726);
nor U2309 (N_2309,N_1662,N_1630);
nor U2310 (N_2310,N_1627,N_1903);
nor U2311 (N_2311,N_1902,N_1832);
and U2312 (N_2312,N_1872,N_1587);
and U2313 (N_2313,N_1806,N_1959);
nor U2314 (N_2314,N_1532,N_1839);
or U2315 (N_2315,N_1750,N_1670);
nand U2316 (N_2316,N_1774,N_1887);
and U2317 (N_2317,N_1899,N_1628);
or U2318 (N_2318,N_1613,N_1861);
and U2319 (N_2319,N_1671,N_1782);
nor U2320 (N_2320,N_1572,N_1575);
nand U2321 (N_2321,N_1652,N_1807);
nand U2322 (N_2322,N_1891,N_1834);
and U2323 (N_2323,N_1943,N_1552);
nand U2324 (N_2324,N_1704,N_1594);
or U2325 (N_2325,N_1557,N_1586);
nor U2326 (N_2326,N_1585,N_1861);
or U2327 (N_2327,N_1914,N_1941);
nor U2328 (N_2328,N_1744,N_1645);
or U2329 (N_2329,N_1665,N_1936);
nor U2330 (N_2330,N_1696,N_1888);
or U2331 (N_2331,N_1524,N_1545);
and U2332 (N_2332,N_1854,N_1818);
and U2333 (N_2333,N_1828,N_1750);
nor U2334 (N_2334,N_1929,N_1571);
or U2335 (N_2335,N_1529,N_1718);
nor U2336 (N_2336,N_1518,N_1502);
and U2337 (N_2337,N_1886,N_1642);
nor U2338 (N_2338,N_1974,N_1791);
and U2339 (N_2339,N_1522,N_1662);
and U2340 (N_2340,N_1784,N_1863);
or U2341 (N_2341,N_1816,N_1989);
or U2342 (N_2342,N_1507,N_1888);
nand U2343 (N_2343,N_1568,N_1795);
and U2344 (N_2344,N_1624,N_1595);
or U2345 (N_2345,N_1640,N_1777);
and U2346 (N_2346,N_1778,N_1782);
or U2347 (N_2347,N_1656,N_1851);
nand U2348 (N_2348,N_1894,N_1909);
nand U2349 (N_2349,N_1685,N_1831);
nand U2350 (N_2350,N_1569,N_1671);
nand U2351 (N_2351,N_1690,N_1672);
and U2352 (N_2352,N_1723,N_1673);
nand U2353 (N_2353,N_1653,N_1876);
nor U2354 (N_2354,N_1879,N_1872);
or U2355 (N_2355,N_1851,N_1709);
or U2356 (N_2356,N_1624,N_1832);
or U2357 (N_2357,N_1721,N_1587);
and U2358 (N_2358,N_1639,N_1884);
or U2359 (N_2359,N_1593,N_1801);
nor U2360 (N_2360,N_1564,N_1599);
nand U2361 (N_2361,N_1777,N_1842);
nor U2362 (N_2362,N_1851,N_1692);
or U2363 (N_2363,N_1743,N_1506);
or U2364 (N_2364,N_1623,N_1918);
nor U2365 (N_2365,N_1624,N_1777);
and U2366 (N_2366,N_1888,N_1677);
nand U2367 (N_2367,N_1994,N_1630);
nor U2368 (N_2368,N_1651,N_1691);
nor U2369 (N_2369,N_1731,N_1874);
xnor U2370 (N_2370,N_1556,N_1748);
nor U2371 (N_2371,N_1657,N_1710);
and U2372 (N_2372,N_1988,N_1953);
nor U2373 (N_2373,N_1664,N_1668);
nand U2374 (N_2374,N_1664,N_1555);
or U2375 (N_2375,N_1987,N_1762);
and U2376 (N_2376,N_1942,N_1855);
nor U2377 (N_2377,N_1729,N_1540);
and U2378 (N_2378,N_1609,N_1738);
and U2379 (N_2379,N_1975,N_1797);
or U2380 (N_2380,N_1627,N_1915);
nand U2381 (N_2381,N_1696,N_1855);
nor U2382 (N_2382,N_1766,N_1961);
nand U2383 (N_2383,N_1626,N_1761);
or U2384 (N_2384,N_1887,N_1537);
or U2385 (N_2385,N_1803,N_1564);
nor U2386 (N_2386,N_1523,N_1767);
and U2387 (N_2387,N_1720,N_1655);
nor U2388 (N_2388,N_1558,N_1922);
nor U2389 (N_2389,N_1987,N_1603);
nand U2390 (N_2390,N_1639,N_1974);
and U2391 (N_2391,N_1873,N_1893);
or U2392 (N_2392,N_1876,N_1669);
and U2393 (N_2393,N_1517,N_1962);
nand U2394 (N_2394,N_1688,N_1698);
or U2395 (N_2395,N_1561,N_1780);
or U2396 (N_2396,N_1509,N_1701);
nand U2397 (N_2397,N_1745,N_1590);
and U2398 (N_2398,N_1512,N_1862);
nand U2399 (N_2399,N_1655,N_1652);
or U2400 (N_2400,N_1533,N_1513);
or U2401 (N_2401,N_1618,N_1521);
and U2402 (N_2402,N_1771,N_1704);
nor U2403 (N_2403,N_1697,N_1620);
nor U2404 (N_2404,N_1966,N_1807);
and U2405 (N_2405,N_1853,N_1617);
or U2406 (N_2406,N_1893,N_1780);
nor U2407 (N_2407,N_1961,N_1868);
nand U2408 (N_2408,N_1742,N_1978);
nand U2409 (N_2409,N_1549,N_1864);
or U2410 (N_2410,N_1666,N_1520);
or U2411 (N_2411,N_1896,N_1689);
nand U2412 (N_2412,N_1747,N_1978);
or U2413 (N_2413,N_1609,N_1747);
xor U2414 (N_2414,N_1872,N_1566);
nand U2415 (N_2415,N_1715,N_1844);
nor U2416 (N_2416,N_1704,N_1524);
and U2417 (N_2417,N_1908,N_1537);
and U2418 (N_2418,N_1863,N_1878);
nand U2419 (N_2419,N_1554,N_1903);
or U2420 (N_2420,N_1913,N_1937);
nand U2421 (N_2421,N_1648,N_1781);
nor U2422 (N_2422,N_1923,N_1715);
nand U2423 (N_2423,N_1717,N_1775);
and U2424 (N_2424,N_1860,N_1789);
or U2425 (N_2425,N_1778,N_1741);
and U2426 (N_2426,N_1999,N_1503);
nor U2427 (N_2427,N_1757,N_1725);
and U2428 (N_2428,N_1705,N_1608);
nor U2429 (N_2429,N_1807,N_1789);
nor U2430 (N_2430,N_1812,N_1818);
and U2431 (N_2431,N_1741,N_1797);
and U2432 (N_2432,N_1540,N_1538);
nand U2433 (N_2433,N_1775,N_1542);
and U2434 (N_2434,N_1675,N_1821);
or U2435 (N_2435,N_1567,N_1831);
nor U2436 (N_2436,N_1512,N_1504);
nor U2437 (N_2437,N_1627,N_1992);
nor U2438 (N_2438,N_1746,N_1872);
nor U2439 (N_2439,N_1962,N_1839);
and U2440 (N_2440,N_1860,N_1821);
and U2441 (N_2441,N_1835,N_1880);
or U2442 (N_2442,N_1864,N_1550);
and U2443 (N_2443,N_1829,N_1876);
nor U2444 (N_2444,N_1676,N_1923);
nand U2445 (N_2445,N_1535,N_1716);
and U2446 (N_2446,N_1570,N_1508);
and U2447 (N_2447,N_1628,N_1812);
or U2448 (N_2448,N_1917,N_1604);
or U2449 (N_2449,N_1967,N_1950);
xor U2450 (N_2450,N_1825,N_1562);
nor U2451 (N_2451,N_1658,N_1770);
and U2452 (N_2452,N_1666,N_1567);
and U2453 (N_2453,N_1768,N_1973);
nand U2454 (N_2454,N_1887,N_1516);
or U2455 (N_2455,N_1758,N_1836);
and U2456 (N_2456,N_1799,N_1951);
and U2457 (N_2457,N_1705,N_1699);
or U2458 (N_2458,N_1793,N_1759);
nor U2459 (N_2459,N_1573,N_1964);
or U2460 (N_2460,N_1640,N_1513);
or U2461 (N_2461,N_1830,N_1755);
nor U2462 (N_2462,N_1710,N_1670);
nor U2463 (N_2463,N_1661,N_1999);
nand U2464 (N_2464,N_1538,N_1861);
nand U2465 (N_2465,N_1696,N_1602);
nand U2466 (N_2466,N_1579,N_1759);
nor U2467 (N_2467,N_1617,N_1578);
or U2468 (N_2468,N_1730,N_1922);
nor U2469 (N_2469,N_1545,N_1694);
and U2470 (N_2470,N_1792,N_1752);
or U2471 (N_2471,N_1821,N_1604);
nand U2472 (N_2472,N_1736,N_1620);
nor U2473 (N_2473,N_1869,N_1587);
or U2474 (N_2474,N_1738,N_1905);
or U2475 (N_2475,N_1527,N_1582);
nor U2476 (N_2476,N_1965,N_1735);
nor U2477 (N_2477,N_1777,N_1516);
or U2478 (N_2478,N_1512,N_1861);
and U2479 (N_2479,N_1935,N_1692);
nand U2480 (N_2480,N_1627,N_1991);
and U2481 (N_2481,N_1872,N_1548);
and U2482 (N_2482,N_1535,N_1809);
nand U2483 (N_2483,N_1578,N_1606);
nand U2484 (N_2484,N_1651,N_1654);
or U2485 (N_2485,N_1856,N_1705);
and U2486 (N_2486,N_1589,N_1906);
and U2487 (N_2487,N_1730,N_1761);
and U2488 (N_2488,N_1824,N_1949);
and U2489 (N_2489,N_1616,N_1506);
nor U2490 (N_2490,N_1550,N_1509);
nand U2491 (N_2491,N_1867,N_1557);
or U2492 (N_2492,N_1807,N_1685);
and U2493 (N_2493,N_1615,N_1694);
and U2494 (N_2494,N_1728,N_1887);
nand U2495 (N_2495,N_1672,N_1958);
and U2496 (N_2496,N_1720,N_1617);
nand U2497 (N_2497,N_1813,N_1782);
xnor U2498 (N_2498,N_1785,N_1745);
or U2499 (N_2499,N_1617,N_1545);
and U2500 (N_2500,N_2331,N_2190);
or U2501 (N_2501,N_2090,N_2189);
nand U2502 (N_2502,N_2218,N_2269);
or U2503 (N_2503,N_2290,N_2182);
nor U2504 (N_2504,N_2326,N_2068);
and U2505 (N_2505,N_2052,N_2373);
or U2506 (N_2506,N_2493,N_2003);
and U2507 (N_2507,N_2295,N_2399);
nand U2508 (N_2508,N_2154,N_2332);
or U2509 (N_2509,N_2431,N_2359);
nor U2510 (N_2510,N_2026,N_2265);
and U2511 (N_2511,N_2004,N_2042);
and U2512 (N_2512,N_2089,N_2352);
or U2513 (N_2513,N_2279,N_2071);
nand U2514 (N_2514,N_2175,N_2039);
nor U2515 (N_2515,N_2215,N_2479);
or U2516 (N_2516,N_2064,N_2210);
or U2517 (N_2517,N_2448,N_2402);
or U2518 (N_2518,N_2292,N_2214);
nor U2519 (N_2519,N_2081,N_2335);
or U2520 (N_2520,N_2405,N_2488);
or U2521 (N_2521,N_2296,N_2418);
nand U2522 (N_2522,N_2145,N_2456);
nor U2523 (N_2523,N_2103,N_2420);
nand U2524 (N_2524,N_2419,N_2391);
nand U2525 (N_2525,N_2112,N_2208);
and U2526 (N_2526,N_2494,N_2077);
and U2527 (N_2527,N_2166,N_2370);
nor U2528 (N_2528,N_2430,N_2375);
and U2529 (N_2529,N_2293,N_2165);
nor U2530 (N_2530,N_2246,N_2294);
or U2531 (N_2531,N_2378,N_2065);
and U2532 (N_2532,N_2091,N_2106);
nand U2533 (N_2533,N_2137,N_2180);
nand U2534 (N_2534,N_2357,N_2084);
nand U2535 (N_2535,N_2327,N_2118);
xnor U2536 (N_2536,N_2035,N_2440);
nand U2537 (N_2537,N_2238,N_2413);
and U2538 (N_2538,N_2219,N_2186);
and U2539 (N_2539,N_2450,N_2049);
or U2540 (N_2540,N_2025,N_2453);
and U2541 (N_2541,N_2364,N_2038);
nor U2542 (N_2542,N_2342,N_2428);
nand U2543 (N_2543,N_2429,N_2369);
nand U2544 (N_2544,N_2347,N_2385);
or U2545 (N_2545,N_2462,N_2015);
nor U2546 (N_2546,N_2236,N_2099);
and U2547 (N_2547,N_2427,N_2047);
or U2548 (N_2548,N_2325,N_2121);
nor U2549 (N_2549,N_2339,N_2177);
nor U2550 (N_2550,N_2132,N_2277);
nor U2551 (N_2551,N_2232,N_2379);
or U2552 (N_2552,N_2034,N_2128);
nor U2553 (N_2553,N_2388,N_2434);
or U2554 (N_2554,N_2080,N_2008);
nor U2555 (N_2555,N_2123,N_2174);
or U2556 (N_2556,N_2437,N_2032);
nand U2557 (N_2557,N_2408,N_2087);
and U2558 (N_2558,N_2260,N_2486);
nand U2559 (N_2559,N_2116,N_2130);
nor U2560 (N_2560,N_2253,N_2381);
and U2561 (N_2561,N_2017,N_2110);
or U2562 (N_2562,N_2005,N_2138);
and U2563 (N_2563,N_2351,N_2368);
nand U2564 (N_2564,N_2241,N_2348);
nor U2565 (N_2565,N_2029,N_2200);
nor U2566 (N_2566,N_2308,N_2247);
nor U2567 (N_2567,N_2148,N_2129);
and U2568 (N_2568,N_2316,N_2484);
nor U2569 (N_2569,N_2044,N_2157);
nor U2570 (N_2570,N_2237,N_2257);
nor U2571 (N_2571,N_2187,N_2449);
nor U2572 (N_2572,N_2113,N_2060);
nor U2573 (N_2573,N_2036,N_2027);
nand U2574 (N_2574,N_2248,N_2377);
and U2575 (N_2575,N_2171,N_2014);
nand U2576 (N_2576,N_2161,N_2389);
nor U2577 (N_2577,N_2336,N_2487);
or U2578 (N_2578,N_2376,N_2019);
nor U2579 (N_2579,N_2082,N_2196);
or U2580 (N_2580,N_2392,N_2315);
nor U2581 (N_2581,N_2333,N_2345);
nor U2582 (N_2582,N_2184,N_2134);
nor U2583 (N_2583,N_2188,N_2202);
or U2584 (N_2584,N_2023,N_2105);
nor U2585 (N_2585,N_2270,N_2020);
nand U2586 (N_2586,N_2122,N_2466);
and U2587 (N_2587,N_2281,N_2193);
nor U2588 (N_2588,N_2021,N_2255);
nor U2589 (N_2589,N_2299,N_2474);
or U2590 (N_2590,N_2282,N_2362);
or U2591 (N_2591,N_2179,N_2258);
nor U2592 (N_2592,N_2421,N_2114);
and U2593 (N_2593,N_2322,N_2457);
nand U2594 (N_2594,N_2176,N_2168);
nor U2595 (N_2595,N_2300,N_2483);
or U2596 (N_2596,N_2143,N_2152);
nor U2597 (N_2597,N_2076,N_2056);
and U2598 (N_2598,N_2229,N_2334);
nand U2599 (N_2599,N_2464,N_2473);
nor U2600 (N_2600,N_2183,N_2367);
nor U2601 (N_2601,N_2226,N_2201);
nor U2602 (N_2602,N_2040,N_2446);
and U2603 (N_2603,N_2463,N_2140);
or U2604 (N_2604,N_2412,N_2361);
nor U2605 (N_2605,N_2301,N_2169);
nand U2606 (N_2606,N_2059,N_2415);
and U2607 (N_2607,N_2268,N_2010);
nand U2608 (N_2608,N_2360,N_2289);
nor U2609 (N_2609,N_2125,N_2149);
nor U2610 (N_2610,N_2062,N_2498);
nand U2611 (N_2611,N_2163,N_2382);
or U2612 (N_2612,N_2425,N_2136);
nor U2613 (N_2613,N_2120,N_2205);
nor U2614 (N_2614,N_2374,N_2459);
nor U2615 (N_2615,N_2309,N_2314);
and U2616 (N_2616,N_2159,N_2101);
or U2617 (N_2617,N_2452,N_2444);
nand U2618 (N_2618,N_2400,N_2403);
nand U2619 (N_2619,N_2297,N_2432);
nor U2620 (N_2620,N_2324,N_2079);
nand U2621 (N_2621,N_2280,N_2424);
and U2622 (N_2622,N_2371,N_2051);
nand U2623 (N_2623,N_2073,N_2461);
nor U2624 (N_2624,N_2050,N_2227);
or U2625 (N_2625,N_2206,N_2115);
and U2626 (N_2626,N_2490,N_2097);
and U2627 (N_2627,N_2330,N_2303);
nand U2628 (N_2628,N_2013,N_2234);
or U2629 (N_2629,N_2111,N_2022);
nand U2630 (N_2630,N_2133,N_2158);
nor U2631 (N_2631,N_2142,N_2287);
nand U2632 (N_2632,N_2102,N_2222);
nor U2633 (N_2633,N_2144,N_2497);
nand U2634 (N_2634,N_2092,N_2191);
and U2635 (N_2635,N_2313,N_2061);
or U2636 (N_2636,N_2235,N_2319);
and U2637 (N_2637,N_2387,N_2066);
and U2638 (N_2638,N_2249,N_2285);
nand U2639 (N_2639,N_2291,N_2024);
or U2640 (N_2640,N_2283,N_2386);
or U2641 (N_2641,N_2485,N_2489);
and U2642 (N_2642,N_2383,N_2096);
nor U2643 (N_2643,N_2100,N_2471);
or U2644 (N_2644,N_2094,N_2016);
nand U2645 (N_2645,N_2470,N_2476);
nand U2646 (N_2646,N_2178,N_2302);
or U2647 (N_2647,N_2317,N_2212);
nor U2648 (N_2648,N_2477,N_2321);
nand U2649 (N_2649,N_2438,N_2088);
and U2650 (N_2650,N_2414,N_2467);
and U2651 (N_2651,N_2160,N_2233);
nor U2652 (N_2652,N_2328,N_2455);
nand U2653 (N_2653,N_2155,N_2354);
and U2654 (N_2654,N_2454,N_2213);
and U2655 (N_2655,N_2240,N_2496);
and U2656 (N_2656,N_2198,N_2181);
and U2657 (N_2657,N_2480,N_2119);
nand U2658 (N_2658,N_2482,N_2220);
nor U2659 (N_2659,N_2349,N_2284);
and U2660 (N_2660,N_2054,N_2443);
nor U2661 (N_2661,N_2264,N_2243);
and U2662 (N_2662,N_2346,N_2447);
nand U2663 (N_2663,N_2093,N_2266);
nand U2664 (N_2664,N_2272,N_2104);
and U2665 (N_2665,N_2107,N_2069);
and U2666 (N_2666,N_2338,N_2156);
and U2667 (N_2667,N_2078,N_2007);
or U2668 (N_2668,N_2209,N_2343);
or U2669 (N_2669,N_2067,N_2397);
and U2670 (N_2670,N_2204,N_2126);
nand U2671 (N_2671,N_2310,N_2495);
and U2672 (N_2672,N_2095,N_2288);
nand U2673 (N_2673,N_2207,N_2472);
nor U2674 (N_2674,N_2468,N_2410);
nor U2675 (N_2675,N_2251,N_2394);
or U2676 (N_2676,N_2195,N_2363);
or U2677 (N_2677,N_2341,N_2002);
and U2678 (N_2678,N_2398,N_2147);
and U2679 (N_2679,N_2478,N_2409);
nand U2680 (N_2680,N_2075,N_2298);
or U2681 (N_2681,N_2304,N_2018);
and U2682 (N_2682,N_2221,N_2278);
and U2683 (N_2683,N_2305,N_2262);
xor U2684 (N_2684,N_2380,N_2372);
and U2685 (N_2685,N_2491,N_2337);
nand U2686 (N_2686,N_2000,N_2009);
nand U2687 (N_2687,N_2416,N_2217);
nor U2688 (N_2688,N_2250,N_2261);
and U2689 (N_2689,N_2417,N_2030);
nor U2690 (N_2690,N_2194,N_2216);
nand U2691 (N_2691,N_2242,N_2329);
nand U2692 (N_2692,N_2146,N_2366);
or U2693 (N_2693,N_2117,N_2012);
or U2694 (N_2694,N_2072,N_2451);
nor U2695 (N_2695,N_2344,N_2445);
nand U2696 (N_2696,N_2046,N_2393);
nor U2697 (N_2697,N_2436,N_2127);
or U2698 (N_2698,N_2475,N_2435);
nand U2699 (N_2699,N_2224,N_2230);
nand U2700 (N_2700,N_2108,N_2340);
or U2701 (N_2701,N_2172,N_2252);
nor U2702 (N_2702,N_2263,N_2001);
nand U2703 (N_2703,N_2307,N_2271);
or U2704 (N_2704,N_2053,N_2273);
nand U2705 (N_2705,N_2254,N_2124);
or U2706 (N_2706,N_2406,N_2031);
or U2707 (N_2707,N_2070,N_2048);
and U2708 (N_2708,N_2384,N_2197);
nor U2709 (N_2709,N_2028,N_2063);
nand U2710 (N_2710,N_2286,N_2225);
or U2711 (N_2711,N_2150,N_2492);
or U2712 (N_2712,N_2481,N_2074);
nand U2713 (N_2713,N_2083,N_2356);
nand U2714 (N_2714,N_2045,N_2086);
nand U2715 (N_2715,N_2469,N_2037);
or U2716 (N_2716,N_2244,N_2320);
nand U2717 (N_2717,N_2433,N_2422);
and U2718 (N_2718,N_2256,N_2401);
or U2719 (N_2719,N_2259,N_2426);
and U2720 (N_2720,N_2276,N_2312);
nor U2721 (N_2721,N_2306,N_2223);
nor U2722 (N_2722,N_2318,N_2006);
or U2723 (N_2723,N_2211,N_2239);
nand U2724 (N_2724,N_2442,N_2173);
nand U2725 (N_2725,N_2267,N_2058);
and U2726 (N_2726,N_2323,N_2085);
or U2727 (N_2727,N_2404,N_2228);
nor U2728 (N_2728,N_2043,N_2274);
nand U2729 (N_2729,N_2131,N_2139);
or U2730 (N_2730,N_2353,N_2041);
and U2731 (N_2731,N_2055,N_2411);
and U2732 (N_2732,N_2231,N_2151);
nand U2733 (N_2733,N_2396,N_2109);
nand U2734 (N_2734,N_2458,N_2439);
or U2735 (N_2735,N_2275,N_2098);
nand U2736 (N_2736,N_2167,N_2162);
nand U2737 (N_2737,N_2057,N_2407);
or U2738 (N_2738,N_2170,N_2365);
nor U2739 (N_2739,N_2460,N_2355);
or U2740 (N_2740,N_2199,N_2164);
or U2741 (N_2741,N_2311,N_2358);
or U2742 (N_2742,N_2441,N_2390);
nand U2743 (N_2743,N_2245,N_2423);
nand U2744 (N_2744,N_2350,N_2141);
or U2745 (N_2745,N_2395,N_2011);
nor U2746 (N_2746,N_2192,N_2135);
nor U2747 (N_2747,N_2185,N_2203);
nand U2748 (N_2748,N_2033,N_2499);
nand U2749 (N_2749,N_2465,N_2153);
or U2750 (N_2750,N_2337,N_2130);
or U2751 (N_2751,N_2353,N_2031);
and U2752 (N_2752,N_2295,N_2282);
or U2753 (N_2753,N_2421,N_2115);
or U2754 (N_2754,N_2262,N_2076);
nand U2755 (N_2755,N_2185,N_2186);
and U2756 (N_2756,N_2417,N_2134);
nor U2757 (N_2757,N_2464,N_2360);
nand U2758 (N_2758,N_2002,N_2247);
or U2759 (N_2759,N_2324,N_2366);
and U2760 (N_2760,N_2186,N_2253);
nand U2761 (N_2761,N_2182,N_2378);
nor U2762 (N_2762,N_2078,N_2272);
or U2763 (N_2763,N_2166,N_2269);
or U2764 (N_2764,N_2405,N_2071);
and U2765 (N_2765,N_2073,N_2315);
nand U2766 (N_2766,N_2414,N_2146);
nor U2767 (N_2767,N_2052,N_2097);
nand U2768 (N_2768,N_2301,N_2455);
nand U2769 (N_2769,N_2157,N_2416);
and U2770 (N_2770,N_2409,N_2109);
nor U2771 (N_2771,N_2301,N_2044);
or U2772 (N_2772,N_2256,N_2104);
or U2773 (N_2773,N_2343,N_2400);
and U2774 (N_2774,N_2095,N_2442);
or U2775 (N_2775,N_2220,N_2213);
nand U2776 (N_2776,N_2199,N_2291);
nand U2777 (N_2777,N_2132,N_2092);
or U2778 (N_2778,N_2401,N_2371);
nand U2779 (N_2779,N_2190,N_2363);
nand U2780 (N_2780,N_2415,N_2399);
nor U2781 (N_2781,N_2146,N_2173);
nand U2782 (N_2782,N_2435,N_2169);
nand U2783 (N_2783,N_2064,N_2251);
and U2784 (N_2784,N_2023,N_2329);
and U2785 (N_2785,N_2045,N_2423);
nand U2786 (N_2786,N_2132,N_2065);
and U2787 (N_2787,N_2092,N_2356);
or U2788 (N_2788,N_2025,N_2140);
nand U2789 (N_2789,N_2241,N_2131);
or U2790 (N_2790,N_2081,N_2133);
or U2791 (N_2791,N_2032,N_2078);
and U2792 (N_2792,N_2084,N_2052);
nand U2793 (N_2793,N_2304,N_2464);
nor U2794 (N_2794,N_2471,N_2491);
xor U2795 (N_2795,N_2306,N_2059);
or U2796 (N_2796,N_2083,N_2345);
nand U2797 (N_2797,N_2343,N_2361);
or U2798 (N_2798,N_2183,N_2303);
and U2799 (N_2799,N_2220,N_2230);
nor U2800 (N_2800,N_2455,N_2207);
nor U2801 (N_2801,N_2400,N_2182);
or U2802 (N_2802,N_2352,N_2024);
nor U2803 (N_2803,N_2456,N_2283);
nor U2804 (N_2804,N_2125,N_2025);
or U2805 (N_2805,N_2305,N_2265);
and U2806 (N_2806,N_2338,N_2086);
and U2807 (N_2807,N_2393,N_2097);
and U2808 (N_2808,N_2265,N_2378);
nand U2809 (N_2809,N_2182,N_2175);
or U2810 (N_2810,N_2002,N_2286);
and U2811 (N_2811,N_2264,N_2248);
or U2812 (N_2812,N_2470,N_2010);
nor U2813 (N_2813,N_2266,N_2062);
nor U2814 (N_2814,N_2126,N_2211);
or U2815 (N_2815,N_2047,N_2480);
or U2816 (N_2816,N_2206,N_2329);
and U2817 (N_2817,N_2094,N_2374);
or U2818 (N_2818,N_2294,N_2330);
nand U2819 (N_2819,N_2348,N_2248);
or U2820 (N_2820,N_2374,N_2008);
or U2821 (N_2821,N_2038,N_2188);
or U2822 (N_2822,N_2474,N_2473);
and U2823 (N_2823,N_2387,N_2366);
nand U2824 (N_2824,N_2270,N_2097);
and U2825 (N_2825,N_2277,N_2141);
and U2826 (N_2826,N_2039,N_2280);
nor U2827 (N_2827,N_2040,N_2281);
nor U2828 (N_2828,N_2006,N_2444);
nor U2829 (N_2829,N_2250,N_2286);
and U2830 (N_2830,N_2472,N_2263);
nand U2831 (N_2831,N_2274,N_2135);
or U2832 (N_2832,N_2163,N_2081);
nor U2833 (N_2833,N_2312,N_2022);
nand U2834 (N_2834,N_2058,N_2005);
nor U2835 (N_2835,N_2447,N_2268);
nor U2836 (N_2836,N_2451,N_2206);
or U2837 (N_2837,N_2287,N_2405);
and U2838 (N_2838,N_2184,N_2279);
nand U2839 (N_2839,N_2125,N_2112);
nor U2840 (N_2840,N_2392,N_2205);
xor U2841 (N_2841,N_2051,N_2132);
nand U2842 (N_2842,N_2167,N_2080);
nor U2843 (N_2843,N_2417,N_2121);
and U2844 (N_2844,N_2059,N_2389);
and U2845 (N_2845,N_2074,N_2060);
nand U2846 (N_2846,N_2075,N_2231);
or U2847 (N_2847,N_2340,N_2317);
or U2848 (N_2848,N_2326,N_2243);
nand U2849 (N_2849,N_2042,N_2008);
or U2850 (N_2850,N_2088,N_2416);
or U2851 (N_2851,N_2494,N_2161);
and U2852 (N_2852,N_2431,N_2314);
or U2853 (N_2853,N_2045,N_2386);
nor U2854 (N_2854,N_2287,N_2409);
and U2855 (N_2855,N_2479,N_2001);
nor U2856 (N_2856,N_2453,N_2402);
or U2857 (N_2857,N_2456,N_2044);
nor U2858 (N_2858,N_2191,N_2225);
nand U2859 (N_2859,N_2290,N_2206);
and U2860 (N_2860,N_2276,N_2179);
or U2861 (N_2861,N_2075,N_2141);
or U2862 (N_2862,N_2242,N_2404);
nand U2863 (N_2863,N_2095,N_2222);
nor U2864 (N_2864,N_2079,N_2199);
and U2865 (N_2865,N_2341,N_2387);
and U2866 (N_2866,N_2199,N_2474);
and U2867 (N_2867,N_2369,N_2216);
nand U2868 (N_2868,N_2176,N_2166);
and U2869 (N_2869,N_2239,N_2149);
nand U2870 (N_2870,N_2107,N_2145);
and U2871 (N_2871,N_2178,N_2217);
or U2872 (N_2872,N_2217,N_2114);
and U2873 (N_2873,N_2429,N_2174);
nor U2874 (N_2874,N_2132,N_2387);
xnor U2875 (N_2875,N_2105,N_2072);
or U2876 (N_2876,N_2450,N_2421);
nor U2877 (N_2877,N_2436,N_2277);
nand U2878 (N_2878,N_2048,N_2141);
nor U2879 (N_2879,N_2124,N_2185);
nor U2880 (N_2880,N_2091,N_2234);
and U2881 (N_2881,N_2339,N_2343);
or U2882 (N_2882,N_2245,N_2110);
and U2883 (N_2883,N_2372,N_2004);
or U2884 (N_2884,N_2153,N_2261);
and U2885 (N_2885,N_2089,N_2282);
nand U2886 (N_2886,N_2082,N_2089);
nor U2887 (N_2887,N_2185,N_2354);
and U2888 (N_2888,N_2352,N_2060);
nor U2889 (N_2889,N_2296,N_2286);
nor U2890 (N_2890,N_2273,N_2401);
nor U2891 (N_2891,N_2049,N_2238);
or U2892 (N_2892,N_2176,N_2015);
and U2893 (N_2893,N_2462,N_2218);
nand U2894 (N_2894,N_2316,N_2446);
or U2895 (N_2895,N_2473,N_2071);
nand U2896 (N_2896,N_2164,N_2171);
and U2897 (N_2897,N_2142,N_2194);
or U2898 (N_2898,N_2025,N_2053);
nor U2899 (N_2899,N_2496,N_2271);
and U2900 (N_2900,N_2365,N_2307);
xnor U2901 (N_2901,N_2075,N_2341);
nor U2902 (N_2902,N_2375,N_2064);
or U2903 (N_2903,N_2407,N_2462);
nand U2904 (N_2904,N_2007,N_2424);
nand U2905 (N_2905,N_2078,N_2476);
or U2906 (N_2906,N_2285,N_2377);
or U2907 (N_2907,N_2349,N_2016);
nor U2908 (N_2908,N_2084,N_2022);
nor U2909 (N_2909,N_2163,N_2013);
and U2910 (N_2910,N_2394,N_2120);
or U2911 (N_2911,N_2292,N_2385);
nand U2912 (N_2912,N_2198,N_2452);
and U2913 (N_2913,N_2220,N_2426);
nand U2914 (N_2914,N_2394,N_2157);
nor U2915 (N_2915,N_2362,N_2492);
nor U2916 (N_2916,N_2483,N_2302);
nor U2917 (N_2917,N_2073,N_2090);
nor U2918 (N_2918,N_2314,N_2359);
nand U2919 (N_2919,N_2153,N_2088);
nand U2920 (N_2920,N_2425,N_2456);
and U2921 (N_2921,N_2163,N_2142);
nor U2922 (N_2922,N_2367,N_2017);
nand U2923 (N_2923,N_2380,N_2012);
nand U2924 (N_2924,N_2479,N_2033);
or U2925 (N_2925,N_2408,N_2376);
or U2926 (N_2926,N_2433,N_2160);
nand U2927 (N_2927,N_2315,N_2367);
or U2928 (N_2928,N_2051,N_2156);
nor U2929 (N_2929,N_2191,N_2342);
and U2930 (N_2930,N_2041,N_2275);
or U2931 (N_2931,N_2153,N_2012);
nor U2932 (N_2932,N_2083,N_2301);
or U2933 (N_2933,N_2029,N_2453);
nand U2934 (N_2934,N_2012,N_2366);
or U2935 (N_2935,N_2046,N_2206);
or U2936 (N_2936,N_2141,N_2158);
or U2937 (N_2937,N_2272,N_2185);
or U2938 (N_2938,N_2313,N_2211);
nand U2939 (N_2939,N_2020,N_2271);
and U2940 (N_2940,N_2260,N_2259);
nand U2941 (N_2941,N_2451,N_2364);
xor U2942 (N_2942,N_2064,N_2438);
nor U2943 (N_2943,N_2049,N_2117);
nand U2944 (N_2944,N_2029,N_2233);
nor U2945 (N_2945,N_2198,N_2389);
or U2946 (N_2946,N_2447,N_2136);
nor U2947 (N_2947,N_2450,N_2041);
nor U2948 (N_2948,N_2175,N_2096);
and U2949 (N_2949,N_2006,N_2217);
or U2950 (N_2950,N_2439,N_2231);
nand U2951 (N_2951,N_2302,N_2313);
nor U2952 (N_2952,N_2311,N_2067);
nor U2953 (N_2953,N_2449,N_2076);
and U2954 (N_2954,N_2207,N_2499);
and U2955 (N_2955,N_2205,N_2356);
nand U2956 (N_2956,N_2271,N_2061);
nand U2957 (N_2957,N_2077,N_2381);
nand U2958 (N_2958,N_2363,N_2127);
and U2959 (N_2959,N_2357,N_2154);
nand U2960 (N_2960,N_2413,N_2470);
nand U2961 (N_2961,N_2222,N_2329);
nand U2962 (N_2962,N_2331,N_2261);
and U2963 (N_2963,N_2279,N_2278);
nor U2964 (N_2964,N_2251,N_2220);
nor U2965 (N_2965,N_2126,N_2468);
or U2966 (N_2966,N_2288,N_2402);
nand U2967 (N_2967,N_2288,N_2015);
and U2968 (N_2968,N_2143,N_2000);
nand U2969 (N_2969,N_2387,N_2419);
or U2970 (N_2970,N_2460,N_2243);
or U2971 (N_2971,N_2474,N_2241);
and U2972 (N_2972,N_2423,N_2490);
nand U2973 (N_2973,N_2248,N_2028);
or U2974 (N_2974,N_2287,N_2114);
nand U2975 (N_2975,N_2009,N_2270);
nand U2976 (N_2976,N_2016,N_2393);
and U2977 (N_2977,N_2148,N_2240);
and U2978 (N_2978,N_2050,N_2318);
nor U2979 (N_2979,N_2479,N_2179);
nand U2980 (N_2980,N_2483,N_2335);
nand U2981 (N_2981,N_2202,N_2351);
nor U2982 (N_2982,N_2469,N_2112);
or U2983 (N_2983,N_2263,N_2485);
or U2984 (N_2984,N_2300,N_2274);
nor U2985 (N_2985,N_2438,N_2364);
and U2986 (N_2986,N_2251,N_2283);
or U2987 (N_2987,N_2146,N_2323);
nand U2988 (N_2988,N_2199,N_2437);
and U2989 (N_2989,N_2368,N_2254);
or U2990 (N_2990,N_2265,N_2222);
and U2991 (N_2991,N_2298,N_2062);
nand U2992 (N_2992,N_2313,N_2335);
nor U2993 (N_2993,N_2009,N_2222);
or U2994 (N_2994,N_2265,N_2348);
or U2995 (N_2995,N_2250,N_2144);
and U2996 (N_2996,N_2445,N_2496);
nand U2997 (N_2997,N_2225,N_2143);
or U2998 (N_2998,N_2156,N_2092);
and U2999 (N_2999,N_2343,N_2090);
and U3000 (N_3000,N_2687,N_2838);
or U3001 (N_3001,N_2746,N_2762);
nand U3002 (N_3002,N_2628,N_2938);
and U3003 (N_3003,N_2794,N_2845);
and U3004 (N_3004,N_2995,N_2647);
nor U3005 (N_3005,N_2935,N_2953);
and U3006 (N_3006,N_2779,N_2851);
or U3007 (N_3007,N_2664,N_2524);
nor U3008 (N_3008,N_2690,N_2721);
nand U3009 (N_3009,N_2643,N_2804);
nand U3010 (N_3010,N_2500,N_2785);
or U3011 (N_3011,N_2588,N_2822);
and U3012 (N_3012,N_2559,N_2850);
nor U3013 (N_3013,N_2522,N_2882);
or U3014 (N_3014,N_2554,N_2933);
nand U3015 (N_3015,N_2955,N_2878);
nor U3016 (N_3016,N_2833,N_2678);
and U3017 (N_3017,N_2830,N_2846);
and U3018 (N_3018,N_2709,N_2716);
or U3019 (N_3019,N_2871,N_2914);
nand U3020 (N_3020,N_2787,N_2684);
nand U3021 (N_3021,N_2911,N_2887);
and U3022 (N_3022,N_2579,N_2638);
nor U3023 (N_3023,N_2587,N_2671);
and U3024 (N_3024,N_2580,N_2849);
and U3025 (N_3025,N_2742,N_2738);
and U3026 (N_3026,N_2782,N_2751);
and U3027 (N_3027,N_2897,N_2867);
nand U3028 (N_3028,N_2823,N_2908);
xnor U3029 (N_3029,N_2552,N_2888);
or U3030 (N_3030,N_2784,N_2673);
and U3031 (N_3031,N_2650,N_2926);
and U3032 (N_3032,N_2909,N_2907);
and U3033 (N_3033,N_2863,N_2648);
nand U3034 (N_3034,N_2756,N_2977);
nor U3035 (N_3035,N_2841,N_2791);
nand U3036 (N_3036,N_2959,N_2798);
or U3037 (N_3037,N_2812,N_2665);
and U3038 (N_3038,N_2510,N_2964);
nand U3039 (N_3039,N_2915,N_2570);
or U3040 (N_3040,N_2952,N_2504);
and U3041 (N_3041,N_2624,N_2745);
nor U3042 (N_3042,N_2906,N_2610);
nor U3043 (N_3043,N_2621,N_2797);
and U3044 (N_3044,N_2544,N_2734);
nor U3045 (N_3045,N_2750,N_2567);
or U3046 (N_3046,N_2529,N_2972);
or U3047 (N_3047,N_2800,N_2770);
nand U3048 (N_3048,N_2505,N_2864);
or U3049 (N_3049,N_2825,N_2810);
and U3050 (N_3050,N_2950,N_2715);
nand U3051 (N_3051,N_2836,N_2795);
and U3052 (N_3052,N_2929,N_2605);
nor U3053 (N_3053,N_2555,N_2758);
nand U3054 (N_3054,N_2613,N_2549);
nor U3055 (N_3055,N_2595,N_2862);
and U3056 (N_3056,N_2661,N_2565);
nand U3057 (N_3057,N_2832,N_2821);
and U3058 (N_3058,N_2792,N_2966);
nor U3059 (N_3059,N_2930,N_2969);
nand U3060 (N_3060,N_2655,N_2543);
and U3061 (N_3061,N_2997,N_2847);
nor U3062 (N_3062,N_2598,N_2560);
or U3063 (N_3063,N_2509,N_2536);
and U3064 (N_3064,N_2516,N_2679);
or U3065 (N_3065,N_2582,N_2978);
nor U3066 (N_3066,N_2834,N_2688);
and U3067 (N_3067,N_2557,N_2667);
and U3068 (N_3068,N_2820,N_2828);
xor U3069 (N_3069,N_2521,N_2763);
or U3070 (N_3070,N_2880,N_2534);
nand U3071 (N_3071,N_2700,N_2652);
nor U3072 (N_3072,N_2551,N_2941);
and U3073 (N_3073,N_2723,N_2608);
nor U3074 (N_3074,N_2913,N_2803);
nor U3075 (N_3075,N_2872,N_2731);
or U3076 (N_3076,N_2827,N_2636);
nand U3077 (N_3077,N_2985,N_2818);
or U3078 (N_3078,N_2781,N_2506);
and U3079 (N_3079,N_2895,N_2642);
and U3080 (N_3080,N_2719,N_2732);
nor U3081 (N_3081,N_2829,N_2819);
and U3082 (N_3082,N_2837,N_2681);
or U3083 (N_3083,N_2601,N_2928);
nor U3084 (N_3084,N_2625,N_2835);
nand U3085 (N_3085,N_2620,N_2965);
nand U3086 (N_3086,N_2675,N_2635);
or U3087 (N_3087,N_2617,N_2893);
nand U3088 (N_3088,N_2693,N_2542);
nand U3089 (N_3089,N_2563,N_2607);
nand U3090 (N_3090,N_2736,N_2942);
and U3091 (N_3091,N_2753,N_2901);
nor U3092 (N_3092,N_2998,N_2924);
nand U3093 (N_3093,N_2739,N_2651);
or U3094 (N_3094,N_2912,N_2987);
and U3095 (N_3095,N_2527,N_2609);
and U3096 (N_3096,N_2535,N_2619);
nor U3097 (N_3097,N_2817,N_2511);
nand U3098 (N_3098,N_2986,N_2866);
and U3099 (N_3099,N_2634,N_2839);
nand U3100 (N_3100,N_2984,N_2729);
or U3101 (N_3101,N_2576,N_2712);
or U3102 (N_3102,N_2602,N_2528);
xor U3103 (N_3103,N_2523,N_2658);
and U3104 (N_3104,N_2581,N_2672);
nand U3105 (N_3105,N_2879,N_2730);
or U3106 (N_3106,N_2604,N_2632);
or U3107 (N_3107,N_2954,N_2944);
or U3108 (N_3108,N_2948,N_2532);
and U3109 (N_3109,N_2660,N_2718);
or U3110 (N_3110,N_2859,N_2513);
or U3111 (N_3111,N_2899,N_2512);
or U3112 (N_3112,N_2796,N_2857);
nor U3113 (N_3113,N_2980,N_2591);
and U3114 (N_3114,N_2783,N_2764);
nand U3115 (N_3115,N_2517,N_2889);
or U3116 (N_3116,N_2717,N_2566);
xnor U3117 (N_3117,N_2945,N_2865);
nand U3118 (N_3118,N_2801,N_2920);
or U3119 (N_3119,N_2943,N_2520);
or U3120 (N_3120,N_2577,N_2848);
xnor U3121 (N_3121,N_2724,N_2508);
nor U3122 (N_3122,N_2592,N_2548);
nand U3123 (N_3123,N_2695,N_2670);
nor U3124 (N_3124,N_2514,N_2816);
and U3125 (N_3125,N_2891,N_2640);
nand U3126 (N_3126,N_2844,N_2659);
nor U3127 (N_3127,N_2813,N_2765);
nor U3128 (N_3128,N_2789,N_2622);
or U3129 (N_3129,N_2852,N_2737);
and U3130 (N_3130,N_2776,N_2982);
nor U3131 (N_3131,N_2584,N_2873);
or U3132 (N_3132,N_2843,N_2713);
nand U3133 (N_3133,N_2631,N_2799);
or U3134 (N_3134,N_2708,N_2699);
nor U3135 (N_3135,N_2806,N_2698);
nand U3136 (N_3136,N_2957,N_2720);
and U3137 (N_3137,N_2735,N_2677);
nand U3138 (N_3138,N_2949,N_2627);
or U3139 (N_3139,N_2612,N_2733);
nand U3140 (N_3140,N_2572,N_2868);
nand U3141 (N_3141,N_2669,N_2961);
and U3142 (N_3142,N_2793,N_2975);
or U3143 (N_3143,N_2778,N_2769);
nor U3144 (N_3144,N_2540,N_2531);
nor U3145 (N_3145,N_2714,N_2518);
nor U3146 (N_3146,N_2947,N_2526);
nor U3147 (N_3147,N_2919,N_2749);
nand U3148 (N_3148,N_2855,N_2939);
or U3149 (N_3149,N_2963,N_2936);
or U3150 (N_3150,N_2589,N_2562);
nand U3151 (N_3151,N_2809,N_2663);
or U3152 (N_3152,N_2629,N_2903);
or U3153 (N_3153,N_2774,N_2940);
or U3154 (N_3154,N_2685,N_2722);
nand U3155 (N_3155,N_2645,N_2754);
nor U3156 (N_3156,N_2641,N_2996);
and U3157 (N_3157,N_2788,N_2860);
xor U3158 (N_3158,N_2550,N_2743);
nand U3159 (N_3159,N_2780,N_2777);
or U3160 (N_3160,N_2741,N_2707);
nor U3161 (N_3161,N_2662,N_2988);
or U3162 (N_3162,N_2556,N_2553);
and U3163 (N_3163,N_2680,N_2858);
nand U3164 (N_3164,N_2900,N_2958);
nor U3165 (N_3165,N_2596,N_2697);
nand U3166 (N_3166,N_2585,N_2507);
nor U3167 (N_3167,N_2545,N_2861);
and U3168 (N_3168,N_2918,N_2539);
and U3169 (N_3169,N_2773,N_2696);
or U3170 (N_3170,N_2547,N_2501);
nand U3171 (N_3171,N_2902,N_2842);
nor U3172 (N_3172,N_2759,N_2946);
or U3173 (N_3173,N_2761,N_2711);
nor U3174 (N_3174,N_2884,N_2917);
nand U3175 (N_3175,N_2811,N_2881);
nor U3176 (N_3176,N_2910,N_2686);
and U3177 (N_3177,N_2646,N_2757);
or U3178 (N_3178,N_2877,N_2633);
or U3179 (N_3179,N_2586,N_2979);
and U3180 (N_3180,N_2710,N_2876);
and U3181 (N_3181,N_2921,N_2525);
nor U3182 (N_3182,N_2706,N_2537);
or U3183 (N_3183,N_2649,N_2703);
and U3184 (N_3184,N_2702,N_2676);
and U3185 (N_3185,N_2568,N_2705);
or U3186 (N_3186,N_2771,N_2883);
nand U3187 (N_3187,N_2644,N_2970);
nand U3188 (N_3188,N_2593,N_2807);
nor U3189 (N_3189,N_2870,N_2561);
and U3190 (N_3190,N_2606,N_2668);
or U3191 (N_3191,N_2968,N_2656);
or U3192 (N_3192,N_2573,N_2519);
nand U3193 (N_3193,N_2597,N_2923);
nor U3194 (N_3194,N_2541,N_2981);
nor U3195 (N_3195,N_2875,N_2976);
and U3196 (N_3196,N_2630,N_2569);
or U3197 (N_3197,N_2626,N_2974);
nand U3198 (N_3198,N_2766,N_2682);
nand U3199 (N_3199,N_2775,N_2727);
nand U3200 (N_3200,N_2973,N_2874);
or U3201 (N_3201,N_2683,N_2916);
and U3202 (N_3202,N_2892,N_2932);
and U3203 (N_3203,N_2616,N_2728);
nor U3204 (N_3204,N_2740,N_2760);
and U3205 (N_3205,N_2971,N_2600);
nor U3206 (N_3206,N_2854,N_2993);
and U3207 (N_3207,N_2594,N_2802);
and U3208 (N_3208,N_2704,N_2931);
and U3209 (N_3209,N_2904,N_2960);
or U3210 (N_3210,N_2725,N_2666);
nand U3211 (N_3211,N_2808,N_2922);
nand U3212 (N_3212,N_2614,N_2890);
and U3213 (N_3213,N_2805,N_2815);
nor U3214 (N_3214,N_2654,N_2840);
nor U3215 (N_3215,N_2611,N_2691);
or U3216 (N_3216,N_2639,N_2772);
nand U3217 (N_3217,N_2564,N_2752);
or U3218 (N_3218,N_2885,N_2623);
and U3219 (N_3219,N_2558,N_2618);
nor U3220 (N_3220,N_2999,N_2755);
or U3221 (N_3221,N_2637,N_2994);
and U3222 (N_3222,N_2951,N_2694);
nand U3223 (N_3223,N_2853,N_2701);
or U3224 (N_3224,N_2599,N_2575);
and U3225 (N_3225,N_2992,N_2530);
nor U3226 (N_3226,N_2767,N_2934);
nand U3227 (N_3227,N_2962,N_2927);
or U3228 (N_3228,N_2603,N_2937);
or U3229 (N_3229,N_2896,N_2503);
nand U3230 (N_3230,N_2983,N_2786);
nand U3231 (N_3231,N_2824,N_2515);
nor U3232 (N_3232,N_2747,N_2894);
nand U3233 (N_3233,N_2689,N_2571);
nand U3234 (N_3234,N_2502,N_2925);
nand U3235 (N_3235,N_2989,N_2574);
or U3236 (N_3236,N_2615,N_2991);
and U3237 (N_3237,N_2748,N_2590);
or U3238 (N_3238,N_2653,N_2533);
or U3239 (N_3239,N_2898,N_2956);
xor U3240 (N_3240,N_2692,N_2814);
or U3241 (N_3241,N_2657,N_2538);
xnor U3242 (N_3242,N_2578,N_2856);
nand U3243 (N_3243,N_2583,N_2768);
nor U3244 (N_3244,N_2674,N_2744);
nor U3245 (N_3245,N_2826,N_2967);
nand U3246 (N_3246,N_2869,N_2831);
nor U3247 (N_3247,N_2990,N_2790);
or U3248 (N_3248,N_2546,N_2726);
and U3249 (N_3249,N_2905,N_2886);
and U3250 (N_3250,N_2987,N_2523);
and U3251 (N_3251,N_2586,N_2580);
nand U3252 (N_3252,N_2679,N_2557);
nand U3253 (N_3253,N_2608,N_2912);
nor U3254 (N_3254,N_2969,N_2566);
and U3255 (N_3255,N_2835,N_2871);
nor U3256 (N_3256,N_2530,N_2636);
nand U3257 (N_3257,N_2716,N_2852);
nor U3258 (N_3258,N_2839,N_2813);
nor U3259 (N_3259,N_2785,N_2635);
nand U3260 (N_3260,N_2852,N_2719);
or U3261 (N_3261,N_2672,N_2696);
and U3262 (N_3262,N_2607,N_2877);
nor U3263 (N_3263,N_2886,N_2563);
xor U3264 (N_3264,N_2696,N_2908);
nand U3265 (N_3265,N_2590,N_2710);
and U3266 (N_3266,N_2585,N_2978);
or U3267 (N_3267,N_2534,N_2953);
or U3268 (N_3268,N_2757,N_2989);
nand U3269 (N_3269,N_2985,N_2635);
or U3270 (N_3270,N_2834,N_2936);
nand U3271 (N_3271,N_2848,N_2648);
nand U3272 (N_3272,N_2776,N_2558);
nand U3273 (N_3273,N_2829,N_2603);
nor U3274 (N_3274,N_2587,N_2697);
or U3275 (N_3275,N_2513,N_2570);
and U3276 (N_3276,N_2564,N_2948);
and U3277 (N_3277,N_2697,N_2512);
xor U3278 (N_3278,N_2564,N_2674);
or U3279 (N_3279,N_2661,N_2948);
and U3280 (N_3280,N_2595,N_2656);
nand U3281 (N_3281,N_2806,N_2785);
or U3282 (N_3282,N_2879,N_2822);
nor U3283 (N_3283,N_2529,N_2970);
nor U3284 (N_3284,N_2528,N_2634);
or U3285 (N_3285,N_2845,N_2952);
and U3286 (N_3286,N_2844,N_2515);
and U3287 (N_3287,N_2921,N_2537);
nand U3288 (N_3288,N_2729,N_2745);
nor U3289 (N_3289,N_2922,N_2822);
nand U3290 (N_3290,N_2521,N_2852);
and U3291 (N_3291,N_2660,N_2759);
and U3292 (N_3292,N_2829,N_2617);
nand U3293 (N_3293,N_2553,N_2937);
nor U3294 (N_3294,N_2767,N_2806);
and U3295 (N_3295,N_2706,N_2767);
and U3296 (N_3296,N_2733,N_2679);
and U3297 (N_3297,N_2731,N_2990);
or U3298 (N_3298,N_2887,N_2541);
and U3299 (N_3299,N_2955,N_2874);
or U3300 (N_3300,N_2902,N_2918);
nor U3301 (N_3301,N_2503,N_2869);
and U3302 (N_3302,N_2712,N_2565);
and U3303 (N_3303,N_2889,N_2674);
and U3304 (N_3304,N_2726,N_2575);
and U3305 (N_3305,N_2582,N_2701);
and U3306 (N_3306,N_2921,N_2883);
or U3307 (N_3307,N_2789,N_2871);
or U3308 (N_3308,N_2547,N_2537);
or U3309 (N_3309,N_2875,N_2608);
nor U3310 (N_3310,N_2781,N_2544);
or U3311 (N_3311,N_2793,N_2754);
nand U3312 (N_3312,N_2920,N_2751);
nor U3313 (N_3313,N_2869,N_2906);
and U3314 (N_3314,N_2929,N_2746);
or U3315 (N_3315,N_2755,N_2631);
nand U3316 (N_3316,N_2535,N_2647);
nor U3317 (N_3317,N_2763,N_2788);
or U3318 (N_3318,N_2903,N_2907);
and U3319 (N_3319,N_2587,N_2710);
or U3320 (N_3320,N_2557,N_2695);
and U3321 (N_3321,N_2898,N_2662);
or U3322 (N_3322,N_2633,N_2985);
and U3323 (N_3323,N_2720,N_2663);
and U3324 (N_3324,N_2897,N_2600);
and U3325 (N_3325,N_2808,N_2580);
nand U3326 (N_3326,N_2865,N_2940);
nand U3327 (N_3327,N_2661,N_2810);
nor U3328 (N_3328,N_2794,N_2994);
or U3329 (N_3329,N_2604,N_2703);
nor U3330 (N_3330,N_2516,N_2909);
nand U3331 (N_3331,N_2509,N_2816);
or U3332 (N_3332,N_2946,N_2899);
and U3333 (N_3333,N_2752,N_2551);
xor U3334 (N_3334,N_2940,N_2624);
and U3335 (N_3335,N_2678,N_2970);
xor U3336 (N_3336,N_2543,N_2736);
nor U3337 (N_3337,N_2967,N_2736);
xnor U3338 (N_3338,N_2513,N_2640);
nor U3339 (N_3339,N_2894,N_2880);
nand U3340 (N_3340,N_2720,N_2981);
or U3341 (N_3341,N_2998,N_2620);
nand U3342 (N_3342,N_2882,N_2575);
nand U3343 (N_3343,N_2910,N_2949);
and U3344 (N_3344,N_2946,N_2860);
and U3345 (N_3345,N_2902,N_2816);
or U3346 (N_3346,N_2784,N_2835);
or U3347 (N_3347,N_2741,N_2689);
nand U3348 (N_3348,N_2756,N_2860);
nor U3349 (N_3349,N_2779,N_2614);
and U3350 (N_3350,N_2692,N_2822);
nand U3351 (N_3351,N_2709,N_2720);
xor U3352 (N_3352,N_2601,N_2909);
nor U3353 (N_3353,N_2750,N_2755);
and U3354 (N_3354,N_2645,N_2629);
or U3355 (N_3355,N_2705,N_2581);
nand U3356 (N_3356,N_2708,N_2567);
nand U3357 (N_3357,N_2620,N_2819);
or U3358 (N_3358,N_2781,N_2518);
nand U3359 (N_3359,N_2524,N_2601);
nand U3360 (N_3360,N_2600,N_2560);
nand U3361 (N_3361,N_2648,N_2669);
nor U3362 (N_3362,N_2781,N_2812);
and U3363 (N_3363,N_2737,N_2716);
nor U3364 (N_3364,N_2503,N_2844);
and U3365 (N_3365,N_2942,N_2896);
nand U3366 (N_3366,N_2671,N_2751);
and U3367 (N_3367,N_2548,N_2816);
or U3368 (N_3368,N_2824,N_2566);
or U3369 (N_3369,N_2831,N_2788);
nor U3370 (N_3370,N_2828,N_2572);
nor U3371 (N_3371,N_2917,N_2522);
and U3372 (N_3372,N_2708,N_2575);
and U3373 (N_3373,N_2615,N_2815);
or U3374 (N_3374,N_2954,N_2824);
or U3375 (N_3375,N_2534,N_2676);
and U3376 (N_3376,N_2767,N_2586);
and U3377 (N_3377,N_2568,N_2765);
or U3378 (N_3378,N_2632,N_2822);
and U3379 (N_3379,N_2737,N_2890);
nand U3380 (N_3380,N_2947,N_2892);
nor U3381 (N_3381,N_2725,N_2967);
nor U3382 (N_3382,N_2678,N_2971);
or U3383 (N_3383,N_2684,N_2764);
or U3384 (N_3384,N_2923,N_2512);
nand U3385 (N_3385,N_2849,N_2907);
nand U3386 (N_3386,N_2636,N_2895);
and U3387 (N_3387,N_2840,N_2703);
nand U3388 (N_3388,N_2953,N_2573);
nand U3389 (N_3389,N_2860,N_2678);
nor U3390 (N_3390,N_2580,N_2643);
or U3391 (N_3391,N_2835,N_2813);
and U3392 (N_3392,N_2917,N_2612);
or U3393 (N_3393,N_2544,N_2591);
or U3394 (N_3394,N_2905,N_2661);
or U3395 (N_3395,N_2524,N_2844);
and U3396 (N_3396,N_2810,N_2850);
nand U3397 (N_3397,N_2921,N_2544);
or U3398 (N_3398,N_2555,N_2836);
and U3399 (N_3399,N_2879,N_2751);
and U3400 (N_3400,N_2603,N_2624);
nor U3401 (N_3401,N_2862,N_2914);
and U3402 (N_3402,N_2896,N_2887);
and U3403 (N_3403,N_2714,N_2752);
xor U3404 (N_3404,N_2538,N_2784);
nor U3405 (N_3405,N_2704,N_2607);
nand U3406 (N_3406,N_2936,N_2555);
nor U3407 (N_3407,N_2860,N_2507);
nor U3408 (N_3408,N_2928,N_2513);
or U3409 (N_3409,N_2503,N_2887);
nand U3410 (N_3410,N_2606,N_2864);
and U3411 (N_3411,N_2871,N_2925);
nand U3412 (N_3412,N_2737,N_2573);
and U3413 (N_3413,N_2562,N_2536);
nor U3414 (N_3414,N_2991,N_2910);
nor U3415 (N_3415,N_2794,N_2769);
nor U3416 (N_3416,N_2969,N_2522);
nor U3417 (N_3417,N_2921,N_2972);
and U3418 (N_3418,N_2916,N_2770);
nand U3419 (N_3419,N_2584,N_2741);
nand U3420 (N_3420,N_2886,N_2636);
or U3421 (N_3421,N_2682,N_2626);
nor U3422 (N_3422,N_2716,N_2611);
or U3423 (N_3423,N_2775,N_2620);
and U3424 (N_3424,N_2598,N_2664);
and U3425 (N_3425,N_2825,N_2820);
or U3426 (N_3426,N_2700,N_2846);
nand U3427 (N_3427,N_2574,N_2742);
nand U3428 (N_3428,N_2680,N_2932);
nand U3429 (N_3429,N_2578,N_2724);
nand U3430 (N_3430,N_2994,N_2508);
nor U3431 (N_3431,N_2839,N_2949);
nor U3432 (N_3432,N_2650,N_2960);
or U3433 (N_3433,N_2576,N_2617);
and U3434 (N_3434,N_2924,N_2618);
nand U3435 (N_3435,N_2973,N_2546);
nor U3436 (N_3436,N_2508,N_2680);
nor U3437 (N_3437,N_2803,N_2567);
or U3438 (N_3438,N_2718,N_2929);
and U3439 (N_3439,N_2707,N_2943);
xor U3440 (N_3440,N_2961,N_2835);
or U3441 (N_3441,N_2644,N_2739);
nand U3442 (N_3442,N_2694,N_2541);
or U3443 (N_3443,N_2721,N_2804);
or U3444 (N_3444,N_2865,N_2577);
nand U3445 (N_3445,N_2611,N_2738);
nand U3446 (N_3446,N_2882,N_2847);
or U3447 (N_3447,N_2975,N_2814);
nor U3448 (N_3448,N_2844,N_2958);
or U3449 (N_3449,N_2863,N_2549);
nand U3450 (N_3450,N_2538,N_2579);
or U3451 (N_3451,N_2583,N_2524);
nand U3452 (N_3452,N_2715,N_2640);
or U3453 (N_3453,N_2760,N_2712);
or U3454 (N_3454,N_2510,N_2792);
or U3455 (N_3455,N_2907,N_2794);
nand U3456 (N_3456,N_2569,N_2889);
nand U3457 (N_3457,N_2696,N_2809);
and U3458 (N_3458,N_2587,N_2510);
nand U3459 (N_3459,N_2741,N_2810);
nand U3460 (N_3460,N_2993,N_2789);
nand U3461 (N_3461,N_2892,N_2926);
nor U3462 (N_3462,N_2993,N_2611);
nor U3463 (N_3463,N_2737,N_2671);
xnor U3464 (N_3464,N_2882,N_2670);
or U3465 (N_3465,N_2583,N_2872);
nand U3466 (N_3466,N_2923,N_2972);
nor U3467 (N_3467,N_2829,N_2888);
xor U3468 (N_3468,N_2549,N_2583);
or U3469 (N_3469,N_2998,N_2828);
nor U3470 (N_3470,N_2757,N_2644);
nand U3471 (N_3471,N_2607,N_2959);
or U3472 (N_3472,N_2512,N_2759);
or U3473 (N_3473,N_2772,N_2777);
or U3474 (N_3474,N_2530,N_2907);
or U3475 (N_3475,N_2667,N_2548);
or U3476 (N_3476,N_2645,N_2943);
and U3477 (N_3477,N_2686,N_2780);
nor U3478 (N_3478,N_2872,N_2770);
nand U3479 (N_3479,N_2506,N_2518);
nand U3480 (N_3480,N_2966,N_2605);
nor U3481 (N_3481,N_2640,N_2853);
and U3482 (N_3482,N_2858,N_2780);
nand U3483 (N_3483,N_2781,N_2854);
nor U3484 (N_3484,N_2761,N_2690);
and U3485 (N_3485,N_2962,N_2895);
nor U3486 (N_3486,N_2641,N_2549);
nand U3487 (N_3487,N_2859,N_2906);
nor U3488 (N_3488,N_2865,N_2730);
nand U3489 (N_3489,N_2781,N_2667);
nand U3490 (N_3490,N_2968,N_2993);
xor U3491 (N_3491,N_2911,N_2506);
or U3492 (N_3492,N_2712,N_2746);
nand U3493 (N_3493,N_2833,N_2946);
nand U3494 (N_3494,N_2793,N_2893);
nand U3495 (N_3495,N_2717,N_2638);
nand U3496 (N_3496,N_2772,N_2893);
and U3497 (N_3497,N_2582,N_2779);
nor U3498 (N_3498,N_2526,N_2678);
nor U3499 (N_3499,N_2569,N_2952);
or U3500 (N_3500,N_3416,N_3285);
nand U3501 (N_3501,N_3233,N_3455);
and U3502 (N_3502,N_3030,N_3106);
nor U3503 (N_3503,N_3318,N_3254);
or U3504 (N_3504,N_3368,N_3434);
and U3505 (N_3505,N_3265,N_3066);
nand U3506 (N_3506,N_3350,N_3483);
xnor U3507 (N_3507,N_3495,N_3371);
nor U3508 (N_3508,N_3435,N_3181);
nor U3509 (N_3509,N_3286,N_3305);
or U3510 (N_3510,N_3225,N_3330);
and U3511 (N_3511,N_3232,N_3157);
nand U3512 (N_3512,N_3478,N_3067);
or U3513 (N_3513,N_3464,N_3274);
nand U3514 (N_3514,N_3394,N_3211);
or U3515 (N_3515,N_3255,N_3208);
and U3516 (N_3516,N_3044,N_3325);
nand U3517 (N_3517,N_3117,N_3160);
nand U3518 (N_3518,N_3074,N_3126);
or U3519 (N_3519,N_3087,N_3475);
nor U3520 (N_3520,N_3084,N_3245);
or U3521 (N_3521,N_3467,N_3308);
or U3522 (N_3522,N_3338,N_3003);
and U3523 (N_3523,N_3174,N_3449);
nor U3524 (N_3524,N_3215,N_3111);
nor U3525 (N_3525,N_3257,N_3115);
or U3526 (N_3526,N_3349,N_3360);
nand U3527 (N_3527,N_3147,N_3344);
nor U3528 (N_3528,N_3000,N_3089);
or U3529 (N_3529,N_3304,N_3234);
nor U3530 (N_3530,N_3353,N_3073);
and U3531 (N_3531,N_3006,N_3493);
nor U3532 (N_3532,N_3033,N_3345);
nor U3533 (N_3533,N_3121,N_3322);
nor U3534 (N_3534,N_3410,N_3108);
and U3535 (N_3535,N_3195,N_3316);
nor U3536 (N_3536,N_3097,N_3118);
nor U3537 (N_3537,N_3002,N_3202);
nand U3538 (N_3538,N_3352,N_3240);
nor U3539 (N_3539,N_3071,N_3346);
and U3540 (N_3540,N_3358,N_3239);
and U3541 (N_3541,N_3385,N_3463);
nor U3542 (N_3542,N_3314,N_3259);
and U3543 (N_3543,N_3446,N_3153);
nor U3544 (N_3544,N_3300,N_3020);
or U3545 (N_3545,N_3333,N_3271);
and U3546 (N_3546,N_3065,N_3056);
nor U3547 (N_3547,N_3148,N_3373);
and U3548 (N_3548,N_3123,N_3027);
or U3549 (N_3549,N_3356,N_3445);
and U3550 (N_3550,N_3320,N_3028);
nand U3551 (N_3551,N_3465,N_3399);
nand U3552 (N_3552,N_3243,N_3266);
nand U3553 (N_3553,N_3339,N_3041);
or U3554 (N_3554,N_3223,N_3487);
nand U3555 (N_3555,N_3076,N_3175);
nand U3556 (N_3556,N_3008,N_3143);
nand U3557 (N_3557,N_3100,N_3139);
nand U3558 (N_3558,N_3480,N_3023);
or U3559 (N_3559,N_3354,N_3253);
nand U3560 (N_3560,N_3297,N_3343);
or U3561 (N_3561,N_3161,N_3389);
and U3562 (N_3562,N_3430,N_3079);
nand U3563 (N_3563,N_3311,N_3136);
and U3564 (N_3564,N_3213,N_3229);
nor U3565 (N_3565,N_3321,N_3331);
and U3566 (N_3566,N_3370,N_3107);
and U3567 (N_3567,N_3158,N_3263);
nand U3568 (N_3568,N_3193,N_3357);
xnor U3569 (N_3569,N_3043,N_3280);
nor U3570 (N_3570,N_3277,N_3024);
nor U3571 (N_3571,N_3200,N_3101);
and U3572 (N_3572,N_3196,N_3422);
and U3573 (N_3573,N_3238,N_3273);
nor U3574 (N_3574,N_3194,N_3085);
or U3575 (N_3575,N_3301,N_3429);
nand U3576 (N_3576,N_3461,N_3369);
and U3577 (N_3577,N_3119,N_3319);
nand U3578 (N_3578,N_3359,N_3275);
or U3579 (N_3579,N_3295,N_3454);
or U3580 (N_3580,N_3047,N_3070);
nor U3581 (N_3581,N_3267,N_3269);
or U3582 (N_3582,N_3420,N_3282);
and U3583 (N_3583,N_3127,N_3260);
or U3584 (N_3584,N_3432,N_3362);
nand U3585 (N_3585,N_3062,N_3381);
nor U3586 (N_3586,N_3468,N_3132);
xnor U3587 (N_3587,N_3293,N_3165);
nor U3588 (N_3588,N_3015,N_3090);
or U3589 (N_3589,N_3496,N_3116);
and U3590 (N_3590,N_3452,N_3072);
nand U3591 (N_3591,N_3005,N_3186);
nand U3592 (N_3592,N_3185,N_3110);
nand U3593 (N_3593,N_3479,N_3222);
nand U3594 (N_3594,N_3383,N_3060);
and U3595 (N_3595,N_3207,N_3302);
or U3596 (N_3596,N_3387,N_3492);
and U3597 (N_3597,N_3057,N_3376);
nand U3598 (N_3598,N_3094,N_3182);
nand U3599 (N_3599,N_3201,N_3334);
nor U3600 (N_3600,N_3135,N_3477);
nor U3601 (N_3601,N_3444,N_3247);
nand U3602 (N_3602,N_3283,N_3406);
nand U3603 (N_3603,N_3264,N_3258);
or U3604 (N_3604,N_3235,N_3405);
nor U3605 (N_3605,N_3155,N_3324);
nand U3606 (N_3606,N_3241,N_3279);
or U3607 (N_3607,N_3291,N_3313);
or U3608 (N_3608,N_3173,N_3411);
or U3609 (N_3609,N_3290,N_3372);
nor U3610 (N_3610,N_3425,N_3162);
or U3611 (N_3611,N_3326,N_3388);
or U3612 (N_3612,N_3227,N_3018);
nand U3613 (N_3613,N_3098,N_3191);
nor U3614 (N_3614,N_3337,N_3437);
or U3615 (N_3615,N_3484,N_3138);
and U3616 (N_3616,N_3045,N_3251);
nand U3617 (N_3617,N_3340,N_3159);
nand U3618 (N_3618,N_3113,N_3306);
nor U3619 (N_3619,N_3210,N_3105);
nor U3620 (N_3620,N_3317,N_3268);
and U3621 (N_3621,N_3374,N_3332);
xor U3622 (N_3622,N_3424,N_3055);
nand U3623 (N_3623,N_3114,N_3204);
or U3624 (N_3624,N_3011,N_3052);
nor U3625 (N_3625,N_3236,N_3366);
and U3626 (N_3626,N_3178,N_3365);
or U3627 (N_3627,N_3363,N_3412);
and U3628 (N_3628,N_3379,N_3036);
or U3629 (N_3629,N_3287,N_3403);
nor U3630 (N_3630,N_3054,N_3310);
nor U3631 (N_3631,N_3140,N_3217);
nand U3632 (N_3632,N_3081,N_3262);
or U3633 (N_3633,N_3038,N_3197);
or U3634 (N_3634,N_3099,N_3261);
nor U3635 (N_3635,N_3228,N_3413);
or U3636 (N_3636,N_3309,N_3426);
and U3637 (N_3637,N_3169,N_3401);
or U3638 (N_3638,N_3329,N_3409);
or U3639 (N_3639,N_3294,N_3292);
nor U3640 (N_3640,N_3447,N_3443);
or U3641 (N_3641,N_3029,N_3392);
and U3642 (N_3642,N_3364,N_3377);
nor U3643 (N_3643,N_3237,N_3187);
nor U3644 (N_3644,N_3209,N_3164);
nand U3645 (N_3645,N_3246,N_3198);
and U3646 (N_3646,N_3490,N_3244);
or U3647 (N_3647,N_3250,N_3378);
nand U3648 (N_3648,N_3315,N_3440);
nor U3649 (N_3649,N_3408,N_3145);
and U3650 (N_3650,N_3249,N_3031);
and U3651 (N_3651,N_3231,N_3397);
xor U3652 (N_3652,N_3184,N_3404);
nand U3653 (N_3653,N_3386,N_3288);
and U3654 (N_3654,N_3137,N_3407);
and U3655 (N_3655,N_3384,N_3303);
nor U3656 (N_3656,N_3172,N_3335);
or U3657 (N_3657,N_3048,N_3142);
and U3658 (N_3658,N_3489,N_3451);
nor U3659 (N_3659,N_3088,N_3152);
or U3660 (N_3660,N_3400,N_3336);
nor U3661 (N_3661,N_3486,N_3206);
or U3662 (N_3662,N_3456,N_3242);
or U3663 (N_3663,N_3323,N_3433);
and U3664 (N_3664,N_3391,N_3494);
or U3665 (N_3665,N_3428,N_3009);
or U3666 (N_3666,N_3199,N_3012);
nand U3667 (N_3667,N_3472,N_3216);
nand U3668 (N_3668,N_3039,N_3019);
nor U3669 (N_3669,N_3469,N_3341);
nor U3670 (N_3670,N_3001,N_3393);
nor U3671 (N_3671,N_3183,N_3252);
and U3672 (N_3672,N_3453,N_3007);
or U3673 (N_3673,N_3458,N_3219);
and U3674 (N_3674,N_3080,N_3141);
nand U3675 (N_3675,N_3205,N_3129);
or U3676 (N_3676,N_3224,N_3004);
and U3677 (N_3677,N_3328,N_3382);
nand U3678 (N_3678,N_3281,N_3485);
or U3679 (N_3679,N_3040,N_3083);
or U3680 (N_3680,N_3093,N_3154);
nor U3681 (N_3681,N_3276,N_3396);
nor U3682 (N_3682,N_3498,N_3395);
nand U3683 (N_3683,N_3450,N_3462);
or U3684 (N_3684,N_3298,N_3375);
or U3685 (N_3685,N_3482,N_3168);
nand U3686 (N_3686,N_3166,N_3069);
and U3687 (N_3687,N_3431,N_3156);
or U3688 (N_3688,N_3144,N_3095);
or U3689 (N_3689,N_3421,N_3361);
and U3690 (N_3690,N_3131,N_3417);
or U3691 (N_3691,N_3488,N_3307);
or U3692 (N_3692,N_3058,N_3064);
nand U3693 (N_3693,N_3471,N_3355);
and U3694 (N_3694,N_3016,N_3218);
nor U3695 (N_3695,N_3180,N_3367);
nand U3696 (N_3696,N_3167,N_3436);
or U3697 (N_3697,N_3068,N_3189);
nor U3698 (N_3698,N_3212,N_3092);
nand U3699 (N_3699,N_3457,N_3078);
nand U3700 (N_3700,N_3050,N_3125);
nand U3701 (N_3701,N_3439,N_3284);
and U3702 (N_3702,N_3063,N_3046);
nor U3703 (N_3703,N_3203,N_3256);
nand U3704 (N_3704,N_3013,N_3086);
and U3705 (N_3705,N_3221,N_3026);
or U3706 (N_3706,N_3418,N_3299);
nor U3707 (N_3707,N_3351,N_3312);
nor U3708 (N_3708,N_3230,N_3077);
nor U3709 (N_3709,N_3278,N_3120);
nand U3710 (N_3710,N_3014,N_3053);
or U3711 (N_3711,N_3130,N_3327);
xor U3712 (N_3712,N_3049,N_3104);
nor U3713 (N_3713,N_3150,N_3025);
nor U3714 (N_3714,N_3163,N_3248);
nor U3715 (N_3715,N_3473,N_3438);
nand U3716 (N_3716,N_3146,N_3134);
nor U3717 (N_3717,N_3021,N_3051);
and U3718 (N_3718,N_3214,N_3102);
or U3719 (N_3719,N_3176,N_3442);
nand U3720 (N_3720,N_3188,N_3034);
and U3721 (N_3721,N_3124,N_3476);
or U3722 (N_3722,N_3037,N_3226);
and U3723 (N_3723,N_3220,N_3042);
or U3724 (N_3724,N_3423,N_3151);
and U3725 (N_3725,N_3427,N_3348);
nand U3726 (N_3726,N_3289,N_3075);
nand U3727 (N_3727,N_3491,N_3459);
and U3728 (N_3728,N_3441,N_3390);
nor U3729 (N_3729,N_3177,N_3103);
nand U3730 (N_3730,N_3170,N_3380);
nand U3731 (N_3731,N_3010,N_3112);
nand U3732 (N_3732,N_3481,N_3419);
nand U3733 (N_3733,N_3414,N_3190);
nor U3734 (N_3734,N_3460,N_3109);
and U3735 (N_3735,N_3149,N_3059);
or U3736 (N_3736,N_3128,N_3035);
nor U3737 (N_3737,N_3082,N_3171);
and U3738 (N_3738,N_3032,N_3096);
xnor U3739 (N_3739,N_3474,N_3091);
nand U3740 (N_3740,N_3415,N_3017);
nand U3741 (N_3741,N_3398,N_3466);
nand U3742 (N_3742,N_3122,N_3296);
nand U3743 (N_3743,N_3499,N_3448);
and U3744 (N_3744,N_3061,N_3022);
or U3745 (N_3745,N_3497,N_3470);
and U3746 (N_3746,N_3402,N_3347);
or U3747 (N_3747,N_3342,N_3272);
nor U3748 (N_3748,N_3270,N_3179);
and U3749 (N_3749,N_3192,N_3133);
nor U3750 (N_3750,N_3187,N_3460);
and U3751 (N_3751,N_3007,N_3433);
or U3752 (N_3752,N_3475,N_3395);
or U3753 (N_3753,N_3493,N_3097);
nand U3754 (N_3754,N_3453,N_3317);
nand U3755 (N_3755,N_3364,N_3040);
nor U3756 (N_3756,N_3138,N_3100);
nor U3757 (N_3757,N_3114,N_3362);
nor U3758 (N_3758,N_3151,N_3141);
and U3759 (N_3759,N_3338,N_3286);
nand U3760 (N_3760,N_3264,N_3252);
or U3761 (N_3761,N_3156,N_3212);
nand U3762 (N_3762,N_3170,N_3285);
nand U3763 (N_3763,N_3171,N_3493);
or U3764 (N_3764,N_3095,N_3323);
or U3765 (N_3765,N_3335,N_3104);
nand U3766 (N_3766,N_3352,N_3334);
or U3767 (N_3767,N_3287,N_3001);
and U3768 (N_3768,N_3131,N_3245);
or U3769 (N_3769,N_3065,N_3186);
and U3770 (N_3770,N_3064,N_3316);
or U3771 (N_3771,N_3443,N_3309);
nand U3772 (N_3772,N_3053,N_3360);
nor U3773 (N_3773,N_3496,N_3349);
xor U3774 (N_3774,N_3430,N_3335);
or U3775 (N_3775,N_3066,N_3411);
nand U3776 (N_3776,N_3346,N_3048);
and U3777 (N_3777,N_3150,N_3078);
or U3778 (N_3778,N_3314,N_3297);
nor U3779 (N_3779,N_3432,N_3253);
nand U3780 (N_3780,N_3406,N_3373);
nor U3781 (N_3781,N_3034,N_3462);
or U3782 (N_3782,N_3045,N_3269);
and U3783 (N_3783,N_3464,N_3197);
and U3784 (N_3784,N_3277,N_3093);
or U3785 (N_3785,N_3088,N_3340);
and U3786 (N_3786,N_3359,N_3440);
or U3787 (N_3787,N_3481,N_3423);
or U3788 (N_3788,N_3011,N_3157);
xnor U3789 (N_3789,N_3470,N_3015);
nor U3790 (N_3790,N_3404,N_3110);
nor U3791 (N_3791,N_3226,N_3085);
and U3792 (N_3792,N_3046,N_3086);
nand U3793 (N_3793,N_3186,N_3075);
and U3794 (N_3794,N_3430,N_3318);
and U3795 (N_3795,N_3253,N_3077);
and U3796 (N_3796,N_3206,N_3282);
nor U3797 (N_3797,N_3308,N_3172);
nor U3798 (N_3798,N_3012,N_3243);
or U3799 (N_3799,N_3123,N_3021);
nor U3800 (N_3800,N_3101,N_3265);
and U3801 (N_3801,N_3453,N_3086);
or U3802 (N_3802,N_3073,N_3444);
nor U3803 (N_3803,N_3228,N_3031);
nor U3804 (N_3804,N_3289,N_3295);
or U3805 (N_3805,N_3429,N_3347);
nor U3806 (N_3806,N_3168,N_3242);
nor U3807 (N_3807,N_3067,N_3055);
and U3808 (N_3808,N_3068,N_3368);
or U3809 (N_3809,N_3149,N_3260);
nor U3810 (N_3810,N_3434,N_3070);
or U3811 (N_3811,N_3462,N_3120);
and U3812 (N_3812,N_3263,N_3455);
or U3813 (N_3813,N_3026,N_3032);
or U3814 (N_3814,N_3402,N_3113);
and U3815 (N_3815,N_3405,N_3363);
nor U3816 (N_3816,N_3443,N_3469);
or U3817 (N_3817,N_3361,N_3330);
or U3818 (N_3818,N_3244,N_3308);
and U3819 (N_3819,N_3341,N_3160);
or U3820 (N_3820,N_3418,N_3470);
or U3821 (N_3821,N_3365,N_3463);
and U3822 (N_3822,N_3472,N_3076);
nor U3823 (N_3823,N_3213,N_3160);
nand U3824 (N_3824,N_3379,N_3179);
or U3825 (N_3825,N_3150,N_3377);
nor U3826 (N_3826,N_3323,N_3321);
and U3827 (N_3827,N_3212,N_3235);
or U3828 (N_3828,N_3405,N_3398);
or U3829 (N_3829,N_3497,N_3453);
or U3830 (N_3830,N_3117,N_3250);
and U3831 (N_3831,N_3050,N_3272);
nand U3832 (N_3832,N_3411,N_3418);
or U3833 (N_3833,N_3418,N_3020);
nor U3834 (N_3834,N_3288,N_3243);
nor U3835 (N_3835,N_3306,N_3186);
nand U3836 (N_3836,N_3090,N_3183);
and U3837 (N_3837,N_3268,N_3353);
nor U3838 (N_3838,N_3270,N_3109);
or U3839 (N_3839,N_3235,N_3342);
nand U3840 (N_3840,N_3339,N_3324);
nand U3841 (N_3841,N_3116,N_3184);
nor U3842 (N_3842,N_3301,N_3233);
and U3843 (N_3843,N_3381,N_3129);
or U3844 (N_3844,N_3092,N_3057);
and U3845 (N_3845,N_3290,N_3453);
nor U3846 (N_3846,N_3413,N_3247);
nand U3847 (N_3847,N_3362,N_3000);
nand U3848 (N_3848,N_3105,N_3050);
nand U3849 (N_3849,N_3279,N_3399);
nor U3850 (N_3850,N_3402,N_3125);
or U3851 (N_3851,N_3128,N_3038);
nor U3852 (N_3852,N_3372,N_3438);
nand U3853 (N_3853,N_3421,N_3146);
and U3854 (N_3854,N_3002,N_3470);
and U3855 (N_3855,N_3424,N_3038);
and U3856 (N_3856,N_3490,N_3365);
nor U3857 (N_3857,N_3493,N_3042);
or U3858 (N_3858,N_3212,N_3086);
nor U3859 (N_3859,N_3456,N_3085);
and U3860 (N_3860,N_3086,N_3402);
and U3861 (N_3861,N_3214,N_3431);
nand U3862 (N_3862,N_3312,N_3479);
or U3863 (N_3863,N_3221,N_3235);
nor U3864 (N_3864,N_3374,N_3265);
or U3865 (N_3865,N_3264,N_3246);
and U3866 (N_3866,N_3389,N_3237);
nand U3867 (N_3867,N_3231,N_3484);
nand U3868 (N_3868,N_3386,N_3383);
nand U3869 (N_3869,N_3119,N_3197);
or U3870 (N_3870,N_3438,N_3122);
and U3871 (N_3871,N_3241,N_3183);
nand U3872 (N_3872,N_3219,N_3433);
nand U3873 (N_3873,N_3153,N_3020);
or U3874 (N_3874,N_3119,N_3065);
or U3875 (N_3875,N_3476,N_3056);
nor U3876 (N_3876,N_3162,N_3178);
nand U3877 (N_3877,N_3377,N_3203);
nand U3878 (N_3878,N_3239,N_3116);
nor U3879 (N_3879,N_3408,N_3088);
or U3880 (N_3880,N_3494,N_3340);
nor U3881 (N_3881,N_3148,N_3165);
or U3882 (N_3882,N_3376,N_3001);
and U3883 (N_3883,N_3008,N_3315);
and U3884 (N_3884,N_3250,N_3284);
nor U3885 (N_3885,N_3354,N_3052);
or U3886 (N_3886,N_3034,N_3374);
xnor U3887 (N_3887,N_3299,N_3220);
nand U3888 (N_3888,N_3193,N_3196);
nor U3889 (N_3889,N_3158,N_3090);
nor U3890 (N_3890,N_3256,N_3202);
nor U3891 (N_3891,N_3425,N_3492);
nand U3892 (N_3892,N_3291,N_3307);
nor U3893 (N_3893,N_3469,N_3472);
nand U3894 (N_3894,N_3479,N_3159);
nand U3895 (N_3895,N_3195,N_3447);
and U3896 (N_3896,N_3049,N_3018);
or U3897 (N_3897,N_3159,N_3488);
nand U3898 (N_3898,N_3219,N_3333);
and U3899 (N_3899,N_3021,N_3024);
nand U3900 (N_3900,N_3409,N_3007);
nand U3901 (N_3901,N_3344,N_3014);
nor U3902 (N_3902,N_3258,N_3354);
and U3903 (N_3903,N_3079,N_3074);
or U3904 (N_3904,N_3238,N_3326);
or U3905 (N_3905,N_3046,N_3100);
nand U3906 (N_3906,N_3357,N_3065);
nor U3907 (N_3907,N_3456,N_3125);
nand U3908 (N_3908,N_3015,N_3464);
or U3909 (N_3909,N_3279,N_3016);
nor U3910 (N_3910,N_3006,N_3305);
nand U3911 (N_3911,N_3493,N_3124);
nor U3912 (N_3912,N_3256,N_3479);
nand U3913 (N_3913,N_3073,N_3074);
and U3914 (N_3914,N_3049,N_3198);
nor U3915 (N_3915,N_3104,N_3007);
nor U3916 (N_3916,N_3368,N_3196);
nor U3917 (N_3917,N_3403,N_3425);
nor U3918 (N_3918,N_3176,N_3212);
or U3919 (N_3919,N_3342,N_3436);
nor U3920 (N_3920,N_3231,N_3236);
or U3921 (N_3921,N_3383,N_3075);
nor U3922 (N_3922,N_3149,N_3259);
and U3923 (N_3923,N_3428,N_3489);
or U3924 (N_3924,N_3454,N_3467);
nand U3925 (N_3925,N_3254,N_3384);
nand U3926 (N_3926,N_3249,N_3424);
and U3927 (N_3927,N_3126,N_3449);
or U3928 (N_3928,N_3495,N_3218);
nand U3929 (N_3929,N_3194,N_3089);
or U3930 (N_3930,N_3411,N_3424);
nand U3931 (N_3931,N_3346,N_3446);
and U3932 (N_3932,N_3019,N_3494);
or U3933 (N_3933,N_3305,N_3096);
nor U3934 (N_3934,N_3411,N_3442);
or U3935 (N_3935,N_3263,N_3212);
nor U3936 (N_3936,N_3432,N_3383);
or U3937 (N_3937,N_3285,N_3053);
nand U3938 (N_3938,N_3271,N_3446);
or U3939 (N_3939,N_3009,N_3183);
nand U3940 (N_3940,N_3258,N_3221);
and U3941 (N_3941,N_3052,N_3270);
and U3942 (N_3942,N_3325,N_3358);
or U3943 (N_3943,N_3321,N_3087);
and U3944 (N_3944,N_3371,N_3245);
nand U3945 (N_3945,N_3480,N_3151);
nand U3946 (N_3946,N_3183,N_3467);
and U3947 (N_3947,N_3398,N_3232);
or U3948 (N_3948,N_3429,N_3117);
nand U3949 (N_3949,N_3383,N_3299);
nand U3950 (N_3950,N_3478,N_3483);
or U3951 (N_3951,N_3064,N_3089);
or U3952 (N_3952,N_3082,N_3085);
and U3953 (N_3953,N_3410,N_3199);
and U3954 (N_3954,N_3002,N_3452);
nand U3955 (N_3955,N_3477,N_3286);
or U3956 (N_3956,N_3127,N_3484);
nand U3957 (N_3957,N_3297,N_3448);
nor U3958 (N_3958,N_3341,N_3401);
nor U3959 (N_3959,N_3014,N_3140);
nand U3960 (N_3960,N_3248,N_3489);
nor U3961 (N_3961,N_3451,N_3438);
nor U3962 (N_3962,N_3271,N_3473);
and U3963 (N_3963,N_3423,N_3229);
nor U3964 (N_3964,N_3393,N_3437);
nand U3965 (N_3965,N_3259,N_3400);
nand U3966 (N_3966,N_3203,N_3118);
or U3967 (N_3967,N_3330,N_3290);
nand U3968 (N_3968,N_3348,N_3001);
or U3969 (N_3969,N_3242,N_3237);
nor U3970 (N_3970,N_3359,N_3458);
or U3971 (N_3971,N_3052,N_3102);
and U3972 (N_3972,N_3052,N_3483);
and U3973 (N_3973,N_3451,N_3348);
nor U3974 (N_3974,N_3444,N_3053);
nor U3975 (N_3975,N_3410,N_3019);
nor U3976 (N_3976,N_3076,N_3345);
and U3977 (N_3977,N_3138,N_3468);
and U3978 (N_3978,N_3251,N_3282);
nor U3979 (N_3979,N_3073,N_3186);
and U3980 (N_3980,N_3169,N_3246);
or U3981 (N_3981,N_3033,N_3346);
and U3982 (N_3982,N_3199,N_3254);
and U3983 (N_3983,N_3327,N_3215);
nand U3984 (N_3984,N_3376,N_3094);
or U3985 (N_3985,N_3040,N_3370);
or U3986 (N_3986,N_3190,N_3250);
or U3987 (N_3987,N_3210,N_3435);
nand U3988 (N_3988,N_3101,N_3136);
and U3989 (N_3989,N_3322,N_3048);
and U3990 (N_3990,N_3375,N_3383);
or U3991 (N_3991,N_3343,N_3435);
nand U3992 (N_3992,N_3433,N_3336);
and U3993 (N_3993,N_3035,N_3183);
nand U3994 (N_3994,N_3142,N_3146);
nand U3995 (N_3995,N_3078,N_3026);
or U3996 (N_3996,N_3469,N_3404);
or U3997 (N_3997,N_3445,N_3140);
nor U3998 (N_3998,N_3274,N_3334);
or U3999 (N_3999,N_3020,N_3121);
and U4000 (N_4000,N_3573,N_3934);
and U4001 (N_4001,N_3524,N_3958);
xnor U4002 (N_4002,N_3689,N_3578);
nor U4003 (N_4003,N_3835,N_3621);
or U4004 (N_4004,N_3556,N_3932);
or U4005 (N_4005,N_3552,N_3572);
nand U4006 (N_4006,N_3724,N_3534);
nand U4007 (N_4007,N_3865,N_3655);
or U4008 (N_4008,N_3959,N_3570);
nor U4009 (N_4009,N_3577,N_3583);
and U4010 (N_4010,N_3988,N_3858);
or U4011 (N_4011,N_3823,N_3997);
or U4012 (N_4012,N_3853,N_3783);
nand U4013 (N_4013,N_3543,N_3864);
nor U4014 (N_4014,N_3935,N_3920);
and U4015 (N_4015,N_3993,N_3923);
nand U4016 (N_4016,N_3698,N_3947);
and U4017 (N_4017,N_3620,N_3944);
and U4018 (N_4018,N_3593,N_3643);
or U4019 (N_4019,N_3841,N_3764);
or U4020 (N_4020,N_3897,N_3697);
or U4021 (N_4021,N_3690,N_3852);
and U4022 (N_4022,N_3527,N_3905);
nand U4023 (N_4023,N_3792,N_3508);
nand U4024 (N_4024,N_3733,N_3972);
and U4025 (N_4025,N_3804,N_3712);
nor U4026 (N_4026,N_3629,N_3706);
nor U4027 (N_4027,N_3674,N_3505);
and U4028 (N_4028,N_3633,N_3693);
or U4029 (N_4029,N_3607,N_3774);
nor U4030 (N_4030,N_3576,N_3631);
nor U4031 (N_4031,N_3555,N_3710);
or U4032 (N_4032,N_3761,N_3654);
nor U4033 (N_4033,N_3845,N_3789);
or U4034 (N_4034,N_3554,N_3960);
or U4035 (N_4035,N_3821,N_3614);
nor U4036 (N_4036,N_3588,N_3688);
nand U4037 (N_4037,N_3784,N_3538);
or U4038 (N_4038,N_3564,N_3591);
or U4039 (N_4039,N_3989,N_3684);
nand U4040 (N_4040,N_3998,N_3877);
or U4041 (N_4041,N_3969,N_3600);
nand U4042 (N_4042,N_3545,N_3904);
nor U4043 (N_4043,N_3682,N_3863);
nor U4044 (N_4044,N_3504,N_3879);
or U4045 (N_4045,N_3541,N_3994);
or U4046 (N_4046,N_3736,N_3616);
nand U4047 (N_4047,N_3916,N_3762);
and U4048 (N_4048,N_3756,N_3531);
and U4049 (N_4049,N_3526,N_3748);
nor U4050 (N_4050,N_3846,N_3670);
nand U4051 (N_4051,N_3899,N_3651);
or U4052 (N_4052,N_3919,N_3780);
nand U4053 (N_4053,N_3601,N_3820);
or U4054 (N_4054,N_3833,N_3940);
nand U4055 (N_4055,N_3608,N_3847);
and U4056 (N_4056,N_3642,N_3788);
or U4057 (N_4057,N_3571,N_3721);
and U4058 (N_4058,N_3796,N_3895);
and U4059 (N_4059,N_3778,N_3671);
and U4060 (N_4060,N_3569,N_3917);
nor U4061 (N_4061,N_3525,N_3799);
nor U4062 (N_4062,N_3943,N_3679);
nand U4063 (N_4063,N_3903,N_3647);
or U4064 (N_4064,N_3968,N_3992);
or U4065 (N_4065,N_3518,N_3735);
or U4066 (N_4066,N_3834,N_3645);
nand U4067 (N_4067,N_3510,N_3530);
or U4068 (N_4068,N_3840,N_3549);
and U4069 (N_4069,N_3507,N_3560);
nand U4070 (N_4070,N_3786,N_3639);
nor U4071 (N_4071,N_3941,N_3626);
nor U4072 (N_4072,N_3907,N_3584);
and U4073 (N_4073,N_3597,N_3665);
nand U4074 (N_4074,N_3758,N_3886);
or U4075 (N_4075,N_3949,N_3668);
or U4076 (N_4076,N_3678,N_3807);
nor U4077 (N_4077,N_3815,N_3950);
nor U4078 (N_4078,N_3759,N_3811);
nor U4079 (N_4079,N_3791,N_3962);
or U4080 (N_4080,N_3876,N_3715);
nand U4081 (N_4081,N_3767,N_3931);
and U4082 (N_4082,N_3635,N_3661);
nand U4083 (N_4083,N_3930,N_3888);
or U4084 (N_4084,N_3768,N_3825);
nand U4085 (N_4085,N_3836,N_3869);
nor U4086 (N_4086,N_3656,N_3704);
nand U4087 (N_4087,N_3596,N_3963);
or U4088 (N_4088,N_3727,N_3937);
and U4089 (N_4089,N_3967,N_3819);
or U4090 (N_4090,N_3892,N_3535);
nor U4091 (N_4091,N_3641,N_3649);
or U4092 (N_4092,N_3782,N_3831);
nor U4093 (N_4093,N_3722,N_3632);
or U4094 (N_4094,N_3622,N_3906);
nor U4095 (N_4095,N_3559,N_3849);
or U4096 (N_4096,N_3884,N_3734);
or U4097 (N_4097,N_3924,N_3516);
and U4098 (N_4098,N_3702,N_3514);
or U4099 (N_4099,N_3680,N_3793);
and U4100 (N_4100,N_3775,N_3961);
and U4101 (N_4101,N_3856,N_3982);
and U4102 (N_4102,N_3589,N_3829);
nand U4103 (N_4103,N_3558,N_3760);
nor U4104 (N_4104,N_3540,N_3598);
nor U4105 (N_4105,N_3539,N_3557);
or U4106 (N_4106,N_3746,N_3754);
and U4107 (N_4107,N_3975,N_3658);
or U4108 (N_4108,N_3817,N_3749);
or U4109 (N_4109,N_3851,N_3609);
and U4110 (N_4110,N_3602,N_3615);
or U4111 (N_4111,N_3826,N_3890);
and U4112 (N_4112,N_3562,N_3563);
nor U4113 (N_4113,N_3717,N_3725);
or U4114 (N_4114,N_3750,N_3536);
nand U4115 (N_4115,N_3805,N_3716);
or U4116 (N_4116,N_3999,N_3741);
and U4117 (N_4117,N_3870,N_3878);
and U4118 (N_4118,N_3981,N_3914);
or U4119 (N_4119,N_3985,N_3520);
nand U4120 (N_4120,N_3973,N_3648);
nand U4121 (N_4121,N_3942,N_3787);
and U4122 (N_4122,N_3695,N_3585);
and U4123 (N_4123,N_3785,N_3548);
or U4124 (N_4124,N_3922,N_3744);
nor U4125 (N_4125,N_3995,N_3737);
or U4126 (N_4126,N_3669,N_3844);
or U4127 (N_4127,N_3883,N_3551);
or U4128 (N_4128,N_3984,N_3765);
nor U4129 (N_4129,N_3537,N_3705);
nand U4130 (N_4130,N_3606,N_3955);
and U4131 (N_4131,N_3986,N_3766);
nand U4132 (N_4132,N_3664,N_3732);
and U4133 (N_4133,N_3723,N_3842);
nor U4134 (N_4134,N_3553,N_3751);
nand U4135 (N_4135,N_3757,N_3595);
nor U4136 (N_4136,N_3918,N_3798);
and U4137 (N_4137,N_3719,N_3567);
nand U4138 (N_4138,N_3954,N_3681);
nor U4139 (N_4139,N_3740,N_3806);
nand U4140 (N_4140,N_3763,N_3590);
nand U4141 (N_4141,N_3827,N_3859);
and U4142 (N_4142,N_3685,N_3953);
nand U4143 (N_4143,N_3855,N_3575);
and U4144 (N_4144,N_3979,N_3566);
or U4145 (N_4145,N_3794,N_3709);
nand U4146 (N_4146,N_3512,N_3627);
and U4147 (N_4147,N_3933,N_3987);
and U4148 (N_4148,N_3854,N_3901);
and U4149 (N_4149,N_3700,N_3708);
or U4150 (N_4150,N_3502,N_3701);
nand U4151 (N_4151,N_3580,N_3657);
nor U4152 (N_4152,N_3728,N_3718);
nand U4153 (N_4153,N_3739,N_3713);
nor U4154 (N_4154,N_3503,N_3771);
or U4155 (N_4155,N_3662,N_3909);
nand U4156 (N_4156,N_3848,N_3747);
nor U4157 (N_4157,N_3946,N_3686);
nand U4158 (N_4158,N_3521,N_3519);
nor U4159 (N_4159,N_3714,N_3637);
nor U4160 (N_4160,N_3911,N_3824);
and U4161 (N_4161,N_3653,N_3673);
and U4162 (N_4162,N_3683,N_3898);
nand U4163 (N_4163,N_3777,N_3921);
or U4164 (N_4164,N_3547,N_3612);
nand U4165 (N_4165,N_3636,N_3929);
nor U4166 (N_4166,N_3980,N_3753);
nor U4167 (N_4167,N_3644,N_3666);
nand U4168 (N_4168,N_3965,N_3506);
or U4169 (N_4169,N_3990,N_3818);
nand U4170 (N_4170,N_3896,N_3581);
and U4171 (N_4171,N_3692,N_3816);
or U4172 (N_4172,N_3707,N_3880);
nor U4173 (N_4173,N_3945,N_3522);
and U4174 (N_4174,N_3592,N_3887);
or U4175 (N_4175,N_3731,N_3977);
or U4176 (N_4176,N_3875,N_3638);
nor U4177 (N_4177,N_3663,N_3971);
and U4178 (N_4178,N_3574,N_3660);
nand U4179 (N_4179,N_3861,N_3927);
nand U4180 (N_4180,N_3772,N_3532);
and U4181 (N_4181,N_3889,N_3915);
or U4182 (N_4182,N_3752,N_3565);
nor U4183 (N_4183,N_3675,N_3938);
and U4184 (N_4184,N_3813,N_3640);
nand U4185 (N_4185,N_3797,N_3857);
nand U4186 (N_4186,N_3568,N_3885);
or U4187 (N_4187,N_3509,N_3970);
nor U4188 (N_4188,N_3810,N_3513);
or U4189 (N_4189,N_3561,N_3978);
nor U4190 (N_4190,N_3745,N_3925);
nor U4191 (N_4191,N_3605,N_3617);
or U4192 (N_4192,N_3511,N_3528);
or U4193 (N_4193,N_3822,N_3730);
and U4194 (N_4194,N_3866,N_3579);
nand U4195 (N_4195,N_3501,N_3948);
and U4196 (N_4196,N_3881,N_3613);
and U4197 (N_4197,N_3770,N_3726);
nor U4198 (N_4198,N_3743,N_3646);
nor U4199 (N_4199,N_3630,N_3913);
and U4200 (N_4200,N_3802,N_3809);
and U4201 (N_4201,N_3515,N_3800);
nor U4202 (N_4202,N_3983,N_3603);
and U4203 (N_4203,N_3618,N_3843);
nor U4204 (N_4204,N_3974,N_3957);
and U4205 (N_4205,N_3667,N_3703);
or U4206 (N_4206,N_3839,N_3828);
nor U4207 (N_4207,N_3623,N_3659);
or U4208 (N_4208,N_3544,N_3860);
xor U4209 (N_4209,N_3517,N_3996);
and U4210 (N_4210,N_3594,N_3781);
and U4211 (N_4211,N_3742,N_3599);
nand U4212 (N_4212,N_3910,N_3720);
and U4213 (N_4213,N_3868,N_3893);
nor U4214 (N_4214,N_3550,N_3976);
nor U4215 (N_4215,N_3894,N_3650);
or U4216 (N_4216,N_3687,N_3779);
and U4217 (N_4217,N_3873,N_3776);
nor U4218 (N_4218,N_3790,N_3832);
or U4219 (N_4219,N_3500,N_3625);
or U4220 (N_4220,N_3523,N_3610);
xor U4221 (N_4221,N_3830,N_3769);
and U4222 (N_4222,N_3964,N_3634);
nand U4223 (N_4223,N_3956,N_3738);
or U4224 (N_4224,N_3628,N_3533);
and U4225 (N_4225,N_3926,N_3755);
nand U4226 (N_4226,N_3872,N_3729);
and U4227 (N_4227,N_3795,N_3966);
nand U4228 (N_4228,N_3808,N_3773);
and U4229 (N_4229,N_3672,N_3676);
or U4230 (N_4230,N_3587,N_3546);
nor U4231 (N_4231,N_3542,N_3912);
and U4232 (N_4232,N_3604,N_3952);
nor U4233 (N_4233,N_3812,N_3801);
or U4234 (N_4234,N_3652,N_3837);
nor U4235 (N_4235,N_3902,N_3951);
and U4236 (N_4236,N_3691,N_3882);
or U4237 (N_4237,N_3611,N_3803);
or U4238 (N_4238,N_3862,N_3908);
nand U4239 (N_4239,N_3838,N_3928);
and U4240 (N_4240,N_3624,N_3867);
nand U4241 (N_4241,N_3814,N_3939);
and U4242 (N_4242,N_3619,N_3874);
or U4243 (N_4243,N_3696,N_3582);
nor U4244 (N_4244,N_3699,N_3711);
and U4245 (N_4245,N_3586,N_3991);
or U4246 (N_4246,N_3529,N_3850);
or U4247 (N_4247,N_3677,N_3936);
nand U4248 (N_4248,N_3871,N_3900);
or U4249 (N_4249,N_3694,N_3891);
and U4250 (N_4250,N_3881,N_3855);
nand U4251 (N_4251,N_3555,N_3638);
and U4252 (N_4252,N_3619,N_3739);
and U4253 (N_4253,N_3651,N_3763);
nor U4254 (N_4254,N_3614,N_3506);
nand U4255 (N_4255,N_3791,N_3805);
or U4256 (N_4256,N_3750,N_3795);
nand U4257 (N_4257,N_3628,N_3830);
nand U4258 (N_4258,N_3909,N_3661);
and U4259 (N_4259,N_3745,N_3597);
nor U4260 (N_4260,N_3672,N_3753);
or U4261 (N_4261,N_3977,N_3862);
or U4262 (N_4262,N_3832,N_3500);
nand U4263 (N_4263,N_3891,N_3756);
nand U4264 (N_4264,N_3831,N_3501);
nand U4265 (N_4265,N_3637,N_3540);
or U4266 (N_4266,N_3689,N_3551);
or U4267 (N_4267,N_3889,N_3710);
nand U4268 (N_4268,N_3750,N_3950);
nand U4269 (N_4269,N_3812,N_3529);
and U4270 (N_4270,N_3627,N_3539);
and U4271 (N_4271,N_3838,N_3778);
and U4272 (N_4272,N_3957,N_3777);
nor U4273 (N_4273,N_3793,N_3910);
or U4274 (N_4274,N_3681,N_3875);
nor U4275 (N_4275,N_3913,N_3941);
nand U4276 (N_4276,N_3572,N_3864);
nand U4277 (N_4277,N_3628,N_3673);
or U4278 (N_4278,N_3914,N_3645);
nor U4279 (N_4279,N_3597,N_3541);
and U4280 (N_4280,N_3915,N_3570);
xnor U4281 (N_4281,N_3737,N_3846);
nor U4282 (N_4282,N_3757,N_3637);
nand U4283 (N_4283,N_3612,N_3542);
or U4284 (N_4284,N_3525,N_3829);
nor U4285 (N_4285,N_3842,N_3952);
nand U4286 (N_4286,N_3713,N_3944);
or U4287 (N_4287,N_3566,N_3732);
nor U4288 (N_4288,N_3549,N_3784);
or U4289 (N_4289,N_3606,N_3747);
nor U4290 (N_4290,N_3888,N_3957);
and U4291 (N_4291,N_3758,N_3696);
or U4292 (N_4292,N_3963,N_3826);
and U4293 (N_4293,N_3620,N_3813);
nand U4294 (N_4294,N_3533,N_3734);
xor U4295 (N_4295,N_3715,N_3593);
or U4296 (N_4296,N_3965,N_3773);
nor U4297 (N_4297,N_3858,N_3891);
and U4298 (N_4298,N_3971,N_3732);
nor U4299 (N_4299,N_3966,N_3689);
and U4300 (N_4300,N_3502,N_3915);
nand U4301 (N_4301,N_3877,N_3756);
and U4302 (N_4302,N_3744,N_3662);
or U4303 (N_4303,N_3657,N_3732);
nor U4304 (N_4304,N_3581,N_3518);
nor U4305 (N_4305,N_3564,N_3997);
or U4306 (N_4306,N_3948,N_3630);
and U4307 (N_4307,N_3610,N_3759);
or U4308 (N_4308,N_3822,N_3946);
and U4309 (N_4309,N_3845,N_3934);
and U4310 (N_4310,N_3863,N_3687);
or U4311 (N_4311,N_3575,N_3951);
or U4312 (N_4312,N_3895,N_3602);
nand U4313 (N_4313,N_3884,N_3829);
nand U4314 (N_4314,N_3929,N_3539);
nand U4315 (N_4315,N_3963,N_3503);
or U4316 (N_4316,N_3773,N_3525);
nor U4317 (N_4317,N_3752,N_3822);
or U4318 (N_4318,N_3687,N_3608);
and U4319 (N_4319,N_3691,N_3957);
and U4320 (N_4320,N_3505,N_3739);
nor U4321 (N_4321,N_3510,N_3751);
and U4322 (N_4322,N_3870,N_3845);
or U4323 (N_4323,N_3660,N_3705);
or U4324 (N_4324,N_3526,N_3597);
or U4325 (N_4325,N_3767,N_3871);
or U4326 (N_4326,N_3767,N_3534);
nand U4327 (N_4327,N_3611,N_3846);
nor U4328 (N_4328,N_3611,N_3671);
nand U4329 (N_4329,N_3554,N_3963);
nand U4330 (N_4330,N_3569,N_3702);
nand U4331 (N_4331,N_3843,N_3795);
nor U4332 (N_4332,N_3715,N_3989);
nor U4333 (N_4333,N_3561,N_3695);
and U4334 (N_4334,N_3641,N_3524);
nor U4335 (N_4335,N_3830,N_3956);
or U4336 (N_4336,N_3644,N_3854);
nand U4337 (N_4337,N_3840,N_3933);
nand U4338 (N_4338,N_3850,N_3856);
and U4339 (N_4339,N_3581,N_3547);
or U4340 (N_4340,N_3931,N_3773);
or U4341 (N_4341,N_3556,N_3543);
and U4342 (N_4342,N_3793,N_3906);
and U4343 (N_4343,N_3670,N_3957);
and U4344 (N_4344,N_3510,N_3987);
and U4345 (N_4345,N_3858,N_3868);
nand U4346 (N_4346,N_3509,N_3592);
or U4347 (N_4347,N_3557,N_3970);
or U4348 (N_4348,N_3901,N_3707);
or U4349 (N_4349,N_3828,N_3690);
and U4350 (N_4350,N_3763,N_3945);
nor U4351 (N_4351,N_3624,N_3797);
nand U4352 (N_4352,N_3952,N_3955);
nand U4353 (N_4353,N_3509,N_3945);
nor U4354 (N_4354,N_3988,N_3847);
nor U4355 (N_4355,N_3851,N_3984);
nor U4356 (N_4356,N_3761,N_3626);
and U4357 (N_4357,N_3516,N_3941);
or U4358 (N_4358,N_3693,N_3617);
and U4359 (N_4359,N_3603,N_3547);
nor U4360 (N_4360,N_3739,N_3994);
and U4361 (N_4361,N_3570,N_3866);
and U4362 (N_4362,N_3720,N_3878);
and U4363 (N_4363,N_3788,N_3638);
nand U4364 (N_4364,N_3595,N_3767);
and U4365 (N_4365,N_3977,N_3627);
or U4366 (N_4366,N_3959,N_3682);
or U4367 (N_4367,N_3957,N_3840);
nand U4368 (N_4368,N_3572,N_3508);
and U4369 (N_4369,N_3598,N_3588);
and U4370 (N_4370,N_3872,N_3945);
xor U4371 (N_4371,N_3963,N_3745);
or U4372 (N_4372,N_3648,N_3630);
nand U4373 (N_4373,N_3522,N_3905);
or U4374 (N_4374,N_3532,N_3862);
or U4375 (N_4375,N_3941,N_3852);
and U4376 (N_4376,N_3772,N_3858);
and U4377 (N_4377,N_3857,N_3659);
and U4378 (N_4378,N_3719,N_3753);
or U4379 (N_4379,N_3638,N_3879);
and U4380 (N_4380,N_3924,N_3659);
nand U4381 (N_4381,N_3988,N_3998);
nor U4382 (N_4382,N_3524,N_3622);
nor U4383 (N_4383,N_3758,N_3568);
and U4384 (N_4384,N_3507,N_3860);
or U4385 (N_4385,N_3664,N_3837);
and U4386 (N_4386,N_3950,N_3996);
nor U4387 (N_4387,N_3713,N_3678);
nor U4388 (N_4388,N_3631,N_3954);
nor U4389 (N_4389,N_3765,N_3519);
nor U4390 (N_4390,N_3677,N_3986);
or U4391 (N_4391,N_3624,N_3664);
and U4392 (N_4392,N_3674,N_3809);
or U4393 (N_4393,N_3986,N_3990);
or U4394 (N_4394,N_3541,N_3859);
nor U4395 (N_4395,N_3979,N_3686);
xor U4396 (N_4396,N_3882,N_3889);
and U4397 (N_4397,N_3530,N_3652);
xor U4398 (N_4398,N_3594,N_3747);
and U4399 (N_4399,N_3817,N_3971);
nand U4400 (N_4400,N_3779,N_3515);
and U4401 (N_4401,N_3632,N_3716);
and U4402 (N_4402,N_3561,N_3954);
and U4403 (N_4403,N_3986,N_3512);
nor U4404 (N_4404,N_3846,N_3703);
or U4405 (N_4405,N_3677,N_3780);
nand U4406 (N_4406,N_3525,N_3801);
nand U4407 (N_4407,N_3976,N_3524);
or U4408 (N_4408,N_3941,N_3819);
nor U4409 (N_4409,N_3897,N_3801);
or U4410 (N_4410,N_3674,N_3511);
and U4411 (N_4411,N_3550,N_3598);
nand U4412 (N_4412,N_3521,N_3850);
and U4413 (N_4413,N_3888,N_3864);
or U4414 (N_4414,N_3997,N_3609);
nand U4415 (N_4415,N_3603,N_3539);
nor U4416 (N_4416,N_3648,N_3777);
nor U4417 (N_4417,N_3901,N_3841);
nor U4418 (N_4418,N_3854,N_3827);
nor U4419 (N_4419,N_3642,N_3626);
nor U4420 (N_4420,N_3603,N_3559);
nor U4421 (N_4421,N_3567,N_3620);
nand U4422 (N_4422,N_3923,N_3590);
or U4423 (N_4423,N_3910,N_3832);
nand U4424 (N_4424,N_3510,N_3967);
or U4425 (N_4425,N_3522,N_3671);
nand U4426 (N_4426,N_3900,N_3929);
and U4427 (N_4427,N_3856,N_3611);
and U4428 (N_4428,N_3795,N_3514);
or U4429 (N_4429,N_3895,N_3509);
and U4430 (N_4430,N_3696,N_3843);
nor U4431 (N_4431,N_3617,N_3930);
and U4432 (N_4432,N_3737,N_3866);
and U4433 (N_4433,N_3993,N_3786);
nor U4434 (N_4434,N_3521,N_3841);
or U4435 (N_4435,N_3503,N_3836);
and U4436 (N_4436,N_3556,N_3746);
nand U4437 (N_4437,N_3842,N_3805);
or U4438 (N_4438,N_3878,N_3659);
nor U4439 (N_4439,N_3526,N_3707);
and U4440 (N_4440,N_3914,N_3977);
or U4441 (N_4441,N_3933,N_3754);
nor U4442 (N_4442,N_3793,N_3755);
and U4443 (N_4443,N_3660,N_3980);
nand U4444 (N_4444,N_3680,N_3526);
or U4445 (N_4445,N_3778,N_3988);
nand U4446 (N_4446,N_3670,N_3595);
nor U4447 (N_4447,N_3679,N_3657);
nand U4448 (N_4448,N_3808,N_3834);
and U4449 (N_4449,N_3547,N_3664);
nand U4450 (N_4450,N_3936,N_3799);
nor U4451 (N_4451,N_3662,N_3749);
or U4452 (N_4452,N_3528,N_3809);
nor U4453 (N_4453,N_3718,N_3963);
nand U4454 (N_4454,N_3812,N_3922);
or U4455 (N_4455,N_3815,N_3809);
nand U4456 (N_4456,N_3964,N_3613);
nand U4457 (N_4457,N_3758,N_3503);
nand U4458 (N_4458,N_3768,N_3939);
nand U4459 (N_4459,N_3506,N_3891);
nor U4460 (N_4460,N_3720,N_3581);
or U4461 (N_4461,N_3684,N_3886);
nor U4462 (N_4462,N_3594,N_3871);
nand U4463 (N_4463,N_3587,N_3974);
nor U4464 (N_4464,N_3788,N_3542);
nor U4465 (N_4465,N_3957,N_3770);
and U4466 (N_4466,N_3895,N_3700);
or U4467 (N_4467,N_3732,N_3570);
nor U4468 (N_4468,N_3688,N_3738);
or U4469 (N_4469,N_3862,N_3597);
nand U4470 (N_4470,N_3600,N_3576);
nand U4471 (N_4471,N_3723,N_3804);
nand U4472 (N_4472,N_3986,N_3517);
nor U4473 (N_4473,N_3546,N_3873);
or U4474 (N_4474,N_3653,N_3576);
and U4475 (N_4475,N_3893,N_3706);
or U4476 (N_4476,N_3555,N_3878);
and U4477 (N_4477,N_3843,N_3995);
nand U4478 (N_4478,N_3752,N_3756);
nand U4479 (N_4479,N_3533,N_3690);
or U4480 (N_4480,N_3958,N_3655);
nand U4481 (N_4481,N_3528,N_3934);
xor U4482 (N_4482,N_3802,N_3704);
nand U4483 (N_4483,N_3925,N_3978);
nand U4484 (N_4484,N_3851,N_3844);
nand U4485 (N_4485,N_3765,N_3897);
nor U4486 (N_4486,N_3629,N_3581);
or U4487 (N_4487,N_3608,N_3936);
and U4488 (N_4488,N_3532,N_3552);
and U4489 (N_4489,N_3680,N_3545);
nor U4490 (N_4490,N_3979,N_3939);
nor U4491 (N_4491,N_3861,N_3642);
and U4492 (N_4492,N_3841,N_3554);
or U4493 (N_4493,N_3729,N_3532);
xnor U4494 (N_4494,N_3994,N_3981);
and U4495 (N_4495,N_3976,N_3804);
or U4496 (N_4496,N_3556,N_3565);
nand U4497 (N_4497,N_3582,N_3702);
nor U4498 (N_4498,N_3815,N_3755);
and U4499 (N_4499,N_3786,N_3929);
nand U4500 (N_4500,N_4007,N_4273);
nand U4501 (N_4501,N_4039,N_4049);
nand U4502 (N_4502,N_4401,N_4416);
and U4503 (N_4503,N_4335,N_4323);
or U4504 (N_4504,N_4241,N_4358);
and U4505 (N_4505,N_4352,N_4446);
and U4506 (N_4506,N_4353,N_4231);
and U4507 (N_4507,N_4002,N_4332);
and U4508 (N_4508,N_4220,N_4208);
and U4509 (N_4509,N_4479,N_4067);
nor U4510 (N_4510,N_4382,N_4414);
and U4511 (N_4511,N_4019,N_4480);
nand U4512 (N_4512,N_4020,N_4330);
and U4513 (N_4513,N_4272,N_4177);
nand U4514 (N_4514,N_4126,N_4334);
nand U4515 (N_4515,N_4322,N_4472);
nand U4516 (N_4516,N_4439,N_4034);
and U4517 (N_4517,N_4193,N_4143);
or U4518 (N_4518,N_4174,N_4035);
and U4519 (N_4519,N_4385,N_4054);
or U4520 (N_4520,N_4190,N_4417);
and U4521 (N_4521,N_4235,N_4453);
and U4522 (N_4522,N_4087,N_4394);
and U4523 (N_4523,N_4074,N_4121);
nor U4524 (N_4524,N_4469,N_4141);
nand U4525 (N_4525,N_4227,N_4349);
and U4526 (N_4526,N_4366,N_4304);
nand U4527 (N_4527,N_4425,N_4102);
and U4528 (N_4528,N_4426,N_4159);
or U4529 (N_4529,N_4259,N_4195);
and U4530 (N_4530,N_4355,N_4176);
xnor U4531 (N_4531,N_4033,N_4068);
or U4532 (N_4532,N_4093,N_4085);
nand U4533 (N_4533,N_4058,N_4015);
and U4534 (N_4534,N_4199,N_4045);
nor U4535 (N_4535,N_4278,N_4247);
nor U4536 (N_4536,N_4456,N_4402);
or U4537 (N_4537,N_4254,N_4044);
nand U4538 (N_4538,N_4265,N_4441);
and U4539 (N_4539,N_4282,N_4269);
or U4540 (N_4540,N_4092,N_4160);
nor U4541 (N_4541,N_4233,N_4270);
and U4542 (N_4542,N_4229,N_4368);
nor U4543 (N_4543,N_4369,N_4042);
nor U4544 (N_4544,N_4072,N_4413);
and U4545 (N_4545,N_4228,N_4482);
nand U4546 (N_4546,N_4277,N_4154);
nor U4547 (N_4547,N_4333,N_4292);
and U4548 (N_4548,N_4040,N_4225);
nor U4549 (N_4549,N_4476,N_4217);
nor U4550 (N_4550,N_4161,N_4065);
nand U4551 (N_4551,N_4314,N_4100);
nor U4552 (N_4552,N_4418,N_4279);
nand U4553 (N_4553,N_4041,N_4274);
nor U4554 (N_4554,N_4275,N_4169);
nor U4555 (N_4555,N_4116,N_4242);
nor U4556 (N_4556,N_4250,N_4158);
nand U4557 (N_4557,N_4205,N_4427);
nand U4558 (N_4558,N_4184,N_4059);
nor U4559 (N_4559,N_4080,N_4108);
nand U4560 (N_4560,N_4130,N_4120);
nor U4561 (N_4561,N_4050,N_4471);
and U4562 (N_4562,N_4110,N_4263);
or U4563 (N_4563,N_4462,N_4051);
nand U4564 (N_4564,N_4447,N_4389);
nor U4565 (N_4565,N_4290,N_4434);
or U4566 (N_4566,N_4312,N_4474);
or U4567 (N_4567,N_4477,N_4098);
nand U4568 (N_4568,N_4397,N_4387);
nand U4569 (N_4569,N_4128,N_4187);
nor U4570 (N_4570,N_4498,N_4201);
and U4571 (N_4571,N_4399,N_4197);
or U4572 (N_4572,N_4010,N_4112);
nor U4573 (N_4573,N_4478,N_4252);
and U4574 (N_4574,N_4094,N_4428);
and U4575 (N_4575,N_4367,N_4014);
and U4576 (N_4576,N_4057,N_4483);
nand U4577 (N_4577,N_4357,N_4203);
nand U4578 (N_4578,N_4200,N_4324);
nand U4579 (N_4579,N_4156,N_4144);
or U4580 (N_4580,N_4155,N_4489);
nand U4581 (N_4581,N_4244,N_4013);
nand U4582 (N_4582,N_4029,N_4017);
and U4583 (N_4583,N_4374,N_4223);
or U4584 (N_4584,N_4097,N_4262);
nor U4585 (N_4585,N_4444,N_4056);
nand U4586 (N_4586,N_4243,N_4175);
and U4587 (N_4587,N_4379,N_4037);
nor U4588 (N_4588,N_4302,N_4255);
and U4589 (N_4589,N_4157,N_4071);
nor U4590 (N_4590,N_4211,N_4105);
nor U4591 (N_4591,N_4404,N_4099);
nand U4592 (N_4592,N_4248,N_4083);
nor U4593 (N_4593,N_4125,N_4053);
and U4594 (N_4594,N_4487,N_4329);
or U4595 (N_4595,N_4484,N_4343);
nor U4596 (N_4596,N_4025,N_4189);
nor U4597 (N_4597,N_4179,N_4308);
nand U4598 (N_4598,N_4468,N_4070);
nor U4599 (N_4599,N_4463,N_4342);
nor U4600 (N_4600,N_4490,N_4060);
nand U4601 (N_4601,N_4152,N_4359);
and U4602 (N_4602,N_4403,N_4104);
nand U4603 (N_4603,N_4214,N_4412);
nand U4604 (N_4604,N_4151,N_4305);
xnor U4605 (N_4605,N_4137,N_4436);
nor U4606 (N_4606,N_4139,N_4069);
or U4607 (N_4607,N_4351,N_4240);
or U4608 (N_4608,N_4493,N_4153);
nor U4609 (N_4609,N_4488,N_4146);
xnor U4610 (N_4610,N_4295,N_4318);
nor U4611 (N_4611,N_4400,N_4192);
and U4612 (N_4612,N_4030,N_4222);
xnor U4613 (N_4613,N_4196,N_4321);
and U4614 (N_4614,N_4317,N_4260);
and U4615 (N_4615,N_4331,N_4454);
nand U4616 (N_4616,N_4234,N_4089);
or U4617 (N_4617,N_4285,N_4380);
nor U4618 (N_4618,N_4003,N_4445);
nor U4619 (N_4619,N_4491,N_4396);
and U4620 (N_4620,N_4362,N_4170);
nand U4621 (N_4621,N_4264,N_4494);
nor U4622 (N_4622,N_4073,N_4496);
or U4623 (N_4623,N_4344,N_4319);
nand U4624 (N_4624,N_4230,N_4326);
or U4625 (N_4625,N_4415,N_4164);
xnor U4626 (N_4626,N_4226,N_4076);
nor U4627 (N_4627,N_4466,N_4119);
and U4628 (N_4628,N_4364,N_4027);
and U4629 (N_4629,N_4420,N_4109);
nand U4630 (N_4630,N_4470,N_4341);
nand U4631 (N_4631,N_4113,N_4467);
nand U4632 (N_4632,N_4438,N_4320);
or U4633 (N_4633,N_4063,N_4009);
nand U4634 (N_4634,N_4188,N_4210);
nor U4635 (N_4635,N_4450,N_4061);
or U4636 (N_4636,N_4457,N_4309);
or U4637 (N_4637,N_4219,N_4107);
and U4638 (N_4638,N_4303,N_4082);
and U4639 (N_4639,N_4392,N_4306);
or U4640 (N_4640,N_4202,N_4345);
nand U4641 (N_4641,N_4300,N_4391);
or U4642 (N_4642,N_4132,N_4168);
nor U4643 (N_4643,N_4216,N_4361);
nor U4644 (N_4644,N_4348,N_4249);
or U4645 (N_4645,N_4142,N_4307);
nor U4646 (N_4646,N_4461,N_4129);
or U4647 (N_4647,N_4442,N_4424);
or U4648 (N_4648,N_4298,N_4464);
and U4649 (N_4649,N_4451,N_4390);
nor U4650 (N_4650,N_4339,N_4232);
and U4651 (N_4651,N_4111,N_4409);
nand U4652 (N_4652,N_4291,N_4328);
or U4653 (N_4653,N_4492,N_4499);
nor U4654 (N_4654,N_4360,N_4388);
or U4655 (N_4655,N_4384,N_4336);
or U4656 (N_4656,N_4131,N_4149);
or U4657 (N_4657,N_4432,N_4383);
or U4658 (N_4658,N_4101,N_4431);
and U4659 (N_4659,N_4117,N_4410);
or U4660 (N_4660,N_4327,N_4147);
nand U4661 (N_4661,N_4036,N_4148);
and U4662 (N_4662,N_4062,N_4221);
and U4663 (N_4663,N_4018,N_4140);
or U4664 (N_4664,N_4088,N_4091);
nor U4665 (N_4665,N_4411,N_4204);
and U4666 (N_4666,N_4354,N_4251);
or U4667 (N_4667,N_4378,N_4377);
nor U4668 (N_4668,N_4449,N_4261);
nand U4669 (N_4669,N_4038,N_4114);
nor U4670 (N_4670,N_4381,N_4180);
nand U4671 (N_4671,N_4408,N_4268);
or U4672 (N_4672,N_4310,N_4165);
and U4673 (N_4673,N_4266,N_4315);
or U4674 (N_4674,N_4347,N_4173);
nor U4675 (N_4675,N_4256,N_4271);
and U4676 (N_4676,N_4458,N_4372);
or U4677 (N_4677,N_4301,N_4122);
nor U4678 (N_4678,N_4455,N_4055);
nand U4679 (N_4679,N_4398,N_4134);
nand U4680 (N_4680,N_4473,N_4150);
nand U4681 (N_4681,N_4001,N_4375);
nand U4682 (N_4682,N_4284,N_4365);
or U4683 (N_4683,N_4376,N_4437);
nand U4684 (N_4684,N_4135,N_4005);
or U4685 (N_4685,N_4452,N_4136);
nor U4686 (N_4686,N_4024,N_4386);
or U4687 (N_4687,N_4253,N_4198);
or U4688 (N_4688,N_4166,N_4224);
or U4689 (N_4689,N_4337,N_4340);
nand U4690 (N_4690,N_4206,N_4448);
or U4691 (N_4691,N_4373,N_4346);
and U4692 (N_4692,N_4172,N_4423);
nand U4693 (N_4693,N_4371,N_4276);
or U4694 (N_4694,N_4239,N_4429);
xnor U4695 (N_4695,N_4460,N_4194);
and U4696 (N_4696,N_4021,N_4026);
or U4697 (N_4697,N_4103,N_4350);
or U4698 (N_4698,N_4338,N_4075);
or U4699 (N_4699,N_4213,N_4052);
and U4700 (N_4700,N_4422,N_4212);
nand U4701 (N_4701,N_4430,N_4023);
or U4702 (N_4702,N_4363,N_4012);
and U4703 (N_4703,N_4405,N_4011);
and U4704 (N_4704,N_4433,N_4419);
nor U4705 (N_4705,N_4095,N_4465);
xnor U4706 (N_4706,N_4115,N_4182);
nor U4707 (N_4707,N_4407,N_4181);
or U4708 (N_4708,N_4481,N_4299);
nor U4709 (N_4709,N_4245,N_4123);
and U4710 (N_4710,N_4495,N_4004);
nor U4711 (N_4711,N_4293,N_4475);
or U4712 (N_4712,N_4163,N_4325);
or U4713 (N_4713,N_4296,N_4167);
or U4714 (N_4714,N_4106,N_4162);
or U4715 (N_4715,N_4287,N_4000);
nor U4716 (N_4716,N_4046,N_4288);
nor U4717 (N_4717,N_4031,N_4145);
or U4718 (N_4718,N_4443,N_4280);
nand U4719 (N_4719,N_4238,N_4138);
and U4720 (N_4720,N_4079,N_4171);
nor U4721 (N_4721,N_4133,N_4090);
nand U4722 (N_4722,N_4246,N_4406);
nor U4723 (N_4723,N_4008,N_4078);
nor U4724 (N_4724,N_4022,N_4313);
nand U4725 (N_4725,N_4258,N_4191);
and U4726 (N_4726,N_4048,N_4066);
nand U4727 (N_4727,N_4006,N_4297);
nand U4728 (N_4728,N_4267,N_4257);
nand U4729 (N_4729,N_4497,N_4356);
nor U4730 (N_4730,N_4370,N_4316);
nand U4731 (N_4731,N_4185,N_4032);
nor U4732 (N_4732,N_4283,N_4178);
nand U4733 (N_4733,N_4311,N_4118);
nand U4734 (N_4734,N_4096,N_4084);
nor U4735 (N_4735,N_4028,N_4127);
or U4736 (N_4736,N_4081,N_4047);
nand U4737 (N_4737,N_4421,N_4237);
or U4738 (N_4738,N_4393,N_4064);
and U4739 (N_4739,N_4486,N_4215);
and U4740 (N_4740,N_4435,N_4086);
or U4741 (N_4741,N_4218,N_4281);
or U4742 (N_4742,N_4440,N_4207);
and U4743 (N_4743,N_4186,N_4043);
or U4744 (N_4744,N_4016,N_4183);
and U4745 (N_4745,N_4236,N_4124);
or U4746 (N_4746,N_4077,N_4459);
or U4747 (N_4747,N_4294,N_4395);
or U4748 (N_4748,N_4485,N_4209);
or U4749 (N_4749,N_4286,N_4289);
nand U4750 (N_4750,N_4375,N_4306);
xor U4751 (N_4751,N_4332,N_4263);
nand U4752 (N_4752,N_4365,N_4327);
or U4753 (N_4753,N_4047,N_4045);
nor U4754 (N_4754,N_4472,N_4465);
and U4755 (N_4755,N_4281,N_4260);
or U4756 (N_4756,N_4149,N_4199);
nand U4757 (N_4757,N_4182,N_4210);
or U4758 (N_4758,N_4357,N_4363);
nor U4759 (N_4759,N_4186,N_4229);
and U4760 (N_4760,N_4209,N_4337);
or U4761 (N_4761,N_4398,N_4183);
nand U4762 (N_4762,N_4109,N_4276);
nor U4763 (N_4763,N_4224,N_4154);
nand U4764 (N_4764,N_4212,N_4125);
nand U4765 (N_4765,N_4273,N_4349);
nor U4766 (N_4766,N_4336,N_4204);
and U4767 (N_4767,N_4436,N_4006);
nor U4768 (N_4768,N_4197,N_4464);
or U4769 (N_4769,N_4286,N_4306);
xnor U4770 (N_4770,N_4367,N_4030);
nand U4771 (N_4771,N_4187,N_4314);
nor U4772 (N_4772,N_4378,N_4164);
and U4773 (N_4773,N_4228,N_4261);
and U4774 (N_4774,N_4048,N_4195);
nor U4775 (N_4775,N_4149,N_4418);
nor U4776 (N_4776,N_4006,N_4015);
nand U4777 (N_4777,N_4208,N_4484);
and U4778 (N_4778,N_4199,N_4364);
or U4779 (N_4779,N_4240,N_4376);
nand U4780 (N_4780,N_4299,N_4471);
nor U4781 (N_4781,N_4170,N_4145);
and U4782 (N_4782,N_4112,N_4348);
and U4783 (N_4783,N_4372,N_4312);
or U4784 (N_4784,N_4157,N_4373);
nor U4785 (N_4785,N_4120,N_4395);
and U4786 (N_4786,N_4350,N_4026);
nand U4787 (N_4787,N_4373,N_4449);
and U4788 (N_4788,N_4194,N_4170);
or U4789 (N_4789,N_4113,N_4189);
or U4790 (N_4790,N_4310,N_4097);
or U4791 (N_4791,N_4109,N_4016);
or U4792 (N_4792,N_4039,N_4078);
or U4793 (N_4793,N_4042,N_4095);
nor U4794 (N_4794,N_4492,N_4268);
nor U4795 (N_4795,N_4133,N_4490);
nor U4796 (N_4796,N_4073,N_4334);
or U4797 (N_4797,N_4018,N_4097);
and U4798 (N_4798,N_4187,N_4494);
or U4799 (N_4799,N_4251,N_4318);
nor U4800 (N_4800,N_4422,N_4441);
and U4801 (N_4801,N_4326,N_4345);
or U4802 (N_4802,N_4216,N_4341);
nand U4803 (N_4803,N_4371,N_4166);
nand U4804 (N_4804,N_4073,N_4217);
nor U4805 (N_4805,N_4020,N_4302);
nor U4806 (N_4806,N_4335,N_4235);
or U4807 (N_4807,N_4221,N_4163);
or U4808 (N_4808,N_4109,N_4345);
or U4809 (N_4809,N_4030,N_4086);
or U4810 (N_4810,N_4083,N_4271);
nor U4811 (N_4811,N_4105,N_4379);
or U4812 (N_4812,N_4105,N_4015);
nand U4813 (N_4813,N_4048,N_4253);
nor U4814 (N_4814,N_4499,N_4135);
and U4815 (N_4815,N_4307,N_4448);
nand U4816 (N_4816,N_4174,N_4292);
or U4817 (N_4817,N_4393,N_4065);
nor U4818 (N_4818,N_4022,N_4029);
nor U4819 (N_4819,N_4185,N_4471);
or U4820 (N_4820,N_4168,N_4333);
and U4821 (N_4821,N_4157,N_4152);
nand U4822 (N_4822,N_4197,N_4282);
or U4823 (N_4823,N_4005,N_4283);
or U4824 (N_4824,N_4377,N_4371);
and U4825 (N_4825,N_4214,N_4212);
nand U4826 (N_4826,N_4035,N_4137);
or U4827 (N_4827,N_4116,N_4329);
and U4828 (N_4828,N_4266,N_4143);
nor U4829 (N_4829,N_4439,N_4072);
or U4830 (N_4830,N_4360,N_4447);
nor U4831 (N_4831,N_4245,N_4373);
nand U4832 (N_4832,N_4266,N_4161);
nor U4833 (N_4833,N_4424,N_4016);
nand U4834 (N_4834,N_4021,N_4398);
and U4835 (N_4835,N_4011,N_4107);
or U4836 (N_4836,N_4104,N_4000);
or U4837 (N_4837,N_4031,N_4303);
nor U4838 (N_4838,N_4330,N_4419);
and U4839 (N_4839,N_4122,N_4047);
and U4840 (N_4840,N_4148,N_4496);
or U4841 (N_4841,N_4294,N_4398);
or U4842 (N_4842,N_4451,N_4126);
nor U4843 (N_4843,N_4139,N_4058);
or U4844 (N_4844,N_4301,N_4081);
nand U4845 (N_4845,N_4180,N_4283);
and U4846 (N_4846,N_4429,N_4060);
nand U4847 (N_4847,N_4094,N_4091);
nor U4848 (N_4848,N_4494,N_4342);
nand U4849 (N_4849,N_4223,N_4190);
xnor U4850 (N_4850,N_4164,N_4194);
nand U4851 (N_4851,N_4299,N_4267);
nor U4852 (N_4852,N_4374,N_4110);
and U4853 (N_4853,N_4380,N_4317);
nand U4854 (N_4854,N_4134,N_4334);
and U4855 (N_4855,N_4295,N_4460);
nor U4856 (N_4856,N_4257,N_4078);
nand U4857 (N_4857,N_4061,N_4051);
nor U4858 (N_4858,N_4253,N_4326);
nand U4859 (N_4859,N_4379,N_4275);
nor U4860 (N_4860,N_4142,N_4453);
and U4861 (N_4861,N_4082,N_4316);
and U4862 (N_4862,N_4287,N_4326);
and U4863 (N_4863,N_4455,N_4129);
nor U4864 (N_4864,N_4476,N_4354);
nor U4865 (N_4865,N_4456,N_4263);
and U4866 (N_4866,N_4370,N_4106);
or U4867 (N_4867,N_4203,N_4195);
and U4868 (N_4868,N_4006,N_4069);
nor U4869 (N_4869,N_4453,N_4217);
and U4870 (N_4870,N_4434,N_4166);
nor U4871 (N_4871,N_4479,N_4012);
and U4872 (N_4872,N_4027,N_4220);
nand U4873 (N_4873,N_4299,N_4465);
and U4874 (N_4874,N_4158,N_4469);
and U4875 (N_4875,N_4486,N_4190);
or U4876 (N_4876,N_4082,N_4213);
nand U4877 (N_4877,N_4151,N_4145);
nor U4878 (N_4878,N_4374,N_4404);
nand U4879 (N_4879,N_4124,N_4436);
and U4880 (N_4880,N_4469,N_4165);
nand U4881 (N_4881,N_4390,N_4393);
or U4882 (N_4882,N_4416,N_4221);
or U4883 (N_4883,N_4268,N_4150);
nand U4884 (N_4884,N_4096,N_4071);
nand U4885 (N_4885,N_4049,N_4222);
or U4886 (N_4886,N_4472,N_4291);
nor U4887 (N_4887,N_4470,N_4081);
or U4888 (N_4888,N_4051,N_4085);
nand U4889 (N_4889,N_4153,N_4430);
nand U4890 (N_4890,N_4213,N_4268);
nand U4891 (N_4891,N_4008,N_4209);
or U4892 (N_4892,N_4040,N_4248);
or U4893 (N_4893,N_4495,N_4084);
or U4894 (N_4894,N_4396,N_4274);
nor U4895 (N_4895,N_4028,N_4409);
and U4896 (N_4896,N_4476,N_4383);
nor U4897 (N_4897,N_4448,N_4440);
nand U4898 (N_4898,N_4277,N_4333);
nor U4899 (N_4899,N_4062,N_4246);
nor U4900 (N_4900,N_4425,N_4417);
and U4901 (N_4901,N_4105,N_4252);
or U4902 (N_4902,N_4416,N_4439);
and U4903 (N_4903,N_4445,N_4130);
or U4904 (N_4904,N_4464,N_4378);
or U4905 (N_4905,N_4452,N_4000);
and U4906 (N_4906,N_4370,N_4062);
or U4907 (N_4907,N_4495,N_4223);
or U4908 (N_4908,N_4347,N_4384);
nand U4909 (N_4909,N_4211,N_4019);
nand U4910 (N_4910,N_4492,N_4020);
or U4911 (N_4911,N_4033,N_4463);
nor U4912 (N_4912,N_4131,N_4498);
nand U4913 (N_4913,N_4333,N_4097);
nor U4914 (N_4914,N_4355,N_4408);
or U4915 (N_4915,N_4149,N_4005);
or U4916 (N_4916,N_4300,N_4166);
or U4917 (N_4917,N_4098,N_4164);
and U4918 (N_4918,N_4120,N_4309);
or U4919 (N_4919,N_4192,N_4300);
and U4920 (N_4920,N_4364,N_4370);
and U4921 (N_4921,N_4011,N_4016);
nor U4922 (N_4922,N_4069,N_4296);
nor U4923 (N_4923,N_4205,N_4170);
nand U4924 (N_4924,N_4415,N_4309);
and U4925 (N_4925,N_4010,N_4310);
and U4926 (N_4926,N_4288,N_4345);
nor U4927 (N_4927,N_4249,N_4091);
nand U4928 (N_4928,N_4146,N_4308);
or U4929 (N_4929,N_4129,N_4146);
or U4930 (N_4930,N_4160,N_4317);
and U4931 (N_4931,N_4364,N_4212);
nor U4932 (N_4932,N_4282,N_4494);
and U4933 (N_4933,N_4376,N_4052);
nor U4934 (N_4934,N_4051,N_4291);
nand U4935 (N_4935,N_4346,N_4485);
nor U4936 (N_4936,N_4041,N_4011);
nor U4937 (N_4937,N_4233,N_4289);
or U4938 (N_4938,N_4485,N_4432);
or U4939 (N_4939,N_4387,N_4486);
or U4940 (N_4940,N_4167,N_4393);
nand U4941 (N_4941,N_4080,N_4343);
nand U4942 (N_4942,N_4459,N_4494);
or U4943 (N_4943,N_4129,N_4439);
and U4944 (N_4944,N_4145,N_4227);
or U4945 (N_4945,N_4418,N_4224);
or U4946 (N_4946,N_4094,N_4127);
nand U4947 (N_4947,N_4433,N_4393);
nand U4948 (N_4948,N_4186,N_4083);
nor U4949 (N_4949,N_4379,N_4221);
or U4950 (N_4950,N_4338,N_4284);
nand U4951 (N_4951,N_4191,N_4196);
nor U4952 (N_4952,N_4289,N_4325);
nor U4953 (N_4953,N_4409,N_4465);
or U4954 (N_4954,N_4141,N_4220);
or U4955 (N_4955,N_4125,N_4204);
or U4956 (N_4956,N_4043,N_4159);
and U4957 (N_4957,N_4168,N_4338);
or U4958 (N_4958,N_4193,N_4033);
or U4959 (N_4959,N_4250,N_4182);
nor U4960 (N_4960,N_4066,N_4155);
nand U4961 (N_4961,N_4295,N_4491);
and U4962 (N_4962,N_4053,N_4173);
nor U4963 (N_4963,N_4496,N_4396);
nand U4964 (N_4964,N_4012,N_4027);
nor U4965 (N_4965,N_4043,N_4203);
or U4966 (N_4966,N_4322,N_4036);
nand U4967 (N_4967,N_4155,N_4114);
and U4968 (N_4968,N_4425,N_4122);
nand U4969 (N_4969,N_4365,N_4063);
nor U4970 (N_4970,N_4102,N_4052);
nor U4971 (N_4971,N_4198,N_4234);
or U4972 (N_4972,N_4257,N_4445);
or U4973 (N_4973,N_4024,N_4287);
or U4974 (N_4974,N_4263,N_4155);
nor U4975 (N_4975,N_4269,N_4453);
nor U4976 (N_4976,N_4185,N_4263);
and U4977 (N_4977,N_4201,N_4082);
nor U4978 (N_4978,N_4013,N_4130);
nor U4979 (N_4979,N_4208,N_4083);
or U4980 (N_4980,N_4437,N_4003);
or U4981 (N_4981,N_4135,N_4411);
nor U4982 (N_4982,N_4101,N_4212);
and U4983 (N_4983,N_4025,N_4051);
nor U4984 (N_4984,N_4460,N_4228);
nand U4985 (N_4985,N_4199,N_4293);
nand U4986 (N_4986,N_4093,N_4176);
nand U4987 (N_4987,N_4201,N_4071);
and U4988 (N_4988,N_4339,N_4472);
or U4989 (N_4989,N_4428,N_4137);
or U4990 (N_4990,N_4368,N_4479);
nor U4991 (N_4991,N_4094,N_4222);
or U4992 (N_4992,N_4215,N_4408);
nand U4993 (N_4993,N_4402,N_4050);
and U4994 (N_4994,N_4306,N_4143);
nor U4995 (N_4995,N_4315,N_4409);
nand U4996 (N_4996,N_4474,N_4241);
nand U4997 (N_4997,N_4473,N_4298);
and U4998 (N_4998,N_4463,N_4038);
nand U4999 (N_4999,N_4111,N_4430);
and U5000 (N_5000,N_4616,N_4942);
and U5001 (N_5001,N_4660,N_4501);
and U5002 (N_5002,N_4530,N_4540);
or U5003 (N_5003,N_4598,N_4988);
and U5004 (N_5004,N_4747,N_4821);
and U5005 (N_5005,N_4930,N_4828);
or U5006 (N_5006,N_4799,N_4698);
xor U5007 (N_5007,N_4597,N_4759);
or U5008 (N_5008,N_4631,N_4771);
and U5009 (N_5009,N_4937,N_4869);
nor U5010 (N_5010,N_4628,N_4979);
or U5011 (N_5011,N_4800,N_4753);
nor U5012 (N_5012,N_4559,N_4814);
or U5013 (N_5013,N_4645,N_4613);
nand U5014 (N_5014,N_4849,N_4543);
or U5015 (N_5015,N_4641,N_4579);
and U5016 (N_5016,N_4842,N_4734);
nor U5017 (N_5017,N_4554,N_4743);
or U5018 (N_5018,N_4615,N_4907);
nand U5019 (N_5019,N_4954,N_4636);
or U5020 (N_5020,N_4866,N_4600);
or U5021 (N_5021,N_4592,N_4701);
nor U5022 (N_5022,N_4845,N_4656);
nand U5023 (N_5023,N_4726,N_4716);
and U5024 (N_5024,N_4815,N_4647);
xor U5025 (N_5025,N_4865,N_4978);
nor U5026 (N_5026,N_4620,N_4870);
or U5027 (N_5027,N_4793,N_4776);
and U5028 (N_5028,N_4603,N_4695);
nand U5029 (N_5029,N_4512,N_4707);
nand U5030 (N_5030,N_4722,N_4706);
nand U5031 (N_5031,N_4632,N_4682);
xor U5032 (N_5032,N_4503,N_4843);
xnor U5033 (N_5033,N_4638,N_4783);
nor U5034 (N_5034,N_4801,N_4609);
nand U5035 (N_5035,N_4663,N_4792);
nor U5036 (N_5036,N_4547,N_4635);
nand U5037 (N_5037,N_4898,N_4577);
and U5038 (N_5038,N_4568,N_4673);
or U5039 (N_5039,N_4982,N_4969);
or U5040 (N_5040,N_4502,N_4590);
and U5041 (N_5041,N_4816,N_4857);
nor U5042 (N_5042,N_4725,N_4583);
or U5043 (N_5043,N_4626,N_4996);
and U5044 (N_5044,N_4961,N_4888);
nor U5045 (N_5045,N_4894,N_4901);
nand U5046 (N_5046,N_4912,N_4885);
or U5047 (N_5047,N_4697,N_4710);
nor U5048 (N_5048,N_4522,N_4584);
nand U5049 (N_5049,N_4593,N_4675);
nand U5050 (N_5050,N_4708,N_4826);
nor U5051 (N_5051,N_4651,N_4691);
nand U5052 (N_5052,N_4995,N_4863);
and U5053 (N_5053,N_4694,N_4892);
and U5054 (N_5054,N_4602,N_4860);
or U5055 (N_5055,N_4830,N_4947);
and U5056 (N_5056,N_4719,N_4987);
and U5057 (N_5057,N_4891,N_4546);
nor U5058 (N_5058,N_4509,N_4606);
and U5059 (N_5059,N_4976,N_4850);
xor U5060 (N_5060,N_4764,N_4571);
nor U5061 (N_5061,N_4505,N_4856);
or U5062 (N_5062,N_4835,N_4671);
or U5063 (N_5063,N_4795,N_4745);
and U5064 (N_5064,N_4925,N_4810);
and U5065 (N_5065,N_4789,N_4871);
and U5066 (N_5066,N_4744,N_4762);
and U5067 (N_5067,N_4922,N_4855);
and U5068 (N_5068,N_4825,N_4627);
nor U5069 (N_5069,N_4882,N_4713);
nor U5070 (N_5070,N_4802,N_4629);
nor U5071 (N_5071,N_4610,N_4909);
nand U5072 (N_5072,N_4986,N_4761);
nand U5073 (N_5073,N_4643,N_4808);
nor U5074 (N_5074,N_4659,N_4720);
nand U5075 (N_5075,N_4848,N_4974);
and U5076 (N_5076,N_4665,N_4834);
and U5077 (N_5077,N_4596,N_4576);
nand U5078 (N_5078,N_4785,N_4934);
or U5079 (N_5079,N_4867,N_4536);
or U5080 (N_5080,N_4548,N_4605);
nor U5081 (N_5081,N_4562,N_4724);
or U5082 (N_5082,N_4539,N_4798);
nor U5083 (N_5083,N_4964,N_4889);
nor U5084 (N_5084,N_4965,N_4985);
nand U5085 (N_5085,N_4578,N_4607);
nor U5086 (N_5086,N_4723,N_4791);
nor U5087 (N_5087,N_4941,N_4511);
nand U5088 (N_5088,N_4787,N_4972);
nand U5089 (N_5089,N_4962,N_4840);
and U5090 (N_5090,N_4977,N_4657);
nand U5091 (N_5091,N_4526,N_4681);
nand U5092 (N_5092,N_4997,N_4847);
or U5093 (N_5093,N_4741,N_4858);
nand U5094 (N_5094,N_4939,N_4971);
or U5095 (N_5095,N_4737,N_4839);
nand U5096 (N_5096,N_4919,N_4938);
or U5097 (N_5097,N_4773,N_4959);
and U5098 (N_5098,N_4932,N_4832);
nand U5099 (N_5099,N_4960,N_4705);
nand U5100 (N_5100,N_4796,N_4900);
nand U5101 (N_5101,N_4994,N_4837);
nand U5102 (N_5102,N_4589,N_4550);
nor U5103 (N_5103,N_4684,N_4914);
nor U5104 (N_5104,N_4736,N_4558);
nand U5105 (N_5105,N_4668,N_4967);
xnor U5106 (N_5106,N_4715,N_4893);
and U5107 (N_5107,N_4742,N_4824);
xnor U5108 (N_5108,N_4926,N_4670);
nand U5109 (N_5109,N_4523,N_4696);
nor U5110 (N_5110,N_4794,N_4667);
and U5111 (N_5111,N_4945,N_4763);
and U5112 (N_5112,N_4756,N_4709);
nor U5113 (N_5113,N_4819,N_4803);
or U5114 (N_5114,N_4731,N_4879);
nand U5115 (N_5115,N_4672,N_4630);
and U5116 (N_5116,N_4999,N_4983);
and U5117 (N_5117,N_4545,N_4608);
nor U5118 (N_5118,N_4676,N_4618);
nor U5119 (N_5119,N_4507,N_4784);
or U5120 (N_5120,N_4654,N_4746);
nor U5121 (N_5121,N_4662,N_4872);
or U5122 (N_5122,N_4968,N_4781);
nor U5123 (N_5123,N_4679,N_4859);
nand U5124 (N_5124,N_4903,N_4758);
nor U5125 (N_5125,N_4683,N_4807);
nand U5126 (N_5126,N_4556,N_4527);
nand U5127 (N_5127,N_4884,N_4797);
or U5128 (N_5128,N_4658,N_4581);
nor U5129 (N_5129,N_4648,N_4544);
nand U5130 (N_5130,N_4703,N_4998);
and U5131 (N_5131,N_4680,N_4655);
nand U5132 (N_5132,N_4864,N_4990);
nor U5133 (N_5133,N_4664,N_4678);
nor U5134 (N_5134,N_4642,N_4563);
or U5135 (N_5135,N_4931,N_4686);
nor U5136 (N_5136,N_4833,N_4588);
or U5137 (N_5137,N_4873,N_4533);
or U5138 (N_5138,N_4897,N_4878);
or U5139 (N_5139,N_4693,N_4537);
nand U5140 (N_5140,N_4519,N_4923);
nand U5141 (N_5141,N_4517,N_4565);
and U5142 (N_5142,N_4951,N_4874);
nor U5143 (N_5143,N_4980,N_4779);
nand U5144 (N_5144,N_4920,N_4560);
or U5145 (N_5145,N_4886,N_4567);
nand U5146 (N_5146,N_4940,N_4838);
nor U5147 (N_5147,N_4817,N_4538);
nand U5148 (N_5148,N_4587,N_4809);
nand U5149 (N_5149,N_4625,N_4646);
nand U5150 (N_5150,N_4757,N_4529);
nand U5151 (N_5151,N_4573,N_4700);
nand U5152 (N_5152,N_4575,N_4572);
or U5153 (N_5153,N_4738,N_4570);
or U5154 (N_5154,N_4750,N_4765);
nor U5155 (N_5155,N_4521,N_4591);
nor U5156 (N_5156,N_4666,N_4692);
nand U5157 (N_5157,N_4890,N_4790);
nand U5158 (N_5158,N_4846,N_4906);
and U5159 (N_5159,N_4649,N_4580);
nor U5160 (N_5160,N_4748,N_4896);
or U5161 (N_5161,N_4624,N_4574);
nor U5162 (N_5162,N_4822,N_4729);
and U5163 (N_5163,N_4535,N_4728);
or U5164 (N_5164,N_4599,N_4929);
or U5165 (N_5165,N_4780,N_4669);
nand U5166 (N_5166,N_4514,N_4910);
and U5167 (N_5167,N_4677,N_4853);
nand U5168 (N_5168,N_4944,N_4594);
nor U5169 (N_5169,N_4955,N_4689);
nor U5170 (N_5170,N_4513,N_4927);
and U5171 (N_5171,N_4953,N_4516);
or U5172 (N_5172,N_4989,N_4504);
nor U5173 (N_5173,N_4611,N_4908);
or U5174 (N_5174,N_4862,N_4569);
xnor U5175 (N_5175,N_4688,N_4704);
nor U5176 (N_5176,N_4904,N_4751);
or U5177 (N_5177,N_4935,N_4541);
nand U5178 (N_5178,N_4690,N_4633);
and U5179 (N_5179,N_4949,N_4727);
or U5180 (N_5180,N_4924,N_4614);
nand U5181 (N_5181,N_4601,N_4827);
nand U5182 (N_5182,N_4621,N_4561);
nand U5183 (N_5183,N_4948,N_4818);
and U5184 (N_5184,N_4721,N_4739);
or U5185 (N_5185,N_4774,N_4564);
xnor U5186 (N_5186,N_4918,N_4619);
or U5187 (N_5187,N_4851,N_4531);
and U5188 (N_5188,N_4880,N_4981);
and U5189 (N_5189,N_4740,N_4687);
and U5190 (N_5190,N_4661,N_4778);
or U5191 (N_5191,N_4623,N_4844);
nand U5192 (N_5192,N_4813,N_4950);
nor U5193 (N_5193,N_4975,N_4732);
and U5194 (N_5194,N_4854,N_4902);
or U5195 (N_5195,N_4520,N_4508);
and U5196 (N_5196,N_4542,N_4993);
nor U5197 (N_5197,N_4769,N_4836);
or U5198 (N_5198,N_4717,N_4804);
or U5199 (N_5199,N_4730,N_4823);
nor U5200 (N_5200,N_4552,N_4515);
or U5201 (N_5201,N_4674,N_4956);
and U5202 (N_5202,N_4534,N_4777);
nand U5203 (N_5203,N_4852,N_4916);
nand U5204 (N_5204,N_4952,N_4555);
nor U5205 (N_5205,N_4650,N_4805);
or U5206 (N_5206,N_4752,N_4911);
and U5207 (N_5207,N_4566,N_4991);
or U5208 (N_5208,N_4877,N_4699);
or U5209 (N_5209,N_4622,N_4549);
nand U5210 (N_5210,N_4551,N_4966);
or U5211 (N_5211,N_4528,N_4524);
nor U5212 (N_5212,N_4714,N_4782);
and U5213 (N_5213,N_4766,N_4749);
or U5214 (N_5214,N_4786,N_4812);
or U5215 (N_5215,N_4506,N_4702);
and U5216 (N_5216,N_4718,N_4585);
and U5217 (N_5217,N_4604,N_4881);
or U5218 (N_5218,N_4936,N_4760);
and U5219 (N_5219,N_4943,N_4711);
xnor U5220 (N_5220,N_4640,N_4652);
or U5221 (N_5221,N_4868,N_4770);
nand U5222 (N_5222,N_4685,N_4946);
nand U5223 (N_5223,N_4733,N_4788);
nor U5224 (N_5224,N_4899,N_4595);
nand U5225 (N_5225,N_4806,N_4915);
nor U5226 (N_5226,N_4992,N_4905);
or U5227 (N_5227,N_4525,N_4754);
and U5228 (N_5228,N_4767,N_4500);
nand U5229 (N_5229,N_4518,N_4883);
nand U5230 (N_5230,N_4612,N_4653);
nor U5231 (N_5231,N_4917,N_4970);
and U5232 (N_5232,N_4984,N_4820);
nand U5233 (N_5233,N_4887,N_4921);
or U5234 (N_5234,N_4829,N_4876);
and U5235 (N_5235,N_4768,N_4532);
and U5236 (N_5236,N_4557,N_4973);
nand U5237 (N_5237,N_4775,N_4755);
or U5238 (N_5238,N_4712,N_4637);
nand U5239 (N_5239,N_4841,N_4639);
nand U5240 (N_5240,N_4510,N_4831);
xnor U5241 (N_5241,N_4957,N_4963);
or U5242 (N_5242,N_4617,N_4553);
nor U5243 (N_5243,N_4928,N_4634);
nor U5244 (N_5244,N_4582,N_4933);
and U5245 (N_5245,N_4772,N_4861);
and U5246 (N_5246,N_4958,N_4586);
and U5247 (N_5247,N_4644,N_4913);
nor U5248 (N_5248,N_4735,N_4811);
or U5249 (N_5249,N_4875,N_4895);
or U5250 (N_5250,N_4804,N_4718);
or U5251 (N_5251,N_4788,N_4686);
and U5252 (N_5252,N_4728,N_4664);
and U5253 (N_5253,N_4509,N_4517);
or U5254 (N_5254,N_4633,N_4668);
nand U5255 (N_5255,N_4672,N_4948);
nor U5256 (N_5256,N_4967,N_4553);
or U5257 (N_5257,N_4806,N_4890);
nor U5258 (N_5258,N_4944,N_4666);
or U5259 (N_5259,N_4515,N_4605);
nor U5260 (N_5260,N_4580,N_4877);
nand U5261 (N_5261,N_4538,N_4658);
nor U5262 (N_5262,N_4697,N_4539);
and U5263 (N_5263,N_4870,N_4581);
or U5264 (N_5264,N_4937,N_4800);
or U5265 (N_5265,N_4771,N_4679);
and U5266 (N_5266,N_4890,N_4670);
nand U5267 (N_5267,N_4647,N_4819);
nor U5268 (N_5268,N_4596,N_4727);
nand U5269 (N_5269,N_4856,N_4990);
nand U5270 (N_5270,N_4630,N_4840);
nor U5271 (N_5271,N_4717,N_4639);
or U5272 (N_5272,N_4786,N_4660);
nor U5273 (N_5273,N_4591,N_4779);
nor U5274 (N_5274,N_4761,N_4899);
nand U5275 (N_5275,N_4544,N_4767);
and U5276 (N_5276,N_4710,N_4855);
nor U5277 (N_5277,N_4968,N_4994);
or U5278 (N_5278,N_4756,N_4794);
or U5279 (N_5279,N_4542,N_4715);
or U5280 (N_5280,N_4652,N_4966);
nor U5281 (N_5281,N_4936,N_4636);
nand U5282 (N_5282,N_4615,N_4597);
nor U5283 (N_5283,N_4608,N_4642);
or U5284 (N_5284,N_4994,N_4690);
nand U5285 (N_5285,N_4520,N_4791);
and U5286 (N_5286,N_4689,N_4515);
xor U5287 (N_5287,N_4856,N_4871);
or U5288 (N_5288,N_4996,N_4771);
nor U5289 (N_5289,N_4933,N_4838);
nand U5290 (N_5290,N_4540,N_4964);
and U5291 (N_5291,N_4769,N_4772);
nor U5292 (N_5292,N_4520,N_4970);
nand U5293 (N_5293,N_4845,N_4922);
nor U5294 (N_5294,N_4637,N_4509);
or U5295 (N_5295,N_4524,N_4523);
nor U5296 (N_5296,N_4774,N_4957);
or U5297 (N_5297,N_4562,N_4983);
or U5298 (N_5298,N_4891,N_4709);
or U5299 (N_5299,N_4704,N_4537);
nor U5300 (N_5300,N_4826,N_4848);
nand U5301 (N_5301,N_4921,N_4925);
nor U5302 (N_5302,N_4865,N_4828);
nor U5303 (N_5303,N_4580,N_4847);
and U5304 (N_5304,N_4848,N_4810);
nor U5305 (N_5305,N_4802,N_4731);
and U5306 (N_5306,N_4597,N_4515);
and U5307 (N_5307,N_4626,N_4527);
and U5308 (N_5308,N_4796,N_4822);
and U5309 (N_5309,N_4670,N_4981);
or U5310 (N_5310,N_4637,N_4816);
nor U5311 (N_5311,N_4899,N_4741);
and U5312 (N_5312,N_4854,N_4965);
or U5313 (N_5313,N_4821,N_4836);
and U5314 (N_5314,N_4551,N_4735);
xor U5315 (N_5315,N_4877,N_4952);
nor U5316 (N_5316,N_4560,N_4826);
nor U5317 (N_5317,N_4683,N_4833);
nor U5318 (N_5318,N_4815,N_4615);
or U5319 (N_5319,N_4507,N_4631);
or U5320 (N_5320,N_4817,N_4936);
nand U5321 (N_5321,N_4531,N_4572);
nor U5322 (N_5322,N_4879,N_4714);
nor U5323 (N_5323,N_4916,N_4586);
nor U5324 (N_5324,N_4670,N_4675);
or U5325 (N_5325,N_4995,N_4836);
and U5326 (N_5326,N_4946,N_4819);
and U5327 (N_5327,N_4728,N_4777);
nand U5328 (N_5328,N_4634,N_4541);
nor U5329 (N_5329,N_4738,N_4955);
and U5330 (N_5330,N_4771,N_4556);
nor U5331 (N_5331,N_4509,N_4939);
and U5332 (N_5332,N_4712,N_4735);
nor U5333 (N_5333,N_4842,N_4933);
nor U5334 (N_5334,N_4907,N_4506);
nor U5335 (N_5335,N_4697,N_4642);
nand U5336 (N_5336,N_4523,N_4534);
nor U5337 (N_5337,N_4849,N_4899);
nor U5338 (N_5338,N_4762,N_4560);
nand U5339 (N_5339,N_4720,N_4792);
and U5340 (N_5340,N_4568,N_4897);
or U5341 (N_5341,N_4565,N_4618);
xor U5342 (N_5342,N_4793,N_4818);
nand U5343 (N_5343,N_4985,N_4715);
or U5344 (N_5344,N_4992,N_4828);
nor U5345 (N_5345,N_4681,N_4623);
nor U5346 (N_5346,N_4955,N_4942);
or U5347 (N_5347,N_4546,N_4660);
nor U5348 (N_5348,N_4899,N_4971);
nand U5349 (N_5349,N_4600,N_4689);
nor U5350 (N_5350,N_4757,N_4750);
nand U5351 (N_5351,N_4683,N_4525);
nand U5352 (N_5352,N_4983,N_4938);
and U5353 (N_5353,N_4598,N_4816);
nand U5354 (N_5354,N_4798,N_4995);
and U5355 (N_5355,N_4790,N_4889);
and U5356 (N_5356,N_4819,N_4936);
nor U5357 (N_5357,N_4821,N_4749);
nand U5358 (N_5358,N_4925,N_4796);
and U5359 (N_5359,N_4780,N_4970);
nor U5360 (N_5360,N_4562,N_4762);
nand U5361 (N_5361,N_4792,N_4847);
nor U5362 (N_5362,N_4508,N_4843);
nor U5363 (N_5363,N_4772,N_4882);
or U5364 (N_5364,N_4688,N_4587);
nor U5365 (N_5365,N_4788,N_4998);
nor U5366 (N_5366,N_4703,N_4894);
or U5367 (N_5367,N_4649,N_4939);
nor U5368 (N_5368,N_4845,N_4554);
nor U5369 (N_5369,N_4909,N_4705);
or U5370 (N_5370,N_4613,N_4883);
and U5371 (N_5371,N_4623,N_4760);
or U5372 (N_5372,N_4908,N_4759);
and U5373 (N_5373,N_4814,N_4600);
and U5374 (N_5374,N_4802,N_4549);
nand U5375 (N_5375,N_4751,N_4962);
or U5376 (N_5376,N_4742,N_4860);
or U5377 (N_5377,N_4758,N_4880);
and U5378 (N_5378,N_4979,N_4515);
nand U5379 (N_5379,N_4630,N_4722);
nand U5380 (N_5380,N_4707,N_4890);
or U5381 (N_5381,N_4747,N_4606);
and U5382 (N_5382,N_4506,N_4866);
nand U5383 (N_5383,N_4843,N_4705);
or U5384 (N_5384,N_4514,N_4985);
and U5385 (N_5385,N_4648,N_4806);
nand U5386 (N_5386,N_4987,N_4592);
nand U5387 (N_5387,N_4562,N_4601);
and U5388 (N_5388,N_4509,N_4797);
nand U5389 (N_5389,N_4536,N_4968);
nand U5390 (N_5390,N_4936,N_4654);
and U5391 (N_5391,N_4803,N_4971);
nor U5392 (N_5392,N_4690,N_4619);
nand U5393 (N_5393,N_4742,N_4770);
and U5394 (N_5394,N_4875,N_4845);
or U5395 (N_5395,N_4912,N_4602);
nand U5396 (N_5396,N_4782,N_4661);
or U5397 (N_5397,N_4648,N_4711);
xnor U5398 (N_5398,N_4789,N_4660);
nor U5399 (N_5399,N_4670,N_4712);
and U5400 (N_5400,N_4626,N_4943);
and U5401 (N_5401,N_4683,N_4991);
or U5402 (N_5402,N_4558,N_4821);
nor U5403 (N_5403,N_4708,N_4614);
nand U5404 (N_5404,N_4969,N_4553);
or U5405 (N_5405,N_4900,N_4627);
nand U5406 (N_5406,N_4530,N_4677);
nor U5407 (N_5407,N_4872,N_4655);
nand U5408 (N_5408,N_4941,N_4929);
or U5409 (N_5409,N_4681,N_4611);
nor U5410 (N_5410,N_4694,N_4633);
or U5411 (N_5411,N_4520,N_4857);
nand U5412 (N_5412,N_4761,N_4997);
and U5413 (N_5413,N_4962,N_4696);
nor U5414 (N_5414,N_4555,N_4831);
or U5415 (N_5415,N_4897,N_4678);
xor U5416 (N_5416,N_4652,N_4772);
nor U5417 (N_5417,N_4757,N_4588);
or U5418 (N_5418,N_4919,N_4986);
nor U5419 (N_5419,N_4722,N_4679);
or U5420 (N_5420,N_4628,N_4552);
or U5421 (N_5421,N_4990,N_4556);
and U5422 (N_5422,N_4820,N_4940);
and U5423 (N_5423,N_4735,N_4510);
and U5424 (N_5424,N_4709,N_4648);
nand U5425 (N_5425,N_4867,N_4810);
nor U5426 (N_5426,N_4874,N_4897);
nor U5427 (N_5427,N_4519,N_4750);
and U5428 (N_5428,N_4872,N_4826);
or U5429 (N_5429,N_4756,N_4811);
or U5430 (N_5430,N_4793,N_4610);
nor U5431 (N_5431,N_4510,N_4893);
or U5432 (N_5432,N_4544,N_4846);
nor U5433 (N_5433,N_4711,N_4986);
nor U5434 (N_5434,N_4858,N_4605);
xor U5435 (N_5435,N_4961,N_4890);
or U5436 (N_5436,N_4913,N_4607);
xor U5437 (N_5437,N_4721,N_4987);
or U5438 (N_5438,N_4545,N_4762);
nor U5439 (N_5439,N_4811,N_4595);
nor U5440 (N_5440,N_4660,N_4844);
or U5441 (N_5441,N_4851,N_4874);
nand U5442 (N_5442,N_4998,N_4815);
nor U5443 (N_5443,N_4687,N_4635);
and U5444 (N_5444,N_4610,N_4743);
xor U5445 (N_5445,N_4793,N_4899);
nor U5446 (N_5446,N_4798,N_4922);
nand U5447 (N_5447,N_4782,N_4532);
and U5448 (N_5448,N_4961,N_4934);
nand U5449 (N_5449,N_4884,N_4967);
and U5450 (N_5450,N_4634,N_4787);
or U5451 (N_5451,N_4534,N_4699);
and U5452 (N_5452,N_4817,N_4545);
nand U5453 (N_5453,N_4665,N_4777);
or U5454 (N_5454,N_4786,N_4934);
or U5455 (N_5455,N_4560,N_4858);
nor U5456 (N_5456,N_4744,N_4794);
or U5457 (N_5457,N_4718,N_4721);
nor U5458 (N_5458,N_4774,N_4863);
and U5459 (N_5459,N_4773,N_4906);
nor U5460 (N_5460,N_4684,N_4867);
nand U5461 (N_5461,N_4845,N_4947);
and U5462 (N_5462,N_4590,N_4615);
nand U5463 (N_5463,N_4893,N_4660);
and U5464 (N_5464,N_4603,N_4552);
and U5465 (N_5465,N_4610,N_4701);
or U5466 (N_5466,N_4597,N_4514);
or U5467 (N_5467,N_4689,N_4609);
or U5468 (N_5468,N_4649,N_4799);
and U5469 (N_5469,N_4865,N_4678);
nor U5470 (N_5470,N_4751,N_4770);
nor U5471 (N_5471,N_4931,N_4992);
nor U5472 (N_5472,N_4997,N_4804);
nand U5473 (N_5473,N_4745,N_4762);
nor U5474 (N_5474,N_4856,N_4954);
or U5475 (N_5475,N_4896,N_4516);
nand U5476 (N_5476,N_4682,N_4668);
or U5477 (N_5477,N_4951,N_4876);
and U5478 (N_5478,N_4783,N_4521);
nor U5479 (N_5479,N_4503,N_4771);
nor U5480 (N_5480,N_4874,N_4786);
nand U5481 (N_5481,N_4500,N_4772);
nand U5482 (N_5482,N_4830,N_4743);
nor U5483 (N_5483,N_4690,N_4813);
nor U5484 (N_5484,N_4873,N_4627);
or U5485 (N_5485,N_4932,N_4906);
or U5486 (N_5486,N_4619,N_4686);
and U5487 (N_5487,N_4932,N_4604);
nand U5488 (N_5488,N_4752,N_4986);
nand U5489 (N_5489,N_4590,N_4682);
or U5490 (N_5490,N_4515,N_4753);
nand U5491 (N_5491,N_4990,N_4638);
or U5492 (N_5492,N_4783,N_4854);
and U5493 (N_5493,N_4613,N_4987);
nor U5494 (N_5494,N_4731,N_4658);
nor U5495 (N_5495,N_4946,N_4613);
nor U5496 (N_5496,N_4522,N_4796);
nor U5497 (N_5497,N_4575,N_4957);
or U5498 (N_5498,N_4545,N_4848);
or U5499 (N_5499,N_4865,N_4570);
or U5500 (N_5500,N_5398,N_5051);
nor U5501 (N_5501,N_5056,N_5392);
and U5502 (N_5502,N_5302,N_5492);
and U5503 (N_5503,N_5463,N_5275);
nor U5504 (N_5504,N_5004,N_5216);
nand U5505 (N_5505,N_5022,N_5193);
or U5506 (N_5506,N_5116,N_5285);
and U5507 (N_5507,N_5094,N_5209);
nand U5508 (N_5508,N_5395,N_5461);
nor U5509 (N_5509,N_5254,N_5021);
nand U5510 (N_5510,N_5493,N_5199);
and U5511 (N_5511,N_5150,N_5298);
and U5512 (N_5512,N_5367,N_5432);
nand U5513 (N_5513,N_5165,N_5273);
nand U5514 (N_5514,N_5326,N_5419);
or U5515 (N_5515,N_5427,N_5351);
or U5516 (N_5516,N_5450,N_5341);
nand U5517 (N_5517,N_5031,N_5189);
or U5518 (N_5518,N_5194,N_5460);
nand U5519 (N_5519,N_5304,N_5289);
and U5520 (N_5520,N_5019,N_5484);
and U5521 (N_5521,N_5203,N_5205);
and U5522 (N_5522,N_5343,N_5368);
or U5523 (N_5523,N_5401,N_5356);
nand U5524 (N_5524,N_5267,N_5312);
nor U5525 (N_5525,N_5457,N_5244);
and U5526 (N_5526,N_5067,N_5123);
and U5527 (N_5527,N_5434,N_5293);
nand U5528 (N_5528,N_5237,N_5075);
and U5529 (N_5529,N_5308,N_5465);
and U5530 (N_5530,N_5352,N_5410);
nand U5531 (N_5531,N_5174,N_5062);
nand U5532 (N_5532,N_5256,N_5339);
or U5533 (N_5533,N_5278,N_5486);
and U5534 (N_5534,N_5230,N_5160);
nand U5535 (N_5535,N_5133,N_5043);
nand U5536 (N_5536,N_5489,N_5321);
nand U5537 (N_5537,N_5126,N_5477);
and U5538 (N_5538,N_5444,N_5498);
nand U5539 (N_5539,N_5111,N_5242);
and U5540 (N_5540,N_5142,N_5191);
nor U5541 (N_5541,N_5228,N_5496);
or U5542 (N_5542,N_5272,N_5329);
nor U5543 (N_5543,N_5381,N_5200);
or U5544 (N_5544,N_5172,N_5140);
or U5545 (N_5545,N_5249,N_5421);
nor U5546 (N_5546,N_5316,N_5383);
and U5547 (N_5547,N_5462,N_5428);
nand U5548 (N_5548,N_5088,N_5181);
nor U5549 (N_5549,N_5436,N_5045);
and U5550 (N_5550,N_5417,N_5217);
and U5551 (N_5551,N_5214,N_5277);
and U5552 (N_5552,N_5154,N_5349);
or U5553 (N_5553,N_5451,N_5481);
nand U5554 (N_5554,N_5141,N_5286);
or U5555 (N_5555,N_5017,N_5033);
nor U5556 (N_5556,N_5358,N_5151);
nand U5557 (N_5557,N_5466,N_5030);
nor U5558 (N_5558,N_5208,N_5029);
nand U5559 (N_5559,N_5282,N_5008);
nor U5560 (N_5560,N_5429,N_5037);
and U5561 (N_5561,N_5185,N_5259);
nand U5562 (N_5562,N_5206,N_5370);
nand U5563 (N_5563,N_5005,N_5234);
and U5564 (N_5564,N_5309,N_5317);
nor U5565 (N_5565,N_5082,N_5310);
nand U5566 (N_5566,N_5028,N_5120);
or U5567 (N_5567,N_5283,N_5485);
nand U5568 (N_5568,N_5439,N_5188);
and U5569 (N_5569,N_5219,N_5240);
or U5570 (N_5570,N_5161,N_5355);
or U5571 (N_5571,N_5110,N_5246);
nand U5572 (N_5572,N_5162,N_5041);
or U5573 (N_5573,N_5117,N_5290);
nand U5574 (N_5574,N_5297,N_5132);
or U5575 (N_5575,N_5458,N_5099);
or U5576 (N_5576,N_5404,N_5121);
nand U5577 (N_5577,N_5006,N_5125);
or U5578 (N_5578,N_5258,N_5057);
and U5579 (N_5579,N_5324,N_5414);
nor U5580 (N_5580,N_5320,N_5109);
nand U5581 (N_5581,N_5371,N_5475);
and U5582 (N_5582,N_5063,N_5332);
or U5583 (N_5583,N_5023,N_5119);
nand U5584 (N_5584,N_5291,N_5479);
or U5585 (N_5585,N_5229,N_5402);
and U5586 (N_5586,N_5337,N_5470);
nor U5587 (N_5587,N_5168,N_5134);
nand U5588 (N_5588,N_5202,N_5480);
nor U5589 (N_5589,N_5012,N_5148);
and U5590 (N_5590,N_5350,N_5182);
or U5591 (N_5591,N_5103,N_5261);
nand U5592 (N_5592,N_5157,N_5345);
and U5593 (N_5593,N_5059,N_5036);
or U5594 (N_5594,N_5014,N_5388);
and U5595 (N_5595,N_5338,N_5243);
and U5596 (N_5596,N_5076,N_5169);
or U5597 (N_5597,N_5319,N_5306);
nand U5598 (N_5598,N_5274,N_5476);
nand U5599 (N_5599,N_5074,N_5026);
and U5600 (N_5600,N_5292,N_5016);
nor U5601 (N_5601,N_5369,N_5173);
or U5602 (N_5602,N_5003,N_5129);
or U5603 (N_5603,N_5072,N_5212);
xnor U5604 (N_5604,N_5250,N_5265);
nand U5605 (N_5605,N_5374,N_5397);
nand U5606 (N_5606,N_5342,N_5105);
or U5607 (N_5607,N_5391,N_5112);
nor U5608 (N_5608,N_5394,N_5336);
nor U5609 (N_5609,N_5166,N_5459);
and U5610 (N_5610,N_5180,N_5251);
nand U5611 (N_5611,N_5420,N_5366);
and U5612 (N_5612,N_5423,N_5376);
nand U5613 (N_5613,N_5416,N_5195);
nor U5614 (N_5614,N_5415,N_5011);
nor U5615 (N_5615,N_5054,N_5340);
or U5616 (N_5616,N_5077,N_5437);
nand U5617 (N_5617,N_5070,N_5046);
nand U5618 (N_5618,N_5020,N_5107);
nor U5619 (N_5619,N_5472,N_5281);
nand U5620 (N_5620,N_5474,N_5106);
nor U5621 (N_5621,N_5178,N_5495);
or U5622 (N_5622,N_5307,N_5433);
nand U5623 (N_5623,N_5325,N_5255);
nor U5624 (N_5624,N_5002,N_5163);
and U5625 (N_5625,N_5221,N_5405);
nand U5626 (N_5626,N_5380,N_5233);
and U5627 (N_5627,N_5201,N_5048);
or U5628 (N_5628,N_5393,N_5018);
nand U5629 (N_5629,N_5090,N_5487);
nor U5630 (N_5630,N_5149,N_5176);
nor U5631 (N_5631,N_5066,N_5333);
nor U5632 (N_5632,N_5038,N_5295);
and U5633 (N_5633,N_5471,N_5353);
xor U5634 (N_5634,N_5236,N_5085);
nor U5635 (N_5635,N_5186,N_5050);
nor U5636 (N_5636,N_5053,N_5001);
and U5637 (N_5637,N_5138,N_5287);
nor U5638 (N_5638,N_5280,N_5431);
nor U5639 (N_5639,N_5210,N_5078);
and U5640 (N_5640,N_5080,N_5266);
or U5641 (N_5641,N_5296,N_5323);
and U5642 (N_5642,N_5390,N_5049);
nor U5643 (N_5643,N_5412,N_5382);
nand U5644 (N_5644,N_5055,N_5102);
nand U5645 (N_5645,N_5257,N_5362);
nand U5646 (N_5646,N_5127,N_5024);
nand U5647 (N_5647,N_5311,N_5315);
or U5648 (N_5648,N_5443,N_5378);
nor U5649 (N_5649,N_5087,N_5299);
or U5650 (N_5650,N_5318,N_5007);
nand U5651 (N_5651,N_5327,N_5071);
nand U5652 (N_5652,N_5425,N_5198);
nor U5653 (N_5653,N_5136,N_5288);
and U5654 (N_5654,N_5027,N_5042);
nand U5655 (N_5655,N_5122,N_5406);
and U5656 (N_5656,N_5190,N_5407);
nor U5657 (N_5657,N_5032,N_5093);
nor U5658 (N_5658,N_5035,N_5396);
nor U5659 (N_5659,N_5491,N_5204);
or U5660 (N_5660,N_5238,N_5235);
nand U5661 (N_5661,N_5081,N_5096);
nand U5662 (N_5662,N_5124,N_5411);
and U5663 (N_5663,N_5101,N_5455);
or U5664 (N_5664,N_5441,N_5060);
nor U5665 (N_5665,N_5473,N_5079);
and U5666 (N_5666,N_5365,N_5314);
and U5667 (N_5667,N_5490,N_5155);
nand U5668 (N_5668,N_5322,N_5488);
nor U5669 (N_5669,N_5346,N_5260);
nor U5670 (N_5670,N_5248,N_5100);
or U5671 (N_5671,N_5331,N_5167);
nor U5672 (N_5672,N_5245,N_5262);
nand U5673 (N_5673,N_5034,N_5211);
or U5674 (N_5674,N_5224,N_5399);
and U5675 (N_5675,N_5156,N_5226);
or U5676 (N_5676,N_5497,N_5084);
and U5677 (N_5677,N_5426,N_5264);
nor U5678 (N_5678,N_5453,N_5114);
and U5679 (N_5679,N_5061,N_5357);
or U5680 (N_5680,N_5301,N_5440);
nor U5681 (N_5681,N_5387,N_5268);
and U5682 (N_5682,N_5231,N_5448);
nand U5683 (N_5683,N_5247,N_5089);
or U5684 (N_5684,N_5241,N_5145);
nand U5685 (N_5685,N_5385,N_5058);
nor U5686 (N_5686,N_5108,N_5184);
nor U5687 (N_5687,N_5373,N_5025);
nor U5688 (N_5688,N_5335,N_5098);
and U5689 (N_5689,N_5386,N_5069);
nand U5690 (N_5690,N_5073,N_5364);
nor U5691 (N_5691,N_5478,N_5213);
nor U5692 (N_5692,N_5044,N_5348);
or U5693 (N_5693,N_5192,N_5179);
nand U5694 (N_5694,N_5065,N_5409);
xnor U5695 (N_5695,N_5147,N_5271);
or U5696 (N_5696,N_5276,N_5068);
nand U5697 (N_5697,N_5118,N_5253);
nand U5698 (N_5698,N_5449,N_5445);
nor U5699 (N_5699,N_5207,N_5239);
nor U5700 (N_5700,N_5400,N_5010);
nor U5701 (N_5701,N_5215,N_5359);
and U5702 (N_5702,N_5130,N_5424);
or U5703 (N_5703,N_5131,N_5334);
or U5704 (N_5704,N_5435,N_5389);
nor U5705 (N_5705,N_5135,N_5009);
nand U5706 (N_5706,N_5052,N_5363);
or U5707 (N_5707,N_5218,N_5223);
nor U5708 (N_5708,N_5153,N_5442);
nor U5709 (N_5709,N_5159,N_5361);
or U5710 (N_5710,N_5284,N_5456);
nor U5711 (N_5711,N_5305,N_5377);
nor U5712 (N_5712,N_5454,N_5438);
or U5713 (N_5713,N_5384,N_5279);
nand U5714 (N_5714,N_5499,N_5418);
nand U5715 (N_5715,N_5000,N_5013);
and U5716 (N_5716,N_5413,N_5403);
and U5717 (N_5717,N_5344,N_5128);
nor U5718 (N_5718,N_5047,N_5452);
nor U5719 (N_5719,N_5483,N_5467);
nor U5720 (N_5720,N_5294,N_5095);
nor U5721 (N_5721,N_5328,N_5197);
nand U5722 (N_5722,N_5144,N_5115);
and U5723 (N_5723,N_5177,N_5225);
nor U5724 (N_5724,N_5430,N_5252);
nor U5725 (N_5725,N_5347,N_5104);
nor U5726 (N_5726,N_5379,N_5354);
nor U5727 (N_5727,N_5039,N_5040);
and U5728 (N_5728,N_5232,N_5139);
and U5729 (N_5729,N_5482,N_5170);
nand U5730 (N_5730,N_5313,N_5227);
or U5731 (N_5731,N_5064,N_5360);
or U5732 (N_5732,N_5146,N_5171);
nor U5733 (N_5733,N_5300,N_5330);
nor U5734 (N_5734,N_5303,N_5164);
or U5735 (N_5735,N_5152,N_5187);
nor U5736 (N_5736,N_5175,N_5446);
nor U5737 (N_5737,N_5469,N_5375);
nand U5738 (N_5738,N_5183,N_5092);
or U5739 (N_5739,N_5113,N_5269);
and U5740 (N_5740,N_5137,N_5408);
nor U5741 (N_5741,N_5447,N_5372);
and U5742 (N_5742,N_5494,N_5270);
nor U5743 (N_5743,N_5097,N_5220);
nand U5744 (N_5744,N_5464,N_5263);
and U5745 (N_5745,N_5158,N_5083);
or U5746 (N_5746,N_5091,N_5015);
and U5747 (N_5747,N_5422,N_5222);
nor U5748 (N_5748,N_5143,N_5468);
and U5749 (N_5749,N_5086,N_5196);
nand U5750 (N_5750,N_5465,N_5398);
or U5751 (N_5751,N_5386,N_5373);
nor U5752 (N_5752,N_5087,N_5331);
nor U5753 (N_5753,N_5048,N_5241);
nand U5754 (N_5754,N_5151,N_5458);
nand U5755 (N_5755,N_5220,N_5430);
nor U5756 (N_5756,N_5266,N_5209);
nor U5757 (N_5757,N_5352,N_5232);
nor U5758 (N_5758,N_5344,N_5000);
nand U5759 (N_5759,N_5434,N_5229);
and U5760 (N_5760,N_5198,N_5378);
nor U5761 (N_5761,N_5443,N_5213);
nand U5762 (N_5762,N_5115,N_5259);
and U5763 (N_5763,N_5089,N_5447);
nor U5764 (N_5764,N_5411,N_5461);
nand U5765 (N_5765,N_5241,N_5267);
or U5766 (N_5766,N_5052,N_5152);
nand U5767 (N_5767,N_5312,N_5407);
or U5768 (N_5768,N_5043,N_5036);
or U5769 (N_5769,N_5483,N_5405);
and U5770 (N_5770,N_5343,N_5137);
nand U5771 (N_5771,N_5275,N_5490);
nand U5772 (N_5772,N_5414,N_5375);
nand U5773 (N_5773,N_5426,N_5249);
nor U5774 (N_5774,N_5347,N_5275);
or U5775 (N_5775,N_5438,N_5226);
and U5776 (N_5776,N_5290,N_5170);
nor U5777 (N_5777,N_5099,N_5081);
and U5778 (N_5778,N_5242,N_5359);
and U5779 (N_5779,N_5202,N_5301);
nor U5780 (N_5780,N_5037,N_5211);
or U5781 (N_5781,N_5141,N_5089);
or U5782 (N_5782,N_5250,N_5380);
nor U5783 (N_5783,N_5212,N_5215);
and U5784 (N_5784,N_5258,N_5187);
nor U5785 (N_5785,N_5097,N_5281);
nand U5786 (N_5786,N_5373,N_5299);
nor U5787 (N_5787,N_5000,N_5336);
xor U5788 (N_5788,N_5134,N_5396);
nor U5789 (N_5789,N_5435,N_5421);
nor U5790 (N_5790,N_5120,N_5458);
or U5791 (N_5791,N_5293,N_5198);
and U5792 (N_5792,N_5185,N_5393);
and U5793 (N_5793,N_5085,N_5419);
nand U5794 (N_5794,N_5209,N_5257);
or U5795 (N_5795,N_5446,N_5253);
or U5796 (N_5796,N_5059,N_5200);
and U5797 (N_5797,N_5401,N_5385);
xnor U5798 (N_5798,N_5334,N_5315);
nor U5799 (N_5799,N_5274,N_5169);
and U5800 (N_5800,N_5262,N_5209);
or U5801 (N_5801,N_5331,N_5138);
nor U5802 (N_5802,N_5264,N_5011);
or U5803 (N_5803,N_5389,N_5398);
or U5804 (N_5804,N_5355,N_5453);
nand U5805 (N_5805,N_5472,N_5256);
or U5806 (N_5806,N_5339,N_5316);
or U5807 (N_5807,N_5442,N_5309);
nor U5808 (N_5808,N_5222,N_5212);
nand U5809 (N_5809,N_5053,N_5461);
and U5810 (N_5810,N_5309,N_5464);
nor U5811 (N_5811,N_5124,N_5187);
nand U5812 (N_5812,N_5227,N_5428);
or U5813 (N_5813,N_5359,N_5205);
or U5814 (N_5814,N_5354,N_5480);
or U5815 (N_5815,N_5455,N_5476);
nor U5816 (N_5816,N_5443,N_5148);
nor U5817 (N_5817,N_5081,N_5379);
and U5818 (N_5818,N_5219,N_5178);
nand U5819 (N_5819,N_5439,N_5421);
nand U5820 (N_5820,N_5416,N_5255);
nand U5821 (N_5821,N_5293,N_5370);
or U5822 (N_5822,N_5074,N_5006);
and U5823 (N_5823,N_5260,N_5157);
or U5824 (N_5824,N_5085,N_5084);
and U5825 (N_5825,N_5046,N_5115);
nand U5826 (N_5826,N_5009,N_5052);
nor U5827 (N_5827,N_5455,N_5032);
and U5828 (N_5828,N_5063,N_5362);
or U5829 (N_5829,N_5428,N_5226);
or U5830 (N_5830,N_5044,N_5049);
or U5831 (N_5831,N_5261,N_5257);
and U5832 (N_5832,N_5382,N_5041);
or U5833 (N_5833,N_5130,N_5353);
xnor U5834 (N_5834,N_5166,N_5393);
and U5835 (N_5835,N_5220,N_5206);
and U5836 (N_5836,N_5020,N_5410);
or U5837 (N_5837,N_5450,N_5185);
nand U5838 (N_5838,N_5273,N_5096);
nand U5839 (N_5839,N_5054,N_5277);
nand U5840 (N_5840,N_5368,N_5336);
nand U5841 (N_5841,N_5034,N_5065);
nand U5842 (N_5842,N_5205,N_5234);
or U5843 (N_5843,N_5404,N_5402);
nor U5844 (N_5844,N_5421,N_5028);
nor U5845 (N_5845,N_5145,N_5480);
nor U5846 (N_5846,N_5461,N_5490);
nor U5847 (N_5847,N_5155,N_5373);
or U5848 (N_5848,N_5152,N_5062);
nor U5849 (N_5849,N_5220,N_5155);
or U5850 (N_5850,N_5077,N_5068);
and U5851 (N_5851,N_5068,N_5198);
or U5852 (N_5852,N_5407,N_5240);
nor U5853 (N_5853,N_5326,N_5135);
and U5854 (N_5854,N_5072,N_5374);
nand U5855 (N_5855,N_5340,N_5217);
nand U5856 (N_5856,N_5374,N_5179);
nor U5857 (N_5857,N_5352,N_5246);
nand U5858 (N_5858,N_5252,N_5214);
nand U5859 (N_5859,N_5360,N_5109);
or U5860 (N_5860,N_5367,N_5420);
nor U5861 (N_5861,N_5493,N_5098);
nand U5862 (N_5862,N_5446,N_5203);
nand U5863 (N_5863,N_5296,N_5483);
or U5864 (N_5864,N_5162,N_5211);
nand U5865 (N_5865,N_5141,N_5014);
and U5866 (N_5866,N_5067,N_5177);
or U5867 (N_5867,N_5433,N_5200);
and U5868 (N_5868,N_5369,N_5035);
or U5869 (N_5869,N_5001,N_5330);
or U5870 (N_5870,N_5285,N_5339);
nor U5871 (N_5871,N_5271,N_5139);
nor U5872 (N_5872,N_5150,N_5272);
nor U5873 (N_5873,N_5473,N_5443);
nor U5874 (N_5874,N_5335,N_5171);
nand U5875 (N_5875,N_5198,N_5452);
or U5876 (N_5876,N_5089,N_5130);
and U5877 (N_5877,N_5272,N_5391);
and U5878 (N_5878,N_5196,N_5122);
or U5879 (N_5879,N_5268,N_5043);
nand U5880 (N_5880,N_5052,N_5262);
nand U5881 (N_5881,N_5382,N_5149);
nor U5882 (N_5882,N_5067,N_5043);
and U5883 (N_5883,N_5325,N_5093);
nor U5884 (N_5884,N_5210,N_5470);
and U5885 (N_5885,N_5440,N_5123);
nor U5886 (N_5886,N_5192,N_5128);
or U5887 (N_5887,N_5153,N_5411);
or U5888 (N_5888,N_5138,N_5461);
nand U5889 (N_5889,N_5413,N_5019);
nand U5890 (N_5890,N_5430,N_5129);
or U5891 (N_5891,N_5111,N_5467);
nand U5892 (N_5892,N_5403,N_5334);
nor U5893 (N_5893,N_5284,N_5437);
and U5894 (N_5894,N_5027,N_5450);
or U5895 (N_5895,N_5144,N_5353);
nand U5896 (N_5896,N_5275,N_5043);
and U5897 (N_5897,N_5193,N_5305);
or U5898 (N_5898,N_5083,N_5464);
or U5899 (N_5899,N_5459,N_5333);
nand U5900 (N_5900,N_5050,N_5476);
and U5901 (N_5901,N_5201,N_5127);
and U5902 (N_5902,N_5431,N_5316);
nand U5903 (N_5903,N_5035,N_5310);
nor U5904 (N_5904,N_5483,N_5104);
nand U5905 (N_5905,N_5111,N_5070);
nor U5906 (N_5906,N_5360,N_5217);
nand U5907 (N_5907,N_5476,N_5219);
and U5908 (N_5908,N_5004,N_5405);
or U5909 (N_5909,N_5363,N_5398);
and U5910 (N_5910,N_5207,N_5080);
nor U5911 (N_5911,N_5108,N_5132);
or U5912 (N_5912,N_5499,N_5099);
nand U5913 (N_5913,N_5399,N_5336);
nand U5914 (N_5914,N_5011,N_5069);
nor U5915 (N_5915,N_5333,N_5318);
nand U5916 (N_5916,N_5037,N_5016);
and U5917 (N_5917,N_5237,N_5065);
nor U5918 (N_5918,N_5456,N_5057);
nor U5919 (N_5919,N_5058,N_5462);
or U5920 (N_5920,N_5414,N_5429);
and U5921 (N_5921,N_5302,N_5030);
or U5922 (N_5922,N_5498,N_5428);
and U5923 (N_5923,N_5068,N_5382);
nand U5924 (N_5924,N_5368,N_5344);
and U5925 (N_5925,N_5263,N_5244);
nor U5926 (N_5926,N_5404,N_5449);
or U5927 (N_5927,N_5056,N_5092);
nand U5928 (N_5928,N_5308,N_5304);
nand U5929 (N_5929,N_5321,N_5330);
or U5930 (N_5930,N_5335,N_5052);
nand U5931 (N_5931,N_5166,N_5298);
nand U5932 (N_5932,N_5243,N_5028);
nor U5933 (N_5933,N_5342,N_5135);
xnor U5934 (N_5934,N_5407,N_5218);
or U5935 (N_5935,N_5483,N_5270);
nand U5936 (N_5936,N_5024,N_5426);
xor U5937 (N_5937,N_5338,N_5493);
and U5938 (N_5938,N_5244,N_5310);
and U5939 (N_5939,N_5063,N_5480);
nand U5940 (N_5940,N_5184,N_5348);
nor U5941 (N_5941,N_5376,N_5355);
nor U5942 (N_5942,N_5332,N_5495);
nor U5943 (N_5943,N_5098,N_5337);
nor U5944 (N_5944,N_5244,N_5080);
nand U5945 (N_5945,N_5174,N_5241);
nor U5946 (N_5946,N_5062,N_5031);
nor U5947 (N_5947,N_5201,N_5481);
or U5948 (N_5948,N_5123,N_5330);
nand U5949 (N_5949,N_5148,N_5390);
or U5950 (N_5950,N_5350,N_5228);
or U5951 (N_5951,N_5373,N_5317);
and U5952 (N_5952,N_5248,N_5023);
and U5953 (N_5953,N_5177,N_5073);
and U5954 (N_5954,N_5495,N_5090);
nor U5955 (N_5955,N_5391,N_5394);
nand U5956 (N_5956,N_5439,N_5159);
or U5957 (N_5957,N_5311,N_5096);
and U5958 (N_5958,N_5320,N_5040);
nor U5959 (N_5959,N_5258,N_5460);
nor U5960 (N_5960,N_5064,N_5434);
and U5961 (N_5961,N_5280,N_5042);
nand U5962 (N_5962,N_5255,N_5297);
nand U5963 (N_5963,N_5140,N_5220);
or U5964 (N_5964,N_5457,N_5354);
nor U5965 (N_5965,N_5066,N_5026);
nor U5966 (N_5966,N_5144,N_5458);
nor U5967 (N_5967,N_5410,N_5095);
and U5968 (N_5968,N_5098,N_5246);
and U5969 (N_5969,N_5111,N_5245);
or U5970 (N_5970,N_5231,N_5358);
and U5971 (N_5971,N_5146,N_5307);
nor U5972 (N_5972,N_5490,N_5445);
xor U5973 (N_5973,N_5002,N_5339);
nor U5974 (N_5974,N_5009,N_5075);
nor U5975 (N_5975,N_5399,N_5390);
and U5976 (N_5976,N_5310,N_5407);
or U5977 (N_5977,N_5267,N_5026);
nand U5978 (N_5978,N_5494,N_5331);
nand U5979 (N_5979,N_5373,N_5495);
and U5980 (N_5980,N_5018,N_5362);
nor U5981 (N_5981,N_5147,N_5057);
and U5982 (N_5982,N_5367,N_5358);
or U5983 (N_5983,N_5226,N_5267);
nand U5984 (N_5984,N_5273,N_5258);
or U5985 (N_5985,N_5080,N_5131);
and U5986 (N_5986,N_5377,N_5037);
nor U5987 (N_5987,N_5218,N_5180);
nor U5988 (N_5988,N_5253,N_5364);
or U5989 (N_5989,N_5017,N_5217);
nand U5990 (N_5990,N_5424,N_5245);
and U5991 (N_5991,N_5005,N_5196);
nand U5992 (N_5992,N_5427,N_5110);
nor U5993 (N_5993,N_5047,N_5486);
nand U5994 (N_5994,N_5077,N_5292);
and U5995 (N_5995,N_5356,N_5063);
nand U5996 (N_5996,N_5494,N_5443);
nor U5997 (N_5997,N_5251,N_5127);
nand U5998 (N_5998,N_5271,N_5090);
nor U5999 (N_5999,N_5057,N_5024);
nand U6000 (N_6000,N_5809,N_5824);
nand U6001 (N_6001,N_5542,N_5604);
or U6002 (N_6002,N_5936,N_5525);
or U6003 (N_6003,N_5933,N_5541);
and U6004 (N_6004,N_5747,N_5917);
and U6005 (N_6005,N_5757,N_5504);
or U6006 (N_6006,N_5856,N_5527);
nand U6007 (N_6007,N_5590,N_5907);
and U6008 (N_6008,N_5644,N_5659);
nand U6009 (N_6009,N_5761,N_5599);
nor U6010 (N_6010,N_5502,N_5686);
and U6011 (N_6011,N_5973,N_5526);
and U6012 (N_6012,N_5988,N_5895);
nand U6013 (N_6013,N_5974,N_5626);
or U6014 (N_6014,N_5847,N_5744);
and U6015 (N_6015,N_5547,N_5964);
nor U6016 (N_6016,N_5536,N_5645);
nor U6017 (N_6017,N_5717,N_5913);
nand U6018 (N_6018,N_5636,N_5788);
nand U6019 (N_6019,N_5773,N_5726);
and U6020 (N_6020,N_5520,N_5640);
nand U6021 (N_6021,N_5909,N_5681);
nand U6022 (N_6022,N_5700,N_5997);
or U6023 (N_6023,N_5946,N_5537);
nor U6024 (N_6024,N_5969,N_5678);
or U6025 (N_6025,N_5822,N_5945);
nor U6026 (N_6026,N_5524,N_5957);
nor U6027 (N_6027,N_5554,N_5736);
and U6028 (N_6028,N_5820,N_5924);
and U6029 (N_6029,N_5768,N_5797);
or U6030 (N_6030,N_5707,N_5955);
nand U6031 (N_6031,N_5885,N_5980);
or U6032 (N_6032,N_5549,N_5690);
nand U6033 (N_6033,N_5656,N_5697);
nand U6034 (N_6034,N_5635,N_5649);
nand U6035 (N_6035,N_5662,N_5647);
nand U6036 (N_6036,N_5865,N_5778);
and U6037 (N_6037,N_5993,N_5598);
nand U6038 (N_6038,N_5722,N_5953);
nor U6039 (N_6039,N_5651,N_5854);
nor U6040 (N_6040,N_5733,N_5560);
nand U6041 (N_6041,N_5996,N_5511);
nor U6042 (N_6042,N_5978,N_5658);
and U6043 (N_6043,N_5588,N_5515);
and U6044 (N_6044,N_5634,N_5838);
and U6045 (N_6045,N_5593,N_5800);
nor U6046 (N_6046,N_5639,N_5523);
nand U6047 (N_6047,N_5614,N_5836);
nand U6048 (N_6048,N_5591,N_5804);
nor U6049 (N_6049,N_5742,N_5948);
nor U6050 (N_6050,N_5812,N_5643);
nand U6051 (N_6051,N_5713,N_5971);
nor U6052 (N_6052,N_5951,N_5507);
nor U6053 (N_6053,N_5687,N_5540);
nand U6054 (N_6054,N_5671,N_5840);
and U6055 (N_6055,N_5558,N_5683);
and U6056 (N_6056,N_5528,N_5921);
or U6057 (N_6057,N_5926,N_5689);
nand U6058 (N_6058,N_5825,N_5663);
and U6059 (N_6059,N_5762,N_5694);
or U6060 (N_6060,N_5503,N_5810);
and U6061 (N_6061,N_5914,N_5595);
or U6062 (N_6062,N_5811,N_5753);
and U6063 (N_6063,N_5594,N_5780);
nand U6064 (N_6064,N_5652,N_5602);
or U6065 (N_6065,N_5918,N_5606);
nand U6066 (N_6066,N_5620,N_5764);
nor U6067 (N_6067,N_5863,N_5706);
nor U6068 (N_6068,N_5986,N_5877);
and U6069 (N_6069,N_5880,N_5719);
nand U6070 (N_6070,N_5774,N_5879);
nor U6071 (N_6071,N_5585,N_5559);
and U6072 (N_6072,N_5741,N_5514);
nand U6073 (N_6073,N_5956,N_5961);
nand U6074 (N_6074,N_5912,N_5965);
nand U6075 (N_6075,N_5871,N_5579);
or U6076 (N_6076,N_5600,N_5786);
nand U6077 (N_6077,N_5740,N_5545);
and U6078 (N_6078,N_5710,N_5884);
nand U6079 (N_6079,N_5860,N_5702);
nand U6080 (N_6080,N_5882,N_5805);
or U6081 (N_6081,N_5543,N_5967);
nand U6082 (N_6082,N_5699,N_5839);
nand U6083 (N_6083,N_5894,N_5738);
or U6084 (N_6084,N_5775,N_5883);
and U6085 (N_6085,N_5653,N_5931);
or U6086 (N_6086,N_5798,N_5760);
or U6087 (N_6087,N_5958,N_5556);
nor U6088 (N_6088,N_5670,N_5848);
nor U6089 (N_6089,N_5872,N_5928);
or U6090 (N_6090,N_5565,N_5782);
and U6091 (N_6091,N_5675,N_5596);
nand U6092 (N_6092,N_5517,N_5954);
or U6093 (N_6093,N_5938,N_5712);
nor U6094 (N_6094,N_5785,N_5570);
or U6095 (N_6095,N_5576,N_5770);
or U6096 (N_6096,N_5501,N_5818);
or U6097 (N_6097,N_5716,N_5533);
nand U6098 (N_6098,N_5679,N_5637);
or U6099 (N_6099,N_5897,N_5845);
and U6100 (N_6100,N_5718,N_5915);
and U6101 (N_6101,N_5698,N_5830);
nor U6102 (N_6102,N_5841,N_5641);
nor U6103 (N_6103,N_5597,N_5688);
nor U6104 (N_6104,N_5939,N_5842);
nor U6105 (N_6105,N_5564,N_5925);
and U6106 (N_6106,N_5513,N_5942);
nand U6107 (N_6107,N_5844,N_5756);
nand U6108 (N_6108,N_5586,N_5783);
nor U6109 (N_6109,N_5630,N_5544);
or U6110 (N_6110,N_5771,N_5563);
nand U6111 (N_6111,N_5720,N_5896);
xor U6112 (N_6112,N_5566,N_5843);
nand U6113 (N_6113,N_5900,N_5869);
or U6114 (N_6114,N_5500,N_5927);
nand U6115 (N_6115,N_5669,N_5932);
nand U6116 (N_6116,N_5629,N_5616);
and U6117 (N_6117,N_5592,N_5801);
nand U6118 (N_6118,N_5734,N_5911);
nor U6119 (N_6119,N_5803,N_5920);
and U6120 (N_6120,N_5849,N_5518);
nor U6121 (N_6121,N_5555,N_5923);
nand U6122 (N_6122,N_5569,N_5512);
and U6123 (N_6123,N_5799,N_5750);
nor U6124 (N_6124,N_5919,N_5705);
or U6125 (N_6125,N_5519,N_5963);
nand U6126 (N_6126,N_5767,N_5562);
nand U6127 (N_6127,N_5832,N_5892);
or U6128 (N_6128,N_5711,N_5763);
or U6129 (N_6129,N_5866,N_5834);
or U6130 (N_6130,N_5721,N_5949);
nand U6131 (N_6131,N_5660,N_5608);
nor U6132 (N_6132,N_5508,N_5772);
or U6133 (N_6133,N_5612,N_5692);
or U6134 (N_6134,N_5682,N_5935);
or U6135 (N_6135,N_5846,N_5850);
and U6136 (N_6136,N_5724,N_5580);
nand U6137 (N_6137,N_5633,N_5950);
nand U6138 (N_6138,N_5960,N_5561);
or U6139 (N_6139,N_5858,N_5899);
nand U6140 (N_6140,N_5793,N_5759);
nor U6141 (N_6141,N_5708,N_5813);
xor U6142 (N_6142,N_5769,N_5781);
and U6143 (N_6143,N_5779,N_5859);
nand U6144 (N_6144,N_5685,N_5638);
nor U6145 (N_6145,N_5992,N_5864);
nand U6146 (N_6146,N_5615,N_5827);
or U6147 (N_6147,N_5725,N_5796);
nand U6148 (N_6148,N_5703,N_5823);
nor U6149 (N_6149,N_5867,N_5989);
and U6150 (N_6150,N_5607,N_5968);
nor U6151 (N_6151,N_5790,N_5617);
and U6152 (N_6152,N_5521,N_5904);
nand U6153 (N_6153,N_5619,N_5765);
nor U6154 (N_6154,N_5622,N_5970);
and U6155 (N_6155,N_5603,N_5819);
and U6156 (N_6156,N_5731,N_5777);
nand U6157 (N_6157,N_5618,N_5876);
nand U6158 (N_6158,N_5693,N_5966);
nand U6159 (N_6159,N_5582,N_5655);
nor U6160 (N_6160,N_5878,N_5976);
or U6161 (N_6161,N_5611,N_5623);
and U6162 (N_6162,N_5539,N_5905);
and U6163 (N_6163,N_5922,N_5530);
or U6164 (N_6164,N_5665,N_5696);
or U6165 (N_6165,N_5552,N_5704);
nor U6166 (N_6166,N_5940,N_5728);
and U6167 (N_6167,N_5743,N_5601);
or U6168 (N_6168,N_5751,N_5929);
nand U6169 (N_6169,N_5735,N_5794);
nand U6170 (N_6170,N_5862,N_5852);
and U6171 (N_6171,N_5529,N_5982);
nor U6172 (N_6172,N_5646,N_5573);
nand U6173 (N_6173,N_5755,N_5857);
nor U6174 (N_6174,N_5908,N_5701);
nor U6175 (N_6175,N_5959,N_5583);
and U6176 (N_6176,N_5505,N_5837);
nand U6177 (N_6177,N_5972,N_5510);
or U6178 (N_6178,N_5817,N_5890);
xor U6179 (N_6179,N_5998,N_5715);
nand U6180 (N_6180,N_5806,N_5546);
and U6181 (N_6181,N_5826,N_5991);
and U6182 (N_6182,N_5985,N_5535);
or U6183 (N_6183,N_5833,N_5509);
and U6184 (N_6184,N_5983,N_5621);
nand U6185 (N_6185,N_5661,N_5821);
and U6186 (N_6186,N_5934,N_5752);
and U6187 (N_6187,N_5589,N_5672);
xnor U6188 (N_6188,N_5791,N_5916);
or U6189 (N_6189,N_5714,N_5538);
and U6190 (N_6190,N_5684,N_5903);
or U6191 (N_6191,N_5572,N_5881);
or U6192 (N_6192,N_5668,N_5676);
and U6193 (N_6193,N_5990,N_5650);
or U6194 (N_6194,N_5888,N_5975);
or U6195 (N_6195,N_5674,N_5613);
and U6196 (N_6196,N_5680,N_5930);
or U6197 (N_6197,N_5808,N_5861);
nand U6198 (N_6198,N_5677,N_5667);
nor U6199 (N_6199,N_5814,N_5816);
nand U6200 (N_6200,N_5624,N_5746);
nor U6201 (N_6201,N_5789,N_5910);
nand U6202 (N_6202,N_5893,N_5732);
or U6203 (N_6203,N_5522,N_5947);
or U6204 (N_6204,N_5657,N_5835);
nor U6205 (N_6205,N_5748,N_5901);
nand U6206 (N_6206,N_5792,N_5875);
nor U6207 (N_6207,N_5962,N_5851);
nand U6208 (N_6208,N_5952,N_5737);
or U6209 (N_6209,N_5506,N_5906);
or U6210 (N_6210,N_5587,N_5627);
nand U6211 (N_6211,N_5673,N_5831);
and U6212 (N_6212,N_5979,N_5723);
and U6213 (N_6213,N_5625,N_5532);
or U6214 (N_6214,N_5666,N_5550);
nand U6215 (N_6215,N_5758,N_5886);
nand U6216 (N_6216,N_5632,N_5654);
nand U6217 (N_6217,N_5887,N_5874);
nand U6218 (N_6218,N_5575,N_5609);
or U6219 (N_6219,N_5557,N_5944);
or U6220 (N_6220,N_5941,N_5766);
or U6221 (N_6221,N_5891,N_5553);
nand U6222 (N_6222,N_5531,N_5853);
nand U6223 (N_6223,N_5995,N_5902);
or U6224 (N_6224,N_5691,N_5829);
nor U6225 (N_6225,N_5574,N_5729);
nand U6226 (N_6226,N_5610,N_5695);
or U6227 (N_6227,N_5648,N_5548);
or U6228 (N_6228,N_5749,N_5642);
nand U6229 (N_6229,N_5802,N_5994);
and U6230 (N_6230,N_5977,N_5815);
or U6231 (N_6231,N_5870,N_5631);
or U6232 (N_6232,N_5943,N_5981);
and U6233 (N_6233,N_5937,N_5568);
and U6234 (N_6234,N_5754,N_5889);
or U6235 (N_6235,N_5551,N_5628);
and U6236 (N_6236,N_5584,N_5571);
nor U6237 (N_6237,N_5855,N_5567);
and U6238 (N_6238,N_5581,N_5578);
and U6239 (N_6239,N_5787,N_5730);
nor U6240 (N_6240,N_5873,N_5828);
or U6241 (N_6241,N_5807,N_5577);
nor U6242 (N_6242,N_5664,N_5727);
nand U6243 (N_6243,N_5709,N_5987);
and U6244 (N_6244,N_5776,N_5784);
nor U6245 (N_6245,N_5739,N_5898);
nand U6246 (N_6246,N_5605,N_5516);
nor U6247 (N_6247,N_5745,N_5534);
nand U6248 (N_6248,N_5984,N_5795);
nor U6249 (N_6249,N_5999,N_5868);
nand U6250 (N_6250,N_5856,N_5854);
nor U6251 (N_6251,N_5548,N_5573);
nor U6252 (N_6252,N_5854,N_5860);
nand U6253 (N_6253,N_5812,N_5838);
nand U6254 (N_6254,N_5876,N_5857);
or U6255 (N_6255,N_5858,N_5669);
and U6256 (N_6256,N_5623,N_5653);
or U6257 (N_6257,N_5842,N_5898);
or U6258 (N_6258,N_5713,N_5845);
nand U6259 (N_6259,N_5752,N_5893);
or U6260 (N_6260,N_5559,N_5614);
nor U6261 (N_6261,N_5879,N_5790);
and U6262 (N_6262,N_5622,N_5518);
nor U6263 (N_6263,N_5636,N_5800);
nor U6264 (N_6264,N_5586,N_5883);
or U6265 (N_6265,N_5601,N_5973);
and U6266 (N_6266,N_5589,N_5853);
nand U6267 (N_6267,N_5740,N_5628);
and U6268 (N_6268,N_5738,N_5530);
and U6269 (N_6269,N_5814,N_5680);
xnor U6270 (N_6270,N_5577,N_5835);
nand U6271 (N_6271,N_5640,N_5515);
nor U6272 (N_6272,N_5520,N_5601);
or U6273 (N_6273,N_5682,N_5949);
and U6274 (N_6274,N_5841,N_5948);
and U6275 (N_6275,N_5882,N_5500);
or U6276 (N_6276,N_5565,N_5672);
nand U6277 (N_6277,N_5634,N_5921);
and U6278 (N_6278,N_5819,N_5976);
and U6279 (N_6279,N_5997,N_5629);
and U6280 (N_6280,N_5704,N_5917);
or U6281 (N_6281,N_5975,N_5675);
and U6282 (N_6282,N_5849,N_5779);
nand U6283 (N_6283,N_5905,N_5803);
nand U6284 (N_6284,N_5881,N_5604);
or U6285 (N_6285,N_5996,N_5583);
nand U6286 (N_6286,N_5542,N_5676);
nand U6287 (N_6287,N_5512,N_5613);
nand U6288 (N_6288,N_5586,N_5728);
and U6289 (N_6289,N_5748,N_5914);
and U6290 (N_6290,N_5629,N_5642);
nand U6291 (N_6291,N_5614,N_5672);
or U6292 (N_6292,N_5658,N_5896);
nand U6293 (N_6293,N_5510,N_5705);
or U6294 (N_6294,N_5584,N_5650);
nor U6295 (N_6295,N_5883,N_5776);
and U6296 (N_6296,N_5977,N_5643);
and U6297 (N_6297,N_5741,N_5537);
or U6298 (N_6298,N_5572,N_5535);
or U6299 (N_6299,N_5981,N_5920);
nand U6300 (N_6300,N_5807,N_5539);
and U6301 (N_6301,N_5704,N_5679);
nand U6302 (N_6302,N_5713,N_5744);
or U6303 (N_6303,N_5688,N_5550);
nand U6304 (N_6304,N_5546,N_5588);
or U6305 (N_6305,N_5660,N_5891);
nand U6306 (N_6306,N_5648,N_5644);
or U6307 (N_6307,N_5862,N_5872);
or U6308 (N_6308,N_5832,N_5860);
or U6309 (N_6309,N_5594,N_5740);
and U6310 (N_6310,N_5679,N_5949);
xor U6311 (N_6311,N_5580,N_5727);
nor U6312 (N_6312,N_5788,N_5912);
or U6313 (N_6313,N_5941,N_5633);
or U6314 (N_6314,N_5641,N_5726);
nand U6315 (N_6315,N_5804,N_5643);
or U6316 (N_6316,N_5624,N_5896);
or U6317 (N_6317,N_5948,N_5865);
or U6318 (N_6318,N_5846,N_5899);
nand U6319 (N_6319,N_5518,N_5565);
nor U6320 (N_6320,N_5567,N_5789);
or U6321 (N_6321,N_5518,N_5806);
or U6322 (N_6322,N_5742,N_5879);
nor U6323 (N_6323,N_5977,N_5861);
nor U6324 (N_6324,N_5572,N_5523);
and U6325 (N_6325,N_5655,N_5508);
or U6326 (N_6326,N_5904,N_5658);
or U6327 (N_6327,N_5964,N_5629);
nand U6328 (N_6328,N_5951,N_5624);
and U6329 (N_6329,N_5528,N_5925);
nor U6330 (N_6330,N_5852,N_5770);
nor U6331 (N_6331,N_5549,N_5556);
or U6332 (N_6332,N_5537,N_5812);
nand U6333 (N_6333,N_5865,N_5799);
and U6334 (N_6334,N_5683,N_5938);
nand U6335 (N_6335,N_5872,N_5787);
nor U6336 (N_6336,N_5752,N_5982);
or U6337 (N_6337,N_5602,N_5927);
or U6338 (N_6338,N_5782,N_5805);
nor U6339 (N_6339,N_5785,N_5754);
or U6340 (N_6340,N_5613,N_5976);
and U6341 (N_6341,N_5823,N_5560);
and U6342 (N_6342,N_5628,N_5899);
nor U6343 (N_6343,N_5573,N_5774);
and U6344 (N_6344,N_5713,N_5542);
and U6345 (N_6345,N_5755,N_5548);
nor U6346 (N_6346,N_5685,N_5565);
and U6347 (N_6347,N_5893,N_5773);
or U6348 (N_6348,N_5797,N_5997);
and U6349 (N_6349,N_5656,N_5995);
nor U6350 (N_6350,N_5961,N_5962);
and U6351 (N_6351,N_5718,N_5505);
or U6352 (N_6352,N_5689,N_5589);
nand U6353 (N_6353,N_5718,N_5792);
and U6354 (N_6354,N_5855,N_5986);
or U6355 (N_6355,N_5558,N_5782);
nor U6356 (N_6356,N_5593,N_5594);
nor U6357 (N_6357,N_5775,N_5924);
nand U6358 (N_6358,N_5813,N_5676);
and U6359 (N_6359,N_5897,N_5973);
nor U6360 (N_6360,N_5883,N_5984);
and U6361 (N_6361,N_5682,N_5700);
and U6362 (N_6362,N_5555,N_5527);
nand U6363 (N_6363,N_5919,N_5538);
and U6364 (N_6364,N_5550,N_5806);
nand U6365 (N_6365,N_5834,N_5779);
or U6366 (N_6366,N_5633,N_5682);
and U6367 (N_6367,N_5573,N_5819);
nor U6368 (N_6368,N_5904,N_5777);
and U6369 (N_6369,N_5960,N_5768);
and U6370 (N_6370,N_5980,N_5611);
and U6371 (N_6371,N_5967,N_5603);
nand U6372 (N_6372,N_5532,N_5890);
nand U6373 (N_6373,N_5751,N_5838);
nand U6374 (N_6374,N_5572,N_5617);
or U6375 (N_6375,N_5654,N_5518);
and U6376 (N_6376,N_5982,N_5861);
nand U6377 (N_6377,N_5503,N_5898);
and U6378 (N_6378,N_5534,N_5920);
nor U6379 (N_6379,N_5858,N_5827);
nor U6380 (N_6380,N_5547,N_5566);
or U6381 (N_6381,N_5693,N_5843);
or U6382 (N_6382,N_5662,N_5670);
nor U6383 (N_6383,N_5685,N_5960);
nor U6384 (N_6384,N_5543,N_5628);
or U6385 (N_6385,N_5889,N_5939);
nor U6386 (N_6386,N_5918,N_5774);
nor U6387 (N_6387,N_5782,N_5932);
or U6388 (N_6388,N_5977,N_5615);
or U6389 (N_6389,N_5962,N_5577);
and U6390 (N_6390,N_5535,N_5623);
and U6391 (N_6391,N_5564,N_5966);
and U6392 (N_6392,N_5712,N_5803);
nor U6393 (N_6393,N_5682,N_5692);
nor U6394 (N_6394,N_5542,N_5628);
nand U6395 (N_6395,N_5690,N_5550);
or U6396 (N_6396,N_5847,N_5944);
and U6397 (N_6397,N_5540,N_5548);
and U6398 (N_6398,N_5578,N_5558);
nand U6399 (N_6399,N_5733,N_5918);
nor U6400 (N_6400,N_5969,N_5699);
nor U6401 (N_6401,N_5572,N_5794);
nand U6402 (N_6402,N_5649,N_5549);
nand U6403 (N_6403,N_5699,N_5941);
or U6404 (N_6404,N_5516,N_5685);
nand U6405 (N_6405,N_5940,N_5979);
nand U6406 (N_6406,N_5703,N_5952);
nor U6407 (N_6407,N_5874,N_5753);
and U6408 (N_6408,N_5699,N_5923);
nor U6409 (N_6409,N_5509,N_5623);
and U6410 (N_6410,N_5784,N_5571);
or U6411 (N_6411,N_5574,N_5843);
nor U6412 (N_6412,N_5656,N_5991);
nand U6413 (N_6413,N_5949,N_5661);
nor U6414 (N_6414,N_5978,N_5607);
and U6415 (N_6415,N_5650,N_5849);
or U6416 (N_6416,N_5929,N_5675);
nand U6417 (N_6417,N_5907,N_5963);
nor U6418 (N_6418,N_5592,N_5513);
nand U6419 (N_6419,N_5685,N_5938);
and U6420 (N_6420,N_5785,N_5867);
nor U6421 (N_6421,N_5820,N_5638);
nor U6422 (N_6422,N_5510,N_5571);
or U6423 (N_6423,N_5519,N_5632);
nand U6424 (N_6424,N_5726,N_5784);
nor U6425 (N_6425,N_5734,N_5559);
nand U6426 (N_6426,N_5788,N_5871);
nand U6427 (N_6427,N_5816,N_5683);
and U6428 (N_6428,N_5774,N_5892);
and U6429 (N_6429,N_5651,N_5935);
or U6430 (N_6430,N_5843,N_5828);
and U6431 (N_6431,N_5563,N_5690);
or U6432 (N_6432,N_5862,N_5545);
and U6433 (N_6433,N_5594,N_5783);
and U6434 (N_6434,N_5537,N_5984);
nor U6435 (N_6435,N_5740,N_5516);
nor U6436 (N_6436,N_5535,N_5846);
nand U6437 (N_6437,N_5802,N_5988);
or U6438 (N_6438,N_5528,N_5936);
or U6439 (N_6439,N_5601,N_5962);
nor U6440 (N_6440,N_5628,N_5749);
nand U6441 (N_6441,N_5901,N_5841);
nand U6442 (N_6442,N_5526,N_5649);
or U6443 (N_6443,N_5574,N_5539);
nor U6444 (N_6444,N_5859,N_5858);
nand U6445 (N_6445,N_5902,N_5918);
nor U6446 (N_6446,N_5953,N_5596);
nand U6447 (N_6447,N_5644,N_5904);
or U6448 (N_6448,N_5805,N_5985);
nor U6449 (N_6449,N_5913,N_5714);
nor U6450 (N_6450,N_5641,N_5558);
nand U6451 (N_6451,N_5502,N_5813);
nand U6452 (N_6452,N_5837,N_5858);
nand U6453 (N_6453,N_5908,N_5561);
nand U6454 (N_6454,N_5892,N_5764);
and U6455 (N_6455,N_5569,N_5927);
nand U6456 (N_6456,N_5965,N_5540);
nor U6457 (N_6457,N_5965,N_5806);
or U6458 (N_6458,N_5501,N_5897);
or U6459 (N_6459,N_5629,N_5774);
nand U6460 (N_6460,N_5854,N_5869);
nor U6461 (N_6461,N_5725,N_5825);
nor U6462 (N_6462,N_5671,N_5975);
and U6463 (N_6463,N_5676,N_5681);
nand U6464 (N_6464,N_5965,N_5646);
or U6465 (N_6465,N_5591,N_5633);
and U6466 (N_6466,N_5548,N_5682);
and U6467 (N_6467,N_5955,N_5921);
nor U6468 (N_6468,N_5956,N_5664);
nor U6469 (N_6469,N_5857,N_5786);
xor U6470 (N_6470,N_5658,N_5611);
or U6471 (N_6471,N_5832,N_5590);
nand U6472 (N_6472,N_5887,N_5598);
nor U6473 (N_6473,N_5675,N_5930);
nand U6474 (N_6474,N_5622,N_5841);
or U6475 (N_6475,N_5571,N_5729);
nand U6476 (N_6476,N_5512,N_5771);
nor U6477 (N_6477,N_5912,N_5517);
and U6478 (N_6478,N_5806,N_5907);
nand U6479 (N_6479,N_5865,N_5915);
nor U6480 (N_6480,N_5910,N_5999);
nor U6481 (N_6481,N_5840,N_5934);
nand U6482 (N_6482,N_5907,N_5802);
nand U6483 (N_6483,N_5987,N_5787);
nand U6484 (N_6484,N_5793,N_5506);
and U6485 (N_6485,N_5806,N_5676);
xor U6486 (N_6486,N_5967,N_5767);
and U6487 (N_6487,N_5960,N_5556);
nor U6488 (N_6488,N_5635,N_5804);
nor U6489 (N_6489,N_5605,N_5638);
nor U6490 (N_6490,N_5984,N_5820);
nor U6491 (N_6491,N_5987,N_5842);
or U6492 (N_6492,N_5790,N_5997);
nand U6493 (N_6493,N_5792,N_5533);
and U6494 (N_6494,N_5931,N_5793);
and U6495 (N_6495,N_5975,N_5935);
nand U6496 (N_6496,N_5641,N_5655);
nand U6497 (N_6497,N_5729,N_5780);
and U6498 (N_6498,N_5507,N_5954);
or U6499 (N_6499,N_5712,N_5745);
and U6500 (N_6500,N_6099,N_6139);
nand U6501 (N_6501,N_6260,N_6225);
or U6502 (N_6502,N_6465,N_6487);
nor U6503 (N_6503,N_6146,N_6042);
or U6504 (N_6504,N_6114,N_6408);
nor U6505 (N_6505,N_6327,N_6000);
nand U6506 (N_6506,N_6073,N_6119);
or U6507 (N_6507,N_6253,N_6125);
and U6508 (N_6508,N_6353,N_6392);
nand U6509 (N_6509,N_6076,N_6012);
or U6510 (N_6510,N_6231,N_6469);
nand U6511 (N_6511,N_6266,N_6357);
nor U6512 (N_6512,N_6177,N_6223);
or U6513 (N_6513,N_6300,N_6341);
nor U6514 (N_6514,N_6192,N_6206);
and U6515 (N_6515,N_6136,N_6133);
nand U6516 (N_6516,N_6460,N_6093);
nand U6517 (N_6517,N_6482,N_6490);
nor U6518 (N_6518,N_6017,N_6080);
nor U6519 (N_6519,N_6150,N_6023);
nand U6520 (N_6520,N_6005,N_6098);
nor U6521 (N_6521,N_6387,N_6288);
and U6522 (N_6522,N_6440,N_6238);
nor U6523 (N_6523,N_6191,N_6089);
nor U6524 (N_6524,N_6097,N_6091);
or U6525 (N_6525,N_6046,N_6468);
nor U6526 (N_6526,N_6228,N_6412);
or U6527 (N_6527,N_6250,N_6145);
nand U6528 (N_6528,N_6101,N_6361);
or U6529 (N_6529,N_6245,N_6371);
nand U6530 (N_6530,N_6486,N_6416);
nand U6531 (N_6531,N_6355,N_6386);
nand U6532 (N_6532,N_6442,N_6335);
nor U6533 (N_6533,N_6441,N_6003);
nand U6534 (N_6534,N_6421,N_6033);
nor U6535 (N_6535,N_6188,N_6029);
and U6536 (N_6536,N_6088,N_6430);
and U6537 (N_6537,N_6171,N_6013);
and U6538 (N_6538,N_6247,N_6103);
or U6539 (N_6539,N_6261,N_6109);
and U6540 (N_6540,N_6481,N_6384);
and U6541 (N_6541,N_6165,N_6281);
and U6542 (N_6542,N_6218,N_6105);
nand U6543 (N_6543,N_6362,N_6167);
nand U6544 (N_6544,N_6276,N_6257);
nor U6545 (N_6545,N_6142,N_6462);
nand U6546 (N_6546,N_6354,N_6219);
or U6547 (N_6547,N_6369,N_6235);
nand U6548 (N_6548,N_6001,N_6108);
or U6549 (N_6549,N_6026,N_6246);
nand U6550 (N_6550,N_6488,N_6208);
nor U6551 (N_6551,N_6397,N_6347);
and U6552 (N_6552,N_6311,N_6022);
and U6553 (N_6553,N_6217,N_6199);
nor U6554 (N_6554,N_6379,N_6072);
nand U6555 (N_6555,N_6318,N_6415);
nand U6556 (N_6556,N_6472,N_6489);
or U6557 (N_6557,N_6485,N_6410);
and U6558 (N_6558,N_6444,N_6158);
nor U6559 (N_6559,N_6367,N_6278);
nand U6560 (N_6560,N_6140,N_6148);
xor U6561 (N_6561,N_6233,N_6376);
nand U6562 (N_6562,N_6306,N_6370);
and U6563 (N_6563,N_6198,N_6248);
nand U6564 (N_6564,N_6385,N_6273);
or U6565 (N_6565,N_6409,N_6317);
nand U6566 (N_6566,N_6036,N_6252);
and U6567 (N_6567,N_6068,N_6106);
nand U6568 (N_6568,N_6458,N_6197);
nor U6569 (N_6569,N_6423,N_6459);
nand U6570 (N_6570,N_6304,N_6346);
nand U6571 (N_6571,N_6396,N_6393);
or U6572 (N_6572,N_6259,N_6181);
xnor U6573 (N_6573,N_6478,N_6284);
nand U6574 (N_6574,N_6411,N_6417);
and U6575 (N_6575,N_6141,N_6209);
or U6576 (N_6576,N_6110,N_6004);
and U6577 (N_6577,N_6289,N_6244);
and U6578 (N_6578,N_6014,N_6302);
or U6579 (N_6579,N_6405,N_6449);
nand U6580 (N_6580,N_6085,N_6390);
nand U6581 (N_6581,N_6323,N_6314);
or U6582 (N_6582,N_6180,N_6154);
xnor U6583 (N_6583,N_6120,N_6360);
or U6584 (N_6584,N_6187,N_6185);
nand U6585 (N_6585,N_6475,N_6342);
nor U6586 (N_6586,N_6083,N_6499);
xnor U6587 (N_6587,N_6100,N_6075);
and U6588 (N_6588,N_6035,N_6236);
nor U6589 (N_6589,N_6443,N_6243);
nand U6590 (N_6590,N_6316,N_6320);
nand U6591 (N_6591,N_6404,N_6315);
nand U6592 (N_6592,N_6258,N_6414);
nor U6593 (N_6593,N_6179,N_6117);
nand U6594 (N_6594,N_6473,N_6319);
and U6595 (N_6595,N_6377,N_6184);
nand U6596 (N_6596,N_6153,N_6049);
and U6597 (N_6597,N_6204,N_6052);
nand U6598 (N_6598,N_6336,N_6143);
nor U6599 (N_6599,N_6427,N_6127);
or U6600 (N_6600,N_6104,N_6028);
or U6601 (N_6601,N_6020,N_6356);
or U6602 (N_6602,N_6493,N_6166);
or U6603 (N_6603,N_6178,N_6403);
nor U6604 (N_6604,N_6368,N_6113);
and U6605 (N_6605,N_6293,N_6064);
nand U6606 (N_6606,N_6438,N_6173);
and U6607 (N_6607,N_6265,N_6329);
nand U6608 (N_6608,N_6321,N_6275);
nor U6609 (N_6609,N_6374,N_6366);
nand U6610 (N_6610,N_6463,N_6196);
and U6611 (N_6611,N_6169,N_6305);
nand U6612 (N_6612,N_6431,N_6292);
nor U6613 (N_6613,N_6092,N_6161);
nor U6614 (N_6614,N_6494,N_6309);
nor U6615 (N_6615,N_6242,N_6340);
nand U6616 (N_6616,N_6118,N_6194);
nand U6617 (N_6617,N_6450,N_6102);
and U6618 (N_6618,N_6285,N_6131);
or U6619 (N_6619,N_6437,N_6263);
nand U6620 (N_6620,N_6388,N_6451);
nand U6621 (N_6621,N_6174,N_6121);
xor U6622 (N_6622,N_6399,N_6071);
nand U6623 (N_6623,N_6254,N_6394);
and U6624 (N_6624,N_6137,N_6447);
or U6625 (N_6625,N_6332,N_6349);
nand U6626 (N_6626,N_6380,N_6229);
nand U6627 (N_6627,N_6348,N_6215);
or U6628 (N_6628,N_6381,N_6331);
or U6629 (N_6629,N_6337,N_6291);
and U6630 (N_6630,N_6270,N_6018);
nor U6631 (N_6631,N_6081,N_6226);
and U6632 (N_6632,N_6310,N_6077);
or U6633 (N_6633,N_6160,N_6452);
nand U6634 (N_6634,N_6152,N_6457);
nand U6635 (N_6635,N_6445,N_6008);
xor U6636 (N_6636,N_6201,N_6062);
or U6637 (N_6637,N_6359,N_6419);
and U6638 (N_6638,N_6299,N_6112);
or U6639 (N_6639,N_6406,N_6221);
and U6640 (N_6640,N_6124,N_6267);
or U6641 (N_6641,N_6497,N_6144);
or U6642 (N_6642,N_6389,N_6476);
and U6643 (N_6643,N_6290,N_6294);
nand U6644 (N_6644,N_6009,N_6059);
nor U6645 (N_6645,N_6186,N_6163);
or U6646 (N_6646,N_6395,N_6477);
and U6647 (N_6647,N_6067,N_6070);
nand U6648 (N_6648,N_6128,N_6372);
and U6649 (N_6649,N_6115,N_6279);
and U6650 (N_6650,N_6183,N_6344);
nor U6651 (N_6651,N_6429,N_6205);
nand U6652 (N_6652,N_6021,N_6043);
and U6653 (N_6653,N_6065,N_6230);
nor U6654 (N_6654,N_6339,N_6413);
or U6655 (N_6655,N_6363,N_6287);
or U6656 (N_6656,N_6491,N_6138);
or U6657 (N_6657,N_6040,N_6474);
nor U6658 (N_6658,N_6031,N_6375);
nor U6659 (N_6659,N_6297,N_6239);
nor U6660 (N_6660,N_6338,N_6203);
nand U6661 (N_6661,N_6313,N_6135);
or U6662 (N_6662,N_6007,N_6400);
nor U6663 (N_6663,N_6495,N_6333);
or U6664 (N_6664,N_6050,N_6448);
or U6665 (N_6665,N_6157,N_6496);
nand U6666 (N_6666,N_6216,N_6498);
nor U6667 (N_6667,N_6434,N_6082);
or U6668 (N_6668,N_6129,N_6039);
nand U6669 (N_6669,N_6041,N_6358);
and U6670 (N_6670,N_6195,N_6132);
nand U6671 (N_6671,N_6011,N_6303);
nor U6672 (N_6672,N_6054,N_6432);
nand U6673 (N_6673,N_6364,N_6224);
and U6674 (N_6674,N_6325,N_6079);
nand U6675 (N_6675,N_6352,N_6038);
or U6676 (N_6676,N_6471,N_6383);
nand U6677 (N_6677,N_6237,N_6326);
nor U6678 (N_6678,N_6466,N_6240);
nor U6679 (N_6679,N_6467,N_6048);
and U6680 (N_6680,N_6182,N_6433);
nand U6681 (N_6681,N_6024,N_6200);
nand U6682 (N_6682,N_6277,N_6308);
nor U6683 (N_6683,N_6268,N_6061);
nor U6684 (N_6684,N_6175,N_6095);
or U6685 (N_6685,N_6087,N_6249);
nor U6686 (N_6686,N_6032,N_6030);
nor U6687 (N_6687,N_6151,N_6210);
nand U6688 (N_6688,N_6365,N_6483);
and U6689 (N_6689,N_6420,N_6213);
nor U6690 (N_6690,N_6010,N_6155);
or U6691 (N_6691,N_6424,N_6162);
or U6692 (N_6692,N_6189,N_6168);
or U6693 (N_6693,N_6207,N_6453);
and U6694 (N_6694,N_6222,N_6063);
and U6695 (N_6695,N_6090,N_6002);
and U6696 (N_6696,N_6006,N_6428);
nor U6697 (N_6697,N_6251,N_6456);
nor U6698 (N_6698,N_6147,N_6398);
nor U6699 (N_6699,N_6402,N_6149);
nand U6700 (N_6700,N_6351,N_6492);
and U6701 (N_6701,N_6283,N_6066);
or U6702 (N_6702,N_6401,N_6034);
or U6703 (N_6703,N_6373,N_6312);
xor U6704 (N_6704,N_6422,N_6202);
nand U6705 (N_6705,N_6272,N_6391);
or U6706 (N_6706,N_6055,N_6126);
nand U6707 (N_6707,N_6274,N_6096);
nor U6708 (N_6708,N_6296,N_6123);
nor U6709 (N_6709,N_6382,N_6345);
or U6710 (N_6710,N_6211,N_6045);
or U6711 (N_6711,N_6269,N_6107);
nor U6712 (N_6712,N_6464,N_6069);
nor U6713 (N_6713,N_6086,N_6407);
nand U6714 (N_6714,N_6324,N_6480);
or U6715 (N_6715,N_6328,N_6074);
or U6716 (N_6716,N_6461,N_6134);
nor U6717 (N_6717,N_6280,N_6271);
nand U6718 (N_6718,N_6295,N_6193);
and U6719 (N_6719,N_6454,N_6426);
nand U6720 (N_6720,N_6170,N_6025);
and U6721 (N_6721,N_6058,N_6255);
or U6722 (N_6722,N_6084,N_6307);
nand U6723 (N_6723,N_6418,N_6262);
or U6724 (N_6724,N_6435,N_6220);
nand U6725 (N_6725,N_6057,N_6056);
nand U6726 (N_6726,N_6130,N_6425);
and U6727 (N_6727,N_6122,N_6037);
xor U6728 (N_6728,N_6172,N_6164);
and U6729 (N_6729,N_6214,N_6016);
nand U6730 (N_6730,N_6027,N_6111);
xor U6731 (N_6731,N_6078,N_6439);
and U6732 (N_6732,N_6286,N_6479);
and U6733 (N_6733,N_6334,N_6301);
nand U6734 (N_6734,N_6156,N_6015);
nand U6735 (N_6735,N_6241,N_6232);
nand U6736 (N_6736,N_6446,N_6212);
nand U6737 (N_6737,N_6051,N_6350);
or U6738 (N_6738,N_6044,N_6264);
nor U6739 (N_6739,N_6322,N_6298);
nand U6740 (N_6740,N_6234,N_6436);
nor U6741 (N_6741,N_6227,N_6094);
nand U6742 (N_6742,N_6378,N_6116);
or U6743 (N_6743,N_6455,N_6282);
nand U6744 (N_6744,N_6019,N_6256);
nor U6745 (N_6745,N_6484,N_6047);
nor U6746 (N_6746,N_6190,N_6159);
nor U6747 (N_6747,N_6470,N_6330);
or U6748 (N_6748,N_6053,N_6343);
or U6749 (N_6749,N_6176,N_6060);
and U6750 (N_6750,N_6381,N_6036);
nor U6751 (N_6751,N_6476,N_6201);
or U6752 (N_6752,N_6093,N_6272);
and U6753 (N_6753,N_6187,N_6150);
or U6754 (N_6754,N_6462,N_6296);
nor U6755 (N_6755,N_6283,N_6010);
and U6756 (N_6756,N_6402,N_6347);
nor U6757 (N_6757,N_6434,N_6206);
or U6758 (N_6758,N_6357,N_6030);
and U6759 (N_6759,N_6262,N_6271);
or U6760 (N_6760,N_6120,N_6190);
and U6761 (N_6761,N_6195,N_6470);
nand U6762 (N_6762,N_6310,N_6127);
or U6763 (N_6763,N_6041,N_6286);
and U6764 (N_6764,N_6290,N_6236);
nor U6765 (N_6765,N_6166,N_6351);
and U6766 (N_6766,N_6278,N_6235);
or U6767 (N_6767,N_6230,N_6381);
or U6768 (N_6768,N_6320,N_6011);
nor U6769 (N_6769,N_6259,N_6044);
and U6770 (N_6770,N_6063,N_6005);
nor U6771 (N_6771,N_6358,N_6277);
nand U6772 (N_6772,N_6367,N_6229);
nand U6773 (N_6773,N_6133,N_6401);
or U6774 (N_6774,N_6190,N_6385);
and U6775 (N_6775,N_6201,N_6029);
nand U6776 (N_6776,N_6051,N_6378);
or U6777 (N_6777,N_6379,N_6175);
or U6778 (N_6778,N_6363,N_6137);
nor U6779 (N_6779,N_6337,N_6278);
and U6780 (N_6780,N_6014,N_6185);
nor U6781 (N_6781,N_6063,N_6485);
and U6782 (N_6782,N_6031,N_6367);
or U6783 (N_6783,N_6372,N_6083);
and U6784 (N_6784,N_6198,N_6100);
nor U6785 (N_6785,N_6322,N_6413);
nor U6786 (N_6786,N_6193,N_6297);
and U6787 (N_6787,N_6215,N_6396);
nand U6788 (N_6788,N_6133,N_6405);
nand U6789 (N_6789,N_6326,N_6196);
or U6790 (N_6790,N_6197,N_6329);
nand U6791 (N_6791,N_6234,N_6142);
nor U6792 (N_6792,N_6030,N_6116);
nand U6793 (N_6793,N_6364,N_6407);
or U6794 (N_6794,N_6049,N_6286);
nand U6795 (N_6795,N_6341,N_6393);
or U6796 (N_6796,N_6031,N_6004);
and U6797 (N_6797,N_6319,N_6048);
nor U6798 (N_6798,N_6383,N_6124);
or U6799 (N_6799,N_6342,N_6330);
nor U6800 (N_6800,N_6481,N_6130);
and U6801 (N_6801,N_6242,N_6454);
and U6802 (N_6802,N_6255,N_6492);
and U6803 (N_6803,N_6088,N_6483);
nor U6804 (N_6804,N_6233,N_6404);
nor U6805 (N_6805,N_6299,N_6418);
and U6806 (N_6806,N_6476,N_6320);
and U6807 (N_6807,N_6302,N_6393);
nor U6808 (N_6808,N_6175,N_6018);
or U6809 (N_6809,N_6400,N_6393);
and U6810 (N_6810,N_6065,N_6040);
nor U6811 (N_6811,N_6308,N_6360);
nor U6812 (N_6812,N_6316,N_6099);
nand U6813 (N_6813,N_6388,N_6039);
and U6814 (N_6814,N_6111,N_6493);
nand U6815 (N_6815,N_6302,N_6419);
or U6816 (N_6816,N_6331,N_6443);
and U6817 (N_6817,N_6496,N_6212);
or U6818 (N_6818,N_6388,N_6329);
nor U6819 (N_6819,N_6411,N_6230);
or U6820 (N_6820,N_6359,N_6325);
and U6821 (N_6821,N_6122,N_6351);
nor U6822 (N_6822,N_6283,N_6001);
and U6823 (N_6823,N_6273,N_6058);
and U6824 (N_6824,N_6264,N_6371);
nor U6825 (N_6825,N_6463,N_6078);
and U6826 (N_6826,N_6146,N_6316);
or U6827 (N_6827,N_6331,N_6345);
or U6828 (N_6828,N_6489,N_6326);
nor U6829 (N_6829,N_6168,N_6077);
nor U6830 (N_6830,N_6478,N_6322);
or U6831 (N_6831,N_6229,N_6144);
and U6832 (N_6832,N_6057,N_6407);
nor U6833 (N_6833,N_6306,N_6429);
nand U6834 (N_6834,N_6198,N_6292);
or U6835 (N_6835,N_6378,N_6431);
or U6836 (N_6836,N_6010,N_6368);
and U6837 (N_6837,N_6421,N_6308);
or U6838 (N_6838,N_6035,N_6245);
nand U6839 (N_6839,N_6235,N_6163);
and U6840 (N_6840,N_6436,N_6459);
nand U6841 (N_6841,N_6167,N_6087);
or U6842 (N_6842,N_6374,N_6419);
nor U6843 (N_6843,N_6087,N_6473);
nor U6844 (N_6844,N_6297,N_6171);
nand U6845 (N_6845,N_6183,N_6024);
nand U6846 (N_6846,N_6242,N_6329);
and U6847 (N_6847,N_6013,N_6059);
or U6848 (N_6848,N_6383,N_6499);
nand U6849 (N_6849,N_6475,N_6405);
nor U6850 (N_6850,N_6179,N_6291);
nand U6851 (N_6851,N_6442,N_6176);
nor U6852 (N_6852,N_6386,N_6004);
and U6853 (N_6853,N_6399,N_6197);
or U6854 (N_6854,N_6437,N_6431);
or U6855 (N_6855,N_6476,N_6491);
nor U6856 (N_6856,N_6116,N_6044);
nor U6857 (N_6857,N_6326,N_6211);
nand U6858 (N_6858,N_6388,N_6033);
nor U6859 (N_6859,N_6430,N_6332);
and U6860 (N_6860,N_6345,N_6259);
and U6861 (N_6861,N_6485,N_6084);
nor U6862 (N_6862,N_6219,N_6083);
or U6863 (N_6863,N_6324,N_6333);
nand U6864 (N_6864,N_6126,N_6471);
and U6865 (N_6865,N_6084,N_6409);
and U6866 (N_6866,N_6374,N_6068);
nand U6867 (N_6867,N_6218,N_6230);
and U6868 (N_6868,N_6314,N_6192);
or U6869 (N_6869,N_6338,N_6297);
nand U6870 (N_6870,N_6078,N_6288);
and U6871 (N_6871,N_6162,N_6310);
nand U6872 (N_6872,N_6268,N_6489);
and U6873 (N_6873,N_6074,N_6047);
nand U6874 (N_6874,N_6381,N_6072);
nor U6875 (N_6875,N_6495,N_6207);
and U6876 (N_6876,N_6443,N_6150);
nor U6877 (N_6877,N_6250,N_6198);
nand U6878 (N_6878,N_6333,N_6309);
and U6879 (N_6879,N_6388,N_6275);
or U6880 (N_6880,N_6464,N_6425);
nand U6881 (N_6881,N_6441,N_6119);
or U6882 (N_6882,N_6027,N_6313);
nand U6883 (N_6883,N_6492,N_6242);
and U6884 (N_6884,N_6300,N_6234);
and U6885 (N_6885,N_6275,N_6302);
and U6886 (N_6886,N_6000,N_6095);
nand U6887 (N_6887,N_6248,N_6375);
nand U6888 (N_6888,N_6110,N_6481);
or U6889 (N_6889,N_6181,N_6273);
nor U6890 (N_6890,N_6291,N_6313);
and U6891 (N_6891,N_6075,N_6448);
or U6892 (N_6892,N_6182,N_6357);
nor U6893 (N_6893,N_6213,N_6315);
and U6894 (N_6894,N_6105,N_6061);
nand U6895 (N_6895,N_6063,N_6462);
or U6896 (N_6896,N_6433,N_6066);
or U6897 (N_6897,N_6389,N_6414);
nor U6898 (N_6898,N_6064,N_6133);
and U6899 (N_6899,N_6292,N_6345);
nand U6900 (N_6900,N_6274,N_6225);
nor U6901 (N_6901,N_6424,N_6198);
nand U6902 (N_6902,N_6125,N_6240);
and U6903 (N_6903,N_6309,N_6344);
nor U6904 (N_6904,N_6063,N_6014);
nand U6905 (N_6905,N_6322,N_6157);
or U6906 (N_6906,N_6484,N_6086);
nand U6907 (N_6907,N_6073,N_6420);
nand U6908 (N_6908,N_6324,N_6205);
or U6909 (N_6909,N_6361,N_6087);
nand U6910 (N_6910,N_6137,N_6499);
nor U6911 (N_6911,N_6476,N_6368);
nor U6912 (N_6912,N_6002,N_6253);
and U6913 (N_6913,N_6136,N_6217);
or U6914 (N_6914,N_6310,N_6407);
nand U6915 (N_6915,N_6392,N_6134);
nor U6916 (N_6916,N_6324,N_6031);
and U6917 (N_6917,N_6358,N_6071);
nor U6918 (N_6918,N_6288,N_6249);
and U6919 (N_6919,N_6273,N_6271);
or U6920 (N_6920,N_6313,N_6331);
nand U6921 (N_6921,N_6173,N_6477);
nor U6922 (N_6922,N_6298,N_6066);
and U6923 (N_6923,N_6451,N_6019);
nor U6924 (N_6924,N_6453,N_6205);
and U6925 (N_6925,N_6321,N_6092);
nor U6926 (N_6926,N_6225,N_6262);
or U6927 (N_6927,N_6486,N_6188);
nand U6928 (N_6928,N_6242,N_6138);
nor U6929 (N_6929,N_6286,N_6388);
nor U6930 (N_6930,N_6272,N_6417);
and U6931 (N_6931,N_6436,N_6012);
nand U6932 (N_6932,N_6383,N_6276);
nor U6933 (N_6933,N_6108,N_6022);
and U6934 (N_6934,N_6263,N_6118);
nand U6935 (N_6935,N_6053,N_6121);
and U6936 (N_6936,N_6331,N_6071);
and U6937 (N_6937,N_6345,N_6142);
and U6938 (N_6938,N_6156,N_6122);
nand U6939 (N_6939,N_6016,N_6390);
nor U6940 (N_6940,N_6327,N_6179);
nor U6941 (N_6941,N_6270,N_6283);
and U6942 (N_6942,N_6355,N_6062);
or U6943 (N_6943,N_6420,N_6191);
nand U6944 (N_6944,N_6499,N_6133);
or U6945 (N_6945,N_6132,N_6090);
nor U6946 (N_6946,N_6375,N_6012);
nor U6947 (N_6947,N_6337,N_6117);
nor U6948 (N_6948,N_6400,N_6135);
nor U6949 (N_6949,N_6259,N_6021);
or U6950 (N_6950,N_6405,N_6289);
nand U6951 (N_6951,N_6470,N_6084);
and U6952 (N_6952,N_6490,N_6379);
or U6953 (N_6953,N_6250,N_6106);
nor U6954 (N_6954,N_6229,N_6035);
and U6955 (N_6955,N_6025,N_6332);
or U6956 (N_6956,N_6393,N_6023);
xor U6957 (N_6957,N_6465,N_6228);
nand U6958 (N_6958,N_6158,N_6182);
nand U6959 (N_6959,N_6479,N_6145);
nor U6960 (N_6960,N_6441,N_6183);
or U6961 (N_6961,N_6057,N_6278);
or U6962 (N_6962,N_6457,N_6048);
nand U6963 (N_6963,N_6198,N_6383);
or U6964 (N_6964,N_6483,N_6399);
nor U6965 (N_6965,N_6172,N_6328);
or U6966 (N_6966,N_6002,N_6445);
or U6967 (N_6967,N_6354,N_6216);
and U6968 (N_6968,N_6424,N_6059);
nand U6969 (N_6969,N_6046,N_6179);
or U6970 (N_6970,N_6320,N_6068);
nor U6971 (N_6971,N_6239,N_6123);
and U6972 (N_6972,N_6110,N_6212);
and U6973 (N_6973,N_6061,N_6461);
and U6974 (N_6974,N_6175,N_6019);
or U6975 (N_6975,N_6109,N_6315);
or U6976 (N_6976,N_6293,N_6352);
nand U6977 (N_6977,N_6161,N_6355);
or U6978 (N_6978,N_6043,N_6475);
nand U6979 (N_6979,N_6158,N_6051);
and U6980 (N_6980,N_6267,N_6415);
nand U6981 (N_6981,N_6471,N_6371);
or U6982 (N_6982,N_6181,N_6117);
xor U6983 (N_6983,N_6289,N_6457);
nand U6984 (N_6984,N_6077,N_6126);
nand U6985 (N_6985,N_6004,N_6248);
nand U6986 (N_6986,N_6220,N_6398);
and U6987 (N_6987,N_6102,N_6051);
or U6988 (N_6988,N_6225,N_6144);
nand U6989 (N_6989,N_6025,N_6200);
nand U6990 (N_6990,N_6478,N_6389);
nor U6991 (N_6991,N_6308,N_6399);
nand U6992 (N_6992,N_6333,N_6314);
nand U6993 (N_6993,N_6324,N_6491);
and U6994 (N_6994,N_6000,N_6198);
nor U6995 (N_6995,N_6079,N_6078);
nand U6996 (N_6996,N_6431,N_6186);
nand U6997 (N_6997,N_6419,N_6088);
or U6998 (N_6998,N_6166,N_6466);
or U6999 (N_6999,N_6232,N_6463);
or U7000 (N_7000,N_6842,N_6965);
or U7001 (N_7001,N_6608,N_6695);
nor U7002 (N_7002,N_6687,N_6854);
and U7003 (N_7003,N_6989,N_6894);
or U7004 (N_7004,N_6865,N_6612);
or U7005 (N_7005,N_6868,N_6838);
or U7006 (N_7006,N_6554,N_6658);
nor U7007 (N_7007,N_6729,N_6970);
and U7008 (N_7008,N_6947,N_6665);
nand U7009 (N_7009,N_6964,N_6768);
nand U7010 (N_7010,N_6872,N_6821);
nor U7011 (N_7011,N_6938,N_6848);
nor U7012 (N_7012,N_6591,N_6693);
nor U7013 (N_7013,N_6756,N_6589);
and U7014 (N_7014,N_6962,N_6992);
or U7015 (N_7015,N_6610,N_6611);
nor U7016 (N_7016,N_6902,N_6883);
and U7017 (N_7017,N_6727,N_6792);
nor U7018 (N_7018,N_6579,N_6606);
and U7019 (N_7019,N_6900,N_6532);
and U7020 (N_7020,N_6956,N_6661);
or U7021 (N_7021,N_6567,N_6908);
nor U7022 (N_7022,N_6997,N_6577);
or U7023 (N_7023,N_6820,N_6582);
nor U7024 (N_7024,N_6599,N_6887);
or U7025 (N_7025,N_6690,N_6776);
and U7026 (N_7026,N_6588,N_6939);
or U7027 (N_7027,N_6761,N_6773);
and U7028 (N_7028,N_6736,N_6853);
nand U7029 (N_7029,N_6787,N_6858);
nand U7030 (N_7030,N_6814,N_6988);
or U7031 (N_7031,N_6668,N_6779);
xnor U7032 (N_7032,N_6638,N_6518);
nor U7033 (N_7033,N_6824,N_6837);
nand U7034 (N_7034,N_6869,N_6609);
or U7035 (N_7035,N_6874,N_6969);
nand U7036 (N_7036,N_6831,N_6981);
or U7037 (N_7037,N_6598,N_6728);
and U7038 (N_7038,N_6948,N_6982);
nor U7039 (N_7039,N_6734,N_6985);
or U7040 (N_7040,N_6507,N_6559);
or U7041 (N_7041,N_6927,N_6644);
xnor U7042 (N_7042,N_6651,N_6841);
or U7043 (N_7043,N_6688,N_6917);
or U7044 (N_7044,N_6685,N_6891);
nand U7045 (N_7045,N_6654,N_6556);
nand U7046 (N_7046,N_6692,N_6862);
nand U7047 (N_7047,N_6595,N_6944);
and U7048 (N_7048,N_6694,N_6603);
nor U7049 (N_7049,N_6528,N_6839);
nor U7050 (N_7050,N_6583,N_6635);
nor U7051 (N_7051,N_6879,N_6666);
or U7052 (N_7052,N_6797,N_6571);
nor U7053 (N_7053,N_6664,N_6790);
nor U7054 (N_7054,N_6924,N_6500);
or U7055 (N_7055,N_6758,N_6830);
nand U7056 (N_7056,N_6735,N_6524);
and U7057 (N_7057,N_6557,N_6513);
nor U7058 (N_7058,N_6523,N_6561);
nand U7059 (N_7059,N_6960,N_6684);
nor U7060 (N_7060,N_6984,N_6630);
nand U7061 (N_7061,N_6922,N_6877);
nor U7062 (N_7062,N_6604,N_6569);
nand U7063 (N_7063,N_6551,N_6618);
or U7064 (N_7064,N_6657,N_6520);
and U7065 (N_7065,N_6995,N_6601);
and U7066 (N_7066,N_6913,N_6763);
or U7067 (N_7067,N_6809,N_6623);
and U7068 (N_7068,N_6961,N_6748);
and U7069 (N_7069,N_6752,N_6896);
nor U7070 (N_7070,N_6680,N_6574);
and U7071 (N_7071,N_6732,N_6682);
nor U7072 (N_7072,N_6505,N_6808);
or U7073 (N_7073,N_6542,N_6713);
and U7074 (N_7074,N_6619,N_6867);
nand U7075 (N_7075,N_6875,N_6674);
nor U7076 (N_7076,N_6593,N_6765);
nand U7077 (N_7077,N_6503,N_6940);
or U7078 (N_7078,N_6564,N_6570);
nor U7079 (N_7079,N_6585,N_6640);
nor U7080 (N_7080,N_6725,N_6681);
nand U7081 (N_7081,N_6886,N_6718);
nor U7082 (N_7082,N_6671,N_6760);
and U7083 (N_7083,N_6866,N_6861);
and U7084 (N_7084,N_6791,N_6555);
or U7085 (N_7085,N_6535,N_6749);
nor U7086 (N_7086,N_6815,N_6798);
nand U7087 (N_7087,N_6504,N_6967);
or U7088 (N_7088,N_6534,N_6803);
nor U7089 (N_7089,N_6807,N_6942);
nand U7090 (N_7090,N_6538,N_6907);
and U7091 (N_7091,N_6953,N_6702);
or U7092 (N_7092,N_6525,N_6719);
or U7093 (N_7093,N_6622,N_6785);
nor U7094 (N_7094,N_6515,N_6512);
nand U7095 (N_7095,N_6627,N_6678);
nand U7096 (N_7096,N_6899,N_6882);
nand U7097 (N_7097,N_6739,N_6508);
or U7098 (N_7098,N_6950,N_6552);
or U7099 (N_7099,N_6783,N_6592);
nand U7100 (N_7100,N_6918,N_6714);
nand U7101 (N_7101,N_6716,N_6636);
and U7102 (N_7102,N_6597,N_6539);
nand U7103 (N_7103,N_6537,N_6823);
and U7104 (N_7104,N_6708,N_6700);
nand U7105 (N_7105,N_6626,N_6957);
nand U7106 (N_7106,N_6793,N_6977);
or U7107 (N_7107,N_6613,N_6740);
nor U7108 (N_7108,N_6717,N_6715);
and U7109 (N_7109,N_6655,N_6946);
xnor U7110 (N_7110,N_6549,N_6851);
nand U7111 (N_7111,N_6802,N_6796);
and U7112 (N_7112,N_6706,N_6852);
nor U7113 (N_7113,N_6544,N_6782);
or U7114 (N_7114,N_6971,N_6526);
nor U7115 (N_7115,N_6911,N_6634);
nor U7116 (N_7116,N_6605,N_6677);
nor U7117 (N_7117,N_6986,N_6683);
nor U7118 (N_7118,N_6701,N_6774);
nand U7119 (N_7119,N_6553,N_6843);
nor U7120 (N_7120,N_6993,N_6958);
nand U7121 (N_7121,N_6712,N_6963);
nor U7122 (N_7122,N_6932,N_6943);
nand U7123 (N_7123,N_6772,N_6705);
nand U7124 (N_7124,N_6836,N_6696);
nor U7125 (N_7125,N_6864,N_6855);
or U7126 (N_7126,N_6607,N_6898);
and U7127 (N_7127,N_6781,N_6813);
or U7128 (N_7128,N_6745,N_6722);
nand U7129 (N_7129,N_6777,N_6594);
nand U7130 (N_7130,N_6691,N_6656);
and U7131 (N_7131,N_6757,N_6901);
nand U7132 (N_7132,N_6983,N_6633);
nor U7133 (N_7133,N_6949,N_6751);
nor U7134 (N_7134,N_6876,N_6895);
and U7135 (N_7135,N_6990,N_6642);
or U7136 (N_7136,N_6572,N_6662);
or U7137 (N_7137,N_6543,N_6966);
nand U7138 (N_7138,N_6580,N_6889);
and U7139 (N_7139,N_6936,N_6522);
nor U7140 (N_7140,N_6778,N_6743);
xnor U7141 (N_7141,N_6923,N_6780);
nor U7142 (N_7142,N_6560,N_6650);
nand U7143 (N_7143,N_6675,N_6649);
or U7144 (N_7144,N_6999,N_6912);
nor U7145 (N_7145,N_6873,N_6514);
and U7146 (N_7146,N_6738,N_6941);
or U7147 (N_7147,N_6646,N_6670);
or U7148 (N_7148,N_6850,N_6741);
and U7149 (N_7149,N_6653,N_6976);
and U7150 (N_7150,N_6721,N_6914);
and U7151 (N_7151,N_6925,N_6531);
nor U7152 (N_7152,N_6737,N_6615);
and U7153 (N_7153,N_6632,N_6698);
or U7154 (N_7154,N_6786,N_6659);
nand U7155 (N_7155,N_6959,N_6910);
nor U7156 (N_7156,N_6770,N_6517);
or U7157 (N_7157,N_6581,N_6952);
nand U7158 (N_7158,N_6699,N_6998);
or U7159 (N_7159,N_6935,N_6587);
or U7160 (N_7160,N_6974,N_6929);
and U7161 (N_7161,N_6529,N_6903);
and U7162 (N_7162,N_6906,N_6972);
or U7163 (N_7163,N_6816,N_6643);
or U7164 (N_7164,N_6915,N_6616);
or U7165 (N_7165,N_6931,N_6568);
nand U7166 (N_7166,N_6759,N_6527);
and U7167 (N_7167,N_6926,N_6870);
nor U7168 (N_7168,N_6892,N_6928);
and U7169 (N_7169,N_6955,N_6888);
nand U7170 (N_7170,N_6600,N_6794);
nor U7171 (N_7171,N_6881,N_6686);
or U7172 (N_7172,N_6663,N_6614);
nand U7173 (N_7173,N_6510,N_6835);
nand U7174 (N_7174,N_6822,N_6769);
nor U7175 (N_7175,N_6673,N_6720);
nand U7176 (N_7176,N_6826,N_6921);
and U7177 (N_7177,N_6885,N_6847);
and U7178 (N_7178,N_6904,N_6652);
and U7179 (N_7179,N_6845,N_6711);
and U7180 (N_7180,N_6704,N_6707);
nor U7181 (N_7181,N_6819,N_6540);
or U7182 (N_7182,N_6934,N_6825);
nor U7183 (N_7183,N_6754,N_6536);
xnor U7184 (N_7184,N_6755,N_6775);
nand U7185 (N_7185,N_6811,N_6506);
and U7186 (N_7186,N_6679,N_6550);
nor U7187 (N_7187,N_6629,N_6624);
and U7188 (N_7188,N_6799,N_6753);
and U7189 (N_7189,N_6501,N_6689);
and U7190 (N_7190,N_6788,N_6833);
nand U7191 (N_7191,N_6849,N_6558);
nand U7192 (N_7192,N_6509,N_6631);
nand U7193 (N_7193,N_6897,N_6733);
nor U7194 (N_7194,N_6817,N_6994);
nor U7195 (N_7195,N_6909,N_6951);
or U7196 (N_7196,N_6731,N_6810);
xor U7197 (N_7197,N_6546,N_6795);
nor U7198 (N_7198,N_6893,N_6647);
and U7199 (N_7199,N_6625,N_6703);
or U7200 (N_7200,N_6933,N_6829);
nand U7201 (N_7201,N_6562,N_6547);
nand U7202 (N_7202,N_6828,N_6863);
or U7203 (N_7203,N_6639,N_6937);
or U7204 (N_7204,N_6519,N_6533);
and U7205 (N_7205,N_6857,N_6846);
and U7206 (N_7206,N_6516,N_6784);
and U7207 (N_7207,N_6596,N_6919);
nor U7208 (N_7208,N_6945,N_6805);
nand U7209 (N_7209,N_6860,N_6521);
nand U7210 (N_7210,N_6672,N_6832);
and U7211 (N_7211,N_6996,N_6767);
or U7212 (N_7212,N_6812,N_6575);
and U7213 (N_7213,N_6742,N_6676);
or U7214 (N_7214,N_6954,N_6730);
or U7215 (N_7215,N_6884,N_6744);
xor U7216 (N_7216,N_6800,N_6916);
nand U7217 (N_7217,N_6804,N_6801);
nand U7218 (N_7218,N_6871,N_6697);
and U7219 (N_7219,N_6645,N_6709);
nor U7220 (N_7220,N_6750,N_6973);
nor U7221 (N_7221,N_6621,N_6590);
nor U7222 (N_7222,N_6578,N_6764);
or U7223 (N_7223,N_6840,N_6566);
nand U7224 (N_7224,N_6920,N_6620);
or U7225 (N_7225,N_6980,N_6541);
and U7226 (N_7226,N_6545,N_6905);
or U7227 (N_7227,N_6576,N_6834);
nor U7228 (N_7228,N_6979,N_6806);
and U7229 (N_7229,N_6648,N_6747);
and U7230 (N_7230,N_6511,N_6844);
nand U7231 (N_7231,N_6530,N_6584);
or U7232 (N_7232,N_6978,N_6766);
nand U7233 (N_7233,N_6502,N_6991);
and U7234 (N_7234,N_6930,N_6573);
and U7235 (N_7235,N_6968,N_6762);
nand U7236 (N_7236,N_6818,N_6880);
xor U7237 (N_7237,N_6602,N_6771);
nand U7238 (N_7238,N_6726,N_6637);
and U7239 (N_7239,N_6565,N_6859);
nand U7240 (N_7240,N_6827,N_6878);
or U7241 (N_7241,N_6667,N_6975);
or U7242 (N_7242,N_6617,N_6641);
nor U7243 (N_7243,N_6660,N_6890);
and U7244 (N_7244,N_6548,N_6563);
and U7245 (N_7245,N_6628,N_6586);
and U7246 (N_7246,N_6746,N_6723);
nand U7247 (N_7247,N_6856,N_6987);
nand U7248 (N_7248,N_6724,N_6669);
nor U7249 (N_7249,N_6710,N_6789);
nand U7250 (N_7250,N_6655,N_6754);
and U7251 (N_7251,N_6643,N_6516);
and U7252 (N_7252,N_6501,N_6989);
and U7253 (N_7253,N_6561,N_6612);
and U7254 (N_7254,N_6633,N_6544);
and U7255 (N_7255,N_6811,N_6862);
nor U7256 (N_7256,N_6793,N_6856);
xnor U7257 (N_7257,N_6585,N_6696);
or U7258 (N_7258,N_6687,N_6592);
or U7259 (N_7259,N_6649,N_6535);
and U7260 (N_7260,N_6939,N_6712);
nand U7261 (N_7261,N_6961,N_6702);
or U7262 (N_7262,N_6517,N_6596);
nor U7263 (N_7263,N_6606,N_6591);
or U7264 (N_7264,N_6617,N_6902);
nor U7265 (N_7265,N_6832,N_6562);
nand U7266 (N_7266,N_6642,N_6659);
and U7267 (N_7267,N_6980,N_6632);
nand U7268 (N_7268,N_6763,N_6745);
and U7269 (N_7269,N_6584,N_6794);
and U7270 (N_7270,N_6513,N_6632);
nor U7271 (N_7271,N_6877,N_6915);
and U7272 (N_7272,N_6714,N_6624);
nand U7273 (N_7273,N_6712,N_6915);
nor U7274 (N_7274,N_6760,N_6846);
nand U7275 (N_7275,N_6987,N_6898);
and U7276 (N_7276,N_6785,N_6516);
and U7277 (N_7277,N_6686,N_6599);
and U7278 (N_7278,N_6536,N_6953);
nand U7279 (N_7279,N_6894,N_6625);
and U7280 (N_7280,N_6837,N_6798);
or U7281 (N_7281,N_6802,N_6974);
and U7282 (N_7282,N_6595,N_6699);
or U7283 (N_7283,N_6561,N_6563);
nand U7284 (N_7284,N_6988,N_6550);
and U7285 (N_7285,N_6979,N_6577);
nand U7286 (N_7286,N_6620,N_6551);
or U7287 (N_7287,N_6855,N_6592);
nand U7288 (N_7288,N_6622,N_6689);
and U7289 (N_7289,N_6786,N_6855);
nor U7290 (N_7290,N_6808,N_6860);
nor U7291 (N_7291,N_6981,N_6813);
nor U7292 (N_7292,N_6576,N_6671);
nand U7293 (N_7293,N_6569,N_6531);
and U7294 (N_7294,N_6974,N_6852);
or U7295 (N_7295,N_6516,N_6548);
and U7296 (N_7296,N_6741,N_6544);
or U7297 (N_7297,N_6689,N_6943);
nand U7298 (N_7298,N_6500,N_6522);
or U7299 (N_7299,N_6679,N_6646);
nor U7300 (N_7300,N_6835,N_6750);
nand U7301 (N_7301,N_6927,N_6898);
nand U7302 (N_7302,N_6699,N_6506);
nor U7303 (N_7303,N_6922,N_6837);
nor U7304 (N_7304,N_6948,N_6514);
nand U7305 (N_7305,N_6943,N_6754);
or U7306 (N_7306,N_6759,N_6890);
xor U7307 (N_7307,N_6612,N_6542);
or U7308 (N_7308,N_6923,N_6939);
nand U7309 (N_7309,N_6933,N_6769);
and U7310 (N_7310,N_6865,N_6781);
and U7311 (N_7311,N_6581,N_6919);
and U7312 (N_7312,N_6928,N_6919);
or U7313 (N_7313,N_6877,N_6949);
and U7314 (N_7314,N_6977,N_6759);
or U7315 (N_7315,N_6912,N_6750);
nand U7316 (N_7316,N_6558,N_6640);
or U7317 (N_7317,N_6881,N_6590);
nor U7318 (N_7318,N_6522,N_6756);
or U7319 (N_7319,N_6656,N_6846);
nor U7320 (N_7320,N_6797,N_6821);
and U7321 (N_7321,N_6999,N_6752);
and U7322 (N_7322,N_6676,N_6577);
and U7323 (N_7323,N_6507,N_6814);
or U7324 (N_7324,N_6805,N_6722);
nor U7325 (N_7325,N_6648,N_6943);
xor U7326 (N_7326,N_6783,N_6589);
nand U7327 (N_7327,N_6867,N_6687);
nor U7328 (N_7328,N_6933,N_6994);
and U7329 (N_7329,N_6949,N_6995);
nor U7330 (N_7330,N_6569,N_6688);
or U7331 (N_7331,N_6925,N_6611);
and U7332 (N_7332,N_6676,N_6699);
nand U7333 (N_7333,N_6563,N_6532);
or U7334 (N_7334,N_6790,N_6630);
nand U7335 (N_7335,N_6944,N_6808);
nor U7336 (N_7336,N_6883,N_6579);
or U7337 (N_7337,N_6728,N_6963);
or U7338 (N_7338,N_6794,N_6707);
and U7339 (N_7339,N_6610,N_6738);
and U7340 (N_7340,N_6912,N_6786);
nand U7341 (N_7341,N_6512,N_6692);
nand U7342 (N_7342,N_6644,N_6950);
and U7343 (N_7343,N_6758,N_6981);
or U7344 (N_7344,N_6667,N_6785);
or U7345 (N_7345,N_6545,N_6576);
nand U7346 (N_7346,N_6644,N_6634);
and U7347 (N_7347,N_6616,N_6908);
xnor U7348 (N_7348,N_6733,N_6978);
or U7349 (N_7349,N_6746,N_6900);
nand U7350 (N_7350,N_6517,N_6888);
and U7351 (N_7351,N_6786,N_6731);
and U7352 (N_7352,N_6694,N_6854);
or U7353 (N_7353,N_6721,N_6576);
or U7354 (N_7354,N_6665,N_6847);
nor U7355 (N_7355,N_6752,N_6516);
nor U7356 (N_7356,N_6670,N_6845);
nor U7357 (N_7357,N_6915,N_6983);
nor U7358 (N_7358,N_6504,N_6763);
or U7359 (N_7359,N_6752,N_6840);
or U7360 (N_7360,N_6918,N_6988);
nand U7361 (N_7361,N_6521,N_6916);
and U7362 (N_7362,N_6594,N_6762);
or U7363 (N_7363,N_6543,N_6651);
and U7364 (N_7364,N_6712,N_6826);
nand U7365 (N_7365,N_6622,N_6987);
and U7366 (N_7366,N_6577,N_6683);
nor U7367 (N_7367,N_6742,N_6725);
xnor U7368 (N_7368,N_6932,N_6556);
and U7369 (N_7369,N_6511,N_6990);
or U7370 (N_7370,N_6974,N_6512);
and U7371 (N_7371,N_6661,N_6997);
nand U7372 (N_7372,N_6783,N_6942);
and U7373 (N_7373,N_6914,N_6746);
or U7374 (N_7374,N_6999,N_6570);
nor U7375 (N_7375,N_6939,N_6899);
nand U7376 (N_7376,N_6965,N_6650);
or U7377 (N_7377,N_6943,N_6988);
nand U7378 (N_7378,N_6598,N_6759);
nor U7379 (N_7379,N_6579,N_6761);
nor U7380 (N_7380,N_6837,N_6534);
or U7381 (N_7381,N_6932,N_6625);
nor U7382 (N_7382,N_6854,N_6960);
or U7383 (N_7383,N_6516,N_6829);
or U7384 (N_7384,N_6515,N_6878);
nor U7385 (N_7385,N_6837,N_6884);
nor U7386 (N_7386,N_6631,N_6713);
nand U7387 (N_7387,N_6517,N_6521);
or U7388 (N_7388,N_6872,N_6879);
nand U7389 (N_7389,N_6528,N_6847);
or U7390 (N_7390,N_6962,N_6862);
nand U7391 (N_7391,N_6537,N_6680);
or U7392 (N_7392,N_6974,N_6660);
and U7393 (N_7393,N_6701,N_6916);
or U7394 (N_7394,N_6811,N_6537);
or U7395 (N_7395,N_6927,N_6596);
and U7396 (N_7396,N_6813,N_6507);
and U7397 (N_7397,N_6547,N_6553);
nor U7398 (N_7398,N_6552,N_6724);
nand U7399 (N_7399,N_6686,N_6571);
nor U7400 (N_7400,N_6730,N_6678);
nand U7401 (N_7401,N_6906,N_6752);
and U7402 (N_7402,N_6847,N_6930);
nor U7403 (N_7403,N_6945,N_6517);
or U7404 (N_7404,N_6713,N_6960);
nor U7405 (N_7405,N_6834,N_6743);
nand U7406 (N_7406,N_6874,N_6658);
or U7407 (N_7407,N_6724,N_6524);
nor U7408 (N_7408,N_6752,N_6560);
or U7409 (N_7409,N_6930,N_6690);
and U7410 (N_7410,N_6617,N_6831);
nor U7411 (N_7411,N_6547,N_6996);
or U7412 (N_7412,N_6646,N_6517);
or U7413 (N_7413,N_6791,N_6596);
or U7414 (N_7414,N_6876,N_6960);
or U7415 (N_7415,N_6571,N_6841);
nor U7416 (N_7416,N_6580,N_6840);
or U7417 (N_7417,N_6936,N_6821);
nor U7418 (N_7418,N_6639,N_6660);
nor U7419 (N_7419,N_6839,N_6754);
nand U7420 (N_7420,N_6596,N_6607);
and U7421 (N_7421,N_6681,N_6793);
nand U7422 (N_7422,N_6513,N_6950);
and U7423 (N_7423,N_6691,N_6655);
or U7424 (N_7424,N_6761,N_6758);
and U7425 (N_7425,N_6764,N_6732);
or U7426 (N_7426,N_6666,N_6738);
nand U7427 (N_7427,N_6986,N_6735);
nor U7428 (N_7428,N_6675,N_6945);
or U7429 (N_7429,N_6925,N_6594);
or U7430 (N_7430,N_6811,N_6671);
and U7431 (N_7431,N_6881,N_6606);
nor U7432 (N_7432,N_6695,N_6801);
or U7433 (N_7433,N_6874,N_6558);
nand U7434 (N_7434,N_6701,N_6630);
nand U7435 (N_7435,N_6693,N_6986);
or U7436 (N_7436,N_6828,N_6989);
and U7437 (N_7437,N_6693,N_6588);
nand U7438 (N_7438,N_6963,N_6631);
or U7439 (N_7439,N_6828,N_6906);
and U7440 (N_7440,N_6915,N_6553);
and U7441 (N_7441,N_6855,N_6964);
nor U7442 (N_7442,N_6611,N_6603);
nand U7443 (N_7443,N_6892,N_6750);
and U7444 (N_7444,N_6775,N_6971);
nand U7445 (N_7445,N_6657,N_6941);
xor U7446 (N_7446,N_6941,N_6919);
nand U7447 (N_7447,N_6920,N_6579);
nand U7448 (N_7448,N_6783,N_6512);
and U7449 (N_7449,N_6934,N_6722);
nand U7450 (N_7450,N_6652,N_6835);
and U7451 (N_7451,N_6876,N_6952);
nor U7452 (N_7452,N_6566,N_6745);
and U7453 (N_7453,N_6808,N_6721);
nor U7454 (N_7454,N_6531,N_6511);
and U7455 (N_7455,N_6950,N_6890);
and U7456 (N_7456,N_6772,N_6866);
or U7457 (N_7457,N_6758,N_6705);
nand U7458 (N_7458,N_6919,N_6861);
or U7459 (N_7459,N_6792,N_6985);
nor U7460 (N_7460,N_6552,N_6753);
nand U7461 (N_7461,N_6506,N_6540);
nand U7462 (N_7462,N_6525,N_6928);
and U7463 (N_7463,N_6512,N_6625);
nand U7464 (N_7464,N_6589,N_6973);
and U7465 (N_7465,N_6679,N_6964);
nand U7466 (N_7466,N_6911,N_6858);
nor U7467 (N_7467,N_6724,N_6584);
xnor U7468 (N_7468,N_6771,N_6569);
or U7469 (N_7469,N_6680,N_6820);
or U7470 (N_7470,N_6743,N_6916);
and U7471 (N_7471,N_6956,N_6693);
nor U7472 (N_7472,N_6820,N_6892);
nand U7473 (N_7473,N_6527,N_6636);
nand U7474 (N_7474,N_6765,N_6737);
and U7475 (N_7475,N_6966,N_6742);
nand U7476 (N_7476,N_6610,N_6770);
nor U7477 (N_7477,N_6622,N_6833);
or U7478 (N_7478,N_6760,N_6654);
and U7479 (N_7479,N_6714,N_6656);
nor U7480 (N_7480,N_6917,N_6818);
nor U7481 (N_7481,N_6916,N_6667);
nor U7482 (N_7482,N_6654,N_6749);
and U7483 (N_7483,N_6840,N_6868);
and U7484 (N_7484,N_6699,N_6863);
or U7485 (N_7485,N_6758,N_6540);
or U7486 (N_7486,N_6882,N_6655);
nor U7487 (N_7487,N_6611,N_6797);
and U7488 (N_7488,N_6974,N_6567);
nor U7489 (N_7489,N_6610,N_6779);
nor U7490 (N_7490,N_6984,N_6661);
or U7491 (N_7491,N_6966,N_6986);
or U7492 (N_7492,N_6887,N_6897);
or U7493 (N_7493,N_6706,N_6741);
nor U7494 (N_7494,N_6898,N_6593);
and U7495 (N_7495,N_6559,N_6654);
or U7496 (N_7496,N_6594,N_6826);
nand U7497 (N_7497,N_6661,N_6738);
and U7498 (N_7498,N_6539,N_6787);
nor U7499 (N_7499,N_6983,N_6543);
nand U7500 (N_7500,N_7321,N_7226);
or U7501 (N_7501,N_7106,N_7182);
nor U7502 (N_7502,N_7480,N_7407);
nor U7503 (N_7503,N_7108,N_7103);
or U7504 (N_7504,N_7389,N_7039);
nor U7505 (N_7505,N_7285,N_7175);
nor U7506 (N_7506,N_7490,N_7016);
or U7507 (N_7507,N_7339,N_7334);
nand U7508 (N_7508,N_7277,N_7195);
or U7509 (N_7509,N_7345,N_7032);
or U7510 (N_7510,N_7161,N_7413);
nor U7511 (N_7511,N_7074,N_7299);
nand U7512 (N_7512,N_7030,N_7488);
nor U7513 (N_7513,N_7427,N_7440);
nor U7514 (N_7514,N_7010,N_7383);
and U7515 (N_7515,N_7014,N_7150);
nor U7516 (N_7516,N_7335,N_7063);
nor U7517 (N_7517,N_7061,N_7128);
nor U7518 (N_7518,N_7243,N_7473);
nand U7519 (N_7519,N_7127,N_7369);
nor U7520 (N_7520,N_7362,N_7192);
and U7521 (N_7521,N_7004,N_7100);
or U7522 (N_7522,N_7188,N_7041);
or U7523 (N_7523,N_7380,N_7303);
or U7524 (N_7524,N_7002,N_7123);
nand U7525 (N_7525,N_7351,N_7023);
and U7526 (N_7526,N_7064,N_7348);
xnor U7527 (N_7527,N_7132,N_7395);
nor U7528 (N_7528,N_7283,N_7073);
or U7529 (N_7529,N_7008,N_7086);
nand U7530 (N_7530,N_7246,N_7305);
nand U7531 (N_7531,N_7329,N_7197);
nand U7532 (N_7532,N_7149,N_7385);
nand U7533 (N_7533,N_7430,N_7379);
nand U7534 (N_7534,N_7051,N_7291);
nor U7535 (N_7535,N_7131,N_7204);
or U7536 (N_7536,N_7317,N_7095);
or U7537 (N_7537,N_7360,N_7109);
nor U7538 (N_7538,N_7025,N_7286);
or U7539 (N_7539,N_7475,N_7057);
and U7540 (N_7540,N_7352,N_7183);
and U7541 (N_7541,N_7459,N_7037);
nor U7542 (N_7542,N_7212,N_7478);
and U7543 (N_7543,N_7412,N_7307);
and U7544 (N_7544,N_7337,N_7089);
nand U7545 (N_7545,N_7194,N_7421);
and U7546 (N_7546,N_7258,N_7232);
nand U7547 (N_7547,N_7423,N_7444);
or U7548 (N_7548,N_7468,N_7117);
nor U7549 (N_7549,N_7294,N_7198);
nand U7550 (N_7550,N_7304,N_7152);
or U7551 (N_7551,N_7404,N_7344);
and U7552 (N_7552,N_7071,N_7469);
or U7553 (N_7553,N_7203,N_7267);
nor U7554 (N_7554,N_7021,N_7067);
and U7555 (N_7555,N_7436,N_7176);
nand U7556 (N_7556,N_7055,N_7009);
nand U7557 (N_7557,N_7287,N_7392);
nor U7558 (N_7558,N_7384,N_7433);
nand U7559 (N_7559,N_7489,N_7406);
nand U7560 (N_7560,N_7442,N_7264);
or U7561 (N_7561,N_7144,N_7429);
nor U7562 (N_7562,N_7324,N_7330);
or U7563 (N_7563,N_7054,N_7001);
or U7564 (N_7564,N_7116,N_7217);
and U7565 (N_7565,N_7431,N_7377);
nor U7566 (N_7566,N_7015,N_7465);
and U7567 (N_7567,N_7234,N_7235);
or U7568 (N_7568,N_7328,N_7166);
and U7569 (N_7569,N_7457,N_7276);
nand U7570 (N_7570,N_7078,N_7481);
nand U7571 (N_7571,N_7314,N_7419);
nor U7572 (N_7572,N_7196,N_7254);
and U7573 (N_7573,N_7279,N_7233);
nor U7574 (N_7574,N_7134,N_7099);
or U7575 (N_7575,N_7062,N_7047);
or U7576 (N_7576,N_7326,N_7347);
nor U7577 (N_7577,N_7472,N_7027);
nand U7578 (N_7578,N_7318,N_7160);
and U7579 (N_7579,N_7215,N_7236);
nand U7580 (N_7580,N_7292,N_7220);
nor U7581 (N_7581,N_7136,N_7129);
or U7582 (N_7582,N_7297,N_7311);
or U7583 (N_7583,N_7260,N_7340);
nand U7584 (N_7584,N_7388,N_7119);
nor U7585 (N_7585,N_7491,N_7365);
and U7586 (N_7586,N_7155,N_7443);
and U7587 (N_7587,N_7240,N_7168);
nand U7588 (N_7588,N_7088,N_7118);
xor U7589 (N_7589,N_7300,N_7274);
and U7590 (N_7590,N_7044,N_7393);
nand U7591 (N_7591,N_7438,N_7072);
and U7592 (N_7592,N_7474,N_7087);
xor U7593 (N_7593,N_7425,N_7376);
nor U7594 (N_7594,N_7271,N_7422);
nand U7595 (N_7595,N_7482,N_7173);
nor U7596 (N_7596,N_7302,N_7439);
or U7597 (N_7597,N_7239,N_7043);
nor U7598 (N_7598,N_7282,N_7111);
nand U7599 (N_7599,N_7179,N_7206);
nand U7600 (N_7600,N_7202,N_7358);
nor U7601 (N_7601,N_7081,N_7418);
nand U7602 (N_7602,N_7237,N_7434);
or U7603 (N_7603,N_7169,N_7493);
nand U7604 (N_7604,N_7346,N_7060);
and U7605 (N_7605,N_7093,N_7448);
nor U7606 (N_7606,N_7200,N_7333);
nor U7607 (N_7607,N_7479,N_7445);
and U7608 (N_7608,N_7371,N_7091);
nand U7609 (N_7609,N_7263,N_7464);
or U7610 (N_7610,N_7024,N_7193);
and U7611 (N_7611,N_7184,N_7224);
nand U7612 (N_7612,N_7035,N_7484);
nor U7613 (N_7613,N_7495,N_7222);
or U7614 (N_7614,N_7456,N_7415);
and U7615 (N_7615,N_7270,N_7364);
or U7616 (N_7616,N_7387,N_7112);
nor U7617 (N_7617,N_7181,N_7139);
and U7618 (N_7618,N_7363,N_7096);
or U7619 (N_7619,N_7242,N_7293);
or U7620 (N_7620,N_7101,N_7005);
nor U7621 (N_7621,N_7000,N_7121);
or U7622 (N_7622,N_7174,N_7207);
nor U7623 (N_7623,N_7402,N_7244);
nand U7624 (N_7624,N_7467,N_7048);
nand U7625 (N_7625,N_7281,N_7312);
nor U7626 (N_7626,N_7250,N_7097);
or U7627 (N_7627,N_7308,N_7451);
nand U7628 (N_7628,N_7435,N_7114);
nor U7629 (N_7629,N_7403,N_7315);
nand U7630 (N_7630,N_7426,N_7133);
or U7631 (N_7631,N_7007,N_7373);
and U7632 (N_7632,N_7463,N_7447);
or U7633 (N_7633,N_7070,N_7248);
or U7634 (N_7634,N_7449,N_7485);
nor U7635 (N_7635,N_7375,N_7115);
nand U7636 (N_7636,N_7428,N_7068);
nor U7637 (N_7637,N_7390,N_7177);
nand U7638 (N_7638,N_7228,N_7361);
nand U7639 (N_7639,N_7411,N_7147);
and U7640 (N_7640,N_7247,N_7309);
nand U7641 (N_7641,N_7356,N_7110);
and U7642 (N_7642,N_7420,N_7386);
nand U7643 (N_7643,N_7017,N_7408);
nand U7644 (N_7644,N_7059,N_7498);
xor U7645 (N_7645,N_7298,N_7137);
or U7646 (N_7646,N_7381,N_7185);
and U7647 (N_7647,N_7288,N_7049);
and U7648 (N_7648,N_7031,N_7280);
or U7649 (N_7649,N_7083,N_7245);
or U7650 (N_7650,N_7486,N_7253);
nor U7651 (N_7651,N_7320,N_7201);
nand U7652 (N_7652,N_7499,N_7124);
nand U7653 (N_7653,N_7462,N_7210);
nor U7654 (N_7654,N_7125,N_7325);
nand U7655 (N_7655,N_7076,N_7126);
or U7656 (N_7656,N_7350,N_7400);
nand U7657 (N_7657,N_7255,N_7167);
nand U7658 (N_7658,N_7306,N_7164);
or U7659 (N_7659,N_7033,N_7018);
and U7660 (N_7660,N_7045,N_7011);
nor U7661 (N_7661,N_7257,N_7399);
or U7662 (N_7662,N_7209,N_7424);
or U7663 (N_7663,N_7159,N_7322);
nor U7664 (N_7664,N_7343,N_7020);
nand U7665 (N_7665,N_7219,N_7158);
and U7666 (N_7666,N_7432,N_7275);
and U7667 (N_7667,N_7251,N_7278);
or U7668 (N_7668,N_7261,N_7187);
or U7669 (N_7669,N_7476,N_7098);
nand U7670 (N_7670,N_7441,N_7289);
and U7671 (N_7671,N_7122,N_7437);
nand U7672 (N_7672,N_7148,N_7162);
and U7673 (N_7673,N_7466,N_7138);
nor U7674 (N_7674,N_7120,N_7417);
nand U7675 (N_7675,N_7310,N_7113);
or U7676 (N_7676,N_7216,N_7256);
nand U7677 (N_7677,N_7022,N_7229);
nand U7678 (N_7678,N_7266,N_7370);
or U7679 (N_7679,N_7178,N_7130);
and U7680 (N_7680,N_7084,N_7382);
and U7681 (N_7681,N_7012,N_7050);
nand U7682 (N_7682,N_7218,N_7401);
and U7683 (N_7683,N_7273,N_7367);
nand U7684 (N_7684,N_7189,N_7082);
or U7685 (N_7685,N_7191,N_7378);
nor U7686 (N_7686,N_7213,N_7461);
nand U7687 (N_7687,N_7156,N_7231);
and U7688 (N_7688,N_7042,N_7446);
and U7689 (N_7689,N_7332,N_7496);
or U7690 (N_7690,N_7450,N_7214);
or U7691 (N_7691,N_7006,N_7301);
nor U7692 (N_7692,N_7165,N_7066);
nor U7693 (N_7693,N_7470,N_7458);
and U7694 (N_7694,N_7397,N_7105);
and U7695 (N_7695,N_7336,N_7368);
nand U7696 (N_7696,N_7157,N_7085);
nor U7697 (N_7697,N_7092,N_7452);
nand U7698 (N_7698,N_7026,N_7040);
or U7699 (N_7699,N_7141,N_7034);
or U7700 (N_7700,N_7142,N_7268);
nand U7701 (N_7701,N_7455,N_7259);
nor U7702 (N_7702,N_7038,N_7241);
nand U7703 (N_7703,N_7075,N_7205);
nand U7704 (N_7704,N_7230,N_7028);
nor U7705 (N_7705,N_7341,N_7372);
and U7706 (N_7706,N_7331,N_7225);
and U7707 (N_7707,N_7079,N_7053);
or U7708 (N_7708,N_7353,N_7077);
or U7709 (N_7709,N_7454,N_7180);
nor U7710 (N_7710,N_7190,N_7398);
and U7711 (N_7711,N_7410,N_7252);
and U7712 (N_7712,N_7477,N_7327);
nor U7713 (N_7713,N_7295,N_7163);
nor U7714 (N_7714,N_7223,N_7296);
nor U7715 (N_7715,N_7227,N_7019);
nor U7716 (N_7716,N_7265,N_7069);
nand U7717 (N_7717,N_7357,N_7140);
nor U7718 (N_7718,N_7453,N_7284);
nor U7719 (N_7719,N_7396,N_7354);
nor U7720 (N_7720,N_7094,N_7414);
nor U7721 (N_7721,N_7013,N_7374);
nand U7722 (N_7722,N_7146,N_7221);
nand U7723 (N_7723,N_7366,N_7153);
or U7724 (N_7724,N_7080,N_7065);
nor U7725 (N_7725,N_7409,N_7143);
or U7726 (N_7726,N_7186,N_7391);
nand U7727 (N_7727,N_7249,N_7211);
nor U7728 (N_7728,N_7290,N_7172);
nor U7729 (N_7729,N_7170,N_7262);
nor U7730 (N_7730,N_7171,N_7056);
nor U7731 (N_7731,N_7349,N_7208);
nor U7732 (N_7732,N_7046,N_7102);
nor U7733 (N_7733,N_7497,N_7003);
nor U7734 (N_7734,N_7272,N_7145);
or U7735 (N_7735,N_7492,N_7342);
or U7736 (N_7736,N_7323,N_7107);
nor U7737 (N_7737,N_7316,N_7487);
or U7738 (N_7738,N_7394,N_7338);
or U7739 (N_7739,N_7052,N_7460);
nor U7740 (N_7740,N_7029,N_7355);
or U7741 (N_7741,N_7319,N_7416);
or U7742 (N_7742,N_7199,N_7483);
or U7743 (N_7743,N_7154,N_7090);
nor U7744 (N_7744,N_7359,N_7238);
or U7745 (N_7745,N_7036,N_7151);
and U7746 (N_7746,N_7104,N_7135);
nand U7747 (N_7747,N_7313,N_7471);
or U7748 (N_7748,N_7494,N_7058);
or U7749 (N_7749,N_7269,N_7405);
nor U7750 (N_7750,N_7330,N_7174);
and U7751 (N_7751,N_7092,N_7082);
or U7752 (N_7752,N_7137,N_7251);
nand U7753 (N_7753,N_7360,N_7182);
and U7754 (N_7754,N_7286,N_7181);
and U7755 (N_7755,N_7112,N_7371);
nand U7756 (N_7756,N_7306,N_7213);
nand U7757 (N_7757,N_7092,N_7233);
or U7758 (N_7758,N_7154,N_7331);
and U7759 (N_7759,N_7498,N_7322);
nor U7760 (N_7760,N_7052,N_7423);
nand U7761 (N_7761,N_7041,N_7301);
nor U7762 (N_7762,N_7166,N_7366);
nor U7763 (N_7763,N_7001,N_7216);
nand U7764 (N_7764,N_7113,N_7454);
or U7765 (N_7765,N_7013,N_7159);
nand U7766 (N_7766,N_7372,N_7036);
or U7767 (N_7767,N_7257,N_7444);
and U7768 (N_7768,N_7149,N_7283);
nor U7769 (N_7769,N_7038,N_7406);
nand U7770 (N_7770,N_7456,N_7203);
or U7771 (N_7771,N_7126,N_7281);
or U7772 (N_7772,N_7041,N_7316);
and U7773 (N_7773,N_7048,N_7292);
nand U7774 (N_7774,N_7437,N_7213);
nor U7775 (N_7775,N_7275,N_7391);
or U7776 (N_7776,N_7099,N_7422);
or U7777 (N_7777,N_7156,N_7254);
nor U7778 (N_7778,N_7158,N_7194);
or U7779 (N_7779,N_7391,N_7193);
and U7780 (N_7780,N_7310,N_7464);
nand U7781 (N_7781,N_7451,N_7145);
nor U7782 (N_7782,N_7350,N_7394);
nand U7783 (N_7783,N_7484,N_7415);
nand U7784 (N_7784,N_7336,N_7077);
nand U7785 (N_7785,N_7242,N_7364);
nor U7786 (N_7786,N_7134,N_7284);
nand U7787 (N_7787,N_7286,N_7247);
nand U7788 (N_7788,N_7133,N_7321);
and U7789 (N_7789,N_7468,N_7429);
nor U7790 (N_7790,N_7135,N_7368);
and U7791 (N_7791,N_7057,N_7409);
or U7792 (N_7792,N_7317,N_7222);
nor U7793 (N_7793,N_7168,N_7305);
and U7794 (N_7794,N_7455,N_7358);
nand U7795 (N_7795,N_7174,N_7115);
nor U7796 (N_7796,N_7080,N_7331);
and U7797 (N_7797,N_7311,N_7209);
nor U7798 (N_7798,N_7131,N_7180);
nand U7799 (N_7799,N_7364,N_7000);
nor U7800 (N_7800,N_7471,N_7331);
and U7801 (N_7801,N_7161,N_7094);
or U7802 (N_7802,N_7297,N_7072);
nand U7803 (N_7803,N_7488,N_7086);
and U7804 (N_7804,N_7111,N_7083);
nor U7805 (N_7805,N_7188,N_7444);
nor U7806 (N_7806,N_7257,N_7483);
and U7807 (N_7807,N_7302,N_7498);
or U7808 (N_7808,N_7355,N_7119);
nor U7809 (N_7809,N_7455,N_7395);
and U7810 (N_7810,N_7265,N_7161);
nor U7811 (N_7811,N_7257,N_7392);
and U7812 (N_7812,N_7084,N_7398);
nor U7813 (N_7813,N_7257,N_7404);
xor U7814 (N_7814,N_7179,N_7061);
or U7815 (N_7815,N_7150,N_7277);
and U7816 (N_7816,N_7254,N_7242);
or U7817 (N_7817,N_7247,N_7362);
nand U7818 (N_7818,N_7114,N_7348);
or U7819 (N_7819,N_7023,N_7062);
nor U7820 (N_7820,N_7225,N_7418);
nor U7821 (N_7821,N_7320,N_7168);
and U7822 (N_7822,N_7486,N_7162);
nand U7823 (N_7823,N_7388,N_7167);
and U7824 (N_7824,N_7392,N_7110);
nand U7825 (N_7825,N_7085,N_7337);
nor U7826 (N_7826,N_7352,N_7267);
nand U7827 (N_7827,N_7412,N_7133);
and U7828 (N_7828,N_7462,N_7192);
or U7829 (N_7829,N_7397,N_7125);
nor U7830 (N_7830,N_7027,N_7250);
and U7831 (N_7831,N_7269,N_7191);
nor U7832 (N_7832,N_7158,N_7112);
or U7833 (N_7833,N_7428,N_7298);
or U7834 (N_7834,N_7100,N_7279);
nor U7835 (N_7835,N_7320,N_7025);
or U7836 (N_7836,N_7286,N_7329);
nor U7837 (N_7837,N_7244,N_7397);
nor U7838 (N_7838,N_7413,N_7256);
or U7839 (N_7839,N_7136,N_7108);
or U7840 (N_7840,N_7354,N_7276);
nor U7841 (N_7841,N_7453,N_7426);
and U7842 (N_7842,N_7274,N_7178);
nor U7843 (N_7843,N_7080,N_7308);
nand U7844 (N_7844,N_7078,N_7141);
nand U7845 (N_7845,N_7419,N_7020);
nor U7846 (N_7846,N_7096,N_7150);
or U7847 (N_7847,N_7398,N_7086);
nor U7848 (N_7848,N_7010,N_7020);
nand U7849 (N_7849,N_7248,N_7456);
and U7850 (N_7850,N_7252,N_7036);
nor U7851 (N_7851,N_7447,N_7087);
nand U7852 (N_7852,N_7173,N_7198);
or U7853 (N_7853,N_7054,N_7162);
nor U7854 (N_7854,N_7483,N_7466);
nand U7855 (N_7855,N_7141,N_7239);
nor U7856 (N_7856,N_7466,N_7210);
nor U7857 (N_7857,N_7219,N_7427);
and U7858 (N_7858,N_7055,N_7358);
and U7859 (N_7859,N_7063,N_7491);
nand U7860 (N_7860,N_7215,N_7396);
and U7861 (N_7861,N_7361,N_7359);
nor U7862 (N_7862,N_7167,N_7353);
and U7863 (N_7863,N_7200,N_7164);
nand U7864 (N_7864,N_7032,N_7001);
or U7865 (N_7865,N_7178,N_7374);
or U7866 (N_7866,N_7229,N_7039);
or U7867 (N_7867,N_7172,N_7104);
nand U7868 (N_7868,N_7368,N_7406);
nand U7869 (N_7869,N_7381,N_7297);
nor U7870 (N_7870,N_7082,N_7004);
nor U7871 (N_7871,N_7422,N_7214);
or U7872 (N_7872,N_7499,N_7210);
or U7873 (N_7873,N_7145,N_7291);
or U7874 (N_7874,N_7178,N_7263);
nand U7875 (N_7875,N_7450,N_7408);
nor U7876 (N_7876,N_7014,N_7445);
or U7877 (N_7877,N_7454,N_7199);
nand U7878 (N_7878,N_7092,N_7102);
or U7879 (N_7879,N_7186,N_7416);
nor U7880 (N_7880,N_7211,N_7159);
or U7881 (N_7881,N_7495,N_7045);
nor U7882 (N_7882,N_7238,N_7017);
or U7883 (N_7883,N_7044,N_7319);
or U7884 (N_7884,N_7054,N_7400);
nor U7885 (N_7885,N_7238,N_7164);
nor U7886 (N_7886,N_7284,N_7430);
nand U7887 (N_7887,N_7404,N_7037);
or U7888 (N_7888,N_7267,N_7122);
nor U7889 (N_7889,N_7376,N_7347);
or U7890 (N_7890,N_7439,N_7077);
nor U7891 (N_7891,N_7003,N_7221);
nand U7892 (N_7892,N_7246,N_7227);
nor U7893 (N_7893,N_7489,N_7445);
nor U7894 (N_7894,N_7003,N_7030);
and U7895 (N_7895,N_7292,N_7343);
or U7896 (N_7896,N_7020,N_7477);
nand U7897 (N_7897,N_7342,N_7041);
nor U7898 (N_7898,N_7325,N_7414);
and U7899 (N_7899,N_7166,N_7193);
nor U7900 (N_7900,N_7482,N_7204);
nor U7901 (N_7901,N_7005,N_7113);
and U7902 (N_7902,N_7467,N_7339);
or U7903 (N_7903,N_7162,N_7361);
and U7904 (N_7904,N_7092,N_7404);
or U7905 (N_7905,N_7247,N_7377);
nand U7906 (N_7906,N_7362,N_7184);
nand U7907 (N_7907,N_7080,N_7105);
or U7908 (N_7908,N_7492,N_7069);
nand U7909 (N_7909,N_7305,N_7091);
or U7910 (N_7910,N_7285,N_7382);
or U7911 (N_7911,N_7279,N_7204);
or U7912 (N_7912,N_7370,N_7393);
or U7913 (N_7913,N_7177,N_7234);
nand U7914 (N_7914,N_7131,N_7396);
nand U7915 (N_7915,N_7174,N_7249);
or U7916 (N_7916,N_7091,N_7245);
nor U7917 (N_7917,N_7167,N_7470);
or U7918 (N_7918,N_7380,N_7455);
nand U7919 (N_7919,N_7220,N_7360);
or U7920 (N_7920,N_7313,N_7457);
nor U7921 (N_7921,N_7005,N_7356);
nor U7922 (N_7922,N_7187,N_7424);
or U7923 (N_7923,N_7003,N_7224);
nor U7924 (N_7924,N_7055,N_7208);
and U7925 (N_7925,N_7057,N_7111);
nor U7926 (N_7926,N_7471,N_7172);
nand U7927 (N_7927,N_7159,N_7106);
and U7928 (N_7928,N_7488,N_7492);
and U7929 (N_7929,N_7259,N_7210);
nor U7930 (N_7930,N_7015,N_7277);
nand U7931 (N_7931,N_7376,N_7387);
or U7932 (N_7932,N_7086,N_7074);
or U7933 (N_7933,N_7172,N_7226);
nor U7934 (N_7934,N_7476,N_7287);
nor U7935 (N_7935,N_7436,N_7020);
or U7936 (N_7936,N_7278,N_7138);
or U7937 (N_7937,N_7271,N_7364);
nor U7938 (N_7938,N_7027,N_7110);
or U7939 (N_7939,N_7088,N_7349);
nand U7940 (N_7940,N_7434,N_7265);
nor U7941 (N_7941,N_7292,N_7172);
nand U7942 (N_7942,N_7369,N_7088);
nand U7943 (N_7943,N_7327,N_7391);
and U7944 (N_7944,N_7139,N_7082);
or U7945 (N_7945,N_7248,N_7462);
and U7946 (N_7946,N_7282,N_7377);
or U7947 (N_7947,N_7302,N_7191);
nand U7948 (N_7948,N_7438,N_7138);
and U7949 (N_7949,N_7204,N_7038);
nor U7950 (N_7950,N_7424,N_7031);
nor U7951 (N_7951,N_7351,N_7266);
nand U7952 (N_7952,N_7102,N_7458);
or U7953 (N_7953,N_7038,N_7095);
or U7954 (N_7954,N_7199,N_7263);
and U7955 (N_7955,N_7424,N_7296);
xnor U7956 (N_7956,N_7239,N_7277);
or U7957 (N_7957,N_7092,N_7492);
and U7958 (N_7958,N_7155,N_7389);
nand U7959 (N_7959,N_7264,N_7448);
or U7960 (N_7960,N_7084,N_7165);
nand U7961 (N_7961,N_7493,N_7033);
or U7962 (N_7962,N_7152,N_7498);
nand U7963 (N_7963,N_7362,N_7155);
nor U7964 (N_7964,N_7034,N_7086);
or U7965 (N_7965,N_7157,N_7480);
nor U7966 (N_7966,N_7450,N_7466);
and U7967 (N_7967,N_7109,N_7034);
and U7968 (N_7968,N_7187,N_7297);
or U7969 (N_7969,N_7416,N_7080);
nand U7970 (N_7970,N_7041,N_7165);
nand U7971 (N_7971,N_7098,N_7191);
or U7972 (N_7972,N_7122,N_7013);
and U7973 (N_7973,N_7074,N_7104);
nor U7974 (N_7974,N_7207,N_7049);
or U7975 (N_7975,N_7458,N_7261);
and U7976 (N_7976,N_7246,N_7383);
or U7977 (N_7977,N_7013,N_7021);
or U7978 (N_7978,N_7103,N_7181);
nand U7979 (N_7979,N_7228,N_7063);
or U7980 (N_7980,N_7372,N_7163);
nor U7981 (N_7981,N_7397,N_7216);
and U7982 (N_7982,N_7324,N_7076);
nor U7983 (N_7983,N_7451,N_7282);
nand U7984 (N_7984,N_7221,N_7338);
nand U7985 (N_7985,N_7335,N_7385);
nor U7986 (N_7986,N_7002,N_7154);
or U7987 (N_7987,N_7293,N_7165);
and U7988 (N_7988,N_7490,N_7359);
nor U7989 (N_7989,N_7402,N_7263);
and U7990 (N_7990,N_7132,N_7443);
nor U7991 (N_7991,N_7470,N_7129);
nor U7992 (N_7992,N_7151,N_7056);
or U7993 (N_7993,N_7328,N_7385);
or U7994 (N_7994,N_7078,N_7443);
or U7995 (N_7995,N_7265,N_7255);
nor U7996 (N_7996,N_7211,N_7305);
nor U7997 (N_7997,N_7329,N_7470);
xor U7998 (N_7998,N_7144,N_7448);
nor U7999 (N_7999,N_7152,N_7038);
nand U8000 (N_8000,N_7645,N_7769);
nor U8001 (N_8001,N_7929,N_7750);
nor U8002 (N_8002,N_7790,N_7913);
nand U8003 (N_8003,N_7702,N_7888);
nor U8004 (N_8004,N_7744,N_7643);
or U8005 (N_8005,N_7547,N_7897);
and U8006 (N_8006,N_7555,N_7705);
and U8007 (N_8007,N_7628,N_7746);
and U8008 (N_8008,N_7821,N_7610);
or U8009 (N_8009,N_7721,N_7908);
nor U8010 (N_8010,N_7654,N_7681);
and U8011 (N_8011,N_7999,N_7672);
nand U8012 (N_8012,N_7581,N_7983);
or U8013 (N_8013,N_7567,N_7529);
and U8014 (N_8014,N_7539,N_7737);
or U8015 (N_8015,N_7520,N_7509);
or U8016 (N_8016,N_7601,N_7896);
and U8017 (N_8017,N_7798,N_7950);
or U8018 (N_8018,N_7851,N_7518);
or U8019 (N_8019,N_7876,N_7587);
or U8020 (N_8020,N_7638,N_7833);
and U8021 (N_8021,N_7840,N_7611);
or U8022 (N_8022,N_7909,N_7505);
nor U8023 (N_8023,N_7782,N_7847);
nor U8024 (N_8024,N_7716,N_7531);
nand U8025 (N_8025,N_7685,N_7934);
or U8026 (N_8026,N_7784,N_7937);
or U8027 (N_8027,N_7859,N_7642);
nand U8028 (N_8028,N_7893,N_7964);
nand U8029 (N_8029,N_7920,N_7626);
nor U8030 (N_8030,N_7924,N_7959);
or U8031 (N_8031,N_7836,N_7564);
nor U8032 (N_8032,N_7513,N_7571);
and U8033 (N_8033,N_7994,N_7582);
nand U8034 (N_8034,N_7646,N_7624);
or U8035 (N_8035,N_7771,N_7886);
nor U8036 (N_8036,N_7917,N_7770);
nand U8037 (N_8037,N_7548,N_7939);
and U8038 (N_8038,N_7807,N_7993);
nor U8039 (N_8039,N_7545,N_7900);
nor U8040 (N_8040,N_7868,N_7933);
nand U8041 (N_8041,N_7714,N_7965);
and U8042 (N_8042,N_7560,N_7764);
and U8043 (N_8043,N_7891,N_7528);
and U8044 (N_8044,N_7941,N_7792);
nor U8045 (N_8045,N_7542,N_7992);
and U8046 (N_8046,N_7817,N_7752);
and U8047 (N_8047,N_7818,N_7748);
nand U8048 (N_8048,N_7967,N_7803);
or U8049 (N_8049,N_7627,N_7591);
or U8050 (N_8050,N_7565,N_7892);
or U8051 (N_8051,N_7780,N_7802);
and U8052 (N_8052,N_7641,N_7691);
and U8053 (N_8053,N_7731,N_7856);
nor U8054 (N_8054,N_7887,N_7980);
or U8055 (N_8055,N_7953,N_7512);
nor U8056 (N_8056,N_7905,N_7594);
and U8057 (N_8057,N_7596,N_7569);
nor U8058 (N_8058,N_7867,N_7903);
or U8059 (N_8059,N_7898,N_7508);
xor U8060 (N_8060,N_7558,N_7753);
or U8061 (N_8061,N_7864,N_7546);
and U8062 (N_8062,N_7741,N_7614);
nand U8063 (N_8063,N_7515,N_7830);
nand U8064 (N_8064,N_7815,N_7604);
nor U8065 (N_8065,N_7541,N_7793);
nand U8066 (N_8066,N_7609,N_7843);
nor U8067 (N_8067,N_7969,N_7580);
or U8068 (N_8068,N_7814,N_7561);
and U8069 (N_8069,N_7837,N_7944);
or U8070 (N_8070,N_7577,N_7701);
and U8071 (N_8071,N_7844,N_7592);
nor U8072 (N_8072,N_7789,N_7975);
and U8073 (N_8073,N_7633,N_7979);
and U8074 (N_8074,N_7772,N_7831);
and U8075 (N_8075,N_7668,N_7507);
or U8076 (N_8076,N_7730,N_7940);
or U8077 (N_8077,N_7958,N_7535);
or U8078 (N_8078,N_7576,N_7689);
and U8079 (N_8079,N_7516,N_7514);
or U8080 (N_8080,N_7759,N_7679);
or U8081 (N_8081,N_7754,N_7718);
or U8082 (N_8082,N_7931,N_7922);
or U8083 (N_8083,N_7595,N_7794);
or U8084 (N_8084,N_7726,N_7823);
and U8085 (N_8085,N_7534,N_7540);
nand U8086 (N_8086,N_7848,N_7796);
or U8087 (N_8087,N_7707,N_7862);
or U8088 (N_8088,N_7630,N_7998);
xor U8089 (N_8089,N_7544,N_7727);
nand U8090 (N_8090,N_7952,N_7563);
and U8091 (N_8091,N_7788,N_7625);
nor U8092 (N_8092,N_7733,N_7756);
nor U8093 (N_8093,N_7674,N_7678);
nor U8094 (N_8094,N_7620,N_7504);
nand U8095 (N_8095,N_7890,N_7957);
and U8096 (N_8096,N_7901,N_7760);
and U8097 (N_8097,N_7751,N_7656);
and U8098 (N_8098,N_7666,N_7910);
nand U8099 (N_8099,N_7526,N_7806);
nor U8100 (N_8100,N_7974,N_7826);
nand U8101 (N_8101,N_7524,N_7570);
and U8102 (N_8102,N_7602,N_7961);
nor U8103 (N_8103,N_7574,N_7631);
and U8104 (N_8104,N_7945,N_7606);
nor U8105 (N_8105,N_7568,N_7828);
xor U8106 (N_8106,N_7774,N_7777);
nor U8107 (N_8107,N_7522,N_7651);
or U8108 (N_8108,N_7849,N_7720);
and U8109 (N_8109,N_7935,N_7942);
and U8110 (N_8110,N_7882,N_7584);
and U8111 (N_8111,N_7525,N_7805);
nor U8112 (N_8112,N_7763,N_7977);
or U8113 (N_8113,N_7676,N_7599);
and U8114 (N_8114,N_7981,N_7600);
and U8115 (N_8115,N_7928,N_7550);
and U8116 (N_8116,N_7842,N_7855);
and U8117 (N_8117,N_7879,N_7801);
nand U8118 (N_8118,N_7682,N_7517);
nor U8119 (N_8119,N_7543,N_7810);
and U8120 (N_8120,N_7578,N_7736);
or U8121 (N_8121,N_7549,N_7621);
nand U8122 (N_8122,N_7647,N_7809);
nand U8123 (N_8123,N_7659,N_7838);
nand U8124 (N_8124,N_7966,N_7503);
nand U8125 (N_8125,N_7527,N_7575);
or U8126 (N_8126,N_7846,N_7536);
nand U8127 (N_8127,N_7991,N_7749);
nor U8128 (N_8128,N_7811,N_7692);
nand U8129 (N_8129,N_7703,N_7704);
and U8130 (N_8130,N_7747,N_7552);
and U8131 (N_8131,N_7938,N_7834);
nor U8132 (N_8132,N_7743,N_7955);
and U8133 (N_8133,N_7853,N_7972);
and U8134 (N_8134,N_7661,N_7889);
and U8135 (N_8135,N_7664,N_7511);
nor U8136 (N_8136,N_7779,N_7786);
nand U8137 (N_8137,N_7962,N_7634);
nand U8138 (N_8138,N_7717,N_7783);
or U8139 (N_8139,N_7916,N_7655);
and U8140 (N_8140,N_7841,N_7884);
nor U8141 (N_8141,N_7919,N_7506);
and U8142 (N_8142,N_7878,N_7537);
and U8143 (N_8143,N_7532,N_7554);
or U8144 (N_8144,N_7766,N_7662);
or U8145 (N_8145,N_7861,N_7593);
nand U8146 (N_8146,N_7925,N_7835);
or U8147 (N_8147,N_7694,N_7711);
nand U8148 (N_8148,N_7735,N_7700);
nor U8149 (N_8149,N_7715,N_7710);
nor U8150 (N_8150,N_7667,N_7758);
nand U8151 (N_8151,N_7765,N_7573);
and U8152 (N_8152,N_7871,N_7971);
nand U8153 (N_8153,N_7649,N_7881);
and U8154 (N_8154,N_7684,N_7800);
nor U8155 (N_8155,N_7985,N_7742);
nand U8156 (N_8156,N_7899,N_7616);
and U8157 (N_8157,N_7644,N_7869);
and U8158 (N_8158,N_7551,N_7995);
and U8159 (N_8159,N_7686,N_7812);
or U8160 (N_8160,N_7724,N_7530);
or U8161 (N_8161,N_7863,N_7822);
nand U8162 (N_8162,N_7617,N_7894);
nand U8163 (N_8163,N_7956,N_7732);
nor U8164 (N_8164,N_7845,N_7880);
or U8165 (N_8165,N_7926,N_7865);
nor U8166 (N_8166,N_7559,N_7723);
nand U8167 (N_8167,N_7619,N_7607);
or U8168 (N_8168,N_7671,N_7603);
nor U8169 (N_8169,N_7728,N_7739);
or U8170 (N_8170,N_7875,N_7585);
or U8171 (N_8171,N_7708,N_7658);
nand U8172 (N_8172,N_7930,N_7990);
nor U8173 (N_8173,N_7857,N_7533);
and U8174 (N_8174,N_7827,N_7829);
nor U8175 (N_8175,N_7706,N_7820);
and U8176 (N_8176,N_7877,N_7768);
or U8177 (N_8177,N_7523,N_7698);
or U8178 (N_8178,N_7673,N_7885);
nor U8179 (N_8179,N_7612,N_7590);
or U8180 (N_8180,N_7816,N_7874);
nor U8181 (N_8181,N_7613,N_7761);
nand U8182 (N_8182,N_7745,N_7623);
or U8183 (N_8183,N_7914,N_7648);
nand U8184 (N_8184,N_7719,N_7615);
nand U8185 (N_8185,N_7781,N_7813);
nor U8186 (N_8186,N_7997,N_7787);
nor U8187 (N_8187,N_7932,N_7713);
nand U8188 (N_8188,N_7973,N_7819);
or U8189 (N_8189,N_7947,N_7553);
and U8190 (N_8190,N_7943,N_7677);
nand U8191 (N_8191,N_7775,N_7968);
nor U8192 (N_8192,N_7636,N_7688);
nor U8193 (N_8193,N_7669,N_7722);
and U8194 (N_8194,N_7776,N_7556);
or U8195 (N_8195,N_7767,N_7906);
nor U8196 (N_8196,N_7927,N_7637);
or U8197 (N_8197,N_7911,N_7665);
nand U8198 (N_8198,N_7653,N_7699);
nor U8199 (N_8199,N_7895,N_7729);
and U8200 (N_8200,N_7912,N_7832);
nor U8201 (N_8201,N_7663,N_7850);
xor U8202 (N_8202,N_7650,N_7954);
or U8203 (N_8203,N_7687,N_7936);
and U8204 (N_8204,N_7709,N_7510);
nor U8205 (N_8205,N_7618,N_7680);
nand U8206 (N_8206,N_7872,N_7635);
and U8207 (N_8207,N_7629,N_7639);
or U8208 (N_8208,N_7572,N_7923);
nor U8209 (N_8209,N_7566,N_7597);
nor U8210 (N_8210,N_7799,N_7740);
or U8211 (N_8211,N_7873,N_7804);
nor U8212 (N_8212,N_7948,N_7984);
nor U8213 (N_8213,N_7502,N_7734);
nor U8214 (N_8214,N_7946,N_7963);
nand U8215 (N_8215,N_7951,N_7918);
nand U8216 (N_8216,N_7996,N_7632);
nand U8217 (N_8217,N_7660,N_7583);
nand U8218 (N_8218,N_7738,N_7670);
nand U8219 (N_8219,N_7852,N_7622);
or U8220 (N_8220,N_7712,N_7683);
or U8221 (N_8221,N_7960,N_7860);
or U8222 (N_8222,N_7608,N_7725);
or U8223 (N_8223,N_7989,N_7640);
nand U8224 (N_8224,N_7588,N_7825);
and U8225 (N_8225,N_7988,N_7866);
nor U8226 (N_8226,N_7824,N_7986);
nor U8227 (N_8227,N_7605,N_7907);
nor U8228 (N_8228,N_7778,N_7755);
and U8229 (N_8229,N_7652,N_7538);
or U8230 (N_8230,N_7675,N_7902);
nand U8231 (N_8231,N_7987,N_7795);
nand U8232 (N_8232,N_7808,N_7501);
and U8233 (N_8233,N_7904,N_7978);
nand U8234 (N_8234,N_7970,N_7690);
and U8235 (N_8235,N_7949,N_7839);
and U8236 (N_8236,N_7773,N_7695);
and U8237 (N_8237,N_7757,N_7521);
and U8238 (N_8238,N_7797,N_7915);
nor U8239 (N_8239,N_7589,N_7982);
nand U8240 (N_8240,N_7693,N_7598);
and U8241 (N_8241,N_7562,N_7785);
and U8242 (N_8242,N_7791,N_7519);
and U8243 (N_8243,N_7657,N_7500);
or U8244 (N_8244,N_7854,N_7762);
and U8245 (N_8245,N_7858,N_7696);
or U8246 (N_8246,N_7870,N_7697);
nor U8247 (N_8247,N_7976,N_7883);
or U8248 (N_8248,N_7579,N_7557);
nor U8249 (N_8249,N_7921,N_7586);
nor U8250 (N_8250,N_7711,N_7988);
xor U8251 (N_8251,N_7545,N_7996);
nand U8252 (N_8252,N_7517,N_7550);
and U8253 (N_8253,N_7657,N_7853);
nand U8254 (N_8254,N_7842,N_7957);
or U8255 (N_8255,N_7609,N_7723);
nor U8256 (N_8256,N_7545,N_7642);
nor U8257 (N_8257,N_7595,N_7752);
nand U8258 (N_8258,N_7796,N_7611);
and U8259 (N_8259,N_7800,N_7825);
or U8260 (N_8260,N_7875,N_7725);
and U8261 (N_8261,N_7525,N_7915);
nor U8262 (N_8262,N_7656,N_7604);
nand U8263 (N_8263,N_7581,N_7885);
nand U8264 (N_8264,N_7965,N_7647);
nor U8265 (N_8265,N_7602,N_7683);
and U8266 (N_8266,N_7842,N_7909);
and U8267 (N_8267,N_7732,N_7867);
nor U8268 (N_8268,N_7745,N_7509);
or U8269 (N_8269,N_7697,N_7696);
or U8270 (N_8270,N_7701,N_7906);
nand U8271 (N_8271,N_7616,N_7602);
and U8272 (N_8272,N_7958,N_7926);
nor U8273 (N_8273,N_7963,N_7558);
or U8274 (N_8274,N_7637,N_7815);
nor U8275 (N_8275,N_7627,N_7812);
nand U8276 (N_8276,N_7505,N_7969);
nand U8277 (N_8277,N_7525,N_7737);
nor U8278 (N_8278,N_7731,N_7532);
and U8279 (N_8279,N_7765,N_7770);
and U8280 (N_8280,N_7889,N_7594);
and U8281 (N_8281,N_7805,N_7990);
and U8282 (N_8282,N_7731,N_7582);
nand U8283 (N_8283,N_7803,N_7664);
and U8284 (N_8284,N_7544,N_7887);
and U8285 (N_8285,N_7738,N_7741);
nor U8286 (N_8286,N_7949,N_7519);
or U8287 (N_8287,N_7516,N_7571);
nor U8288 (N_8288,N_7912,N_7693);
or U8289 (N_8289,N_7773,N_7734);
nand U8290 (N_8290,N_7786,N_7653);
nand U8291 (N_8291,N_7775,N_7700);
nor U8292 (N_8292,N_7923,N_7629);
nand U8293 (N_8293,N_7700,N_7965);
or U8294 (N_8294,N_7685,N_7966);
or U8295 (N_8295,N_7545,N_7584);
nor U8296 (N_8296,N_7680,N_7518);
nand U8297 (N_8297,N_7664,N_7793);
and U8298 (N_8298,N_7981,N_7987);
nand U8299 (N_8299,N_7783,N_7810);
nand U8300 (N_8300,N_7637,N_7534);
and U8301 (N_8301,N_7806,N_7729);
and U8302 (N_8302,N_7878,N_7581);
or U8303 (N_8303,N_7854,N_7608);
and U8304 (N_8304,N_7554,N_7675);
or U8305 (N_8305,N_7839,N_7961);
or U8306 (N_8306,N_7853,N_7518);
and U8307 (N_8307,N_7986,N_7594);
nand U8308 (N_8308,N_7689,N_7603);
nor U8309 (N_8309,N_7709,N_7557);
nor U8310 (N_8310,N_7525,N_7610);
nand U8311 (N_8311,N_7691,N_7964);
nand U8312 (N_8312,N_7957,N_7930);
nand U8313 (N_8313,N_7658,N_7809);
or U8314 (N_8314,N_7949,N_7730);
or U8315 (N_8315,N_7517,N_7904);
nor U8316 (N_8316,N_7548,N_7946);
nor U8317 (N_8317,N_7623,N_7879);
or U8318 (N_8318,N_7996,N_7826);
nor U8319 (N_8319,N_7565,N_7920);
and U8320 (N_8320,N_7917,N_7672);
nor U8321 (N_8321,N_7836,N_7806);
nand U8322 (N_8322,N_7677,N_7795);
nand U8323 (N_8323,N_7535,N_7885);
nand U8324 (N_8324,N_7771,N_7729);
nor U8325 (N_8325,N_7734,N_7653);
nor U8326 (N_8326,N_7594,N_7763);
or U8327 (N_8327,N_7730,N_7847);
or U8328 (N_8328,N_7590,N_7966);
and U8329 (N_8329,N_7658,N_7850);
and U8330 (N_8330,N_7698,N_7773);
nor U8331 (N_8331,N_7753,N_7584);
or U8332 (N_8332,N_7752,N_7609);
nor U8333 (N_8333,N_7640,N_7568);
or U8334 (N_8334,N_7617,N_7682);
and U8335 (N_8335,N_7863,N_7883);
nand U8336 (N_8336,N_7695,N_7698);
nor U8337 (N_8337,N_7656,N_7624);
nand U8338 (N_8338,N_7904,N_7649);
or U8339 (N_8339,N_7889,N_7656);
nand U8340 (N_8340,N_7510,N_7970);
xor U8341 (N_8341,N_7862,N_7795);
or U8342 (N_8342,N_7728,N_7551);
nor U8343 (N_8343,N_7986,N_7851);
and U8344 (N_8344,N_7773,N_7646);
and U8345 (N_8345,N_7701,N_7543);
nor U8346 (N_8346,N_7923,N_7817);
nand U8347 (N_8347,N_7818,N_7793);
or U8348 (N_8348,N_7852,N_7750);
nand U8349 (N_8349,N_7774,N_7795);
or U8350 (N_8350,N_7690,N_7716);
nor U8351 (N_8351,N_7785,N_7730);
or U8352 (N_8352,N_7558,N_7691);
or U8353 (N_8353,N_7678,N_7824);
and U8354 (N_8354,N_7891,N_7552);
xnor U8355 (N_8355,N_7523,N_7581);
and U8356 (N_8356,N_7969,N_7686);
and U8357 (N_8357,N_7804,N_7718);
nand U8358 (N_8358,N_7744,N_7700);
and U8359 (N_8359,N_7743,N_7965);
and U8360 (N_8360,N_7661,N_7891);
nor U8361 (N_8361,N_7970,N_7506);
or U8362 (N_8362,N_7570,N_7832);
and U8363 (N_8363,N_7634,N_7864);
and U8364 (N_8364,N_7713,N_7968);
nand U8365 (N_8365,N_7757,N_7683);
nand U8366 (N_8366,N_7793,N_7872);
xnor U8367 (N_8367,N_7896,N_7956);
xnor U8368 (N_8368,N_7912,N_7609);
nand U8369 (N_8369,N_7731,N_7716);
nand U8370 (N_8370,N_7881,N_7707);
or U8371 (N_8371,N_7680,N_7507);
and U8372 (N_8372,N_7925,N_7622);
nand U8373 (N_8373,N_7696,N_7941);
and U8374 (N_8374,N_7962,N_7697);
or U8375 (N_8375,N_7993,N_7594);
and U8376 (N_8376,N_7841,N_7623);
and U8377 (N_8377,N_7746,N_7540);
nand U8378 (N_8378,N_7971,N_7799);
or U8379 (N_8379,N_7800,N_7836);
and U8380 (N_8380,N_7727,N_7921);
or U8381 (N_8381,N_7553,N_7810);
nor U8382 (N_8382,N_7908,N_7927);
or U8383 (N_8383,N_7710,N_7905);
and U8384 (N_8384,N_7878,N_7992);
and U8385 (N_8385,N_7867,N_7598);
and U8386 (N_8386,N_7637,N_7995);
and U8387 (N_8387,N_7604,N_7929);
or U8388 (N_8388,N_7940,N_7760);
or U8389 (N_8389,N_7798,N_7710);
and U8390 (N_8390,N_7805,N_7618);
and U8391 (N_8391,N_7784,N_7618);
nor U8392 (N_8392,N_7900,N_7652);
nand U8393 (N_8393,N_7610,N_7687);
and U8394 (N_8394,N_7697,N_7811);
nand U8395 (N_8395,N_7611,N_7596);
nor U8396 (N_8396,N_7939,N_7710);
and U8397 (N_8397,N_7902,N_7513);
nand U8398 (N_8398,N_7808,N_7604);
nor U8399 (N_8399,N_7896,N_7960);
or U8400 (N_8400,N_7936,N_7841);
nor U8401 (N_8401,N_7819,N_7551);
nor U8402 (N_8402,N_7994,N_7948);
nand U8403 (N_8403,N_7895,N_7846);
nor U8404 (N_8404,N_7848,N_7963);
or U8405 (N_8405,N_7500,N_7888);
or U8406 (N_8406,N_7902,N_7941);
nor U8407 (N_8407,N_7534,N_7854);
nor U8408 (N_8408,N_7660,N_7743);
nand U8409 (N_8409,N_7807,N_7983);
nand U8410 (N_8410,N_7525,N_7529);
nand U8411 (N_8411,N_7915,N_7893);
and U8412 (N_8412,N_7836,N_7549);
nor U8413 (N_8413,N_7985,N_7951);
nand U8414 (N_8414,N_7987,N_7685);
and U8415 (N_8415,N_7741,N_7907);
nor U8416 (N_8416,N_7561,N_7944);
nor U8417 (N_8417,N_7748,N_7768);
or U8418 (N_8418,N_7568,N_7674);
and U8419 (N_8419,N_7561,N_7993);
and U8420 (N_8420,N_7512,N_7733);
nand U8421 (N_8421,N_7849,N_7776);
nor U8422 (N_8422,N_7510,N_7929);
or U8423 (N_8423,N_7886,N_7698);
and U8424 (N_8424,N_7809,N_7856);
or U8425 (N_8425,N_7786,N_7721);
and U8426 (N_8426,N_7506,N_7686);
and U8427 (N_8427,N_7645,N_7641);
nand U8428 (N_8428,N_7987,N_7748);
nand U8429 (N_8429,N_7715,N_7586);
or U8430 (N_8430,N_7661,N_7719);
nand U8431 (N_8431,N_7753,N_7545);
and U8432 (N_8432,N_7820,N_7948);
or U8433 (N_8433,N_7688,N_7515);
and U8434 (N_8434,N_7906,N_7994);
and U8435 (N_8435,N_7904,N_7944);
or U8436 (N_8436,N_7622,N_7829);
or U8437 (N_8437,N_7587,N_7851);
or U8438 (N_8438,N_7852,N_7722);
or U8439 (N_8439,N_7868,N_7666);
nand U8440 (N_8440,N_7644,N_7963);
and U8441 (N_8441,N_7677,N_7742);
or U8442 (N_8442,N_7865,N_7586);
nand U8443 (N_8443,N_7841,N_7535);
nand U8444 (N_8444,N_7549,N_7523);
and U8445 (N_8445,N_7838,N_7547);
nand U8446 (N_8446,N_7687,N_7667);
nand U8447 (N_8447,N_7743,N_7719);
nand U8448 (N_8448,N_7612,N_7606);
or U8449 (N_8449,N_7906,N_7621);
nand U8450 (N_8450,N_7962,N_7615);
and U8451 (N_8451,N_7633,N_7995);
nor U8452 (N_8452,N_7565,N_7706);
nor U8453 (N_8453,N_7513,N_7807);
nand U8454 (N_8454,N_7938,N_7882);
nor U8455 (N_8455,N_7774,N_7893);
or U8456 (N_8456,N_7861,N_7812);
and U8457 (N_8457,N_7751,N_7938);
or U8458 (N_8458,N_7503,N_7827);
and U8459 (N_8459,N_7825,N_7636);
or U8460 (N_8460,N_7619,N_7704);
or U8461 (N_8461,N_7558,N_7828);
or U8462 (N_8462,N_7780,N_7940);
nor U8463 (N_8463,N_7561,N_7689);
nor U8464 (N_8464,N_7621,N_7655);
nor U8465 (N_8465,N_7787,N_7651);
and U8466 (N_8466,N_7827,N_7574);
nand U8467 (N_8467,N_7887,N_7576);
and U8468 (N_8468,N_7617,N_7995);
nor U8469 (N_8469,N_7989,N_7714);
or U8470 (N_8470,N_7503,N_7510);
and U8471 (N_8471,N_7798,N_7605);
nand U8472 (N_8472,N_7584,N_7571);
nor U8473 (N_8473,N_7694,N_7838);
nand U8474 (N_8474,N_7616,N_7806);
or U8475 (N_8475,N_7876,N_7577);
or U8476 (N_8476,N_7881,N_7704);
nand U8477 (N_8477,N_7540,N_7807);
nor U8478 (N_8478,N_7914,N_7813);
nor U8479 (N_8479,N_7811,N_7650);
nand U8480 (N_8480,N_7859,N_7535);
nor U8481 (N_8481,N_7642,N_7654);
nor U8482 (N_8482,N_7504,N_7991);
nand U8483 (N_8483,N_7596,N_7538);
nand U8484 (N_8484,N_7760,N_7769);
nor U8485 (N_8485,N_7936,N_7773);
nand U8486 (N_8486,N_7672,N_7751);
nor U8487 (N_8487,N_7644,N_7916);
nand U8488 (N_8488,N_7661,N_7853);
or U8489 (N_8489,N_7995,N_7568);
nand U8490 (N_8490,N_7837,N_7656);
nor U8491 (N_8491,N_7639,N_7994);
nand U8492 (N_8492,N_7960,N_7621);
and U8493 (N_8493,N_7776,N_7735);
and U8494 (N_8494,N_7620,N_7695);
nor U8495 (N_8495,N_7622,N_7835);
or U8496 (N_8496,N_7711,N_7610);
and U8497 (N_8497,N_7623,N_7765);
or U8498 (N_8498,N_7726,N_7929);
and U8499 (N_8499,N_7722,N_7627);
or U8500 (N_8500,N_8113,N_8014);
nor U8501 (N_8501,N_8194,N_8489);
nor U8502 (N_8502,N_8129,N_8171);
nand U8503 (N_8503,N_8230,N_8247);
and U8504 (N_8504,N_8432,N_8237);
nor U8505 (N_8505,N_8181,N_8413);
nor U8506 (N_8506,N_8033,N_8179);
nand U8507 (N_8507,N_8150,N_8177);
or U8508 (N_8508,N_8259,N_8254);
nand U8509 (N_8509,N_8483,N_8137);
and U8510 (N_8510,N_8332,N_8309);
nand U8511 (N_8511,N_8322,N_8243);
or U8512 (N_8512,N_8458,N_8303);
nand U8513 (N_8513,N_8477,N_8214);
nand U8514 (N_8514,N_8045,N_8337);
nor U8515 (N_8515,N_8233,N_8154);
and U8516 (N_8516,N_8258,N_8425);
and U8517 (N_8517,N_8152,N_8397);
and U8518 (N_8518,N_8128,N_8291);
nor U8519 (N_8519,N_8136,N_8357);
nor U8520 (N_8520,N_8111,N_8427);
or U8521 (N_8521,N_8069,N_8020);
and U8522 (N_8522,N_8249,N_8202);
and U8523 (N_8523,N_8324,N_8015);
and U8524 (N_8524,N_8294,N_8109);
or U8525 (N_8525,N_8000,N_8048);
or U8526 (N_8526,N_8132,N_8464);
nor U8527 (N_8527,N_8143,N_8384);
nand U8528 (N_8528,N_8223,N_8238);
nor U8529 (N_8529,N_8066,N_8327);
or U8530 (N_8530,N_8366,N_8484);
nand U8531 (N_8531,N_8036,N_8110);
or U8532 (N_8532,N_8054,N_8242);
or U8533 (N_8533,N_8326,N_8103);
nor U8534 (N_8534,N_8245,N_8052);
and U8535 (N_8535,N_8408,N_8006);
and U8536 (N_8536,N_8368,N_8467);
and U8537 (N_8537,N_8279,N_8151);
nor U8538 (N_8538,N_8466,N_8211);
nand U8539 (N_8539,N_8418,N_8399);
nand U8540 (N_8540,N_8076,N_8450);
nor U8541 (N_8541,N_8356,N_8341);
or U8542 (N_8542,N_8272,N_8264);
nand U8543 (N_8543,N_8117,N_8406);
nand U8544 (N_8544,N_8454,N_8301);
nand U8545 (N_8545,N_8371,N_8157);
or U8546 (N_8546,N_8459,N_8486);
or U8547 (N_8547,N_8082,N_8363);
nor U8548 (N_8548,N_8479,N_8044);
or U8549 (N_8549,N_8049,N_8472);
and U8550 (N_8550,N_8426,N_8126);
nand U8551 (N_8551,N_8490,N_8059);
nor U8552 (N_8552,N_8160,N_8283);
nand U8553 (N_8553,N_8053,N_8163);
nand U8554 (N_8554,N_8393,N_8091);
or U8555 (N_8555,N_8289,N_8423);
nor U8556 (N_8556,N_8265,N_8164);
and U8557 (N_8557,N_8481,N_8496);
nand U8558 (N_8558,N_8145,N_8431);
and U8559 (N_8559,N_8354,N_8468);
nor U8560 (N_8560,N_8175,N_8394);
or U8561 (N_8561,N_8170,N_8224);
nor U8562 (N_8562,N_8282,N_8402);
and U8563 (N_8563,N_8051,N_8446);
nand U8564 (N_8564,N_8353,N_8414);
and U8565 (N_8565,N_8046,N_8021);
xor U8566 (N_8566,N_8307,N_8293);
nand U8567 (N_8567,N_8209,N_8005);
and U8568 (N_8568,N_8096,N_8144);
nor U8569 (N_8569,N_8106,N_8186);
nand U8570 (N_8570,N_8205,N_8148);
and U8571 (N_8571,N_8198,N_8158);
nand U8572 (N_8572,N_8038,N_8365);
nor U8573 (N_8573,N_8424,N_8348);
nand U8574 (N_8574,N_8032,N_8093);
xor U8575 (N_8575,N_8379,N_8314);
nor U8576 (N_8576,N_8167,N_8183);
or U8577 (N_8577,N_8457,N_8491);
nor U8578 (N_8578,N_8041,N_8063);
nand U8579 (N_8579,N_8018,N_8057);
nor U8580 (N_8580,N_8391,N_8275);
and U8581 (N_8581,N_8473,N_8039);
or U8582 (N_8582,N_8452,N_8002);
and U8583 (N_8583,N_8058,N_8405);
nand U8584 (N_8584,N_8462,N_8292);
nand U8585 (N_8585,N_8390,N_8100);
and U8586 (N_8586,N_8409,N_8429);
or U8587 (N_8587,N_8221,N_8396);
and U8588 (N_8588,N_8085,N_8026);
or U8589 (N_8589,N_8274,N_8090);
nor U8590 (N_8590,N_8122,N_8206);
nor U8591 (N_8591,N_8193,N_8027);
and U8592 (N_8592,N_8493,N_8334);
or U8593 (N_8593,N_8299,N_8461);
nor U8594 (N_8594,N_8439,N_8192);
or U8595 (N_8595,N_8287,N_8138);
and U8596 (N_8596,N_8469,N_8300);
nand U8597 (N_8597,N_8433,N_8013);
nor U8598 (N_8598,N_8407,N_8311);
or U8599 (N_8599,N_8362,N_8412);
and U8600 (N_8600,N_8404,N_8448);
nand U8601 (N_8601,N_8342,N_8403);
and U8602 (N_8602,N_8313,N_8153);
nor U8603 (N_8603,N_8280,N_8270);
or U8604 (N_8604,N_8298,N_8174);
or U8605 (N_8605,N_8141,N_8127);
or U8606 (N_8606,N_8331,N_8430);
and U8607 (N_8607,N_8031,N_8182);
nand U8608 (N_8608,N_8343,N_8072);
nor U8609 (N_8609,N_8352,N_8361);
nor U8610 (N_8610,N_8217,N_8201);
or U8611 (N_8611,N_8135,N_8101);
or U8612 (N_8612,N_8008,N_8315);
and U8613 (N_8613,N_8378,N_8304);
nand U8614 (N_8614,N_8350,N_8239);
nor U8615 (N_8615,N_8386,N_8277);
and U8616 (N_8616,N_8207,N_8107);
and U8617 (N_8617,N_8329,N_8478);
or U8618 (N_8618,N_8095,N_8081);
nand U8619 (N_8619,N_8176,N_8438);
nor U8620 (N_8620,N_8050,N_8218);
and U8621 (N_8621,N_8121,N_8389);
nor U8622 (N_8622,N_8415,N_8024);
and U8623 (N_8623,N_8437,N_8411);
nor U8624 (N_8624,N_8112,N_8351);
nand U8625 (N_8625,N_8364,N_8263);
nor U8626 (N_8626,N_8480,N_8001);
or U8627 (N_8627,N_8323,N_8248);
and U8628 (N_8628,N_8215,N_8269);
nor U8629 (N_8629,N_8133,N_8213);
nor U8630 (N_8630,N_8199,N_8125);
nand U8631 (N_8631,N_8310,N_8382);
nor U8632 (N_8632,N_8234,N_8102);
nor U8633 (N_8633,N_8078,N_8312);
and U8634 (N_8634,N_8440,N_8184);
and U8635 (N_8635,N_8022,N_8492);
nor U8636 (N_8636,N_8344,N_8019);
nand U8637 (N_8637,N_8268,N_8004);
nor U8638 (N_8638,N_8320,N_8062);
xor U8639 (N_8639,N_8043,N_8498);
nor U8640 (N_8640,N_8098,N_8476);
xor U8641 (N_8641,N_8358,N_8318);
nand U8642 (N_8642,N_8104,N_8497);
or U8643 (N_8643,N_8338,N_8114);
and U8644 (N_8644,N_8253,N_8204);
nand U8645 (N_8645,N_8267,N_8040);
and U8646 (N_8646,N_8395,N_8017);
nand U8647 (N_8647,N_8488,N_8190);
nand U8648 (N_8648,N_8197,N_8271);
nand U8649 (N_8649,N_8453,N_8042);
nor U8650 (N_8650,N_8422,N_8097);
and U8651 (N_8651,N_8037,N_8385);
nor U8652 (N_8652,N_8079,N_8165);
or U8653 (N_8653,N_8149,N_8435);
nand U8654 (N_8654,N_8225,N_8372);
or U8655 (N_8655,N_8229,N_8346);
nand U8656 (N_8656,N_8187,N_8130);
nor U8657 (N_8657,N_8266,N_8220);
nand U8658 (N_8658,N_8392,N_8060);
nand U8659 (N_8659,N_8495,N_8281);
or U8660 (N_8660,N_8131,N_8231);
nor U8661 (N_8661,N_8118,N_8071);
or U8662 (N_8662,N_8116,N_8288);
nand U8663 (N_8663,N_8169,N_8055);
and U8664 (N_8664,N_8068,N_8035);
nand U8665 (N_8665,N_8200,N_8336);
or U8666 (N_8666,N_8123,N_8189);
nor U8667 (N_8667,N_8308,N_8428);
nor U8668 (N_8668,N_8380,N_8061);
or U8669 (N_8669,N_8124,N_8030);
and U8670 (N_8670,N_8067,N_8494);
and U8671 (N_8671,N_8359,N_8155);
nor U8672 (N_8672,N_8485,N_8369);
nor U8673 (N_8673,N_8256,N_8244);
nor U8674 (N_8674,N_8261,N_8142);
or U8675 (N_8675,N_8162,N_8222);
nor U8676 (N_8676,N_8023,N_8456);
and U8677 (N_8677,N_8442,N_8073);
and U8678 (N_8678,N_8262,N_8075);
nor U8679 (N_8679,N_8381,N_8108);
and U8680 (N_8680,N_8115,N_8306);
nand U8681 (N_8681,N_8195,N_8203);
nand U8682 (N_8682,N_8447,N_8325);
nor U8683 (N_8683,N_8376,N_8007);
or U8684 (N_8684,N_8420,N_8316);
nand U8685 (N_8685,N_8286,N_8011);
nor U8686 (N_8686,N_8296,N_8185);
or U8687 (N_8687,N_8094,N_8463);
nand U8688 (N_8688,N_8470,N_8375);
and U8689 (N_8689,N_8216,N_8499);
nand U8690 (N_8690,N_8319,N_8227);
and U8691 (N_8691,N_8047,N_8373);
nand U8692 (N_8692,N_8297,N_8250);
nor U8693 (N_8693,N_8347,N_8099);
or U8694 (N_8694,N_8482,N_8180);
nand U8695 (N_8695,N_8178,N_8172);
nor U8696 (N_8696,N_8370,N_8159);
or U8697 (N_8697,N_8134,N_8240);
nor U8698 (N_8698,N_8449,N_8173);
nor U8699 (N_8699,N_8360,N_8290);
and U8700 (N_8700,N_8252,N_8444);
and U8701 (N_8701,N_8228,N_8105);
nand U8702 (N_8702,N_8445,N_8339);
xor U8703 (N_8703,N_8305,N_8355);
or U8704 (N_8704,N_8410,N_8156);
or U8705 (N_8705,N_8421,N_8188);
nand U8706 (N_8706,N_8487,N_8475);
and U8707 (N_8707,N_8302,N_8070);
and U8708 (N_8708,N_8443,N_8398);
and U8709 (N_8709,N_8087,N_8285);
and U8710 (N_8710,N_8367,N_8092);
nor U8711 (N_8711,N_8084,N_8471);
nand U8712 (N_8712,N_8273,N_8328);
nor U8713 (N_8713,N_8003,N_8089);
nand U8714 (N_8714,N_8417,N_8196);
nor U8715 (N_8715,N_8139,N_8345);
nand U8716 (N_8716,N_8056,N_8257);
nor U8717 (N_8717,N_8147,N_8434);
nand U8718 (N_8718,N_8377,N_8333);
xnor U8719 (N_8719,N_8383,N_8009);
nor U8720 (N_8720,N_8065,N_8120);
nand U8721 (N_8721,N_8119,N_8086);
or U8722 (N_8722,N_8083,N_8064);
nand U8723 (N_8723,N_8168,N_8232);
nor U8724 (N_8724,N_8208,N_8235);
or U8725 (N_8725,N_8387,N_8321);
nand U8726 (N_8726,N_8340,N_8349);
nor U8727 (N_8727,N_8010,N_8400);
nand U8728 (N_8728,N_8025,N_8161);
or U8729 (N_8729,N_8335,N_8455);
and U8730 (N_8730,N_8401,N_8140);
nor U8731 (N_8731,N_8080,N_8441);
nand U8732 (N_8732,N_8416,N_8012);
and U8733 (N_8733,N_8088,N_8077);
nand U8734 (N_8734,N_8212,N_8251);
nor U8735 (N_8735,N_8278,N_8241);
nor U8736 (N_8736,N_8460,N_8074);
and U8737 (N_8737,N_8034,N_8317);
and U8738 (N_8738,N_8284,N_8451);
or U8739 (N_8739,N_8374,N_8028);
nand U8740 (N_8740,N_8295,N_8474);
and U8741 (N_8741,N_8388,N_8029);
or U8742 (N_8742,N_8219,N_8260);
nor U8743 (N_8743,N_8226,N_8146);
nor U8744 (N_8744,N_8166,N_8276);
nand U8745 (N_8745,N_8246,N_8436);
nor U8746 (N_8746,N_8465,N_8330);
nand U8747 (N_8747,N_8191,N_8236);
nor U8748 (N_8748,N_8419,N_8210);
nor U8749 (N_8749,N_8016,N_8255);
nor U8750 (N_8750,N_8332,N_8183);
and U8751 (N_8751,N_8155,N_8336);
nand U8752 (N_8752,N_8070,N_8003);
nand U8753 (N_8753,N_8478,N_8372);
and U8754 (N_8754,N_8280,N_8233);
or U8755 (N_8755,N_8218,N_8493);
nor U8756 (N_8756,N_8001,N_8320);
nor U8757 (N_8757,N_8052,N_8269);
and U8758 (N_8758,N_8300,N_8287);
nor U8759 (N_8759,N_8174,N_8197);
nor U8760 (N_8760,N_8385,N_8396);
and U8761 (N_8761,N_8290,N_8291);
nand U8762 (N_8762,N_8189,N_8057);
and U8763 (N_8763,N_8404,N_8280);
nand U8764 (N_8764,N_8195,N_8275);
nand U8765 (N_8765,N_8465,N_8441);
nor U8766 (N_8766,N_8390,N_8194);
nand U8767 (N_8767,N_8316,N_8124);
or U8768 (N_8768,N_8457,N_8186);
nand U8769 (N_8769,N_8343,N_8381);
and U8770 (N_8770,N_8319,N_8442);
nor U8771 (N_8771,N_8456,N_8301);
nand U8772 (N_8772,N_8186,N_8347);
or U8773 (N_8773,N_8086,N_8497);
or U8774 (N_8774,N_8151,N_8497);
or U8775 (N_8775,N_8386,N_8270);
nand U8776 (N_8776,N_8383,N_8230);
nand U8777 (N_8777,N_8261,N_8499);
and U8778 (N_8778,N_8353,N_8324);
and U8779 (N_8779,N_8121,N_8091);
nor U8780 (N_8780,N_8094,N_8071);
nor U8781 (N_8781,N_8241,N_8413);
nor U8782 (N_8782,N_8166,N_8263);
nand U8783 (N_8783,N_8368,N_8458);
and U8784 (N_8784,N_8418,N_8000);
and U8785 (N_8785,N_8067,N_8474);
or U8786 (N_8786,N_8203,N_8019);
nor U8787 (N_8787,N_8091,N_8303);
and U8788 (N_8788,N_8236,N_8255);
nor U8789 (N_8789,N_8031,N_8371);
and U8790 (N_8790,N_8298,N_8492);
nand U8791 (N_8791,N_8072,N_8188);
or U8792 (N_8792,N_8189,N_8200);
and U8793 (N_8793,N_8265,N_8010);
and U8794 (N_8794,N_8143,N_8106);
nor U8795 (N_8795,N_8043,N_8256);
and U8796 (N_8796,N_8162,N_8191);
nor U8797 (N_8797,N_8492,N_8341);
nor U8798 (N_8798,N_8452,N_8123);
nand U8799 (N_8799,N_8217,N_8275);
or U8800 (N_8800,N_8024,N_8459);
nand U8801 (N_8801,N_8238,N_8215);
and U8802 (N_8802,N_8185,N_8016);
and U8803 (N_8803,N_8006,N_8230);
nor U8804 (N_8804,N_8265,N_8319);
and U8805 (N_8805,N_8293,N_8125);
nand U8806 (N_8806,N_8048,N_8014);
nor U8807 (N_8807,N_8435,N_8410);
and U8808 (N_8808,N_8281,N_8440);
nand U8809 (N_8809,N_8314,N_8002);
nand U8810 (N_8810,N_8053,N_8250);
nand U8811 (N_8811,N_8359,N_8058);
nor U8812 (N_8812,N_8445,N_8304);
and U8813 (N_8813,N_8307,N_8406);
nor U8814 (N_8814,N_8029,N_8280);
or U8815 (N_8815,N_8018,N_8397);
and U8816 (N_8816,N_8349,N_8052);
nor U8817 (N_8817,N_8479,N_8305);
or U8818 (N_8818,N_8045,N_8000);
nand U8819 (N_8819,N_8066,N_8043);
nand U8820 (N_8820,N_8184,N_8106);
nor U8821 (N_8821,N_8099,N_8410);
nor U8822 (N_8822,N_8092,N_8151);
nand U8823 (N_8823,N_8302,N_8432);
nor U8824 (N_8824,N_8113,N_8355);
nor U8825 (N_8825,N_8176,N_8462);
or U8826 (N_8826,N_8144,N_8468);
and U8827 (N_8827,N_8033,N_8074);
or U8828 (N_8828,N_8106,N_8482);
or U8829 (N_8829,N_8456,N_8099);
nand U8830 (N_8830,N_8220,N_8346);
xnor U8831 (N_8831,N_8025,N_8457);
and U8832 (N_8832,N_8378,N_8279);
or U8833 (N_8833,N_8086,N_8212);
nand U8834 (N_8834,N_8101,N_8178);
xnor U8835 (N_8835,N_8342,N_8353);
and U8836 (N_8836,N_8376,N_8321);
and U8837 (N_8837,N_8123,N_8105);
nor U8838 (N_8838,N_8125,N_8453);
nor U8839 (N_8839,N_8001,N_8086);
and U8840 (N_8840,N_8268,N_8195);
nand U8841 (N_8841,N_8300,N_8284);
nor U8842 (N_8842,N_8173,N_8477);
or U8843 (N_8843,N_8102,N_8036);
or U8844 (N_8844,N_8356,N_8067);
or U8845 (N_8845,N_8488,N_8449);
or U8846 (N_8846,N_8387,N_8114);
nor U8847 (N_8847,N_8198,N_8343);
or U8848 (N_8848,N_8167,N_8182);
or U8849 (N_8849,N_8018,N_8094);
nor U8850 (N_8850,N_8085,N_8081);
nor U8851 (N_8851,N_8353,N_8212);
and U8852 (N_8852,N_8268,N_8207);
xnor U8853 (N_8853,N_8451,N_8132);
or U8854 (N_8854,N_8411,N_8247);
nor U8855 (N_8855,N_8122,N_8007);
or U8856 (N_8856,N_8064,N_8151);
nand U8857 (N_8857,N_8416,N_8065);
nor U8858 (N_8858,N_8337,N_8470);
nand U8859 (N_8859,N_8375,N_8432);
or U8860 (N_8860,N_8289,N_8220);
nor U8861 (N_8861,N_8444,N_8353);
nor U8862 (N_8862,N_8253,N_8035);
nand U8863 (N_8863,N_8063,N_8175);
or U8864 (N_8864,N_8224,N_8164);
nand U8865 (N_8865,N_8323,N_8157);
or U8866 (N_8866,N_8192,N_8482);
nor U8867 (N_8867,N_8053,N_8452);
nand U8868 (N_8868,N_8020,N_8229);
or U8869 (N_8869,N_8332,N_8499);
nand U8870 (N_8870,N_8135,N_8066);
and U8871 (N_8871,N_8331,N_8330);
or U8872 (N_8872,N_8199,N_8329);
and U8873 (N_8873,N_8311,N_8494);
nand U8874 (N_8874,N_8478,N_8474);
and U8875 (N_8875,N_8026,N_8037);
nand U8876 (N_8876,N_8188,N_8104);
and U8877 (N_8877,N_8392,N_8282);
and U8878 (N_8878,N_8227,N_8363);
and U8879 (N_8879,N_8268,N_8095);
nand U8880 (N_8880,N_8318,N_8403);
nor U8881 (N_8881,N_8170,N_8237);
or U8882 (N_8882,N_8394,N_8235);
or U8883 (N_8883,N_8050,N_8081);
and U8884 (N_8884,N_8004,N_8408);
or U8885 (N_8885,N_8028,N_8070);
or U8886 (N_8886,N_8260,N_8247);
and U8887 (N_8887,N_8017,N_8119);
nand U8888 (N_8888,N_8151,N_8464);
and U8889 (N_8889,N_8001,N_8293);
and U8890 (N_8890,N_8209,N_8196);
nor U8891 (N_8891,N_8087,N_8122);
and U8892 (N_8892,N_8163,N_8487);
and U8893 (N_8893,N_8429,N_8384);
nand U8894 (N_8894,N_8211,N_8490);
nor U8895 (N_8895,N_8210,N_8372);
nor U8896 (N_8896,N_8371,N_8163);
nand U8897 (N_8897,N_8247,N_8345);
nand U8898 (N_8898,N_8495,N_8286);
nor U8899 (N_8899,N_8269,N_8333);
or U8900 (N_8900,N_8104,N_8040);
and U8901 (N_8901,N_8007,N_8072);
or U8902 (N_8902,N_8417,N_8164);
nand U8903 (N_8903,N_8361,N_8323);
nor U8904 (N_8904,N_8019,N_8157);
nand U8905 (N_8905,N_8435,N_8469);
nand U8906 (N_8906,N_8488,N_8160);
nor U8907 (N_8907,N_8009,N_8492);
and U8908 (N_8908,N_8381,N_8207);
or U8909 (N_8909,N_8485,N_8226);
xor U8910 (N_8910,N_8218,N_8098);
or U8911 (N_8911,N_8282,N_8486);
nor U8912 (N_8912,N_8464,N_8456);
nand U8913 (N_8913,N_8112,N_8255);
nand U8914 (N_8914,N_8260,N_8379);
nand U8915 (N_8915,N_8156,N_8377);
and U8916 (N_8916,N_8319,N_8332);
or U8917 (N_8917,N_8388,N_8038);
and U8918 (N_8918,N_8331,N_8128);
xor U8919 (N_8919,N_8065,N_8312);
and U8920 (N_8920,N_8219,N_8396);
and U8921 (N_8921,N_8366,N_8487);
and U8922 (N_8922,N_8133,N_8163);
or U8923 (N_8923,N_8254,N_8317);
or U8924 (N_8924,N_8085,N_8166);
and U8925 (N_8925,N_8253,N_8181);
and U8926 (N_8926,N_8159,N_8219);
and U8927 (N_8927,N_8047,N_8098);
nor U8928 (N_8928,N_8266,N_8359);
or U8929 (N_8929,N_8062,N_8410);
xnor U8930 (N_8930,N_8248,N_8174);
nor U8931 (N_8931,N_8404,N_8164);
and U8932 (N_8932,N_8149,N_8396);
or U8933 (N_8933,N_8093,N_8036);
and U8934 (N_8934,N_8012,N_8315);
and U8935 (N_8935,N_8097,N_8098);
and U8936 (N_8936,N_8365,N_8207);
or U8937 (N_8937,N_8473,N_8170);
nor U8938 (N_8938,N_8047,N_8237);
nand U8939 (N_8939,N_8282,N_8121);
and U8940 (N_8940,N_8280,N_8269);
nand U8941 (N_8941,N_8444,N_8356);
or U8942 (N_8942,N_8304,N_8381);
nand U8943 (N_8943,N_8469,N_8106);
nand U8944 (N_8944,N_8453,N_8422);
nor U8945 (N_8945,N_8447,N_8222);
nand U8946 (N_8946,N_8072,N_8250);
or U8947 (N_8947,N_8052,N_8085);
nor U8948 (N_8948,N_8192,N_8046);
nand U8949 (N_8949,N_8158,N_8466);
nor U8950 (N_8950,N_8173,N_8483);
or U8951 (N_8951,N_8166,N_8187);
nand U8952 (N_8952,N_8463,N_8192);
or U8953 (N_8953,N_8359,N_8220);
nor U8954 (N_8954,N_8322,N_8048);
and U8955 (N_8955,N_8475,N_8398);
nand U8956 (N_8956,N_8455,N_8375);
nand U8957 (N_8957,N_8388,N_8242);
or U8958 (N_8958,N_8388,N_8238);
or U8959 (N_8959,N_8457,N_8423);
or U8960 (N_8960,N_8031,N_8158);
nand U8961 (N_8961,N_8180,N_8395);
or U8962 (N_8962,N_8159,N_8029);
or U8963 (N_8963,N_8417,N_8145);
nand U8964 (N_8964,N_8146,N_8305);
and U8965 (N_8965,N_8183,N_8084);
nor U8966 (N_8966,N_8148,N_8153);
or U8967 (N_8967,N_8043,N_8337);
or U8968 (N_8968,N_8032,N_8439);
nor U8969 (N_8969,N_8496,N_8484);
nor U8970 (N_8970,N_8100,N_8141);
nand U8971 (N_8971,N_8398,N_8147);
nand U8972 (N_8972,N_8139,N_8130);
and U8973 (N_8973,N_8160,N_8133);
or U8974 (N_8974,N_8457,N_8007);
nor U8975 (N_8975,N_8460,N_8106);
and U8976 (N_8976,N_8085,N_8269);
and U8977 (N_8977,N_8148,N_8070);
or U8978 (N_8978,N_8216,N_8196);
and U8979 (N_8979,N_8154,N_8130);
or U8980 (N_8980,N_8216,N_8065);
xnor U8981 (N_8981,N_8195,N_8415);
and U8982 (N_8982,N_8339,N_8401);
xor U8983 (N_8983,N_8066,N_8405);
and U8984 (N_8984,N_8085,N_8365);
nand U8985 (N_8985,N_8250,N_8459);
nand U8986 (N_8986,N_8150,N_8224);
nor U8987 (N_8987,N_8421,N_8237);
nand U8988 (N_8988,N_8169,N_8237);
nand U8989 (N_8989,N_8324,N_8300);
and U8990 (N_8990,N_8273,N_8205);
or U8991 (N_8991,N_8005,N_8177);
nand U8992 (N_8992,N_8347,N_8311);
and U8993 (N_8993,N_8122,N_8004);
nand U8994 (N_8994,N_8418,N_8330);
or U8995 (N_8995,N_8499,N_8498);
nand U8996 (N_8996,N_8116,N_8388);
and U8997 (N_8997,N_8116,N_8164);
and U8998 (N_8998,N_8115,N_8475);
or U8999 (N_8999,N_8487,N_8280);
or U9000 (N_9000,N_8674,N_8928);
and U9001 (N_9001,N_8629,N_8570);
nor U9002 (N_9002,N_8553,N_8528);
and U9003 (N_9003,N_8620,N_8686);
nand U9004 (N_9004,N_8860,N_8821);
nor U9005 (N_9005,N_8594,N_8929);
nand U9006 (N_9006,N_8654,N_8632);
or U9007 (N_9007,N_8783,N_8934);
and U9008 (N_9008,N_8905,N_8679);
or U9009 (N_9009,N_8542,N_8795);
or U9010 (N_9010,N_8742,N_8562);
xor U9011 (N_9011,N_8622,N_8628);
nand U9012 (N_9012,N_8663,N_8705);
and U9013 (N_9013,N_8541,N_8819);
or U9014 (N_9014,N_8978,N_8513);
or U9015 (N_9015,N_8973,N_8558);
nor U9016 (N_9016,N_8587,N_8900);
and U9017 (N_9017,N_8918,N_8915);
nor U9018 (N_9018,N_8621,N_8883);
nor U9019 (N_9019,N_8569,N_8511);
and U9020 (N_9020,N_8617,N_8745);
nor U9021 (N_9021,N_8760,N_8687);
and U9022 (N_9022,N_8965,N_8815);
nor U9023 (N_9023,N_8573,N_8908);
or U9024 (N_9024,N_8680,N_8703);
or U9025 (N_9025,N_8560,N_8980);
and U9026 (N_9026,N_8649,N_8563);
and U9027 (N_9027,N_8549,N_8986);
nor U9028 (N_9028,N_8575,N_8724);
or U9029 (N_9029,N_8976,N_8502);
and U9030 (N_9030,N_8579,N_8864);
and U9031 (N_9031,N_8597,N_8598);
nand U9032 (N_9032,N_8503,N_8737);
and U9033 (N_9033,N_8556,N_8999);
and U9034 (N_9034,N_8704,N_8892);
and U9035 (N_9035,N_8770,N_8518);
and U9036 (N_9036,N_8987,N_8989);
or U9037 (N_9037,N_8521,N_8675);
and U9038 (N_9038,N_8559,N_8804);
nor U9039 (N_9039,N_8958,N_8733);
or U9040 (N_9040,N_8938,N_8792);
nand U9041 (N_9041,N_8710,N_8802);
and U9042 (N_9042,N_8719,N_8896);
nand U9043 (N_9043,N_8699,N_8685);
nor U9044 (N_9044,N_8626,N_8669);
nand U9045 (N_9045,N_8778,N_8960);
or U9046 (N_9046,N_8913,N_8810);
nor U9047 (N_9047,N_8906,N_8727);
nor U9048 (N_9048,N_8867,N_8803);
or U9049 (N_9049,N_8645,N_8646);
or U9050 (N_9050,N_8641,N_8523);
nor U9051 (N_9051,N_8977,N_8774);
nand U9052 (N_9052,N_8666,N_8584);
and U9053 (N_9053,N_8624,N_8577);
or U9054 (N_9054,N_8949,N_8614);
nor U9055 (N_9055,N_8950,N_8941);
nor U9056 (N_9056,N_8970,N_8817);
or U9057 (N_9057,N_8608,N_8638);
or U9058 (N_9058,N_8557,N_8859);
and U9059 (N_9059,N_8758,N_8762);
nor U9060 (N_9060,N_8937,N_8532);
and U9061 (N_9061,N_8717,N_8512);
or U9062 (N_9062,N_8777,N_8902);
and U9063 (N_9063,N_8828,N_8767);
or U9064 (N_9064,N_8891,N_8789);
nor U9065 (N_9065,N_8870,N_8967);
and U9066 (N_9066,N_8855,N_8940);
nand U9067 (N_9067,N_8730,N_8567);
nand U9068 (N_9068,N_8882,N_8837);
nor U9069 (N_9069,N_8946,N_8725);
nor U9070 (N_9070,N_8874,N_8684);
and U9071 (N_9071,N_8786,N_8681);
and U9072 (N_9072,N_8580,N_8634);
and U9073 (N_9073,N_8526,N_8591);
or U9074 (N_9074,N_8827,N_8531);
nand U9075 (N_9075,N_8765,N_8854);
or U9076 (N_9076,N_8747,N_8939);
nor U9077 (N_9077,N_8947,N_8662);
nand U9078 (N_9078,N_8726,N_8933);
nand U9079 (N_9079,N_8793,N_8881);
and U9080 (N_9080,N_8930,N_8734);
and U9081 (N_9081,N_8613,N_8616);
and U9082 (N_9082,N_8981,N_8964);
nor U9083 (N_9083,N_8656,N_8856);
nand U9084 (N_9084,N_8923,N_8722);
nor U9085 (N_9085,N_8974,N_8651);
or U9086 (N_9086,N_8788,N_8691);
or U9087 (N_9087,N_8890,N_8944);
or U9088 (N_9088,N_8873,N_8971);
nand U9089 (N_9089,N_8612,N_8811);
nor U9090 (N_9090,N_8713,N_8901);
or U9091 (N_9091,N_8849,N_8667);
and U9092 (N_9092,N_8875,N_8748);
xor U9093 (N_9093,N_8903,N_8658);
nand U9094 (N_9094,N_8625,N_8838);
or U9095 (N_9095,N_8909,N_8990);
nor U9096 (N_9096,N_8853,N_8500);
nand U9097 (N_9097,N_8914,N_8566);
nor U9098 (N_9098,N_8768,N_8552);
nor U9099 (N_9099,N_8879,N_8682);
nor U9100 (N_9100,N_8657,N_8529);
and U9101 (N_9101,N_8863,N_8721);
nor U9102 (N_9102,N_8787,N_8785);
or U9103 (N_9103,N_8955,N_8547);
xnor U9104 (N_9104,N_8781,N_8865);
nor U9105 (N_9105,N_8732,N_8780);
and U9106 (N_9106,N_8919,N_8887);
and U9107 (N_9107,N_8602,N_8850);
nand U9108 (N_9108,N_8731,N_8991);
and U9109 (N_9109,N_8688,N_8535);
and U9110 (N_9110,N_8522,N_8678);
nand U9111 (N_9111,N_8800,N_8993);
and U9112 (N_9112,N_8581,N_8631);
or U9113 (N_9113,N_8872,N_8809);
and U9114 (N_9114,N_8953,N_8582);
nand U9115 (N_9115,N_8808,N_8884);
nor U9116 (N_9116,N_8668,N_8766);
and U9117 (N_9117,N_8673,N_8606);
nor U9118 (N_9118,N_8593,N_8520);
and U9119 (N_9119,N_8982,N_8985);
and U9120 (N_9120,N_8711,N_8832);
nor U9121 (N_9121,N_8655,N_8718);
and U9122 (N_9122,N_8861,N_8642);
or U9123 (N_9123,N_8565,N_8871);
nand U9124 (N_9124,N_8639,N_8611);
or U9125 (N_9125,N_8689,N_8755);
or U9126 (N_9126,N_8504,N_8508);
or U9127 (N_9127,N_8690,N_8515);
and U9128 (N_9128,N_8630,N_8885);
or U9129 (N_9129,N_8618,N_8866);
nand U9130 (N_9130,N_8844,N_8650);
nor U9131 (N_9131,N_8840,N_8664);
or U9132 (N_9132,N_8589,N_8633);
nor U9133 (N_9133,N_8596,N_8869);
or U9134 (N_9134,N_8701,N_8935);
and U9135 (N_9135,N_8665,N_8776);
and U9136 (N_9136,N_8551,N_8583);
nor U9137 (N_9137,N_8697,N_8898);
nand U9138 (N_9138,N_8886,N_8992);
nor U9139 (N_9139,N_8907,N_8979);
or U9140 (N_9140,N_8763,N_8961);
and U9141 (N_9141,N_8683,N_8839);
xor U9142 (N_9142,N_8835,N_8533);
nor U9143 (N_9143,N_8794,N_8706);
or U9144 (N_9144,N_8852,N_8525);
and U9145 (N_9145,N_8501,N_8897);
nor U9146 (N_9146,N_8670,N_8942);
nor U9147 (N_9147,N_8538,N_8696);
and U9148 (N_9148,N_8693,N_8752);
or U9149 (N_9149,N_8648,N_8814);
and U9150 (N_9150,N_8707,N_8539);
or U9151 (N_9151,N_8889,N_8769);
nand U9152 (N_9152,N_8695,N_8920);
or U9153 (N_9153,N_8833,N_8607);
nand U9154 (N_9154,N_8820,N_8729);
nand U9155 (N_9155,N_8997,N_8761);
or U9156 (N_9156,N_8895,N_8507);
and U9157 (N_9157,N_8983,N_8829);
or U9158 (N_9158,N_8652,N_8739);
nor U9159 (N_9159,N_8893,N_8824);
nand U9160 (N_9160,N_8806,N_8544);
nor U9161 (N_9161,N_8995,N_8694);
nand U9162 (N_9162,N_8534,N_8888);
or U9163 (N_9163,N_8599,N_8957);
nand U9164 (N_9164,N_8797,N_8975);
nor U9165 (N_9165,N_8555,N_8561);
and U9166 (N_9166,N_8925,N_8813);
or U9167 (N_9167,N_8831,N_8927);
and U9168 (N_9168,N_8543,N_8595);
nand U9169 (N_9169,N_8604,N_8917);
nand U9170 (N_9170,N_8659,N_8926);
and U9171 (N_9171,N_8848,N_8677);
and U9172 (N_9172,N_8799,N_8640);
nand U9173 (N_9173,N_8994,N_8728);
and U9174 (N_9174,N_8771,N_8753);
and U9175 (N_9175,N_8924,N_8572);
nor U9176 (N_9176,N_8880,N_8744);
or U9177 (N_9177,N_8635,N_8517);
or U9178 (N_9178,N_8530,N_8818);
nor U9179 (N_9179,N_8962,N_8796);
and U9180 (N_9180,N_8943,N_8894);
nor U9181 (N_9181,N_8904,N_8816);
and U9182 (N_9182,N_8972,N_8830);
or U9183 (N_9183,N_8931,N_8600);
and U9184 (N_9184,N_8603,N_8858);
nor U9185 (N_9185,N_8545,N_8911);
or U9186 (N_9186,N_8506,N_8609);
nor U9187 (N_9187,N_8812,N_8782);
nor U9188 (N_9188,N_8959,N_8956);
nand U9189 (N_9189,N_8822,N_8750);
nor U9190 (N_9190,N_8536,N_8951);
and U9191 (N_9191,N_8743,N_8672);
nor U9192 (N_9192,N_8825,N_8823);
and U9193 (N_9193,N_8524,N_8676);
and U9194 (N_9194,N_8736,N_8546);
nor U9195 (N_9195,N_8740,N_8554);
or U9196 (N_9196,N_8548,N_8636);
nor U9197 (N_9197,N_8968,N_8790);
nand U9198 (N_9198,N_8637,N_8945);
nand U9199 (N_9199,N_8592,N_8510);
and U9200 (N_9200,N_8574,N_8984);
or U9201 (N_9201,N_8836,N_8708);
and U9202 (N_9202,N_8916,N_8712);
nor U9203 (N_9203,N_8910,N_8537);
nor U9204 (N_9204,N_8988,N_8954);
and U9205 (N_9205,N_8805,N_8643);
and U9206 (N_9206,N_8723,N_8847);
nor U9207 (N_9207,N_8671,N_8702);
nor U9208 (N_9208,N_8784,N_8936);
nor U9209 (N_9209,N_8807,N_8615);
or U9210 (N_9210,N_8514,N_8627);
or U9211 (N_9211,N_8568,N_8516);
and U9212 (N_9212,N_8756,N_8899);
and U9213 (N_9213,N_8698,N_8772);
nand U9214 (N_9214,N_8741,N_8952);
and U9215 (N_9215,N_8834,N_8912);
nor U9216 (N_9216,N_8715,N_8714);
or U9217 (N_9217,N_8564,N_8826);
nor U9218 (N_9218,N_8749,N_8692);
and U9219 (N_9219,N_8751,N_8845);
nand U9220 (N_9220,N_8846,N_8966);
nor U9221 (N_9221,N_8505,N_8757);
nand U9222 (N_9222,N_8590,N_8843);
and U9223 (N_9223,N_8623,N_8709);
nand U9224 (N_9224,N_8996,N_8610);
nor U9225 (N_9225,N_8791,N_8653);
nand U9226 (N_9226,N_8588,N_8921);
and U9227 (N_9227,N_8775,N_8661);
nand U9228 (N_9228,N_8700,N_8932);
or U9229 (N_9229,N_8759,N_8754);
nand U9230 (N_9230,N_8842,N_8922);
nand U9231 (N_9231,N_8963,N_8660);
or U9232 (N_9232,N_8779,N_8868);
nand U9233 (N_9233,N_8841,N_8586);
nand U9234 (N_9234,N_8735,N_8605);
nor U9235 (N_9235,N_8877,N_8969);
nand U9236 (N_9236,N_8998,N_8716);
nand U9237 (N_9237,N_8876,N_8798);
and U9238 (N_9238,N_8509,N_8519);
and U9239 (N_9239,N_8540,N_8851);
and U9240 (N_9240,N_8578,N_8738);
nor U9241 (N_9241,N_8527,N_8720);
nand U9242 (N_9242,N_8571,N_8644);
nor U9243 (N_9243,N_8878,N_8948);
or U9244 (N_9244,N_8862,N_8647);
and U9245 (N_9245,N_8857,N_8619);
or U9246 (N_9246,N_8773,N_8801);
and U9247 (N_9247,N_8746,N_8550);
nor U9248 (N_9248,N_8764,N_8601);
nand U9249 (N_9249,N_8585,N_8576);
nor U9250 (N_9250,N_8629,N_8683);
nor U9251 (N_9251,N_8929,N_8604);
or U9252 (N_9252,N_8912,N_8697);
nand U9253 (N_9253,N_8681,N_8843);
nor U9254 (N_9254,N_8741,N_8923);
xnor U9255 (N_9255,N_8651,N_8674);
and U9256 (N_9256,N_8582,N_8813);
or U9257 (N_9257,N_8788,N_8931);
nand U9258 (N_9258,N_8624,N_8559);
nor U9259 (N_9259,N_8611,N_8997);
nor U9260 (N_9260,N_8504,N_8822);
or U9261 (N_9261,N_8936,N_8606);
or U9262 (N_9262,N_8629,N_8833);
and U9263 (N_9263,N_8825,N_8876);
and U9264 (N_9264,N_8727,N_8596);
or U9265 (N_9265,N_8750,N_8567);
and U9266 (N_9266,N_8904,N_8856);
nand U9267 (N_9267,N_8877,N_8648);
or U9268 (N_9268,N_8990,N_8626);
nand U9269 (N_9269,N_8779,N_8601);
or U9270 (N_9270,N_8990,N_8546);
nand U9271 (N_9271,N_8705,N_8563);
nor U9272 (N_9272,N_8745,N_8533);
or U9273 (N_9273,N_8651,N_8856);
and U9274 (N_9274,N_8872,N_8617);
xnor U9275 (N_9275,N_8994,N_8995);
xor U9276 (N_9276,N_8753,N_8756);
or U9277 (N_9277,N_8692,N_8883);
or U9278 (N_9278,N_8693,N_8699);
nor U9279 (N_9279,N_8978,N_8977);
and U9280 (N_9280,N_8616,N_8507);
nor U9281 (N_9281,N_8761,N_8921);
nor U9282 (N_9282,N_8972,N_8594);
nor U9283 (N_9283,N_8950,N_8827);
and U9284 (N_9284,N_8510,N_8570);
nand U9285 (N_9285,N_8655,N_8699);
and U9286 (N_9286,N_8517,N_8691);
nand U9287 (N_9287,N_8524,N_8842);
or U9288 (N_9288,N_8661,N_8977);
and U9289 (N_9289,N_8545,N_8717);
nand U9290 (N_9290,N_8794,N_8859);
and U9291 (N_9291,N_8622,N_8731);
nor U9292 (N_9292,N_8718,N_8712);
and U9293 (N_9293,N_8791,N_8614);
nand U9294 (N_9294,N_8728,N_8563);
or U9295 (N_9295,N_8604,N_8538);
and U9296 (N_9296,N_8765,N_8993);
nand U9297 (N_9297,N_8914,N_8538);
nand U9298 (N_9298,N_8758,N_8537);
nor U9299 (N_9299,N_8876,N_8950);
or U9300 (N_9300,N_8689,N_8945);
nand U9301 (N_9301,N_8577,N_8962);
or U9302 (N_9302,N_8636,N_8595);
nand U9303 (N_9303,N_8772,N_8749);
nor U9304 (N_9304,N_8740,N_8641);
or U9305 (N_9305,N_8520,N_8658);
and U9306 (N_9306,N_8554,N_8715);
nand U9307 (N_9307,N_8862,N_8939);
or U9308 (N_9308,N_8759,N_8888);
nor U9309 (N_9309,N_8792,N_8567);
nand U9310 (N_9310,N_8988,N_8967);
nand U9311 (N_9311,N_8909,N_8666);
nand U9312 (N_9312,N_8568,N_8639);
nand U9313 (N_9313,N_8811,N_8689);
and U9314 (N_9314,N_8924,N_8615);
and U9315 (N_9315,N_8982,N_8511);
nor U9316 (N_9316,N_8831,N_8863);
nand U9317 (N_9317,N_8887,N_8628);
or U9318 (N_9318,N_8873,N_8795);
nor U9319 (N_9319,N_8918,N_8670);
nand U9320 (N_9320,N_8858,N_8501);
nor U9321 (N_9321,N_8524,N_8615);
or U9322 (N_9322,N_8794,N_8690);
and U9323 (N_9323,N_8885,N_8619);
or U9324 (N_9324,N_8620,N_8683);
and U9325 (N_9325,N_8984,N_8641);
nor U9326 (N_9326,N_8768,N_8513);
nor U9327 (N_9327,N_8726,N_8518);
xnor U9328 (N_9328,N_8851,N_8759);
or U9329 (N_9329,N_8588,N_8510);
or U9330 (N_9330,N_8734,N_8951);
nand U9331 (N_9331,N_8727,N_8803);
or U9332 (N_9332,N_8644,N_8511);
nor U9333 (N_9333,N_8515,N_8791);
or U9334 (N_9334,N_8919,N_8685);
nand U9335 (N_9335,N_8576,N_8746);
and U9336 (N_9336,N_8806,N_8623);
nand U9337 (N_9337,N_8844,N_8596);
or U9338 (N_9338,N_8828,N_8755);
nor U9339 (N_9339,N_8989,N_8713);
nand U9340 (N_9340,N_8541,N_8922);
nand U9341 (N_9341,N_8607,N_8804);
nor U9342 (N_9342,N_8591,N_8593);
nand U9343 (N_9343,N_8664,N_8998);
and U9344 (N_9344,N_8704,N_8716);
nand U9345 (N_9345,N_8806,N_8561);
xor U9346 (N_9346,N_8773,N_8504);
or U9347 (N_9347,N_8738,N_8879);
nand U9348 (N_9348,N_8870,N_8894);
nor U9349 (N_9349,N_8520,N_8849);
and U9350 (N_9350,N_8587,N_8991);
and U9351 (N_9351,N_8840,N_8742);
nor U9352 (N_9352,N_8847,N_8925);
and U9353 (N_9353,N_8821,N_8514);
and U9354 (N_9354,N_8518,N_8941);
and U9355 (N_9355,N_8787,N_8769);
nor U9356 (N_9356,N_8776,N_8974);
and U9357 (N_9357,N_8958,N_8804);
nand U9358 (N_9358,N_8549,N_8811);
nand U9359 (N_9359,N_8951,N_8695);
and U9360 (N_9360,N_8633,N_8710);
and U9361 (N_9361,N_8948,N_8901);
nand U9362 (N_9362,N_8924,N_8825);
or U9363 (N_9363,N_8741,N_8616);
and U9364 (N_9364,N_8681,N_8769);
nand U9365 (N_9365,N_8716,N_8842);
nor U9366 (N_9366,N_8680,N_8903);
or U9367 (N_9367,N_8706,N_8721);
and U9368 (N_9368,N_8774,N_8918);
or U9369 (N_9369,N_8997,N_8820);
nand U9370 (N_9370,N_8796,N_8512);
or U9371 (N_9371,N_8982,N_8820);
and U9372 (N_9372,N_8662,N_8981);
or U9373 (N_9373,N_8957,N_8933);
and U9374 (N_9374,N_8875,N_8599);
and U9375 (N_9375,N_8972,N_8918);
and U9376 (N_9376,N_8549,N_8673);
nor U9377 (N_9377,N_8536,N_8960);
nand U9378 (N_9378,N_8506,N_8780);
and U9379 (N_9379,N_8608,N_8947);
and U9380 (N_9380,N_8509,N_8762);
nand U9381 (N_9381,N_8819,N_8700);
and U9382 (N_9382,N_8791,N_8953);
or U9383 (N_9383,N_8519,N_8540);
and U9384 (N_9384,N_8559,N_8825);
or U9385 (N_9385,N_8951,N_8941);
or U9386 (N_9386,N_8725,N_8945);
or U9387 (N_9387,N_8872,N_8749);
and U9388 (N_9388,N_8649,N_8797);
and U9389 (N_9389,N_8558,N_8863);
and U9390 (N_9390,N_8693,N_8846);
nand U9391 (N_9391,N_8922,N_8591);
and U9392 (N_9392,N_8939,N_8954);
nand U9393 (N_9393,N_8954,N_8744);
nand U9394 (N_9394,N_8836,N_8717);
and U9395 (N_9395,N_8963,N_8745);
and U9396 (N_9396,N_8644,N_8528);
and U9397 (N_9397,N_8731,N_8523);
nand U9398 (N_9398,N_8792,N_8610);
nor U9399 (N_9399,N_8820,N_8935);
nor U9400 (N_9400,N_8625,N_8589);
and U9401 (N_9401,N_8608,N_8992);
or U9402 (N_9402,N_8778,N_8614);
nor U9403 (N_9403,N_8763,N_8832);
or U9404 (N_9404,N_8837,N_8986);
and U9405 (N_9405,N_8530,N_8591);
nand U9406 (N_9406,N_8719,N_8999);
nand U9407 (N_9407,N_8536,N_8993);
or U9408 (N_9408,N_8824,N_8921);
nor U9409 (N_9409,N_8510,N_8797);
or U9410 (N_9410,N_8763,N_8632);
nor U9411 (N_9411,N_8718,N_8792);
or U9412 (N_9412,N_8813,N_8946);
or U9413 (N_9413,N_8669,N_8869);
and U9414 (N_9414,N_8810,N_8886);
nand U9415 (N_9415,N_8788,N_8958);
or U9416 (N_9416,N_8936,N_8594);
nor U9417 (N_9417,N_8634,N_8952);
or U9418 (N_9418,N_8831,N_8610);
and U9419 (N_9419,N_8722,N_8845);
nor U9420 (N_9420,N_8835,N_8715);
nand U9421 (N_9421,N_8682,N_8785);
or U9422 (N_9422,N_8824,N_8539);
or U9423 (N_9423,N_8902,N_8726);
nand U9424 (N_9424,N_8710,N_8532);
xor U9425 (N_9425,N_8756,N_8530);
nand U9426 (N_9426,N_8546,N_8611);
xor U9427 (N_9427,N_8853,N_8803);
nor U9428 (N_9428,N_8752,N_8827);
or U9429 (N_9429,N_8685,N_8848);
or U9430 (N_9430,N_8919,N_8869);
and U9431 (N_9431,N_8989,N_8801);
and U9432 (N_9432,N_8751,N_8754);
nor U9433 (N_9433,N_8971,N_8560);
nor U9434 (N_9434,N_8575,N_8760);
nor U9435 (N_9435,N_8799,N_8606);
nor U9436 (N_9436,N_8956,N_8718);
or U9437 (N_9437,N_8994,N_8744);
or U9438 (N_9438,N_8837,N_8617);
nor U9439 (N_9439,N_8822,N_8644);
and U9440 (N_9440,N_8772,N_8542);
xnor U9441 (N_9441,N_8963,N_8844);
nor U9442 (N_9442,N_8840,N_8997);
and U9443 (N_9443,N_8723,N_8681);
nand U9444 (N_9444,N_8833,N_8625);
nor U9445 (N_9445,N_8988,N_8892);
or U9446 (N_9446,N_8806,N_8660);
nand U9447 (N_9447,N_8942,N_8931);
or U9448 (N_9448,N_8816,N_8538);
nor U9449 (N_9449,N_8608,N_8581);
and U9450 (N_9450,N_8837,N_8917);
and U9451 (N_9451,N_8834,N_8793);
and U9452 (N_9452,N_8732,N_8508);
nor U9453 (N_9453,N_8566,N_8963);
nor U9454 (N_9454,N_8864,N_8921);
and U9455 (N_9455,N_8693,N_8972);
nor U9456 (N_9456,N_8883,N_8586);
nor U9457 (N_9457,N_8927,N_8693);
nand U9458 (N_9458,N_8823,N_8798);
nor U9459 (N_9459,N_8821,N_8837);
nand U9460 (N_9460,N_8901,N_8547);
and U9461 (N_9461,N_8822,N_8500);
or U9462 (N_9462,N_8811,N_8974);
nand U9463 (N_9463,N_8739,N_8576);
nand U9464 (N_9464,N_8674,N_8976);
or U9465 (N_9465,N_8641,N_8552);
nand U9466 (N_9466,N_8603,N_8924);
and U9467 (N_9467,N_8892,N_8523);
nor U9468 (N_9468,N_8929,N_8978);
nor U9469 (N_9469,N_8887,N_8975);
or U9470 (N_9470,N_8993,N_8532);
and U9471 (N_9471,N_8806,N_8612);
or U9472 (N_9472,N_8952,N_8770);
nor U9473 (N_9473,N_8661,N_8958);
or U9474 (N_9474,N_8950,N_8772);
and U9475 (N_9475,N_8536,N_8548);
or U9476 (N_9476,N_8635,N_8634);
or U9477 (N_9477,N_8903,N_8824);
nor U9478 (N_9478,N_8974,N_8828);
nor U9479 (N_9479,N_8821,N_8710);
and U9480 (N_9480,N_8644,N_8840);
and U9481 (N_9481,N_8723,N_8617);
nand U9482 (N_9482,N_8921,N_8573);
and U9483 (N_9483,N_8786,N_8877);
nor U9484 (N_9484,N_8664,N_8945);
nand U9485 (N_9485,N_8876,N_8989);
nand U9486 (N_9486,N_8555,N_8863);
or U9487 (N_9487,N_8785,N_8729);
and U9488 (N_9488,N_8578,N_8950);
or U9489 (N_9489,N_8790,N_8791);
nand U9490 (N_9490,N_8553,N_8629);
or U9491 (N_9491,N_8743,N_8816);
nand U9492 (N_9492,N_8714,N_8652);
nor U9493 (N_9493,N_8867,N_8598);
nor U9494 (N_9494,N_8691,N_8674);
nand U9495 (N_9495,N_8749,N_8625);
nand U9496 (N_9496,N_8594,N_8607);
nor U9497 (N_9497,N_8893,N_8670);
nand U9498 (N_9498,N_8763,N_8859);
or U9499 (N_9499,N_8615,N_8691);
and U9500 (N_9500,N_9230,N_9273);
or U9501 (N_9501,N_9205,N_9247);
or U9502 (N_9502,N_9019,N_9180);
nand U9503 (N_9503,N_9049,N_9415);
or U9504 (N_9504,N_9025,N_9393);
nor U9505 (N_9505,N_9052,N_9171);
or U9506 (N_9506,N_9182,N_9351);
nor U9507 (N_9507,N_9360,N_9407);
nor U9508 (N_9508,N_9280,N_9163);
and U9509 (N_9509,N_9367,N_9057);
and U9510 (N_9510,N_9154,N_9045);
nor U9511 (N_9511,N_9353,N_9161);
and U9512 (N_9512,N_9439,N_9391);
nor U9513 (N_9513,N_9189,N_9333);
and U9514 (N_9514,N_9251,N_9417);
and U9515 (N_9515,N_9158,N_9093);
nor U9516 (N_9516,N_9235,N_9159);
and U9517 (N_9517,N_9341,N_9226);
and U9518 (N_9518,N_9347,N_9033);
nand U9519 (N_9519,N_9398,N_9186);
or U9520 (N_9520,N_9084,N_9430);
xor U9521 (N_9521,N_9438,N_9232);
or U9522 (N_9522,N_9266,N_9244);
nand U9523 (N_9523,N_9043,N_9324);
or U9524 (N_9524,N_9326,N_9485);
or U9525 (N_9525,N_9488,N_9175);
or U9526 (N_9526,N_9318,N_9047);
nor U9527 (N_9527,N_9078,N_9113);
nand U9528 (N_9528,N_9443,N_9060);
and U9529 (N_9529,N_9050,N_9123);
and U9530 (N_9530,N_9164,N_9011);
nor U9531 (N_9531,N_9480,N_9356);
and U9532 (N_9532,N_9167,N_9269);
nand U9533 (N_9533,N_9003,N_9392);
and U9534 (N_9534,N_9172,N_9343);
and U9535 (N_9535,N_9075,N_9453);
and U9536 (N_9536,N_9127,N_9272);
nand U9537 (N_9537,N_9174,N_9424);
nand U9538 (N_9538,N_9065,N_9059);
or U9539 (N_9539,N_9320,N_9370);
or U9540 (N_9540,N_9109,N_9130);
nor U9541 (N_9541,N_9100,N_9498);
nand U9542 (N_9542,N_9128,N_9355);
or U9543 (N_9543,N_9384,N_9215);
or U9544 (N_9544,N_9067,N_9069);
nand U9545 (N_9545,N_9371,N_9148);
and U9546 (N_9546,N_9440,N_9144);
and U9547 (N_9547,N_9181,N_9039);
nor U9548 (N_9548,N_9002,N_9283);
or U9549 (N_9549,N_9395,N_9041);
nand U9550 (N_9550,N_9170,N_9124);
or U9551 (N_9551,N_9221,N_9137);
and U9552 (N_9552,N_9151,N_9292);
nor U9553 (N_9553,N_9289,N_9310);
nand U9554 (N_9554,N_9029,N_9473);
or U9555 (N_9555,N_9467,N_9420);
nor U9556 (N_9556,N_9012,N_9284);
nand U9557 (N_9557,N_9135,N_9162);
nand U9558 (N_9558,N_9404,N_9132);
nor U9559 (N_9559,N_9241,N_9242);
and U9560 (N_9560,N_9243,N_9297);
and U9561 (N_9561,N_9452,N_9111);
nand U9562 (N_9562,N_9032,N_9224);
or U9563 (N_9563,N_9455,N_9362);
nand U9564 (N_9564,N_9133,N_9074);
nor U9565 (N_9565,N_9462,N_9028);
and U9566 (N_9566,N_9116,N_9330);
and U9567 (N_9567,N_9304,N_9448);
and U9568 (N_9568,N_9290,N_9293);
or U9569 (N_9569,N_9139,N_9416);
nand U9570 (N_9570,N_9449,N_9193);
nand U9571 (N_9571,N_9344,N_9478);
or U9572 (N_9572,N_9007,N_9489);
nor U9573 (N_9573,N_9345,N_9044);
and U9574 (N_9574,N_9436,N_9017);
nand U9575 (N_9575,N_9357,N_9222);
nor U9576 (N_9576,N_9267,N_9021);
or U9577 (N_9577,N_9434,N_9218);
or U9578 (N_9578,N_9220,N_9239);
and U9579 (N_9579,N_9444,N_9006);
and U9580 (N_9580,N_9466,N_9114);
nor U9581 (N_9581,N_9143,N_9302);
or U9582 (N_9582,N_9339,N_9046);
nand U9583 (N_9583,N_9223,N_9454);
and U9584 (N_9584,N_9432,N_9372);
and U9585 (N_9585,N_9316,N_9185);
or U9586 (N_9586,N_9248,N_9168);
and U9587 (N_9587,N_9319,N_9173);
nand U9588 (N_9588,N_9388,N_9368);
nand U9589 (N_9589,N_9446,N_9340);
nand U9590 (N_9590,N_9202,N_9134);
or U9591 (N_9591,N_9274,N_9147);
nand U9592 (N_9592,N_9457,N_9107);
or U9593 (N_9593,N_9387,N_9053);
and U9594 (N_9594,N_9321,N_9279);
or U9595 (N_9595,N_9497,N_9258);
and U9596 (N_9596,N_9275,N_9020);
nand U9597 (N_9597,N_9098,N_9265);
or U9598 (N_9598,N_9421,N_9257);
nor U9599 (N_9599,N_9091,N_9027);
nor U9600 (N_9600,N_9264,N_9016);
nor U9601 (N_9601,N_9090,N_9451);
or U9602 (N_9602,N_9270,N_9286);
and U9603 (N_9603,N_9382,N_9227);
and U9604 (N_9604,N_9104,N_9165);
nand U9605 (N_9605,N_9194,N_9217);
nand U9606 (N_9606,N_9307,N_9179);
xnor U9607 (N_9607,N_9299,N_9335);
nand U9608 (N_9608,N_9034,N_9153);
and U9609 (N_9609,N_9350,N_9401);
nor U9610 (N_9610,N_9071,N_9008);
and U9611 (N_9611,N_9411,N_9484);
and U9612 (N_9612,N_9155,N_9169);
nand U9613 (N_9613,N_9058,N_9447);
nand U9614 (N_9614,N_9219,N_9140);
nor U9615 (N_9615,N_9066,N_9429);
and U9616 (N_9616,N_9410,N_9460);
or U9617 (N_9617,N_9073,N_9237);
and U9618 (N_9618,N_9191,N_9352);
or U9619 (N_9619,N_9196,N_9380);
nand U9620 (N_9620,N_9346,N_9470);
or U9621 (N_9621,N_9229,N_9081);
nor U9622 (N_9622,N_9233,N_9492);
or U9623 (N_9623,N_9495,N_9254);
nand U9624 (N_9624,N_9358,N_9231);
nor U9625 (N_9625,N_9082,N_9472);
and U9626 (N_9626,N_9051,N_9010);
or U9627 (N_9627,N_9465,N_9197);
and U9628 (N_9628,N_9262,N_9328);
nand U9629 (N_9629,N_9225,N_9402);
and U9630 (N_9630,N_9418,N_9048);
and U9631 (N_9631,N_9409,N_9150);
nor U9632 (N_9632,N_9322,N_9184);
nand U9633 (N_9633,N_9037,N_9342);
nand U9634 (N_9634,N_9327,N_9177);
nand U9635 (N_9635,N_9192,N_9394);
or U9636 (N_9636,N_9178,N_9129);
or U9637 (N_9637,N_9119,N_9157);
nor U9638 (N_9638,N_9209,N_9332);
nor U9639 (N_9639,N_9433,N_9099);
or U9640 (N_9640,N_9373,N_9379);
and U9641 (N_9641,N_9195,N_9260);
nand U9642 (N_9642,N_9490,N_9022);
and U9643 (N_9643,N_9072,N_9240);
nor U9644 (N_9644,N_9435,N_9259);
nor U9645 (N_9645,N_9001,N_9276);
or U9646 (N_9646,N_9256,N_9375);
or U9647 (N_9647,N_9306,N_9131);
and U9648 (N_9648,N_9252,N_9413);
or U9649 (N_9649,N_9487,N_9101);
and U9650 (N_9650,N_9285,N_9277);
nand U9651 (N_9651,N_9312,N_9294);
or U9652 (N_9652,N_9145,N_9095);
and U9653 (N_9653,N_9477,N_9329);
nand U9654 (N_9654,N_9390,N_9303);
and U9655 (N_9655,N_9009,N_9425);
or U9656 (N_9656,N_9325,N_9088);
and U9657 (N_9657,N_9077,N_9102);
nand U9658 (N_9658,N_9288,N_9281);
nor U9659 (N_9659,N_9450,N_9376);
xnor U9660 (N_9660,N_9491,N_9026);
nor U9661 (N_9661,N_9141,N_9210);
nor U9662 (N_9662,N_9397,N_9377);
nand U9663 (N_9663,N_9408,N_9403);
or U9664 (N_9664,N_9471,N_9004);
nand U9665 (N_9665,N_9361,N_9199);
xnor U9666 (N_9666,N_9054,N_9152);
nand U9667 (N_9667,N_9092,N_9085);
and U9668 (N_9668,N_9461,N_9468);
nor U9669 (N_9669,N_9015,N_9494);
and U9670 (N_9670,N_9187,N_9108);
nand U9671 (N_9671,N_9469,N_9486);
and U9672 (N_9672,N_9476,N_9300);
or U9673 (N_9673,N_9278,N_9366);
nor U9674 (N_9674,N_9369,N_9348);
nand U9675 (N_9675,N_9213,N_9349);
and U9676 (N_9676,N_9309,N_9126);
nand U9677 (N_9677,N_9305,N_9061);
nor U9678 (N_9678,N_9263,N_9030);
or U9679 (N_9679,N_9354,N_9176);
and U9680 (N_9680,N_9253,N_9499);
and U9681 (N_9681,N_9323,N_9018);
nor U9682 (N_9682,N_9214,N_9055);
nand U9683 (N_9683,N_9121,N_9087);
nor U9684 (N_9684,N_9314,N_9334);
nand U9685 (N_9685,N_9261,N_9138);
nand U9686 (N_9686,N_9207,N_9422);
and U9687 (N_9687,N_9198,N_9249);
nor U9688 (N_9688,N_9374,N_9105);
or U9689 (N_9689,N_9493,N_9456);
or U9690 (N_9690,N_9208,N_9441);
or U9691 (N_9691,N_9080,N_9201);
nand U9692 (N_9692,N_9110,N_9359);
or U9693 (N_9693,N_9200,N_9136);
or U9694 (N_9694,N_9381,N_9118);
and U9695 (N_9695,N_9188,N_9203);
nand U9696 (N_9696,N_9282,N_9024);
nand U9697 (N_9697,N_9031,N_9216);
and U9698 (N_9698,N_9399,N_9496);
nor U9699 (N_9699,N_9298,N_9386);
nor U9700 (N_9700,N_9062,N_9042);
nand U9701 (N_9701,N_9183,N_9313);
nand U9702 (N_9702,N_9234,N_9423);
nand U9703 (N_9703,N_9437,N_9035);
and U9704 (N_9704,N_9000,N_9086);
and U9705 (N_9705,N_9315,N_9094);
nor U9706 (N_9706,N_9474,N_9295);
or U9707 (N_9707,N_9149,N_9122);
nor U9708 (N_9708,N_9228,N_9255);
nand U9709 (N_9709,N_9412,N_9317);
nand U9710 (N_9710,N_9442,N_9079);
nand U9711 (N_9711,N_9364,N_9023);
and U9712 (N_9712,N_9096,N_9389);
nor U9713 (N_9713,N_9056,N_9166);
nor U9714 (N_9714,N_9287,N_9481);
and U9715 (N_9715,N_9070,N_9125);
nand U9716 (N_9716,N_9414,N_9482);
and U9717 (N_9717,N_9336,N_9427);
or U9718 (N_9718,N_9268,N_9005);
nand U9719 (N_9719,N_9445,N_9311);
nor U9720 (N_9720,N_9458,N_9246);
or U9721 (N_9721,N_9014,N_9396);
nand U9722 (N_9722,N_9156,N_9112);
nor U9723 (N_9723,N_9308,N_9426);
and U9724 (N_9724,N_9038,N_9365);
and U9725 (N_9725,N_9463,N_9245);
or U9726 (N_9726,N_9206,N_9160);
and U9727 (N_9727,N_9337,N_9190);
or U9728 (N_9728,N_9097,N_9238);
and U9729 (N_9729,N_9405,N_9475);
nor U9730 (N_9730,N_9378,N_9013);
or U9731 (N_9731,N_9271,N_9338);
xnor U9732 (N_9732,N_9431,N_9236);
nor U9733 (N_9733,N_9428,N_9211);
nand U9734 (N_9734,N_9400,N_9301);
nor U9735 (N_9735,N_9106,N_9406);
nor U9736 (N_9736,N_9383,N_9068);
nand U9737 (N_9737,N_9250,N_9212);
or U9738 (N_9738,N_9296,N_9083);
or U9739 (N_9739,N_9204,N_9464);
or U9740 (N_9740,N_9459,N_9063);
and U9741 (N_9741,N_9103,N_9291);
nor U9742 (N_9742,N_9142,N_9117);
and U9743 (N_9743,N_9331,N_9115);
nand U9744 (N_9744,N_9363,N_9120);
or U9745 (N_9745,N_9483,N_9089);
nor U9746 (N_9746,N_9064,N_9076);
or U9747 (N_9747,N_9385,N_9146);
and U9748 (N_9748,N_9479,N_9040);
or U9749 (N_9749,N_9036,N_9419);
and U9750 (N_9750,N_9364,N_9067);
and U9751 (N_9751,N_9018,N_9363);
nor U9752 (N_9752,N_9247,N_9476);
and U9753 (N_9753,N_9138,N_9334);
nand U9754 (N_9754,N_9364,N_9485);
or U9755 (N_9755,N_9435,N_9357);
nor U9756 (N_9756,N_9450,N_9344);
nor U9757 (N_9757,N_9463,N_9004);
or U9758 (N_9758,N_9013,N_9027);
nor U9759 (N_9759,N_9276,N_9305);
nor U9760 (N_9760,N_9074,N_9173);
or U9761 (N_9761,N_9450,N_9145);
or U9762 (N_9762,N_9255,N_9424);
and U9763 (N_9763,N_9386,N_9194);
or U9764 (N_9764,N_9315,N_9001);
nor U9765 (N_9765,N_9184,N_9409);
nand U9766 (N_9766,N_9406,N_9342);
or U9767 (N_9767,N_9052,N_9436);
nor U9768 (N_9768,N_9203,N_9194);
and U9769 (N_9769,N_9194,N_9157);
nor U9770 (N_9770,N_9421,N_9102);
nor U9771 (N_9771,N_9117,N_9357);
nor U9772 (N_9772,N_9371,N_9395);
nand U9773 (N_9773,N_9437,N_9090);
and U9774 (N_9774,N_9353,N_9425);
nor U9775 (N_9775,N_9395,N_9111);
nor U9776 (N_9776,N_9423,N_9412);
or U9777 (N_9777,N_9118,N_9037);
and U9778 (N_9778,N_9459,N_9447);
nand U9779 (N_9779,N_9150,N_9077);
nor U9780 (N_9780,N_9006,N_9483);
or U9781 (N_9781,N_9150,N_9405);
and U9782 (N_9782,N_9447,N_9256);
and U9783 (N_9783,N_9343,N_9463);
nor U9784 (N_9784,N_9076,N_9444);
or U9785 (N_9785,N_9208,N_9046);
or U9786 (N_9786,N_9365,N_9352);
nor U9787 (N_9787,N_9219,N_9114);
nand U9788 (N_9788,N_9220,N_9123);
and U9789 (N_9789,N_9048,N_9327);
nor U9790 (N_9790,N_9377,N_9140);
nor U9791 (N_9791,N_9088,N_9475);
and U9792 (N_9792,N_9110,N_9438);
nor U9793 (N_9793,N_9367,N_9420);
nand U9794 (N_9794,N_9314,N_9263);
nand U9795 (N_9795,N_9342,N_9444);
and U9796 (N_9796,N_9067,N_9350);
or U9797 (N_9797,N_9084,N_9340);
or U9798 (N_9798,N_9454,N_9175);
and U9799 (N_9799,N_9215,N_9266);
and U9800 (N_9800,N_9415,N_9167);
and U9801 (N_9801,N_9307,N_9064);
nand U9802 (N_9802,N_9409,N_9486);
and U9803 (N_9803,N_9202,N_9055);
or U9804 (N_9804,N_9103,N_9041);
and U9805 (N_9805,N_9062,N_9099);
nor U9806 (N_9806,N_9439,N_9041);
nand U9807 (N_9807,N_9105,N_9447);
and U9808 (N_9808,N_9389,N_9080);
nor U9809 (N_9809,N_9468,N_9038);
and U9810 (N_9810,N_9418,N_9388);
or U9811 (N_9811,N_9120,N_9059);
and U9812 (N_9812,N_9236,N_9301);
or U9813 (N_9813,N_9139,N_9254);
nor U9814 (N_9814,N_9464,N_9411);
or U9815 (N_9815,N_9146,N_9105);
or U9816 (N_9816,N_9448,N_9296);
and U9817 (N_9817,N_9009,N_9374);
and U9818 (N_9818,N_9230,N_9309);
nand U9819 (N_9819,N_9384,N_9181);
or U9820 (N_9820,N_9319,N_9408);
and U9821 (N_9821,N_9006,N_9311);
nand U9822 (N_9822,N_9125,N_9327);
nand U9823 (N_9823,N_9283,N_9190);
and U9824 (N_9824,N_9213,N_9401);
nand U9825 (N_9825,N_9228,N_9020);
or U9826 (N_9826,N_9183,N_9200);
or U9827 (N_9827,N_9497,N_9066);
and U9828 (N_9828,N_9195,N_9106);
nor U9829 (N_9829,N_9429,N_9041);
nor U9830 (N_9830,N_9176,N_9005);
nor U9831 (N_9831,N_9390,N_9359);
or U9832 (N_9832,N_9080,N_9428);
and U9833 (N_9833,N_9455,N_9317);
and U9834 (N_9834,N_9224,N_9483);
nand U9835 (N_9835,N_9410,N_9030);
nor U9836 (N_9836,N_9117,N_9444);
nor U9837 (N_9837,N_9039,N_9469);
nor U9838 (N_9838,N_9217,N_9325);
or U9839 (N_9839,N_9308,N_9009);
and U9840 (N_9840,N_9166,N_9276);
and U9841 (N_9841,N_9373,N_9017);
nand U9842 (N_9842,N_9358,N_9044);
and U9843 (N_9843,N_9024,N_9366);
nor U9844 (N_9844,N_9300,N_9162);
nor U9845 (N_9845,N_9170,N_9142);
or U9846 (N_9846,N_9040,N_9489);
nand U9847 (N_9847,N_9295,N_9062);
nand U9848 (N_9848,N_9077,N_9125);
nand U9849 (N_9849,N_9313,N_9332);
nand U9850 (N_9850,N_9468,N_9432);
and U9851 (N_9851,N_9017,N_9346);
and U9852 (N_9852,N_9276,N_9383);
or U9853 (N_9853,N_9187,N_9060);
nor U9854 (N_9854,N_9200,N_9167);
nand U9855 (N_9855,N_9355,N_9003);
and U9856 (N_9856,N_9395,N_9198);
and U9857 (N_9857,N_9296,N_9082);
nand U9858 (N_9858,N_9270,N_9387);
or U9859 (N_9859,N_9489,N_9363);
nor U9860 (N_9860,N_9212,N_9157);
or U9861 (N_9861,N_9105,N_9351);
and U9862 (N_9862,N_9024,N_9276);
nand U9863 (N_9863,N_9397,N_9167);
nand U9864 (N_9864,N_9453,N_9137);
or U9865 (N_9865,N_9014,N_9071);
nor U9866 (N_9866,N_9246,N_9247);
nand U9867 (N_9867,N_9230,N_9320);
or U9868 (N_9868,N_9400,N_9190);
or U9869 (N_9869,N_9264,N_9335);
nor U9870 (N_9870,N_9071,N_9073);
or U9871 (N_9871,N_9275,N_9048);
or U9872 (N_9872,N_9348,N_9211);
nand U9873 (N_9873,N_9214,N_9474);
nor U9874 (N_9874,N_9075,N_9489);
nand U9875 (N_9875,N_9375,N_9498);
nor U9876 (N_9876,N_9404,N_9498);
or U9877 (N_9877,N_9087,N_9173);
and U9878 (N_9878,N_9494,N_9392);
or U9879 (N_9879,N_9165,N_9009);
and U9880 (N_9880,N_9078,N_9253);
nand U9881 (N_9881,N_9124,N_9111);
nand U9882 (N_9882,N_9391,N_9195);
nor U9883 (N_9883,N_9089,N_9454);
or U9884 (N_9884,N_9404,N_9030);
or U9885 (N_9885,N_9428,N_9478);
nand U9886 (N_9886,N_9476,N_9036);
nand U9887 (N_9887,N_9179,N_9452);
and U9888 (N_9888,N_9485,N_9369);
nand U9889 (N_9889,N_9168,N_9297);
or U9890 (N_9890,N_9170,N_9345);
or U9891 (N_9891,N_9384,N_9457);
nand U9892 (N_9892,N_9074,N_9171);
or U9893 (N_9893,N_9074,N_9226);
nor U9894 (N_9894,N_9045,N_9373);
nand U9895 (N_9895,N_9279,N_9133);
xnor U9896 (N_9896,N_9272,N_9047);
nor U9897 (N_9897,N_9100,N_9411);
nor U9898 (N_9898,N_9060,N_9377);
nor U9899 (N_9899,N_9348,N_9074);
or U9900 (N_9900,N_9043,N_9322);
nor U9901 (N_9901,N_9232,N_9045);
or U9902 (N_9902,N_9008,N_9247);
and U9903 (N_9903,N_9088,N_9419);
and U9904 (N_9904,N_9203,N_9138);
or U9905 (N_9905,N_9116,N_9356);
nor U9906 (N_9906,N_9193,N_9233);
nor U9907 (N_9907,N_9004,N_9289);
nor U9908 (N_9908,N_9020,N_9365);
or U9909 (N_9909,N_9046,N_9190);
and U9910 (N_9910,N_9273,N_9177);
and U9911 (N_9911,N_9477,N_9272);
nor U9912 (N_9912,N_9250,N_9445);
or U9913 (N_9913,N_9355,N_9452);
nand U9914 (N_9914,N_9325,N_9494);
nand U9915 (N_9915,N_9427,N_9211);
or U9916 (N_9916,N_9304,N_9007);
or U9917 (N_9917,N_9283,N_9264);
nand U9918 (N_9918,N_9395,N_9203);
or U9919 (N_9919,N_9450,N_9392);
or U9920 (N_9920,N_9325,N_9049);
nor U9921 (N_9921,N_9353,N_9064);
nand U9922 (N_9922,N_9161,N_9035);
nand U9923 (N_9923,N_9452,N_9392);
and U9924 (N_9924,N_9156,N_9439);
and U9925 (N_9925,N_9254,N_9417);
and U9926 (N_9926,N_9180,N_9249);
and U9927 (N_9927,N_9446,N_9479);
nand U9928 (N_9928,N_9338,N_9492);
or U9929 (N_9929,N_9242,N_9427);
and U9930 (N_9930,N_9364,N_9276);
xor U9931 (N_9931,N_9277,N_9263);
or U9932 (N_9932,N_9322,N_9063);
nand U9933 (N_9933,N_9418,N_9177);
nor U9934 (N_9934,N_9167,N_9222);
nor U9935 (N_9935,N_9072,N_9225);
or U9936 (N_9936,N_9228,N_9036);
nand U9937 (N_9937,N_9045,N_9091);
or U9938 (N_9938,N_9457,N_9495);
and U9939 (N_9939,N_9226,N_9264);
and U9940 (N_9940,N_9087,N_9198);
nor U9941 (N_9941,N_9325,N_9393);
nand U9942 (N_9942,N_9325,N_9055);
nor U9943 (N_9943,N_9225,N_9021);
or U9944 (N_9944,N_9031,N_9470);
and U9945 (N_9945,N_9230,N_9308);
and U9946 (N_9946,N_9256,N_9206);
or U9947 (N_9947,N_9114,N_9178);
nand U9948 (N_9948,N_9058,N_9219);
or U9949 (N_9949,N_9123,N_9083);
or U9950 (N_9950,N_9097,N_9193);
nand U9951 (N_9951,N_9240,N_9306);
nand U9952 (N_9952,N_9261,N_9304);
nand U9953 (N_9953,N_9189,N_9030);
nand U9954 (N_9954,N_9132,N_9326);
or U9955 (N_9955,N_9184,N_9062);
or U9956 (N_9956,N_9157,N_9374);
nor U9957 (N_9957,N_9379,N_9233);
nor U9958 (N_9958,N_9471,N_9258);
and U9959 (N_9959,N_9039,N_9336);
or U9960 (N_9960,N_9189,N_9064);
nor U9961 (N_9961,N_9020,N_9114);
or U9962 (N_9962,N_9141,N_9096);
and U9963 (N_9963,N_9019,N_9350);
and U9964 (N_9964,N_9017,N_9354);
and U9965 (N_9965,N_9453,N_9345);
or U9966 (N_9966,N_9187,N_9464);
and U9967 (N_9967,N_9376,N_9250);
or U9968 (N_9968,N_9399,N_9270);
and U9969 (N_9969,N_9142,N_9334);
or U9970 (N_9970,N_9230,N_9316);
nor U9971 (N_9971,N_9048,N_9161);
nor U9972 (N_9972,N_9140,N_9110);
nand U9973 (N_9973,N_9057,N_9175);
or U9974 (N_9974,N_9408,N_9012);
nand U9975 (N_9975,N_9227,N_9466);
nor U9976 (N_9976,N_9099,N_9176);
and U9977 (N_9977,N_9326,N_9056);
or U9978 (N_9978,N_9093,N_9047);
and U9979 (N_9979,N_9352,N_9175);
nor U9980 (N_9980,N_9457,N_9240);
nor U9981 (N_9981,N_9346,N_9080);
and U9982 (N_9982,N_9330,N_9233);
nand U9983 (N_9983,N_9182,N_9109);
nand U9984 (N_9984,N_9026,N_9406);
and U9985 (N_9985,N_9243,N_9007);
and U9986 (N_9986,N_9132,N_9069);
and U9987 (N_9987,N_9466,N_9464);
nand U9988 (N_9988,N_9090,N_9297);
and U9989 (N_9989,N_9262,N_9229);
nand U9990 (N_9990,N_9296,N_9316);
nor U9991 (N_9991,N_9447,N_9168);
or U9992 (N_9992,N_9257,N_9299);
or U9993 (N_9993,N_9135,N_9335);
nor U9994 (N_9994,N_9129,N_9061);
nor U9995 (N_9995,N_9002,N_9028);
nor U9996 (N_9996,N_9075,N_9189);
nor U9997 (N_9997,N_9041,N_9384);
or U9998 (N_9998,N_9211,N_9053);
nand U9999 (N_9999,N_9251,N_9230);
or U10000 (N_10000,N_9745,N_9827);
xnor U10001 (N_10001,N_9604,N_9977);
or U10002 (N_10002,N_9616,N_9509);
nor U10003 (N_10003,N_9626,N_9612);
and U10004 (N_10004,N_9722,N_9605);
or U10005 (N_10005,N_9966,N_9572);
nand U10006 (N_10006,N_9559,N_9922);
nor U10007 (N_10007,N_9746,N_9799);
and U10008 (N_10008,N_9561,N_9554);
nand U10009 (N_10009,N_9601,N_9757);
nand U10010 (N_10010,N_9598,N_9810);
nand U10011 (N_10011,N_9792,N_9649);
or U10012 (N_10012,N_9564,N_9990);
and U10013 (N_10013,N_9943,N_9664);
and U10014 (N_10014,N_9873,N_9883);
or U10015 (N_10015,N_9514,N_9923);
and U10016 (N_10016,N_9661,N_9540);
nor U10017 (N_10017,N_9737,N_9621);
nor U10018 (N_10018,N_9866,N_9813);
and U10019 (N_10019,N_9894,N_9547);
nand U10020 (N_10020,N_9533,N_9761);
and U10021 (N_10021,N_9603,N_9837);
or U10022 (N_10022,N_9955,N_9963);
and U10023 (N_10023,N_9788,N_9997);
or U10024 (N_10024,N_9762,N_9687);
and U10025 (N_10025,N_9717,N_9599);
nand U10026 (N_10026,N_9726,N_9899);
nand U10027 (N_10027,N_9893,N_9663);
or U10028 (N_10028,N_9812,N_9742);
nor U10029 (N_10029,N_9962,N_9868);
nor U10030 (N_10030,N_9732,N_9608);
and U10031 (N_10031,N_9948,N_9713);
nand U10032 (N_10032,N_9674,N_9625);
or U10033 (N_10033,N_9929,N_9536);
nand U10034 (N_10034,N_9716,N_9517);
xor U10035 (N_10035,N_9576,N_9889);
and U10036 (N_10036,N_9821,N_9987);
nor U10037 (N_10037,N_9627,N_9522);
or U10038 (N_10038,N_9708,N_9692);
nand U10039 (N_10039,N_9550,N_9901);
and U10040 (N_10040,N_9871,N_9706);
nand U10041 (N_10041,N_9678,N_9506);
nand U10042 (N_10042,N_9876,N_9562);
and U10043 (N_10043,N_9971,N_9710);
nor U10044 (N_10044,N_9635,N_9681);
nor U10045 (N_10045,N_9507,N_9823);
or U10046 (N_10046,N_9973,N_9778);
nand U10047 (N_10047,N_9927,N_9529);
or U10048 (N_10048,N_9566,N_9758);
nand U10049 (N_10049,N_9691,N_9911);
nor U10050 (N_10050,N_9647,N_9921);
or U10051 (N_10051,N_9685,N_9748);
or U10052 (N_10052,N_9844,N_9865);
nor U10053 (N_10053,N_9546,N_9610);
nor U10054 (N_10054,N_9659,N_9904);
or U10055 (N_10055,N_9944,N_9641);
or U10056 (N_10056,N_9730,N_9819);
or U10057 (N_10057,N_9895,N_9860);
and U10058 (N_10058,N_9829,N_9556);
and U10059 (N_10059,N_9578,N_9539);
or U10060 (N_10060,N_9887,N_9545);
and U10061 (N_10061,N_9916,N_9993);
or U10062 (N_10062,N_9982,N_9655);
or U10063 (N_10063,N_9833,N_9518);
or U10064 (N_10064,N_9932,N_9931);
or U10065 (N_10065,N_9835,N_9841);
and U10066 (N_10066,N_9751,N_9567);
or U10067 (N_10067,N_9679,N_9801);
nand U10068 (N_10068,N_9636,N_9814);
nand U10069 (N_10069,N_9670,N_9861);
or U10070 (N_10070,N_9704,N_9777);
and U10071 (N_10071,N_9872,N_9953);
or U10072 (N_10072,N_9632,N_9839);
nand U10073 (N_10073,N_9620,N_9854);
nand U10074 (N_10074,N_9631,N_9880);
and U10075 (N_10075,N_9719,N_9733);
nor U10076 (N_10076,N_9569,N_9597);
or U10077 (N_10077,N_9945,N_9563);
nand U10078 (N_10078,N_9975,N_9830);
nor U10079 (N_10079,N_9979,N_9648);
nand U10080 (N_10080,N_9644,N_9832);
nor U10081 (N_10081,N_9782,N_9634);
nor U10082 (N_10082,N_9571,N_9581);
and U10083 (N_10083,N_9637,N_9867);
or U10084 (N_10084,N_9729,N_9989);
and U10085 (N_10085,N_9771,N_9542);
or U10086 (N_10086,N_9537,N_9940);
nor U10087 (N_10087,N_9698,N_9557);
or U10088 (N_10088,N_9912,N_9828);
and U10089 (N_10089,N_9891,N_9847);
nand U10090 (N_10090,N_9501,N_9803);
nor U10091 (N_10091,N_9902,N_9958);
nand U10092 (N_10092,N_9642,N_9906);
or U10093 (N_10093,N_9858,N_9853);
and U10094 (N_10094,N_9967,N_9974);
or U10095 (N_10095,N_9702,N_9573);
nand U10096 (N_10096,N_9628,N_9548);
or U10097 (N_10097,N_9511,N_9503);
nor U10098 (N_10098,N_9756,N_9864);
nand U10099 (N_10099,N_9721,N_9960);
nand U10100 (N_10100,N_9505,N_9718);
nor U10101 (N_10101,N_9534,N_9677);
or U10102 (N_10102,N_9918,N_9580);
nand U10103 (N_10103,N_9947,N_9836);
nand U10104 (N_10104,N_9525,N_9798);
nor U10105 (N_10105,N_9747,N_9957);
nand U10106 (N_10106,N_9683,N_9660);
nand U10107 (N_10107,N_9749,N_9651);
nand U10108 (N_10108,N_9807,N_9970);
or U10109 (N_10109,N_9707,N_9753);
or U10110 (N_10110,N_9743,N_9521);
or U10111 (N_10111,N_9976,N_9884);
or U10112 (N_10112,N_9523,N_9988);
or U10113 (N_10113,N_9934,N_9985);
and U10114 (N_10114,N_9815,N_9686);
or U10115 (N_10115,N_9903,N_9705);
nor U10116 (N_10116,N_9696,N_9577);
or U10117 (N_10117,N_9723,N_9790);
and U10118 (N_10118,N_9825,N_9935);
or U10119 (N_10119,N_9796,N_9654);
or U10120 (N_10120,N_9532,N_9838);
nand U10121 (N_10121,N_9639,N_9936);
and U10122 (N_10122,N_9555,N_9986);
nor U10123 (N_10123,N_9671,N_9711);
or U10124 (N_10124,N_9951,N_9898);
or U10125 (N_10125,N_9606,N_9519);
nor U10126 (N_10126,N_9874,N_9956);
or U10127 (N_10127,N_9794,N_9862);
and U10128 (N_10128,N_9926,N_9857);
xnor U10129 (N_10129,N_9781,N_9583);
or U10130 (N_10130,N_9870,N_9816);
nand U10131 (N_10131,N_9972,N_9991);
or U10132 (N_10132,N_9907,N_9849);
xor U10133 (N_10133,N_9512,N_9731);
or U10134 (N_10134,N_9712,N_9544);
or U10135 (N_10135,N_9842,N_9910);
and U10136 (N_10136,N_9558,N_9789);
or U10137 (N_10137,N_9863,N_9767);
or U10138 (N_10138,N_9755,N_9652);
nand U10139 (N_10139,N_9669,N_9797);
nor U10140 (N_10140,N_9508,N_9524);
and U10141 (N_10141,N_9896,N_9667);
nor U10142 (N_10142,N_9996,N_9834);
nand U10143 (N_10143,N_9530,N_9741);
and U10144 (N_10144,N_9510,N_9773);
nand U10145 (N_10145,N_9551,N_9930);
nor U10146 (N_10146,N_9793,N_9805);
or U10147 (N_10147,N_9658,N_9787);
nor U10148 (N_10148,N_9579,N_9630);
or U10149 (N_10149,N_9920,N_9676);
and U10150 (N_10150,N_9694,N_9994);
nand U10151 (N_10151,N_9763,N_9806);
nand U10152 (N_10152,N_9504,N_9969);
and U10153 (N_10153,N_9968,N_9850);
nand U10154 (N_10154,N_9811,N_9984);
nand U10155 (N_10155,N_9882,N_9774);
nand U10156 (N_10156,N_9543,N_9851);
nor U10157 (N_10157,N_9688,N_9961);
or U10158 (N_10158,N_9924,N_9769);
and U10159 (N_10159,N_9584,N_9843);
nand U10160 (N_10160,N_9818,N_9900);
nand U10161 (N_10161,N_9750,N_9856);
nand U10162 (N_10162,N_9728,N_9570);
and U10163 (N_10163,N_9701,N_9673);
nand U10164 (N_10164,N_9808,N_9699);
or U10165 (N_10165,N_9888,N_9999);
nand U10166 (N_10166,N_9846,N_9527);
and U10167 (N_10167,N_9560,N_9638);
or U10168 (N_10168,N_9954,N_9766);
nor U10169 (N_10169,N_9734,N_9675);
and U10170 (N_10170,N_9709,N_9689);
xnor U10171 (N_10171,N_9802,N_9528);
nor U10172 (N_10172,N_9822,N_9852);
nand U10173 (N_10173,N_9582,N_9549);
nor U10174 (N_10174,N_9591,N_9520);
nand U10175 (N_10175,N_9869,N_9587);
nand U10176 (N_10176,N_9568,N_9879);
or U10177 (N_10177,N_9650,N_9859);
and U10178 (N_10178,N_9877,N_9592);
or U10179 (N_10179,N_9772,N_9727);
and U10180 (N_10180,N_9715,N_9680);
and U10181 (N_10181,N_9740,N_9791);
nor U10182 (N_10182,N_9693,N_9624);
and U10183 (N_10183,N_9919,N_9725);
and U10184 (N_10184,N_9905,N_9765);
nand U10185 (N_10185,N_9593,N_9928);
nor U10186 (N_10186,N_9502,N_9939);
nor U10187 (N_10187,N_9995,N_9878);
nand U10188 (N_10188,N_9697,N_9917);
or U10189 (N_10189,N_9662,N_9611);
and U10190 (N_10190,N_9531,N_9602);
nor U10191 (N_10191,N_9764,N_9786);
or U10192 (N_10192,N_9909,N_9574);
nand U10193 (N_10193,N_9890,N_9633);
nor U10194 (N_10194,N_9950,N_9700);
or U10195 (N_10195,N_9752,N_9607);
or U10196 (N_10196,N_9538,N_9586);
or U10197 (N_10197,N_9892,N_9594);
or U10198 (N_10198,N_9617,N_9565);
or U10199 (N_10199,N_9824,N_9619);
nand U10200 (N_10200,N_9779,N_9665);
nand U10201 (N_10201,N_9914,N_9959);
nand U10202 (N_10202,N_9622,N_9585);
and U10203 (N_10203,N_9998,N_9744);
nor U10204 (N_10204,N_9513,N_9809);
nand U10205 (N_10205,N_9684,N_9595);
and U10206 (N_10206,N_9515,N_9609);
nand U10207 (N_10207,N_9596,N_9775);
and U10208 (N_10208,N_9964,N_9615);
or U10209 (N_10209,N_9776,N_9657);
or U10210 (N_10210,N_9885,N_9938);
nand U10211 (N_10211,N_9553,N_9760);
xor U10212 (N_10212,N_9915,N_9820);
nand U10213 (N_10213,N_9981,N_9720);
nor U10214 (N_10214,N_9881,N_9780);
and U10215 (N_10215,N_9600,N_9937);
nor U10216 (N_10216,N_9736,N_9575);
and U10217 (N_10217,N_9614,N_9933);
and U10218 (N_10218,N_9941,N_9897);
nand U10219 (N_10219,N_9643,N_9653);
or U10220 (N_10220,N_9783,N_9589);
or U10221 (N_10221,N_9980,N_9516);
or U10222 (N_10222,N_9908,N_9754);
nor U10223 (N_10223,N_9724,N_9785);
nor U10224 (N_10224,N_9739,N_9848);
nand U10225 (N_10225,N_9768,N_9672);
and U10226 (N_10226,N_9875,N_9831);
nand U10227 (N_10227,N_9666,N_9656);
nor U10228 (N_10228,N_9668,N_9552);
or U10229 (N_10229,N_9784,N_9500);
or U10230 (N_10230,N_9759,N_9526);
or U10231 (N_10231,N_9804,N_9618);
and U10232 (N_10232,N_9913,N_9640);
and U10233 (N_10233,N_9646,N_9682);
nand U10234 (N_10234,N_9590,N_9703);
and U10235 (N_10235,N_9965,N_9795);
or U10236 (N_10236,N_9840,N_9629);
and U10237 (N_10237,N_9826,N_9942);
nand U10238 (N_10238,N_9535,N_9695);
and U10239 (N_10239,N_9541,N_9978);
or U10240 (N_10240,N_9690,N_9817);
nand U10241 (N_10241,N_9952,N_9735);
and U10242 (N_10242,N_9845,N_9645);
and U10243 (N_10243,N_9925,N_9738);
or U10244 (N_10244,N_9992,N_9714);
nor U10245 (N_10245,N_9855,N_9949);
nand U10246 (N_10246,N_9770,N_9946);
nand U10247 (N_10247,N_9983,N_9613);
and U10248 (N_10248,N_9886,N_9800);
and U10249 (N_10249,N_9588,N_9623);
nor U10250 (N_10250,N_9932,N_9811);
nor U10251 (N_10251,N_9642,N_9793);
nor U10252 (N_10252,N_9665,N_9960);
nand U10253 (N_10253,N_9654,N_9908);
and U10254 (N_10254,N_9849,N_9785);
nand U10255 (N_10255,N_9555,N_9715);
or U10256 (N_10256,N_9628,N_9958);
or U10257 (N_10257,N_9501,N_9888);
and U10258 (N_10258,N_9846,N_9588);
or U10259 (N_10259,N_9636,N_9623);
or U10260 (N_10260,N_9873,N_9668);
nor U10261 (N_10261,N_9967,N_9573);
or U10262 (N_10262,N_9991,N_9595);
nor U10263 (N_10263,N_9760,N_9919);
and U10264 (N_10264,N_9942,N_9792);
nor U10265 (N_10265,N_9604,N_9989);
nor U10266 (N_10266,N_9697,N_9920);
nand U10267 (N_10267,N_9557,N_9782);
nor U10268 (N_10268,N_9974,N_9992);
nor U10269 (N_10269,N_9580,N_9995);
or U10270 (N_10270,N_9586,N_9557);
or U10271 (N_10271,N_9735,N_9846);
nand U10272 (N_10272,N_9813,N_9581);
or U10273 (N_10273,N_9520,N_9928);
and U10274 (N_10274,N_9845,N_9953);
and U10275 (N_10275,N_9504,N_9532);
nand U10276 (N_10276,N_9661,N_9785);
nor U10277 (N_10277,N_9735,N_9518);
nand U10278 (N_10278,N_9938,N_9738);
and U10279 (N_10279,N_9671,N_9682);
and U10280 (N_10280,N_9995,N_9514);
and U10281 (N_10281,N_9695,N_9943);
or U10282 (N_10282,N_9896,N_9788);
and U10283 (N_10283,N_9586,N_9671);
nor U10284 (N_10284,N_9800,N_9761);
or U10285 (N_10285,N_9534,N_9978);
or U10286 (N_10286,N_9881,N_9674);
xor U10287 (N_10287,N_9751,N_9587);
nand U10288 (N_10288,N_9501,N_9630);
nand U10289 (N_10289,N_9628,N_9755);
nand U10290 (N_10290,N_9807,N_9983);
nor U10291 (N_10291,N_9562,N_9750);
and U10292 (N_10292,N_9823,N_9877);
and U10293 (N_10293,N_9829,N_9783);
or U10294 (N_10294,N_9947,N_9882);
or U10295 (N_10295,N_9918,N_9556);
nor U10296 (N_10296,N_9742,N_9919);
nand U10297 (N_10297,N_9923,N_9636);
and U10298 (N_10298,N_9869,N_9854);
or U10299 (N_10299,N_9759,N_9613);
nor U10300 (N_10300,N_9764,N_9717);
nand U10301 (N_10301,N_9759,N_9789);
nor U10302 (N_10302,N_9748,N_9594);
nor U10303 (N_10303,N_9961,N_9759);
nand U10304 (N_10304,N_9706,N_9949);
nand U10305 (N_10305,N_9873,N_9816);
or U10306 (N_10306,N_9684,N_9785);
and U10307 (N_10307,N_9677,N_9714);
and U10308 (N_10308,N_9507,N_9850);
and U10309 (N_10309,N_9729,N_9550);
nor U10310 (N_10310,N_9939,N_9832);
and U10311 (N_10311,N_9869,N_9942);
nor U10312 (N_10312,N_9870,N_9896);
nand U10313 (N_10313,N_9550,N_9978);
or U10314 (N_10314,N_9552,N_9921);
or U10315 (N_10315,N_9526,N_9885);
and U10316 (N_10316,N_9912,N_9836);
nand U10317 (N_10317,N_9916,N_9903);
nand U10318 (N_10318,N_9700,N_9719);
or U10319 (N_10319,N_9606,N_9760);
and U10320 (N_10320,N_9683,N_9826);
and U10321 (N_10321,N_9780,N_9749);
and U10322 (N_10322,N_9563,N_9731);
nand U10323 (N_10323,N_9526,N_9663);
and U10324 (N_10324,N_9831,N_9695);
nor U10325 (N_10325,N_9671,N_9812);
or U10326 (N_10326,N_9933,N_9966);
xnor U10327 (N_10327,N_9811,N_9908);
nand U10328 (N_10328,N_9765,N_9565);
nand U10329 (N_10329,N_9930,N_9620);
nand U10330 (N_10330,N_9643,N_9775);
or U10331 (N_10331,N_9554,N_9729);
and U10332 (N_10332,N_9959,N_9912);
and U10333 (N_10333,N_9807,N_9749);
nor U10334 (N_10334,N_9615,N_9875);
or U10335 (N_10335,N_9818,N_9974);
nand U10336 (N_10336,N_9906,N_9593);
nand U10337 (N_10337,N_9755,N_9615);
and U10338 (N_10338,N_9662,N_9513);
or U10339 (N_10339,N_9635,N_9548);
nand U10340 (N_10340,N_9865,N_9752);
nand U10341 (N_10341,N_9752,N_9746);
nor U10342 (N_10342,N_9746,N_9665);
xnor U10343 (N_10343,N_9634,N_9751);
or U10344 (N_10344,N_9758,N_9642);
nand U10345 (N_10345,N_9588,N_9919);
nand U10346 (N_10346,N_9767,N_9937);
and U10347 (N_10347,N_9932,N_9913);
and U10348 (N_10348,N_9587,N_9748);
nand U10349 (N_10349,N_9550,N_9785);
or U10350 (N_10350,N_9807,N_9531);
and U10351 (N_10351,N_9583,N_9983);
nand U10352 (N_10352,N_9935,N_9823);
nand U10353 (N_10353,N_9882,N_9978);
or U10354 (N_10354,N_9778,N_9505);
and U10355 (N_10355,N_9658,N_9566);
nand U10356 (N_10356,N_9666,N_9567);
and U10357 (N_10357,N_9749,N_9792);
or U10358 (N_10358,N_9984,N_9784);
or U10359 (N_10359,N_9734,N_9565);
nand U10360 (N_10360,N_9625,N_9602);
and U10361 (N_10361,N_9853,N_9766);
nor U10362 (N_10362,N_9820,N_9919);
and U10363 (N_10363,N_9766,N_9518);
nand U10364 (N_10364,N_9607,N_9957);
or U10365 (N_10365,N_9877,N_9501);
or U10366 (N_10366,N_9841,N_9621);
and U10367 (N_10367,N_9504,N_9921);
nand U10368 (N_10368,N_9601,N_9649);
or U10369 (N_10369,N_9710,N_9836);
and U10370 (N_10370,N_9824,N_9781);
and U10371 (N_10371,N_9590,N_9696);
or U10372 (N_10372,N_9874,N_9578);
nand U10373 (N_10373,N_9841,N_9910);
or U10374 (N_10374,N_9563,N_9997);
and U10375 (N_10375,N_9534,N_9992);
and U10376 (N_10376,N_9526,N_9725);
and U10377 (N_10377,N_9634,N_9536);
nor U10378 (N_10378,N_9958,N_9616);
or U10379 (N_10379,N_9634,N_9529);
nand U10380 (N_10380,N_9699,N_9556);
nor U10381 (N_10381,N_9530,N_9680);
and U10382 (N_10382,N_9776,N_9501);
nor U10383 (N_10383,N_9693,N_9683);
and U10384 (N_10384,N_9969,N_9593);
nand U10385 (N_10385,N_9539,N_9502);
xnor U10386 (N_10386,N_9647,N_9508);
and U10387 (N_10387,N_9617,N_9788);
and U10388 (N_10388,N_9623,N_9574);
or U10389 (N_10389,N_9687,N_9973);
or U10390 (N_10390,N_9571,N_9891);
nor U10391 (N_10391,N_9976,N_9994);
nor U10392 (N_10392,N_9816,N_9981);
or U10393 (N_10393,N_9509,N_9606);
nand U10394 (N_10394,N_9962,N_9581);
or U10395 (N_10395,N_9952,N_9958);
nor U10396 (N_10396,N_9710,N_9597);
nand U10397 (N_10397,N_9940,N_9862);
or U10398 (N_10398,N_9971,N_9892);
nor U10399 (N_10399,N_9688,N_9783);
or U10400 (N_10400,N_9564,N_9765);
nand U10401 (N_10401,N_9840,N_9622);
nor U10402 (N_10402,N_9781,N_9682);
or U10403 (N_10403,N_9970,N_9694);
nor U10404 (N_10404,N_9831,N_9945);
nand U10405 (N_10405,N_9812,N_9897);
or U10406 (N_10406,N_9778,N_9980);
nand U10407 (N_10407,N_9847,N_9901);
or U10408 (N_10408,N_9883,N_9533);
nand U10409 (N_10409,N_9570,N_9781);
and U10410 (N_10410,N_9576,N_9798);
nor U10411 (N_10411,N_9899,N_9705);
or U10412 (N_10412,N_9651,N_9502);
nand U10413 (N_10413,N_9976,N_9977);
nor U10414 (N_10414,N_9919,N_9861);
and U10415 (N_10415,N_9533,N_9830);
or U10416 (N_10416,N_9746,N_9662);
nor U10417 (N_10417,N_9500,N_9970);
and U10418 (N_10418,N_9705,N_9970);
and U10419 (N_10419,N_9575,N_9952);
or U10420 (N_10420,N_9636,N_9891);
or U10421 (N_10421,N_9799,N_9773);
and U10422 (N_10422,N_9927,N_9557);
or U10423 (N_10423,N_9856,N_9947);
and U10424 (N_10424,N_9871,N_9937);
nand U10425 (N_10425,N_9837,N_9503);
and U10426 (N_10426,N_9823,N_9716);
nand U10427 (N_10427,N_9819,N_9692);
and U10428 (N_10428,N_9920,N_9789);
nand U10429 (N_10429,N_9971,N_9851);
nor U10430 (N_10430,N_9918,N_9874);
or U10431 (N_10431,N_9742,N_9697);
nand U10432 (N_10432,N_9682,N_9538);
nand U10433 (N_10433,N_9944,N_9880);
nor U10434 (N_10434,N_9666,N_9620);
or U10435 (N_10435,N_9651,N_9569);
or U10436 (N_10436,N_9914,N_9699);
nor U10437 (N_10437,N_9957,N_9701);
and U10438 (N_10438,N_9551,N_9605);
nor U10439 (N_10439,N_9993,N_9742);
nor U10440 (N_10440,N_9654,N_9558);
or U10441 (N_10441,N_9512,N_9668);
and U10442 (N_10442,N_9898,N_9631);
nor U10443 (N_10443,N_9694,N_9966);
or U10444 (N_10444,N_9724,N_9813);
and U10445 (N_10445,N_9802,N_9812);
nand U10446 (N_10446,N_9668,N_9581);
nand U10447 (N_10447,N_9751,N_9896);
and U10448 (N_10448,N_9725,N_9843);
nor U10449 (N_10449,N_9819,N_9937);
nor U10450 (N_10450,N_9892,N_9759);
and U10451 (N_10451,N_9744,N_9590);
and U10452 (N_10452,N_9502,N_9952);
and U10453 (N_10453,N_9537,N_9912);
and U10454 (N_10454,N_9653,N_9882);
or U10455 (N_10455,N_9929,N_9869);
nor U10456 (N_10456,N_9739,N_9747);
or U10457 (N_10457,N_9616,N_9553);
nand U10458 (N_10458,N_9954,N_9946);
and U10459 (N_10459,N_9827,N_9838);
or U10460 (N_10460,N_9632,N_9808);
nor U10461 (N_10461,N_9827,N_9599);
nor U10462 (N_10462,N_9970,N_9614);
nor U10463 (N_10463,N_9660,N_9618);
nand U10464 (N_10464,N_9669,N_9604);
nand U10465 (N_10465,N_9518,N_9898);
or U10466 (N_10466,N_9586,N_9911);
nand U10467 (N_10467,N_9722,N_9552);
or U10468 (N_10468,N_9726,N_9764);
nand U10469 (N_10469,N_9972,N_9681);
and U10470 (N_10470,N_9516,N_9685);
or U10471 (N_10471,N_9708,N_9684);
nand U10472 (N_10472,N_9521,N_9735);
or U10473 (N_10473,N_9707,N_9850);
and U10474 (N_10474,N_9676,N_9872);
nor U10475 (N_10475,N_9783,N_9770);
and U10476 (N_10476,N_9705,N_9977);
nand U10477 (N_10477,N_9876,N_9603);
or U10478 (N_10478,N_9684,N_9890);
nand U10479 (N_10479,N_9907,N_9970);
nand U10480 (N_10480,N_9859,N_9889);
or U10481 (N_10481,N_9919,N_9859);
nand U10482 (N_10482,N_9990,N_9707);
or U10483 (N_10483,N_9750,N_9759);
and U10484 (N_10484,N_9936,N_9801);
nor U10485 (N_10485,N_9579,N_9927);
nor U10486 (N_10486,N_9540,N_9788);
and U10487 (N_10487,N_9570,N_9797);
or U10488 (N_10488,N_9592,N_9752);
or U10489 (N_10489,N_9781,N_9911);
and U10490 (N_10490,N_9712,N_9825);
nand U10491 (N_10491,N_9768,N_9871);
nor U10492 (N_10492,N_9647,N_9969);
or U10493 (N_10493,N_9563,N_9669);
nor U10494 (N_10494,N_9555,N_9998);
nand U10495 (N_10495,N_9747,N_9521);
or U10496 (N_10496,N_9940,N_9538);
nand U10497 (N_10497,N_9658,N_9771);
and U10498 (N_10498,N_9757,N_9507);
and U10499 (N_10499,N_9730,N_9776);
or U10500 (N_10500,N_10304,N_10466);
or U10501 (N_10501,N_10452,N_10341);
nor U10502 (N_10502,N_10275,N_10338);
or U10503 (N_10503,N_10451,N_10321);
and U10504 (N_10504,N_10261,N_10032);
or U10505 (N_10505,N_10349,N_10203);
or U10506 (N_10506,N_10394,N_10404);
nand U10507 (N_10507,N_10296,N_10389);
or U10508 (N_10508,N_10298,N_10267);
nor U10509 (N_10509,N_10238,N_10386);
and U10510 (N_10510,N_10206,N_10056);
nand U10511 (N_10511,N_10020,N_10282);
nor U10512 (N_10512,N_10091,N_10196);
or U10513 (N_10513,N_10136,N_10019);
and U10514 (N_10514,N_10325,N_10262);
nand U10515 (N_10515,N_10132,N_10217);
nor U10516 (N_10516,N_10025,N_10215);
nor U10517 (N_10517,N_10312,N_10475);
nor U10518 (N_10518,N_10285,N_10142);
nor U10519 (N_10519,N_10185,N_10375);
or U10520 (N_10520,N_10313,N_10065);
and U10521 (N_10521,N_10301,N_10123);
nor U10522 (N_10522,N_10333,N_10414);
or U10523 (N_10523,N_10074,N_10357);
and U10524 (N_10524,N_10351,N_10278);
nor U10525 (N_10525,N_10226,N_10435);
and U10526 (N_10526,N_10096,N_10376);
and U10527 (N_10527,N_10080,N_10127);
nand U10528 (N_10528,N_10302,N_10399);
nor U10529 (N_10529,N_10381,N_10202);
nand U10530 (N_10530,N_10249,N_10059);
or U10531 (N_10531,N_10128,N_10210);
nand U10532 (N_10532,N_10200,N_10077);
nand U10533 (N_10533,N_10410,N_10244);
and U10534 (N_10534,N_10124,N_10446);
nor U10535 (N_10535,N_10177,N_10075);
nor U10536 (N_10536,N_10237,N_10067);
nand U10537 (N_10537,N_10009,N_10277);
nand U10538 (N_10538,N_10186,N_10078);
and U10539 (N_10539,N_10454,N_10055);
nor U10540 (N_10540,N_10288,N_10476);
and U10541 (N_10541,N_10168,N_10430);
and U10542 (N_10542,N_10489,N_10150);
nand U10543 (N_10543,N_10493,N_10497);
nand U10544 (N_10544,N_10485,N_10233);
nand U10545 (N_10545,N_10195,N_10264);
nand U10546 (N_10546,N_10016,N_10187);
and U10547 (N_10547,N_10022,N_10402);
or U10548 (N_10548,N_10141,N_10122);
or U10549 (N_10549,N_10204,N_10324);
nand U10550 (N_10550,N_10445,N_10212);
or U10551 (N_10551,N_10161,N_10384);
or U10552 (N_10552,N_10382,N_10440);
nor U10553 (N_10553,N_10283,N_10260);
or U10554 (N_10554,N_10052,N_10374);
nor U10555 (N_10555,N_10494,N_10042);
or U10556 (N_10556,N_10027,N_10164);
nand U10557 (N_10557,N_10450,N_10120);
nor U10558 (N_10558,N_10486,N_10295);
or U10559 (N_10559,N_10050,N_10409);
and U10560 (N_10560,N_10329,N_10490);
and U10561 (N_10561,N_10364,N_10099);
nor U10562 (N_10562,N_10255,N_10138);
nor U10563 (N_10563,N_10421,N_10133);
nand U10564 (N_10564,N_10112,N_10179);
or U10565 (N_10565,N_10129,N_10356);
nor U10566 (N_10566,N_10358,N_10343);
and U10567 (N_10567,N_10280,N_10315);
nand U10568 (N_10568,N_10148,N_10337);
nor U10569 (N_10569,N_10416,N_10378);
nand U10570 (N_10570,N_10235,N_10151);
nor U10571 (N_10571,N_10348,N_10170);
nor U10572 (N_10572,N_10095,N_10308);
or U10573 (N_10573,N_10429,N_10182);
nand U10574 (N_10574,N_10113,N_10463);
nor U10575 (N_10575,N_10330,N_10274);
nand U10576 (N_10576,N_10413,N_10455);
and U10577 (N_10577,N_10137,N_10085);
or U10578 (N_10578,N_10299,N_10054);
or U10579 (N_10579,N_10434,N_10039);
nor U10580 (N_10580,N_10420,N_10484);
or U10581 (N_10581,N_10332,N_10383);
and U10582 (N_10582,N_10363,N_10154);
nand U10583 (N_10583,N_10010,N_10201);
nor U10584 (N_10584,N_10172,N_10286);
or U10585 (N_10585,N_10145,N_10487);
nand U10586 (N_10586,N_10347,N_10492);
nor U10587 (N_10587,N_10388,N_10166);
and U10588 (N_10588,N_10232,N_10415);
nor U10589 (N_10589,N_10397,N_10071);
or U10590 (N_10590,N_10439,N_10030);
or U10591 (N_10591,N_10100,N_10335);
nand U10592 (N_10592,N_10360,N_10181);
nor U10593 (N_10593,N_10014,N_10292);
nor U10594 (N_10594,N_10370,N_10184);
xnor U10595 (N_10595,N_10121,N_10084);
nor U10596 (N_10596,N_10068,N_10322);
and U10597 (N_10597,N_10163,N_10005);
or U10598 (N_10598,N_10199,N_10353);
or U10599 (N_10599,N_10083,N_10246);
nor U10600 (N_10600,N_10241,N_10149);
or U10601 (N_10601,N_10218,N_10015);
and U10602 (N_10602,N_10311,N_10380);
or U10603 (N_10603,N_10422,N_10369);
nor U10604 (N_10604,N_10355,N_10104);
and U10605 (N_10605,N_10076,N_10205);
nor U10606 (N_10606,N_10208,N_10270);
nand U10607 (N_10607,N_10344,N_10481);
or U10608 (N_10608,N_10190,N_10222);
nand U10609 (N_10609,N_10368,N_10392);
or U10610 (N_10610,N_10064,N_10037);
nor U10611 (N_10611,N_10146,N_10290);
nand U10612 (N_10612,N_10098,N_10140);
nor U10613 (N_10613,N_10216,N_10488);
nand U10614 (N_10614,N_10066,N_10191);
or U10615 (N_10615,N_10013,N_10107);
and U10616 (N_10616,N_10259,N_10171);
nand U10617 (N_10617,N_10373,N_10437);
and U10618 (N_10618,N_10002,N_10243);
nand U10619 (N_10619,N_10453,N_10153);
nand U10620 (N_10620,N_10387,N_10209);
nor U10621 (N_10621,N_10044,N_10006);
nand U10622 (N_10622,N_10130,N_10183);
nor U10623 (N_10623,N_10478,N_10279);
nand U10624 (N_10624,N_10221,N_10316);
or U10625 (N_10625,N_10436,N_10427);
or U10626 (N_10626,N_10092,N_10155);
and U10627 (N_10627,N_10406,N_10291);
nand U10628 (N_10628,N_10459,N_10334);
and U10629 (N_10629,N_10034,N_10281);
nor U10630 (N_10630,N_10319,N_10362);
xnor U10631 (N_10631,N_10424,N_10371);
nand U10632 (N_10632,N_10496,N_10017);
nand U10633 (N_10633,N_10156,N_10461);
nand U10634 (N_10634,N_10297,N_10023);
nor U10635 (N_10635,N_10135,N_10405);
nor U10636 (N_10636,N_10088,N_10001);
nor U10637 (N_10637,N_10234,N_10167);
and U10638 (N_10638,N_10224,N_10038);
and U10639 (N_10639,N_10467,N_10225);
and U10640 (N_10640,N_10116,N_10284);
and U10641 (N_10641,N_10125,N_10102);
nand U10642 (N_10642,N_10139,N_10118);
or U10643 (N_10643,N_10081,N_10214);
nor U10644 (N_10644,N_10043,N_10331);
nand U10645 (N_10645,N_10131,N_10162);
nor U10646 (N_10646,N_10469,N_10143);
and U10647 (N_10647,N_10287,N_10213);
or U10648 (N_10648,N_10499,N_10060);
or U10649 (N_10649,N_10053,N_10176);
nor U10650 (N_10650,N_10342,N_10035);
and U10651 (N_10651,N_10423,N_10227);
nand U10652 (N_10652,N_10041,N_10008);
or U10653 (N_10653,N_10033,N_10289);
nand U10654 (N_10654,N_10336,N_10328);
and U10655 (N_10655,N_10158,N_10094);
and U10656 (N_10656,N_10411,N_10266);
and U10657 (N_10657,N_10441,N_10093);
or U10658 (N_10658,N_10443,N_10194);
and U10659 (N_10659,N_10385,N_10174);
or U10660 (N_10660,N_10026,N_10231);
or U10661 (N_10661,N_10400,N_10470);
nor U10662 (N_10662,N_10449,N_10219);
and U10663 (N_10663,N_10004,N_10101);
or U10664 (N_10664,N_10152,N_10211);
nand U10665 (N_10665,N_10359,N_10178);
nor U10666 (N_10666,N_10391,N_10007);
nor U10667 (N_10667,N_10103,N_10256);
nand U10668 (N_10668,N_10448,N_10157);
and U10669 (N_10669,N_10165,N_10072);
nand U10670 (N_10670,N_10126,N_10407);
nand U10671 (N_10671,N_10265,N_10117);
nand U10672 (N_10672,N_10310,N_10401);
or U10673 (N_10673,N_10115,N_10040);
nor U10674 (N_10674,N_10021,N_10229);
or U10675 (N_10675,N_10272,N_10498);
nor U10676 (N_10676,N_10079,N_10365);
and U10677 (N_10677,N_10361,N_10012);
and U10678 (N_10678,N_10379,N_10327);
and U10679 (N_10679,N_10108,N_10198);
nand U10680 (N_10680,N_10144,N_10228);
and U10681 (N_10681,N_10134,N_10110);
or U10682 (N_10682,N_10105,N_10058);
nor U10683 (N_10683,N_10390,N_10300);
nor U10684 (N_10684,N_10169,N_10495);
nor U10685 (N_10685,N_10426,N_10082);
or U10686 (N_10686,N_10046,N_10028);
or U10687 (N_10687,N_10097,N_10396);
nor U10688 (N_10688,N_10431,N_10367);
nor U10689 (N_10689,N_10307,N_10428);
nand U10690 (N_10690,N_10269,N_10412);
and U10691 (N_10691,N_10003,N_10048);
or U10692 (N_10692,N_10257,N_10419);
nor U10693 (N_10693,N_10483,N_10061);
or U10694 (N_10694,N_10031,N_10273);
or U10695 (N_10695,N_10073,N_10480);
and U10696 (N_10696,N_10248,N_10220);
or U10697 (N_10697,N_10477,N_10000);
nor U10698 (N_10698,N_10189,N_10377);
nor U10699 (N_10699,N_10447,N_10339);
nor U10700 (N_10700,N_10147,N_10456);
nor U10701 (N_10701,N_10069,N_10294);
and U10702 (N_10702,N_10251,N_10111);
and U10703 (N_10703,N_10045,N_10245);
or U10704 (N_10704,N_10057,N_10063);
and U10705 (N_10705,N_10372,N_10087);
and U10706 (N_10706,N_10395,N_10086);
nor U10707 (N_10707,N_10323,N_10354);
nor U10708 (N_10708,N_10193,N_10305);
nand U10709 (N_10709,N_10047,N_10340);
and U10710 (N_10710,N_10018,N_10403);
xnor U10711 (N_10711,N_10471,N_10114);
and U10712 (N_10712,N_10417,N_10051);
or U10713 (N_10713,N_10464,N_10223);
nand U10714 (N_10714,N_10029,N_10011);
and U10715 (N_10715,N_10036,N_10089);
or U10716 (N_10716,N_10366,N_10460);
nor U10717 (N_10717,N_10458,N_10345);
or U10718 (N_10718,N_10318,N_10254);
nand U10719 (N_10719,N_10293,N_10468);
and U10720 (N_10720,N_10309,N_10457);
or U10721 (N_10721,N_10320,N_10433);
nor U10722 (N_10722,N_10444,N_10062);
and U10723 (N_10723,N_10159,N_10024);
nor U10724 (N_10724,N_10398,N_10239);
nand U10725 (N_10725,N_10160,N_10268);
nor U10726 (N_10726,N_10236,N_10306);
nand U10727 (N_10727,N_10242,N_10109);
nor U10728 (N_10728,N_10326,N_10250);
or U10729 (N_10729,N_10240,N_10192);
nor U10730 (N_10730,N_10197,N_10474);
and U10731 (N_10731,N_10070,N_10393);
nand U10732 (N_10732,N_10090,N_10252);
or U10733 (N_10733,N_10425,N_10173);
nor U10734 (N_10734,N_10207,N_10350);
nand U10735 (N_10735,N_10247,N_10473);
or U10736 (N_10736,N_10253,N_10188);
nor U10737 (N_10737,N_10346,N_10442);
nand U10738 (N_10738,N_10317,N_10352);
or U10739 (N_10739,N_10119,N_10432);
or U10740 (N_10740,N_10418,N_10482);
or U10741 (N_10741,N_10180,N_10491);
or U10742 (N_10742,N_10408,N_10271);
nand U10743 (N_10743,N_10230,N_10258);
or U10744 (N_10744,N_10276,N_10472);
nor U10745 (N_10745,N_10438,N_10263);
nand U10746 (N_10746,N_10175,N_10465);
nand U10747 (N_10747,N_10462,N_10314);
and U10748 (N_10748,N_10479,N_10303);
or U10749 (N_10749,N_10049,N_10106);
and U10750 (N_10750,N_10000,N_10008);
nand U10751 (N_10751,N_10236,N_10328);
or U10752 (N_10752,N_10302,N_10387);
nand U10753 (N_10753,N_10104,N_10148);
nor U10754 (N_10754,N_10175,N_10348);
nor U10755 (N_10755,N_10095,N_10051);
nand U10756 (N_10756,N_10413,N_10456);
nand U10757 (N_10757,N_10097,N_10156);
and U10758 (N_10758,N_10006,N_10012);
or U10759 (N_10759,N_10426,N_10391);
and U10760 (N_10760,N_10202,N_10203);
nand U10761 (N_10761,N_10208,N_10211);
or U10762 (N_10762,N_10247,N_10103);
or U10763 (N_10763,N_10131,N_10199);
nand U10764 (N_10764,N_10027,N_10494);
and U10765 (N_10765,N_10289,N_10457);
nand U10766 (N_10766,N_10264,N_10037);
and U10767 (N_10767,N_10249,N_10024);
and U10768 (N_10768,N_10139,N_10049);
or U10769 (N_10769,N_10346,N_10485);
or U10770 (N_10770,N_10296,N_10409);
nand U10771 (N_10771,N_10478,N_10280);
nor U10772 (N_10772,N_10419,N_10152);
nor U10773 (N_10773,N_10019,N_10058);
nor U10774 (N_10774,N_10334,N_10287);
or U10775 (N_10775,N_10489,N_10038);
and U10776 (N_10776,N_10451,N_10439);
and U10777 (N_10777,N_10348,N_10484);
nand U10778 (N_10778,N_10089,N_10320);
nor U10779 (N_10779,N_10115,N_10308);
and U10780 (N_10780,N_10384,N_10207);
or U10781 (N_10781,N_10456,N_10486);
or U10782 (N_10782,N_10419,N_10453);
and U10783 (N_10783,N_10029,N_10154);
nor U10784 (N_10784,N_10155,N_10434);
nand U10785 (N_10785,N_10418,N_10357);
or U10786 (N_10786,N_10095,N_10024);
nor U10787 (N_10787,N_10059,N_10093);
nor U10788 (N_10788,N_10393,N_10305);
nand U10789 (N_10789,N_10256,N_10407);
and U10790 (N_10790,N_10424,N_10268);
nor U10791 (N_10791,N_10333,N_10446);
nand U10792 (N_10792,N_10394,N_10346);
nand U10793 (N_10793,N_10103,N_10061);
nor U10794 (N_10794,N_10443,N_10130);
nor U10795 (N_10795,N_10300,N_10283);
nand U10796 (N_10796,N_10483,N_10157);
nand U10797 (N_10797,N_10294,N_10471);
nand U10798 (N_10798,N_10197,N_10131);
nor U10799 (N_10799,N_10049,N_10348);
nand U10800 (N_10800,N_10429,N_10234);
nor U10801 (N_10801,N_10472,N_10242);
and U10802 (N_10802,N_10439,N_10048);
nand U10803 (N_10803,N_10230,N_10157);
or U10804 (N_10804,N_10457,N_10490);
and U10805 (N_10805,N_10419,N_10479);
or U10806 (N_10806,N_10031,N_10252);
nand U10807 (N_10807,N_10073,N_10142);
nand U10808 (N_10808,N_10354,N_10285);
nand U10809 (N_10809,N_10477,N_10247);
nor U10810 (N_10810,N_10310,N_10050);
and U10811 (N_10811,N_10342,N_10126);
nor U10812 (N_10812,N_10483,N_10111);
and U10813 (N_10813,N_10472,N_10115);
nor U10814 (N_10814,N_10414,N_10098);
nand U10815 (N_10815,N_10464,N_10321);
and U10816 (N_10816,N_10381,N_10472);
or U10817 (N_10817,N_10398,N_10330);
and U10818 (N_10818,N_10389,N_10468);
and U10819 (N_10819,N_10233,N_10452);
or U10820 (N_10820,N_10077,N_10182);
nor U10821 (N_10821,N_10444,N_10206);
nand U10822 (N_10822,N_10264,N_10029);
or U10823 (N_10823,N_10299,N_10005);
or U10824 (N_10824,N_10407,N_10339);
and U10825 (N_10825,N_10099,N_10037);
or U10826 (N_10826,N_10259,N_10317);
xnor U10827 (N_10827,N_10363,N_10071);
nor U10828 (N_10828,N_10197,N_10186);
or U10829 (N_10829,N_10070,N_10376);
nand U10830 (N_10830,N_10434,N_10294);
nand U10831 (N_10831,N_10329,N_10220);
nor U10832 (N_10832,N_10335,N_10408);
nand U10833 (N_10833,N_10478,N_10317);
nor U10834 (N_10834,N_10366,N_10382);
and U10835 (N_10835,N_10003,N_10171);
or U10836 (N_10836,N_10431,N_10165);
and U10837 (N_10837,N_10179,N_10219);
and U10838 (N_10838,N_10216,N_10226);
or U10839 (N_10839,N_10176,N_10444);
or U10840 (N_10840,N_10122,N_10018);
and U10841 (N_10841,N_10275,N_10331);
or U10842 (N_10842,N_10410,N_10412);
or U10843 (N_10843,N_10179,N_10225);
nand U10844 (N_10844,N_10030,N_10210);
or U10845 (N_10845,N_10200,N_10033);
or U10846 (N_10846,N_10148,N_10293);
and U10847 (N_10847,N_10234,N_10122);
nor U10848 (N_10848,N_10295,N_10499);
or U10849 (N_10849,N_10287,N_10307);
or U10850 (N_10850,N_10109,N_10058);
and U10851 (N_10851,N_10396,N_10198);
nand U10852 (N_10852,N_10144,N_10273);
xor U10853 (N_10853,N_10124,N_10024);
nand U10854 (N_10854,N_10433,N_10099);
nand U10855 (N_10855,N_10417,N_10339);
or U10856 (N_10856,N_10072,N_10058);
nand U10857 (N_10857,N_10254,N_10165);
and U10858 (N_10858,N_10240,N_10457);
and U10859 (N_10859,N_10370,N_10101);
nand U10860 (N_10860,N_10355,N_10196);
nand U10861 (N_10861,N_10115,N_10273);
nor U10862 (N_10862,N_10118,N_10375);
and U10863 (N_10863,N_10062,N_10269);
nor U10864 (N_10864,N_10394,N_10224);
nor U10865 (N_10865,N_10443,N_10396);
nor U10866 (N_10866,N_10457,N_10482);
nor U10867 (N_10867,N_10463,N_10292);
nor U10868 (N_10868,N_10033,N_10480);
or U10869 (N_10869,N_10476,N_10297);
and U10870 (N_10870,N_10078,N_10146);
nor U10871 (N_10871,N_10167,N_10154);
nor U10872 (N_10872,N_10315,N_10361);
nand U10873 (N_10873,N_10157,N_10088);
nand U10874 (N_10874,N_10093,N_10495);
nor U10875 (N_10875,N_10480,N_10001);
or U10876 (N_10876,N_10455,N_10482);
nor U10877 (N_10877,N_10073,N_10384);
nand U10878 (N_10878,N_10353,N_10168);
or U10879 (N_10879,N_10256,N_10298);
and U10880 (N_10880,N_10094,N_10364);
and U10881 (N_10881,N_10249,N_10083);
nor U10882 (N_10882,N_10347,N_10013);
nor U10883 (N_10883,N_10473,N_10119);
nor U10884 (N_10884,N_10265,N_10230);
nand U10885 (N_10885,N_10291,N_10005);
nand U10886 (N_10886,N_10388,N_10099);
nand U10887 (N_10887,N_10150,N_10367);
or U10888 (N_10888,N_10428,N_10275);
nand U10889 (N_10889,N_10463,N_10078);
nor U10890 (N_10890,N_10213,N_10373);
or U10891 (N_10891,N_10036,N_10368);
or U10892 (N_10892,N_10011,N_10466);
or U10893 (N_10893,N_10266,N_10055);
or U10894 (N_10894,N_10131,N_10081);
and U10895 (N_10895,N_10482,N_10478);
and U10896 (N_10896,N_10016,N_10057);
nor U10897 (N_10897,N_10253,N_10062);
nand U10898 (N_10898,N_10311,N_10464);
and U10899 (N_10899,N_10254,N_10123);
and U10900 (N_10900,N_10006,N_10188);
nor U10901 (N_10901,N_10111,N_10075);
nor U10902 (N_10902,N_10142,N_10398);
and U10903 (N_10903,N_10103,N_10166);
nand U10904 (N_10904,N_10471,N_10483);
and U10905 (N_10905,N_10328,N_10200);
nand U10906 (N_10906,N_10441,N_10449);
xor U10907 (N_10907,N_10328,N_10058);
or U10908 (N_10908,N_10214,N_10350);
xor U10909 (N_10909,N_10013,N_10404);
nand U10910 (N_10910,N_10141,N_10406);
nor U10911 (N_10911,N_10159,N_10163);
or U10912 (N_10912,N_10066,N_10480);
nand U10913 (N_10913,N_10276,N_10413);
and U10914 (N_10914,N_10235,N_10126);
and U10915 (N_10915,N_10120,N_10130);
nor U10916 (N_10916,N_10032,N_10122);
and U10917 (N_10917,N_10199,N_10223);
nor U10918 (N_10918,N_10335,N_10158);
and U10919 (N_10919,N_10055,N_10321);
nor U10920 (N_10920,N_10049,N_10426);
or U10921 (N_10921,N_10308,N_10440);
and U10922 (N_10922,N_10077,N_10105);
nor U10923 (N_10923,N_10012,N_10438);
nor U10924 (N_10924,N_10071,N_10320);
and U10925 (N_10925,N_10126,N_10026);
nor U10926 (N_10926,N_10078,N_10072);
or U10927 (N_10927,N_10409,N_10255);
or U10928 (N_10928,N_10499,N_10235);
nand U10929 (N_10929,N_10160,N_10052);
nand U10930 (N_10930,N_10096,N_10046);
nand U10931 (N_10931,N_10394,N_10344);
or U10932 (N_10932,N_10232,N_10389);
nand U10933 (N_10933,N_10482,N_10047);
or U10934 (N_10934,N_10017,N_10265);
or U10935 (N_10935,N_10241,N_10431);
or U10936 (N_10936,N_10116,N_10151);
nor U10937 (N_10937,N_10400,N_10343);
or U10938 (N_10938,N_10365,N_10342);
nand U10939 (N_10939,N_10476,N_10281);
nand U10940 (N_10940,N_10103,N_10454);
nand U10941 (N_10941,N_10477,N_10273);
or U10942 (N_10942,N_10032,N_10129);
nor U10943 (N_10943,N_10359,N_10463);
and U10944 (N_10944,N_10278,N_10177);
or U10945 (N_10945,N_10120,N_10493);
and U10946 (N_10946,N_10334,N_10223);
nand U10947 (N_10947,N_10080,N_10221);
nand U10948 (N_10948,N_10096,N_10224);
nand U10949 (N_10949,N_10310,N_10201);
nor U10950 (N_10950,N_10410,N_10347);
and U10951 (N_10951,N_10480,N_10040);
or U10952 (N_10952,N_10201,N_10258);
nor U10953 (N_10953,N_10036,N_10438);
nand U10954 (N_10954,N_10437,N_10027);
nor U10955 (N_10955,N_10169,N_10115);
and U10956 (N_10956,N_10253,N_10337);
nand U10957 (N_10957,N_10447,N_10280);
and U10958 (N_10958,N_10105,N_10463);
nand U10959 (N_10959,N_10359,N_10222);
or U10960 (N_10960,N_10417,N_10408);
nor U10961 (N_10961,N_10470,N_10244);
or U10962 (N_10962,N_10222,N_10373);
and U10963 (N_10963,N_10410,N_10036);
and U10964 (N_10964,N_10274,N_10182);
nand U10965 (N_10965,N_10145,N_10317);
nor U10966 (N_10966,N_10125,N_10362);
nand U10967 (N_10967,N_10427,N_10195);
and U10968 (N_10968,N_10226,N_10065);
and U10969 (N_10969,N_10182,N_10028);
nor U10970 (N_10970,N_10146,N_10355);
or U10971 (N_10971,N_10286,N_10108);
and U10972 (N_10972,N_10456,N_10250);
and U10973 (N_10973,N_10106,N_10092);
nor U10974 (N_10974,N_10077,N_10479);
and U10975 (N_10975,N_10484,N_10114);
nand U10976 (N_10976,N_10313,N_10188);
nor U10977 (N_10977,N_10383,N_10095);
or U10978 (N_10978,N_10447,N_10463);
nand U10979 (N_10979,N_10203,N_10068);
and U10980 (N_10980,N_10366,N_10049);
and U10981 (N_10981,N_10479,N_10258);
nor U10982 (N_10982,N_10253,N_10007);
and U10983 (N_10983,N_10098,N_10047);
nor U10984 (N_10984,N_10390,N_10362);
and U10985 (N_10985,N_10425,N_10434);
nand U10986 (N_10986,N_10401,N_10074);
nor U10987 (N_10987,N_10075,N_10424);
nand U10988 (N_10988,N_10312,N_10299);
nand U10989 (N_10989,N_10496,N_10183);
nand U10990 (N_10990,N_10451,N_10351);
nand U10991 (N_10991,N_10367,N_10232);
nand U10992 (N_10992,N_10309,N_10201);
or U10993 (N_10993,N_10271,N_10367);
or U10994 (N_10994,N_10271,N_10309);
nor U10995 (N_10995,N_10271,N_10377);
nand U10996 (N_10996,N_10191,N_10195);
or U10997 (N_10997,N_10273,N_10289);
nand U10998 (N_10998,N_10331,N_10026);
or U10999 (N_10999,N_10386,N_10433);
and U11000 (N_11000,N_10861,N_10628);
nand U11001 (N_11001,N_10597,N_10799);
nor U11002 (N_11002,N_10513,N_10981);
or U11003 (N_11003,N_10883,N_10582);
and U11004 (N_11004,N_10857,N_10721);
nand U11005 (N_11005,N_10870,N_10918);
nand U11006 (N_11006,N_10923,N_10874);
nand U11007 (N_11007,N_10932,N_10689);
nand U11008 (N_11008,N_10632,N_10949);
nand U11009 (N_11009,N_10617,N_10655);
or U11010 (N_11010,N_10723,N_10577);
nor U11011 (N_11011,N_10809,N_10562);
or U11012 (N_11012,N_10877,N_10840);
or U11013 (N_11013,N_10630,N_10916);
nor U11014 (N_11014,N_10605,N_10800);
nor U11015 (N_11015,N_10727,N_10853);
or U11016 (N_11016,N_10903,N_10591);
or U11017 (N_11017,N_10604,N_10561);
and U11018 (N_11018,N_10624,N_10671);
nor U11019 (N_11019,N_10948,N_10578);
nand U11020 (N_11020,N_10964,N_10696);
nor U11021 (N_11021,N_10635,N_10784);
nor U11022 (N_11022,N_10838,N_10554);
nand U11023 (N_11023,N_10525,N_10538);
or U11024 (N_11024,N_10622,N_10517);
nand U11025 (N_11025,N_10897,N_10753);
and U11026 (N_11026,N_10703,N_10810);
nor U11027 (N_11027,N_10640,N_10771);
nand U11028 (N_11028,N_10946,N_10669);
nand U11029 (N_11029,N_10894,N_10855);
or U11030 (N_11030,N_10930,N_10712);
nand U11031 (N_11031,N_10869,N_10974);
nor U11032 (N_11032,N_10673,N_10588);
or U11033 (N_11033,N_10720,N_10973);
nand U11034 (N_11034,N_10953,N_10514);
nand U11035 (N_11035,N_10746,N_10748);
nand U11036 (N_11036,N_10831,N_10885);
nor U11037 (N_11037,N_10958,N_10739);
nor U11038 (N_11038,N_10821,N_10917);
nor U11039 (N_11039,N_10965,N_10601);
nand U11040 (N_11040,N_10787,N_10537);
nand U11041 (N_11041,N_10573,N_10995);
and U11042 (N_11042,N_10834,N_10585);
nor U11043 (N_11043,N_10811,N_10820);
and U11044 (N_11044,N_10994,N_10543);
nand U11045 (N_11045,N_10744,N_10891);
nor U11046 (N_11046,N_10901,N_10507);
or U11047 (N_11047,N_10652,N_10825);
nand U11048 (N_11048,N_10716,N_10631);
or U11049 (N_11049,N_10709,N_10590);
or U11050 (N_11050,N_10725,N_10828);
nand U11051 (N_11051,N_10648,N_10523);
nand U11052 (N_11052,N_10895,N_10976);
or U11053 (N_11053,N_10788,N_10541);
or U11054 (N_11054,N_10919,N_10618);
or U11055 (N_11055,N_10553,N_10830);
nor U11056 (N_11056,N_10872,N_10770);
nand U11057 (N_11057,N_10867,N_10627);
nand U11058 (N_11058,N_10643,N_10647);
or U11059 (N_11059,N_10683,N_10697);
and U11060 (N_11060,N_10674,N_10659);
or U11061 (N_11061,N_10583,N_10576);
or U11062 (N_11062,N_10993,N_10778);
nor U11063 (N_11063,N_10760,N_10656);
or U11064 (N_11064,N_10888,N_10847);
or U11065 (N_11065,N_10915,N_10959);
and U11066 (N_11066,N_10592,N_10729);
nand U11067 (N_11067,N_10851,N_10952);
nand U11068 (N_11068,N_10580,N_10556);
nand U11069 (N_11069,N_10774,N_10572);
nor U11070 (N_11070,N_10984,N_10505);
and U11071 (N_11071,N_10661,N_10791);
or U11072 (N_11072,N_10611,N_10693);
and U11073 (N_11073,N_10986,N_10741);
nor U11074 (N_11074,N_10772,N_10910);
nor U11075 (N_11075,N_10531,N_10927);
or U11076 (N_11076,N_10502,N_10710);
or U11077 (N_11077,N_10728,N_10747);
nand U11078 (N_11078,N_10503,N_10719);
and U11079 (N_11079,N_10909,N_10519);
or U11080 (N_11080,N_10680,N_10570);
nor U11081 (N_11081,N_10929,N_10990);
nor U11082 (N_11082,N_10856,N_10908);
nor U11083 (N_11083,N_10650,N_10694);
and U11084 (N_11084,N_10904,N_10567);
and U11085 (N_11085,N_10866,N_10603);
nand U11086 (N_11086,N_10609,N_10718);
nor U11087 (N_11087,N_10623,N_10742);
nand U11088 (N_11088,N_10815,N_10805);
nand U11089 (N_11089,N_10859,N_10688);
and U11090 (N_11090,N_10676,N_10907);
nand U11091 (N_11091,N_10945,N_10599);
and U11092 (N_11092,N_10690,N_10706);
or U11093 (N_11093,N_10947,N_10938);
and U11094 (N_11094,N_10707,N_10510);
nor U11095 (N_11095,N_10657,N_10685);
or U11096 (N_11096,N_10873,N_10566);
nor U11097 (N_11097,N_10983,N_10612);
and U11098 (N_11098,N_10509,N_10698);
nand U11099 (N_11099,N_10822,N_10768);
and U11100 (N_11100,N_10886,N_10996);
nor U11101 (N_11101,N_10782,N_10971);
nor U11102 (N_11102,N_10549,N_10813);
and U11103 (N_11103,N_10975,N_10950);
nand U11104 (N_11104,N_10944,N_10646);
nor U11105 (N_11105,N_10645,N_10881);
and U11106 (N_11106,N_10960,N_10786);
or U11107 (N_11107,N_10559,N_10518);
nand U11108 (N_11108,N_10783,N_10779);
and U11109 (N_11109,N_10878,N_10527);
or U11110 (N_11110,N_10684,N_10569);
or U11111 (N_11111,N_10966,N_10803);
nand U11112 (N_11112,N_10922,N_10763);
and U11113 (N_11113,N_10515,N_10546);
and U11114 (N_11114,N_10890,N_10615);
nand U11115 (N_11115,N_10936,N_10875);
nand U11116 (N_11116,N_10766,N_10846);
nand U11117 (N_11117,N_10662,N_10529);
nor U11118 (N_11118,N_10636,N_10539);
xnor U11119 (N_11119,N_10790,N_10862);
and U11120 (N_11120,N_10621,N_10841);
and U11121 (N_11121,N_10535,N_10731);
or U11122 (N_11122,N_10607,N_10972);
or U11123 (N_11123,N_10668,N_10914);
nor U11124 (N_11124,N_10955,N_10951);
nand U11125 (N_11125,N_10667,N_10776);
nor U11126 (N_11126,N_10963,N_10899);
or U11127 (N_11127,N_10681,N_10620);
nand U11128 (N_11128,N_10928,N_10780);
nor U11129 (N_11129,N_10893,N_10586);
or U11130 (N_11130,N_10797,N_10575);
nor U11131 (N_11131,N_10817,N_10839);
nor U11132 (N_11132,N_10987,N_10924);
nand U11133 (N_11133,N_10902,N_10508);
or U11134 (N_11134,N_10773,N_10702);
or U11135 (N_11135,N_10608,N_10550);
nand U11136 (N_11136,N_10563,N_10602);
nor U11137 (N_11137,N_10835,N_10581);
nand U11138 (N_11138,N_10865,N_10610);
and U11139 (N_11139,N_10935,N_10524);
or U11140 (N_11140,N_10644,N_10734);
and U11141 (N_11141,N_10552,N_10536);
and U11142 (N_11142,N_10584,N_10896);
or U11143 (N_11143,N_10804,N_10695);
and U11144 (N_11144,N_10967,N_10732);
and U11145 (N_11145,N_10794,N_10551);
or U11146 (N_11146,N_10638,N_10977);
nor U11147 (N_11147,N_10724,N_10606);
and U11148 (N_11148,N_10526,N_10943);
nor U11149 (N_11149,N_10837,N_10557);
or U11150 (N_11150,N_10666,N_10845);
nand U11151 (N_11151,N_10547,N_10660);
or U11152 (N_11152,N_10682,N_10767);
or U11153 (N_11153,N_10613,N_10860);
and U11154 (N_11154,N_10769,N_10997);
nand U11155 (N_11155,N_10882,N_10651);
nand U11156 (N_11156,N_10957,N_10989);
and U11157 (N_11157,N_10876,N_10675);
or U11158 (N_11158,N_10740,N_10634);
and U11159 (N_11159,N_10921,N_10812);
nor U11160 (N_11160,N_10992,N_10678);
or U11161 (N_11161,N_10751,N_10900);
and U11162 (N_11162,N_10934,N_10844);
and U11163 (N_11163,N_10642,N_10555);
nor U11164 (N_11164,N_10879,N_10985);
and U11165 (N_11165,N_10755,N_10762);
nand U11166 (N_11166,N_10653,N_10871);
nand U11167 (N_11167,N_10758,N_10991);
nand U11168 (N_11168,N_10892,N_10745);
nor U11169 (N_11169,N_10801,N_10665);
nand U11170 (N_11170,N_10884,N_10558);
nand U11171 (N_11171,N_10864,N_10880);
nand U11172 (N_11172,N_10511,N_10594);
or U11173 (N_11173,N_10789,N_10752);
nor U11174 (N_11174,N_10733,N_10593);
and U11175 (N_11175,N_10616,N_10970);
nor U11176 (N_11176,N_10614,N_10574);
nor U11177 (N_11177,N_10641,N_10564);
or U11178 (N_11178,N_10520,N_10819);
and U11179 (N_11179,N_10625,N_10889);
or U11180 (N_11180,N_10522,N_10629);
nor U11181 (N_11181,N_10824,N_10814);
nor U11182 (N_11182,N_10686,N_10931);
and U11183 (N_11183,N_10670,N_10626);
nor U11184 (N_11184,N_10722,N_10540);
nor U11185 (N_11185,N_10806,N_10761);
and U11186 (N_11186,N_10713,N_10939);
and U11187 (N_11187,N_10836,N_10542);
or U11188 (N_11188,N_10568,N_10595);
and U11189 (N_11189,N_10548,N_10798);
or U11190 (N_11190,N_10600,N_10887);
or U11191 (N_11191,N_10701,N_10749);
and U11192 (N_11192,N_10961,N_10850);
nand U11193 (N_11193,N_10998,N_10726);
and U11194 (N_11194,N_10757,N_10925);
and U11195 (N_11195,N_10793,N_10750);
nor U11196 (N_11196,N_10905,N_10705);
and U11197 (N_11197,N_10823,N_10692);
nand U11198 (N_11198,N_10735,N_10565);
nor U11199 (N_11199,N_10979,N_10544);
and U11200 (N_11200,N_10816,N_10940);
and U11201 (N_11201,N_10598,N_10920);
nor U11202 (N_11202,N_10933,N_10663);
nor U11203 (N_11203,N_10699,N_10639);
and U11204 (N_11204,N_10765,N_10978);
nor U11205 (N_11205,N_10802,N_10738);
nor U11206 (N_11206,N_10528,N_10937);
nand U11207 (N_11207,N_10941,N_10818);
nand U11208 (N_11208,N_10504,N_10516);
or U11209 (N_11209,N_10730,N_10827);
nor U11210 (N_11210,N_10980,N_10579);
nor U11211 (N_11211,N_10808,N_10700);
nor U11212 (N_11212,N_10832,N_10911);
nand U11213 (N_11213,N_10968,N_10999);
nor U11214 (N_11214,N_10868,N_10795);
nand U11215 (N_11215,N_10781,N_10717);
nand U11216 (N_11216,N_10708,N_10852);
nand U11217 (N_11217,N_10956,N_10654);
or U11218 (N_11218,N_10506,N_10982);
nor U11219 (N_11219,N_10988,N_10842);
and U11220 (N_11220,N_10633,N_10954);
and U11221 (N_11221,N_10545,N_10807);
and U11222 (N_11222,N_10637,N_10926);
nor U11223 (N_11223,N_10658,N_10711);
nand U11224 (N_11224,N_10687,N_10843);
and U11225 (N_11225,N_10596,N_10587);
or U11226 (N_11226,N_10737,N_10619);
nor U11227 (N_11227,N_10826,N_10649);
or U11228 (N_11228,N_10679,N_10533);
nor U11229 (N_11229,N_10500,N_10759);
and U11230 (N_11230,N_10691,N_10942);
nor U11231 (N_11231,N_10530,N_10785);
nand U11232 (N_11232,N_10589,N_10571);
nor U11233 (N_11233,N_10501,N_10792);
nor U11234 (N_11234,N_10672,N_10736);
and U11235 (N_11235,N_10833,N_10898);
nand U11236 (N_11236,N_10863,N_10969);
and U11237 (N_11237,N_10743,N_10677);
nand U11238 (N_11238,N_10777,N_10534);
and U11239 (N_11239,N_10913,N_10560);
and U11240 (N_11240,N_10704,N_10715);
and U11241 (N_11241,N_10796,N_10714);
and U11242 (N_11242,N_10854,N_10764);
nor U11243 (N_11243,N_10858,N_10775);
or U11244 (N_11244,N_10512,N_10829);
nand U11245 (N_11245,N_10756,N_10848);
nor U11246 (N_11246,N_10962,N_10521);
nor U11247 (N_11247,N_10912,N_10532);
nand U11248 (N_11248,N_10849,N_10664);
xnor U11249 (N_11249,N_10906,N_10754);
or U11250 (N_11250,N_10932,N_10860);
nor U11251 (N_11251,N_10566,N_10953);
nand U11252 (N_11252,N_10518,N_10717);
or U11253 (N_11253,N_10523,N_10676);
nor U11254 (N_11254,N_10717,N_10522);
or U11255 (N_11255,N_10877,N_10948);
or U11256 (N_11256,N_10585,N_10954);
nand U11257 (N_11257,N_10922,N_10849);
and U11258 (N_11258,N_10880,N_10701);
nand U11259 (N_11259,N_10688,N_10797);
and U11260 (N_11260,N_10584,N_10845);
nand U11261 (N_11261,N_10793,N_10620);
nand U11262 (N_11262,N_10577,N_10694);
or U11263 (N_11263,N_10579,N_10949);
or U11264 (N_11264,N_10950,N_10730);
nand U11265 (N_11265,N_10928,N_10611);
and U11266 (N_11266,N_10858,N_10844);
or U11267 (N_11267,N_10806,N_10619);
or U11268 (N_11268,N_10912,N_10650);
nand U11269 (N_11269,N_10585,N_10606);
nand U11270 (N_11270,N_10745,N_10999);
and U11271 (N_11271,N_10896,N_10741);
or U11272 (N_11272,N_10583,N_10585);
and U11273 (N_11273,N_10551,N_10695);
nand U11274 (N_11274,N_10771,N_10624);
or U11275 (N_11275,N_10507,N_10738);
or U11276 (N_11276,N_10611,N_10837);
nand U11277 (N_11277,N_10552,N_10871);
xor U11278 (N_11278,N_10591,N_10857);
nand U11279 (N_11279,N_10741,N_10587);
nor U11280 (N_11280,N_10557,N_10706);
or U11281 (N_11281,N_10874,N_10592);
or U11282 (N_11282,N_10556,N_10944);
nand U11283 (N_11283,N_10787,N_10654);
and U11284 (N_11284,N_10581,N_10728);
and U11285 (N_11285,N_10587,N_10646);
and U11286 (N_11286,N_10841,N_10853);
or U11287 (N_11287,N_10864,N_10735);
or U11288 (N_11288,N_10919,N_10527);
nor U11289 (N_11289,N_10526,N_10681);
xnor U11290 (N_11290,N_10893,N_10589);
and U11291 (N_11291,N_10705,N_10815);
nor U11292 (N_11292,N_10787,N_10731);
and U11293 (N_11293,N_10960,N_10690);
nand U11294 (N_11294,N_10754,N_10918);
and U11295 (N_11295,N_10958,N_10678);
nor U11296 (N_11296,N_10825,N_10836);
xnor U11297 (N_11297,N_10567,N_10833);
nor U11298 (N_11298,N_10744,N_10747);
or U11299 (N_11299,N_10700,N_10955);
and U11300 (N_11300,N_10853,N_10707);
and U11301 (N_11301,N_10996,N_10512);
nor U11302 (N_11302,N_10556,N_10927);
nor U11303 (N_11303,N_10856,N_10716);
and U11304 (N_11304,N_10576,N_10691);
and U11305 (N_11305,N_10701,N_10969);
xor U11306 (N_11306,N_10654,N_10930);
or U11307 (N_11307,N_10544,N_10664);
nor U11308 (N_11308,N_10652,N_10921);
nor U11309 (N_11309,N_10915,N_10993);
nor U11310 (N_11310,N_10622,N_10751);
nand U11311 (N_11311,N_10629,N_10849);
or U11312 (N_11312,N_10772,N_10911);
and U11313 (N_11313,N_10954,N_10728);
and U11314 (N_11314,N_10766,N_10672);
or U11315 (N_11315,N_10594,N_10718);
and U11316 (N_11316,N_10633,N_10908);
nor U11317 (N_11317,N_10779,N_10808);
nand U11318 (N_11318,N_10949,N_10602);
or U11319 (N_11319,N_10571,N_10794);
and U11320 (N_11320,N_10695,N_10528);
nor U11321 (N_11321,N_10696,N_10752);
nor U11322 (N_11322,N_10535,N_10907);
and U11323 (N_11323,N_10553,N_10522);
or U11324 (N_11324,N_10761,N_10714);
nor U11325 (N_11325,N_10685,N_10694);
or U11326 (N_11326,N_10744,N_10561);
and U11327 (N_11327,N_10835,N_10974);
nor U11328 (N_11328,N_10756,N_10924);
or U11329 (N_11329,N_10898,N_10647);
nor U11330 (N_11330,N_10533,N_10761);
nor U11331 (N_11331,N_10889,N_10508);
or U11332 (N_11332,N_10987,N_10781);
and U11333 (N_11333,N_10535,N_10760);
or U11334 (N_11334,N_10939,N_10769);
and U11335 (N_11335,N_10954,N_10949);
nor U11336 (N_11336,N_10922,N_10752);
nor U11337 (N_11337,N_10966,N_10797);
and U11338 (N_11338,N_10964,N_10942);
or U11339 (N_11339,N_10698,N_10917);
and U11340 (N_11340,N_10556,N_10989);
nor U11341 (N_11341,N_10503,N_10929);
and U11342 (N_11342,N_10744,N_10880);
or U11343 (N_11343,N_10861,N_10705);
nor U11344 (N_11344,N_10642,N_10608);
and U11345 (N_11345,N_10785,N_10797);
nand U11346 (N_11346,N_10601,N_10682);
and U11347 (N_11347,N_10814,N_10914);
and U11348 (N_11348,N_10963,N_10689);
and U11349 (N_11349,N_10631,N_10590);
nand U11350 (N_11350,N_10933,N_10782);
nor U11351 (N_11351,N_10815,N_10816);
nand U11352 (N_11352,N_10794,N_10527);
or U11353 (N_11353,N_10693,N_10927);
and U11354 (N_11354,N_10546,N_10612);
nor U11355 (N_11355,N_10793,N_10770);
nand U11356 (N_11356,N_10685,N_10777);
or U11357 (N_11357,N_10688,N_10952);
xor U11358 (N_11358,N_10898,N_10825);
and U11359 (N_11359,N_10639,N_10804);
or U11360 (N_11360,N_10747,N_10716);
nand U11361 (N_11361,N_10897,N_10533);
and U11362 (N_11362,N_10601,N_10998);
or U11363 (N_11363,N_10973,N_10878);
nand U11364 (N_11364,N_10622,N_10533);
or U11365 (N_11365,N_10638,N_10598);
nand U11366 (N_11366,N_10757,N_10982);
nor U11367 (N_11367,N_10639,N_10595);
and U11368 (N_11368,N_10739,N_10783);
or U11369 (N_11369,N_10823,N_10875);
and U11370 (N_11370,N_10556,N_10743);
or U11371 (N_11371,N_10766,N_10659);
and U11372 (N_11372,N_10591,N_10992);
nand U11373 (N_11373,N_10589,N_10845);
nor U11374 (N_11374,N_10692,N_10657);
and U11375 (N_11375,N_10690,N_10605);
nand U11376 (N_11376,N_10970,N_10682);
nand U11377 (N_11377,N_10520,N_10573);
nor U11378 (N_11378,N_10606,N_10613);
and U11379 (N_11379,N_10729,N_10771);
and U11380 (N_11380,N_10594,N_10973);
and U11381 (N_11381,N_10925,N_10969);
and U11382 (N_11382,N_10676,N_10925);
nand U11383 (N_11383,N_10766,N_10836);
and U11384 (N_11384,N_10658,N_10916);
nor U11385 (N_11385,N_10808,N_10872);
nand U11386 (N_11386,N_10636,N_10666);
nor U11387 (N_11387,N_10806,N_10827);
or U11388 (N_11388,N_10844,N_10611);
nor U11389 (N_11389,N_10557,N_10764);
nor U11390 (N_11390,N_10764,N_10870);
or U11391 (N_11391,N_10856,N_10617);
xor U11392 (N_11392,N_10930,N_10811);
nand U11393 (N_11393,N_10570,N_10612);
nand U11394 (N_11394,N_10882,N_10739);
nor U11395 (N_11395,N_10985,N_10741);
and U11396 (N_11396,N_10659,N_10959);
nor U11397 (N_11397,N_10571,N_10705);
and U11398 (N_11398,N_10983,N_10795);
or U11399 (N_11399,N_10767,N_10938);
or U11400 (N_11400,N_10555,N_10769);
and U11401 (N_11401,N_10632,N_10520);
nor U11402 (N_11402,N_10797,N_10836);
nand U11403 (N_11403,N_10878,N_10775);
or U11404 (N_11404,N_10831,N_10823);
or U11405 (N_11405,N_10967,N_10903);
and U11406 (N_11406,N_10689,N_10827);
and U11407 (N_11407,N_10502,N_10761);
nand U11408 (N_11408,N_10683,N_10938);
nor U11409 (N_11409,N_10671,N_10526);
nand U11410 (N_11410,N_10849,N_10606);
or U11411 (N_11411,N_10815,N_10507);
or U11412 (N_11412,N_10730,N_10614);
and U11413 (N_11413,N_10657,N_10738);
and U11414 (N_11414,N_10701,N_10868);
xnor U11415 (N_11415,N_10711,N_10962);
nand U11416 (N_11416,N_10575,N_10758);
and U11417 (N_11417,N_10975,N_10767);
nand U11418 (N_11418,N_10619,N_10548);
nor U11419 (N_11419,N_10868,N_10561);
nand U11420 (N_11420,N_10805,N_10611);
and U11421 (N_11421,N_10958,N_10671);
nor U11422 (N_11422,N_10737,N_10717);
and U11423 (N_11423,N_10818,N_10842);
or U11424 (N_11424,N_10951,N_10504);
and U11425 (N_11425,N_10646,N_10669);
nor U11426 (N_11426,N_10739,N_10680);
nand U11427 (N_11427,N_10852,N_10815);
and U11428 (N_11428,N_10798,N_10698);
nand U11429 (N_11429,N_10509,N_10982);
nor U11430 (N_11430,N_10644,N_10741);
nor U11431 (N_11431,N_10553,N_10806);
nand U11432 (N_11432,N_10691,N_10831);
nor U11433 (N_11433,N_10840,N_10713);
nand U11434 (N_11434,N_10844,N_10538);
or U11435 (N_11435,N_10918,N_10996);
and U11436 (N_11436,N_10549,N_10575);
or U11437 (N_11437,N_10628,N_10546);
nand U11438 (N_11438,N_10935,N_10643);
nand U11439 (N_11439,N_10723,N_10896);
and U11440 (N_11440,N_10688,N_10964);
or U11441 (N_11441,N_10501,N_10644);
nor U11442 (N_11442,N_10968,N_10895);
and U11443 (N_11443,N_10979,N_10564);
and U11444 (N_11444,N_10742,N_10610);
and U11445 (N_11445,N_10932,N_10615);
nor U11446 (N_11446,N_10928,N_10781);
nand U11447 (N_11447,N_10830,N_10510);
and U11448 (N_11448,N_10720,N_10864);
nor U11449 (N_11449,N_10807,N_10766);
and U11450 (N_11450,N_10707,N_10504);
nor U11451 (N_11451,N_10863,N_10715);
nor U11452 (N_11452,N_10684,N_10747);
or U11453 (N_11453,N_10876,N_10568);
or U11454 (N_11454,N_10744,N_10679);
and U11455 (N_11455,N_10821,N_10949);
and U11456 (N_11456,N_10708,N_10760);
nand U11457 (N_11457,N_10975,N_10591);
and U11458 (N_11458,N_10731,N_10860);
nor U11459 (N_11459,N_10970,N_10759);
nor U11460 (N_11460,N_10547,N_10969);
nor U11461 (N_11461,N_10723,N_10616);
or U11462 (N_11462,N_10694,N_10990);
xnor U11463 (N_11463,N_10756,N_10845);
nor U11464 (N_11464,N_10750,N_10565);
nor U11465 (N_11465,N_10912,N_10867);
or U11466 (N_11466,N_10904,N_10676);
nand U11467 (N_11467,N_10679,N_10981);
nor U11468 (N_11468,N_10762,N_10928);
nand U11469 (N_11469,N_10685,N_10644);
or U11470 (N_11470,N_10728,N_10865);
and U11471 (N_11471,N_10546,N_10873);
nand U11472 (N_11472,N_10604,N_10658);
and U11473 (N_11473,N_10554,N_10803);
nand U11474 (N_11474,N_10647,N_10720);
or U11475 (N_11475,N_10691,N_10706);
nor U11476 (N_11476,N_10894,N_10886);
and U11477 (N_11477,N_10695,N_10779);
and U11478 (N_11478,N_10806,N_10841);
and U11479 (N_11479,N_10666,N_10953);
nand U11480 (N_11480,N_10931,N_10539);
nor U11481 (N_11481,N_10947,N_10604);
nor U11482 (N_11482,N_10961,N_10602);
and U11483 (N_11483,N_10558,N_10547);
or U11484 (N_11484,N_10985,N_10725);
nand U11485 (N_11485,N_10955,N_10593);
nor U11486 (N_11486,N_10819,N_10566);
nor U11487 (N_11487,N_10531,N_10657);
nor U11488 (N_11488,N_10723,N_10930);
or U11489 (N_11489,N_10868,N_10732);
nor U11490 (N_11490,N_10665,N_10524);
and U11491 (N_11491,N_10755,N_10717);
nand U11492 (N_11492,N_10845,N_10913);
nand U11493 (N_11493,N_10633,N_10695);
or U11494 (N_11494,N_10878,N_10842);
nand U11495 (N_11495,N_10693,N_10765);
nor U11496 (N_11496,N_10818,N_10883);
or U11497 (N_11497,N_10758,N_10768);
or U11498 (N_11498,N_10879,N_10949);
nor U11499 (N_11499,N_10902,N_10556);
nand U11500 (N_11500,N_11481,N_11254);
nand U11501 (N_11501,N_11213,N_11470);
or U11502 (N_11502,N_11471,N_11284);
or U11503 (N_11503,N_11177,N_11396);
and U11504 (N_11504,N_11272,N_11124);
nand U11505 (N_11505,N_11068,N_11455);
nor U11506 (N_11506,N_11050,N_11066);
and U11507 (N_11507,N_11046,N_11473);
nand U11508 (N_11508,N_11435,N_11200);
and U11509 (N_11509,N_11228,N_11147);
nand U11510 (N_11510,N_11163,N_11301);
or U11511 (N_11511,N_11460,N_11113);
nor U11512 (N_11512,N_11164,N_11057);
or U11513 (N_11513,N_11367,N_11197);
and U11514 (N_11514,N_11283,N_11490);
and U11515 (N_11515,N_11065,N_11154);
or U11516 (N_11516,N_11487,N_11445);
nor U11517 (N_11517,N_11220,N_11480);
and U11518 (N_11518,N_11231,N_11184);
nand U11519 (N_11519,N_11450,N_11031);
nor U11520 (N_11520,N_11288,N_11414);
nor U11521 (N_11521,N_11210,N_11499);
nor U11522 (N_11522,N_11214,N_11179);
or U11523 (N_11523,N_11035,N_11243);
and U11524 (N_11524,N_11497,N_11389);
nor U11525 (N_11525,N_11441,N_11298);
xor U11526 (N_11526,N_11010,N_11042);
and U11527 (N_11527,N_11053,N_11119);
or U11528 (N_11528,N_11356,N_11153);
nor U11529 (N_11529,N_11095,N_11238);
nor U11530 (N_11530,N_11223,N_11144);
nor U11531 (N_11531,N_11167,N_11364);
or U11532 (N_11532,N_11032,N_11036);
and U11533 (N_11533,N_11203,N_11334);
nand U11534 (N_11534,N_11131,N_11437);
nor U11535 (N_11535,N_11316,N_11017);
or U11536 (N_11536,N_11263,N_11368);
or U11537 (N_11537,N_11135,N_11067);
nand U11538 (N_11538,N_11279,N_11078);
or U11539 (N_11539,N_11215,N_11173);
nor U11540 (N_11540,N_11488,N_11280);
nor U11541 (N_11541,N_11307,N_11377);
nor U11542 (N_11542,N_11384,N_11161);
and U11543 (N_11543,N_11474,N_11002);
or U11544 (N_11544,N_11343,N_11321);
or U11545 (N_11545,N_11345,N_11338);
and U11546 (N_11546,N_11246,N_11048);
and U11547 (N_11547,N_11077,N_11388);
and U11548 (N_11548,N_11360,N_11402);
or U11549 (N_11549,N_11180,N_11101);
or U11550 (N_11550,N_11462,N_11310);
nand U11551 (N_11551,N_11258,N_11421);
and U11552 (N_11552,N_11052,N_11076);
nand U11553 (N_11553,N_11090,N_11433);
and U11554 (N_11554,N_11121,N_11329);
nor U11555 (N_11555,N_11404,N_11028);
nor U11556 (N_11556,N_11357,N_11439);
and U11557 (N_11557,N_11112,N_11019);
nand U11558 (N_11558,N_11132,N_11271);
nand U11559 (N_11559,N_11047,N_11390);
nor U11560 (N_11560,N_11103,N_11024);
or U11561 (N_11561,N_11296,N_11020);
and U11562 (N_11562,N_11072,N_11461);
or U11563 (N_11563,N_11039,N_11269);
nand U11564 (N_11564,N_11012,N_11413);
or U11565 (N_11565,N_11075,N_11295);
nor U11566 (N_11566,N_11256,N_11313);
and U11567 (N_11567,N_11138,N_11201);
and U11568 (N_11568,N_11085,N_11202);
or U11569 (N_11569,N_11382,N_11171);
nand U11570 (N_11570,N_11089,N_11374);
nand U11571 (N_11571,N_11080,N_11309);
and U11572 (N_11572,N_11142,N_11178);
and U11573 (N_11573,N_11299,N_11423);
nand U11574 (N_11574,N_11328,N_11183);
and U11575 (N_11575,N_11468,N_11411);
or U11576 (N_11576,N_11375,N_11217);
and U11577 (N_11577,N_11140,N_11422);
and U11578 (N_11578,N_11371,N_11442);
and U11579 (N_11579,N_11195,N_11436);
and U11580 (N_11580,N_11348,N_11070);
nand U11581 (N_11581,N_11176,N_11185);
or U11582 (N_11582,N_11380,N_11387);
or U11583 (N_11583,N_11270,N_11102);
or U11584 (N_11584,N_11196,N_11292);
nor U11585 (N_11585,N_11484,N_11114);
nand U11586 (N_11586,N_11449,N_11479);
nor U11587 (N_11587,N_11083,N_11105);
or U11588 (N_11588,N_11150,N_11312);
nor U11589 (N_11589,N_11034,N_11315);
nand U11590 (N_11590,N_11082,N_11230);
nor U11591 (N_11591,N_11236,N_11199);
or U11592 (N_11592,N_11063,N_11306);
nand U11593 (N_11593,N_11006,N_11240);
nor U11594 (N_11594,N_11126,N_11148);
or U11595 (N_11595,N_11420,N_11359);
and U11596 (N_11596,N_11018,N_11169);
nand U11597 (N_11597,N_11275,N_11198);
nand U11598 (N_11598,N_11000,N_11281);
nor U11599 (N_11599,N_11381,N_11257);
or U11600 (N_11600,N_11259,N_11416);
or U11601 (N_11601,N_11123,N_11033);
nand U11602 (N_11602,N_11385,N_11145);
or U11603 (N_11603,N_11454,N_11276);
nand U11604 (N_11604,N_11267,N_11327);
nand U11605 (N_11605,N_11443,N_11398);
nand U11606 (N_11606,N_11026,N_11096);
or U11607 (N_11607,N_11266,N_11193);
nand U11608 (N_11608,N_11426,N_11175);
nand U11609 (N_11609,N_11146,N_11486);
nor U11610 (N_11610,N_11318,N_11244);
and U11611 (N_11611,N_11137,N_11060);
nor U11612 (N_11612,N_11111,N_11250);
nand U11613 (N_11613,N_11346,N_11289);
and U11614 (N_11614,N_11110,N_11333);
nor U11615 (N_11615,N_11134,N_11467);
nor U11616 (N_11616,N_11049,N_11354);
or U11617 (N_11617,N_11409,N_11495);
nand U11618 (N_11618,N_11136,N_11094);
nor U11619 (N_11619,N_11181,N_11400);
and U11620 (N_11620,N_11425,N_11051);
or U11621 (N_11621,N_11030,N_11403);
nor U11622 (N_11622,N_11099,N_11417);
nor U11623 (N_11623,N_11438,N_11013);
nand U11624 (N_11624,N_11242,N_11247);
nor U11625 (N_11625,N_11363,N_11129);
and U11626 (N_11626,N_11005,N_11392);
nor U11627 (N_11627,N_11405,N_11317);
or U11628 (N_11628,N_11191,N_11383);
nor U11629 (N_11629,N_11340,N_11245);
and U11630 (N_11630,N_11274,N_11358);
or U11631 (N_11631,N_11457,N_11108);
nand U11632 (N_11632,N_11170,N_11172);
and U11633 (N_11633,N_11043,N_11353);
and U11634 (N_11634,N_11463,N_11476);
and U11635 (N_11635,N_11118,N_11311);
nand U11636 (N_11636,N_11187,N_11222);
or U11637 (N_11637,N_11361,N_11432);
nand U11638 (N_11638,N_11139,N_11003);
nor U11639 (N_11639,N_11478,N_11022);
nor U11640 (N_11640,N_11227,N_11492);
or U11641 (N_11641,N_11045,N_11379);
or U11642 (N_11642,N_11235,N_11498);
or U11643 (N_11643,N_11128,N_11475);
nand U11644 (N_11644,N_11219,N_11216);
nor U11645 (N_11645,N_11120,N_11302);
and U11646 (N_11646,N_11226,N_11429);
nand U11647 (N_11647,N_11428,N_11395);
nor U11648 (N_11648,N_11248,N_11483);
or U11649 (N_11649,N_11007,N_11001);
or U11650 (N_11650,N_11351,N_11155);
and U11651 (N_11651,N_11320,N_11464);
nor U11652 (N_11652,N_11332,N_11494);
nor U11653 (N_11653,N_11261,N_11015);
nor U11654 (N_11654,N_11293,N_11287);
nor U11655 (N_11655,N_11415,N_11237);
or U11656 (N_11656,N_11251,N_11418);
and U11657 (N_11657,N_11344,N_11190);
and U11658 (N_11658,N_11294,N_11037);
and U11659 (N_11659,N_11125,N_11448);
or U11660 (N_11660,N_11308,N_11365);
nand U11661 (N_11661,N_11084,N_11204);
nor U11662 (N_11662,N_11430,N_11286);
and U11663 (N_11663,N_11192,N_11188);
or U11664 (N_11664,N_11406,N_11054);
nor U11665 (N_11665,N_11249,N_11158);
and U11666 (N_11666,N_11152,N_11482);
nand U11667 (N_11667,N_11174,N_11116);
nor U11668 (N_11668,N_11011,N_11401);
nand U11669 (N_11669,N_11159,N_11014);
nor U11670 (N_11670,N_11291,N_11446);
nor U11671 (N_11671,N_11009,N_11427);
nor U11672 (N_11672,N_11156,N_11373);
or U11673 (N_11673,N_11331,N_11341);
nand U11674 (N_11674,N_11229,N_11335);
nor U11675 (N_11675,N_11025,N_11088);
and U11676 (N_11676,N_11452,N_11378);
or U11677 (N_11677,N_11064,N_11071);
or U11678 (N_11678,N_11297,N_11330);
nor U11679 (N_11679,N_11489,N_11008);
nand U11680 (N_11680,N_11056,N_11234);
nor U11681 (N_11681,N_11151,N_11255);
or U11682 (N_11682,N_11355,N_11456);
nor U11683 (N_11683,N_11491,N_11264);
or U11684 (N_11684,N_11342,N_11336);
and U11685 (N_11685,N_11469,N_11485);
or U11686 (N_11686,N_11087,N_11419);
xor U11687 (N_11687,N_11004,N_11493);
and U11688 (N_11688,N_11466,N_11207);
and U11689 (N_11689,N_11098,N_11376);
or U11690 (N_11690,N_11107,N_11440);
or U11691 (N_11691,N_11016,N_11027);
and U11692 (N_11692,N_11391,N_11038);
and U11693 (N_11693,N_11278,N_11073);
nor U11694 (N_11694,N_11305,N_11431);
nand U11695 (N_11695,N_11062,N_11205);
or U11696 (N_11696,N_11349,N_11300);
or U11697 (N_11697,N_11323,N_11339);
nor U11698 (N_11698,N_11189,N_11241);
nor U11699 (N_11699,N_11225,N_11211);
nand U11700 (N_11700,N_11044,N_11208);
nand U11701 (N_11701,N_11273,N_11397);
or U11702 (N_11702,N_11097,N_11117);
and U11703 (N_11703,N_11218,N_11304);
nand U11704 (N_11704,N_11386,N_11122);
and U11705 (N_11705,N_11130,N_11366);
nor U11706 (N_11706,N_11160,N_11347);
nand U11707 (N_11707,N_11074,N_11362);
nor U11708 (N_11708,N_11233,N_11412);
and U11709 (N_11709,N_11021,N_11399);
nor U11710 (N_11710,N_11212,N_11221);
nor U11711 (N_11711,N_11322,N_11168);
or U11712 (N_11712,N_11059,N_11092);
nor U11713 (N_11713,N_11314,N_11352);
nor U11714 (N_11714,N_11434,N_11194);
and U11715 (N_11715,N_11232,N_11079);
and U11716 (N_11716,N_11394,N_11209);
or U11717 (N_11717,N_11393,N_11093);
or U11718 (N_11718,N_11496,N_11069);
and U11719 (N_11719,N_11115,N_11285);
nor U11720 (N_11720,N_11447,N_11260);
nand U11721 (N_11721,N_11165,N_11133);
nor U11722 (N_11722,N_11477,N_11100);
and U11723 (N_11723,N_11141,N_11029);
or U11724 (N_11724,N_11091,N_11182);
or U11725 (N_11725,N_11350,N_11058);
or U11726 (N_11726,N_11407,N_11453);
or U11727 (N_11727,N_11410,N_11444);
nand U11728 (N_11728,N_11472,N_11324);
and U11729 (N_11729,N_11023,N_11265);
and U11730 (N_11730,N_11337,N_11061);
nand U11731 (N_11731,N_11239,N_11149);
nand U11732 (N_11732,N_11458,N_11040);
or U11733 (N_11733,N_11459,N_11081);
nor U11734 (N_11734,N_11451,N_11369);
nor U11735 (N_11735,N_11157,N_11325);
nand U11736 (N_11736,N_11055,N_11319);
and U11737 (N_11737,N_11206,N_11127);
nor U11738 (N_11738,N_11143,N_11372);
nor U11739 (N_11739,N_11408,N_11109);
nand U11740 (N_11740,N_11162,N_11253);
and U11741 (N_11741,N_11370,N_11290);
or U11742 (N_11742,N_11326,N_11303);
nor U11743 (N_11743,N_11262,N_11252);
or U11744 (N_11744,N_11282,N_11041);
nor U11745 (N_11745,N_11268,N_11104);
and U11746 (N_11746,N_11424,N_11166);
and U11747 (N_11747,N_11277,N_11224);
or U11748 (N_11748,N_11086,N_11106);
nor U11749 (N_11749,N_11186,N_11465);
nand U11750 (N_11750,N_11401,N_11249);
nand U11751 (N_11751,N_11113,N_11164);
nor U11752 (N_11752,N_11404,N_11197);
or U11753 (N_11753,N_11231,N_11261);
and U11754 (N_11754,N_11087,N_11499);
or U11755 (N_11755,N_11134,N_11108);
or U11756 (N_11756,N_11280,N_11261);
or U11757 (N_11757,N_11493,N_11355);
or U11758 (N_11758,N_11439,N_11140);
nor U11759 (N_11759,N_11310,N_11358);
and U11760 (N_11760,N_11168,N_11162);
and U11761 (N_11761,N_11020,N_11488);
nand U11762 (N_11762,N_11385,N_11260);
and U11763 (N_11763,N_11364,N_11464);
and U11764 (N_11764,N_11412,N_11175);
nor U11765 (N_11765,N_11261,N_11312);
nor U11766 (N_11766,N_11101,N_11446);
or U11767 (N_11767,N_11178,N_11064);
and U11768 (N_11768,N_11116,N_11318);
and U11769 (N_11769,N_11095,N_11303);
nand U11770 (N_11770,N_11401,N_11407);
nor U11771 (N_11771,N_11176,N_11106);
nor U11772 (N_11772,N_11116,N_11392);
nor U11773 (N_11773,N_11276,N_11275);
and U11774 (N_11774,N_11038,N_11313);
and U11775 (N_11775,N_11015,N_11042);
or U11776 (N_11776,N_11048,N_11149);
nor U11777 (N_11777,N_11478,N_11420);
and U11778 (N_11778,N_11335,N_11255);
nor U11779 (N_11779,N_11261,N_11197);
nand U11780 (N_11780,N_11163,N_11231);
nand U11781 (N_11781,N_11128,N_11193);
nor U11782 (N_11782,N_11380,N_11425);
nand U11783 (N_11783,N_11017,N_11015);
or U11784 (N_11784,N_11112,N_11225);
or U11785 (N_11785,N_11332,N_11156);
and U11786 (N_11786,N_11151,N_11478);
and U11787 (N_11787,N_11447,N_11058);
nor U11788 (N_11788,N_11310,N_11336);
nor U11789 (N_11789,N_11464,N_11192);
xor U11790 (N_11790,N_11391,N_11292);
nand U11791 (N_11791,N_11277,N_11244);
and U11792 (N_11792,N_11049,N_11248);
nor U11793 (N_11793,N_11380,N_11093);
or U11794 (N_11794,N_11201,N_11375);
xor U11795 (N_11795,N_11453,N_11192);
nand U11796 (N_11796,N_11104,N_11031);
nand U11797 (N_11797,N_11479,N_11174);
and U11798 (N_11798,N_11029,N_11498);
nor U11799 (N_11799,N_11113,N_11248);
nand U11800 (N_11800,N_11120,N_11283);
nor U11801 (N_11801,N_11381,N_11484);
nor U11802 (N_11802,N_11158,N_11271);
nand U11803 (N_11803,N_11282,N_11111);
or U11804 (N_11804,N_11366,N_11028);
nor U11805 (N_11805,N_11134,N_11000);
and U11806 (N_11806,N_11318,N_11016);
or U11807 (N_11807,N_11421,N_11396);
and U11808 (N_11808,N_11190,N_11254);
nand U11809 (N_11809,N_11304,N_11041);
or U11810 (N_11810,N_11146,N_11136);
and U11811 (N_11811,N_11243,N_11196);
or U11812 (N_11812,N_11308,N_11368);
xor U11813 (N_11813,N_11181,N_11051);
nand U11814 (N_11814,N_11058,N_11038);
and U11815 (N_11815,N_11010,N_11240);
or U11816 (N_11816,N_11198,N_11276);
or U11817 (N_11817,N_11029,N_11471);
nand U11818 (N_11818,N_11193,N_11425);
and U11819 (N_11819,N_11068,N_11294);
and U11820 (N_11820,N_11272,N_11248);
or U11821 (N_11821,N_11148,N_11263);
xnor U11822 (N_11822,N_11063,N_11212);
nor U11823 (N_11823,N_11175,N_11176);
nand U11824 (N_11824,N_11036,N_11272);
xnor U11825 (N_11825,N_11286,N_11400);
or U11826 (N_11826,N_11424,N_11234);
nor U11827 (N_11827,N_11240,N_11220);
nand U11828 (N_11828,N_11143,N_11462);
and U11829 (N_11829,N_11131,N_11046);
or U11830 (N_11830,N_11076,N_11379);
or U11831 (N_11831,N_11077,N_11454);
nor U11832 (N_11832,N_11400,N_11251);
or U11833 (N_11833,N_11323,N_11429);
nor U11834 (N_11834,N_11222,N_11410);
or U11835 (N_11835,N_11037,N_11167);
and U11836 (N_11836,N_11372,N_11353);
nor U11837 (N_11837,N_11084,N_11270);
or U11838 (N_11838,N_11057,N_11362);
or U11839 (N_11839,N_11352,N_11306);
and U11840 (N_11840,N_11144,N_11150);
nand U11841 (N_11841,N_11065,N_11377);
nand U11842 (N_11842,N_11463,N_11244);
and U11843 (N_11843,N_11133,N_11471);
nand U11844 (N_11844,N_11015,N_11401);
and U11845 (N_11845,N_11018,N_11042);
nor U11846 (N_11846,N_11247,N_11211);
nand U11847 (N_11847,N_11458,N_11186);
nor U11848 (N_11848,N_11061,N_11057);
nor U11849 (N_11849,N_11199,N_11224);
nor U11850 (N_11850,N_11443,N_11152);
nor U11851 (N_11851,N_11172,N_11048);
nor U11852 (N_11852,N_11467,N_11003);
or U11853 (N_11853,N_11239,N_11294);
and U11854 (N_11854,N_11090,N_11456);
and U11855 (N_11855,N_11352,N_11476);
nor U11856 (N_11856,N_11214,N_11303);
nand U11857 (N_11857,N_11009,N_11082);
nand U11858 (N_11858,N_11403,N_11080);
and U11859 (N_11859,N_11468,N_11093);
and U11860 (N_11860,N_11391,N_11453);
or U11861 (N_11861,N_11030,N_11117);
nand U11862 (N_11862,N_11288,N_11088);
nand U11863 (N_11863,N_11467,N_11220);
and U11864 (N_11864,N_11070,N_11134);
and U11865 (N_11865,N_11233,N_11406);
nand U11866 (N_11866,N_11329,N_11117);
nor U11867 (N_11867,N_11490,N_11023);
and U11868 (N_11868,N_11128,N_11186);
nor U11869 (N_11869,N_11227,N_11470);
and U11870 (N_11870,N_11428,N_11141);
nand U11871 (N_11871,N_11188,N_11459);
or U11872 (N_11872,N_11347,N_11148);
nor U11873 (N_11873,N_11330,N_11097);
or U11874 (N_11874,N_11069,N_11029);
nor U11875 (N_11875,N_11204,N_11491);
nor U11876 (N_11876,N_11182,N_11073);
nand U11877 (N_11877,N_11139,N_11408);
or U11878 (N_11878,N_11073,N_11259);
nor U11879 (N_11879,N_11169,N_11207);
nor U11880 (N_11880,N_11362,N_11163);
nor U11881 (N_11881,N_11363,N_11102);
nor U11882 (N_11882,N_11005,N_11377);
and U11883 (N_11883,N_11402,N_11267);
and U11884 (N_11884,N_11098,N_11002);
and U11885 (N_11885,N_11173,N_11075);
nand U11886 (N_11886,N_11085,N_11412);
and U11887 (N_11887,N_11363,N_11366);
and U11888 (N_11888,N_11073,N_11054);
nor U11889 (N_11889,N_11105,N_11205);
nand U11890 (N_11890,N_11483,N_11391);
and U11891 (N_11891,N_11143,N_11370);
nand U11892 (N_11892,N_11230,N_11197);
or U11893 (N_11893,N_11276,N_11475);
and U11894 (N_11894,N_11194,N_11276);
and U11895 (N_11895,N_11294,N_11127);
or U11896 (N_11896,N_11261,N_11446);
nand U11897 (N_11897,N_11273,N_11275);
or U11898 (N_11898,N_11291,N_11311);
and U11899 (N_11899,N_11280,N_11043);
or U11900 (N_11900,N_11142,N_11439);
nor U11901 (N_11901,N_11266,N_11105);
and U11902 (N_11902,N_11025,N_11490);
nand U11903 (N_11903,N_11411,N_11230);
nor U11904 (N_11904,N_11255,N_11285);
or U11905 (N_11905,N_11053,N_11242);
nand U11906 (N_11906,N_11122,N_11433);
or U11907 (N_11907,N_11104,N_11070);
or U11908 (N_11908,N_11110,N_11159);
nand U11909 (N_11909,N_11265,N_11341);
and U11910 (N_11910,N_11013,N_11252);
or U11911 (N_11911,N_11442,N_11476);
nor U11912 (N_11912,N_11300,N_11285);
xnor U11913 (N_11913,N_11271,N_11151);
nand U11914 (N_11914,N_11213,N_11029);
nor U11915 (N_11915,N_11190,N_11277);
nor U11916 (N_11916,N_11110,N_11028);
and U11917 (N_11917,N_11281,N_11386);
nand U11918 (N_11918,N_11119,N_11298);
nand U11919 (N_11919,N_11194,N_11316);
or U11920 (N_11920,N_11098,N_11470);
and U11921 (N_11921,N_11342,N_11289);
and U11922 (N_11922,N_11411,N_11252);
nand U11923 (N_11923,N_11032,N_11429);
nand U11924 (N_11924,N_11014,N_11090);
or U11925 (N_11925,N_11217,N_11316);
nor U11926 (N_11926,N_11110,N_11000);
nand U11927 (N_11927,N_11472,N_11145);
or U11928 (N_11928,N_11459,N_11477);
or U11929 (N_11929,N_11247,N_11303);
nand U11930 (N_11930,N_11445,N_11489);
nand U11931 (N_11931,N_11153,N_11043);
nand U11932 (N_11932,N_11426,N_11040);
nand U11933 (N_11933,N_11453,N_11255);
and U11934 (N_11934,N_11061,N_11035);
or U11935 (N_11935,N_11275,N_11107);
or U11936 (N_11936,N_11122,N_11155);
nand U11937 (N_11937,N_11234,N_11398);
nor U11938 (N_11938,N_11298,N_11215);
nor U11939 (N_11939,N_11108,N_11363);
and U11940 (N_11940,N_11115,N_11384);
or U11941 (N_11941,N_11142,N_11301);
xnor U11942 (N_11942,N_11283,N_11261);
and U11943 (N_11943,N_11029,N_11018);
or U11944 (N_11944,N_11295,N_11083);
nor U11945 (N_11945,N_11204,N_11163);
and U11946 (N_11946,N_11211,N_11446);
nand U11947 (N_11947,N_11146,N_11169);
nand U11948 (N_11948,N_11199,N_11125);
nand U11949 (N_11949,N_11132,N_11304);
or U11950 (N_11950,N_11463,N_11218);
nor U11951 (N_11951,N_11491,N_11374);
nor U11952 (N_11952,N_11181,N_11473);
nand U11953 (N_11953,N_11491,N_11220);
or U11954 (N_11954,N_11008,N_11268);
nand U11955 (N_11955,N_11186,N_11483);
or U11956 (N_11956,N_11118,N_11019);
nand U11957 (N_11957,N_11482,N_11246);
or U11958 (N_11958,N_11250,N_11411);
or U11959 (N_11959,N_11358,N_11437);
nor U11960 (N_11960,N_11093,N_11125);
and U11961 (N_11961,N_11172,N_11386);
and U11962 (N_11962,N_11320,N_11059);
nand U11963 (N_11963,N_11040,N_11060);
and U11964 (N_11964,N_11358,N_11409);
nor U11965 (N_11965,N_11081,N_11153);
or U11966 (N_11966,N_11285,N_11346);
nand U11967 (N_11967,N_11379,N_11156);
nor U11968 (N_11968,N_11046,N_11347);
nand U11969 (N_11969,N_11272,N_11093);
and U11970 (N_11970,N_11228,N_11041);
nand U11971 (N_11971,N_11024,N_11208);
or U11972 (N_11972,N_11298,N_11267);
nor U11973 (N_11973,N_11002,N_11074);
and U11974 (N_11974,N_11435,N_11483);
and U11975 (N_11975,N_11317,N_11346);
and U11976 (N_11976,N_11179,N_11277);
nor U11977 (N_11977,N_11000,N_11392);
nor U11978 (N_11978,N_11105,N_11390);
nand U11979 (N_11979,N_11146,N_11309);
nand U11980 (N_11980,N_11273,N_11142);
or U11981 (N_11981,N_11379,N_11251);
nor U11982 (N_11982,N_11012,N_11072);
nor U11983 (N_11983,N_11037,N_11373);
and U11984 (N_11984,N_11438,N_11432);
nand U11985 (N_11985,N_11433,N_11389);
and U11986 (N_11986,N_11090,N_11081);
or U11987 (N_11987,N_11008,N_11223);
or U11988 (N_11988,N_11224,N_11330);
nor U11989 (N_11989,N_11317,N_11219);
or U11990 (N_11990,N_11335,N_11325);
nand U11991 (N_11991,N_11115,N_11157);
and U11992 (N_11992,N_11021,N_11046);
and U11993 (N_11993,N_11069,N_11422);
nor U11994 (N_11994,N_11312,N_11344);
or U11995 (N_11995,N_11422,N_11164);
and U11996 (N_11996,N_11419,N_11071);
nor U11997 (N_11997,N_11356,N_11241);
nor U11998 (N_11998,N_11107,N_11265);
nor U11999 (N_11999,N_11259,N_11330);
and U12000 (N_12000,N_11952,N_11606);
and U12001 (N_12001,N_11964,N_11845);
nor U12002 (N_12002,N_11996,N_11945);
or U12003 (N_12003,N_11518,N_11679);
nor U12004 (N_12004,N_11803,N_11544);
and U12005 (N_12005,N_11513,N_11502);
or U12006 (N_12006,N_11724,N_11962);
and U12007 (N_12007,N_11727,N_11547);
nor U12008 (N_12008,N_11920,N_11593);
or U12009 (N_12009,N_11682,N_11626);
nand U12010 (N_12010,N_11979,N_11519);
and U12011 (N_12011,N_11919,N_11990);
nand U12012 (N_12012,N_11867,N_11526);
nor U12013 (N_12013,N_11981,N_11609);
nand U12014 (N_12014,N_11720,N_11521);
nor U12015 (N_12015,N_11717,N_11879);
and U12016 (N_12016,N_11758,N_11571);
or U12017 (N_12017,N_11785,N_11937);
xor U12018 (N_12018,N_11853,N_11987);
and U12019 (N_12019,N_11784,N_11949);
or U12020 (N_12020,N_11973,N_11725);
or U12021 (N_12021,N_11868,N_11883);
or U12022 (N_12022,N_11559,N_11833);
or U12023 (N_12023,N_11570,N_11870);
nand U12024 (N_12024,N_11903,N_11786);
nor U12025 (N_12025,N_11957,N_11540);
nand U12026 (N_12026,N_11711,N_11795);
or U12027 (N_12027,N_11931,N_11608);
nor U12028 (N_12028,N_11645,N_11652);
nand U12029 (N_12029,N_11646,N_11779);
nand U12030 (N_12030,N_11542,N_11885);
or U12031 (N_12031,N_11948,N_11848);
or U12032 (N_12032,N_11583,N_11707);
nand U12033 (N_12033,N_11986,N_11689);
nand U12034 (N_12034,N_11854,N_11842);
or U12035 (N_12035,N_11776,N_11680);
and U12036 (N_12036,N_11506,N_11802);
nand U12037 (N_12037,N_11837,N_11993);
nand U12038 (N_12038,N_11796,N_11860);
nor U12039 (N_12039,N_11702,N_11928);
and U12040 (N_12040,N_11751,N_11941);
and U12041 (N_12041,N_11624,N_11976);
or U12042 (N_12042,N_11539,N_11989);
nand U12043 (N_12043,N_11905,N_11761);
or U12044 (N_12044,N_11978,N_11953);
and U12045 (N_12045,N_11618,N_11810);
nor U12046 (N_12046,N_11923,N_11806);
nand U12047 (N_12047,N_11813,N_11824);
nor U12048 (N_12048,N_11632,N_11619);
xnor U12049 (N_12049,N_11822,N_11746);
nand U12050 (N_12050,N_11791,N_11798);
or U12051 (N_12051,N_11704,N_11734);
or U12052 (N_12052,N_11759,N_11744);
nand U12053 (N_12053,N_11561,N_11777);
or U12054 (N_12054,N_11788,N_11535);
nand U12055 (N_12055,N_11829,N_11718);
nand U12056 (N_12056,N_11590,N_11847);
nor U12057 (N_12057,N_11596,N_11657);
nand U12058 (N_12058,N_11631,N_11782);
or U12059 (N_12059,N_11850,N_11617);
and U12060 (N_12060,N_11697,N_11956);
nor U12061 (N_12061,N_11792,N_11588);
nand U12062 (N_12062,N_11816,N_11505);
nand U12063 (N_12063,N_11935,N_11886);
or U12064 (N_12064,N_11705,N_11563);
nand U12065 (N_12065,N_11528,N_11980);
nand U12066 (N_12066,N_11736,N_11669);
nor U12067 (N_12067,N_11753,N_11660);
or U12068 (N_12068,N_11844,N_11749);
or U12069 (N_12069,N_11983,N_11527);
or U12070 (N_12070,N_11898,N_11774);
nor U12071 (N_12071,N_11805,N_11698);
nand U12072 (N_12072,N_11656,N_11871);
and U12073 (N_12073,N_11650,N_11515);
and U12074 (N_12074,N_11579,N_11647);
and U12075 (N_12075,N_11819,N_11830);
and U12076 (N_12076,N_11875,N_11742);
nor U12077 (N_12077,N_11881,N_11991);
nor U12078 (N_12078,N_11926,N_11884);
and U12079 (N_12079,N_11825,N_11797);
nor U12080 (N_12080,N_11752,N_11536);
or U12081 (N_12081,N_11787,N_11548);
and U12082 (N_12082,N_11684,N_11582);
or U12083 (N_12083,N_11686,N_11770);
nand U12084 (N_12084,N_11740,N_11573);
nor U12085 (N_12085,N_11858,N_11633);
or U12086 (N_12086,N_11932,N_11700);
nand U12087 (N_12087,N_11627,N_11500);
nand U12088 (N_12088,N_11667,N_11814);
or U12089 (N_12089,N_11572,N_11567);
or U12090 (N_12090,N_11511,N_11872);
nor U12091 (N_12091,N_11866,N_11899);
nor U12092 (N_12092,N_11874,N_11721);
nor U12093 (N_12093,N_11600,N_11611);
nor U12094 (N_12094,N_11654,N_11509);
nor U12095 (N_12095,N_11781,N_11739);
and U12096 (N_12096,N_11900,N_11925);
or U12097 (N_12097,N_11581,N_11963);
nand U12098 (N_12098,N_11706,N_11818);
or U12099 (N_12099,N_11930,N_11914);
nor U12100 (N_12100,N_11726,N_11970);
nor U12101 (N_12101,N_11672,N_11901);
or U12102 (N_12102,N_11732,N_11807);
nand U12103 (N_12103,N_11675,N_11566);
nand U12104 (N_12104,N_11530,N_11940);
or U12105 (N_12105,N_11594,N_11944);
or U12106 (N_12106,N_11613,N_11630);
nand U12107 (N_12107,N_11938,N_11864);
or U12108 (N_12108,N_11694,N_11737);
nor U12109 (N_12109,N_11741,N_11557);
or U12110 (N_12110,N_11743,N_11550);
or U12111 (N_12111,N_11701,N_11893);
and U12112 (N_12112,N_11565,N_11889);
and U12113 (N_12113,N_11673,N_11934);
nor U12114 (N_12114,N_11936,N_11560);
or U12115 (N_12115,N_11768,N_11649);
nor U12116 (N_12116,N_11766,N_11662);
nor U12117 (N_12117,N_11773,N_11832);
nand U12118 (N_12118,N_11754,N_11841);
or U12119 (N_12119,N_11757,N_11895);
and U12120 (N_12120,N_11843,N_11562);
nand U12121 (N_12121,N_11554,N_11531);
and U12122 (N_12122,N_11681,N_11729);
nand U12123 (N_12123,N_11551,N_11569);
nor U12124 (N_12124,N_11549,N_11954);
nand U12125 (N_12125,N_11876,N_11541);
and U12126 (N_12126,N_11877,N_11644);
nand U12127 (N_12127,N_11762,N_11508);
and U12128 (N_12128,N_11998,N_11912);
and U12129 (N_12129,N_11719,N_11933);
nand U12130 (N_12130,N_11648,N_11894);
xnor U12131 (N_12131,N_11638,N_11851);
nor U12132 (N_12132,N_11887,N_11747);
and U12133 (N_12133,N_11951,N_11728);
or U12134 (N_12134,N_11826,N_11537);
nor U12135 (N_12135,N_11852,N_11605);
nand U12136 (N_12136,N_11615,N_11603);
or U12137 (N_12137,N_11915,N_11985);
nand U12138 (N_12138,N_11659,N_11677);
nand U12139 (N_12139,N_11780,N_11827);
and U12140 (N_12140,N_11969,N_11817);
nor U12141 (N_12141,N_11862,N_11775);
or U12142 (N_12142,N_11623,N_11636);
or U12143 (N_12143,N_11589,N_11815);
or U12144 (N_12144,N_11799,N_11713);
nand U12145 (N_12145,N_11664,N_11688);
nand U12146 (N_12146,N_11909,N_11918);
or U12147 (N_12147,N_11663,N_11863);
nand U12148 (N_12148,N_11599,N_11553);
nor U12149 (N_12149,N_11997,N_11999);
nor U12150 (N_12150,N_11873,N_11601);
or U12151 (N_12151,N_11735,N_11516);
nor U12152 (N_12152,N_11577,N_11564);
or U12153 (N_12153,N_11512,N_11917);
and U12154 (N_12154,N_11856,N_11738);
nand U12155 (N_12155,N_11576,N_11913);
nor U12156 (N_12156,N_11592,N_11622);
nor U12157 (N_12157,N_11756,N_11586);
nand U12158 (N_12158,N_11835,N_11836);
or U12159 (N_12159,N_11767,N_11961);
nor U12160 (N_12160,N_11965,N_11959);
or U12161 (N_12161,N_11598,N_11823);
nor U12162 (N_12162,N_11927,N_11995);
nor U12163 (N_12163,N_11533,N_11882);
and U12164 (N_12164,N_11520,N_11828);
or U12165 (N_12165,N_11809,N_11974);
nor U12166 (N_12166,N_11878,N_11730);
or U12167 (N_12167,N_11699,N_11703);
and U12168 (N_12168,N_11733,N_11676);
nor U12169 (N_12169,N_11545,N_11693);
nor U12170 (N_12170,N_11789,N_11574);
nand U12171 (N_12171,N_11865,N_11943);
or U12172 (N_12172,N_11950,N_11800);
nand U12173 (N_12173,N_11670,N_11678);
and U12174 (N_12174,N_11532,N_11665);
and U12175 (N_12175,N_11831,N_11745);
nand U12176 (N_12176,N_11838,N_11857);
nand U12177 (N_12177,N_11640,N_11604);
nor U12178 (N_12178,N_11910,N_11628);
nor U12179 (N_12179,N_11639,N_11992);
nor U12180 (N_12180,N_11523,N_11510);
nor U12181 (N_12181,N_11890,N_11546);
nor U12182 (N_12182,N_11760,N_11616);
nand U12183 (N_12183,N_11793,N_11655);
nor U12184 (N_12184,N_11514,N_11661);
or U12185 (N_12185,N_11902,N_11960);
nand U12186 (N_12186,N_11501,N_11610);
or U12187 (N_12187,N_11929,N_11924);
nor U12188 (N_12188,N_11790,N_11524);
nor U12189 (N_12189,N_11804,N_11896);
and U12190 (N_12190,N_11911,N_11692);
nand U12191 (N_12191,N_11888,N_11556);
and U12192 (N_12192,N_11955,N_11812);
nor U12193 (N_12193,N_11916,N_11723);
or U12194 (N_12194,N_11748,N_11968);
or U12195 (N_12195,N_11771,N_11614);
and U12196 (N_12196,N_11861,N_11620);
or U12197 (N_12197,N_11869,N_11907);
nand U12198 (N_12198,N_11722,N_11716);
and U12199 (N_12199,N_11769,N_11971);
nand U12200 (N_12200,N_11683,N_11584);
nand U12201 (N_12201,N_11685,N_11690);
or U12202 (N_12202,N_11503,N_11585);
nand U12203 (N_12203,N_11834,N_11947);
and U12204 (N_12204,N_11607,N_11906);
nor U12205 (N_12205,N_11658,N_11772);
nor U12206 (N_12206,N_11921,N_11859);
and U12207 (N_12207,N_11525,N_11811);
or U12208 (N_12208,N_11765,N_11783);
and U12209 (N_12209,N_11522,N_11691);
nor U12210 (N_12210,N_11982,N_11763);
or U12211 (N_12211,N_11849,N_11840);
nand U12212 (N_12212,N_11755,N_11629);
and U12213 (N_12213,N_11750,N_11731);
nand U12214 (N_12214,N_11634,N_11666);
nor U12215 (N_12215,N_11904,N_11575);
and U12216 (N_12216,N_11892,N_11696);
or U12217 (N_12217,N_11714,N_11687);
nor U12218 (N_12218,N_11621,N_11625);
nand U12219 (N_12219,N_11977,N_11587);
or U12220 (N_12220,N_11942,N_11695);
or U12221 (N_12221,N_11504,N_11591);
and U12222 (N_12222,N_11653,N_11674);
and U12223 (N_12223,N_11908,N_11642);
and U12224 (N_12224,N_11641,N_11715);
or U12225 (N_12225,N_11651,N_11988);
and U12226 (N_12226,N_11558,N_11820);
nand U12227 (N_12227,N_11946,N_11612);
nand U12228 (N_12228,N_11821,N_11764);
nor U12229 (N_12229,N_11994,N_11708);
nand U12230 (N_12230,N_11543,N_11635);
nand U12231 (N_12231,N_11846,N_11984);
and U12232 (N_12232,N_11808,N_11709);
nand U12233 (N_12233,N_11897,N_11517);
or U12234 (N_12234,N_11891,N_11637);
or U12235 (N_12235,N_11529,N_11643);
xnor U12236 (N_12236,N_11880,N_11839);
and U12237 (N_12237,N_11671,N_11778);
or U12238 (N_12238,N_11939,N_11972);
nand U12239 (N_12239,N_11552,N_11507);
or U12240 (N_12240,N_11801,N_11922);
nand U12241 (N_12241,N_11712,N_11534);
nor U12242 (N_12242,N_11958,N_11580);
nand U12243 (N_12243,N_11568,N_11602);
nor U12244 (N_12244,N_11966,N_11595);
xnor U12245 (N_12245,N_11668,N_11975);
nand U12246 (N_12246,N_11855,N_11597);
and U12247 (N_12247,N_11794,N_11538);
and U12248 (N_12248,N_11578,N_11555);
and U12249 (N_12249,N_11967,N_11710);
nand U12250 (N_12250,N_11811,N_11813);
nor U12251 (N_12251,N_11650,N_11525);
nor U12252 (N_12252,N_11933,N_11914);
and U12253 (N_12253,N_11784,N_11905);
nor U12254 (N_12254,N_11693,N_11993);
nor U12255 (N_12255,N_11681,N_11704);
nor U12256 (N_12256,N_11832,N_11970);
or U12257 (N_12257,N_11922,N_11684);
or U12258 (N_12258,N_11940,N_11528);
nand U12259 (N_12259,N_11666,N_11697);
nand U12260 (N_12260,N_11874,N_11915);
nand U12261 (N_12261,N_11914,N_11903);
and U12262 (N_12262,N_11972,N_11960);
nor U12263 (N_12263,N_11785,N_11645);
xnor U12264 (N_12264,N_11792,N_11836);
nand U12265 (N_12265,N_11958,N_11980);
or U12266 (N_12266,N_11550,N_11672);
and U12267 (N_12267,N_11964,N_11812);
and U12268 (N_12268,N_11669,N_11564);
nand U12269 (N_12269,N_11989,N_11692);
nand U12270 (N_12270,N_11559,N_11509);
and U12271 (N_12271,N_11670,N_11880);
xnor U12272 (N_12272,N_11746,N_11889);
nand U12273 (N_12273,N_11950,N_11742);
and U12274 (N_12274,N_11708,N_11851);
nor U12275 (N_12275,N_11838,N_11780);
or U12276 (N_12276,N_11749,N_11557);
nor U12277 (N_12277,N_11552,N_11765);
nor U12278 (N_12278,N_11527,N_11873);
or U12279 (N_12279,N_11956,N_11768);
and U12280 (N_12280,N_11713,N_11686);
nor U12281 (N_12281,N_11964,N_11584);
nor U12282 (N_12282,N_11886,N_11746);
or U12283 (N_12283,N_11605,N_11700);
nand U12284 (N_12284,N_11602,N_11929);
and U12285 (N_12285,N_11569,N_11600);
or U12286 (N_12286,N_11696,N_11582);
nor U12287 (N_12287,N_11945,N_11763);
and U12288 (N_12288,N_11969,N_11874);
or U12289 (N_12289,N_11748,N_11742);
nand U12290 (N_12290,N_11767,N_11903);
and U12291 (N_12291,N_11956,N_11707);
or U12292 (N_12292,N_11960,N_11667);
nor U12293 (N_12293,N_11857,N_11940);
nand U12294 (N_12294,N_11828,N_11981);
or U12295 (N_12295,N_11589,N_11727);
and U12296 (N_12296,N_11570,N_11960);
nand U12297 (N_12297,N_11668,N_11550);
nor U12298 (N_12298,N_11603,N_11695);
or U12299 (N_12299,N_11538,N_11758);
nand U12300 (N_12300,N_11528,N_11822);
and U12301 (N_12301,N_11748,N_11673);
nand U12302 (N_12302,N_11982,N_11877);
or U12303 (N_12303,N_11645,N_11561);
or U12304 (N_12304,N_11612,N_11790);
nand U12305 (N_12305,N_11834,N_11823);
nor U12306 (N_12306,N_11974,N_11784);
nor U12307 (N_12307,N_11777,N_11952);
xor U12308 (N_12308,N_11846,N_11696);
and U12309 (N_12309,N_11603,N_11659);
and U12310 (N_12310,N_11942,N_11951);
nor U12311 (N_12311,N_11690,N_11649);
and U12312 (N_12312,N_11738,N_11916);
nor U12313 (N_12313,N_11926,N_11624);
or U12314 (N_12314,N_11760,N_11652);
nor U12315 (N_12315,N_11607,N_11702);
nand U12316 (N_12316,N_11560,N_11932);
and U12317 (N_12317,N_11926,N_11801);
and U12318 (N_12318,N_11568,N_11678);
and U12319 (N_12319,N_11519,N_11969);
nor U12320 (N_12320,N_11898,N_11638);
and U12321 (N_12321,N_11507,N_11556);
or U12322 (N_12322,N_11851,N_11902);
nand U12323 (N_12323,N_11960,N_11980);
nor U12324 (N_12324,N_11823,N_11738);
or U12325 (N_12325,N_11711,N_11713);
nor U12326 (N_12326,N_11890,N_11658);
and U12327 (N_12327,N_11793,N_11916);
nand U12328 (N_12328,N_11576,N_11535);
nor U12329 (N_12329,N_11903,N_11657);
and U12330 (N_12330,N_11592,N_11962);
and U12331 (N_12331,N_11656,N_11897);
nor U12332 (N_12332,N_11709,N_11898);
nand U12333 (N_12333,N_11711,N_11847);
nor U12334 (N_12334,N_11944,N_11669);
or U12335 (N_12335,N_11677,N_11554);
nor U12336 (N_12336,N_11567,N_11900);
nor U12337 (N_12337,N_11861,N_11533);
nand U12338 (N_12338,N_11598,N_11521);
and U12339 (N_12339,N_11908,N_11771);
nor U12340 (N_12340,N_11618,N_11995);
nand U12341 (N_12341,N_11598,N_11535);
or U12342 (N_12342,N_11906,N_11839);
nor U12343 (N_12343,N_11578,N_11876);
nand U12344 (N_12344,N_11913,N_11653);
nand U12345 (N_12345,N_11582,N_11562);
nand U12346 (N_12346,N_11578,N_11791);
xor U12347 (N_12347,N_11759,N_11588);
nor U12348 (N_12348,N_11955,N_11735);
nor U12349 (N_12349,N_11684,N_11744);
and U12350 (N_12350,N_11881,N_11858);
nand U12351 (N_12351,N_11658,N_11589);
nand U12352 (N_12352,N_11750,N_11657);
and U12353 (N_12353,N_11978,N_11581);
or U12354 (N_12354,N_11770,N_11805);
and U12355 (N_12355,N_11716,N_11972);
and U12356 (N_12356,N_11590,N_11539);
or U12357 (N_12357,N_11692,N_11567);
nor U12358 (N_12358,N_11971,N_11864);
or U12359 (N_12359,N_11803,N_11859);
nor U12360 (N_12360,N_11970,N_11848);
nand U12361 (N_12361,N_11502,N_11849);
or U12362 (N_12362,N_11886,N_11576);
and U12363 (N_12363,N_11824,N_11938);
and U12364 (N_12364,N_11535,N_11980);
nand U12365 (N_12365,N_11694,N_11564);
nand U12366 (N_12366,N_11929,N_11940);
nor U12367 (N_12367,N_11678,N_11754);
and U12368 (N_12368,N_11635,N_11907);
nand U12369 (N_12369,N_11964,N_11778);
nand U12370 (N_12370,N_11995,N_11605);
or U12371 (N_12371,N_11511,N_11575);
or U12372 (N_12372,N_11974,N_11858);
or U12373 (N_12373,N_11866,N_11512);
or U12374 (N_12374,N_11900,N_11858);
nor U12375 (N_12375,N_11971,N_11798);
nand U12376 (N_12376,N_11876,N_11738);
and U12377 (N_12377,N_11946,N_11900);
nor U12378 (N_12378,N_11849,N_11531);
nor U12379 (N_12379,N_11752,N_11887);
and U12380 (N_12380,N_11938,N_11754);
nor U12381 (N_12381,N_11985,N_11972);
nand U12382 (N_12382,N_11813,N_11685);
and U12383 (N_12383,N_11693,N_11666);
or U12384 (N_12384,N_11660,N_11902);
and U12385 (N_12385,N_11853,N_11664);
nor U12386 (N_12386,N_11918,N_11533);
and U12387 (N_12387,N_11877,N_11711);
or U12388 (N_12388,N_11598,N_11862);
nand U12389 (N_12389,N_11518,N_11814);
nor U12390 (N_12390,N_11848,N_11647);
and U12391 (N_12391,N_11554,N_11969);
or U12392 (N_12392,N_11616,N_11710);
nor U12393 (N_12393,N_11523,N_11552);
or U12394 (N_12394,N_11708,N_11559);
nor U12395 (N_12395,N_11763,N_11558);
or U12396 (N_12396,N_11757,N_11952);
nand U12397 (N_12397,N_11533,N_11679);
and U12398 (N_12398,N_11927,N_11924);
nor U12399 (N_12399,N_11673,N_11801);
and U12400 (N_12400,N_11762,N_11577);
or U12401 (N_12401,N_11963,N_11628);
nand U12402 (N_12402,N_11541,N_11957);
nor U12403 (N_12403,N_11707,N_11738);
nor U12404 (N_12404,N_11595,N_11797);
nand U12405 (N_12405,N_11531,N_11986);
nand U12406 (N_12406,N_11810,N_11995);
or U12407 (N_12407,N_11620,N_11770);
nor U12408 (N_12408,N_11737,N_11596);
nand U12409 (N_12409,N_11971,N_11744);
nand U12410 (N_12410,N_11810,N_11723);
or U12411 (N_12411,N_11625,N_11651);
nand U12412 (N_12412,N_11527,N_11971);
and U12413 (N_12413,N_11883,N_11762);
and U12414 (N_12414,N_11653,N_11815);
or U12415 (N_12415,N_11656,N_11914);
or U12416 (N_12416,N_11718,N_11741);
and U12417 (N_12417,N_11705,N_11606);
nand U12418 (N_12418,N_11869,N_11598);
nor U12419 (N_12419,N_11739,N_11890);
nand U12420 (N_12420,N_11623,N_11872);
nand U12421 (N_12421,N_11675,N_11841);
nand U12422 (N_12422,N_11817,N_11763);
nor U12423 (N_12423,N_11563,N_11988);
or U12424 (N_12424,N_11765,N_11566);
nand U12425 (N_12425,N_11881,N_11567);
nor U12426 (N_12426,N_11639,N_11598);
nor U12427 (N_12427,N_11617,N_11831);
or U12428 (N_12428,N_11538,N_11760);
and U12429 (N_12429,N_11884,N_11832);
nand U12430 (N_12430,N_11790,N_11706);
or U12431 (N_12431,N_11603,N_11663);
or U12432 (N_12432,N_11721,N_11704);
xor U12433 (N_12433,N_11611,N_11661);
nor U12434 (N_12434,N_11680,N_11932);
and U12435 (N_12435,N_11854,N_11669);
nand U12436 (N_12436,N_11608,N_11653);
or U12437 (N_12437,N_11665,N_11879);
nor U12438 (N_12438,N_11669,N_11623);
or U12439 (N_12439,N_11858,N_11527);
and U12440 (N_12440,N_11953,N_11579);
and U12441 (N_12441,N_11767,N_11783);
nand U12442 (N_12442,N_11846,N_11742);
or U12443 (N_12443,N_11788,N_11514);
or U12444 (N_12444,N_11856,N_11811);
nand U12445 (N_12445,N_11796,N_11565);
and U12446 (N_12446,N_11559,N_11788);
or U12447 (N_12447,N_11589,N_11841);
and U12448 (N_12448,N_11503,N_11889);
nor U12449 (N_12449,N_11976,N_11625);
or U12450 (N_12450,N_11804,N_11905);
nand U12451 (N_12451,N_11723,N_11777);
nor U12452 (N_12452,N_11658,N_11967);
nand U12453 (N_12453,N_11699,N_11644);
or U12454 (N_12454,N_11847,N_11812);
and U12455 (N_12455,N_11697,N_11800);
nor U12456 (N_12456,N_11845,N_11836);
nor U12457 (N_12457,N_11742,N_11802);
or U12458 (N_12458,N_11616,N_11530);
nand U12459 (N_12459,N_11718,N_11742);
nand U12460 (N_12460,N_11979,N_11589);
nor U12461 (N_12461,N_11801,N_11797);
or U12462 (N_12462,N_11802,N_11719);
or U12463 (N_12463,N_11817,N_11676);
and U12464 (N_12464,N_11730,N_11796);
nand U12465 (N_12465,N_11752,N_11529);
and U12466 (N_12466,N_11714,N_11804);
or U12467 (N_12467,N_11517,N_11745);
or U12468 (N_12468,N_11799,N_11736);
or U12469 (N_12469,N_11707,N_11853);
nor U12470 (N_12470,N_11508,N_11631);
or U12471 (N_12471,N_11804,N_11589);
and U12472 (N_12472,N_11797,N_11575);
or U12473 (N_12473,N_11650,N_11558);
nor U12474 (N_12474,N_11583,N_11796);
or U12475 (N_12475,N_11535,N_11853);
or U12476 (N_12476,N_11908,N_11860);
and U12477 (N_12477,N_11756,N_11685);
or U12478 (N_12478,N_11536,N_11614);
nor U12479 (N_12479,N_11863,N_11534);
and U12480 (N_12480,N_11829,N_11621);
or U12481 (N_12481,N_11774,N_11716);
or U12482 (N_12482,N_11907,N_11804);
nand U12483 (N_12483,N_11725,N_11894);
and U12484 (N_12484,N_11639,N_11926);
or U12485 (N_12485,N_11516,N_11615);
or U12486 (N_12486,N_11727,N_11840);
or U12487 (N_12487,N_11541,N_11935);
and U12488 (N_12488,N_11909,N_11931);
nor U12489 (N_12489,N_11897,N_11781);
and U12490 (N_12490,N_11673,N_11852);
nor U12491 (N_12491,N_11591,N_11821);
nor U12492 (N_12492,N_11891,N_11574);
nor U12493 (N_12493,N_11501,N_11733);
or U12494 (N_12494,N_11550,N_11661);
nand U12495 (N_12495,N_11681,N_11742);
nor U12496 (N_12496,N_11598,N_11534);
or U12497 (N_12497,N_11973,N_11665);
or U12498 (N_12498,N_11756,N_11721);
and U12499 (N_12499,N_11625,N_11969);
and U12500 (N_12500,N_12229,N_12436);
or U12501 (N_12501,N_12126,N_12145);
nor U12502 (N_12502,N_12369,N_12475);
nor U12503 (N_12503,N_12357,N_12127);
and U12504 (N_12504,N_12134,N_12457);
and U12505 (N_12505,N_12249,N_12302);
or U12506 (N_12506,N_12059,N_12190);
nand U12507 (N_12507,N_12052,N_12409);
nand U12508 (N_12508,N_12375,N_12431);
and U12509 (N_12509,N_12020,N_12403);
and U12510 (N_12510,N_12480,N_12494);
or U12511 (N_12511,N_12049,N_12407);
xnor U12512 (N_12512,N_12439,N_12138);
and U12513 (N_12513,N_12488,N_12055);
nand U12514 (N_12514,N_12043,N_12322);
or U12515 (N_12515,N_12114,N_12191);
and U12516 (N_12516,N_12474,N_12282);
nand U12517 (N_12517,N_12413,N_12180);
nand U12518 (N_12518,N_12223,N_12228);
nand U12519 (N_12519,N_12258,N_12365);
and U12520 (N_12520,N_12017,N_12124);
or U12521 (N_12521,N_12288,N_12495);
xnor U12522 (N_12522,N_12356,N_12433);
or U12523 (N_12523,N_12351,N_12056);
nor U12524 (N_12524,N_12364,N_12455);
or U12525 (N_12525,N_12283,N_12247);
or U12526 (N_12526,N_12107,N_12158);
nor U12527 (N_12527,N_12081,N_12168);
or U12528 (N_12528,N_12421,N_12316);
nor U12529 (N_12529,N_12267,N_12401);
nor U12530 (N_12530,N_12404,N_12149);
or U12531 (N_12531,N_12153,N_12281);
and U12532 (N_12532,N_12370,N_12230);
or U12533 (N_12533,N_12254,N_12184);
or U12534 (N_12534,N_12027,N_12262);
or U12535 (N_12535,N_12006,N_12132);
and U12536 (N_12536,N_12263,N_12019);
or U12537 (N_12537,N_12358,N_12074);
nand U12538 (N_12538,N_12306,N_12154);
and U12539 (N_12539,N_12050,N_12186);
and U12540 (N_12540,N_12447,N_12312);
nor U12541 (N_12541,N_12151,N_12148);
and U12542 (N_12542,N_12402,N_12164);
or U12543 (N_12543,N_12057,N_12422);
nand U12544 (N_12544,N_12325,N_12389);
or U12545 (N_12545,N_12060,N_12156);
nand U12546 (N_12546,N_12441,N_12205);
and U12547 (N_12547,N_12317,N_12061);
nand U12548 (N_12548,N_12011,N_12384);
or U12549 (N_12549,N_12347,N_12286);
or U12550 (N_12550,N_12348,N_12147);
nand U12551 (N_12551,N_12159,N_12106);
nand U12552 (N_12552,N_12329,N_12116);
or U12553 (N_12553,N_12160,N_12387);
nand U12554 (N_12554,N_12386,N_12220);
and U12555 (N_12555,N_12424,N_12453);
nor U12556 (N_12556,N_12451,N_12082);
nand U12557 (N_12557,N_12385,N_12236);
nand U12558 (N_12558,N_12174,N_12465);
nand U12559 (N_12559,N_12008,N_12244);
and U12560 (N_12560,N_12496,N_12499);
or U12561 (N_12561,N_12349,N_12371);
nand U12562 (N_12562,N_12115,N_12048);
or U12563 (N_12563,N_12498,N_12266);
nor U12564 (N_12564,N_12064,N_12095);
nand U12565 (N_12565,N_12437,N_12289);
nor U12566 (N_12566,N_12084,N_12233);
nor U12567 (N_12567,N_12171,N_12333);
and U12568 (N_12568,N_12343,N_12121);
and U12569 (N_12569,N_12467,N_12217);
or U12570 (N_12570,N_12321,N_12260);
and U12571 (N_12571,N_12368,N_12099);
and U12572 (N_12572,N_12486,N_12328);
and U12573 (N_12573,N_12014,N_12037);
nor U12574 (N_12574,N_12477,N_12080);
nor U12575 (N_12575,N_12314,N_12198);
nor U12576 (N_12576,N_12323,N_12462);
xnor U12577 (N_12577,N_12133,N_12226);
nand U12578 (N_12578,N_12419,N_12416);
nand U12579 (N_12579,N_12259,N_12243);
nand U12580 (N_12580,N_12461,N_12327);
and U12581 (N_12581,N_12192,N_12309);
or U12582 (N_12582,N_12468,N_12382);
nand U12583 (N_12583,N_12010,N_12346);
or U12584 (N_12584,N_12079,N_12204);
nor U12585 (N_12585,N_12277,N_12446);
nand U12586 (N_12586,N_12025,N_12235);
nor U12587 (N_12587,N_12030,N_12458);
and U12588 (N_12588,N_12435,N_12090);
and U12589 (N_12589,N_12108,N_12278);
or U12590 (N_12590,N_12303,N_12058);
or U12591 (N_12591,N_12352,N_12215);
or U12592 (N_12592,N_12097,N_12344);
and U12593 (N_12593,N_12428,N_12113);
and U12594 (N_12594,N_12213,N_12004);
nor U12595 (N_12595,N_12367,N_12045);
and U12596 (N_12596,N_12181,N_12062);
and U12597 (N_12597,N_12152,N_12194);
nor U12598 (N_12598,N_12381,N_12342);
and U12599 (N_12599,N_12285,N_12473);
xor U12600 (N_12600,N_12326,N_12391);
xnor U12601 (N_12601,N_12227,N_12340);
nor U12602 (N_12602,N_12219,N_12373);
nand U12603 (N_12603,N_12432,N_12290);
nor U12604 (N_12604,N_12456,N_12112);
and U12605 (N_12605,N_12253,N_12234);
nand U12606 (N_12606,N_12143,N_12430);
or U12607 (N_12607,N_12040,N_12165);
nor U12608 (N_12608,N_12176,N_12144);
and U12609 (N_12609,N_12245,N_12221);
and U12610 (N_12610,N_12140,N_12295);
nor U12611 (N_12611,N_12031,N_12076);
and U12612 (N_12612,N_12086,N_12197);
or U12613 (N_12613,N_12257,N_12293);
or U12614 (N_12614,N_12232,N_12360);
nand U12615 (N_12615,N_12066,N_12212);
or U12616 (N_12616,N_12398,N_12395);
or U12617 (N_12617,N_12318,N_12070);
and U12618 (N_12618,N_12202,N_12497);
and U12619 (N_12619,N_12311,N_12482);
nor U12620 (N_12620,N_12101,N_12069);
nand U12621 (N_12621,N_12361,N_12033);
and U12622 (N_12622,N_12463,N_12334);
nand U12623 (N_12623,N_12359,N_12015);
or U12624 (N_12624,N_12122,N_12300);
nand U12625 (N_12625,N_12196,N_12117);
nand U12626 (N_12626,N_12085,N_12023);
nand U12627 (N_12627,N_12125,N_12479);
and U12628 (N_12628,N_12175,N_12423);
or U12629 (N_12629,N_12355,N_12250);
and U12630 (N_12630,N_12071,N_12362);
nand U12631 (N_12631,N_12018,N_12150);
and U12632 (N_12632,N_12083,N_12053);
and U12633 (N_12633,N_12310,N_12274);
nor U12634 (N_12634,N_12272,N_12450);
nand U12635 (N_12635,N_12073,N_12276);
nor U12636 (N_12636,N_12142,N_12354);
nor U12637 (N_12637,N_12096,N_12378);
nor U12638 (N_12638,N_12054,N_12393);
or U12639 (N_12639,N_12039,N_12291);
or U12640 (N_12640,N_12067,N_12214);
nor U12641 (N_12641,N_12490,N_12324);
or U12642 (N_12642,N_12211,N_12105);
and U12643 (N_12643,N_12100,N_12162);
nand U12644 (N_12644,N_12021,N_12392);
nor U12645 (N_12645,N_12047,N_12454);
and U12646 (N_12646,N_12009,N_12264);
xnor U12647 (N_12647,N_12161,N_12208);
and U12648 (N_12648,N_12131,N_12363);
nand U12649 (N_12649,N_12301,N_12476);
nand U12650 (N_12650,N_12237,N_12438);
nand U12651 (N_12651,N_12163,N_12315);
nand U12652 (N_12652,N_12248,N_12270);
nand U12653 (N_12653,N_12210,N_12345);
nand U12654 (N_12654,N_12353,N_12170);
or U12655 (N_12655,N_12418,N_12380);
or U12656 (N_12656,N_12225,N_12297);
and U12657 (N_12657,N_12222,N_12051);
and U12658 (N_12658,N_12307,N_12075);
and U12659 (N_12659,N_12199,N_12135);
and U12660 (N_12660,N_12089,N_12022);
and U12661 (N_12661,N_12137,N_12207);
nand U12662 (N_12662,N_12078,N_12129);
nor U12663 (N_12663,N_12445,N_12173);
nand U12664 (N_12664,N_12136,N_12188);
nand U12665 (N_12665,N_12119,N_12251);
or U12666 (N_12666,N_12201,N_12185);
nor U12667 (N_12667,N_12109,N_12118);
or U12668 (N_12668,N_12087,N_12157);
nand U12669 (N_12669,N_12492,N_12093);
nand U12670 (N_12670,N_12414,N_12330);
nor U12671 (N_12671,N_12035,N_12252);
or U12672 (N_12672,N_12002,N_12464);
nor U12673 (N_12673,N_12337,N_12013);
nand U12674 (N_12674,N_12338,N_12331);
nor U12675 (N_12675,N_12376,N_12141);
and U12676 (N_12676,N_12026,N_12489);
and U12677 (N_12677,N_12146,N_12183);
nor U12678 (N_12678,N_12139,N_12110);
nor U12679 (N_12679,N_12000,N_12187);
nand U12680 (N_12680,N_12400,N_12094);
nand U12681 (N_12681,N_12412,N_12296);
or U12682 (N_12682,N_12195,N_12044);
or U12683 (N_12683,N_12396,N_12292);
nand U12684 (N_12684,N_12304,N_12275);
and U12685 (N_12685,N_12460,N_12238);
nand U12686 (N_12686,N_12449,N_12265);
and U12687 (N_12687,N_12332,N_12072);
xnor U12688 (N_12688,N_12478,N_12372);
and U12689 (N_12689,N_12397,N_12484);
nor U12690 (N_12690,N_12007,N_12231);
or U12691 (N_12691,N_12405,N_12068);
and U12692 (N_12692,N_12128,N_12336);
or U12693 (N_12693,N_12028,N_12169);
nor U12694 (N_12694,N_12374,N_12287);
and U12695 (N_12695,N_12209,N_12426);
or U12696 (N_12696,N_12481,N_12166);
or U12697 (N_12697,N_12394,N_12120);
nor U12698 (N_12698,N_12042,N_12472);
nand U12699 (N_12699,N_12298,N_12417);
or U12700 (N_12700,N_12123,N_12379);
nor U12701 (N_12701,N_12448,N_12241);
nor U12702 (N_12702,N_12001,N_12155);
nor U12703 (N_12703,N_12493,N_12452);
nor U12704 (N_12704,N_12034,N_12408);
or U12705 (N_12705,N_12065,N_12299);
nor U12706 (N_12706,N_12240,N_12320);
or U12707 (N_12707,N_12103,N_12271);
and U12708 (N_12708,N_12440,N_12366);
nor U12709 (N_12709,N_12182,N_12280);
and U12710 (N_12710,N_12032,N_12411);
and U12711 (N_12711,N_12088,N_12036);
or U12712 (N_12712,N_12485,N_12341);
nand U12713 (N_12713,N_12284,N_12092);
or U12714 (N_12714,N_12218,N_12203);
or U12715 (N_12715,N_12470,N_12308);
nor U12716 (N_12716,N_12005,N_12410);
or U12717 (N_12717,N_12273,N_12206);
and U12718 (N_12718,N_12246,N_12104);
or U12719 (N_12719,N_12279,N_12242);
nand U12720 (N_12720,N_12487,N_12167);
and U12721 (N_12721,N_12024,N_12172);
and U12722 (N_12722,N_12077,N_12041);
nor U12723 (N_12723,N_12256,N_12268);
and U12724 (N_12724,N_12012,N_12255);
or U12725 (N_12725,N_12269,N_12429);
or U12726 (N_12726,N_12420,N_12383);
nor U12727 (N_12727,N_12224,N_12216);
nor U12728 (N_12728,N_12469,N_12098);
or U12729 (N_12729,N_12016,N_12471);
and U12730 (N_12730,N_12444,N_12200);
nand U12731 (N_12731,N_12111,N_12483);
nand U12732 (N_12732,N_12335,N_12046);
nor U12733 (N_12733,N_12313,N_12179);
or U12734 (N_12734,N_12350,N_12390);
nand U12735 (N_12735,N_12399,N_12319);
nor U12736 (N_12736,N_12029,N_12178);
or U12737 (N_12737,N_12339,N_12425);
and U12738 (N_12738,N_12442,N_12193);
nor U12739 (N_12739,N_12406,N_12491);
or U12740 (N_12740,N_12415,N_12063);
or U12741 (N_12741,N_12003,N_12466);
and U12742 (N_12742,N_12261,N_12091);
nand U12743 (N_12743,N_12189,N_12427);
and U12744 (N_12744,N_12388,N_12038);
nand U12745 (N_12745,N_12434,N_12239);
and U12746 (N_12746,N_12294,N_12102);
nor U12747 (N_12747,N_12305,N_12177);
and U12748 (N_12748,N_12459,N_12443);
and U12749 (N_12749,N_12377,N_12130);
nor U12750 (N_12750,N_12150,N_12306);
or U12751 (N_12751,N_12112,N_12274);
and U12752 (N_12752,N_12004,N_12299);
nor U12753 (N_12753,N_12173,N_12123);
or U12754 (N_12754,N_12024,N_12124);
or U12755 (N_12755,N_12029,N_12133);
or U12756 (N_12756,N_12049,N_12110);
and U12757 (N_12757,N_12145,N_12132);
nand U12758 (N_12758,N_12340,N_12022);
and U12759 (N_12759,N_12305,N_12173);
and U12760 (N_12760,N_12185,N_12317);
nor U12761 (N_12761,N_12443,N_12474);
and U12762 (N_12762,N_12363,N_12256);
nand U12763 (N_12763,N_12428,N_12156);
and U12764 (N_12764,N_12122,N_12304);
and U12765 (N_12765,N_12305,N_12388);
or U12766 (N_12766,N_12327,N_12274);
or U12767 (N_12767,N_12137,N_12005);
nor U12768 (N_12768,N_12478,N_12214);
nand U12769 (N_12769,N_12273,N_12310);
nor U12770 (N_12770,N_12006,N_12347);
nor U12771 (N_12771,N_12034,N_12059);
and U12772 (N_12772,N_12326,N_12260);
and U12773 (N_12773,N_12304,N_12408);
and U12774 (N_12774,N_12302,N_12149);
or U12775 (N_12775,N_12114,N_12188);
or U12776 (N_12776,N_12492,N_12462);
or U12777 (N_12777,N_12381,N_12228);
nand U12778 (N_12778,N_12437,N_12418);
nand U12779 (N_12779,N_12202,N_12246);
nor U12780 (N_12780,N_12027,N_12455);
nand U12781 (N_12781,N_12210,N_12357);
or U12782 (N_12782,N_12462,N_12427);
or U12783 (N_12783,N_12491,N_12379);
or U12784 (N_12784,N_12009,N_12064);
or U12785 (N_12785,N_12274,N_12362);
and U12786 (N_12786,N_12386,N_12136);
and U12787 (N_12787,N_12046,N_12394);
nand U12788 (N_12788,N_12102,N_12050);
or U12789 (N_12789,N_12346,N_12438);
nor U12790 (N_12790,N_12132,N_12407);
or U12791 (N_12791,N_12375,N_12359);
nand U12792 (N_12792,N_12043,N_12407);
nand U12793 (N_12793,N_12200,N_12098);
nor U12794 (N_12794,N_12453,N_12264);
nand U12795 (N_12795,N_12434,N_12124);
nor U12796 (N_12796,N_12378,N_12104);
nor U12797 (N_12797,N_12101,N_12280);
or U12798 (N_12798,N_12028,N_12124);
nand U12799 (N_12799,N_12456,N_12261);
and U12800 (N_12800,N_12094,N_12454);
nand U12801 (N_12801,N_12469,N_12281);
nand U12802 (N_12802,N_12365,N_12215);
nor U12803 (N_12803,N_12052,N_12026);
nor U12804 (N_12804,N_12153,N_12252);
nor U12805 (N_12805,N_12356,N_12453);
nand U12806 (N_12806,N_12282,N_12425);
and U12807 (N_12807,N_12178,N_12280);
nor U12808 (N_12808,N_12211,N_12489);
or U12809 (N_12809,N_12091,N_12095);
and U12810 (N_12810,N_12404,N_12245);
and U12811 (N_12811,N_12408,N_12240);
or U12812 (N_12812,N_12050,N_12170);
or U12813 (N_12813,N_12328,N_12086);
or U12814 (N_12814,N_12187,N_12454);
nand U12815 (N_12815,N_12194,N_12337);
nor U12816 (N_12816,N_12160,N_12118);
or U12817 (N_12817,N_12234,N_12293);
nand U12818 (N_12818,N_12463,N_12391);
nand U12819 (N_12819,N_12200,N_12223);
or U12820 (N_12820,N_12284,N_12215);
nor U12821 (N_12821,N_12435,N_12003);
nor U12822 (N_12822,N_12287,N_12306);
nor U12823 (N_12823,N_12027,N_12057);
nand U12824 (N_12824,N_12286,N_12168);
nor U12825 (N_12825,N_12194,N_12384);
and U12826 (N_12826,N_12076,N_12266);
and U12827 (N_12827,N_12276,N_12151);
and U12828 (N_12828,N_12265,N_12482);
nand U12829 (N_12829,N_12316,N_12395);
and U12830 (N_12830,N_12289,N_12445);
or U12831 (N_12831,N_12019,N_12476);
nand U12832 (N_12832,N_12414,N_12395);
nand U12833 (N_12833,N_12324,N_12087);
nand U12834 (N_12834,N_12239,N_12338);
and U12835 (N_12835,N_12041,N_12467);
nand U12836 (N_12836,N_12403,N_12457);
nor U12837 (N_12837,N_12356,N_12039);
nand U12838 (N_12838,N_12406,N_12134);
or U12839 (N_12839,N_12248,N_12163);
nand U12840 (N_12840,N_12319,N_12042);
or U12841 (N_12841,N_12293,N_12402);
nor U12842 (N_12842,N_12085,N_12127);
or U12843 (N_12843,N_12481,N_12145);
nand U12844 (N_12844,N_12072,N_12407);
and U12845 (N_12845,N_12315,N_12088);
nor U12846 (N_12846,N_12024,N_12059);
and U12847 (N_12847,N_12423,N_12209);
nor U12848 (N_12848,N_12023,N_12144);
or U12849 (N_12849,N_12216,N_12439);
or U12850 (N_12850,N_12419,N_12087);
nor U12851 (N_12851,N_12144,N_12194);
or U12852 (N_12852,N_12312,N_12113);
nand U12853 (N_12853,N_12217,N_12436);
or U12854 (N_12854,N_12289,N_12243);
and U12855 (N_12855,N_12496,N_12042);
nor U12856 (N_12856,N_12099,N_12433);
or U12857 (N_12857,N_12013,N_12401);
nand U12858 (N_12858,N_12473,N_12289);
and U12859 (N_12859,N_12422,N_12354);
nor U12860 (N_12860,N_12274,N_12482);
nor U12861 (N_12861,N_12350,N_12021);
or U12862 (N_12862,N_12229,N_12431);
nor U12863 (N_12863,N_12216,N_12234);
or U12864 (N_12864,N_12183,N_12462);
nand U12865 (N_12865,N_12472,N_12021);
or U12866 (N_12866,N_12160,N_12219);
and U12867 (N_12867,N_12226,N_12195);
or U12868 (N_12868,N_12416,N_12237);
nor U12869 (N_12869,N_12457,N_12123);
nor U12870 (N_12870,N_12160,N_12157);
and U12871 (N_12871,N_12371,N_12077);
nand U12872 (N_12872,N_12357,N_12193);
xnor U12873 (N_12873,N_12434,N_12365);
and U12874 (N_12874,N_12155,N_12368);
or U12875 (N_12875,N_12147,N_12059);
and U12876 (N_12876,N_12109,N_12084);
nand U12877 (N_12877,N_12151,N_12393);
and U12878 (N_12878,N_12024,N_12414);
or U12879 (N_12879,N_12301,N_12358);
or U12880 (N_12880,N_12027,N_12114);
nor U12881 (N_12881,N_12265,N_12397);
and U12882 (N_12882,N_12275,N_12136);
nor U12883 (N_12883,N_12191,N_12399);
or U12884 (N_12884,N_12240,N_12238);
and U12885 (N_12885,N_12227,N_12497);
and U12886 (N_12886,N_12022,N_12202);
nor U12887 (N_12887,N_12270,N_12274);
nor U12888 (N_12888,N_12380,N_12372);
xnor U12889 (N_12889,N_12326,N_12352);
nor U12890 (N_12890,N_12057,N_12028);
and U12891 (N_12891,N_12442,N_12238);
or U12892 (N_12892,N_12095,N_12094);
nand U12893 (N_12893,N_12161,N_12303);
or U12894 (N_12894,N_12261,N_12347);
or U12895 (N_12895,N_12166,N_12274);
nor U12896 (N_12896,N_12072,N_12080);
nor U12897 (N_12897,N_12195,N_12021);
nor U12898 (N_12898,N_12221,N_12256);
or U12899 (N_12899,N_12247,N_12004);
and U12900 (N_12900,N_12275,N_12045);
or U12901 (N_12901,N_12161,N_12403);
and U12902 (N_12902,N_12033,N_12338);
or U12903 (N_12903,N_12004,N_12390);
or U12904 (N_12904,N_12007,N_12329);
nand U12905 (N_12905,N_12434,N_12430);
nand U12906 (N_12906,N_12390,N_12444);
nor U12907 (N_12907,N_12421,N_12256);
nand U12908 (N_12908,N_12344,N_12260);
or U12909 (N_12909,N_12291,N_12290);
nand U12910 (N_12910,N_12414,N_12235);
nand U12911 (N_12911,N_12309,N_12340);
and U12912 (N_12912,N_12041,N_12495);
nor U12913 (N_12913,N_12177,N_12468);
nor U12914 (N_12914,N_12324,N_12413);
nand U12915 (N_12915,N_12346,N_12181);
nand U12916 (N_12916,N_12136,N_12094);
nor U12917 (N_12917,N_12234,N_12138);
nand U12918 (N_12918,N_12057,N_12002);
nor U12919 (N_12919,N_12443,N_12064);
nor U12920 (N_12920,N_12438,N_12332);
or U12921 (N_12921,N_12263,N_12095);
and U12922 (N_12922,N_12418,N_12028);
or U12923 (N_12923,N_12103,N_12442);
or U12924 (N_12924,N_12199,N_12027);
or U12925 (N_12925,N_12121,N_12243);
and U12926 (N_12926,N_12303,N_12216);
nor U12927 (N_12927,N_12469,N_12267);
or U12928 (N_12928,N_12042,N_12300);
nand U12929 (N_12929,N_12205,N_12038);
nor U12930 (N_12930,N_12234,N_12213);
or U12931 (N_12931,N_12059,N_12205);
and U12932 (N_12932,N_12147,N_12318);
nor U12933 (N_12933,N_12366,N_12074);
or U12934 (N_12934,N_12264,N_12485);
nor U12935 (N_12935,N_12330,N_12488);
nand U12936 (N_12936,N_12166,N_12455);
nand U12937 (N_12937,N_12353,N_12201);
nor U12938 (N_12938,N_12050,N_12322);
nor U12939 (N_12939,N_12343,N_12490);
or U12940 (N_12940,N_12497,N_12405);
or U12941 (N_12941,N_12221,N_12223);
and U12942 (N_12942,N_12410,N_12460);
or U12943 (N_12943,N_12427,N_12210);
nand U12944 (N_12944,N_12122,N_12029);
nor U12945 (N_12945,N_12195,N_12054);
or U12946 (N_12946,N_12468,N_12315);
nand U12947 (N_12947,N_12116,N_12272);
and U12948 (N_12948,N_12285,N_12255);
and U12949 (N_12949,N_12173,N_12048);
nand U12950 (N_12950,N_12095,N_12355);
nand U12951 (N_12951,N_12320,N_12112);
nor U12952 (N_12952,N_12213,N_12201);
or U12953 (N_12953,N_12185,N_12278);
and U12954 (N_12954,N_12227,N_12445);
nand U12955 (N_12955,N_12026,N_12162);
nand U12956 (N_12956,N_12019,N_12379);
or U12957 (N_12957,N_12112,N_12305);
nor U12958 (N_12958,N_12315,N_12046);
and U12959 (N_12959,N_12181,N_12038);
nand U12960 (N_12960,N_12366,N_12199);
nor U12961 (N_12961,N_12081,N_12385);
and U12962 (N_12962,N_12333,N_12391);
nand U12963 (N_12963,N_12124,N_12224);
nand U12964 (N_12964,N_12204,N_12001);
nor U12965 (N_12965,N_12028,N_12084);
and U12966 (N_12966,N_12289,N_12234);
and U12967 (N_12967,N_12097,N_12314);
nand U12968 (N_12968,N_12262,N_12182);
and U12969 (N_12969,N_12443,N_12122);
nor U12970 (N_12970,N_12199,N_12372);
and U12971 (N_12971,N_12388,N_12136);
nand U12972 (N_12972,N_12023,N_12012);
and U12973 (N_12973,N_12357,N_12071);
nor U12974 (N_12974,N_12483,N_12108);
nand U12975 (N_12975,N_12174,N_12213);
nor U12976 (N_12976,N_12008,N_12132);
and U12977 (N_12977,N_12088,N_12243);
nand U12978 (N_12978,N_12016,N_12269);
or U12979 (N_12979,N_12446,N_12163);
and U12980 (N_12980,N_12117,N_12092);
and U12981 (N_12981,N_12252,N_12199);
and U12982 (N_12982,N_12494,N_12100);
or U12983 (N_12983,N_12456,N_12402);
and U12984 (N_12984,N_12107,N_12003);
nor U12985 (N_12985,N_12258,N_12382);
nor U12986 (N_12986,N_12276,N_12304);
and U12987 (N_12987,N_12152,N_12073);
nand U12988 (N_12988,N_12488,N_12256);
or U12989 (N_12989,N_12395,N_12157);
nand U12990 (N_12990,N_12208,N_12138);
nand U12991 (N_12991,N_12280,N_12076);
and U12992 (N_12992,N_12483,N_12190);
and U12993 (N_12993,N_12024,N_12181);
and U12994 (N_12994,N_12446,N_12443);
or U12995 (N_12995,N_12226,N_12016);
nand U12996 (N_12996,N_12375,N_12256);
or U12997 (N_12997,N_12001,N_12196);
nand U12998 (N_12998,N_12149,N_12087);
nand U12999 (N_12999,N_12081,N_12158);
nand U13000 (N_13000,N_12659,N_12742);
and U13001 (N_13001,N_12584,N_12967);
xnor U13002 (N_13002,N_12518,N_12725);
nor U13003 (N_13003,N_12551,N_12624);
or U13004 (N_13004,N_12524,N_12996);
nor U13005 (N_13005,N_12707,N_12912);
nor U13006 (N_13006,N_12515,N_12739);
nand U13007 (N_13007,N_12962,N_12648);
nand U13008 (N_13008,N_12928,N_12651);
nor U13009 (N_13009,N_12708,N_12669);
and U13010 (N_13010,N_12621,N_12630);
nor U13011 (N_13011,N_12597,N_12709);
nand U13012 (N_13012,N_12803,N_12658);
nor U13013 (N_13013,N_12687,N_12556);
nor U13014 (N_13014,N_12570,N_12843);
and U13015 (N_13015,N_12649,N_12741);
or U13016 (N_13016,N_12797,N_12559);
or U13017 (N_13017,N_12922,N_12886);
nor U13018 (N_13018,N_12506,N_12854);
or U13019 (N_13019,N_12729,N_12665);
nor U13020 (N_13020,N_12527,N_12593);
nor U13021 (N_13021,N_12523,N_12986);
and U13022 (N_13022,N_12587,N_12892);
nand U13023 (N_13023,N_12756,N_12948);
and U13024 (N_13024,N_12606,N_12664);
nor U13025 (N_13025,N_12757,N_12615);
and U13026 (N_13026,N_12623,N_12572);
or U13027 (N_13027,N_12857,N_12504);
nand U13028 (N_13028,N_12601,N_12957);
and U13029 (N_13029,N_12812,N_12721);
nor U13030 (N_13030,N_12530,N_12543);
or U13031 (N_13031,N_12550,N_12746);
nor U13032 (N_13032,N_12531,N_12848);
or U13033 (N_13033,N_12813,N_12569);
nand U13034 (N_13034,N_12824,N_12532);
or U13035 (N_13035,N_12882,N_12685);
and U13036 (N_13036,N_12937,N_12804);
nand U13037 (N_13037,N_12971,N_12560);
nand U13038 (N_13038,N_12642,N_12655);
or U13039 (N_13039,N_12865,N_12952);
nand U13040 (N_13040,N_12613,N_12701);
nand U13041 (N_13041,N_12713,N_12686);
nor U13042 (N_13042,N_12696,N_12694);
nand U13043 (N_13043,N_12977,N_12808);
nor U13044 (N_13044,N_12974,N_12590);
nor U13045 (N_13045,N_12941,N_12810);
nor U13046 (N_13046,N_12512,N_12575);
nand U13047 (N_13047,N_12945,N_12950);
nor U13048 (N_13048,N_12825,N_12517);
nor U13049 (N_13049,N_12548,N_12960);
nor U13050 (N_13050,N_12722,N_12758);
and U13051 (N_13051,N_12975,N_12700);
or U13052 (N_13052,N_12862,N_12902);
nand U13053 (N_13053,N_12919,N_12732);
and U13054 (N_13054,N_12782,N_12763);
nand U13055 (N_13055,N_12987,N_12993);
nor U13056 (N_13056,N_12896,N_12586);
nand U13057 (N_13057,N_12540,N_12958);
or U13058 (N_13058,N_12894,N_12784);
or U13059 (N_13059,N_12925,N_12851);
nor U13060 (N_13060,N_12616,N_12985);
and U13061 (N_13061,N_12668,N_12845);
and U13062 (N_13062,N_12650,N_12682);
nor U13063 (N_13063,N_12944,N_12787);
or U13064 (N_13064,N_12995,N_12869);
nand U13065 (N_13065,N_12988,N_12814);
nor U13066 (N_13066,N_12726,N_12927);
and U13067 (N_13067,N_12728,N_12744);
or U13068 (N_13068,N_12695,N_12521);
nand U13069 (N_13069,N_12968,N_12806);
nor U13070 (N_13070,N_12895,N_12963);
xnor U13071 (N_13071,N_12724,N_12915);
nand U13072 (N_13072,N_12893,N_12541);
nand U13073 (N_13073,N_12760,N_12641);
and U13074 (N_13074,N_12508,N_12583);
nor U13075 (N_13075,N_12637,N_12536);
and U13076 (N_13076,N_12863,N_12979);
nor U13077 (N_13077,N_12612,N_12589);
or U13078 (N_13078,N_12594,N_12991);
and U13079 (N_13079,N_12692,N_12826);
or U13080 (N_13080,N_12513,N_12846);
or U13081 (N_13081,N_12801,N_12940);
and U13082 (N_13082,N_12961,N_12998);
nand U13083 (N_13083,N_12720,N_12627);
and U13084 (N_13084,N_12938,N_12926);
or U13085 (N_13085,N_12535,N_12835);
nor U13086 (N_13086,N_12982,N_12607);
xor U13087 (N_13087,N_12661,N_12534);
nor U13088 (N_13088,N_12533,N_12605);
nor U13089 (N_13089,N_12753,N_12883);
or U13090 (N_13090,N_12680,N_12514);
and U13091 (N_13091,N_12859,N_12888);
and U13092 (N_13092,N_12809,N_12678);
xnor U13093 (N_13093,N_12547,N_12703);
or U13094 (N_13094,N_12916,N_12672);
or U13095 (N_13095,N_12702,N_12891);
and U13096 (N_13096,N_12983,N_12574);
nor U13097 (N_13097,N_12749,N_12614);
or U13098 (N_13098,N_12887,N_12565);
nand U13099 (N_13099,N_12914,N_12617);
and U13100 (N_13100,N_12629,N_12830);
or U13101 (N_13101,N_12766,N_12640);
nand U13102 (N_13102,N_12666,N_12779);
nand U13103 (N_13103,N_12662,N_12807);
nor U13104 (N_13104,N_12880,N_12834);
nand U13105 (N_13105,N_12647,N_12871);
nor U13106 (N_13106,N_12727,N_12520);
nor U13107 (N_13107,N_12820,N_12679);
and U13108 (N_13108,N_12546,N_12599);
or U13109 (N_13109,N_12505,N_12833);
or U13110 (N_13110,N_12821,N_12767);
or U13111 (N_13111,N_12693,N_12885);
nor U13112 (N_13112,N_12849,N_12762);
nand U13113 (N_13113,N_12837,N_12622);
and U13114 (N_13114,N_12785,N_12811);
or U13115 (N_13115,N_12911,N_12774);
nor U13116 (N_13116,N_12873,N_12799);
nand U13117 (N_13117,N_12608,N_12566);
nand U13118 (N_13118,N_12596,N_12643);
and U13119 (N_13119,N_12691,N_12549);
or U13120 (N_13120,N_12690,N_12769);
nor U13121 (N_13121,N_12778,N_12832);
and U13122 (N_13122,N_12656,N_12576);
nor U13123 (N_13123,N_12562,N_12924);
nand U13124 (N_13124,N_12723,N_12936);
nand U13125 (N_13125,N_12964,N_12516);
and U13126 (N_13126,N_12667,N_12973);
nor U13127 (N_13127,N_12618,N_12731);
and U13128 (N_13128,N_12852,N_12828);
nand U13129 (N_13129,N_12840,N_12636);
or U13130 (N_13130,N_12634,N_12877);
nor U13131 (N_13131,N_12903,N_12509);
nor U13132 (N_13132,N_12609,N_12639);
and U13133 (N_13133,N_12718,N_12552);
nor U13134 (N_13134,N_12847,N_12684);
and U13135 (N_13135,N_12764,N_12719);
nor U13136 (N_13136,N_12949,N_12561);
and U13137 (N_13137,N_12734,N_12783);
nor U13138 (N_13138,N_12775,N_12717);
nor U13139 (N_13139,N_12573,N_12750);
nor U13140 (N_13140,N_12580,N_12653);
and U13141 (N_13141,N_12677,N_12805);
and U13142 (N_13142,N_12644,N_12878);
or U13143 (N_13143,N_12951,N_12972);
nor U13144 (N_13144,N_12981,N_12999);
or U13145 (N_13145,N_12591,N_12761);
and U13146 (N_13146,N_12676,N_12554);
and U13147 (N_13147,N_12841,N_12781);
nor U13148 (N_13148,N_12595,N_12598);
nor U13149 (N_13149,N_12776,N_12571);
or U13150 (N_13150,N_12542,N_12602);
nor U13151 (N_13151,N_12698,N_12934);
nor U13152 (N_13152,N_12539,N_12681);
nor U13153 (N_13153,N_12791,N_12953);
or U13154 (N_13154,N_12800,N_12790);
and U13155 (N_13155,N_12789,N_12798);
nand U13156 (N_13156,N_12500,N_12836);
and U13157 (N_13157,N_12853,N_12777);
nand U13158 (N_13158,N_12673,N_12923);
nor U13159 (N_13159,N_12752,N_12969);
nor U13160 (N_13160,N_12568,N_12631);
or U13161 (N_13161,N_12646,N_12545);
nor U13162 (N_13162,N_12699,N_12733);
and U13163 (N_13163,N_12970,N_12652);
or U13164 (N_13164,N_12829,N_12959);
or U13165 (N_13165,N_12844,N_12994);
or U13166 (N_13166,N_12992,N_12772);
or U13167 (N_13167,N_12619,N_12870);
or U13168 (N_13168,N_12557,N_12908);
and U13169 (N_13169,N_12933,N_12737);
and U13170 (N_13170,N_12511,N_12989);
and U13171 (N_13171,N_12831,N_12827);
and U13172 (N_13172,N_12850,N_12564);
and U13173 (N_13173,N_12906,N_12946);
nand U13174 (N_13174,N_12671,N_12660);
and U13175 (N_13175,N_12966,N_12978);
or U13176 (N_13176,N_12984,N_12918);
and U13177 (N_13177,N_12884,N_12526);
nand U13178 (N_13178,N_12899,N_12567);
and U13179 (N_13179,N_12954,N_12604);
nor U13180 (N_13180,N_12910,N_12881);
nand U13181 (N_13181,N_12502,N_12901);
nor U13182 (N_13182,N_12751,N_12705);
and U13183 (N_13183,N_12755,N_12558);
and U13184 (N_13184,N_12710,N_12579);
nand U13185 (N_13185,N_12628,N_12633);
nor U13186 (N_13186,N_12675,N_12802);
nor U13187 (N_13187,N_12955,N_12585);
nand U13188 (N_13188,N_12842,N_12905);
or U13189 (N_13189,N_12503,N_12715);
nand U13190 (N_13190,N_12654,N_12889);
nand U13191 (N_13191,N_12942,N_12563);
or U13192 (N_13192,N_12716,N_12839);
and U13193 (N_13193,N_12704,N_12935);
nor U13194 (N_13194,N_12712,N_12822);
or U13195 (N_13195,N_12537,N_12620);
nand U13196 (N_13196,N_12793,N_12578);
or U13197 (N_13197,N_12976,N_12759);
nor U13198 (N_13198,N_12765,N_12610);
and U13199 (N_13199,N_12697,N_12900);
nor U13200 (N_13200,N_12929,N_12625);
nand U13201 (N_13201,N_12740,N_12795);
nor U13202 (N_13202,N_12528,N_12943);
and U13203 (N_13203,N_12507,N_12921);
nor U13204 (N_13204,N_12861,N_12711);
and U13205 (N_13205,N_12754,N_12786);
and U13206 (N_13206,N_12768,N_12730);
nand U13207 (N_13207,N_12815,N_12931);
or U13208 (N_13208,N_12626,N_12980);
nand U13209 (N_13209,N_12674,N_12510);
or U13210 (N_13210,N_12736,N_12773);
and U13211 (N_13211,N_12868,N_12688);
and U13212 (N_13212,N_12907,N_12747);
and U13213 (N_13213,N_12600,N_12816);
nor U13214 (N_13214,N_12932,N_12683);
nand U13215 (N_13215,N_12838,N_12663);
nor U13216 (N_13216,N_12582,N_12738);
nor U13217 (N_13217,N_12522,N_12909);
or U13218 (N_13218,N_12858,N_12920);
nand U13219 (N_13219,N_12792,N_12897);
and U13220 (N_13220,N_12866,N_12771);
nor U13221 (N_13221,N_12670,N_12917);
and U13222 (N_13222,N_12544,N_12947);
nor U13223 (N_13223,N_12635,N_12898);
nor U13224 (N_13224,N_12529,N_12872);
nand U13225 (N_13225,N_12525,N_12611);
and U13226 (N_13226,N_12745,N_12904);
nor U13227 (N_13227,N_12875,N_12519);
nor U13228 (N_13228,N_12735,N_12788);
or U13229 (N_13229,N_12657,N_12879);
or U13230 (N_13230,N_12714,N_12770);
nand U13231 (N_13231,N_12553,N_12939);
nor U13232 (N_13232,N_12796,N_12603);
and U13233 (N_13233,N_12689,N_12577);
or U13234 (N_13234,N_12588,N_12743);
nor U13235 (N_13235,N_12632,N_12638);
nor U13236 (N_13236,N_12956,N_12890);
or U13237 (N_13237,N_12965,N_12748);
nand U13238 (N_13238,N_12581,N_12818);
nor U13239 (N_13239,N_12538,N_12706);
and U13240 (N_13240,N_12794,N_12930);
or U13241 (N_13241,N_12819,N_12867);
or U13242 (N_13242,N_12780,N_12817);
or U13243 (N_13243,N_12645,N_12874);
nor U13244 (N_13244,N_12990,N_12997);
and U13245 (N_13245,N_12501,N_12555);
nand U13246 (N_13246,N_12876,N_12864);
nor U13247 (N_13247,N_12856,N_12823);
nand U13248 (N_13248,N_12860,N_12592);
nor U13249 (N_13249,N_12855,N_12913);
or U13250 (N_13250,N_12716,N_12678);
or U13251 (N_13251,N_12827,N_12721);
and U13252 (N_13252,N_12527,N_12953);
nand U13253 (N_13253,N_12928,N_12810);
and U13254 (N_13254,N_12723,N_12637);
nor U13255 (N_13255,N_12500,N_12945);
or U13256 (N_13256,N_12744,N_12905);
or U13257 (N_13257,N_12623,N_12514);
nand U13258 (N_13258,N_12825,N_12797);
or U13259 (N_13259,N_12981,N_12727);
nor U13260 (N_13260,N_12876,N_12974);
nor U13261 (N_13261,N_12636,N_12967);
and U13262 (N_13262,N_12572,N_12667);
nor U13263 (N_13263,N_12869,N_12619);
nor U13264 (N_13264,N_12899,N_12894);
nor U13265 (N_13265,N_12927,N_12887);
nand U13266 (N_13266,N_12829,N_12504);
nor U13267 (N_13267,N_12739,N_12844);
nor U13268 (N_13268,N_12851,N_12820);
nor U13269 (N_13269,N_12913,N_12503);
nor U13270 (N_13270,N_12901,N_12781);
or U13271 (N_13271,N_12816,N_12529);
or U13272 (N_13272,N_12973,N_12586);
and U13273 (N_13273,N_12824,N_12630);
nand U13274 (N_13274,N_12512,N_12866);
or U13275 (N_13275,N_12511,N_12940);
and U13276 (N_13276,N_12823,N_12719);
and U13277 (N_13277,N_12926,N_12969);
nand U13278 (N_13278,N_12552,N_12985);
nand U13279 (N_13279,N_12733,N_12589);
or U13280 (N_13280,N_12773,N_12921);
and U13281 (N_13281,N_12662,N_12602);
nand U13282 (N_13282,N_12527,N_12588);
nand U13283 (N_13283,N_12840,N_12519);
and U13284 (N_13284,N_12646,N_12862);
nor U13285 (N_13285,N_12562,N_12589);
nor U13286 (N_13286,N_12549,N_12982);
nor U13287 (N_13287,N_12809,N_12915);
xnor U13288 (N_13288,N_12779,N_12543);
nand U13289 (N_13289,N_12785,N_12711);
nor U13290 (N_13290,N_12795,N_12515);
or U13291 (N_13291,N_12534,N_12697);
and U13292 (N_13292,N_12618,N_12637);
nand U13293 (N_13293,N_12546,N_12796);
nor U13294 (N_13294,N_12967,N_12553);
and U13295 (N_13295,N_12544,N_12811);
and U13296 (N_13296,N_12932,N_12638);
and U13297 (N_13297,N_12679,N_12532);
and U13298 (N_13298,N_12812,N_12906);
and U13299 (N_13299,N_12925,N_12547);
or U13300 (N_13300,N_12568,N_12663);
and U13301 (N_13301,N_12602,N_12882);
nand U13302 (N_13302,N_12513,N_12803);
or U13303 (N_13303,N_12911,N_12931);
and U13304 (N_13304,N_12642,N_12855);
nand U13305 (N_13305,N_12819,N_12966);
or U13306 (N_13306,N_12679,N_12872);
nor U13307 (N_13307,N_12721,N_12915);
or U13308 (N_13308,N_12772,N_12615);
or U13309 (N_13309,N_12933,N_12864);
or U13310 (N_13310,N_12894,N_12793);
and U13311 (N_13311,N_12840,N_12987);
or U13312 (N_13312,N_12613,N_12648);
or U13313 (N_13313,N_12839,N_12996);
nor U13314 (N_13314,N_12786,N_12654);
nand U13315 (N_13315,N_12619,N_12670);
or U13316 (N_13316,N_12541,N_12918);
and U13317 (N_13317,N_12890,N_12532);
or U13318 (N_13318,N_12753,N_12917);
or U13319 (N_13319,N_12508,N_12840);
nand U13320 (N_13320,N_12713,N_12707);
and U13321 (N_13321,N_12713,N_12822);
nand U13322 (N_13322,N_12979,N_12779);
and U13323 (N_13323,N_12579,N_12748);
and U13324 (N_13324,N_12549,N_12889);
or U13325 (N_13325,N_12609,N_12637);
or U13326 (N_13326,N_12615,N_12636);
nand U13327 (N_13327,N_12804,N_12693);
nor U13328 (N_13328,N_12785,N_12896);
and U13329 (N_13329,N_12868,N_12539);
nor U13330 (N_13330,N_12650,N_12729);
nand U13331 (N_13331,N_12697,N_12782);
nor U13332 (N_13332,N_12730,N_12859);
and U13333 (N_13333,N_12661,N_12978);
nor U13334 (N_13334,N_12671,N_12566);
or U13335 (N_13335,N_12701,N_12644);
nand U13336 (N_13336,N_12729,N_12981);
or U13337 (N_13337,N_12681,N_12925);
nand U13338 (N_13338,N_12532,N_12913);
nand U13339 (N_13339,N_12780,N_12543);
and U13340 (N_13340,N_12950,N_12877);
nor U13341 (N_13341,N_12666,N_12938);
xnor U13342 (N_13342,N_12624,N_12943);
and U13343 (N_13343,N_12876,N_12613);
and U13344 (N_13344,N_12596,N_12808);
nand U13345 (N_13345,N_12681,N_12654);
nand U13346 (N_13346,N_12695,N_12618);
nor U13347 (N_13347,N_12628,N_12766);
nor U13348 (N_13348,N_12619,N_12880);
nand U13349 (N_13349,N_12506,N_12600);
nand U13350 (N_13350,N_12529,N_12571);
or U13351 (N_13351,N_12678,N_12821);
and U13352 (N_13352,N_12692,N_12545);
and U13353 (N_13353,N_12500,N_12766);
nand U13354 (N_13354,N_12621,N_12787);
nand U13355 (N_13355,N_12567,N_12645);
and U13356 (N_13356,N_12917,N_12727);
nand U13357 (N_13357,N_12594,N_12961);
or U13358 (N_13358,N_12513,N_12706);
and U13359 (N_13359,N_12885,N_12771);
nand U13360 (N_13360,N_12845,N_12968);
and U13361 (N_13361,N_12910,N_12569);
nand U13362 (N_13362,N_12976,N_12998);
or U13363 (N_13363,N_12976,N_12916);
and U13364 (N_13364,N_12934,N_12858);
nor U13365 (N_13365,N_12638,N_12816);
nand U13366 (N_13366,N_12771,N_12828);
or U13367 (N_13367,N_12751,N_12858);
nor U13368 (N_13368,N_12568,N_12625);
and U13369 (N_13369,N_12920,N_12770);
nor U13370 (N_13370,N_12796,N_12999);
and U13371 (N_13371,N_12938,N_12942);
nor U13372 (N_13372,N_12598,N_12849);
nor U13373 (N_13373,N_12813,N_12580);
nor U13374 (N_13374,N_12774,N_12659);
and U13375 (N_13375,N_12619,N_12618);
or U13376 (N_13376,N_12862,N_12823);
and U13377 (N_13377,N_12524,N_12859);
or U13378 (N_13378,N_12687,N_12778);
or U13379 (N_13379,N_12605,N_12674);
nand U13380 (N_13380,N_12566,N_12697);
nor U13381 (N_13381,N_12656,N_12689);
nand U13382 (N_13382,N_12740,N_12531);
and U13383 (N_13383,N_12722,N_12735);
and U13384 (N_13384,N_12998,N_12552);
or U13385 (N_13385,N_12519,N_12539);
and U13386 (N_13386,N_12619,N_12886);
nor U13387 (N_13387,N_12872,N_12861);
nand U13388 (N_13388,N_12952,N_12828);
or U13389 (N_13389,N_12771,N_12620);
nor U13390 (N_13390,N_12609,N_12516);
or U13391 (N_13391,N_12730,N_12613);
or U13392 (N_13392,N_12852,N_12608);
and U13393 (N_13393,N_12575,N_12663);
nand U13394 (N_13394,N_12790,N_12801);
or U13395 (N_13395,N_12904,N_12608);
or U13396 (N_13396,N_12892,N_12836);
or U13397 (N_13397,N_12737,N_12628);
and U13398 (N_13398,N_12607,N_12555);
nand U13399 (N_13399,N_12679,N_12885);
and U13400 (N_13400,N_12528,N_12643);
or U13401 (N_13401,N_12809,N_12565);
or U13402 (N_13402,N_12645,N_12563);
or U13403 (N_13403,N_12580,N_12816);
nand U13404 (N_13404,N_12831,N_12810);
and U13405 (N_13405,N_12718,N_12528);
nor U13406 (N_13406,N_12586,N_12803);
nand U13407 (N_13407,N_12670,N_12510);
or U13408 (N_13408,N_12850,N_12680);
nand U13409 (N_13409,N_12533,N_12886);
or U13410 (N_13410,N_12971,N_12681);
and U13411 (N_13411,N_12964,N_12510);
nand U13412 (N_13412,N_12630,N_12821);
and U13413 (N_13413,N_12661,N_12567);
and U13414 (N_13414,N_12653,N_12704);
and U13415 (N_13415,N_12910,N_12719);
nand U13416 (N_13416,N_12895,N_12664);
and U13417 (N_13417,N_12552,N_12578);
nand U13418 (N_13418,N_12526,N_12897);
and U13419 (N_13419,N_12564,N_12710);
nand U13420 (N_13420,N_12725,N_12814);
and U13421 (N_13421,N_12850,N_12615);
nand U13422 (N_13422,N_12612,N_12933);
or U13423 (N_13423,N_12731,N_12560);
nor U13424 (N_13424,N_12595,N_12753);
or U13425 (N_13425,N_12818,N_12861);
or U13426 (N_13426,N_12808,N_12761);
nor U13427 (N_13427,N_12550,N_12645);
nor U13428 (N_13428,N_12545,N_12822);
and U13429 (N_13429,N_12739,N_12906);
xor U13430 (N_13430,N_12543,N_12950);
and U13431 (N_13431,N_12918,N_12698);
nor U13432 (N_13432,N_12625,N_12793);
and U13433 (N_13433,N_12742,N_12744);
or U13434 (N_13434,N_12667,N_12808);
nor U13435 (N_13435,N_12897,N_12711);
nor U13436 (N_13436,N_12636,N_12810);
nand U13437 (N_13437,N_12978,N_12603);
nand U13438 (N_13438,N_12613,N_12758);
nand U13439 (N_13439,N_12828,N_12727);
nor U13440 (N_13440,N_12630,N_12858);
and U13441 (N_13441,N_12932,N_12935);
xnor U13442 (N_13442,N_12531,N_12764);
and U13443 (N_13443,N_12874,N_12831);
nand U13444 (N_13444,N_12869,N_12835);
and U13445 (N_13445,N_12698,N_12887);
nand U13446 (N_13446,N_12769,N_12795);
or U13447 (N_13447,N_12577,N_12541);
or U13448 (N_13448,N_12904,N_12774);
and U13449 (N_13449,N_12919,N_12926);
and U13450 (N_13450,N_12534,N_12682);
nor U13451 (N_13451,N_12613,N_12709);
nand U13452 (N_13452,N_12979,N_12923);
nor U13453 (N_13453,N_12771,N_12766);
nand U13454 (N_13454,N_12981,N_12774);
or U13455 (N_13455,N_12632,N_12639);
and U13456 (N_13456,N_12863,N_12725);
nand U13457 (N_13457,N_12857,N_12672);
nor U13458 (N_13458,N_12515,N_12755);
and U13459 (N_13459,N_12560,N_12872);
and U13460 (N_13460,N_12686,N_12585);
nand U13461 (N_13461,N_12772,N_12855);
and U13462 (N_13462,N_12508,N_12750);
and U13463 (N_13463,N_12878,N_12769);
or U13464 (N_13464,N_12599,N_12795);
and U13465 (N_13465,N_12779,N_12695);
nand U13466 (N_13466,N_12510,N_12785);
nand U13467 (N_13467,N_12883,N_12754);
or U13468 (N_13468,N_12511,N_12981);
nand U13469 (N_13469,N_12503,N_12915);
nand U13470 (N_13470,N_12983,N_12720);
nor U13471 (N_13471,N_12986,N_12730);
nor U13472 (N_13472,N_12550,N_12739);
or U13473 (N_13473,N_12876,N_12758);
nor U13474 (N_13474,N_12539,N_12635);
or U13475 (N_13475,N_12881,N_12610);
nand U13476 (N_13476,N_12876,N_12536);
nand U13477 (N_13477,N_12515,N_12767);
nor U13478 (N_13478,N_12577,N_12892);
nand U13479 (N_13479,N_12691,N_12562);
and U13480 (N_13480,N_12832,N_12962);
nand U13481 (N_13481,N_12806,N_12629);
nand U13482 (N_13482,N_12857,N_12902);
nor U13483 (N_13483,N_12826,N_12591);
nand U13484 (N_13484,N_12958,N_12551);
or U13485 (N_13485,N_12582,N_12541);
nor U13486 (N_13486,N_12727,N_12883);
nand U13487 (N_13487,N_12909,N_12505);
or U13488 (N_13488,N_12806,N_12959);
nor U13489 (N_13489,N_12964,N_12676);
and U13490 (N_13490,N_12636,N_12802);
or U13491 (N_13491,N_12988,N_12675);
nor U13492 (N_13492,N_12717,N_12530);
and U13493 (N_13493,N_12826,N_12614);
or U13494 (N_13494,N_12503,N_12765);
or U13495 (N_13495,N_12995,N_12504);
nand U13496 (N_13496,N_12833,N_12634);
or U13497 (N_13497,N_12920,N_12588);
and U13498 (N_13498,N_12633,N_12809);
nand U13499 (N_13499,N_12987,N_12896);
nor U13500 (N_13500,N_13066,N_13385);
nor U13501 (N_13501,N_13040,N_13470);
and U13502 (N_13502,N_13498,N_13301);
and U13503 (N_13503,N_13446,N_13126);
and U13504 (N_13504,N_13319,N_13044);
nor U13505 (N_13505,N_13071,N_13339);
nand U13506 (N_13506,N_13018,N_13223);
or U13507 (N_13507,N_13341,N_13442);
nor U13508 (N_13508,N_13037,N_13233);
nor U13509 (N_13509,N_13101,N_13127);
and U13510 (N_13510,N_13267,N_13202);
nand U13511 (N_13511,N_13343,N_13479);
or U13512 (N_13512,N_13312,N_13140);
and U13513 (N_13513,N_13191,N_13156);
and U13514 (N_13514,N_13180,N_13175);
or U13515 (N_13515,N_13457,N_13057);
or U13516 (N_13516,N_13437,N_13496);
or U13517 (N_13517,N_13225,N_13328);
nor U13518 (N_13518,N_13441,N_13025);
and U13519 (N_13519,N_13234,N_13253);
and U13520 (N_13520,N_13295,N_13249);
or U13521 (N_13521,N_13224,N_13222);
or U13522 (N_13522,N_13240,N_13390);
nor U13523 (N_13523,N_13483,N_13229);
and U13524 (N_13524,N_13375,N_13347);
nand U13525 (N_13525,N_13230,N_13004);
and U13526 (N_13526,N_13166,N_13227);
or U13527 (N_13527,N_13274,N_13194);
or U13528 (N_13528,N_13102,N_13411);
xor U13529 (N_13529,N_13370,N_13447);
or U13530 (N_13530,N_13334,N_13491);
nand U13531 (N_13531,N_13268,N_13056);
nand U13532 (N_13532,N_13368,N_13184);
and U13533 (N_13533,N_13177,N_13336);
nor U13534 (N_13534,N_13287,N_13303);
nand U13535 (N_13535,N_13367,N_13129);
and U13536 (N_13536,N_13389,N_13392);
nor U13537 (N_13537,N_13193,N_13260);
and U13538 (N_13538,N_13484,N_13103);
nand U13539 (N_13539,N_13373,N_13123);
nor U13540 (N_13540,N_13108,N_13073);
nand U13541 (N_13541,N_13308,N_13247);
and U13542 (N_13542,N_13313,N_13409);
nand U13543 (N_13543,N_13391,N_13054);
and U13544 (N_13544,N_13284,N_13176);
nand U13545 (N_13545,N_13246,N_13497);
and U13546 (N_13546,N_13179,N_13417);
and U13547 (N_13547,N_13088,N_13350);
and U13548 (N_13548,N_13327,N_13183);
nand U13549 (N_13549,N_13135,N_13262);
or U13550 (N_13550,N_13003,N_13119);
nand U13551 (N_13551,N_13038,N_13243);
nor U13552 (N_13552,N_13173,N_13265);
nand U13553 (N_13553,N_13214,N_13236);
and U13554 (N_13554,N_13374,N_13257);
and U13555 (N_13555,N_13200,N_13043);
nand U13556 (N_13556,N_13144,N_13450);
or U13557 (N_13557,N_13077,N_13329);
and U13558 (N_13558,N_13047,N_13134);
nor U13559 (N_13559,N_13104,N_13172);
or U13560 (N_13560,N_13460,N_13288);
or U13561 (N_13561,N_13046,N_13415);
and U13562 (N_13562,N_13089,N_13245);
nand U13563 (N_13563,N_13439,N_13051);
nand U13564 (N_13564,N_13143,N_13009);
nor U13565 (N_13565,N_13008,N_13394);
nor U13566 (N_13566,N_13403,N_13205);
or U13567 (N_13567,N_13235,N_13393);
and U13568 (N_13568,N_13293,N_13396);
and U13569 (N_13569,N_13167,N_13091);
or U13570 (N_13570,N_13217,N_13019);
nor U13571 (N_13571,N_13305,N_13399);
or U13572 (N_13572,N_13443,N_13357);
nor U13573 (N_13573,N_13157,N_13188);
and U13574 (N_13574,N_13363,N_13079);
or U13575 (N_13575,N_13386,N_13153);
and U13576 (N_13576,N_13187,N_13307);
or U13577 (N_13577,N_13418,N_13259);
nor U13578 (N_13578,N_13408,N_13416);
or U13579 (N_13579,N_13076,N_13482);
nor U13580 (N_13580,N_13033,N_13467);
and U13581 (N_13581,N_13158,N_13421);
or U13582 (N_13582,N_13364,N_13100);
or U13583 (N_13583,N_13298,N_13142);
nor U13584 (N_13584,N_13139,N_13435);
nor U13585 (N_13585,N_13494,N_13097);
or U13586 (N_13586,N_13039,N_13168);
and U13587 (N_13587,N_13074,N_13318);
nor U13588 (N_13588,N_13086,N_13174);
nor U13589 (N_13589,N_13382,N_13237);
and U13590 (N_13590,N_13053,N_13406);
nand U13591 (N_13591,N_13451,N_13306);
nand U13592 (N_13592,N_13203,N_13152);
nand U13593 (N_13593,N_13349,N_13159);
nand U13594 (N_13594,N_13190,N_13352);
and U13595 (N_13595,N_13321,N_13232);
and U13596 (N_13596,N_13070,N_13407);
nor U13597 (N_13597,N_13429,N_13380);
nor U13598 (N_13598,N_13197,N_13331);
and U13599 (N_13599,N_13252,N_13337);
nand U13600 (N_13600,N_13469,N_13461);
and U13601 (N_13601,N_13000,N_13462);
and U13602 (N_13602,N_13060,N_13058);
or U13603 (N_13603,N_13115,N_13015);
nor U13604 (N_13604,N_13422,N_13304);
nand U13605 (N_13605,N_13125,N_13064);
and U13606 (N_13606,N_13032,N_13261);
or U13607 (N_13607,N_13322,N_13324);
xor U13608 (N_13608,N_13106,N_13006);
or U13609 (N_13609,N_13366,N_13189);
and U13610 (N_13610,N_13419,N_13436);
nand U13611 (N_13611,N_13081,N_13354);
or U13612 (N_13612,N_13198,N_13472);
nor U13613 (N_13613,N_13493,N_13241);
and U13614 (N_13614,N_13445,N_13400);
and U13615 (N_13615,N_13291,N_13340);
nand U13616 (N_13616,N_13438,N_13178);
and U13617 (N_13617,N_13454,N_13210);
and U13618 (N_13618,N_13093,N_13151);
or U13619 (N_13619,N_13365,N_13080);
and U13620 (N_13620,N_13376,N_13410);
nand U13621 (N_13621,N_13464,N_13083);
and U13622 (N_13622,N_13353,N_13286);
or U13623 (N_13623,N_13078,N_13338);
xnor U13624 (N_13624,N_13121,N_13239);
or U13625 (N_13625,N_13024,N_13112);
or U13626 (N_13626,N_13473,N_13300);
and U13627 (N_13627,N_13315,N_13278);
or U13628 (N_13628,N_13448,N_13309);
or U13629 (N_13629,N_13316,N_13122);
or U13630 (N_13630,N_13326,N_13250);
and U13631 (N_13631,N_13030,N_13061);
and U13632 (N_13632,N_13154,N_13413);
nand U13633 (N_13633,N_13013,N_13269);
or U13634 (N_13634,N_13226,N_13397);
nor U13635 (N_13635,N_13209,N_13016);
nor U13636 (N_13636,N_13029,N_13118);
nor U13637 (N_13637,N_13351,N_13317);
nand U13638 (N_13638,N_13490,N_13330);
or U13639 (N_13639,N_13275,N_13186);
nand U13640 (N_13640,N_13036,N_13213);
or U13641 (N_13641,N_13280,N_13358);
or U13642 (N_13642,N_13434,N_13359);
or U13643 (N_13643,N_13345,N_13199);
nand U13644 (N_13644,N_13137,N_13492);
nand U13645 (N_13645,N_13423,N_13480);
nand U13646 (N_13646,N_13474,N_13116);
and U13647 (N_13647,N_13150,N_13310);
or U13648 (N_13648,N_13147,N_13465);
or U13649 (N_13649,N_13201,N_13185);
or U13650 (N_13650,N_13440,N_13132);
and U13651 (N_13651,N_13272,N_13302);
nor U13652 (N_13652,N_13495,N_13471);
and U13653 (N_13653,N_13136,N_13082);
or U13654 (N_13654,N_13485,N_13068);
nand U13655 (N_13655,N_13049,N_13220);
or U13656 (N_13656,N_13022,N_13433);
and U13657 (N_13657,N_13067,N_13196);
and U13658 (N_13658,N_13377,N_13361);
and U13659 (N_13659,N_13042,N_13001);
nor U13660 (N_13660,N_13387,N_13055);
or U13661 (N_13661,N_13065,N_13412);
and U13662 (N_13662,N_13146,N_13458);
or U13663 (N_13663,N_13131,N_13005);
nand U13664 (N_13664,N_13401,N_13320);
nor U13665 (N_13665,N_13105,N_13475);
and U13666 (N_13666,N_13425,N_13251);
nor U13667 (N_13667,N_13087,N_13356);
and U13668 (N_13668,N_13398,N_13052);
and U13669 (N_13669,N_13242,N_13041);
nor U13670 (N_13670,N_13026,N_13372);
nand U13671 (N_13671,N_13459,N_13355);
and U13672 (N_13672,N_13430,N_13164);
and U13673 (N_13673,N_13130,N_13271);
and U13674 (N_13674,N_13427,N_13050);
and U13675 (N_13675,N_13145,N_13362);
nor U13676 (N_13676,N_13133,N_13023);
or U13677 (N_13677,N_13455,N_13325);
nor U13678 (N_13678,N_13273,N_13282);
nand U13679 (N_13679,N_13084,N_13211);
and U13680 (N_13680,N_13072,N_13099);
or U13681 (N_13681,N_13020,N_13010);
nand U13682 (N_13682,N_13170,N_13216);
and U13683 (N_13683,N_13481,N_13276);
nor U13684 (N_13684,N_13031,N_13414);
or U13685 (N_13685,N_13468,N_13110);
nor U13686 (N_13686,N_13169,N_13096);
and U13687 (N_13687,N_13405,N_13378);
nand U13688 (N_13688,N_13486,N_13277);
nor U13689 (N_13689,N_13012,N_13333);
nand U13690 (N_13690,N_13290,N_13212);
or U13691 (N_13691,N_13335,N_13466);
and U13692 (N_13692,N_13182,N_13279);
nor U13693 (N_13693,N_13171,N_13281);
or U13694 (N_13694,N_13141,N_13346);
or U13695 (N_13695,N_13283,N_13007);
or U13696 (N_13696,N_13138,N_13219);
nand U13697 (N_13697,N_13332,N_13034);
or U13698 (N_13698,N_13478,N_13124);
nand U13699 (N_13699,N_13452,N_13014);
nand U13700 (N_13700,N_13092,N_13296);
nor U13701 (N_13701,N_13258,N_13395);
nor U13702 (N_13702,N_13292,N_13476);
and U13703 (N_13703,N_13161,N_13270);
nand U13704 (N_13704,N_13075,N_13059);
and U13705 (N_13705,N_13128,N_13085);
nor U13706 (N_13706,N_13027,N_13488);
and U13707 (N_13707,N_13192,N_13109);
or U13708 (N_13708,N_13255,N_13360);
and U13709 (N_13709,N_13449,N_13371);
and U13710 (N_13710,N_13095,N_13107);
nor U13711 (N_13711,N_13379,N_13113);
nor U13712 (N_13712,N_13221,N_13094);
nand U13713 (N_13713,N_13489,N_13181);
and U13714 (N_13714,N_13456,N_13063);
or U13715 (N_13715,N_13299,N_13155);
nand U13716 (N_13716,N_13297,N_13028);
nand U13717 (N_13717,N_13264,N_13238);
and U13718 (N_13718,N_13424,N_13165);
nand U13719 (N_13719,N_13285,N_13244);
and U13720 (N_13720,N_13149,N_13160);
or U13721 (N_13721,N_13263,N_13289);
nand U13722 (N_13722,N_13311,N_13420);
nand U13723 (N_13723,N_13090,N_13428);
nor U13724 (N_13724,N_13111,N_13195);
nand U13725 (N_13725,N_13404,N_13011);
or U13726 (N_13726,N_13002,N_13402);
nor U13727 (N_13727,N_13477,N_13463);
and U13728 (N_13728,N_13206,N_13062);
nor U13729 (N_13729,N_13444,N_13426);
and U13730 (N_13730,N_13048,N_13388);
nor U13731 (N_13731,N_13021,N_13294);
and U13732 (N_13732,N_13148,N_13314);
nor U13733 (N_13733,N_13323,N_13228);
nand U13734 (N_13734,N_13114,N_13487);
nor U13735 (N_13735,N_13254,N_13208);
nand U13736 (N_13736,N_13499,N_13069);
nor U13737 (N_13737,N_13163,N_13218);
and U13738 (N_13738,N_13045,N_13348);
nand U13739 (N_13739,N_13117,N_13384);
and U13740 (N_13740,N_13035,N_13207);
nand U13741 (N_13741,N_13120,N_13256);
or U13742 (N_13742,N_13381,N_13098);
and U13743 (N_13743,N_13369,N_13231);
and U13744 (N_13744,N_13266,N_13248);
or U13745 (N_13745,N_13162,N_13342);
or U13746 (N_13746,N_13017,N_13431);
nor U13747 (N_13747,N_13204,N_13453);
or U13748 (N_13748,N_13383,N_13215);
nor U13749 (N_13749,N_13432,N_13344);
nand U13750 (N_13750,N_13222,N_13477);
nor U13751 (N_13751,N_13169,N_13163);
xnor U13752 (N_13752,N_13229,N_13493);
or U13753 (N_13753,N_13358,N_13235);
nor U13754 (N_13754,N_13366,N_13222);
nor U13755 (N_13755,N_13055,N_13357);
nor U13756 (N_13756,N_13022,N_13106);
and U13757 (N_13757,N_13350,N_13321);
or U13758 (N_13758,N_13103,N_13358);
nand U13759 (N_13759,N_13488,N_13434);
nand U13760 (N_13760,N_13309,N_13161);
nor U13761 (N_13761,N_13498,N_13177);
and U13762 (N_13762,N_13415,N_13371);
or U13763 (N_13763,N_13386,N_13286);
nand U13764 (N_13764,N_13204,N_13222);
and U13765 (N_13765,N_13032,N_13018);
nand U13766 (N_13766,N_13022,N_13302);
and U13767 (N_13767,N_13190,N_13112);
nor U13768 (N_13768,N_13454,N_13314);
nand U13769 (N_13769,N_13499,N_13178);
and U13770 (N_13770,N_13144,N_13195);
nor U13771 (N_13771,N_13147,N_13088);
or U13772 (N_13772,N_13091,N_13292);
or U13773 (N_13773,N_13076,N_13432);
and U13774 (N_13774,N_13255,N_13086);
and U13775 (N_13775,N_13346,N_13145);
or U13776 (N_13776,N_13009,N_13131);
nand U13777 (N_13777,N_13052,N_13306);
and U13778 (N_13778,N_13008,N_13093);
nand U13779 (N_13779,N_13275,N_13407);
and U13780 (N_13780,N_13498,N_13020);
nor U13781 (N_13781,N_13214,N_13252);
or U13782 (N_13782,N_13017,N_13363);
and U13783 (N_13783,N_13307,N_13127);
nor U13784 (N_13784,N_13455,N_13128);
nand U13785 (N_13785,N_13300,N_13070);
nor U13786 (N_13786,N_13312,N_13421);
and U13787 (N_13787,N_13140,N_13384);
or U13788 (N_13788,N_13220,N_13002);
and U13789 (N_13789,N_13138,N_13007);
or U13790 (N_13790,N_13492,N_13170);
or U13791 (N_13791,N_13451,N_13092);
nor U13792 (N_13792,N_13144,N_13186);
and U13793 (N_13793,N_13141,N_13024);
or U13794 (N_13794,N_13463,N_13484);
or U13795 (N_13795,N_13241,N_13381);
nand U13796 (N_13796,N_13393,N_13352);
nor U13797 (N_13797,N_13294,N_13102);
and U13798 (N_13798,N_13418,N_13010);
or U13799 (N_13799,N_13170,N_13489);
nand U13800 (N_13800,N_13397,N_13058);
or U13801 (N_13801,N_13227,N_13278);
or U13802 (N_13802,N_13112,N_13212);
and U13803 (N_13803,N_13115,N_13162);
and U13804 (N_13804,N_13345,N_13207);
and U13805 (N_13805,N_13351,N_13092);
and U13806 (N_13806,N_13019,N_13259);
nand U13807 (N_13807,N_13119,N_13332);
nand U13808 (N_13808,N_13220,N_13459);
nor U13809 (N_13809,N_13402,N_13305);
and U13810 (N_13810,N_13355,N_13058);
or U13811 (N_13811,N_13112,N_13201);
or U13812 (N_13812,N_13133,N_13277);
or U13813 (N_13813,N_13029,N_13103);
and U13814 (N_13814,N_13337,N_13323);
and U13815 (N_13815,N_13370,N_13358);
and U13816 (N_13816,N_13053,N_13495);
nor U13817 (N_13817,N_13297,N_13324);
or U13818 (N_13818,N_13010,N_13027);
and U13819 (N_13819,N_13014,N_13298);
or U13820 (N_13820,N_13346,N_13148);
nand U13821 (N_13821,N_13302,N_13160);
nand U13822 (N_13822,N_13014,N_13488);
nor U13823 (N_13823,N_13135,N_13487);
and U13824 (N_13824,N_13380,N_13464);
or U13825 (N_13825,N_13492,N_13085);
nor U13826 (N_13826,N_13335,N_13268);
and U13827 (N_13827,N_13375,N_13373);
nand U13828 (N_13828,N_13044,N_13003);
nor U13829 (N_13829,N_13025,N_13035);
nand U13830 (N_13830,N_13447,N_13035);
nand U13831 (N_13831,N_13100,N_13448);
nand U13832 (N_13832,N_13438,N_13044);
nor U13833 (N_13833,N_13249,N_13179);
nor U13834 (N_13834,N_13473,N_13478);
and U13835 (N_13835,N_13291,N_13253);
or U13836 (N_13836,N_13417,N_13169);
nor U13837 (N_13837,N_13495,N_13239);
and U13838 (N_13838,N_13166,N_13427);
xor U13839 (N_13839,N_13207,N_13200);
nand U13840 (N_13840,N_13449,N_13024);
nand U13841 (N_13841,N_13396,N_13376);
and U13842 (N_13842,N_13053,N_13211);
nand U13843 (N_13843,N_13162,N_13393);
or U13844 (N_13844,N_13224,N_13042);
nand U13845 (N_13845,N_13475,N_13259);
nor U13846 (N_13846,N_13013,N_13266);
nor U13847 (N_13847,N_13333,N_13265);
xor U13848 (N_13848,N_13055,N_13098);
or U13849 (N_13849,N_13019,N_13434);
or U13850 (N_13850,N_13161,N_13384);
nor U13851 (N_13851,N_13170,N_13313);
nand U13852 (N_13852,N_13368,N_13259);
or U13853 (N_13853,N_13127,N_13115);
and U13854 (N_13854,N_13070,N_13322);
or U13855 (N_13855,N_13374,N_13212);
or U13856 (N_13856,N_13341,N_13413);
nand U13857 (N_13857,N_13415,N_13207);
or U13858 (N_13858,N_13454,N_13462);
and U13859 (N_13859,N_13084,N_13210);
nand U13860 (N_13860,N_13068,N_13268);
or U13861 (N_13861,N_13017,N_13085);
nor U13862 (N_13862,N_13342,N_13165);
and U13863 (N_13863,N_13127,N_13379);
and U13864 (N_13864,N_13067,N_13271);
nand U13865 (N_13865,N_13312,N_13083);
and U13866 (N_13866,N_13271,N_13367);
or U13867 (N_13867,N_13170,N_13360);
nor U13868 (N_13868,N_13418,N_13496);
or U13869 (N_13869,N_13184,N_13384);
or U13870 (N_13870,N_13126,N_13109);
xor U13871 (N_13871,N_13132,N_13265);
and U13872 (N_13872,N_13365,N_13151);
nand U13873 (N_13873,N_13335,N_13015);
nor U13874 (N_13874,N_13039,N_13343);
nand U13875 (N_13875,N_13217,N_13361);
nand U13876 (N_13876,N_13324,N_13299);
nor U13877 (N_13877,N_13140,N_13479);
nor U13878 (N_13878,N_13019,N_13255);
and U13879 (N_13879,N_13095,N_13337);
or U13880 (N_13880,N_13286,N_13403);
and U13881 (N_13881,N_13411,N_13393);
xnor U13882 (N_13882,N_13384,N_13273);
nor U13883 (N_13883,N_13496,N_13466);
nand U13884 (N_13884,N_13480,N_13481);
nand U13885 (N_13885,N_13121,N_13165);
or U13886 (N_13886,N_13045,N_13415);
and U13887 (N_13887,N_13397,N_13366);
or U13888 (N_13888,N_13074,N_13056);
and U13889 (N_13889,N_13027,N_13472);
or U13890 (N_13890,N_13358,N_13136);
or U13891 (N_13891,N_13308,N_13148);
nor U13892 (N_13892,N_13165,N_13354);
nand U13893 (N_13893,N_13326,N_13412);
nor U13894 (N_13894,N_13310,N_13482);
or U13895 (N_13895,N_13240,N_13073);
and U13896 (N_13896,N_13209,N_13484);
xnor U13897 (N_13897,N_13242,N_13405);
nand U13898 (N_13898,N_13438,N_13304);
and U13899 (N_13899,N_13037,N_13122);
nand U13900 (N_13900,N_13067,N_13084);
and U13901 (N_13901,N_13353,N_13153);
nand U13902 (N_13902,N_13063,N_13227);
and U13903 (N_13903,N_13433,N_13475);
and U13904 (N_13904,N_13158,N_13431);
or U13905 (N_13905,N_13424,N_13039);
nor U13906 (N_13906,N_13402,N_13018);
or U13907 (N_13907,N_13337,N_13273);
nor U13908 (N_13908,N_13020,N_13191);
or U13909 (N_13909,N_13383,N_13032);
nand U13910 (N_13910,N_13441,N_13241);
and U13911 (N_13911,N_13270,N_13455);
nor U13912 (N_13912,N_13061,N_13300);
nand U13913 (N_13913,N_13452,N_13070);
and U13914 (N_13914,N_13406,N_13113);
or U13915 (N_13915,N_13011,N_13479);
and U13916 (N_13916,N_13494,N_13387);
nor U13917 (N_13917,N_13264,N_13338);
and U13918 (N_13918,N_13321,N_13072);
and U13919 (N_13919,N_13238,N_13173);
or U13920 (N_13920,N_13445,N_13006);
nor U13921 (N_13921,N_13276,N_13009);
or U13922 (N_13922,N_13321,N_13124);
and U13923 (N_13923,N_13217,N_13061);
nand U13924 (N_13924,N_13459,N_13474);
nand U13925 (N_13925,N_13081,N_13392);
nand U13926 (N_13926,N_13018,N_13325);
nor U13927 (N_13927,N_13257,N_13307);
nor U13928 (N_13928,N_13495,N_13241);
nor U13929 (N_13929,N_13367,N_13283);
nor U13930 (N_13930,N_13342,N_13113);
nand U13931 (N_13931,N_13050,N_13348);
or U13932 (N_13932,N_13212,N_13123);
or U13933 (N_13933,N_13137,N_13027);
and U13934 (N_13934,N_13438,N_13411);
or U13935 (N_13935,N_13228,N_13498);
nand U13936 (N_13936,N_13072,N_13225);
and U13937 (N_13937,N_13308,N_13398);
nor U13938 (N_13938,N_13288,N_13264);
or U13939 (N_13939,N_13051,N_13108);
and U13940 (N_13940,N_13316,N_13224);
or U13941 (N_13941,N_13499,N_13090);
nand U13942 (N_13942,N_13256,N_13183);
nand U13943 (N_13943,N_13349,N_13211);
and U13944 (N_13944,N_13029,N_13114);
or U13945 (N_13945,N_13400,N_13121);
and U13946 (N_13946,N_13154,N_13466);
nand U13947 (N_13947,N_13447,N_13101);
nand U13948 (N_13948,N_13305,N_13193);
and U13949 (N_13949,N_13120,N_13042);
nand U13950 (N_13950,N_13211,N_13241);
nand U13951 (N_13951,N_13419,N_13307);
and U13952 (N_13952,N_13219,N_13475);
and U13953 (N_13953,N_13304,N_13180);
xor U13954 (N_13954,N_13474,N_13218);
or U13955 (N_13955,N_13335,N_13072);
or U13956 (N_13956,N_13151,N_13282);
nor U13957 (N_13957,N_13209,N_13117);
nand U13958 (N_13958,N_13397,N_13225);
nand U13959 (N_13959,N_13344,N_13494);
or U13960 (N_13960,N_13194,N_13002);
nand U13961 (N_13961,N_13085,N_13219);
nand U13962 (N_13962,N_13496,N_13357);
nor U13963 (N_13963,N_13332,N_13045);
and U13964 (N_13964,N_13231,N_13459);
and U13965 (N_13965,N_13325,N_13125);
or U13966 (N_13966,N_13027,N_13148);
nand U13967 (N_13967,N_13373,N_13059);
nor U13968 (N_13968,N_13239,N_13197);
and U13969 (N_13969,N_13234,N_13148);
or U13970 (N_13970,N_13477,N_13004);
and U13971 (N_13971,N_13439,N_13312);
nor U13972 (N_13972,N_13498,N_13453);
or U13973 (N_13973,N_13095,N_13255);
nand U13974 (N_13974,N_13172,N_13135);
xor U13975 (N_13975,N_13234,N_13362);
or U13976 (N_13976,N_13022,N_13446);
nand U13977 (N_13977,N_13480,N_13363);
nor U13978 (N_13978,N_13311,N_13342);
and U13979 (N_13979,N_13164,N_13381);
nand U13980 (N_13980,N_13443,N_13473);
or U13981 (N_13981,N_13347,N_13358);
or U13982 (N_13982,N_13352,N_13424);
or U13983 (N_13983,N_13203,N_13348);
and U13984 (N_13984,N_13471,N_13113);
and U13985 (N_13985,N_13401,N_13193);
nand U13986 (N_13986,N_13358,N_13279);
or U13987 (N_13987,N_13062,N_13013);
and U13988 (N_13988,N_13452,N_13461);
nand U13989 (N_13989,N_13480,N_13163);
nor U13990 (N_13990,N_13082,N_13363);
nand U13991 (N_13991,N_13019,N_13395);
nor U13992 (N_13992,N_13014,N_13158);
or U13993 (N_13993,N_13452,N_13288);
or U13994 (N_13994,N_13456,N_13332);
or U13995 (N_13995,N_13445,N_13113);
or U13996 (N_13996,N_13095,N_13233);
nand U13997 (N_13997,N_13104,N_13296);
nor U13998 (N_13998,N_13430,N_13361);
nor U13999 (N_13999,N_13069,N_13372);
nor U14000 (N_14000,N_13543,N_13799);
or U14001 (N_14001,N_13531,N_13953);
and U14002 (N_14002,N_13541,N_13998);
nand U14003 (N_14003,N_13978,N_13704);
nand U14004 (N_14004,N_13602,N_13701);
or U14005 (N_14005,N_13526,N_13837);
and U14006 (N_14006,N_13950,N_13999);
and U14007 (N_14007,N_13776,N_13994);
or U14008 (N_14008,N_13655,N_13935);
nor U14009 (N_14009,N_13598,N_13943);
nor U14010 (N_14010,N_13840,N_13679);
or U14011 (N_14011,N_13795,N_13737);
nor U14012 (N_14012,N_13565,N_13981);
nor U14013 (N_14013,N_13549,N_13609);
or U14014 (N_14014,N_13832,N_13826);
and U14015 (N_14015,N_13607,N_13592);
or U14016 (N_14016,N_13856,N_13848);
nor U14017 (N_14017,N_13570,N_13977);
nand U14018 (N_14018,N_13673,N_13796);
or U14019 (N_14019,N_13610,N_13867);
or U14020 (N_14020,N_13813,N_13545);
nor U14021 (N_14021,N_13616,N_13846);
nand U14022 (N_14022,N_13523,N_13972);
nor U14023 (N_14023,N_13730,N_13926);
nand U14024 (N_14024,N_13951,N_13783);
nand U14025 (N_14025,N_13642,N_13690);
or U14026 (N_14026,N_13939,N_13591);
and U14027 (N_14027,N_13711,N_13747);
nand U14028 (N_14028,N_13877,N_13718);
or U14029 (N_14029,N_13640,N_13868);
or U14030 (N_14030,N_13965,N_13924);
nand U14031 (N_14031,N_13956,N_13736);
nand U14032 (N_14032,N_13741,N_13585);
nand U14033 (N_14033,N_13643,N_13656);
nand U14034 (N_14034,N_13993,N_13819);
nor U14035 (N_14035,N_13768,N_13902);
nand U14036 (N_14036,N_13560,N_13687);
nand U14037 (N_14037,N_13641,N_13705);
and U14038 (N_14038,N_13725,N_13806);
nor U14039 (N_14039,N_13734,N_13786);
or U14040 (N_14040,N_13880,N_13992);
and U14041 (N_14041,N_13727,N_13574);
and U14042 (N_14042,N_13818,N_13780);
nand U14043 (N_14043,N_13594,N_13986);
nor U14044 (N_14044,N_13859,N_13851);
nand U14045 (N_14045,N_13675,N_13692);
nand U14046 (N_14046,N_13534,N_13723);
or U14047 (N_14047,N_13724,N_13653);
and U14048 (N_14048,N_13893,N_13948);
nand U14049 (N_14049,N_13683,N_13661);
nand U14050 (N_14050,N_13581,N_13710);
and U14051 (N_14051,N_13929,N_13630);
nand U14052 (N_14052,N_13546,N_13984);
nand U14053 (N_14053,N_13794,N_13936);
or U14054 (N_14054,N_13513,N_13589);
xnor U14055 (N_14055,N_13932,N_13595);
nor U14056 (N_14056,N_13587,N_13918);
nor U14057 (N_14057,N_13674,N_13666);
or U14058 (N_14058,N_13904,N_13584);
or U14059 (N_14059,N_13652,N_13945);
nand U14060 (N_14060,N_13812,N_13957);
nor U14061 (N_14061,N_13831,N_13510);
nor U14062 (N_14062,N_13588,N_13599);
nor U14063 (N_14063,N_13878,N_13760);
or U14064 (N_14064,N_13561,N_13586);
nand U14065 (N_14065,N_13572,N_13919);
nand U14066 (N_14066,N_13767,N_13600);
or U14067 (N_14067,N_13562,N_13608);
or U14068 (N_14068,N_13664,N_13920);
nand U14069 (N_14069,N_13973,N_13805);
or U14070 (N_14070,N_13772,N_13928);
nor U14071 (N_14071,N_13961,N_13964);
nand U14072 (N_14072,N_13931,N_13915);
and U14073 (N_14073,N_13744,N_13644);
or U14074 (N_14074,N_13763,N_13810);
or U14075 (N_14075,N_13621,N_13770);
xor U14076 (N_14076,N_13825,N_13921);
nor U14077 (N_14077,N_13847,N_13971);
or U14078 (N_14078,N_13693,N_13532);
and U14079 (N_14079,N_13548,N_13686);
nand U14080 (N_14080,N_13942,N_13991);
or U14081 (N_14081,N_13547,N_13703);
xnor U14082 (N_14082,N_13870,N_13885);
nand U14083 (N_14083,N_13959,N_13952);
and U14084 (N_14084,N_13726,N_13521);
or U14085 (N_14085,N_13540,N_13835);
and U14086 (N_14086,N_13804,N_13782);
nor U14087 (N_14087,N_13754,N_13769);
or U14088 (N_14088,N_13612,N_13564);
nor U14089 (N_14089,N_13974,N_13892);
nor U14090 (N_14090,N_13535,N_13544);
nand U14091 (N_14091,N_13755,N_13891);
nor U14092 (N_14092,N_13901,N_13910);
nand U14093 (N_14093,N_13707,N_13504);
nand U14094 (N_14094,N_13721,N_13728);
nand U14095 (N_14095,N_13751,N_13750);
nor U14096 (N_14096,N_13551,N_13646);
and U14097 (N_14097,N_13636,N_13712);
or U14098 (N_14098,N_13735,N_13759);
nor U14099 (N_14099,N_13719,N_13625);
and U14100 (N_14100,N_13722,N_13648);
and U14101 (N_14101,N_13963,N_13527);
nor U14102 (N_14102,N_13514,N_13862);
nor U14103 (N_14103,N_13708,N_13842);
or U14104 (N_14104,N_13511,N_13808);
or U14105 (N_14105,N_13872,N_13659);
nor U14106 (N_14106,N_13863,N_13528);
nor U14107 (N_14107,N_13605,N_13619);
nor U14108 (N_14108,N_13784,N_13916);
nand U14109 (N_14109,N_13658,N_13903);
xor U14110 (N_14110,N_13669,N_13512);
xor U14111 (N_14111,N_13700,N_13828);
or U14112 (N_14112,N_13895,N_13756);
or U14113 (N_14113,N_13777,N_13732);
or U14114 (N_14114,N_13567,N_13855);
nand U14115 (N_14115,N_13522,N_13601);
nand U14116 (N_14116,N_13717,N_13580);
and U14117 (N_14117,N_13678,N_13634);
nor U14118 (N_14118,N_13883,N_13890);
nand U14119 (N_14119,N_13740,N_13906);
and U14120 (N_14120,N_13573,N_13762);
nor U14121 (N_14121,N_13614,N_13876);
nor U14122 (N_14122,N_13995,N_13729);
nand U14123 (N_14123,N_13817,N_13766);
nor U14124 (N_14124,N_13888,N_13507);
nor U14125 (N_14125,N_13542,N_13749);
nand U14126 (N_14126,N_13628,N_13829);
and U14127 (N_14127,N_13887,N_13923);
nand U14128 (N_14128,N_13623,N_13566);
and U14129 (N_14129,N_13650,N_13898);
nand U14130 (N_14130,N_13590,N_13550);
nor U14131 (N_14131,N_13871,N_13603);
nand U14132 (N_14132,N_13637,N_13866);
nand U14133 (N_14133,N_13861,N_13765);
nor U14134 (N_14134,N_13660,N_13533);
or U14135 (N_14135,N_13873,N_13520);
and U14136 (N_14136,N_13997,N_13934);
or U14137 (N_14137,N_13823,N_13685);
and U14138 (N_14138,N_13559,N_13716);
or U14139 (N_14139,N_13954,N_13793);
nand U14140 (N_14140,N_13654,N_13731);
nor U14141 (N_14141,N_13820,N_13622);
or U14142 (N_14142,N_13938,N_13501);
and U14143 (N_14143,N_13774,N_13665);
xor U14144 (N_14144,N_13790,N_13852);
nand U14145 (N_14145,N_13518,N_13684);
nand U14146 (N_14146,N_13814,N_13631);
and U14147 (N_14147,N_13982,N_13967);
and U14148 (N_14148,N_13989,N_13975);
and U14149 (N_14149,N_13530,N_13517);
and U14150 (N_14150,N_13983,N_13937);
nor U14151 (N_14151,N_13836,N_13638);
nand U14152 (N_14152,N_13671,N_13881);
nand U14153 (N_14153,N_13663,N_13899);
nor U14154 (N_14154,N_13645,N_13557);
nor U14155 (N_14155,N_13801,N_13715);
or U14156 (N_14156,N_13917,N_13912);
and U14157 (N_14157,N_13583,N_13875);
nand U14158 (N_14158,N_13976,N_13537);
nand U14159 (N_14159,N_13787,N_13670);
nor U14160 (N_14160,N_13913,N_13985);
nor U14161 (N_14161,N_13955,N_13778);
nor U14162 (N_14162,N_13761,N_13933);
and U14163 (N_14163,N_13558,N_13988);
or U14164 (N_14164,N_13834,N_13742);
nor U14165 (N_14165,N_13713,N_13706);
or U14166 (N_14166,N_13925,N_13830);
and U14167 (N_14167,N_13627,N_13694);
and U14168 (N_14168,N_13516,N_13552);
nor U14169 (N_14169,N_13958,N_13940);
nor U14170 (N_14170,N_13941,N_13811);
nor U14171 (N_14171,N_13629,N_13563);
and U14172 (N_14172,N_13839,N_13709);
or U14173 (N_14173,N_13779,N_13695);
nor U14174 (N_14174,N_13905,N_13889);
or U14175 (N_14175,N_13894,N_13968);
nand U14176 (N_14176,N_13879,N_13886);
nor U14177 (N_14177,N_13815,N_13822);
and U14178 (N_14178,N_13529,N_13896);
and U14179 (N_14179,N_13539,N_13858);
or U14180 (N_14180,N_13569,N_13946);
nand U14181 (N_14181,N_13947,N_13843);
nor U14182 (N_14182,N_13792,N_13927);
nor U14183 (N_14183,N_13509,N_13618);
nand U14184 (N_14184,N_13672,N_13688);
and U14185 (N_14185,N_13752,N_13575);
nand U14186 (N_14186,N_13809,N_13606);
or U14187 (N_14187,N_13647,N_13980);
or U14188 (N_14188,N_13508,N_13775);
or U14189 (N_14189,N_13554,N_13738);
and U14190 (N_14190,N_13816,N_13908);
and U14191 (N_14191,N_13668,N_13733);
nand U14192 (N_14192,N_13914,N_13930);
nand U14193 (N_14193,N_13966,N_13969);
nor U14194 (N_14194,N_13613,N_13500);
nor U14195 (N_14195,N_13911,N_13604);
nand U14196 (N_14196,N_13699,N_13773);
or U14197 (N_14197,N_13536,N_13745);
or U14198 (N_14198,N_13597,N_13691);
nand U14199 (N_14199,N_13502,N_13857);
and U14200 (N_14200,N_13624,N_13757);
or U14201 (N_14201,N_13781,N_13748);
or U14202 (N_14202,N_13571,N_13785);
nor U14203 (N_14203,N_13576,N_13807);
and U14204 (N_14204,N_13556,N_13578);
nand U14205 (N_14205,N_13525,N_13802);
nor U14206 (N_14206,N_13900,N_13680);
nand U14207 (N_14207,N_13962,N_13667);
xnor U14208 (N_14208,N_13789,N_13821);
or U14209 (N_14209,N_13844,N_13702);
or U14210 (N_14210,N_13860,N_13698);
or U14211 (N_14211,N_13696,N_13996);
and U14212 (N_14212,N_13970,N_13791);
nand U14213 (N_14213,N_13681,N_13949);
and U14214 (N_14214,N_13798,N_13596);
or U14215 (N_14215,N_13990,N_13909);
nor U14216 (N_14216,N_13635,N_13626);
and U14217 (N_14217,N_13649,N_13676);
and U14218 (N_14218,N_13897,N_13662);
and U14219 (N_14219,N_13582,N_13746);
nand U14220 (N_14220,N_13803,N_13771);
and U14221 (N_14221,N_13651,N_13850);
nor U14222 (N_14222,N_13505,N_13845);
nor U14223 (N_14223,N_13800,N_13884);
nand U14224 (N_14224,N_13593,N_13579);
or U14225 (N_14225,N_13519,N_13714);
nor U14226 (N_14226,N_13689,N_13849);
or U14227 (N_14227,N_13833,N_13907);
or U14228 (N_14228,N_13788,N_13944);
nor U14229 (N_14229,N_13853,N_13506);
or U14230 (N_14230,N_13743,N_13854);
and U14231 (N_14231,N_13617,N_13555);
nor U14232 (N_14232,N_13865,N_13987);
or U14233 (N_14233,N_13657,N_13758);
nor U14234 (N_14234,N_13864,N_13568);
nor U14235 (N_14235,N_13515,N_13697);
and U14236 (N_14236,N_13827,N_13882);
and U14237 (N_14237,N_13922,N_13869);
nor U14238 (N_14238,N_13632,N_13538);
nand U14239 (N_14239,N_13764,N_13553);
nor U14240 (N_14240,N_13577,N_13753);
and U14241 (N_14241,N_13611,N_13639);
nand U14242 (N_14242,N_13524,N_13677);
or U14243 (N_14243,N_13797,N_13838);
and U14244 (N_14244,N_13615,N_13841);
and U14245 (N_14245,N_13874,N_13960);
nand U14246 (N_14246,N_13503,N_13739);
or U14247 (N_14247,N_13620,N_13682);
and U14248 (N_14248,N_13633,N_13824);
and U14249 (N_14249,N_13979,N_13720);
nor U14250 (N_14250,N_13580,N_13978);
nor U14251 (N_14251,N_13957,N_13924);
nor U14252 (N_14252,N_13879,N_13767);
and U14253 (N_14253,N_13715,N_13523);
nor U14254 (N_14254,N_13831,N_13939);
and U14255 (N_14255,N_13745,N_13579);
and U14256 (N_14256,N_13783,N_13656);
nor U14257 (N_14257,N_13629,N_13554);
nor U14258 (N_14258,N_13723,N_13601);
nand U14259 (N_14259,N_13607,N_13998);
or U14260 (N_14260,N_13894,N_13781);
nand U14261 (N_14261,N_13843,N_13988);
nor U14262 (N_14262,N_13613,N_13716);
and U14263 (N_14263,N_13944,N_13521);
nor U14264 (N_14264,N_13689,N_13918);
nor U14265 (N_14265,N_13989,N_13780);
nor U14266 (N_14266,N_13684,N_13736);
nor U14267 (N_14267,N_13518,N_13923);
xnor U14268 (N_14268,N_13889,N_13626);
nor U14269 (N_14269,N_13652,N_13977);
nand U14270 (N_14270,N_13772,N_13877);
or U14271 (N_14271,N_13641,N_13969);
and U14272 (N_14272,N_13808,N_13740);
and U14273 (N_14273,N_13724,N_13537);
nor U14274 (N_14274,N_13618,N_13657);
nor U14275 (N_14275,N_13653,N_13801);
nor U14276 (N_14276,N_13751,N_13960);
or U14277 (N_14277,N_13822,N_13717);
nor U14278 (N_14278,N_13623,N_13621);
and U14279 (N_14279,N_13533,N_13608);
or U14280 (N_14280,N_13665,N_13830);
and U14281 (N_14281,N_13992,N_13877);
or U14282 (N_14282,N_13755,N_13680);
nand U14283 (N_14283,N_13833,N_13905);
or U14284 (N_14284,N_13533,N_13676);
nor U14285 (N_14285,N_13741,N_13651);
nand U14286 (N_14286,N_13761,N_13823);
xnor U14287 (N_14287,N_13706,N_13768);
and U14288 (N_14288,N_13975,N_13893);
nor U14289 (N_14289,N_13840,N_13623);
nand U14290 (N_14290,N_13684,N_13635);
nor U14291 (N_14291,N_13597,N_13995);
or U14292 (N_14292,N_13962,N_13749);
and U14293 (N_14293,N_13844,N_13858);
nor U14294 (N_14294,N_13756,N_13849);
nand U14295 (N_14295,N_13632,N_13511);
nor U14296 (N_14296,N_13629,N_13923);
and U14297 (N_14297,N_13633,N_13657);
nand U14298 (N_14298,N_13522,N_13898);
nand U14299 (N_14299,N_13825,N_13518);
nor U14300 (N_14300,N_13643,N_13646);
nand U14301 (N_14301,N_13638,N_13897);
and U14302 (N_14302,N_13746,N_13962);
and U14303 (N_14303,N_13785,N_13592);
nor U14304 (N_14304,N_13970,N_13815);
and U14305 (N_14305,N_13755,N_13807);
and U14306 (N_14306,N_13746,N_13917);
nand U14307 (N_14307,N_13817,N_13606);
nand U14308 (N_14308,N_13732,N_13884);
xor U14309 (N_14309,N_13695,N_13994);
or U14310 (N_14310,N_13572,N_13527);
nor U14311 (N_14311,N_13921,N_13798);
nand U14312 (N_14312,N_13967,N_13929);
nor U14313 (N_14313,N_13920,N_13578);
nor U14314 (N_14314,N_13537,N_13527);
and U14315 (N_14315,N_13512,N_13556);
and U14316 (N_14316,N_13532,N_13845);
or U14317 (N_14317,N_13593,N_13879);
or U14318 (N_14318,N_13827,N_13593);
nand U14319 (N_14319,N_13743,N_13584);
nand U14320 (N_14320,N_13523,N_13924);
and U14321 (N_14321,N_13576,N_13787);
nor U14322 (N_14322,N_13998,N_13688);
nor U14323 (N_14323,N_13978,N_13995);
or U14324 (N_14324,N_13900,N_13951);
nor U14325 (N_14325,N_13900,N_13788);
nor U14326 (N_14326,N_13639,N_13532);
nand U14327 (N_14327,N_13902,N_13803);
or U14328 (N_14328,N_13922,N_13521);
and U14329 (N_14329,N_13767,N_13575);
nand U14330 (N_14330,N_13852,N_13514);
nor U14331 (N_14331,N_13577,N_13661);
nand U14332 (N_14332,N_13858,N_13737);
or U14333 (N_14333,N_13762,N_13716);
and U14334 (N_14334,N_13639,N_13843);
or U14335 (N_14335,N_13545,N_13620);
nor U14336 (N_14336,N_13944,N_13672);
nand U14337 (N_14337,N_13709,N_13637);
nor U14338 (N_14338,N_13690,N_13717);
and U14339 (N_14339,N_13674,N_13996);
and U14340 (N_14340,N_13606,N_13974);
nor U14341 (N_14341,N_13778,N_13779);
or U14342 (N_14342,N_13608,N_13952);
nor U14343 (N_14343,N_13777,N_13575);
nor U14344 (N_14344,N_13504,N_13851);
or U14345 (N_14345,N_13927,N_13545);
and U14346 (N_14346,N_13626,N_13959);
and U14347 (N_14347,N_13506,N_13637);
or U14348 (N_14348,N_13910,N_13953);
nor U14349 (N_14349,N_13985,N_13576);
or U14350 (N_14350,N_13982,N_13899);
nor U14351 (N_14351,N_13644,N_13990);
and U14352 (N_14352,N_13882,N_13971);
nand U14353 (N_14353,N_13843,N_13538);
nand U14354 (N_14354,N_13937,N_13801);
nand U14355 (N_14355,N_13810,N_13933);
or U14356 (N_14356,N_13738,N_13794);
nor U14357 (N_14357,N_13568,N_13916);
nand U14358 (N_14358,N_13583,N_13611);
or U14359 (N_14359,N_13598,N_13872);
nor U14360 (N_14360,N_13780,N_13748);
and U14361 (N_14361,N_13727,N_13545);
xnor U14362 (N_14362,N_13754,N_13782);
and U14363 (N_14363,N_13704,N_13558);
nor U14364 (N_14364,N_13501,N_13652);
or U14365 (N_14365,N_13885,N_13851);
nand U14366 (N_14366,N_13958,N_13598);
and U14367 (N_14367,N_13529,N_13867);
or U14368 (N_14368,N_13554,N_13680);
or U14369 (N_14369,N_13828,N_13996);
and U14370 (N_14370,N_13726,N_13580);
nor U14371 (N_14371,N_13794,N_13968);
xnor U14372 (N_14372,N_13851,N_13630);
or U14373 (N_14373,N_13666,N_13899);
or U14374 (N_14374,N_13796,N_13913);
nor U14375 (N_14375,N_13655,N_13625);
nand U14376 (N_14376,N_13772,N_13597);
or U14377 (N_14377,N_13634,N_13924);
and U14378 (N_14378,N_13998,N_13674);
nand U14379 (N_14379,N_13515,N_13966);
nand U14380 (N_14380,N_13523,N_13958);
nor U14381 (N_14381,N_13761,N_13840);
and U14382 (N_14382,N_13621,N_13622);
and U14383 (N_14383,N_13840,N_13630);
nor U14384 (N_14384,N_13572,N_13750);
nor U14385 (N_14385,N_13719,N_13536);
nand U14386 (N_14386,N_13937,N_13580);
or U14387 (N_14387,N_13676,N_13696);
and U14388 (N_14388,N_13889,N_13756);
nand U14389 (N_14389,N_13796,N_13777);
and U14390 (N_14390,N_13859,N_13871);
nand U14391 (N_14391,N_13506,N_13857);
and U14392 (N_14392,N_13666,N_13999);
nor U14393 (N_14393,N_13734,N_13528);
and U14394 (N_14394,N_13782,N_13785);
and U14395 (N_14395,N_13656,N_13574);
nand U14396 (N_14396,N_13616,N_13998);
nand U14397 (N_14397,N_13906,N_13886);
or U14398 (N_14398,N_13655,N_13721);
and U14399 (N_14399,N_13836,N_13821);
nand U14400 (N_14400,N_13626,N_13634);
or U14401 (N_14401,N_13667,N_13825);
nor U14402 (N_14402,N_13615,N_13851);
xor U14403 (N_14403,N_13987,N_13840);
and U14404 (N_14404,N_13720,N_13746);
nand U14405 (N_14405,N_13972,N_13543);
nand U14406 (N_14406,N_13900,N_13938);
or U14407 (N_14407,N_13710,N_13793);
nor U14408 (N_14408,N_13990,N_13889);
and U14409 (N_14409,N_13927,N_13743);
or U14410 (N_14410,N_13924,N_13569);
or U14411 (N_14411,N_13954,N_13929);
and U14412 (N_14412,N_13505,N_13970);
nand U14413 (N_14413,N_13969,N_13508);
and U14414 (N_14414,N_13841,N_13836);
or U14415 (N_14415,N_13698,N_13521);
or U14416 (N_14416,N_13514,N_13807);
or U14417 (N_14417,N_13956,N_13997);
nor U14418 (N_14418,N_13756,N_13950);
and U14419 (N_14419,N_13844,N_13801);
and U14420 (N_14420,N_13812,N_13977);
and U14421 (N_14421,N_13881,N_13716);
and U14422 (N_14422,N_13839,N_13686);
and U14423 (N_14423,N_13835,N_13595);
and U14424 (N_14424,N_13853,N_13809);
or U14425 (N_14425,N_13911,N_13694);
and U14426 (N_14426,N_13581,N_13968);
or U14427 (N_14427,N_13729,N_13590);
nand U14428 (N_14428,N_13536,N_13679);
nor U14429 (N_14429,N_13872,N_13695);
or U14430 (N_14430,N_13635,N_13876);
or U14431 (N_14431,N_13610,N_13842);
and U14432 (N_14432,N_13997,N_13906);
or U14433 (N_14433,N_13643,N_13827);
and U14434 (N_14434,N_13975,N_13887);
or U14435 (N_14435,N_13840,N_13822);
nand U14436 (N_14436,N_13892,N_13845);
and U14437 (N_14437,N_13537,N_13857);
nand U14438 (N_14438,N_13833,N_13519);
nand U14439 (N_14439,N_13968,N_13704);
nor U14440 (N_14440,N_13919,N_13726);
and U14441 (N_14441,N_13624,N_13878);
nor U14442 (N_14442,N_13540,N_13699);
xnor U14443 (N_14443,N_13764,N_13538);
nand U14444 (N_14444,N_13848,N_13930);
and U14445 (N_14445,N_13899,N_13830);
nor U14446 (N_14446,N_13615,N_13647);
nand U14447 (N_14447,N_13703,N_13914);
nand U14448 (N_14448,N_13823,N_13665);
nor U14449 (N_14449,N_13734,N_13828);
xnor U14450 (N_14450,N_13654,N_13544);
and U14451 (N_14451,N_13632,N_13640);
and U14452 (N_14452,N_13600,N_13539);
or U14453 (N_14453,N_13701,N_13632);
nor U14454 (N_14454,N_13933,N_13734);
or U14455 (N_14455,N_13700,N_13972);
or U14456 (N_14456,N_13889,N_13677);
nand U14457 (N_14457,N_13957,N_13943);
nor U14458 (N_14458,N_13955,N_13520);
and U14459 (N_14459,N_13665,N_13519);
nand U14460 (N_14460,N_13837,N_13620);
or U14461 (N_14461,N_13616,N_13551);
or U14462 (N_14462,N_13577,N_13601);
nor U14463 (N_14463,N_13636,N_13585);
nand U14464 (N_14464,N_13944,N_13870);
or U14465 (N_14465,N_13768,N_13569);
nor U14466 (N_14466,N_13575,N_13917);
or U14467 (N_14467,N_13634,N_13816);
nor U14468 (N_14468,N_13922,N_13700);
and U14469 (N_14469,N_13712,N_13547);
and U14470 (N_14470,N_13933,N_13851);
and U14471 (N_14471,N_13625,N_13609);
or U14472 (N_14472,N_13618,N_13549);
nand U14473 (N_14473,N_13519,N_13982);
nand U14474 (N_14474,N_13595,N_13646);
nand U14475 (N_14475,N_13516,N_13542);
nor U14476 (N_14476,N_13673,N_13980);
or U14477 (N_14477,N_13810,N_13607);
nor U14478 (N_14478,N_13759,N_13990);
or U14479 (N_14479,N_13544,N_13649);
nand U14480 (N_14480,N_13831,N_13506);
nor U14481 (N_14481,N_13904,N_13532);
nor U14482 (N_14482,N_13848,N_13810);
nand U14483 (N_14483,N_13515,N_13580);
nand U14484 (N_14484,N_13785,N_13534);
and U14485 (N_14485,N_13874,N_13611);
nor U14486 (N_14486,N_13514,N_13647);
nor U14487 (N_14487,N_13775,N_13584);
and U14488 (N_14488,N_13960,N_13908);
and U14489 (N_14489,N_13754,N_13637);
or U14490 (N_14490,N_13542,N_13555);
nand U14491 (N_14491,N_13634,N_13853);
nand U14492 (N_14492,N_13749,N_13859);
or U14493 (N_14493,N_13678,N_13546);
and U14494 (N_14494,N_13783,N_13778);
and U14495 (N_14495,N_13552,N_13824);
nand U14496 (N_14496,N_13908,N_13860);
nor U14497 (N_14497,N_13702,N_13712);
nor U14498 (N_14498,N_13598,N_13636);
nand U14499 (N_14499,N_13961,N_13707);
and U14500 (N_14500,N_14253,N_14421);
nor U14501 (N_14501,N_14234,N_14211);
and U14502 (N_14502,N_14056,N_14348);
nor U14503 (N_14503,N_14210,N_14424);
nand U14504 (N_14504,N_14046,N_14302);
and U14505 (N_14505,N_14237,N_14411);
nor U14506 (N_14506,N_14485,N_14361);
nand U14507 (N_14507,N_14216,N_14468);
nor U14508 (N_14508,N_14489,N_14274);
and U14509 (N_14509,N_14410,N_14183);
nand U14510 (N_14510,N_14231,N_14435);
nor U14511 (N_14511,N_14197,N_14202);
nand U14512 (N_14512,N_14493,N_14409);
and U14513 (N_14513,N_14205,N_14329);
and U14514 (N_14514,N_14073,N_14428);
nand U14515 (N_14515,N_14229,N_14219);
nand U14516 (N_14516,N_14037,N_14288);
and U14517 (N_14517,N_14173,N_14097);
nand U14518 (N_14518,N_14133,N_14232);
nand U14519 (N_14519,N_14137,N_14112);
or U14520 (N_14520,N_14284,N_14289);
and U14521 (N_14521,N_14432,N_14151);
nor U14522 (N_14522,N_14312,N_14221);
xor U14523 (N_14523,N_14095,N_14327);
or U14524 (N_14524,N_14271,N_14474);
and U14525 (N_14525,N_14132,N_14047);
nand U14526 (N_14526,N_14248,N_14399);
or U14527 (N_14527,N_14473,N_14308);
nor U14528 (N_14528,N_14490,N_14142);
or U14529 (N_14529,N_14452,N_14094);
nor U14530 (N_14530,N_14355,N_14012);
and U14531 (N_14531,N_14444,N_14093);
and U14532 (N_14532,N_14321,N_14195);
nand U14533 (N_14533,N_14344,N_14125);
nand U14534 (N_14534,N_14225,N_14260);
nor U14535 (N_14535,N_14446,N_14364);
and U14536 (N_14536,N_14077,N_14157);
and U14537 (N_14537,N_14465,N_14486);
and U14538 (N_14538,N_14401,N_14051);
and U14539 (N_14539,N_14438,N_14005);
or U14540 (N_14540,N_14346,N_14412);
and U14541 (N_14541,N_14144,N_14086);
nor U14542 (N_14542,N_14407,N_14109);
and U14543 (N_14543,N_14298,N_14362);
nor U14544 (N_14544,N_14233,N_14480);
nand U14545 (N_14545,N_14007,N_14196);
and U14546 (N_14546,N_14460,N_14251);
nor U14547 (N_14547,N_14273,N_14240);
and U14548 (N_14548,N_14416,N_14224);
or U14549 (N_14549,N_14266,N_14050);
or U14550 (N_14550,N_14207,N_14246);
nor U14551 (N_14551,N_14105,N_14127);
nand U14552 (N_14552,N_14040,N_14376);
xnor U14553 (N_14553,N_14322,N_14433);
and U14554 (N_14554,N_14034,N_14400);
nor U14555 (N_14555,N_14179,N_14429);
nor U14556 (N_14556,N_14472,N_14345);
and U14557 (N_14557,N_14031,N_14128);
and U14558 (N_14558,N_14186,N_14120);
or U14559 (N_14559,N_14100,N_14140);
or U14560 (N_14560,N_14264,N_14134);
and U14561 (N_14561,N_14098,N_14442);
or U14562 (N_14562,N_14358,N_14417);
or U14563 (N_14563,N_14340,N_14153);
nor U14564 (N_14564,N_14124,N_14415);
nor U14565 (N_14565,N_14278,N_14038);
nor U14566 (N_14566,N_14019,N_14218);
nor U14567 (N_14567,N_14061,N_14152);
or U14568 (N_14568,N_14117,N_14369);
or U14569 (N_14569,N_14377,N_14239);
and U14570 (N_14570,N_14022,N_14135);
nand U14571 (N_14571,N_14041,N_14226);
nand U14572 (N_14572,N_14074,N_14174);
nor U14573 (N_14573,N_14150,N_14083);
nand U14574 (N_14574,N_14108,N_14395);
or U14575 (N_14575,N_14430,N_14420);
nor U14576 (N_14576,N_14043,N_14350);
and U14577 (N_14577,N_14475,N_14497);
nand U14578 (N_14578,N_14491,N_14423);
or U14579 (N_14579,N_14367,N_14147);
or U14580 (N_14580,N_14082,N_14060);
and U14581 (N_14581,N_14089,N_14070);
or U14582 (N_14582,N_14326,N_14425);
and U14583 (N_14583,N_14275,N_14102);
or U14584 (N_14584,N_14148,N_14198);
nand U14585 (N_14585,N_14126,N_14352);
nor U14586 (N_14586,N_14011,N_14431);
nand U14587 (N_14587,N_14213,N_14470);
and U14588 (N_14588,N_14455,N_14299);
or U14589 (N_14589,N_14319,N_14182);
and U14590 (N_14590,N_14055,N_14335);
and U14591 (N_14591,N_14437,N_14334);
and U14592 (N_14592,N_14149,N_14008);
or U14593 (N_14593,N_14014,N_14466);
nor U14594 (N_14594,N_14293,N_14027);
or U14595 (N_14595,N_14408,N_14405);
and U14596 (N_14596,N_14227,N_14208);
nand U14597 (N_14597,N_14013,N_14110);
or U14598 (N_14598,N_14230,N_14018);
and U14599 (N_14599,N_14010,N_14178);
nand U14600 (N_14600,N_14249,N_14309);
or U14601 (N_14601,N_14297,N_14192);
nand U14602 (N_14602,N_14080,N_14016);
nor U14603 (N_14603,N_14366,N_14397);
nand U14604 (N_14604,N_14262,N_14305);
nor U14605 (N_14605,N_14068,N_14169);
nor U14606 (N_14606,N_14347,N_14467);
or U14607 (N_14607,N_14270,N_14081);
nand U14608 (N_14608,N_14447,N_14045);
or U14609 (N_14609,N_14206,N_14156);
or U14610 (N_14610,N_14277,N_14296);
or U14611 (N_14611,N_14009,N_14357);
nor U14612 (N_14612,N_14184,N_14311);
or U14613 (N_14613,N_14252,N_14382);
nand U14614 (N_14614,N_14223,N_14035);
or U14615 (N_14615,N_14341,N_14049);
and U14616 (N_14616,N_14028,N_14315);
and U14617 (N_14617,N_14263,N_14123);
and U14618 (N_14618,N_14443,N_14313);
or U14619 (N_14619,N_14255,N_14163);
or U14620 (N_14620,N_14303,N_14257);
nand U14621 (N_14621,N_14419,N_14294);
or U14622 (N_14622,N_14388,N_14242);
and U14623 (N_14623,N_14067,N_14199);
nor U14624 (N_14624,N_14440,N_14141);
and U14625 (N_14625,N_14371,N_14404);
or U14626 (N_14626,N_14414,N_14333);
and U14627 (N_14627,N_14373,N_14272);
nand U14628 (N_14628,N_14393,N_14402);
and U14629 (N_14629,N_14427,N_14238);
and U14630 (N_14630,N_14451,N_14032);
or U14631 (N_14631,N_14261,N_14279);
or U14632 (N_14632,N_14488,N_14469);
or U14633 (N_14633,N_14418,N_14200);
nor U14634 (N_14634,N_14104,N_14090);
nand U14635 (N_14635,N_14129,N_14462);
nand U14636 (N_14636,N_14063,N_14471);
or U14637 (N_14637,N_14101,N_14386);
nand U14638 (N_14638,N_14064,N_14209);
nand U14639 (N_14639,N_14314,N_14413);
nor U14640 (N_14640,N_14062,N_14331);
or U14641 (N_14641,N_14039,N_14441);
or U14642 (N_14642,N_14087,N_14079);
or U14643 (N_14643,N_14456,N_14057);
nand U14644 (N_14644,N_14172,N_14044);
nor U14645 (N_14645,N_14190,N_14434);
and U14646 (N_14646,N_14389,N_14436);
or U14647 (N_14647,N_14482,N_14380);
and U14648 (N_14648,N_14164,N_14076);
nand U14649 (N_14649,N_14075,N_14145);
and U14650 (N_14650,N_14286,N_14483);
nand U14651 (N_14651,N_14338,N_14241);
nand U14652 (N_14652,N_14360,N_14191);
nand U14653 (N_14653,N_14454,N_14143);
nand U14654 (N_14654,N_14496,N_14301);
nand U14655 (N_14655,N_14258,N_14487);
xor U14656 (N_14656,N_14176,N_14323);
nor U14657 (N_14657,N_14300,N_14188);
nand U14658 (N_14658,N_14159,N_14464);
nand U14659 (N_14659,N_14021,N_14351);
or U14660 (N_14660,N_14290,N_14282);
and U14661 (N_14661,N_14316,N_14307);
nand U14662 (N_14662,N_14103,N_14265);
nand U14663 (N_14663,N_14484,N_14269);
nor U14664 (N_14664,N_14194,N_14114);
nor U14665 (N_14665,N_14459,N_14214);
or U14666 (N_14666,N_14212,N_14072);
nor U14667 (N_14667,N_14387,N_14167);
nand U14668 (N_14668,N_14162,N_14003);
and U14669 (N_14669,N_14177,N_14030);
or U14670 (N_14670,N_14276,N_14390);
and U14671 (N_14671,N_14398,N_14381);
nand U14672 (N_14672,N_14122,N_14268);
or U14673 (N_14673,N_14091,N_14295);
nor U14674 (N_14674,N_14113,N_14058);
or U14675 (N_14675,N_14138,N_14450);
or U14676 (N_14676,N_14026,N_14025);
nor U14677 (N_14677,N_14383,N_14175);
nand U14678 (N_14678,N_14317,N_14071);
or U14679 (N_14679,N_14343,N_14494);
and U14680 (N_14680,N_14391,N_14353);
or U14681 (N_14681,N_14054,N_14379);
or U14682 (N_14682,N_14365,N_14403);
and U14683 (N_14683,N_14131,N_14171);
and U14684 (N_14684,N_14374,N_14479);
nor U14685 (N_14685,N_14115,N_14259);
and U14686 (N_14686,N_14359,N_14168);
nor U14687 (N_14687,N_14372,N_14332);
nand U14688 (N_14688,N_14392,N_14180);
nor U14689 (N_14689,N_14106,N_14328);
nand U14690 (N_14690,N_14339,N_14004);
or U14691 (N_14691,N_14461,N_14304);
nand U14692 (N_14692,N_14111,N_14222);
or U14693 (N_14693,N_14236,N_14445);
nand U14694 (N_14694,N_14457,N_14155);
or U14695 (N_14695,N_14154,N_14463);
and U14696 (N_14696,N_14285,N_14291);
nand U14697 (N_14697,N_14052,N_14243);
or U14698 (N_14698,N_14349,N_14024);
nor U14699 (N_14699,N_14187,N_14069);
nor U14700 (N_14700,N_14499,N_14029);
or U14701 (N_14701,N_14020,N_14439);
or U14702 (N_14702,N_14354,N_14477);
nor U14703 (N_14703,N_14324,N_14165);
nor U14704 (N_14704,N_14396,N_14495);
and U14705 (N_14705,N_14001,N_14267);
and U14706 (N_14706,N_14139,N_14121);
and U14707 (N_14707,N_14107,N_14498);
nand U14708 (N_14708,N_14170,N_14119);
nand U14709 (N_14709,N_14065,N_14181);
or U14710 (N_14710,N_14330,N_14228);
nor U14711 (N_14711,N_14130,N_14250);
nand U14712 (N_14712,N_14002,N_14099);
nand U14713 (N_14713,N_14096,N_14481);
or U14714 (N_14714,N_14306,N_14160);
and U14715 (N_14715,N_14006,N_14310);
nand U14716 (N_14716,N_14136,N_14203);
and U14717 (N_14717,N_14478,N_14292);
nand U14718 (N_14718,N_14078,N_14426);
nor U14719 (N_14719,N_14320,N_14247);
nor U14720 (N_14720,N_14342,N_14492);
nor U14721 (N_14721,N_14422,N_14204);
nor U14722 (N_14722,N_14256,N_14161);
nand U14723 (N_14723,N_14189,N_14217);
nor U14724 (N_14724,N_14476,N_14449);
nor U14725 (N_14725,N_14325,N_14215);
and U14726 (N_14726,N_14368,N_14287);
or U14727 (N_14727,N_14384,N_14084);
nand U14728 (N_14728,N_14448,N_14166);
nand U14729 (N_14729,N_14023,N_14088);
xnor U14730 (N_14730,N_14042,N_14385);
nor U14731 (N_14731,N_14283,N_14146);
nor U14732 (N_14732,N_14185,N_14245);
or U14733 (N_14733,N_14370,N_14033);
nor U14734 (N_14734,N_14015,N_14254);
nor U14735 (N_14735,N_14336,N_14406);
xnor U14736 (N_14736,N_14453,N_14318);
nor U14737 (N_14737,N_14235,N_14337);
nor U14738 (N_14738,N_14118,N_14281);
or U14739 (N_14739,N_14375,N_14201);
nor U14740 (N_14740,N_14066,N_14280);
nor U14741 (N_14741,N_14059,N_14092);
and U14742 (N_14742,N_14356,N_14378);
nor U14743 (N_14743,N_14458,N_14158);
nor U14744 (N_14744,N_14394,N_14048);
or U14745 (N_14745,N_14017,N_14036);
nand U14746 (N_14746,N_14363,N_14220);
nor U14747 (N_14747,N_14085,N_14193);
nand U14748 (N_14748,N_14244,N_14116);
or U14749 (N_14749,N_14000,N_14053);
or U14750 (N_14750,N_14146,N_14462);
nand U14751 (N_14751,N_14423,N_14301);
and U14752 (N_14752,N_14217,N_14014);
nor U14753 (N_14753,N_14347,N_14096);
or U14754 (N_14754,N_14152,N_14345);
or U14755 (N_14755,N_14064,N_14076);
nor U14756 (N_14756,N_14124,N_14012);
and U14757 (N_14757,N_14003,N_14074);
or U14758 (N_14758,N_14228,N_14363);
and U14759 (N_14759,N_14206,N_14231);
and U14760 (N_14760,N_14493,N_14437);
and U14761 (N_14761,N_14236,N_14315);
nand U14762 (N_14762,N_14251,N_14241);
nand U14763 (N_14763,N_14417,N_14011);
or U14764 (N_14764,N_14148,N_14072);
nand U14765 (N_14765,N_14074,N_14244);
nor U14766 (N_14766,N_14455,N_14135);
or U14767 (N_14767,N_14380,N_14325);
nor U14768 (N_14768,N_14203,N_14382);
nand U14769 (N_14769,N_14212,N_14176);
nor U14770 (N_14770,N_14029,N_14470);
nand U14771 (N_14771,N_14013,N_14484);
or U14772 (N_14772,N_14495,N_14431);
nand U14773 (N_14773,N_14222,N_14446);
nand U14774 (N_14774,N_14041,N_14155);
and U14775 (N_14775,N_14317,N_14190);
or U14776 (N_14776,N_14383,N_14354);
nand U14777 (N_14777,N_14388,N_14173);
nor U14778 (N_14778,N_14409,N_14291);
and U14779 (N_14779,N_14053,N_14490);
and U14780 (N_14780,N_14089,N_14411);
nand U14781 (N_14781,N_14176,N_14403);
nand U14782 (N_14782,N_14330,N_14369);
or U14783 (N_14783,N_14470,N_14382);
nand U14784 (N_14784,N_14252,N_14291);
nand U14785 (N_14785,N_14207,N_14202);
nand U14786 (N_14786,N_14186,N_14307);
nand U14787 (N_14787,N_14346,N_14168);
nor U14788 (N_14788,N_14247,N_14179);
and U14789 (N_14789,N_14306,N_14056);
or U14790 (N_14790,N_14155,N_14298);
and U14791 (N_14791,N_14213,N_14475);
nor U14792 (N_14792,N_14463,N_14079);
and U14793 (N_14793,N_14272,N_14264);
nand U14794 (N_14794,N_14009,N_14421);
and U14795 (N_14795,N_14030,N_14302);
nor U14796 (N_14796,N_14383,N_14255);
or U14797 (N_14797,N_14422,N_14011);
or U14798 (N_14798,N_14411,N_14199);
and U14799 (N_14799,N_14311,N_14073);
and U14800 (N_14800,N_14450,N_14053);
nor U14801 (N_14801,N_14102,N_14177);
nor U14802 (N_14802,N_14420,N_14334);
nor U14803 (N_14803,N_14204,N_14207);
or U14804 (N_14804,N_14494,N_14383);
nor U14805 (N_14805,N_14171,N_14058);
nand U14806 (N_14806,N_14197,N_14272);
xnor U14807 (N_14807,N_14157,N_14264);
nand U14808 (N_14808,N_14366,N_14266);
and U14809 (N_14809,N_14398,N_14232);
nand U14810 (N_14810,N_14240,N_14494);
or U14811 (N_14811,N_14493,N_14463);
nor U14812 (N_14812,N_14320,N_14350);
and U14813 (N_14813,N_14022,N_14349);
or U14814 (N_14814,N_14101,N_14341);
nand U14815 (N_14815,N_14227,N_14436);
nand U14816 (N_14816,N_14076,N_14383);
or U14817 (N_14817,N_14381,N_14168);
nand U14818 (N_14818,N_14090,N_14095);
and U14819 (N_14819,N_14314,N_14375);
and U14820 (N_14820,N_14219,N_14114);
or U14821 (N_14821,N_14265,N_14360);
or U14822 (N_14822,N_14253,N_14314);
nand U14823 (N_14823,N_14038,N_14299);
and U14824 (N_14824,N_14225,N_14055);
or U14825 (N_14825,N_14443,N_14091);
or U14826 (N_14826,N_14134,N_14339);
and U14827 (N_14827,N_14318,N_14139);
nor U14828 (N_14828,N_14190,N_14100);
and U14829 (N_14829,N_14458,N_14130);
or U14830 (N_14830,N_14493,N_14429);
and U14831 (N_14831,N_14193,N_14430);
nand U14832 (N_14832,N_14465,N_14323);
and U14833 (N_14833,N_14193,N_14278);
xor U14834 (N_14834,N_14281,N_14410);
nor U14835 (N_14835,N_14098,N_14340);
nor U14836 (N_14836,N_14253,N_14029);
and U14837 (N_14837,N_14416,N_14136);
nand U14838 (N_14838,N_14008,N_14374);
or U14839 (N_14839,N_14061,N_14173);
and U14840 (N_14840,N_14353,N_14160);
or U14841 (N_14841,N_14071,N_14176);
nor U14842 (N_14842,N_14443,N_14437);
nand U14843 (N_14843,N_14038,N_14177);
or U14844 (N_14844,N_14342,N_14245);
or U14845 (N_14845,N_14334,N_14018);
and U14846 (N_14846,N_14403,N_14070);
and U14847 (N_14847,N_14046,N_14000);
nand U14848 (N_14848,N_14356,N_14271);
nand U14849 (N_14849,N_14136,N_14151);
nor U14850 (N_14850,N_14158,N_14371);
nor U14851 (N_14851,N_14173,N_14295);
and U14852 (N_14852,N_14062,N_14424);
nor U14853 (N_14853,N_14130,N_14486);
and U14854 (N_14854,N_14281,N_14411);
nor U14855 (N_14855,N_14189,N_14437);
or U14856 (N_14856,N_14315,N_14004);
nand U14857 (N_14857,N_14238,N_14477);
and U14858 (N_14858,N_14104,N_14318);
or U14859 (N_14859,N_14220,N_14036);
and U14860 (N_14860,N_14293,N_14490);
nand U14861 (N_14861,N_14148,N_14051);
nor U14862 (N_14862,N_14338,N_14275);
or U14863 (N_14863,N_14284,N_14383);
nand U14864 (N_14864,N_14442,N_14394);
or U14865 (N_14865,N_14345,N_14350);
and U14866 (N_14866,N_14460,N_14103);
nor U14867 (N_14867,N_14339,N_14466);
nor U14868 (N_14868,N_14128,N_14443);
nand U14869 (N_14869,N_14348,N_14283);
nand U14870 (N_14870,N_14442,N_14226);
nand U14871 (N_14871,N_14145,N_14187);
or U14872 (N_14872,N_14186,N_14297);
nor U14873 (N_14873,N_14018,N_14483);
and U14874 (N_14874,N_14064,N_14264);
nand U14875 (N_14875,N_14229,N_14347);
nand U14876 (N_14876,N_14329,N_14097);
nand U14877 (N_14877,N_14031,N_14316);
or U14878 (N_14878,N_14009,N_14325);
or U14879 (N_14879,N_14435,N_14242);
nor U14880 (N_14880,N_14297,N_14214);
and U14881 (N_14881,N_14460,N_14253);
nor U14882 (N_14882,N_14071,N_14192);
and U14883 (N_14883,N_14205,N_14430);
nor U14884 (N_14884,N_14199,N_14227);
or U14885 (N_14885,N_14236,N_14009);
nand U14886 (N_14886,N_14046,N_14330);
and U14887 (N_14887,N_14435,N_14393);
and U14888 (N_14888,N_14015,N_14221);
or U14889 (N_14889,N_14010,N_14219);
or U14890 (N_14890,N_14303,N_14363);
and U14891 (N_14891,N_14313,N_14018);
and U14892 (N_14892,N_14415,N_14015);
nor U14893 (N_14893,N_14444,N_14061);
or U14894 (N_14894,N_14191,N_14407);
nand U14895 (N_14895,N_14478,N_14061);
nor U14896 (N_14896,N_14458,N_14374);
and U14897 (N_14897,N_14495,N_14033);
nor U14898 (N_14898,N_14477,N_14250);
nand U14899 (N_14899,N_14189,N_14161);
nor U14900 (N_14900,N_14456,N_14437);
nand U14901 (N_14901,N_14439,N_14166);
nor U14902 (N_14902,N_14439,N_14148);
or U14903 (N_14903,N_14205,N_14192);
or U14904 (N_14904,N_14074,N_14261);
nand U14905 (N_14905,N_14451,N_14400);
or U14906 (N_14906,N_14472,N_14127);
and U14907 (N_14907,N_14262,N_14153);
nand U14908 (N_14908,N_14465,N_14476);
and U14909 (N_14909,N_14229,N_14000);
nor U14910 (N_14910,N_14171,N_14181);
xnor U14911 (N_14911,N_14237,N_14303);
nand U14912 (N_14912,N_14444,N_14298);
or U14913 (N_14913,N_14087,N_14478);
nand U14914 (N_14914,N_14033,N_14011);
nand U14915 (N_14915,N_14151,N_14377);
and U14916 (N_14916,N_14359,N_14453);
or U14917 (N_14917,N_14016,N_14015);
nand U14918 (N_14918,N_14045,N_14138);
or U14919 (N_14919,N_14375,N_14009);
or U14920 (N_14920,N_14380,N_14042);
nand U14921 (N_14921,N_14423,N_14045);
nand U14922 (N_14922,N_14486,N_14463);
or U14923 (N_14923,N_14364,N_14454);
or U14924 (N_14924,N_14423,N_14107);
and U14925 (N_14925,N_14069,N_14249);
and U14926 (N_14926,N_14402,N_14454);
or U14927 (N_14927,N_14120,N_14411);
and U14928 (N_14928,N_14261,N_14400);
nor U14929 (N_14929,N_14490,N_14055);
and U14930 (N_14930,N_14413,N_14200);
or U14931 (N_14931,N_14473,N_14467);
and U14932 (N_14932,N_14409,N_14160);
nand U14933 (N_14933,N_14170,N_14281);
and U14934 (N_14934,N_14241,N_14419);
and U14935 (N_14935,N_14028,N_14109);
and U14936 (N_14936,N_14442,N_14388);
xnor U14937 (N_14937,N_14455,N_14127);
and U14938 (N_14938,N_14067,N_14387);
nor U14939 (N_14939,N_14402,N_14254);
nor U14940 (N_14940,N_14455,N_14016);
nand U14941 (N_14941,N_14456,N_14259);
nand U14942 (N_14942,N_14042,N_14181);
and U14943 (N_14943,N_14181,N_14104);
and U14944 (N_14944,N_14052,N_14054);
or U14945 (N_14945,N_14103,N_14143);
nor U14946 (N_14946,N_14275,N_14295);
nor U14947 (N_14947,N_14317,N_14349);
or U14948 (N_14948,N_14011,N_14435);
and U14949 (N_14949,N_14176,N_14086);
nor U14950 (N_14950,N_14302,N_14443);
nand U14951 (N_14951,N_14127,N_14390);
nand U14952 (N_14952,N_14155,N_14367);
or U14953 (N_14953,N_14326,N_14145);
and U14954 (N_14954,N_14416,N_14365);
nand U14955 (N_14955,N_14344,N_14287);
or U14956 (N_14956,N_14478,N_14057);
and U14957 (N_14957,N_14208,N_14305);
nand U14958 (N_14958,N_14171,N_14265);
nand U14959 (N_14959,N_14428,N_14112);
nor U14960 (N_14960,N_14178,N_14470);
and U14961 (N_14961,N_14224,N_14297);
or U14962 (N_14962,N_14357,N_14475);
or U14963 (N_14963,N_14465,N_14364);
nand U14964 (N_14964,N_14103,N_14095);
or U14965 (N_14965,N_14264,N_14081);
or U14966 (N_14966,N_14480,N_14126);
nor U14967 (N_14967,N_14165,N_14189);
nor U14968 (N_14968,N_14321,N_14169);
nand U14969 (N_14969,N_14487,N_14138);
nand U14970 (N_14970,N_14350,N_14011);
nor U14971 (N_14971,N_14297,N_14191);
or U14972 (N_14972,N_14121,N_14269);
nor U14973 (N_14973,N_14106,N_14156);
or U14974 (N_14974,N_14030,N_14268);
and U14975 (N_14975,N_14086,N_14082);
nor U14976 (N_14976,N_14032,N_14426);
nor U14977 (N_14977,N_14233,N_14094);
nand U14978 (N_14978,N_14147,N_14436);
and U14979 (N_14979,N_14063,N_14428);
and U14980 (N_14980,N_14312,N_14462);
and U14981 (N_14981,N_14318,N_14165);
nand U14982 (N_14982,N_14214,N_14224);
and U14983 (N_14983,N_14060,N_14133);
and U14984 (N_14984,N_14430,N_14226);
nand U14985 (N_14985,N_14063,N_14077);
or U14986 (N_14986,N_14340,N_14251);
and U14987 (N_14987,N_14332,N_14180);
nand U14988 (N_14988,N_14407,N_14402);
nor U14989 (N_14989,N_14277,N_14016);
or U14990 (N_14990,N_14229,N_14150);
nand U14991 (N_14991,N_14376,N_14211);
or U14992 (N_14992,N_14411,N_14488);
nand U14993 (N_14993,N_14242,N_14266);
nand U14994 (N_14994,N_14140,N_14253);
and U14995 (N_14995,N_14074,N_14341);
nand U14996 (N_14996,N_14459,N_14424);
and U14997 (N_14997,N_14289,N_14096);
nor U14998 (N_14998,N_14038,N_14135);
nand U14999 (N_14999,N_14292,N_14296);
nand U15000 (N_15000,N_14942,N_14917);
xnor U15001 (N_15001,N_14657,N_14559);
and U15002 (N_15002,N_14759,N_14505);
nor U15003 (N_15003,N_14563,N_14592);
or U15004 (N_15004,N_14808,N_14969);
or U15005 (N_15005,N_14647,N_14513);
nand U15006 (N_15006,N_14807,N_14701);
and U15007 (N_15007,N_14736,N_14791);
nand U15008 (N_15008,N_14790,N_14678);
nor U15009 (N_15009,N_14768,N_14504);
nand U15010 (N_15010,N_14507,N_14685);
nor U15011 (N_15011,N_14605,N_14508);
or U15012 (N_15012,N_14755,N_14985);
and U15013 (N_15013,N_14749,N_14772);
nand U15014 (N_15014,N_14882,N_14547);
nand U15015 (N_15015,N_14855,N_14517);
xor U15016 (N_15016,N_14959,N_14528);
or U15017 (N_15017,N_14918,N_14745);
nand U15018 (N_15018,N_14949,N_14624);
and U15019 (N_15019,N_14860,N_14621);
nor U15020 (N_15020,N_14981,N_14620);
and U15021 (N_15021,N_14703,N_14560);
and U15022 (N_15022,N_14904,N_14512);
nor U15023 (N_15023,N_14966,N_14570);
and U15024 (N_15024,N_14540,N_14670);
and U15025 (N_15025,N_14608,N_14542);
nor U15026 (N_15026,N_14932,N_14683);
or U15027 (N_15027,N_14919,N_14561);
nand U15028 (N_15028,N_14973,N_14899);
and U15029 (N_15029,N_14688,N_14668);
and U15030 (N_15030,N_14631,N_14632);
or U15031 (N_15031,N_14622,N_14723);
nand U15032 (N_15032,N_14835,N_14720);
or U15033 (N_15033,N_14609,N_14963);
and U15034 (N_15034,N_14789,N_14849);
or U15035 (N_15035,N_14618,N_14617);
and U15036 (N_15036,N_14898,N_14660);
nand U15037 (N_15037,N_14572,N_14937);
or U15038 (N_15038,N_14598,N_14602);
nor U15039 (N_15039,N_14953,N_14874);
nor U15040 (N_15040,N_14801,N_14551);
or U15041 (N_15041,N_14708,N_14532);
or U15042 (N_15042,N_14521,N_14838);
nor U15043 (N_15043,N_14591,N_14848);
nor U15044 (N_15044,N_14730,N_14948);
or U15045 (N_15045,N_14506,N_14748);
nor U15046 (N_15046,N_14763,N_14765);
nor U15047 (N_15047,N_14941,N_14788);
or U15048 (N_15048,N_14646,N_14533);
nand U15049 (N_15049,N_14641,N_14696);
nor U15050 (N_15050,N_14672,N_14691);
nor U15051 (N_15051,N_14950,N_14722);
nand U15052 (N_15052,N_14803,N_14821);
and U15053 (N_15053,N_14663,N_14931);
nor U15054 (N_15054,N_14721,N_14929);
nor U15055 (N_15055,N_14690,N_14869);
nor U15056 (N_15056,N_14589,N_14792);
nand U15057 (N_15057,N_14652,N_14576);
or U15058 (N_15058,N_14524,N_14968);
nor U15059 (N_15059,N_14771,N_14800);
and U15060 (N_15060,N_14778,N_14897);
and U15061 (N_15061,N_14541,N_14654);
and U15062 (N_15062,N_14908,N_14662);
nand U15063 (N_15063,N_14735,N_14747);
and U15064 (N_15064,N_14834,N_14579);
nand U15065 (N_15065,N_14550,N_14704);
and U15066 (N_15066,N_14638,N_14593);
nor U15067 (N_15067,N_14554,N_14694);
nor U15068 (N_15068,N_14862,N_14852);
nor U15069 (N_15069,N_14676,N_14828);
and U15070 (N_15070,N_14961,N_14752);
nand U15071 (N_15071,N_14984,N_14920);
or U15072 (N_15072,N_14590,N_14956);
and U15073 (N_15073,N_14876,N_14910);
or U15074 (N_15074,N_14830,N_14965);
nor U15075 (N_15075,N_14500,N_14717);
nand U15076 (N_15076,N_14846,N_14831);
nand U15077 (N_15077,N_14843,N_14601);
nor U15078 (N_15078,N_14725,N_14999);
or U15079 (N_15079,N_14659,N_14728);
or U15080 (N_15080,N_14727,N_14635);
nand U15081 (N_15081,N_14986,N_14992);
or U15082 (N_15082,N_14861,N_14509);
nand U15083 (N_15083,N_14557,N_14648);
nor U15084 (N_15084,N_14753,N_14653);
or U15085 (N_15085,N_14630,N_14603);
or U15086 (N_15086,N_14502,N_14955);
or U15087 (N_15087,N_14640,N_14594);
nor U15088 (N_15088,N_14583,N_14614);
nor U15089 (N_15089,N_14825,N_14582);
and U15090 (N_15090,N_14935,N_14675);
and U15091 (N_15091,N_14894,N_14545);
or U15092 (N_15092,N_14684,N_14799);
nand U15093 (N_15093,N_14851,N_14581);
or U15094 (N_15094,N_14510,N_14567);
nor U15095 (N_15095,N_14809,N_14650);
nor U15096 (N_15096,N_14889,N_14895);
nand U15097 (N_15097,N_14795,N_14850);
and U15098 (N_15098,N_14548,N_14818);
nor U15099 (N_15099,N_14974,N_14964);
nor U15100 (N_15100,N_14661,N_14740);
and U15101 (N_15101,N_14700,N_14979);
nor U15102 (N_15102,N_14742,N_14756);
or U15103 (N_15103,N_14766,N_14936);
or U15104 (N_15104,N_14833,N_14892);
xnor U15105 (N_15105,N_14751,N_14757);
and U15106 (N_15106,N_14868,N_14805);
and U15107 (N_15107,N_14698,N_14724);
or U15108 (N_15108,N_14867,N_14633);
and U15109 (N_15109,N_14875,N_14534);
nand U15110 (N_15110,N_14655,N_14713);
or U15111 (N_15111,N_14926,N_14909);
xor U15112 (N_15112,N_14954,N_14893);
or U15113 (N_15113,N_14546,N_14812);
or U15114 (N_15114,N_14970,N_14604);
and U15115 (N_15115,N_14770,N_14938);
and U15116 (N_15116,N_14613,N_14634);
nand U15117 (N_15117,N_14880,N_14944);
nor U15118 (N_15118,N_14832,N_14535);
and U15119 (N_15119,N_14775,N_14706);
and U15120 (N_15120,N_14967,N_14923);
and U15121 (N_15121,N_14989,N_14962);
nand U15122 (N_15122,N_14529,N_14527);
or U15123 (N_15123,N_14573,N_14764);
and U15124 (N_15124,N_14612,N_14743);
and U15125 (N_15125,N_14837,N_14939);
or U15126 (N_15126,N_14811,N_14896);
and U15127 (N_15127,N_14731,N_14983);
nor U15128 (N_15128,N_14695,N_14519);
nor U15129 (N_15129,N_14710,N_14958);
or U15130 (N_15130,N_14726,N_14794);
and U15131 (N_15131,N_14997,N_14879);
and U15132 (N_15132,N_14991,N_14623);
nor U15133 (N_15133,N_14530,N_14993);
nand U15134 (N_15134,N_14697,N_14577);
and U15135 (N_15135,N_14565,N_14681);
or U15136 (N_15136,N_14819,N_14943);
nor U15137 (N_15137,N_14522,N_14569);
xnor U15138 (N_15138,N_14972,N_14520);
or U15139 (N_15139,N_14785,N_14739);
or U15140 (N_15140,N_14568,N_14586);
nand U15141 (N_15141,N_14587,N_14976);
xor U15142 (N_15142,N_14501,N_14922);
and U15143 (N_15143,N_14995,N_14544);
and U15144 (N_15144,N_14715,N_14610);
nor U15145 (N_15145,N_14796,N_14656);
or U15146 (N_15146,N_14616,N_14885);
and U15147 (N_15147,N_14864,N_14978);
and U15148 (N_15148,N_14824,N_14716);
or U15149 (N_15149,N_14606,N_14921);
and U15150 (N_15150,N_14626,N_14729);
nand U15151 (N_15151,N_14556,N_14671);
or U15152 (N_15152,N_14754,N_14669);
nand U15153 (N_15153,N_14679,N_14947);
xnor U15154 (N_15154,N_14625,N_14552);
or U15155 (N_15155,N_14890,N_14866);
or U15156 (N_15156,N_14627,N_14906);
or U15157 (N_15157,N_14977,N_14971);
or U15158 (N_15158,N_14913,N_14711);
nor U15159 (N_15159,N_14523,N_14856);
nor U15160 (N_15160,N_14928,N_14699);
nand U15161 (N_15161,N_14607,N_14859);
and U15162 (N_15162,N_14930,N_14637);
or U15163 (N_15163,N_14871,N_14649);
nor U15164 (N_15164,N_14596,N_14718);
or U15165 (N_15165,N_14780,N_14538);
or U15166 (N_15166,N_14836,N_14826);
and U15167 (N_15167,N_14998,N_14934);
or U15168 (N_15168,N_14903,N_14776);
nor U15169 (N_15169,N_14762,N_14797);
or U15170 (N_15170,N_14705,N_14777);
nor U15171 (N_15171,N_14677,N_14597);
and U15172 (N_15172,N_14750,N_14584);
and U15173 (N_15173,N_14628,N_14719);
or U15174 (N_15174,N_14940,N_14709);
nand U15175 (N_15175,N_14925,N_14829);
nor U15176 (N_15176,N_14839,N_14987);
nor U15177 (N_15177,N_14863,N_14806);
and U15178 (N_15178,N_14526,N_14916);
and U15179 (N_15179,N_14845,N_14870);
and U15180 (N_15180,N_14813,N_14562);
nor U15181 (N_15181,N_14732,N_14642);
nand U15182 (N_15182,N_14802,N_14664);
nor U15183 (N_15183,N_14782,N_14674);
and U15184 (N_15184,N_14884,N_14888);
nand U15185 (N_15185,N_14927,N_14975);
nand U15186 (N_15186,N_14536,N_14798);
nor U15187 (N_15187,N_14687,N_14553);
nand U15188 (N_15188,N_14600,N_14636);
and U15189 (N_15189,N_14911,N_14957);
and U15190 (N_15190,N_14692,N_14815);
and U15191 (N_15191,N_14810,N_14666);
and U15192 (N_15192,N_14878,N_14822);
and U15193 (N_15193,N_14644,N_14639);
or U15194 (N_15194,N_14629,N_14575);
nand U15195 (N_15195,N_14881,N_14571);
nor U15196 (N_15196,N_14865,N_14531);
nand U15197 (N_15197,N_14980,N_14816);
or U15198 (N_15198,N_14566,N_14945);
nor U15199 (N_15199,N_14645,N_14537);
nand U15200 (N_15200,N_14996,N_14702);
nor U15201 (N_15201,N_14595,N_14854);
or U15202 (N_15202,N_14673,N_14518);
nor U15203 (N_15203,N_14886,N_14787);
nand U15204 (N_15204,N_14574,N_14817);
or U15205 (N_15205,N_14901,N_14611);
nand U15206 (N_15206,N_14902,N_14990);
or U15207 (N_15207,N_14781,N_14667);
nand U15208 (N_15208,N_14912,N_14853);
and U15209 (N_15209,N_14651,N_14914);
xor U15210 (N_15210,N_14516,N_14712);
nand U15211 (N_15211,N_14555,N_14841);
nor U15212 (N_15212,N_14786,N_14820);
and U15213 (N_15213,N_14599,N_14767);
nand U15214 (N_15214,N_14744,N_14827);
and U15215 (N_15215,N_14814,N_14951);
or U15216 (N_15216,N_14804,N_14769);
nor U15217 (N_15217,N_14946,N_14511);
or U15218 (N_15218,N_14883,N_14741);
nand U15219 (N_15219,N_14761,N_14924);
nor U15220 (N_15220,N_14907,N_14714);
nor U15221 (N_15221,N_14564,N_14686);
xor U15222 (N_15222,N_14994,N_14858);
or U15223 (N_15223,N_14689,N_14515);
or U15224 (N_15224,N_14707,N_14842);
or U15225 (N_15225,N_14737,N_14774);
nand U15226 (N_15226,N_14844,N_14988);
and U15227 (N_15227,N_14952,N_14847);
nor U15228 (N_15228,N_14760,N_14734);
nand U15229 (N_15229,N_14873,N_14680);
nor U15230 (N_15230,N_14887,N_14877);
nor U15231 (N_15231,N_14960,N_14578);
or U15232 (N_15232,N_14915,N_14840);
nand U15233 (N_15233,N_14588,N_14783);
nand U15234 (N_15234,N_14738,N_14543);
or U15235 (N_15235,N_14558,N_14900);
and U15236 (N_15236,N_14615,N_14933);
and U15237 (N_15237,N_14682,N_14580);
or U15238 (N_15238,N_14779,N_14693);
and U15239 (N_15239,N_14773,N_14619);
nor U15240 (N_15240,N_14746,N_14503);
nand U15241 (N_15241,N_14733,N_14857);
nand U15242 (N_15242,N_14585,N_14823);
nor U15243 (N_15243,N_14514,N_14525);
nor U15244 (N_15244,N_14549,N_14891);
nor U15245 (N_15245,N_14665,N_14539);
nand U15246 (N_15246,N_14793,N_14982);
or U15247 (N_15247,N_14658,N_14643);
or U15248 (N_15248,N_14872,N_14784);
and U15249 (N_15249,N_14758,N_14905);
or U15250 (N_15250,N_14521,N_14891);
nand U15251 (N_15251,N_14780,N_14725);
and U15252 (N_15252,N_14965,N_14735);
and U15253 (N_15253,N_14958,N_14618);
or U15254 (N_15254,N_14625,N_14922);
nand U15255 (N_15255,N_14621,N_14582);
nor U15256 (N_15256,N_14768,N_14541);
xor U15257 (N_15257,N_14636,N_14524);
and U15258 (N_15258,N_14978,N_14754);
nand U15259 (N_15259,N_14770,N_14516);
or U15260 (N_15260,N_14691,N_14623);
and U15261 (N_15261,N_14590,N_14819);
nand U15262 (N_15262,N_14598,N_14851);
or U15263 (N_15263,N_14724,N_14652);
nand U15264 (N_15264,N_14751,N_14721);
or U15265 (N_15265,N_14645,N_14891);
nand U15266 (N_15266,N_14806,N_14585);
and U15267 (N_15267,N_14696,N_14646);
or U15268 (N_15268,N_14624,N_14538);
nor U15269 (N_15269,N_14566,N_14744);
nand U15270 (N_15270,N_14827,N_14921);
and U15271 (N_15271,N_14759,N_14955);
and U15272 (N_15272,N_14813,N_14899);
or U15273 (N_15273,N_14977,N_14613);
or U15274 (N_15274,N_14529,N_14761);
nand U15275 (N_15275,N_14739,N_14513);
nand U15276 (N_15276,N_14668,N_14956);
nor U15277 (N_15277,N_14840,N_14560);
and U15278 (N_15278,N_14814,N_14874);
or U15279 (N_15279,N_14516,N_14900);
or U15280 (N_15280,N_14938,N_14750);
or U15281 (N_15281,N_14713,N_14775);
or U15282 (N_15282,N_14811,N_14552);
or U15283 (N_15283,N_14618,N_14998);
nand U15284 (N_15284,N_14982,N_14635);
nand U15285 (N_15285,N_14801,N_14851);
and U15286 (N_15286,N_14596,N_14861);
nor U15287 (N_15287,N_14738,N_14781);
nand U15288 (N_15288,N_14877,N_14981);
nand U15289 (N_15289,N_14937,N_14959);
nand U15290 (N_15290,N_14907,N_14748);
and U15291 (N_15291,N_14886,N_14732);
or U15292 (N_15292,N_14893,N_14771);
nand U15293 (N_15293,N_14539,N_14888);
nor U15294 (N_15294,N_14852,N_14517);
nand U15295 (N_15295,N_14917,N_14681);
nor U15296 (N_15296,N_14665,N_14777);
nand U15297 (N_15297,N_14606,N_14888);
nand U15298 (N_15298,N_14700,N_14973);
nand U15299 (N_15299,N_14638,N_14960);
nor U15300 (N_15300,N_14730,N_14958);
nor U15301 (N_15301,N_14534,N_14892);
or U15302 (N_15302,N_14553,N_14768);
nor U15303 (N_15303,N_14913,N_14510);
nor U15304 (N_15304,N_14535,N_14887);
nand U15305 (N_15305,N_14925,N_14975);
or U15306 (N_15306,N_14620,N_14595);
nor U15307 (N_15307,N_14898,N_14525);
nor U15308 (N_15308,N_14530,N_14958);
and U15309 (N_15309,N_14753,N_14855);
nor U15310 (N_15310,N_14533,N_14607);
nor U15311 (N_15311,N_14934,N_14919);
and U15312 (N_15312,N_14846,N_14732);
or U15313 (N_15313,N_14632,N_14759);
or U15314 (N_15314,N_14831,N_14668);
or U15315 (N_15315,N_14684,N_14732);
nand U15316 (N_15316,N_14535,N_14646);
and U15317 (N_15317,N_14655,N_14763);
and U15318 (N_15318,N_14901,N_14555);
and U15319 (N_15319,N_14935,N_14596);
nor U15320 (N_15320,N_14593,N_14911);
and U15321 (N_15321,N_14749,N_14654);
nand U15322 (N_15322,N_14539,N_14709);
or U15323 (N_15323,N_14810,N_14888);
or U15324 (N_15324,N_14923,N_14890);
nor U15325 (N_15325,N_14543,N_14871);
nand U15326 (N_15326,N_14762,N_14503);
nor U15327 (N_15327,N_14798,N_14955);
nand U15328 (N_15328,N_14666,N_14563);
nand U15329 (N_15329,N_14905,N_14752);
nand U15330 (N_15330,N_14688,N_14555);
nand U15331 (N_15331,N_14653,N_14683);
and U15332 (N_15332,N_14726,N_14820);
nor U15333 (N_15333,N_14649,N_14596);
and U15334 (N_15334,N_14964,N_14646);
and U15335 (N_15335,N_14860,N_14979);
nor U15336 (N_15336,N_14556,N_14587);
or U15337 (N_15337,N_14994,N_14883);
and U15338 (N_15338,N_14601,N_14757);
nor U15339 (N_15339,N_14584,N_14713);
or U15340 (N_15340,N_14784,N_14665);
or U15341 (N_15341,N_14556,N_14856);
and U15342 (N_15342,N_14603,N_14838);
or U15343 (N_15343,N_14707,N_14591);
and U15344 (N_15344,N_14540,N_14999);
nor U15345 (N_15345,N_14722,N_14802);
and U15346 (N_15346,N_14847,N_14762);
and U15347 (N_15347,N_14813,N_14652);
nor U15348 (N_15348,N_14737,N_14662);
nand U15349 (N_15349,N_14603,N_14878);
nor U15350 (N_15350,N_14563,N_14749);
nor U15351 (N_15351,N_14528,N_14922);
and U15352 (N_15352,N_14676,N_14608);
and U15353 (N_15353,N_14899,N_14951);
and U15354 (N_15354,N_14583,N_14960);
nor U15355 (N_15355,N_14953,N_14743);
and U15356 (N_15356,N_14617,N_14937);
and U15357 (N_15357,N_14768,N_14687);
nand U15358 (N_15358,N_14804,N_14628);
nand U15359 (N_15359,N_14503,N_14697);
nand U15360 (N_15360,N_14714,N_14764);
and U15361 (N_15361,N_14862,N_14915);
or U15362 (N_15362,N_14565,N_14917);
and U15363 (N_15363,N_14537,N_14768);
and U15364 (N_15364,N_14910,N_14506);
and U15365 (N_15365,N_14827,N_14807);
nor U15366 (N_15366,N_14737,N_14712);
nand U15367 (N_15367,N_14780,N_14873);
nand U15368 (N_15368,N_14553,N_14691);
and U15369 (N_15369,N_14574,N_14955);
or U15370 (N_15370,N_14720,N_14628);
and U15371 (N_15371,N_14561,N_14734);
and U15372 (N_15372,N_14827,N_14760);
nand U15373 (N_15373,N_14878,N_14521);
nor U15374 (N_15374,N_14704,N_14607);
nand U15375 (N_15375,N_14617,N_14507);
nand U15376 (N_15376,N_14562,N_14884);
xnor U15377 (N_15377,N_14754,N_14508);
nor U15378 (N_15378,N_14806,N_14793);
and U15379 (N_15379,N_14959,N_14818);
nor U15380 (N_15380,N_14842,N_14989);
nor U15381 (N_15381,N_14525,N_14814);
or U15382 (N_15382,N_14615,N_14875);
nor U15383 (N_15383,N_14626,N_14648);
nor U15384 (N_15384,N_14805,N_14741);
nand U15385 (N_15385,N_14986,N_14830);
nand U15386 (N_15386,N_14678,N_14639);
and U15387 (N_15387,N_14736,N_14725);
nor U15388 (N_15388,N_14848,N_14798);
and U15389 (N_15389,N_14882,N_14788);
and U15390 (N_15390,N_14819,N_14981);
and U15391 (N_15391,N_14826,N_14892);
nand U15392 (N_15392,N_14536,N_14757);
nand U15393 (N_15393,N_14672,N_14893);
nand U15394 (N_15394,N_14782,N_14548);
nand U15395 (N_15395,N_14538,N_14587);
nand U15396 (N_15396,N_14574,N_14802);
nand U15397 (N_15397,N_14598,N_14555);
nand U15398 (N_15398,N_14573,N_14905);
or U15399 (N_15399,N_14562,N_14724);
nor U15400 (N_15400,N_14828,N_14571);
or U15401 (N_15401,N_14961,N_14815);
nand U15402 (N_15402,N_14796,N_14727);
or U15403 (N_15403,N_14986,N_14847);
nor U15404 (N_15404,N_14581,N_14538);
or U15405 (N_15405,N_14616,N_14962);
or U15406 (N_15406,N_14893,N_14502);
nand U15407 (N_15407,N_14636,N_14733);
and U15408 (N_15408,N_14751,N_14611);
and U15409 (N_15409,N_14738,N_14801);
and U15410 (N_15410,N_14516,N_14634);
nand U15411 (N_15411,N_14516,N_14668);
nor U15412 (N_15412,N_14559,N_14879);
nand U15413 (N_15413,N_14919,N_14976);
nor U15414 (N_15414,N_14833,N_14700);
or U15415 (N_15415,N_14783,N_14805);
xor U15416 (N_15416,N_14924,N_14694);
nor U15417 (N_15417,N_14811,N_14668);
nand U15418 (N_15418,N_14547,N_14775);
nor U15419 (N_15419,N_14571,N_14600);
nand U15420 (N_15420,N_14552,N_14638);
or U15421 (N_15421,N_14829,N_14646);
nand U15422 (N_15422,N_14759,N_14510);
nor U15423 (N_15423,N_14741,N_14603);
and U15424 (N_15424,N_14752,N_14648);
or U15425 (N_15425,N_14604,N_14686);
or U15426 (N_15426,N_14886,N_14881);
or U15427 (N_15427,N_14990,N_14963);
nor U15428 (N_15428,N_14520,N_14794);
nor U15429 (N_15429,N_14877,N_14745);
and U15430 (N_15430,N_14712,N_14653);
xor U15431 (N_15431,N_14545,N_14672);
and U15432 (N_15432,N_14585,N_14636);
and U15433 (N_15433,N_14660,N_14862);
nor U15434 (N_15434,N_14980,N_14947);
nor U15435 (N_15435,N_14643,N_14988);
or U15436 (N_15436,N_14800,N_14722);
or U15437 (N_15437,N_14562,N_14921);
nor U15438 (N_15438,N_14534,N_14638);
nand U15439 (N_15439,N_14723,N_14504);
nor U15440 (N_15440,N_14777,N_14706);
nor U15441 (N_15441,N_14832,N_14606);
nand U15442 (N_15442,N_14759,N_14881);
nor U15443 (N_15443,N_14869,N_14804);
nor U15444 (N_15444,N_14859,N_14690);
nor U15445 (N_15445,N_14955,N_14549);
or U15446 (N_15446,N_14550,N_14637);
nor U15447 (N_15447,N_14901,N_14595);
nor U15448 (N_15448,N_14755,N_14930);
xnor U15449 (N_15449,N_14835,N_14825);
nor U15450 (N_15450,N_14937,N_14768);
or U15451 (N_15451,N_14536,N_14892);
or U15452 (N_15452,N_14652,N_14840);
nand U15453 (N_15453,N_14613,N_14638);
nand U15454 (N_15454,N_14671,N_14979);
or U15455 (N_15455,N_14793,N_14650);
nor U15456 (N_15456,N_14668,N_14605);
and U15457 (N_15457,N_14721,N_14564);
nor U15458 (N_15458,N_14582,N_14631);
nand U15459 (N_15459,N_14931,N_14526);
nand U15460 (N_15460,N_14578,N_14739);
or U15461 (N_15461,N_14716,N_14515);
nand U15462 (N_15462,N_14928,N_14871);
nand U15463 (N_15463,N_14866,N_14807);
or U15464 (N_15464,N_14696,N_14910);
and U15465 (N_15465,N_14856,N_14791);
or U15466 (N_15466,N_14899,N_14570);
or U15467 (N_15467,N_14521,N_14932);
nor U15468 (N_15468,N_14614,N_14559);
or U15469 (N_15469,N_14806,N_14670);
and U15470 (N_15470,N_14925,N_14769);
or U15471 (N_15471,N_14602,N_14528);
nor U15472 (N_15472,N_14614,N_14784);
nor U15473 (N_15473,N_14537,N_14709);
and U15474 (N_15474,N_14712,N_14658);
and U15475 (N_15475,N_14555,N_14785);
or U15476 (N_15476,N_14675,N_14722);
or U15477 (N_15477,N_14766,N_14845);
nor U15478 (N_15478,N_14565,N_14550);
or U15479 (N_15479,N_14964,N_14623);
nand U15480 (N_15480,N_14572,N_14664);
or U15481 (N_15481,N_14673,N_14970);
nand U15482 (N_15482,N_14956,N_14600);
nand U15483 (N_15483,N_14945,N_14794);
nand U15484 (N_15484,N_14878,N_14513);
nor U15485 (N_15485,N_14824,N_14643);
and U15486 (N_15486,N_14606,N_14896);
xnor U15487 (N_15487,N_14568,N_14970);
nand U15488 (N_15488,N_14799,N_14674);
nor U15489 (N_15489,N_14909,N_14856);
and U15490 (N_15490,N_14929,N_14855);
nor U15491 (N_15491,N_14875,N_14993);
nor U15492 (N_15492,N_14848,N_14560);
or U15493 (N_15493,N_14541,N_14582);
nand U15494 (N_15494,N_14721,N_14508);
nand U15495 (N_15495,N_14998,N_14895);
and U15496 (N_15496,N_14751,N_14676);
and U15497 (N_15497,N_14841,N_14610);
or U15498 (N_15498,N_14637,N_14902);
nand U15499 (N_15499,N_14953,N_14726);
or U15500 (N_15500,N_15024,N_15015);
and U15501 (N_15501,N_15014,N_15251);
or U15502 (N_15502,N_15248,N_15061);
nand U15503 (N_15503,N_15123,N_15441);
or U15504 (N_15504,N_15259,N_15361);
nor U15505 (N_15505,N_15241,N_15352);
and U15506 (N_15506,N_15082,N_15207);
and U15507 (N_15507,N_15171,N_15358);
or U15508 (N_15508,N_15111,N_15119);
xor U15509 (N_15509,N_15197,N_15282);
or U15510 (N_15510,N_15449,N_15365);
and U15511 (N_15511,N_15401,N_15329);
nor U15512 (N_15512,N_15287,N_15332);
nand U15513 (N_15513,N_15188,N_15093);
nand U15514 (N_15514,N_15369,N_15027);
and U15515 (N_15515,N_15388,N_15047);
or U15516 (N_15516,N_15295,N_15190);
nand U15517 (N_15517,N_15017,N_15258);
and U15518 (N_15518,N_15398,N_15499);
nor U15519 (N_15519,N_15083,N_15243);
or U15520 (N_15520,N_15336,N_15231);
nand U15521 (N_15521,N_15405,N_15096);
and U15522 (N_15522,N_15163,N_15305);
and U15523 (N_15523,N_15403,N_15060);
and U15524 (N_15524,N_15363,N_15367);
nor U15525 (N_15525,N_15113,N_15025);
nand U15526 (N_15526,N_15051,N_15364);
nor U15527 (N_15527,N_15340,N_15433);
or U15528 (N_15528,N_15186,N_15384);
and U15529 (N_15529,N_15232,N_15319);
and U15530 (N_15530,N_15423,N_15218);
or U15531 (N_15531,N_15318,N_15302);
nand U15532 (N_15532,N_15478,N_15337);
nor U15533 (N_15533,N_15154,N_15010);
and U15534 (N_15534,N_15135,N_15090);
or U15535 (N_15535,N_15124,N_15267);
nand U15536 (N_15536,N_15049,N_15125);
and U15537 (N_15537,N_15469,N_15357);
nor U15538 (N_15538,N_15008,N_15289);
or U15539 (N_15539,N_15048,N_15476);
and U15540 (N_15540,N_15293,N_15290);
nand U15541 (N_15541,N_15372,N_15417);
nor U15542 (N_15542,N_15345,N_15198);
or U15543 (N_15543,N_15274,N_15373);
nor U15544 (N_15544,N_15456,N_15344);
nor U15545 (N_15545,N_15247,N_15300);
nand U15546 (N_15546,N_15346,N_15185);
and U15547 (N_15547,N_15483,N_15443);
or U15548 (N_15548,N_15129,N_15054);
or U15549 (N_15549,N_15296,N_15331);
nand U15550 (N_15550,N_15165,N_15042);
and U15551 (N_15551,N_15005,N_15438);
and U15552 (N_15552,N_15058,N_15084);
nand U15553 (N_15553,N_15159,N_15236);
nand U15554 (N_15554,N_15238,N_15276);
nor U15555 (N_15555,N_15203,N_15204);
or U15556 (N_15556,N_15145,N_15172);
nand U15557 (N_15557,N_15088,N_15155);
or U15558 (N_15558,N_15069,N_15177);
and U15559 (N_15559,N_15130,N_15050);
xor U15560 (N_15560,N_15037,N_15448);
nor U15561 (N_15561,N_15407,N_15487);
and U15562 (N_15562,N_15235,N_15339);
and U15563 (N_15563,N_15180,N_15304);
nand U15564 (N_15564,N_15484,N_15467);
and U15565 (N_15565,N_15034,N_15189);
or U15566 (N_15566,N_15019,N_15271);
nand U15567 (N_15567,N_15098,N_15206);
and U15568 (N_15568,N_15440,N_15000);
nor U15569 (N_15569,N_15110,N_15288);
and U15570 (N_15570,N_15278,N_15408);
or U15571 (N_15571,N_15310,N_15269);
nor U15572 (N_15572,N_15077,N_15261);
or U15573 (N_15573,N_15263,N_15316);
and U15574 (N_15574,N_15488,N_15161);
or U15575 (N_15575,N_15201,N_15078);
nor U15576 (N_15576,N_15033,N_15459);
nand U15577 (N_15577,N_15396,N_15052);
and U15578 (N_15578,N_15064,N_15209);
xor U15579 (N_15579,N_15018,N_15230);
nor U15580 (N_15580,N_15292,N_15118);
nand U15581 (N_15581,N_15097,N_15450);
nand U15582 (N_15582,N_15260,N_15425);
or U15583 (N_15583,N_15285,N_15141);
nor U15584 (N_15584,N_15391,N_15157);
and U15585 (N_15585,N_15240,N_15112);
nor U15586 (N_15586,N_15315,N_15181);
nor U15587 (N_15587,N_15477,N_15076);
nand U15588 (N_15588,N_15224,N_15210);
or U15589 (N_15589,N_15242,N_15256);
and U15590 (N_15590,N_15115,N_15133);
nor U15591 (N_15591,N_15351,N_15320);
or U15592 (N_15592,N_15166,N_15187);
nand U15593 (N_15593,N_15321,N_15496);
or U15594 (N_15594,N_15108,N_15265);
nor U15595 (N_15595,N_15043,N_15360);
or U15596 (N_15596,N_15359,N_15453);
nand U15597 (N_15597,N_15193,N_15011);
and U15598 (N_15598,N_15120,N_15040);
and U15599 (N_15599,N_15341,N_15137);
nand U15600 (N_15600,N_15176,N_15264);
nor U15601 (N_15601,N_15021,N_15091);
nor U15602 (N_15602,N_15106,N_15291);
nor U15603 (N_15603,N_15307,N_15192);
and U15604 (N_15604,N_15452,N_15479);
nor U15605 (N_15605,N_15462,N_15109);
nor U15606 (N_15606,N_15143,N_15080);
nor U15607 (N_15607,N_15086,N_15480);
nand U15608 (N_15608,N_15325,N_15099);
and U15609 (N_15609,N_15226,N_15200);
nand U15610 (N_15610,N_15056,N_15087);
nand U15611 (N_15611,N_15308,N_15322);
and U15612 (N_15612,N_15128,N_15392);
nand U15613 (N_15613,N_15436,N_15495);
nand U15614 (N_15614,N_15168,N_15013);
and U15615 (N_15615,N_15347,N_15220);
or U15616 (N_15616,N_15342,N_15374);
or U15617 (N_15617,N_15164,N_15006);
nor U15618 (N_15618,N_15073,N_15009);
or U15619 (N_15619,N_15184,N_15039);
nor U15620 (N_15620,N_15221,N_15280);
nor U15621 (N_15621,N_15022,N_15323);
nor U15622 (N_15622,N_15400,N_15030);
nand U15623 (N_15623,N_15286,N_15222);
nor U15624 (N_15624,N_15023,N_15327);
nand U15625 (N_15625,N_15399,N_15065);
or U15626 (N_15626,N_15306,N_15212);
and U15627 (N_15627,N_15252,N_15205);
nor U15628 (N_15628,N_15378,N_15016);
or U15629 (N_15629,N_15046,N_15284);
and U15630 (N_15630,N_15178,N_15279);
nor U15631 (N_15631,N_15415,N_15196);
nand U15632 (N_15632,N_15167,N_15004);
nor U15633 (N_15633,N_15057,N_15475);
nor U15634 (N_15634,N_15208,N_15041);
nand U15635 (N_15635,N_15416,N_15139);
nor U15636 (N_15636,N_15031,N_15386);
and U15637 (N_15637,N_15102,N_15368);
and U15638 (N_15638,N_15268,N_15348);
nand U15639 (N_15639,N_15397,N_15101);
and U15640 (N_15640,N_15429,N_15362);
or U15641 (N_15641,N_15490,N_15445);
nand U15642 (N_15642,N_15434,N_15149);
and U15643 (N_15643,N_15432,N_15406);
nor U15644 (N_15644,N_15461,N_15217);
and U15645 (N_15645,N_15007,N_15072);
or U15646 (N_15646,N_15328,N_15313);
or U15647 (N_15647,N_15116,N_15094);
and U15648 (N_15648,N_15428,N_15444);
nand U15649 (N_15649,N_15381,N_15103);
and U15650 (N_15650,N_15045,N_15117);
nor U15651 (N_15651,N_15144,N_15349);
or U15652 (N_15652,N_15330,N_15053);
nor U15653 (N_15653,N_15063,N_15385);
nor U15654 (N_15654,N_15160,N_15283);
nor U15655 (N_15655,N_15482,N_15326);
nand U15656 (N_15656,N_15001,N_15114);
or U15657 (N_15657,N_15162,N_15311);
nand U15658 (N_15658,N_15153,N_15173);
or U15659 (N_15659,N_15266,N_15382);
and U15660 (N_15660,N_15472,N_15140);
or U15661 (N_15661,N_15107,N_15297);
and U15662 (N_15662,N_15228,N_15194);
and U15663 (N_15663,N_15383,N_15100);
nand U15664 (N_15664,N_15404,N_15148);
nor U15665 (N_15665,N_15431,N_15175);
nand U15666 (N_15666,N_15427,N_15055);
and U15667 (N_15667,N_15132,N_15253);
and U15668 (N_15668,N_15473,N_15387);
nand U15669 (N_15669,N_15127,N_15442);
or U15670 (N_15670,N_15028,N_15471);
or U15671 (N_15671,N_15317,N_15485);
or U15672 (N_15672,N_15131,N_15169);
or U15673 (N_15673,N_15439,N_15493);
or U15674 (N_15674,N_15262,N_15419);
nor U15675 (N_15675,N_15104,N_15229);
nor U15676 (N_15676,N_15146,N_15085);
or U15677 (N_15677,N_15126,N_15412);
or U15678 (N_15678,N_15150,N_15393);
and U15679 (N_15679,N_15474,N_15366);
nand U15680 (N_15680,N_15275,N_15211);
nand U15681 (N_15681,N_15435,N_15199);
or U15682 (N_15682,N_15244,N_15463);
nor U15683 (N_15683,N_15074,N_15281);
or U15684 (N_15684,N_15219,N_15301);
and U15685 (N_15685,N_15249,N_15250);
xor U15686 (N_15686,N_15066,N_15335);
nor U15687 (N_15687,N_15355,N_15215);
and U15688 (N_15688,N_15234,N_15380);
nor U15689 (N_15689,N_15418,N_15002);
or U15690 (N_15690,N_15121,N_15458);
nor U15691 (N_15691,N_15277,N_15413);
or U15692 (N_15692,N_15223,N_15430);
nand U15693 (N_15693,N_15195,N_15202);
nand U15694 (N_15694,N_15044,N_15298);
nand U15695 (N_15695,N_15376,N_15035);
or U15696 (N_15696,N_15460,N_15414);
nand U15697 (N_15697,N_15354,N_15272);
or U15698 (N_15698,N_15255,N_15454);
or U15699 (N_15699,N_15420,N_15314);
or U15700 (N_15700,N_15095,N_15468);
and U15701 (N_15701,N_15377,N_15402);
and U15702 (N_15702,N_15470,N_15136);
nor U15703 (N_15703,N_15216,N_15092);
nand U15704 (N_15704,N_15067,N_15498);
nand U15705 (N_15705,N_15390,N_15036);
nand U15706 (N_15706,N_15029,N_15156);
nor U15707 (N_15707,N_15182,N_15170);
nor U15708 (N_15708,N_15389,N_15494);
nor U15709 (N_15709,N_15410,N_15451);
or U15710 (N_15710,N_15062,N_15457);
or U15711 (N_15711,N_15089,N_15151);
or U15712 (N_15712,N_15299,N_15481);
nor U15713 (N_15713,N_15422,N_15105);
nor U15714 (N_15714,N_15257,N_15447);
nor U15715 (N_15715,N_15379,N_15246);
nand U15716 (N_15716,N_15038,N_15421);
or U15717 (N_15717,N_15395,N_15411);
nand U15718 (N_15718,N_15070,N_15338);
nor U15719 (N_15719,N_15081,N_15158);
nor U15720 (N_15720,N_15032,N_15071);
nand U15721 (N_15721,N_15370,N_15371);
nor U15722 (N_15722,N_15294,N_15179);
or U15723 (N_15723,N_15270,N_15068);
or U15724 (N_15724,N_15012,N_15134);
nand U15725 (N_15725,N_15464,N_15273);
nand U15726 (N_15726,N_15350,N_15003);
nand U15727 (N_15727,N_15227,N_15312);
and U15728 (N_15728,N_15491,N_15174);
or U15729 (N_15729,N_15455,N_15237);
and U15730 (N_15730,N_15191,N_15409);
nand U15731 (N_15731,N_15426,N_15324);
or U15732 (N_15732,N_15152,N_15183);
nor U15733 (N_15733,N_15138,N_15394);
nand U15734 (N_15734,N_15147,N_15225);
or U15735 (N_15735,N_15122,N_15465);
nor U15736 (N_15736,N_15353,N_15492);
nor U15737 (N_15737,N_15239,N_15309);
nor U15738 (N_15738,N_15497,N_15142);
or U15739 (N_15739,N_15343,N_15026);
nand U15740 (N_15740,N_15437,N_15303);
nor U15741 (N_15741,N_15466,N_15214);
and U15742 (N_15742,N_15075,N_15333);
or U15743 (N_15743,N_15079,N_15375);
nand U15744 (N_15744,N_15254,N_15486);
nand U15745 (N_15745,N_15020,N_15334);
and U15746 (N_15746,N_15059,N_15245);
nand U15747 (N_15747,N_15446,N_15356);
or U15748 (N_15748,N_15213,N_15424);
nand U15749 (N_15749,N_15233,N_15489);
nor U15750 (N_15750,N_15487,N_15159);
and U15751 (N_15751,N_15055,N_15272);
or U15752 (N_15752,N_15097,N_15472);
nand U15753 (N_15753,N_15479,N_15184);
nand U15754 (N_15754,N_15022,N_15097);
or U15755 (N_15755,N_15027,N_15018);
and U15756 (N_15756,N_15373,N_15305);
nor U15757 (N_15757,N_15462,N_15265);
nand U15758 (N_15758,N_15364,N_15350);
nand U15759 (N_15759,N_15195,N_15322);
or U15760 (N_15760,N_15484,N_15002);
and U15761 (N_15761,N_15296,N_15478);
nand U15762 (N_15762,N_15325,N_15253);
nand U15763 (N_15763,N_15129,N_15465);
and U15764 (N_15764,N_15362,N_15001);
nor U15765 (N_15765,N_15274,N_15476);
nor U15766 (N_15766,N_15014,N_15375);
nor U15767 (N_15767,N_15375,N_15158);
and U15768 (N_15768,N_15148,N_15190);
and U15769 (N_15769,N_15301,N_15267);
nand U15770 (N_15770,N_15482,N_15348);
and U15771 (N_15771,N_15484,N_15258);
nor U15772 (N_15772,N_15420,N_15281);
nand U15773 (N_15773,N_15262,N_15212);
or U15774 (N_15774,N_15105,N_15328);
and U15775 (N_15775,N_15111,N_15256);
or U15776 (N_15776,N_15387,N_15383);
nand U15777 (N_15777,N_15484,N_15069);
nor U15778 (N_15778,N_15400,N_15497);
nand U15779 (N_15779,N_15273,N_15297);
nand U15780 (N_15780,N_15296,N_15450);
and U15781 (N_15781,N_15033,N_15100);
nor U15782 (N_15782,N_15246,N_15005);
nand U15783 (N_15783,N_15060,N_15350);
and U15784 (N_15784,N_15272,N_15019);
nor U15785 (N_15785,N_15297,N_15203);
and U15786 (N_15786,N_15011,N_15206);
nand U15787 (N_15787,N_15200,N_15271);
nand U15788 (N_15788,N_15242,N_15402);
nor U15789 (N_15789,N_15461,N_15106);
and U15790 (N_15790,N_15116,N_15370);
and U15791 (N_15791,N_15027,N_15194);
nand U15792 (N_15792,N_15116,N_15088);
nand U15793 (N_15793,N_15018,N_15330);
or U15794 (N_15794,N_15176,N_15454);
and U15795 (N_15795,N_15029,N_15123);
and U15796 (N_15796,N_15103,N_15042);
or U15797 (N_15797,N_15317,N_15140);
nand U15798 (N_15798,N_15074,N_15327);
or U15799 (N_15799,N_15251,N_15267);
and U15800 (N_15800,N_15368,N_15126);
nand U15801 (N_15801,N_15159,N_15028);
xor U15802 (N_15802,N_15371,N_15154);
nand U15803 (N_15803,N_15478,N_15271);
nand U15804 (N_15804,N_15073,N_15365);
or U15805 (N_15805,N_15348,N_15330);
nand U15806 (N_15806,N_15123,N_15385);
and U15807 (N_15807,N_15135,N_15452);
nand U15808 (N_15808,N_15248,N_15345);
or U15809 (N_15809,N_15333,N_15497);
and U15810 (N_15810,N_15288,N_15467);
nand U15811 (N_15811,N_15353,N_15082);
nand U15812 (N_15812,N_15204,N_15344);
or U15813 (N_15813,N_15156,N_15253);
or U15814 (N_15814,N_15067,N_15084);
or U15815 (N_15815,N_15273,N_15392);
and U15816 (N_15816,N_15113,N_15470);
nand U15817 (N_15817,N_15464,N_15007);
nand U15818 (N_15818,N_15045,N_15218);
nand U15819 (N_15819,N_15490,N_15229);
or U15820 (N_15820,N_15438,N_15365);
or U15821 (N_15821,N_15442,N_15011);
nand U15822 (N_15822,N_15365,N_15203);
or U15823 (N_15823,N_15009,N_15114);
nand U15824 (N_15824,N_15097,N_15277);
and U15825 (N_15825,N_15035,N_15075);
or U15826 (N_15826,N_15374,N_15209);
and U15827 (N_15827,N_15483,N_15271);
nand U15828 (N_15828,N_15004,N_15104);
nor U15829 (N_15829,N_15056,N_15277);
nand U15830 (N_15830,N_15396,N_15466);
xor U15831 (N_15831,N_15474,N_15166);
nor U15832 (N_15832,N_15250,N_15438);
and U15833 (N_15833,N_15105,N_15234);
nor U15834 (N_15834,N_15060,N_15014);
nor U15835 (N_15835,N_15427,N_15305);
or U15836 (N_15836,N_15201,N_15276);
and U15837 (N_15837,N_15295,N_15048);
and U15838 (N_15838,N_15296,N_15260);
or U15839 (N_15839,N_15381,N_15399);
nand U15840 (N_15840,N_15142,N_15103);
nor U15841 (N_15841,N_15255,N_15253);
nor U15842 (N_15842,N_15370,N_15283);
nor U15843 (N_15843,N_15225,N_15046);
nor U15844 (N_15844,N_15276,N_15154);
or U15845 (N_15845,N_15370,N_15105);
nor U15846 (N_15846,N_15320,N_15038);
nand U15847 (N_15847,N_15321,N_15119);
nand U15848 (N_15848,N_15354,N_15195);
nor U15849 (N_15849,N_15299,N_15291);
nor U15850 (N_15850,N_15248,N_15037);
nor U15851 (N_15851,N_15268,N_15346);
nand U15852 (N_15852,N_15329,N_15449);
nand U15853 (N_15853,N_15267,N_15158);
and U15854 (N_15854,N_15282,N_15129);
nand U15855 (N_15855,N_15240,N_15268);
nand U15856 (N_15856,N_15412,N_15461);
nor U15857 (N_15857,N_15333,N_15139);
and U15858 (N_15858,N_15122,N_15323);
nand U15859 (N_15859,N_15047,N_15480);
and U15860 (N_15860,N_15133,N_15336);
or U15861 (N_15861,N_15005,N_15096);
or U15862 (N_15862,N_15397,N_15058);
nand U15863 (N_15863,N_15480,N_15358);
nor U15864 (N_15864,N_15472,N_15055);
and U15865 (N_15865,N_15131,N_15075);
or U15866 (N_15866,N_15222,N_15128);
and U15867 (N_15867,N_15449,N_15423);
or U15868 (N_15868,N_15385,N_15382);
and U15869 (N_15869,N_15049,N_15175);
nor U15870 (N_15870,N_15155,N_15082);
and U15871 (N_15871,N_15358,N_15251);
or U15872 (N_15872,N_15164,N_15013);
nand U15873 (N_15873,N_15109,N_15499);
nor U15874 (N_15874,N_15282,N_15031);
and U15875 (N_15875,N_15383,N_15492);
nor U15876 (N_15876,N_15049,N_15345);
or U15877 (N_15877,N_15083,N_15309);
nor U15878 (N_15878,N_15015,N_15088);
nor U15879 (N_15879,N_15261,N_15446);
and U15880 (N_15880,N_15234,N_15284);
and U15881 (N_15881,N_15162,N_15144);
nor U15882 (N_15882,N_15271,N_15076);
and U15883 (N_15883,N_15432,N_15453);
and U15884 (N_15884,N_15002,N_15358);
nor U15885 (N_15885,N_15102,N_15367);
and U15886 (N_15886,N_15197,N_15202);
and U15887 (N_15887,N_15389,N_15056);
or U15888 (N_15888,N_15178,N_15381);
nor U15889 (N_15889,N_15082,N_15397);
nor U15890 (N_15890,N_15118,N_15397);
nor U15891 (N_15891,N_15457,N_15263);
nand U15892 (N_15892,N_15328,N_15128);
or U15893 (N_15893,N_15234,N_15266);
nand U15894 (N_15894,N_15035,N_15150);
or U15895 (N_15895,N_15488,N_15331);
nand U15896 (N_15896,N_15166,N_15420);
nor U15897 (N_15897,N_15444,N_15447);
xnor U15898 (N_15898,N_15256,N_15076);
and U15899 (N_15899,N_15250,N_15308);
nor U15900 (N_15900,N_15167,N_15198);
nor U15901 (N_15901,N_15047,N_15413);
and U15902 (N_15902,N_15146,N_15005);
nor U15903 (N_15903,N_15000,N_15145);
nor U15904 (N_15904,N_15239,N_15330);
nand U15905 (N_15905,N_15446,N_15030);
nand U15906 (N_15906,N_15307,N_15347);
or U15907 (N_15907,N_15309,N_15049);
and U15908 (N_15908,N_15374,N_15335);
nand U15909 (N_15909,N_15221,N_15220);
and U15910 (N_15910,N_15169,N_15330);
or U15911 (N_15911,N_15365,N_15007);
nor U15912 (N_15912,N_15259,N_15147);
nand U15913 (N_15913,N_15448,N_15319);
and U15914 (N_15914,N_15428,N_15440);
nand U15915 (N_15915,N_15338,N_15418);
and U15916 (N_15916,N_15264,N_15361);
nand U15917 (N_15917,N_15030,N_15040);
nand U15918 (N_15918,N_15485,N_15264);
and U15919 (N_15919,N_15002,N_15071);
and U15920 (N_15920,N_15346,N_15246);
or U15921 (N_15921,N_15204,N_15270);
nand U15922 (N_15922,N_15481,N_15148);
nor U15923 (N_15923,N_15122,N_15088);
nor U15924 (N_15924,N_15223,N_15158);
or U15925 (N_15925,N_15463,N_15253);
and U15926 (N_15926,N_15188,N_15120);
or U15927 (N_15927,N_15270,N_15217);
nor U15928 (N_15928,N_15285,N_15027);
and U15929 (N_15929,N_15173,N_15482);
nand U15930 (N_15930,N_15150,N_15448);
nor U15931 (N_15931,N_15179,N_15414);
and U15932 (N_15932,N_15181,N_15125);
nand U15933 (N_15933,N_15261,N_15057);
nand U15934 (N_15934,N_15344,N_15085);
nand U15935 (N_15935,N_15205,N_15166);
or U15936 (N_15936,N_15447,N_15392);
or U15937 (N_15937,N_15223,N_15231);
nand U15938 (N_15938,N_15444,N_15288);
and U15939 (N_15939,N_15300,N_15215);
nor U15940 (N_15940,N_15302,N_15074);
or U15941 (N_15941,N_15420,N_15263);
nor U15942 (N_15942,N_15404,N_15245);
nor U15943 (N_15943,N_15137,N_15037);
and U15944 (N_15944,N_15147,N_15341);
and U15945 (N_15945,N_15215,N_15364);
and U15946 (N_15946,N_15230,N_15051);
and U15947 (N_15947,N_15209,N_15196);
and U15948 (N_15948,N_15319,N_15470);
or U15949 (N_15949,N_15433,N_15102);
nor U15950 (N_15950,N_15106,N_15250);
nand U15951 (N_15951,N_15117,N_15372);
and U15952 (N_15952,N_15482,N_15236);
nor U15953 (N_15953,N_15059,N_15088);
nor U15954 (N_15954,N_15111,N_15204);
or U15955 (N_15955,N_15005,N_15378);
and U15956 (N_15956,N_15009,N_15101);
or U15957 (N_15957,N_15205,N_15091);
and U15958 (N_15958,N_15247,N_15263);
nor U15959 (N_15959,N_15032,N_15308);
and U15960 (N_15960,N_15011,N_15204);
nand U15961 (N_15961,N_15333,N_15104);
nand U15962 (N_15962,N_15135,N_15127);
and U15963 (N_15963,N_15275,N_15003);
xnor U15964 (N_15964,N_15480,N_15207);
or U15965 (N_15965,N_15493,N_15399);
and U15966 (N_15966,N_15449,N_15471);
or U15967 (N_15967,N_15476,N_15266);
nand U15968 (N_15968,N_15009,N_15193);
nor U15969 (N_15969,N_15379,N_15089);
nand U15970 (N_15970,N_15116,N_15211);
and U15971 (N_15971,N_15044,N_15045);
or U15972 (N_15972,N_15107,N_15316);
nor U15973 (N_15973,N_15213,N_15043);
nor U15974 (N_15974,N_15138,N_15055);
or U15975 (N_15975,N_15237,N_15080);
or U15976 (N_15976,N_15104,N_15446);
or U15977 (N_15977,N_15253,N_15356);
or U15978 (N_15978,N_15468,N_15407);
and U15979 (N_15979,N_15375,N_15377);
nor U15980 (N_15980,N_15197,N_15267);
nand U15981 (N_15981,N_15116,N_15033);
or U15982 (N_15982,N_15232,N_15405);
nand U15983 (N_15983,N_15372,N_15158);
nor U15984 (N_15984,N_15031,N_15384);
and U15985 (N_15985,N_15133,N_15234);
or U15986 (N_15986,N_15024,N_15302);
or U15987 (N_15987,N_15083,N_15419);
and U15988 (N_15988,N_15328,N_15014);
nand U15989 (N_15989,N_15074,N_15408);
nor U15990 (N_15990,N_15079,N_15492);
or U15991 (N_15991,N_15376,N_15350);
nor U15992 (N_15992,N_15445,N_15033);
nand U15993 (N_15993,N_15266,N_15185);
nor U15994 (N_15994,N_15021,N_15497);
nor U15995 (N_15995,N_15102,N_15407);
and U15996 (N_15996,N_15327,N_15312);
and U15997 (N_15997,N_15219,N_15161);
nand U15998 (N_15998,N_15371,N_15434);
nand U15999 (N_15999,N_15300,N_15190);
and U16000 (N_16000,N_15531,N_15989);
or U16001 (N_16001,N_15879,N_15836);
xnor U16002 (N_16002,N_15930,N_15596);
and U16003 (N_16003,N_15784,N_15783);
nor U16004 (N_16004,N_15929,N_15740);
nor U16005 (N_16005,N_15881,N_15914);
or U16006 (N_16006,N_15671,N_15703);
nor U16007 (N_16007,N_15593,N_15757);
nor U16008 (N_16008,N_15534,N_15754);
or U16009 (N_16009,N_15667,N_15672);
and U16010 (N_16010,N_15715,N_15705);
nor U16011 (N_16011,N_15562,N_15964);
nor U16012 (N_16012,N_15931,N_15857);
nor U16013 (N_16013,N_15779,N_15641);
nand U16014 (N_16014,N_15628,N_15732);
nand U16015 (N_16015,N_15785,N_15695);
nand U16016 (N_16016,N_15884,N_15626);
or U16017 (N_16017,N_15828,N_15977);
and U16018 (N_16018,N_15567,N_15823);
nand U16019 (N_16019,N_15553,N_15690);
or U16020 (N_16020,N_15699,N_15860);
nor U16021 (N_16021,N_15882,N_15900);
nand U16022 (N_16022,N_15706,N_15662);
nand U16023 (N_16023,N_15885,N_15565);
nor U16024 (N_16024,N_15536,N_15513);
or U16025 (N_16025,N_15861,N_15502);
nand U16026 (N_16026,N_15877,N_15687);
nand U16027 (N_16027,N_15739,N_15846);
and U16028 (N_16028,N_15507,N_15741);
nand U16029 (N_16029,N_15800,N_15924);
nor U16030 (N_16030,N_15995,N_15589);
and U16031 (N_16031,N_15891,N_15901);
nand U16032 (N_16032,N_15804,N_15708);
nand U16033 (N_16033,N_15813,N_15718);
nand U16034 (N_16034,N_15988,N_15967);
nor U16035 (N_16035,N_15873,N_15645);
or U16036 (N_16036,N_15985,N_15782);
and U16037 (N_16037,N_15932,N_15610);
nand U16038 (N_16038,N_15738,N_15733);
or U16039 (N_16039,N_15509,N_15862);
or U16040 (N_16040,N_15642,N_15527);
nor U16041 (N_16041,N_15643,N_15834);
or U16042 (N_16042,N_15632,N_15523);
nand U16043 (N_16043,N_15910,N_15570);
and U16044 (N_16044,N_15559,N_15716);
nand U16045 (N_16045,N_15717,N_15844);
and U16046 (N_16046,N_15994,N_15811);
or U16047 (N_16047,N_15637,N_15809);
nor U16048 (N_16048,N_15826,N_15919);
or U16049 (N_16049,N_15743,N_15688);
nor U16050 (N_16050,N_15710,N_15630);
nor U16051 (N_16051,N_15923,N_15530);
nand U16052 (N_16052,N_15617,N_15801);
or U16053 (N_16053,N_15638,N_15902);
nor U16054 (N_16054,N_15624,N_15622);
and U16055 (N_16055,N_15868,N_15878);
nor U16056 (N_16056,N_15808,N_15554);
nand U16057 (N_16057,N_15555,N_15729);
and U16058 (N_16058,N_15609,N_15944);
nand U16059 (N_16059,N_15971,N_15519);
nor U16060 (N_16060,N_15912,N_15665);
or U16061 (N_16061,N_15763,N_15533);
or U16062 (N_16062,N_15723,N_15520);
or U16063 (N_16063,N_15942,N_15604);
nor U16064 (N_16064,N_15817,N_15644);
and U16065 (N_16065,N_15598,N_15963);
and U16066 (N_16066,N_15529,N_15922);
or U16067 (N_16067,N_15854,N_15525);
nor U16068 (N_16068,N_15939,N_15669);
or U16069 (N_16069,N_15684,N_15657);
nand U16070 (N_16070,N_15611,N_15550);
and U16071 (N_16071,N_15949,N_15731);
or U16072 (N_16072,N_15522,N_15915);
and U16073 (N_16073,N_15750,N_15670);
or U16074 (N_16074,N_15864,N_15614);
or U16075 (N_16075,N_15872,N_15543);
or U16076 (N_16076,N_15696,N_15500);
nor U16077 (N_16077,N_15874,N_15558);
nand U16078 (N_16078,N_15505,N_15560);
nor U16079 (N_16079,N_15992,N_15581);
xor U16080 (N_16080,N_15655,N_15962);
and U16081 (N_16081,N_15906,N_15579);
or U16082 (N_16082,N_15574,N_15587);
and U16083 (N_16083,N_15749,N_15982);
nand U16084 (N_16084,N_15504,N_15952);
and U16085 (N_16085,N_15659,N_15875);
and U16086 (N_16086,N_15585,N_15786);
or U16087 (N_16087,N_15548,N_15721);
nor U16088 (N_16088,N_15599,N_15755);
nand U16089 (N_16089,N_15858,N_15805);
or U16090 (N_16090,N_15516,N_15871);
nor U16091 (N_16091,N_15905,N_15851);
or U16092 (N_16092,N_15578,N_15742);
nor U16093 (N_16093,N_15896,N_15594);
and U16094 (N_16094,N_15815,N_15595);
or U16095 (N_16095,N_15756,N_15908);
or U16096 (N_16096,N_15893,N_15541);
nor U16097 (N_16097,N_15724,N_15676);
nand U16098 (N_16098,N_15955,N_15656);
nand U16099 (N_16099,N_15794,N_15921);
or U16100 (N_16100,N_15532,N_15650);
nor U16101 (N_16101,N_15627,N_15573);
or U16102 (N_16102,N_15652,N_15907);
xor U16103 (N_16103,N_15762,N_15827);
and U16104 (N_16104,N_15588,N_15678);
or U16105 (N_16105,N_15692,N_15897);
nor U16106 (N_16106,N_15661,N_15545);
or U16107 (N_16107,N_15673,N_15984);
nor U16108 (N_16108,N_15727,N_15658);
nor U16109 (N_16109,N_15797,N_15728);
nor U16110 (N_16110,N_15748,N_15904);
and U16111 (N_16111,N_15528,N_15584);
and U16112 (N_16112,N_15777,N_15586);
nor U16113 (N_16113,N_15601,N_15890);
or U16114 (N_16114,N_15653,N_15538);
and U16115 (N_16115,N_15772,N_15590);
nand U16116 (N_16116,N_15713,N_15856);
and U16117 (N_16117,N_15842,N_15758);
and U16118 (N_16118,N_15937,N_15737);
nor U16119 (N_16119,N_15987,N_15966);
or U16120 (N_16120,N_15761,N_15978);
nand U16121 (N_16121,N_15830,N_15511);
nand U16122 (N_16122,N_15566,N_15768);
and U16123 (N_16123,N_15950,N_15799);
and U16124 (N_16124,N_15870,N_15824);
or U16125 (N_16125,N_15773,N_15818);
nand U16126 (N_16126,N_15843,N_15747);
nor U16127 (N_16127,N_15654,N_15795);
and U16128 (N_16128,N_15746,N_15577);
nand U16129 (N_16129,N_15973,N_15814);
nor U16130 (N_16130,N_15635,N_15936);
nor U16131 (N_16131,N_15689,N_15898);
or U16132 (N_16132,N_15668,N_15927);
or U16133 (N_16133,N_15569,N_15619);
nor U16134 (N_16134,N_15582,N_15576);
or U16135 (N_16135,N_15677,N_15865);
nand U16136 (N_16136,N_15888,N_15568);
nor U16137 (N_16137,N_15549,N_15557);
nand U16138 (N_16138,N_15765,N_15709);
nand U16139 (N_16139,N_15852,N_15833);
or U16140 (N_16140,N_15680,N_15951);
nand U16141 (N_16141,N_15928,N_15956);
and U16142 (N_16142,N_15615,N_15542);
or U16143 (N_16143,N_15869,N_15701);
nand U16144 (N_16144,N_15970,N_15957);
or U16145 (N_16145,N_15894,N_15606);
and U16146 (N_16146,N_15938,N_15810);
and U16147 (N_16147,N_15802,N_15774);
nand U16148 (N_16148,N_15521,N_15564);
and U16149 (N_16149,N_15796,N_15691);
or U16150 (N_16150,N_15580,N_15744);
or U16151 (N_16151,N_15812,N_15625);
nand U16152 (N_16152,N_15838,N_15524);
nand U16153 (N_16153,N_15946,N_15997);
nor U16154 (N_16154,N_15648,N_15698);
and U16155 (N_16155,N_15736,N_15603);
nand U16156 (N_16156,N_15633,N_15993);
and U16157 (N_16157,N_15849,N_15892);
nand U16158 (N_16158,N_15848,N_15620);
or U16159 (N_16159,N_15730,N_15602);
or U16160 (N_16160,N_15674,N_15518);
nor U16161 (N_16161,N_15623,N_15702);
and U16162 (N_16162,N_15693,N_15751);
nand U16163 (N_16163,N_15621,N_15798);
and U16164 (N_16164,N_15839,N_15972);
and U16165 (N_16165,N_15734,N_15612);
and U16166 (N_16166,N_15776,N_15613);
or U16167 (N_16167,N_15816,N_15537);
and U16168 (N_16168,N_15781,N_15954);
nand U16169 (N_16169,N_15778,N_15822);
nor U16170 (N_16170,N_15788,N_15859);
nor U16171 (N_16171,N_15685,N_15913);
and U16172 (N_16172,N_15980,N_15832);
and U16173 (N_16173,N_15845,N_15974);
nand U16174 (N_16174,N_15510,N_15683);
and U16175 (N_16175,N_15968,N_15686);
or U16176 (N_16176,N_15722,N_15887);
and U16177 (N_16177,N_15792,N_15759);
and U16178 (N_16178,N_15766,N_15789);
and U16179 (N_16179,N_15681,N_15556);
or U16180 (N_16180,N_15600,N_15629);
and U16181 (N_16181,N_15547,N_15965);
nand U16182 (N_16182,N_15835,N_15508);
nand U16183 (N_16183,N_15666,N_15517);
nor U16184 (N_16184,N_15847,N_15597);
and U16185 (N_16185,N_15506,N_15959);
nand U16186 (N_16186,N_15821,N_15917);
nand U16187 (N_16187,N_15990,N_15775);
nor U16188 (N_16188,N_15618,N_15933);
or U16189 (N_16189,N_15960,N_15753);
nand U16190 (N_16190,N_15840,N_15935);
or U16191 (N_16191,N_15694,N_15712);
nand U16192 (N_16192,N_15720,N_15704);
or U16193 (N_16193,N_15501,N_15679);
nor U16194 (N_16194,N_15918,N_15876);
or U16195 (N_16195,N_15941,N_15855);
nor U16196 (N_16196,N_15850,N_15714);
nor U16197 (N_16197,N_15640,N_15735);
or U16198 (N_16198,N_15526,N_15790);
or U16199 (N_16199,N_15675,N_15976);
or U16200 (N_16200,N_15634,N_15719);
or U16201 (N_16201,N_15911,N_15945);
and U16202 (N_16202,N_15646,N_15663);
nand U16203 (N_16203,N_15592,N_15969);
or U16204 (N_16204,N_15803,N_15660);
or U16205 (N_16205,N_15707,N_15991);
or U16206 (N_16206,N_15607,N_15769);
or U16207 (N_16207,N_15540,N_15571);
and U16208 (N_16208,N_15867,N_15866);
and U16209 (N_16209,N_15764,N_15700);
and U16210 (N_16210,N_15975,N_15711);
and U16211 (N_16211,N_15787,N_15725);
nand U16212 (N_16212,N_15649,N_15880);
nor U16213 (N_16213,N_15591,N_15934);
or U16214 (N_16214,N_15979,N_15983);
and U16215 (N_16215,N_15544,N_15682);
nand U16216 (N_16216,N_15886,N_15793);
nor U16217 (N_16217,N_15503,N_15639);
or U16218 (N_16218,N_15535,N_15752);
or U16219 (N_16219,N_15961,N_15999);
nand U16220 (N_16220,N_15998,N_15605);
nor U16221 (N_16221,N_15981,N_15561);
xnor U16222 (N_16222,N_15883,N_15512);
nand U16223 (N_16223,N_15770,N_15780);
or U16224 (N_16224,N_15583,N_15943);
or U16225 (N_16225,N_15926,N_15948);
and U16226 (N_16226,N_15925,N_15515);
nor U16227 (N_16227,N_15841,N_15760);
nor U16228 (N_16228,N_15909,N_15899);
nand U16229 (N_16229,N_15771,N_15551);
nor U16230 (N_16230,N_15825,N_15889);
nand U16231 (N_16231,N_15575,N_15837);
nand U16232 (N_16232,N_15996,N_15791);
nor U16233 (N_16233,N_15651,N_15953);
nor U16234 (N_16234,N_15829,N_15958);
or U16235 (N_16235,N_15552,N_15916);
nor U16236 (N_16236,N_15986,N_15546);
nand U16237 (N_16237,N_15697,N_15863);
nand U16238 (N_16238,N_15726,N_15745);
and U16239 (N_16239,N_15831,N_15647);
nand U16240 (N_16240,N_15940,N_15820);
and U16241 (N_16241,N_15806,N_15819);
nand U16242 (N_16242,N_15853,N_15920);
and U16243 (N_16243,N_15767,N_15616);
nand U16244 (N_16244,N_15514,N_15664);
nor U16245 (N_16245,N_15572,N_15539);
nor U16246 (N_16246,N_15903,N_15631);
nand U16247 (N_16247,N_15563,N_15636);
nor U16248 (N_16248,N_15895,N_15947);
and U16249 (N_16249,N_15807,N_15608);
nor U16250 (N_16250,N_15539,N_15538);
nor U16251 (N_16251,N_15803,N_15763);
nand U16252 (N_16252,N_15994,N_15797);
or U16253 (N_16253,N_15519,N_15692);
or U16254 (N_16254,N_15712,N_15795);
nor U16255 (N_16255,N_15999,N_15545);
and U16256 (N_16256,N_15745,N_15536);
and U16257 (N_16257,N_15517,N_15583);
or U16258 (N_16258,N_15683,N_15701);
and U16259 (N_16259,N_15656,N_15997);
nor U16260 (N_16260,N_15572,N_15622);
or U16261 (N_16261,N_15875,N_15980);
nor U16262 (N_16262,N_15631,N_15675);
nor U16263 (N_16263,N_15826,N_15845);
nand U16264 (N_16264,N_15907,N_15837);
nor U16265 (N_16265,N_15601,N_15514);
nor U16266 (N_16266,N_15984,N_15566);
or U16267 (N_16267,N_15902,N_15558);
and U16268 (N_16268,N_15597,N_15532);
nor U16269 (N_16269,N_15984,N_15543);
and U16270 (N_16270,N_15640,N_15743);
or U16271 (N_16271,N_15864,N_15884);
nand U16272 (N_16272,N_15634,N_15693);
nor U16273 (N_16273,N_15977,N_15996);
or U16274 (N_16274,N_15788,N_15714);
or U16275 (N_16275,N_15540,N_15676);
nand U16276 (N_16276,N_15908,N_15864);
and U16277 (N_16277,N_15935,N_15730);
or U16278 (N_16278,N_15716,N_15948);
nand U16279 (N_16279,N_15775,N_15815);
nor U16280 (N_16280,N_15941,N_15992);
nand U16281 (N_16281,N_15735,N_15818);
and U16282 (N_16282,N_15969,N_15693);
or U16283 (N_16283,N_15618,N_15949);
or U16284 (N_16284,N_15719,N_15661);
nor U16285 (N_16285,N_15872,N_15592);
and U16286 (N_16286,N_15645,N_15508);
or U16287 (N_16287,N_15597,N_15856);
nor U16288 (N_16288,N_15638,N_15541);
or U16289 (N_16289,N_15702,N_15703);
or U16290 (N_16290,N_15949,N_15856);
nor U16291 (N_16291,N_15528,N_15906);
nand U16292 (N_16292,N_15874,N_15720);
nor U16293 (N_16293,N_15973,N_15666);
nand U16294 (N_16294,N_15630,N_15546);
or U16295 (N_16295,N_15737,N_15612);
and U16296 (N_16296,N_15996,N_15533);
and U16297 (N_16297,N_15685,N_15876);
nand U16298 (N_16298,N_15749,N_15990);
or U16299 (N_16299,N_15548,N_15555);
or U16300 (N_16300,N_15872,N_15985);
nor U16301 (N_16301,N_15616,N_15935);
or U16302 (N_16302,N_15884,N_15881);
or U16303 (N_16303,N_15755,N_15592);
or U16304 (N_16304,N_15781,N_15596);
nor U16305 (N_16305,N_15916,N_15582);
or U16306 (N_16306,N_15904,N_15641);
nand U16307 (N_16307,N_15717,N_15823);
and U16308 (N_16308,N_15581,N_15518);
or U16309 (N_16309,N_15702,N_15934);
xnor U16310 (N_16310,N_15581,N_15861);
nand U16311 (N_16311,N_15772,N_15845);
or U16312 (N_16312,N_15705,N_15506);
or U16313 (N_16313,N_15951,N_15578);
or U16314 (N_16314,N_15604,N_15714);
nor U16315 (N_16315,N_15554,N_15667);
nor U16316 (N_16316,N_15572,N_15779);
xor U16317 (N_16317,N_15926,N_15600);
nor U16318 (N_16318,N_15804,N_15706);
or U16319 (N_16319,N_15771,N_15953);
nor U16320 (N_16320,N_15526,N_15606);
or U16321 (N_16321,N_15937,N_15652);
and U16322 (N_16322,N_15702,N_15655);
nor U16323 (N_16323,N_15683,N_15781);
and U16324 (N_16324,N_15534,N_15541);
or U16325 (N_16325,N_15520,N_15857);
and U16326 (N_16326,N_15859,N_15836);
nand U16327 (N_16327,N_15762,N_15809);
nor U16328 (N_16328,N_15645,N_15617);
and U16329 (N_16329,N_15867,N_15587);
and U16330 (N_16330,N_15759,N_15572);
nor U16331 (N_16331,N_15549,N_15564);
or U16332 (N_16332,N_15570,N_15974);
nand U16333 (N_16333,N_15690,N_15662);
nor U16334 (N_16334,N_15942,N_15905);
or U16335 (N_16335,N_15912,N_15834);
and U16336 (N_16336,N_15992,N_15926);
and U16337 (N_16337,N_15564,N_15662);
or U16338 (N_16338,N_15943,N_15820);
nand U16339 (N_16339,N_15576,N_15820);
and U16340 (N_16340,N_15557,N_15659);
nor U16341 (N_16341,N_15725,N_15898);
nand U16342 (N_16342,N_15734,N_15780);
and U16343 (N_16343,N_15778,N_15706);
nor U16344 (N_16344,N_15558,N_15840);
or U16345 (N_16345,N_15873,N_15949);
or U16346 (N_16346,N_15981,N_15774);
nand U16347 (N_16347,N_15633,N_15695);
nand U16348 (N_16348,N_15606,N_15703);
xnor U16349 (N_16349,N_15800,N_15754);
or U16350 (N_16350,N_15979,N_15541);
or U16351 (N_16351,N_15569,N_15500);
nor U16352 (N_16352,N_15959,N_15765);
nor U16353 (N_16353,N_15726,N_15733);
and U16354 (N_16354,N_15741,N_15555);
or U16355 (N_16355,N_15793,N_15524);
nand U16356 (N_16356,N_15710,N_15816);
and U16357 (N_16357,N_15899,N_15790);
nand U16358 (N_16358,N_15512,N_15599);
nand U16359 (N_16359,N_15936,N_15718);
nor U16360 (N_16360,N_15777,N_15505);
or U16361 (N_16361,N_15631,N_15751);
or U16362 (N_16362,N_15555,N_15549);
or U16363 (N_16363,N_15849,N_15857);
nand U16364 (N_16364,N_15775,N_15741);
or U16365 (N_16365,N_15954,N_15555);
and U16366 (N_16366,N_15759,N_15857);
nand U16367 (N_16367,N_15639,N_15658);
or U16368 (N_16368,N_15517,N_15644);
nor U16369 (N_16369,N_15805,N_15861);
or U16370 (N_16370,N_15541,N_15676);
and U16371 (N_16371,N_15669,N_15626);
nand U16372 (N_16372,N_15506,N_15914);
and U16373 (N_16373,N_15591,N_15901);
nand U16374 (N_16374,N_15701,N_15594);
nor U16375 (N_16375,N_15572,N_15647);
nand U16376 (N_16376,N_15875,N_15672);
or U16377 (N_16377,N_15510,N_15524);
nand U16378 (N_16378,N_15508,N_15830);
nor U16379 (N_16379,N_15645,N_15532);
and U16380 (N_16380,N_15764,N_15938);
nand U16381 (N_16381,N_15933,N_15729);
xor U16382 (N_16382,N_15902,N_15746);
nor U16383 (N_16383,N_15821,N_15720);
and U16384 (N_16384,N_15765,N_15895);
nand U16385 (N_16385,N_15759,N_15886);
or U16386 (N_16386,N_15500,N_15671);
and U16387 (N_16387,N_15602,N_15870);
or U16388 (N_16388,N_15700,N_15603);
nor U16389 (N_16389,N_15757,N_15687);
or U16390 (N_16390,N_15959,N_15553);
or U16391 (N_16391,N_15655,N_15639);
or U16392 (N_16392,N_15631,N_15599);
nand U16393 (N_16393,N_15794,N_15600);
nand U16394 (N_16394,N_15893,N_15701);
or U16395 (N_16395,N_15836,N_15795);
nand U16396 (N_16396,N_15608,N_15916);
or U16397 (N_16397,N_15819,N_15709);
nand U16398 (N_16398,N_15786,N_15855);
nand U16399 (N_16399,N_15865,N_15920);
nand U16400 (N_16400,N_15902,N_15660);
nand U16401 (N_16401,N_15640,N_15950);
nor U16402 (N_16402,N_15645,N_15598);
nor U16403 (N_16403,N_15990,N_15903);
and U16404 (N_16404,N_15615,N_15898);
nand U16405 (N_16405,N_15876,N_15880);
xnor U16406 (N_16406,N_15610,N_15891);
and U16407 (N_16407,N_15766,N_15908);
or U16408 (N_16408,N_15981,N_15581);
and U16409 (N_16409,N_15622,N_15588);
xnor U16410 (N_16410,N_15754,N_15816);
nand U16411 (N_16411,N_15544,N_15675);
nor U16412 (N_16412,N_15848,N_15557);
and U16413 (N_16413,N_15938,N_15834);
and U16414 (N_16414,N_15546,N_15919);
or U16415 (N_16415,N_15813,N_15712);
or U16416 (N_16416,N_15835,N_15620);
nand U16417 (N_16417,N_15582,N_15943);
or U16418 (N_16418,N_15648,N_15641);
nand U16419 (N_16419,N_15997,N_15596);
and U16420 (N_16420,N_15538,N_15837);
nand U16421 (N_16421,N_15700,N_15913);
and U16422 (N_16422,N_15568,N_15835);
nand U16423 (N_16423,N_15946,N_15784);
and U16424 (N_16424,N_15572,N_15739);
or U16425 (N_16425,N_15505,N_15967);
nor U16426 (N_16426,N_15928,N_15666);
and U16427 (N_16427,N_15926,N_15542);
and U16428 (N_16428,N_15594,N_15585);
or U16429 (N_16429,N_15905,N_15908);
nand U16430 (N_16430,N_15560,N_15751);
and U16431 (N_16431,N_15718,N_15755);
nor U16432 (N_16432,N_15692,N_15859);
or U16433 (N_16433,N_15684,N_15745);
nand U16434 (N_16434,N_15564,N_15737);
or U16435 (N_16435,N_15655,N_15909);
xnor U16436 (N_16436,N_15889,N_15891);
nor U16437 (N_16437,N_15789,N_15556);
nor U16438 (N_16438,N_15739,N_15505);
and U16439 (N_16439,N_15670,N_15808);
nor U16440 (N_16440,N_15719,N_15857);
nand U16441 (N_16441,N_15819,N_15637);
nand U16442 (N_16442,N_15666,N_15549);
and U16443 (N_16443,N_15861,N_15956);
and U16444 (N_16444,N_15740,N_15989);
nand U16445 (N_16445,N_15945,N_15923);
nor U16446 (N_16446,N_15867,N_15890);
or U16447 (N_16447,N_15868,N_15564);
nor U16448 (N_16448,N_15530,N_15673);
nand U16449 (N_16449,N_15758,N_15929);
nor U16450 (N_16450,N_15601,N_15798);
nor U16451 (N_16451,N_15527,N_15526);
nor U16452 (N_16452,N_15636,N_15545);
or U16453 (N_16453,N_15683,N_15504);
nor U16454 (N_16454,N_15743,N_15977);
or U16455 (N_16455,N_15866,N_15585);
or U16456 (N_16456,N_15797,N_15940);
nor U16457 (N_16457,N_15761,N_15897);
and U16458 (N_16458,N_15981,N_15583);
or U16459 (N_16459,N_15510,N_15872);
nand U16460 (N_16460,N_15840,N_15830);
nor U16461 (N_16461,N_15760,N_15815);
or U16462 (N_16462,N_15600,N_15754);
or U16463 (N_16463,N_15888,N_15998);
nand U16464 (N_16464,N_15644,N_15601);
or U16465 (N_16465,N_15761,N_15890);
or U16466 (N_16466,N_15773,N_15829);
nand U16467 (N_16467,N_15569,N_15626);
nor U16468 (N_16468,N_15895,N_15564);
and U16469 (N_16469,N_15634,N_15571);
nand U16470 (N_16470,N_15873,N_15928);
and U16471 (N_16471,N_15958,N_15567);
and U16472 (N_16472,N_15954,N_15674);
nor U16473 (N_16473,N_15991,N_15863);
nor U16474 (N_16474,N_15842,N_15600);
or U16475 (N_16475,N_15653,N_15781);
nor U16476 (N_16476,N_15763,N_15618);
or U16477 (N_16477,N_15887,N_15708);
and U16478 (N_16478,N_15959,N_15687);
nand U16479 (N_16479,N_15552,N_15721);
xor U16480 (N_16480,N_15753,N_15905);
or U16481 (N_16481,N_15835,N_15556);
nor U16482 (N_16482,N_15589,N_15685);
and U16483 (N_16483,N_15506,N_15735);
and U16484 (N_16484,N_15920,N_15518);
or U16485 (N_16485,N_15913,N_15966);
and U16486 (N_16486,N_15659,N_15655);
and U16487 (N_16487,N_15758,N_15523);
or U16488 (N_16488,N_15503,N_15615);
and U16489 (N_16489,N_15914,N_15795);
or U16490 (N_16490,N_15904,N_15544);
and U16491 (N_16491,N_15758,N_15905);
and U16492 (N_16492,N_15576,N_15987);
nor U16493 (N_16493,N_15823,N_15512);
nand U16494 (N_16494,N_15646,N_15964);
or U16495 (N_16495,N_15858,N_15633);
and U16496 (N_16496,N_15772,N_15848);
and U16497 (N_16497,N_15913,N_15932);
or U16498 (N_16498,N_15912,N_15767);
or U16499 (N_16499,N_15947,N_15827);
nand U16500 (N_16500,N_16384,N_16481);
or U16501 (N_16501,N_16498,N_16036);
nor U16502 (N_16502,N_16222,N_16361);
nor U16503 (N_16503,N_16285,N_16000);
nand U16504 (N_16504,N_16388,N_16131);
nand U16505 (N_16505,N_16349,N_16041);
or U16506 (N_16506,N_16238,N_16099);
and U16507 (N_16507,N_16400,N_16011);
and U16508 (N_16508,N_16054,N_16287);
or U16509 (N_16509,N_16134,N_16447);
or U16510 (N_16510,N_16120,N_16305);
or U16511 (N_16511,N_16040,N_16272);
nand U16512 (N_16512,N_16480,N_16090);
and U16513 (N_16513,N_16125,N_16462);
or U16514 (N_16514,N_16214,N_16242);
or U16515 (N_16515,N_16237,N_16212);
nor U16516 (N_16516,N_16248,N_16018);
and U16517 (N_16517,N_16363,N_16029);
and U16518 (N_16518,N_16316,N_16091);
nand U16519 (N_16519,N_16342,N_16383);
nor U16520 (N_16520,N_16188,N_16012);
or U16521 (N_16521,N_16302,N_16492);
nor U16522 (N_16522,N_16340,N_16149);
nand U16523 (N_16523,N_16288,N_16034);
nor U16524 (N_16524,N_16482,N_16189);
nor U16525 (N_16525,N_16405,N_16469);
or U16526 (N_16526,N_16471,N_16180);
or U16527 (N_16527,N_16087,N_16420);
and U16528 (N_16528,N_16004,N_16048);
and U16529 (N_16529,N_16357,N_16289);
nand U16530 (N_16530,N_16315,N_16419);
or U16531 (N_16531,N_16255,N_16022);
nand U16532 (N_16532,N_16110,N_16013);
or U16533 (N_16533,N_16064,N_16267);
nor U16534 (N_16534,N_16027,N_16194);
or U16535 (N_16535,N_16228,N_16275);
and U16536 (N_16536,N_16162,N_16331);
and U16537 (N_16537,N_16206,N_16006);
or U16538 (N_16538,N_16453,N_16355);
nor U16539 (N_16539,N_16367,N_16115);
nor U16540 (N_16540,N_16300,N_16283);
nor U16541 (N_16541,N_16274,N_16474);
and U16542 (N_16542,N_16106,N_16170);
or U16543 (N_16543,N_16260,N_16229);
nor U16544 (N_16544,N_16412,N_16215);
nor U16545 (N_16545,N_16205,N_16092);
and U16546 (N_16546,N_16042,N_16244);
and U16547 (N_16547,N_16010,N_16164);
nand U16548 (N_16548,N_16193,N_16485);
nand U16549 (N_16549,N_16160,N_16144);
nor U16550 (N_16550,N_16172,N_16235);
or U16551 (N_16551,N_16204,N_16026);
and U16552 (N_16552,N_16470,N_16252);
and U16553 (N_16553,N_16209,N_16381);
and U16554 (N_16554,N_16208,N_16352);
nor U16555 (N_16555,N_16119,N_16455);
nand U16556 (N_16556,N_16479,N_16397);
or U16557 (N_16557,N_16117,N_16491);
nor U16558 (N_16558,N_16246,N_16376);
nand U16559 (N_16559,N_16251,N_16063);
nor U16560 (N_16560,N_16114,N_16416);
and U16561 (N_16561,N_16444,N_16152);
or U16562 (N_16562,N_16016,N_16337);
nor U16563 (N_16563,N_16043,N_16279);
and U16564 (N_16564,N_16123,N_16418);
or U16565 (N_16565,N_16486,N_16053);
nor U16566 (N_16566,N_16135,N_16295);
and U16567 (N_16567,N_16145,N_16313);
or U16568 (N_16568,N_16232,N_16058);
and U16569 (N_16569,N_16408,N_16192);
nand U16570 (N_16570,N_16231,N_16296);
nand U16571 (N_16571,N_16067,N_16415);
or U16572 (N_16572,N_16157,N_16037);
or U16573 (N_16573,N_16055,N_16345);
or U16574 (N_16574,N_16306,N_16464);
nor U16575 (N_16575,N_16032,N_16326);
nand U16576 (N_16576,N_16082,N_16049);
or U16577 (N_16577,N_16264,N_16089);
or U16578 (N_16578,N_16068,N_16050);
or U16579 (N_16579,N_16138,N_16143);
or U16580 (N_16580,N_16404,N_16395);
and U16581 (N_16581,N_16377,N_16278);
and U16582 (N_16582,N_16309,N_16387);
nor U16583 (N_16583,N_16406,N_16052);
nor U16584 (N_16584,N_16496,N_16182);
or U16585 (N_16585,N_16371,N_16107);
nand U16586 (N_16586,N_16488,N_16028);
or U16587 (N_16587,N_16450,N_16359);
and U16588 (N_16588,N_16437,N_16184);
or U16589 (N_16589,N_16439,N_16169);
or U16590 (N_16590,N_16066,N_16247);
or U16591 (N_16591,N_16465,N_16324);
or U16592 (N_16592,N_16211,N_16057);
nor U16593 (N_16593,N_16281,N_16276);
nand U16594 (N_16594,N_16241,N_16171);
nor U16595 (N_16595,N_16038,N_16103);
or U16596 (N_16596,N_16213,N_16088);
nor U16597 (N_16597,N_16105,N_16176);
or U16598 (N_16598,N_16128,N_16391);
nand U16599 (N_16599,N_16097,N_16158);
nor U16600 (N_16600,N_16432,N_16239);
or U16601 (N_16601,N_16298,N_16060);
or U16602 (N_16602,N_16452,N_16258);
nand U16603 (N_16603,N_16219,N_16148);
and U16604 (N_16604,N_16023,N_16291);
or U16605 (N_16605,N_16421,N_16257);
nand U16606 (N_16606,N_16449,N_16111);
nor U16607 (N_16607,N_16254,N_16159);
and U16608 (N_16608,N_16348,N_16059);
nand U16609 (N_16609,N_16327,N_16095);
or U16610 (N_16610,N_16407,N_16424);
nor U16611 (N_16611,N_16003,N_16386);
and U16612 (N_16612,N_16070,N_16451);
or U16613 (N_16613,N_16354,N_16270);
nand U16614 (N_16614,N_16015,N_16303);
nand U16615 (N_16615,N_16085,N_16375);
and U16616 (N_16616,N_16227,N_16165);
nand U16617 (N_16617,N_16428,N_16382);
and U16618 (N_16618,N_16147,N_16071);
nor U16619 (N_16619,N_16173,N_16021);
or U16620 (N_16620,N_16445,N_16044);
nand U16621 (N_16621,N_16234,N_16366);
or U16622 (N_16622,N_16250,N_16207);
nand U16623 (N_16623,N_16033,N_16369);
nand U16624 (N_16624,N_16132,N_16456);
nor U16625 (N_16625,N_16061,N_16435);
and U16626 (N_16626,N_16423,N_16104);
or U16627 (N_16627,N_16350,N_16045);
and U16628 (N_16628,N_16422,N_16024);
nor U16629 (N_16629,N_16223,N_16074);
or U16630 (N_16630,N_16417,N_16139);
or U16631 (N_16631,N_16080,N_16005);
or U16632 (N_16632,N_16030,N_16484);
nand U16633 (N_16633,N_16191,N_16493);
and U16634 (N_16634,N_16259,N_16076);
nor U16635 (N_16635,N_16472,N_16017);
or U16636 (N_16636,N_16014,N_16442);
nor U16637 (N_16637,N_16393,N_16226);
nor U16638 (N_16638,N_16079,N_16268);
nand U16639 (N_16639,N_16458,N_16286);
and U16640 (N_16640,N_16163,N_16124);
nand U16641 (N_16641,N_16317,N_16368);
or U16642 (N_16642,N_16344,N_16133);
and U16643 (N_16643,N_16333,N_16216);
nor U16644 (N_16644,N_16362,N_16156);
or U16645 (N_16645,N_16343,N_16078);
nand U16646 (N_16646,N_16299,N_16116);
or U16647 (N_16647,N_16200,N_16221);
or U16648 (N_16648,N_16495,N_16186);
and U16649 (N_16649,N_16168,N_16440);
nor U16650 (N_16650,N_16494,N_16233);
nand U16651 (N_16651,N_16122,N_16245);
nand U16652 (N_16652,N_16253,N_16199);
nor U16653 (N_16653,N_16179,N_16220);
nor U16654 (N_16654,N_16126,N_16373);
nor U16655 (N_16655,N_16461,N_16323);
or U16656 (N_16656,N_16463,N_16356);
nor U16657 (N_16657,N_16329,N_16166);
nor U16658 (N_16658,N_16261,N_16321);
and U16659 (N_16659,N_16308,N_16334);
nor U16660 (N_16660,N_16497,N_16039);
and U16661 (N_16661,N_16483,N_16318);
nand U16662 (N_16662,N_16457,N_16392);
or U16663 (N_16663,N_16310,N_16402);
and U16664 (N_16664,N_16083,N_16374);
or U16665 (N_16665,N_16372,N_16346);
nand U16666 (N_16666,N_16140,N_16434);
or U16667 (N_16667,N_16499,N_16389);
nor U16668 (N_16668,N_16297,N_16197);
nand U16669 (N_16669,N_16443,N_16353);
or U16670 (N_16670,N_16454,N_16094);
or U16671 (N_16671,N_16390,N_16396);
or U16672 (N_16672,N_16438,N_16130);
nand U16673 (N_16673,N_16137,N_16129);
or U16674 (N_16674,N_16217,N_16035);
or U16675 (N_16675,N_16118,N_16325);
nand U16676 (N_16676,N_16001,N_16427);
nand U16677 (N_16677,N_16476,N_16151);
or U16678 (N_16678,N_16025,N_16294);
nor U16679 (N_16679,N_16330,N_16339);
or U16680 (N_16680,N_16266,N_16051);
nor U16681 (N_16681,N_16108,N_16282);
nor U16682 (N_16682,N_16273,N_16203);
and U16683 (N_16683,N_16478,N_16460);
nor U16684 (N_16684,N_16475,N_16262);
nand U16685 (N_16685,N_16311,N_16477);
or U16686 (N_16686,N_16425,N_16243);
or U16687 (N_16687,N_16448,N_16084);
or U16688 (N_16688,N_16210,N_16178);
and U16689 (N_16689,N_16102,N_16410);
and U16690 (N_16690,N_16328,N_16224);
and U16691 (N_16691,N_16195,N_16181);
nand U16692 (N_16692,N_16403,N_16414);
nor U16693 (N_16693,N_16399,N_16269);
nor U16694 (N_16694,N_16093,N_16265);
nor U16695 (N_16695,N_16183,N_16358);
and U16696 (N_16696,N_16441,N_16413);
or U16697 (N_16697,N_16161,N_16301);
nand U16698 (N_16698,N_16314,N_16020);
nand U16699 (N_16699,N_16101,N_16304);
nor U16700 (N_16700,N_16098,N_16360);
and U16701 (N_16701,N_16190,N_16489);
and U16702 (N_16702,N_16150,N_16467);
nor U16703 (N_16703,N_16284,N_16154);
nand U16704 (N_16704,N_16411,N_16341);
nand U16705 (N_16705,N_16009,N_16336);
nand U16706 (N_16706,N_16347,N_16174);
nor U16707 (N_16707,N_16271,N_16155);
nor U16708 (N_16708,N_16177,N_16069);
and U16709 (N_16709,N_16112,N_16201);
nor U16710 (N_16710,N_16322,N_16319);
nor U16711 (N_16711,N_16293,N_16077);
and U16712 (N_16712,N_16230,N_16468);
nor U16713 (N_16713,N_16378,N_16007);
or U16714 (N_16714,N_16379,N_16466);
and U16715 (N_16715,N_16236,N_16409);
or U16716 (N_16716,N_16081,N_16142);
nor U16717 (N_16717,N_16072,N_16370);
or U16718 (N_16718,N_16401,N_16096);
nand U16719 (N_16719,N_16198,N_16385);
and U16720 (N_16720,N_16218,N_16002);
nor U16721 (N_16721,N_16225,N_16187);
or U16722 (N_16722,N_16109,N_16086);
or U16723 (N_16723,N_16256,N_16046);
or U16724 (N_16724,N_16146,N_16202);
and U16725 (N_16725,N_16430,N_16019);
nand U16726 (N_16726,N_16335,N_16487);
and U16727 (N_16727,N_16008,N_16332);
or U16728 (N_16728,N_16240,N_16121);
and U16729 (N_16729,N_16351,N_16394);
or U16730 (N_16730,N_16426,N_16075);
and U16731 (N_16731,N_16031,N_16290);
or U16732 (N_16732,N_16446,N_16175);
and U16733 (N_16733,N_16136,N_16141);
nor U16734 (N_16734,N_16062,N_16277);
nand U16735 (N_16735,N_16307,N_16249);
or U16736 (N_16736,N_16153,N_16433);
nor U16737 (N_16737,N_16380,N_16056);
and U16738 (N_16738,N_16312,N_16065);
or U16739 (N_16739,N_16398,N_16431);
nand U16740 (N_16740,N_16292,N_16263);
and U16741 (N_16741,N_16167,N_16429);
nor U16742 (N_16742,N_16196,N_16127);
and U16743 (N_16743,N_16320,N_16073);
nor U16744 (N_16744,N_16364,N_16280);
and U16745 (N_16745,N_16365,N_16113);
nor U16746 (N_16746,N_16490,N_16338);
nand U16747 (N_16747,N_16459,N_16436);
nand U16748 (N_16748,N_16185,N_16047);
and U16749 (N_16749,N_16100,N_16473);
nor U16750 (N_16750,N_16225,N_16123);
or U16751 (N_16751,N_16081,N_16000);
or U16752 (N_16752,N_16446,N_16198);
and U16753 (N_16753,N_16356,N_16325);
and U16754 (N_16754,N_16362,N_16321);
nor U16755 (N_16755,N_16074,N_16439);
nand U16756 (N_16756,N_16491,N_16208);
or U16757 (N_16757,N_16291,N_16213);
nor U16758 (N_16758,N_16346,N_16074);
nand U16759 (N_16759,N_16405,N_16196);
nand U16760 (N_16760,N_16451,N_16135);
nand U16761 (N_16761,N_16187,N_16362);
and U16762 (N_16762,N_16253,N_16006);
or U16763 (N_16763,N_16099,N_16395);
nand U16764 (N_16764,N_16380,N_16428);
and U16765 (N_16765,N_16276,N_16168);
and U16766 (N_16766,N_16433,N_16417);
nor U16767 (N_16767,N_16412,N_16396);
nor U16768 (N_16768,N_16110,N_16234);
or U16769 (N_16769,N_16335,N_16465);
nand U16770 (N_16770,N_16169,N_16425);
nor U16771 (N_16771,N_16040,N_16282);
and U16772 (N_16772,N_16054,N_16379);
nor U16773 (N_16773,N_16241,N_16044);
nand U16774 (N_16774,N_16103,N_16078);
xor U16775 (N_16775,N_16325,N_16146);
nand U16776 (N_16776,N_16157,N_16327);
nand U16777 (N_16777,N_16326,N_16440);
nand U16778 (N_16778,N_16423,N_16096);
nand U16779 (N_16779,N_16416,N_16427);
nor U16780 (N_16780,N_16351,N_16044);
nand U16781 (N_16781,N_16192,N_16385);
and U16782 (N_16782,N_16366,N_16305);
and U16783 (N_16783,N_16206,N_16202);
and U16784 (N_16784,N_16031,N_16194);
or U16785 (N_16785,N_16054,N_16331);
nor U16786 (N_16786,N_16314,N_16417);
nand U16787 (N_16787,N_16069,N_16281);
nor U16788 (N_16788,N_16313,N_16462);
or U16789 (N_16789,N_16365,N_16187);
and U16790 (N_16790,N_16190,N_16312);
nor U16791 (N_16791,N_16403,N_16052);
nand U16792 (N_16792,N_16233,N_16289);
or U16793 (N_16793,N_16199,N_16456);
nor U16794 (N_16794,N_16465,N_16078);
and U16795 (N_16795,N_16362,N_16488);
nand U16796 (N_16796,N_16306,N_16395);
and U16797 (N_16797,N_16279,N_16235);
and U16798 (N_16798,N_16235,N_16065);
or U16799 (N_16799,N_16346,N_16070);
or U16800 (N_16800,N_16396,N_16342);
and U16801 (N_16801,N_16473,N_16259);
nand U16802 (N_16802,N_16139,N_16324);
or U16803 (N_16803,N_16176,N_16249);
and U16804 (N_16804,N_16068,N_16132);
nand U16805 (N_16805,N_16394,N_16339);
nor U16806 (N_16806,N_16302,N_16400);
and U16807 (N_16807,N_16085,N_16259);
nor U16808 (N_16808,N_16402,N_16467);
and U16809 (N_16809,N_16083,N_16336);
nor U16810 (N_16810,N_16377,N_16240);
or U16811 (N_16811,N_16390,N_16468);
or U16812 (N_16812,N_16361,N_16309);
nor U16813 (N_16813,N_16325,N_16218);
nor U16814 (N_16814,N_16332,N_16050);
nand U16815 (N_16815,N_16043,N_16303);
nor U16816 (N_16816,N_16090,N_16135);
and U16817 (N_16817,N_16282,N_16372);
nor U16818 (N_16818,N_16252,N_16022);
nand U16819 (N_16819,N_16215,N_16380);
or U16820 (N_16820,N_16383,N_16388);
and U16821 (N_16821,N_16143,N_16325);
or U16822 (N_16822,N_16218,N_16322);
nor U16823 (N_16823,N_16256,N_16487);
and U16824 (N_16824,N_16249,N_16051);
nand U16825 (N_16825,N_16124,N_16476);
or U16826 (N_16826,N_16368,N_16121);
or U16827 (N_16827,N_16285,N_16009);
or U16828 (N_16828,N_16456,N_16403);
and U16829 (N_16829,N_16417,N_16152);
or U16830 (N_16830,N_16086,N_16105);
or U16831 (N_16831,N_16090,N_16468);
and U16832 (N_16832,N_16022,N_16406);
or U16833 (N_16833,N_16031,N_16069);
and U16834 (N_16834,N_16434,N_16475);
nand U16835 (N_16835,N_16409,N_16311);
nand U16836 (N_16836,N_16321,N_16457);
nor U16837 (N_16837,N_16381,N_16175);
and U16838 (N_16838,N_16248,N_16054);
nand U16839 (N_16839,N_16194,N_16392);
and U16840 (N_16840,N_16481,N_16025);
and U16841 (N_16841,N_16080,N_16237);
or U16842 (N_16842,N_16032,N_16254);
nor U16843 (N_16843,N_16211,N_16307);
or U16844 (N_16844,N_16349,N_16495);
or U16845 (N_16845,N_16158,N_16190);
or U16846 (N_16846,N_16224,N_16253);
and U16847 (N_16847,N_16156,N_16324);
and U16848 (N_16848,N_16048,N_16471);
and U16849 (N_16849,N_16286,N_16380);
and U16850 (N_16850,N_16349,N_16436);
and U16851 (N_16851,N_16499,N_16081);
nor U16852 (N_16852,N_16043,N_16402);
nand U16853 (N_16853,N_16331,N_16477);
nand U16854 (N_16854,N_16463,N_16227);
or U16855 (N_16855,N_16390,N_16184);
nand U16856 (N_16856,N_16413,N_16128);
nor U16857 (N_16857,N_16014,N_16269);
and U16858 (N_16858,N_16067,N_16371);
nand U16859 (N_16859,N_16056,N_16087);
or U16860 (N_16860,N_16117,N_16176);
and U16861 (N_16861,N_16159,N_16425);
or U16862 (N_16862,N_16169,N_16162);
and U16863 (N_16863,N_16109,N_16464);
or U16864 (N_16864,N_16143,N_16034);
or U16865 (N_16865,N_16184,N_16075);
and U16866 (N_16866,N_16339,N_16069);
or U16867 (N_16867,N_16304,N_16129);
nor U16868 (N_16868,N_16444,N_16027);
nand U16869 (N_16869,N_16138,N_16159);
and U16870 (N_16870,N_16080,N_16470);
nor U16871 (N_16871,N_16047,N_16274);
and U16872 (N_16872,N_16057,N_16213);
and U16873 (N_16873,N_16486,N_16224);
nor U16874 (N_16874,N_16463,N_16428);
or U16875 (N_16875,N_16425,N_16094);
or U16876 (N_16876,N_16094,N_16293);
or U16877 (N_16877,N_16332,N_16154);
or U16878 (N_16878,N_16447,N_16011);
and U16879 (N_16879,N_16024,N_16043);
or U16880 (N_16880,N_16473,N_16127);
nor U16881 (N_16881,N_16130,N_16468);
nor U16882 (N_16882,N_16232,N_16012);
nor U16883 (N_16883,N_16101,N_16339);
nand U16884 (N_16884,N_16451,N_16301);
and U16885 (N_16885,N_16416,N_16003);
nand U16886 (N_16886,N_16081,N_16002);
nor U16887 (N_16887,N_16370,N_16457);
and U16888 (N_16888,N_16463,N_16003);
nor U16889 (N_16889,N_16035,N_16394);
and U16890 (N_16890,N_16346,N_16267);
and U16891 (N_16891,N_16385,N_16256);
or U16892 (N_16892,N_16099,N_16267);
and U16893 (N_16893,N_16246,N_16136);
nor U16894 (N_16894,N_16388,N_16101);
or U16895 (N_16895,N_16300,N_16409);
or U16896 (N_16896,N_16481,N_16130);
and U16897 (N_16897,N_16097,N_16321);
or U16898 (N_16898,N_16050,N_16480);
and U16899 (N_16899,N_16030,N_16064);
or U16900 (N_16900,N_16375,N_16014);
and U16901 (N_16901,N_16392,N_16131);
nor U16902 (N_16902,N_16291,N_16352);
and U16903 (N_16903,N_16152,N_16361);
nor U16904 (N_16904,N_16263,N_16348);
and U16905 (N_16905,N_16036,N_16269);
nor U16906 (N_16906,N_16487,N_16447);
nand U16907 (N_16907,N_16028,N_16143);
nand U16908 (N_16908,N_16240,N_16305);
or U16909 (N_16909,N_16438,N_16253);
nand U16910 (N_16910,N_16040,N_16387);
or U16911 (N_16911,N_16356,N_16368);
or U16912 (N_16912,N_16449,N_16478);
and U16913 (N_16913,N_16471,N_16133);
nor U16914 (N_16914,N_16288,N_16326);
and U16915 (N_16915,N_16189,N_16314);
nand U16916 (N_16916,N_16295,N_16140);
xnor U16917 (N_16917,N_16263,N_16036);
or U16918 (N_16918,N_16195,N_16333);
and U16919 (N_16919,N_16085,N_16064);
nand U16920 (N_16920,N_16066,N_16164);
nor U16921 (N_16921,N_16330,N_16001);
and U16922 (N_16922,N_16038,N_16077);
nor U16923 (N_16923,N_16296,N_16009);
nor U16924 (N_16924,N_16480,N_16202);
or U16925 (N_16925,N_16273,N_16149);
nor U16926 (N_16926,N_16480,N_16301);
nor U16927 (N_16927,N_16234,N_16137);
or U16928 (N_16928,N_16482,N_16384);
and U16929 (N_16929,N_16455,N_16029);
nor U16930 (N_16930,N_16277,N_16055);
nor U16931 (N_16931,N_16064,N_16367);
nand U16932 (N_16932,N_16088,N_16487);
nand U16933 (N_16933,N_16204,N_16238);
nor U16934 (N_16934,N_16446,N_16234);
nand U16935 (N_16935,N_16120,N_16432);
or U16936 (N_16936,N_16025,N_16028);
nor U16937 (N_16937,N_16215,N_16010);
or U16938 (N_16938,N_16328,N_16154);
nor U16939 (N_16939,N_16362,N_16224);
and U16940 (N_16940,N_16377,N_16141);
and U16941 (N_16941,N_16182,N_16064);
and U16942 (N_16942,N_16279,N_16332);
or U16943 (N_16943,N_16466,N_16400);
and U16944 (N_16944,N_16197,N_16391);
nand U16945 (N_16945,N_16442,N_16491);
or U16946 (N_16946,N_16494,N_16441);
nand U16947 (N_16947,N_16028,N_16131);
or U16948 (N_16948,N_16408,N_16186);
nand U16949 (N_16949,N_16027,N_16151);
nor U16950 (N_16950,N_16143,N_16016);
and U16951 (N_16951,N_16123,N_16407);
nand U16952 (N_16952,N_16420,N_16182);
or U16953 (N_16953,N_16084,N_16479);
and U16954 (N_16954,N_16438,N_16045);
nand U16955 (N_16955,N_16446,N_16255);
nand U16956 (N_16956,N_16432,N_16191);
and U16957 (N_16957,N_16014,N_16467);
nand U16958 (N_16958,N_16390,N_16255);
or U16959 (N_16959,N_16095,N_16062);
and U16960 (N_16960,N_16024,N_16382);
and U16961 (N_16961,N_16393,N_16137);
and U16962 (N_16962,N_16315,N_16017);
nand U16963 (N_16963,N_16387,N_16275);
and U16964 (N_16964,N_16139,N_16314);
nand U16965 (N_16965,N_16464,N_16268);
or U16966 (N_16966,N_16478,N_16319);
nand U16967 (N_16967,N_16454,N_16284);
and U16968 (N_16968,N_16127,N_16320);
nand U16969 (N_16969,N_16182,N_16185);
nand U16970 (N_16970,N_16187,N_16451);
nor U16971 (N_16971,N_16387,N_16316);
or U16972 (N_16972,N_16154,N_16186);
nor U16973 (N_16973,N_16360,N_16420);
and U16974 (N_16974,N_16032,N_16143);
and U16975 (N_16975,N_16339,N_16238);
nand U16976 (N_16976,N_16425,N_16195);
and U16977 (N_16977,N_16087,N_16233);
nand U16978 (N_16978,N_16092,N_16303);
nand U16979 (N_16979,N_16478,N_16286);
nand U16980 (N_16980,N_16487,N_16117);
and U16981 (N_16981,N_16337,N_16291);
or U16982 (N_16982,N_16224,N_16462);
and U16983 (N_16983,N_16097,N_16431);
nand U16984 (N_16984,N_16297,N_16019);
or U16985 (N_16985,N_16328,N_16161);
nand U16986 (N_16986,N_16320,N_16231);
and U16987 (N_16987,N_16355,N_16233);
nand U16988 (N_16988,N_16297,N_16290);
nand U16989 (N_16989,N_16427,N_16033);
nor U16990 (N_16990,N_16406,N_16037);
nor U16991 (N_16991,N_16319,N_16008);
nor U16992 (N_16992,N_16127,N_16334);
nand U16993 (N_16993,N_16176,N_16140);
or U16994 (N_16994,N_16173,N_16459);
nor U16995 (N_16995,N_16002,N_16454);
xnor U16996 (N_16996,N_16292,N_16382);
and U16997 (N_16997,N_16436,N_16011);
nor U16998 (N_16998,N_16382,N_16492);
or U16999 (N_16999,N_16253,N_16014);
and U17000 (N_17000,N_16831,N_16616);
or U17001 (N_17001,N_16605,N_16766);
nor U17002 (N_17002,N_16537,N_16918);
and U17003 (N_17003,N_16562,N_16998);
and U17004 (N_17004,N_16870,N_16815);
or U17005 (N_17005,N_16536,N_16912);
nand U17006 (N_17006,N_16597,N_16796);
and U17007 (N_17007,N_16784,N_16734);
or U17008 (N_17008,N_16833,N_16798);
nand U17009 (N_17009,N_16924,N_16834);
xnor U17010 (N_17010,N_16602,N_16922);
nor U17011 (N_17011,N_16933,N_16812);
or U17012 (N_17012,N_16808,N_16787);
and U17013 (N_17013,N_16806,N_16719);
nor U17014 (N_17014,N_16532,N_16825);
and U17015 (N_17015,N_16905,N_16611);
and U17016 (N_17016,N_16504,N_16632);
nor U17017 (N_17017,N_16821,N_16722);
or U17018 (N_17018,N_16881,N_16883);
or U17019 (N_17019,N_16691,N_16711);
and U17020 (N_17020,N_16662,N_16548);
nor U17021 (N_17021,N_16989,N_16743);
or U17022 (N_17022,N_16984,N_16811);
or U17023 (N_17023,N_16684,N_16601);
nand U17024 (N_17024,N_16578,N_16680);
and U17025 (N_17025,N_16773,N_16910);
or U17026 (N_17026,N_16664,N_16506);
or U17027 (N_17027,N_16813,N_16539);
nand U17028 (N_17028,N_16976,N_16841);
nor U17029 (N_17029,N_16789,N_16909);
nor U17030 (N_17030,N_16647,N_16614);
nand U17031 (N_17031,N_16519,N_16767);
nor U17032 (N_17032,N_16728,N_16744);
nor U17033 (N_17033,N_16947,N_16669);
and U17034 (N_17034,N_16810,N_16846);
or U17035 (N_17035,N_16964,N_16979);
and U17036 (N_17036,N_16726,N_16627);
and U17037 (N_17037,N_16708,N_16926);
nor U17038 (N_17038,N_16606,N_16770);
or U17039 (N_17039,N_16509,N_16546);
nor U17040 (N_17040,N_16580,N_16668);
and U17041 (N_17041,N_16794,N_16588);
and U17042 (N_17042,N_16761,N_16688);
nor U17043 (N_17043,N_16823,N_16852);
nor U17044 (N_17044,N_16755,N_16582);
and U17045 (N_17045,N_16826,N_16667);
nand U17046 (N_17046,N_16530,N_16779);
nor U17047 (N_17047,N_16855,N_16550);
nand U17048 (N_17048,N_16762,N_16625);
and U17049 (N_17049,N_16746,N_16970);
nand U17050 (N_17050,N_16520,N_16544);
and U17051 (N_17051,N_16753,N_16774);
or U17052 (N_17052,N_16931,N_16879);
and U17053 (N_17053,N_16959,N_16518);
xor U17054 (N_17054,N_16771,N_16685);
nand U17055 (N_17055,N_16945,N_16942);
nand U17056 (N_17056,N_16786,N_16748);
nor U17057 (N_17057,N_16820,N_16844);
nand U17058 (N_17058,N_16732,N_16636);
nor U17059 (N_17059,N_16783,N_16639);
and U17060 (N_17060,N_16987,N_16995);
nand U17061 (N_17061,N_16673,N_16567);
nor U17062 (N_17062,N_16514,N_16788);
nand U17063 (N_17063,N_16862,N_16952);
nand U17064 (N_17064,N_16791,N_16701);
or U17065 (N_17065,N_16955,N_16749);
xor U17066 (N_17066,N_16529,N_16835);
or U17067 (N_17067,N_16534,N_16581);
or U17068 (N_17068,N_16861,N_16928);
nand U17069 (N_17069,N_16859,N_16988);
nor U17070 (N_17070,N_16756,N_16697);
and U17071 (N_17071,N_16535,N_16738);
nor U17072 (N_17072,N_16510,N_16501);
or U17073 (N_17073,N_16948,N_16682);
and U17074 (N_17074,N_16968,N_16842);
or U17075 (N_17075,N_16759,N_16515);
nand U17076 (N_17076,N_16686,N_16698);
nand U17077 (N_17077,N_16814,N_16887);
nand U17078 (N_17078,N_16804,N_16653);
nor U17079 (N_17079,N_16954,N_16594);
nor U17080 (N_17080,N_16752,N_16982);
or U17081 (N_17081,N_16573,N_16713);
nor U17082 (N_17082,N_16974,N_16953);
nor U17083 (N_17083,N_16729,N_16571);
nand U17084 (N_17084,N_16706,N_16750);
and U17085 (N_17085,N_16619,N_16860);
nand U17086 (N_17086,N_16792,N_16890);
and U17087 (N_17087,N_16717,N_16699);
nand U17088 (N_17088,N_16652,N_16695);
or U17089 (N_17089,N_16715,N_16962);
nand U17090 (N_17090,N_16683,N_16888);
or U17091 (N_17091,N_16591,N_16503);
or U17092 (N_17092,N_16949,N_16838);
nor U17093 (N_17093,N_16649,N_16656);
or U17094 (N_17094,N_16843,N_16896);
and U17095 (N_17095,N_16915,N_16644);
nand U17096 (N_17096,N_16527,N_16533);
nand U17097 (N_17097,N_16508,N_16595);
and U17098 (N_17098,N_16568,N_16930);
and U17099 (N_17099,N_16563,N_16723);
and U17100 (N_17100,N_16650,N_16675);
nor U17101 (N_17101,N_16985,N_16872);
nor U17102 (N_17102,N_16589,N_16694);
and U17103 (N_17103,N_16936,N_16598);
and U17104 (N_17104,N_16999,N_16892);
nor U17105 (N_17105,N_16950,N_16642);
nand U17106 (N_17106,N_16781,N_16907);
nor U17107 (N_17107,N_16857,N_16782);
nor U17108 (N_17108,N_16523,N_16564);
nor U17109 (N_17109,N_16615,N_16799);
nand U17110 (N_17110,N_16666,N_16921);
nand U17111 (N_17111,N_16747,N_16967);
and U17112 (N_17112,N_16972,N_16618);
nor U17113 (N_17113,N_16513,N_16724);
nand U17114 (N_17114,N_16898,N_16874);
nand U17115 (N_17115,N_16986,N_16900);
or U17116 (N_17116,N_16853,N_16628);
or U17117 (N_17117,N_16856,N_16911);
and U17118 (N_17118,N_16737,N_16960);
or U17119 (N_17119,N_16740,N_16889);
or U17120 (N_17120,N_16885,N_16512);
and U17121 (N_17121,N_16891,N_16958);
or U17122 (N_17122,N_16661,N_16660);
nand U17123 (N_17123,N_16772,N_16617);
and U17124 (N_17124,N_16648,N_16696);
or U17125 (N_17125,N_16569,N_16693);
nand U17126 (N_17126,N_16754,N_16903);
nor U17127 (N_17127,N_16863,N_16816);
or U17128 (N_17128,N_16961,N_16946);
or U17129 (N_17129,N_16624,N_16765);
xnor U17130 (N_17130,N_16864,N_16681);
nor U17131 (N_17131,N_16689,N_16603);
nand U17132 (N_17132,N_16542,N_16929);
nand U17133 (N_17133,N_16975,N_16585);
nor U17134 (N_17134,N_16604,N_16925);
or U17135 (N_17135,N_16637,N_16654);
nand U17136 (N_17136,N_16600,N_16620);
or U17137 (N_17137,N_16866,N_16801);
or U17138 (N_17138,N_16832,N_16956);
nor U17139 (N_17139,N_16865,N_16780);
and U17140 (N_17140,N_16941,N_16741);
nor U17141 (N_17141,N_16525,N_16797);
or U17142 (N_17142,N_16549,N_16596);
and U17143 (N_17143,N_16802,N_16626);
and U17144 (N_17144,N_16575,N_16908);
and U17145 (N_17145,N_16555,N_16709);
or U17146 (N_17146,N_16920,N_16793);
nor U17147 (N_17147,N_16579,N_16839);
or U17148 (N_17148,N_16655,N_16822);
and U17149 (N_17149,N_16692,N_16731);
nand U17150 (N_17150,N_16511,N_16854);
and U17151 (N_17151,N_16940,N_16521);
and U17152 (N_17152,N_16971,N_16769);
nand U17153 (N_17153,N_16730,N_16676);
nand U17154 (N_17154,N_16674,N_16851);
nor U17155 (N_17155,N_16720,N_16570);
or U17156 (N_17156,N_16612,N_16672);
nor U17157 (N_17157,N_16540,N_16916);
nor U17158 (N_17158,N_16980,N_16845);
or U17159 (N_17159,N_16621,N_16994);
nand U17160 (N_17160,N_16522,N_16914);
nor U17161 (N_17161,N_16704,N_16847);
nor U17162 (N_17162,N_16871,N_16561);
and U17163 (N_17163,N_16643,N_16560);
or U17164 (N_17164,N_16608,N_16776);
xnor U17165 (N_17165,N_16751,N_16705);
nor U17166 (N_17166,N_16700,N_16623);
and U17167 (N_17167,N_16663,N_16500);
nor U17168 (N_17168,N_16742,N_16934);
or U17169 (N_17169,N_16609,N_16923);
or U17170 (N_17170,N_16869,N_16807);
or U17171 (N_17171,N_16651,N_16867);
nand U17172 (N_17172,N_16785,N_16505);
and U17173 (N_17173,N_16757,N_16725);
nor U17174 (N_17174,N_16893,N_16758);
nor U17175 (N_17175,N_16897,N_16531);
and U17176 (N_17176,N_16678,N_16538);
nor U17177 (N_17177,N_16895,N_16583);
or U17178 (N_17178,N_16547,N_16592);
nand U17179 (N_17179,N_16877,N_16703);
and U17180 (N_17180,N_16763,N_16634);
and U17181 (N_17181,N_16640,N_16690);
and U17182 (N_17182,N_16828,N_16795);
nor U17183 (N_17183,N_16516,N_16957);
or U17184 (N_17184,N_16996,N_16944);
nand U17185 (N_17185,N_16727,N_16904);
nor U17186 (N_17186,N_16677,N_16610);
nand U17187 (N_17187,N_16901,N_16665);
and U17188 (N_17188,N_16679,N_16553);
or U17189 (N_17189,N_16764,N_16556);
nor U17190 (N_17190,N_16809,N_16817);
or U17191 (N_17191,N_16951,N_16659);
nand U17192 (N_17192,N_16902,N_16524);
nand U17193 (N_17193,N_16899,N_16827);
nand U17194 (N_17194,N_16830,N_16848);
or U17195 (N_17195,N_16932,N_16966);
and U17196 (N_17196,N_16590,N_16635);
and U17197 (N_17197,N_16850,N_16587);
nand U17198 (N_17198,N_16574,N_16716);
nor U17199 (N_17199,N_16710,N_16990);
or U17200 (N_17200,N_16671,N_16702);
or U17201 (N_17201,N_16735,N_16938);
and U17202 (N_17202,N_16577,N_16778);
and U17203 (N_17203,N_16917,N_16775);
nor U17204 (N_17204,N_16552,N_16593);
and U17205 (N_17205,N_16840,N_16631);
nand U17206 (N_17206,N_16836,N_16565);
or U17207 (N_17207,N_16507,N_16992);
nor U17208 (N_17208,N_16645,N_16829);
nor U17209 (N_17209,N_16559,N_16768);
nand U17210 (N_17210,N_16991,N_16965);
nor U17211 (N_17211,N_16819,N_16993);
nand U17212 (N_17212,N_16586,N_16943);
nor U17213 (N_17213,N_16894,N_16973);
nand U17214 (N_17214,N_16805,N_16541);
or U17215 (N_17215,N_16880,N_16572);
or U17216 (N_17216,N_16760,N_16712);
and U17217 (N_17217,N_16576,N_16670);
nand U17218 (N_17218,N_16613,N_16977);
or U17219 (N_17219,N_16927,N_16849);
nand U17220 (N_17220,N_16543,N_16997);
nor U17221 (N_17221,N_16824,N_16937);
nand U17222 (N_17222,N_16502,N_16718);
or U17223 (N_17223,N_16707,N_16633);
and U17224 (N_17224,N_16558,N_16557);
or U17225 (N_17225,N_16599,N_16528);
nor U17226 (N_17226,N_16721,N_16584);
and U17227 (N_17227,N_16886,N_16906);
and U17228 (N_17228,N_16882,N_16875);
nand U17229 (N_17229,N_16545,N_16733);
nor U17230 (N_17230,N_16745,N_16876);
and U17231 (N_17231,N_16641,N_16630);
and U17232 (N_17232,N_16658,N_16983);
nand U17233 (N_17233,N_16963,N_16714);
nor U17234 (N_17234,N_16935,N_16884);
nand U17235 (N_17235,N_16969,N_16687);
nand U17236 (N_17236,N_16554,N_16873);
nand U17237 (N_17237,N_16790,N_16526);
nand U17238 (N_17238,N_16803,N_16739);
nor U17239 (N_17239,N_16629,N_16736);
and U17240 (N_17240,N_16981,N_16978);
nor U17241 (N_17241,N_16913,N_16607);
nand U17242 (N_17242,N_16777,N_16800);
nor U17243 (N_17243,N_16939,N_16657);
or U17244 (N_17244,N_16878,N_16551);
nor U17245 (N_17245,N_16517,N_16818);
and U17246 (N_17246,N_16858,N_16868);
or U17247 (N_17247,N_16837,N_16638);
or U17248 (N_17248,N_16566,N_16646);
xor U17249 (N_17249,N_16919,N_16622);
and U17250 (N_17250,N_16823,N_16848);
or U17251 (N_17251,N_16551,N_16684);
nand U17252 (N_17252,N_16805,N_16835);
and U17253 (N_17253,N_16980,N_16929);
or U17254 (N_17254,N_16615,N_16998);
xor U17255 (N_17255,N_16541,N_16791);
nand U17256 (N_17256,N_16611,N_16915);
nand U17257 (N_17257,N_16789,N_16517);
nor U17258 (N_17258,N_16699,N_16778);
nor U17259 (N_17259,N_16901,N_16706);
and U17260 (N_17260,N_16528,N_16798);
nand U17261 (N_17261,N_16904,N_16991);
nor U17262 (N_17262,N_16726,N_16821);
nand U17263 (N_17263,N_16995,N_16740);
or U17264 (N_17264,N_16916,N_16532);
nand U17265 (N_17265,N_16708,N_16745);
and U17266 (N_17266,N_16555,N_16638);
nor U17267 (N_17267,N_16810,N_16614);
nor U17268 (N_17268,N_16731,N_16567);
and U17269 (N_17269,N_16752,N_16928);
and U17270 (N_17270,N_16542,N_16532);
nor U17271 (N_17271,N_16760,N_16731);
xor U17272 (N_17272,N_16928,N_16973);
or U17273 (N_17273,N_16753,N_16989);
nand U17274 (N_17274,N_16672,N_16658);
nand U17275 (N_17275,N_16796,N_16797);
nor U17276 (N_17276,N_16545,N_16722);
nor U17277 (N_17277,N_16975,N_16796);
nand U17278 (N_17278,N_16791,N_16972);
nand U17279 (N_17279,N_16668,N_16977);
nor U17280 (N_17280,N_16746,N_16960);
and U17281 (N_17281,N_16512,N_16945);
and U17282 (N_17282,N_16502,N_16643);
nor U17283 (N_17283,N_16527,N_16531);
nor U17284 (N_17284,N_16792,N_16929);
or U17285 (N_17285,N_16806,N_16760);
and U17286 (N_17286,N_16862,N_16566);
nor U17287 (N_17287,N_16799,N_16678);
or U17288 (N_17288,N_16685,N_16687);
and U17289 (N_17289,N_16761,N_16867);
or U17290 (N_17290,N_16799,N_16995);
or U17291 (N_17291,N_16899,N_16806);
or U17292 (N_17292,N_16807,N_16779);
nand U17293 (N_17293,N_16653,N_16989);
nand U17294 (N_17294,N_16586,N_16572);
nor U17295 (N_17295,N_16777,N_16751);
nor U17296 (N_17296,N_16512,N_16903);
or U17297 (N_17297,N_16784,N_16674);
nor U17298 (N_17298,N_16614,N_16611);
or U17299 (N_17299,N_16840,N_16993);
nand U17300 (N_17300,N_16715,N_16631);
xor U17301 (N_17301,N_16636,N_16713);
nand U17302 (N_17302,N_16697,N_16690);
or U17303 (N_17303,N_16600,N_16702);
and U17304 (N_17304,N_16910,N_16520);
nand U17305 (N_17305,N_16607,N_16873);
nor U17306 (N_17306,N_16968,N_16565);
xor U17307 (N_17307,N_16534,N_16526);
and U17308 (N_17308,N_16893,N_16760);
or U17309 (N_17309,N_16759,N_16754);
or U17310 (N_17310,N_16932,N_16832);
and U17311 (N_17311,N_16921,N_16869);
or U17312 (N_17312,N_16877,N_16938);
and U17313 (N_17313,N_16599,N_16980);
or U17314 (N_17314,N_16518,N_16714);
or U17315 (N_17315,N_16731,N_16658);
nor U17316 (N_17316,N_16649,N_16569);
or U17317 (N_17317,N_16593,N_16798);
and U17318 (N_17318,N_16895,N_16618);
or U17319 (N_17319,N_16791,N_16829);
nand U17320 (N_17320,N_16636,N_16882);
and U17321 (N_17321,N_16575,N_16501);
xor U17322 (N_17322,N_16824,N_16882);
nand U17323 (N_17323,N_16747,N_16900);
nand U17324 (N_17324,N_16583,N_16731);
nor U17325 (N_17325,N_16668,N_16824);
and U17326 (N_17326,N_16874,N_16996);
and U17327 (N_17327,N_16664,N_16807);
or U17328 (N_17328,N_16911,N_16925);
nand U17329 (N_17329,N_16925,N_16959);
or U17330 (N_17330,N_16914,N_16802);
nand U17331 (N_17331,N_16853,N_16664);
nand U17332 (N_17332,N_16661,N_16966);
nor U17333 (N_17333,N_16735,N_16945);
or U17334 (N_17334,N_16747,N_16821);
and U17335 (N_17335,N_16647,N_16898);
nor U17336 (N_17336,N_16501,N_16869);
nor U17337 (N_17337,N_16543,N_16940);
nand U17338 (N_17338,N_16956,N_16841);
nand U17339 (N_17339,N_16675,N_16700);
and U17340 (N_17340,N_16834,N_16798);
or U17341 (N_17341,N_16886,N_16827);
nor U17342 (N_17342,N_16723,N_16599);
nor U17343 (N_17343,N_16872,N_16677);
nand U17344 (N_17344,N_16859,N_16770);
nand U17345 (N_17345,N_16770,N_16881);
nand U17346 (N_17346,N_16826,N_16687);
or U17347 (N_17347,N_16892,N_16825);
or U17348 (N_17348,N_16940,N_16846);
nand U17349 (N_17349,N_16788,N_16720);
nand U17350 (N_17350,N_16965,N_16790);
and U17351 (N_17351,N_16723,N_16877);
nand U17352 (N_17352,N_16574,N_16992);
and U17353 (N_17353,N_16930,N_16856);
nand U17354 (N_17354,N_16971,N_16838);
and U17355 (N_17355,N_16568,N_16524);
or U17356 (N_17356,N_16829,N_16674);
nand U17357 (N_17357,N_16511,N_16561);
and U17358 (N_17358,N_16866,N_16840);
or U17359 (N_17359,N_16535,N_16510);
and U17360 (N_17360,N_16827,N_16653);
nor U17361 (N_17361,N_16531,N_16536);
nand U17362 (N_17362,N_16704,N_16672);
or U17363 (N_17363,N_16969,N_16821);
nor U17364 (N_17364,N_16682,N_16710);
nand U17365 (N_17365,N_16874,N_16756);
nand U17366 (N_17366,N_16686,N_16965);
nor U17367 (N_17367,N_16866,N_16709);
nand U17368 (N_17368,N_16714,N_16997);
xor U17369 (N_17369,N_16629,N_16667);
nand U17370 (N_17370,N_16503,N_16856);
nor U17371 (N_17371,N_16833,N_16991);
and U17372 (N_17372,N_16817,N_16866);
nor U17373 (N_17373,N_16768,N_16829);
and U17374 (N_17374,N_16812,N_16738);
and U17375 (N_17375,N_16684,N_16821);
or U17376 (N_17376,N_16764,N_16838);
nand U17377 (N_17377,N_16718,N_16890);
or U17378 (N_17378,N_16687,N_16816);
nor U17379 (N_17379,N_16615,N_16865);
and U17380 (N_17380,N_16998,N_16522);
nor U17381 (N_17381,N_16518,N_16801);
nand U17382 (N_17382,N_16554,N_16881);
or U17383 (N_17383,N_16597,N_16771);
nor U17384 (N_17384,N_16647,N_16508);
or U17385 (N_17385,N_16676,N_16890);
or U17386 (N_17386,N_16570,N_16616);
nand U17387 (N_17387,N_16967,N_16852);
or U17388 (N_17388,N_16983,N_16850);
nor U17389 (N_17389,N_16591,N_16532);
nand U17390 (N_17390,N_16644,N_16917);
nor U17391 (N_17391,N_16861,N_16690);
nor U17392 (N_17392,N_16967,N_16504);
nand U17393 (N_17393,N_16894,N_16726);
or U17394 (N_17394,N_16706,N_16674);
and U17395 (N_17395,N_16821,N_16955);
nand U17396 (N_17396,N_16876,N_16781);
or U17397 (N_17397,N_16819,N_16791);
nand U17398 (N_17398,N_16937,N_16897);
or U17399 (N_17399,N_16696,N_16637);
nor U17400 (N_17400,N_16606,N_16789);
nor U17401 (N_17401,N_16635,N_16724);
nand U17402 (N_17402,N_16962,N_16823);
and U17403 (N_17403,N_16817,N_16752);
and U17404 (N_17404,N_16956,N_16668);
nand U17405 (N_17405,N_16522,N_16911);
or U17406 (N_17406,N_16940,N_16547);
and U17407 (N_17407,N_16795,N_16733);
nor U17408 (N_17408,N_16617,N_16719);
or U17409 (N_17409,N_16990,N_16590);
and U17410 (N_17410,N_16616,N_16776);
xor U17411 (N_17411,N_16951,N_16842);
or U17412 (N_17412,N_16946,N_16599);
nand U17413 (N_17413,N_16729,N_16916);
nor U17414 (N_17414,N_16939,N_16923);
nand U17415 (N_17415,N_16872,N_16737);
or U17416 (N_17416,N_16979,N_16683);
nor U17417 (N_17417,N_16631,N_16819);
or U17418 (N_17418,N_16645,N_16983);
nor U17419 (N_17419,N_16749,N_16992);
or U17420 (N_17420,N_16763,N_16731);
or U17421 (N_17421,N_16881,N_16989);
or U17422 (N_17422,N_16840,N_16642);
nor U17423 (N_17423,N_16982,N_16714);
nor U17424 (N_17424,N_16983,N_16972);
nor U17425 (N_17425,N_16580,N_16952);
nor U17426 (N_17426,N_16742,N_16708);
and U17427 (N_17427,N_16667,N_16963);
nand U17428 (N_17428,N_16816,N_16726);
and U17429 (N_17429,N_16737,N_16707);
nand U17430 (N_17430,N_16612,N_16832);
nor U17431 (N_17431,N_16536,N_16870);
or U17432 (N_17432,N_16601,N_16729);
nand U17433 (N_17433,N_16588,N_16883);
or U17434 (N_17434,N_16618,N_16693);
or U17435 (N_17435,N_16905,N_16842);
nor U17436 (N_17436,N_16975,N_16812);
or U17437 (N_17437,N_16687,N_16860);
nor U17438 (N_17438,N_16896,N_16534);
and U17439 (N_17439,N_16769,N_16887);
nand U17440 (N_17440,N_16755,N_16837);
nor U17441 (N_17441,N_16797,N_16698);
nor U17442 (N_17442,N_16843,N_16519);
and U17443 (N_17443,N_16780,N_16546);
nand U17444 (N_17444,N_16539,N_16952);
and U17445 (N_17445,N_16774,N_16670);
or U17446 (N_17446,N_16641,N_16894);
nor U17447 (N_17447,N_16900,N_16515);
nand U17448 (N_17448,N_16661,N_16569);
and U17449 (N_17449,N_16550,N_16729);
nor U17450 (N_17450,N_16696,N_16543);
and U17451 (N_17451,N_16888,N_16719);
or U17452 (N_17452,N_16923,N_16924);
nand U17453 (N_17453,N_16681,N_16537);
or U17454 (N_17454,N_16778,N_16980);
or U17455 (N_17455,N_16696,N_16763);
nor U17456 (N_17456,N_16530,N_16583);
nor U17457 (N_17457,N_16980,N_16768);
nand U17458 (N_17458,N_16503,N_16595);
and U17459 (N_17459,N_16587,N_16932);
and U17460 (N_17460,N_16739,N_16877);
nand U17461 (N_17461,N_16744,N_16726);
nand U17462 (N_17462,N_16561,N_16772);
nor U17463 (N_17463,N_16529,N_16735);
nand U17464 (N_17464,N_16628,N_16943);
and U17465 (N_17465,N_16557,N_16688);
or U17466 (N_17466,N_16750,N_16664);
and U17467 (N_17467,N_16634,N_16576);
and U17468 (N_17468,N_16706,N_16513);
nand U17469 (N_17469,N_16986,N_16613);
and U17470 (N_17470,N_16901,N_16677);
nor U17471 (N_17471,N_16684,N_16798);
or U17472 (N_17472,N_16991,N_16681);
and U17473 (N_17473,N_16807,N_16847);
xor U17474 (N_17474,N_16834,N_16502);
or U17475 (N_17475,N_16900,N_16525);
nor U17476 (N_17476,N_16860,N_16772);
or U17477 (N_17477,N_16719,N_16543);
nand U17478 (N_17478,N_16602,N_16939);
or U17479 (N_17479,N_16969,N_16933);
nand U17480 (N_17480,N_16595,N_16637);
nor U17481 (N_17481,N_16755,N_16826);
nor U17482 (N_17482,N_16701,N_16556);
and U17483 (N_17483,N_16612,N_16896);
nor U17484 (N_17484,N_16744,N_16851);
xnor U17485 (N_17485,N_16910,N_16803);
and U17486 (N_17486,N_16858,N_16864);
and U17487 (N_17487,N_16898,N_16847);
nand U17488 (N_17488,N_16648,N_16548);
or U17489 (N_17489,N_16903,N_16552);
and U17490 (N_17490,N_16841,N_16717);
or U17491 (N_17491,N_16771,N_16619);
and U17492 (N_17492,N_16601,N_16598);
nand U17493 (N_17493,N_16895,N_16517);
or U17494 (N_17494,N_16946,N_16989);
nand U17495 (N_17495,N_16970,N_16512);
and U17496 (N_17496,N_16717,N_16898);
and U17497 (N_17497,N_16627,N_16848);
and U17498 (N_17498,N_16636,N_16904);
and U17499 (N_17499,N_16708,N_16656);
nand U17500 (N_17500,N_17185,N_17325);
nand U17501 (N_17501,N_17103,N_17483);
and U17502 (N_17502,N_17497,N_17117);
and U17503 (N_17503,N_17213,N_17205);
and U17504 (N_17504,N_17466,N_17287);
and U17505 (N_17505,N_17461,N_17076);
and U17506 (N_17506,N_17209,N_17479);
nand U17507 (N_17507,N_17308,N_17442);
or U17508 (N_17508,N_17046,N_17129);
nor U17509 (N_17509,N_17477,N_17436);
nor U17510 (N_17510,N_17063,N_17239);
nor U17511 (N_17511,N_17266,N_17055);
nor U17512 (N_17512,N_17125,N_17407);
or U17513 (N_17513,N_17165,N_17354);
and U17514 (N_17514,N_17413,N_17023);
or U17515 (N_17515,N_17351,N_17384);
nor U17516 (N_17516,N_17334,N_17356);
nor U17517 (N_17517,N_17134,N_17358);
and U17518 (N_17518,N_17323,N_17018);
nand U17519 (N_17519,N_17460,N_17397);
nand U17520 (N_17520,N_17039,N_17405);
nor U17521 (N_17521,N_17141,N_17142);
nand U17522 (N_17522,N_17448,N_17431);
nand U17523 (N_17523,N_17049,N_17084);
nand U17524 (N_17524,N_17488,N_17077);
or U17525 (N_17525,N_17464,N_17315);
and U17526 (N_17526,N_17302,N_17416);
nand U17527 (N_17527,N_17310,N_17007);
and U17528 (N_17528,N_17143,N_17008);
nor U17529 (N_17529,N_17314,N_17476);
or U17530 (N_17530,N_17158,N_17155);
nor U17531 (N_17531,N_17493,N_17194);
or U17532 (N_17532,N_17475,N_17439);
and U17533 (N_17533,N_17273,N_17121);
nand U17534 (N_17534,N_17449,N_17391);
nor U17535 (N_17535,N_17489,N_17432);
nand U17536 (N_17536,N_17361,N_17051);
and U17537 (N_17537,N_17062,N_17054);
nor U17538 (N_17538,N_17083,N_17374);
nand U17539 (N_17539,N_17094,N_17238);
nor U17540 (N_17540,N_17269,N_17126);
or U17541 (N_17541,N_17138,N_17446);
nor U17542 (N_17542,N_17202,N_17015);
or U17543 (N_17543,N_17048,N_17263);
nor U17544 (N_17544,N_17422,N_17309);
and U17545 (N_17545,N_17324,N_17376);
nor U17546 (N_17546,N_17003,N_17016);
nor U17547 (N_17547,N_17415,N_17445);
or U17548 (N_17548,N_17144,N_17111);
nor U17549 (N_17549,N_17183,N_17187);
nand U17550 (N_17550,N_17276,N_17246);
xor U17551 (N_17551,N_17344,N_17215);
nand U17552 (N_17552,N_17167,N_17406);
nor U17553 (N_17553,N_17359,N_17369);
nand U17554 (N_17554,N_17329,N_17332);
nand U17555 (N_17555,N_17119,N_17226);
or U17556 (N_17556,N_17420,N_17047);
nor U17557 (N_17557,N_17212,N_17345);
nor U17558 (N_17558,N_17087,N_17463);
and U17559 (N_17559,N_17154,N_17395);
and U17560 (N_17560,N_17275,N_17319);
nor U17561 (N_17561,N_17118,N_17434);
nor U17562 (N_17562,N_17452,N_17321);
and U17563 (N_17563,N_17322,N_17453);
nand U17564 (N_17564,N_17081,N_17066);
nor U17565 (N_17565,N_17184,N_17232);
nand U17566 (N_17566,N_17495,N_17256);
nand U17567 (N_17567,N_17365,N_17113);
and U17568 (N_17568,N_17400,N_17485);
and U17569 (N_17569,N_17043,N_17467);
nor U17570 (N_17570,N_17147,N_17450);
nand U17571 (N_17571,N_17274,N_17340);
nor U17572 (N_17572,N_17031,N_17417);
nand U17573 (N_17573,N_17280,N_17120);
and U17574 (N_17574,N_17005,N_17285);
and U17575 (N_17575,N_17425,N_17496);
nand U17576 (N_17576,N_17193,N_17474);
and U17577 (N_17577,N_17326,N_17462);
and U17578 (N_17578,N_17042,N_17045);
or U17579 (N_17579,N_17234,N_17257);
nand U17580 (N_17580,N_17377,N_17207);
and U17581 (N_17581,N_17132,N_17093);
or U17582 (N_17582,N_17097,N_17441);
or U17583 (N_17583,N_17056,N_17244);
nand U17584 (N_17584,N_17494,N_17074);
and U17585 (N_17585,N_17350,N_17170);
nand U17586 (N_17586,N_17072,N_17363);
and U17587 (N_17587,N_17228,N_17089);
nor U17588 (N_17588,N_17253,N_17243);
nand U17589 (N_17589,N_17382,N_17404);
nor U17590 (N_17590,N_17164,N_17311);
or U17591 (N_17591,N_17133,N_17331);
or U17592 (N_17592,N_17386,N_17010);
or U17593 (N_17593,N_17242,N_17271);
nor U17594 (N_17594,N_17053,N_17470);
and U17595 (N_17595,N_17109,N_17487);
nand U17596 (N_17596,N_17073,N_17293);
or U17597 (N_17597,N_17435,N_17333);
and U17598 (N_17598,N_17036,N_17301);
nor U17599 (N_17599,N_17195,N_17027);
or U17600 (N_17600,N_17469,N_17028);
nand U17601 (N_17601,N_17029,N_17300);
nor U17602 (N_17602,N_17380,N_17021);
nand U17603 (N_17603,N_17179,N_17443);
nand U17604 (N_17604,N_17190,N_17498);
nor U17605 (N_17605,N_17423,N_17139);
or U17606 (N_17606,N_17346,N_17251);
and U17607 (N_17607,N_17000,N_17379);
or U17608 (N_17608,N_17116,N_17353);
nor U17609 (N_17609,N_17229,N_17440);
nand U17610 (N_17610,N_17100,N_17286);
and U17611 (N_17611,N_17090,N_17317);
nor U17612 (N_17612,N_17233,N_17260);
or U17613 (N_17613,N_17349,N_17188);
nand U17614 (N_17614,N_17172,N_17067);
and U17615 (N_17615,N_17108,N_17421);
xor U17616 (N_17616,N_17288,N_17282);
and U17617 (N_17617,N_17065,N_17294);
nor U17618 (N_17618,N_17454,N_17082);
nand U17619 (N_17619,N_17347,N_17394);
nor U17620 (N_17620,N_17095,N_17231);
nor U17621 (N_17621,N_17124,N_17298);
nor U17622 (N_17622,N_17012,N_17388);
nand U17623 (N_17623,N_17402,N_17366);
nor U17624 (N_17624,N_17069,N_17372);
nor U17625 (N_17625,N_17412,N_17290);
and U17626 (N_17626,N_17387,N_17424);
nor U17627 (N_17627,N_17303,N_17211);
nand U17628 (N_17628,N_17447,N_17284);
and U17629 (N_17629,N_17057,N_17305);
nor U17630 (N_17630,N_17457,N_17304);
nand U17631 (N_17631,N_17037,N_17360);
or U17632 (N_17632,N_17250,N_17151);
nor U17633 (N_17633,N_17272,N_17465);
and U17634 (N_17634,N_17486,N_17252);
nor U17635 (N_17635,N_17203,N_17035);
and U17636 (N_17636,N_17092,N_17313);
nor U17637 (N_17637,N_17427,N_17022);
or U17638 (N_17638,N_17390,N_17071);
and U17639 (N_17639,N_17289,N_17001);
nand U17640 (N_17640,N_17052,N_17225);
and U17641 (N_17641,N_17255,N_17471);
nor U17642 (N_17642,N_17058,N_17392);
and U17643 (N_17643,N_17107,N_17472);
xnor U17644 (N_17644,N_17398,N_17152);
and U17645 (N_17645,N_17337,N_17490);
and U17646 (N_17646,N_17364,N_17375);
or U17647 (N_17647,N_17403,N_17355);
or U17648 (N_17648,N_17096,N_17075);
nand U17649 (N_17649,N_17197,N_17399);
nor U17650 (N_17650,N_17385,N_17335);
nand U17651 (N_17651,N_17009,N_17123);
nor U17652 (N_17652,N_17070,N_17159);
and U17653 (N_17653,N_17383,N_17091);
and U17654 (N_17654,N_17102,N_17178);
nand U17655 (N_17655,N_17024,N_17378);
and U17656 (N_17656,N_17101,N_17320);
nor U17657 (N_17657,N_17198,N_17222);
nor U17658 (N_17658,N_17214,N_17061);
nand U17659 (N_17659,N_17157,N_17088);
and U17660 (N_17660,N_17160,N_17006);
nand U17661 (N_17661,N_17339,N_17235);
or U17662 (N_17662,N_17254,N_17401);
or U17663 (N_17663,N_17227,N_17484);
or U17664 (N_17664,N_17341,N_17112);
nand U17665 (N_17665,N_17122,N_17156);
nand U17666 (N_17666,N_17307,N_17491);
nand U17667 (N_17667,N_17336,N_17020);
or U17668 (N_17668,N_17451,N_17371);
and U17669 (N_17669,N_17110,N_17411);
nand U17670 (N_17670,N_17292,N_17085);
nor U17671 (N_17671,N_17261,N_17150);
nand U17672 (N_17672,N_17223,N_17419);
nand U17673 (N_17673,N_17174,N_17078);
nor U17674 (N_17674,N_17196,N_17163);
or U17675 (N_17675,N_17131,N_17245);
and U17676 (N_17676,N_17492,N_17459);
or U17677 (N_17677,N_17279,N_17166);
or U17678 (N_17678,N_17348,N_17408);
and U17679 (N_17679,N_17200,N_17145);
or U17680 (N_17680,N_17409,N_17136);
nand U17681 (N_17681,N_17241,N_17328);
or U17682 (N_17682,N_17025,N_17410);
or U17683 (N_17683,N_17299,N_17019);
nand U17684 (N_17684,N_17418,N_17258);
nand U17685 (N_17685,N_17240,N_17060);
nor U17686 (N_17686,N_17201,N_17044);
nor U17687 (N_17687,N_17249,N_17175);
and U17688 (N_17688,N_17034,N_17478);
nor U17689 (N_17689,N_17277,N_17268);
nor U17690 (N_17690,N_17237,N_17080);
nand U17691 (N_17691,N_17014,N_17219);
xor U17692 (N_17692,N_17306,N_17499);
and U17693 (N_17693,N_17396,N_17393);
or U17694 (N_17694,N_17181,N_17148);
or U17695 (N_17695,N_17230,N_17149);
nand U17696 (N_17696,N_17079,N_17040);
nand U17697 (N_17697,N_17456,N_17017);
and U17698 (N_17698,N_17373,N_17468);
and U17699 (N_17699,N_17428,N_17481);
nor U17700 (N_17700,N_17480,N_17291);
or U17701 (N_17701,N_17059,N_17173);
nor U17702 (N_17702,N_17473,N_17186);
nor U17703 (N_17703,N_17199,N_17357);
and U17704 (N_17704,N_17104,N_17270);
and U17705 (N_17705,N_17265,N_17105);
and U17706 (N_17706,N_17161,N_17429);
and U17707 (N_17707,N_17011,N_17327);
nor U17708 (N_17708,N_17296,N_17318);
or U17709 (N_17709,N_17437,N_17208);
nor U17710 (N_17710,N_17026,N_17262);
nor U17711 (N_17711,N_17177,N_17221);
or U17712 (N_17712,N_17004,N_17278);
and U17713 (N_17713,N_17264,N_17224);
nor U17714 (N_17714,N_17192,N_17033);
or U17715 (N_17715,N_17482,N_17086);
nand U17716 (N_17716,N_17128,N_17247);
and U17717 (N_17717,N_17135,N_17362);
and U17718 (N_17718,N_17352,N_17316);
or U17719 (N_17719,N_17218,N_17153);
and U17720 (N_17720,N_17338,N_17312);
or U17721 (N_17721,N_17030,N_17259);
and U17722 (N_17722,N_17210,N_17146);
nand U17723 (N_17723,N_17444,N_17098);
nor U17724 (N_17724,N_17204,N_17099);
nor U17725 (N_17725,N_17169,N_17041);
nor U17726 (N_17726,N_17168,N_17106);
or U17727 (N_17727,N_17220,N_17381);
or U17728 (N_17728,N_17180,N_17032);
and U17729 (N_17729,N_17433,N_17114);
nand U17730 (N_17730,N_17367,N_17176);
nor U17731 (N_17731,N_17171,N_17430);
or U17732 (N_17732,N_17013,N_17248);
nor U17733 (N_17733,N_17370,N_17162);
nand U17734 (N_17734,N_17455,N_17127);
nor U17735 (N_17735,N_17206,N_17368);
and U17736 (N_17736,N_17182,N_17330);
and U17737 (N_17737,N_17236,N_17050);
or U17738 (N_17738,N_17267,N_17038);
or U17739 (N_17739,N_17343,N_17115);
nor U17740 (N_17740,N_17068,N_17216);
nand U17741 (N_17741,N_17458,N_17137);
nand U17742 (N_17742,N_17281,N_17283);
nor U17743 (N_17743,N_17217,N_17438);
nand U17744 (N_17744,N_17189,N_17130);
nor U17745 (N_17745,N_17191,N_17414);
or U17746 (N_17746,N_17064,N_17426);
nand U17747 (N_17747,N_17295,N_17342);
and U17748 (N_17748,N_17297,N_17002);
nand U17749 (N_17749,N_17389,N_17140);
nand U17750 (N_17750,N_17287,N_17066);
or U17751 (N_17751,N_17425,N_17011);
or U17752 (N_17752,N_17195,N_17462);
nor U17753 (N_17753,N_17012,N_17218);
and U17754 (N_17754,N_17456,N_17450);
nor U17755 (N_17755,N_17360,N_17326);
nand U17756 (N_17756,N_17259,N_17396);
and U17757 (N_17757,N_17198,N_17246);
nor U17758 (N_17758,N_17274,N_17334);
or U17759 (N_17759,N_17373,N_17268);
nor U17760 (N_17760,N_17037,N_17222);
or U17761 (N_17761,N_17358,N_17015);
nor U17762 (N_17762,N_17375,N_17085);
and U17763 (N_17763,N_17174,N_17310);
or U17764 (N_17764,N_17093,N_17431);
nor U17765 (N_17765,N_17090,N_17292);
and U17766 (N_17766,N_17228,N_17403);
nand U17767 (N_17767,N_17047,N_17499);
nor U17768 (N_17768,N_17075,N_17231);
and U17769 (N_17769,N_17089,N_17265);
nand U17770 (N_17770,N_17009,N_17030);
nor U17771 (N_17771,N_17175,N_17104);
or U17772 (N_17772,N_17152,N_17180);
nor U17773 (N_17773,N_17131,N_17046);
nor U17774 (N_17774,N_17338,N_17204);
nor U17775 (N_17775,N_17375,N_17293);
and U17776 (N_17776,N_17164,N_17107);
or U17777 (N_17777,N_17004,N_17177);
and U17778 (N_17778,N_17050,N_17068);
or U17779 (N_17779,N_17091,N_17325);
nor U17780 (N_17780,N_17061,N_17113);
and U17781 (N_17781,N_17307,N_17261);
nor U17782 (N_17782,N_17252,N_17226);
and U17783 (N_17783,N_17246,N_17188);
and U17784 (N_17784,N_17217,N_17180);
or U17785 (N_17785,N_17349,N_17420);
nor U17786 (N_17786,N_17143,N_17439);
or U17787 (N_17787,N_17135,N_17368);
or U17788 (N_17788,N_17269,N_17478);
and U17789 (N_17789,N_17057,N_17005);
and U17790 (N_17790,N_17229,N_17228);
nand U17791 (N_17791,N_17232,N_17400);
nor U17792 (N_17792,N_17272,N_17055);
nand U17793 (N_17793,N_17254,N_17351);
or U17794 (N_17794,N_17027,N_17337);
nand U17795 (N_17795,N_17391,N_17113);
or U17796 (N_17796,N_17050,N_17194);
or U17797 (N_17797,N_17295,N_17486);
and U17798 (N_17798,N_17435,N_17285);
or U17799 (N_17799,N_17456,N_17287);
nand U17800 (N_17800,N_17475,N_17072);
nand U17801 (N_17801,N_17111,N_17240);
or U17802 (N_17802,N_17284,N_17005);
or U17803 (N_17803,N_17452,N_17099);
or U17804 (N_17804,N_17206,N_17403);
and U17805 (N_17805,N_17094,N_17160);
nor U17806 (N_17806,N_17037,N_17103);
nor U17807 (N_17807,N_17127,N_17140);
and U17808 (N_17808,N_17245,N_17235);
nand U17809 (N_17809,N_17236,N_17237);
or U17810 (N_17810,N_17091,N_17010);
nor U17811 (N_17811,N_17290,N_17206);
and U17812 (N_17812,N_17455,N_17414);
nor U17813 (N_17813,N_17399,N_17297);
or U17814 (N_17814,N_17071,N_17160);
nand U17815 (N_17815,N_17149,N_17163);
or U17816 (N_17816,N_17203,N_17355);
and U17817 (N_17817,N_17281,N_17324);
nand U17818 (N_17818,N_17440,N_17225);
or U17819 (N_17819,N_17352,N_17288);
nor U17820 (N_17820,N_17446,N_17332);
nor U17821 (N_17821,N_17226,N_17372);
and U17822 (N_17822,N_17495,N_17053);
or U17823 (N_17823,N_17323,N_17376);
nor U17824 (N_17824,N_17186,N_17483);
or U17825 (N_17825,N_17131,N_17346);
nor U17826 (N_17826,N_17411,N_17067);
and U17827 (N_17827,N_17211,N_17206);
nand U17828 (N_17828,N_17098,N_17269);
nand U17829 (N_17829,N_17290,N_17315);
nand U17830 (N_17830,N_17045,N_17167);
and U17831 (N_17831,N_17140,N_17411);
nor U17832 (N_17832,N_17265,N_17115);
nor U17833 (N_17833,N_17098,N_17231);
and U17834 (N_17834,N_17432,N_17098);
nor U17835 (N_17835,N_17192,N_17334);
nor U17836 (N_17836,N_17433,N_17478);
nand U17837 (N_17837,N_17327,N_17203);
nand U17838 (N_17838,N_17004,N_17324);
nand U17839 (N_17839,N_17425,N_17075);
and U17840 (N_17840,N_17361,N_17458);
nand U17841 (N_17841,N_17224,N_17380);
nand U17842 (N_17842,N_17142,N_17018);
nand U17843 (N_17843,N_17492,N_17239);
or U17844 (N_17844,N_17260,N_17084);
nor U17845 (N_17845,N_17041,N_17175);
nand U17846 (N_17846,N_17247,N_17108);
nand U17847 (N_17847,N_17249,N_17183);
or U17848 (N_17848,N_17364,N_17184);
nand U17849 (N_17849,N_17144,N_17192);
nand U17850 (N_17850,N_17377,N_17491);
and U17851 (N_17851,N_17334,N_17353);
nand U17852 (N_17852,N_17381,N_17132);
and U17853 (N_17853,N_17236,N_17178);
and U17854 (N_17854,N_17335,N_17234);
and U17855 (N_17855,N_17214,N_17372);
nor U17856 (N_17856,N_17012,N_17077);
and U17857 (N_17857,N_17358,N_17280);
and U17858 (N_17858,N_17321,N_17220);
and U17859 (N_17859,N_17042,N_17329);
nor U17860 (N_17860,N_17286,N_17452);
nor U17861 (N_17861,N_17494,N_17247);
or U17862 (N_17862,N_17127,N_17418);
nor U17863 (N_17863,N_17418,N_17052);
or U17864 (N_17864,N_17108,N_17369);
and U17865 (N_17865,N_17131,N_17336);
nand U17866 (N_17866,N_17206,N_17318);
nor U17867 (N_17867,N_17433,N_17422);
nor U17868 (N_17868,N_17397,N_17036);
or U17869 (N_17869,N_17074,N_17379);
nand U17870 (N_17870,N_17461,N_17444);
nand U17871 (N_17871,N_17268,N_17119);
nand U17872 (N_17872,N_17328,N_17067);
nand U17873 (N_17873,N_17266,N_17215);
nand U17874 (N_17874,N_17211,N_17326);
and U17875 (N_17875,N_17182,N_17038);
or U17876 (N_17876,N_17295,N_17450);
or U17877 (N_17877,N_17388,N_17227);
nand U17878 (N_17878,N_17046,N_17172);
or U17879 (N_17879,N_17451,N_17348);
and U17880 (N_17880,N_17367,N_17352);
nor U17881 (N_17881,N_17366,N_17121);
nand U17882 (N_17882,N_17224,N_17420);
nor U17883 (N_17883,N_17354,N_17086);
or U17884 (N_17884,N_17338,N_17048);
or U17885 (N_17885,N_17217,N_17457);
nand U17886 (N_17886,N_17297,N_17355);
nand U17887 (N_17887,N_17462,N_17209);
or U17888 (N_17888,N_17016,N_17085);
and U17889 (N_17889,N_17448,N_17453);
or U17890 (N_17890,N_17253,N_17384);
or U17891 (N_17891,N_17192,N_17102);
or U17892 (N_17892,N_17024,N_17133);
nand U17893 (N_17893,N_17266,N_17166);
or U17894 (N_17894,N_17231,N_17021);
or U17895 (N_17895,N_17148,N_17315);
and U17896 (N_17896,N_17373,N_17292);
and U17897 (N_17897,N_17320,N_17293);
nand U17898 (N_17898,N_17079,N_17427);
nand U17899 (N_17899,N_17003,N_17090);
nor U17900 (N_17900,N_17076,N_17435);
nand U17901 (N_17901,N_17322,N_17194);
nand U17902 (N_17902,N_17138,N_17186);
and U17903 (N_17903,N_17377,N_17220);
nand U17904 (N_17904,N_17452,N_17334);
and U17905 (N_17905,N_17352,N_17160);
or U17906 (N_17906,N_17006,N_17266);
or U17907 (N_17907,N_17419,N_17023);
nor U17908 (N_17908,N_17125,N_17412);
nor U17909 (N_17909,N_17395,N_17167);
or U17910 (N_17910,N_17205,N_17171);
and U17911 (N_17911,N_17437,N_17342);
or U17912 (N_17912,N_17201,N_17051);
or U17913 (N_17913,N_17346,N_17060);
nand U17914 (N_17914,N_17177,N_17302);
nand U17915 (N_17915,N_17307,N_17146);
nand U17916 (N_17916,N_17311,N_17002);
or U17917 (N_17917,N_17100,N_17484);
and U17918 (N_17918,N_17122,N_17494);
nor U17919 (N_17919,N_17135,N_17383);
nand U17920 (N_17920,N_17407,N_17225);
or U17921 (N_17921,N_17439,N_17233);
nor U17922 (N_17922,N_17107,N_17274);
nor U17923 (N_17923,N_17314,N_17164);
and U17924 (N_17924,N_17337,N_17379);
or U17925 (N_17925,N_17248,N_17003);
nor U17926 (N_17926,N_17076,N_17283);
nand U17927 (N_17927,N_17102,N_17034);
or U17928 (N_17928,N_17018,N_17442);
nand U17929 (N_17929,N_17124,N_17125);
nand U17930 (N_17930,N_17050,N_17091);
nand U17931 (N_17931,N_17103,N_17450);
nand U17932 (N_17932,N_17279,N_17032);
nand U17933 (N_17933,N_17333,N_17065);
or U17934 (N_17934,N_17409,N_17116);
and U17935 (N_17935,N_17060,N_17082);
and U17936 (N_17936,N_17372,N_17290);
nor U17937 (N_17937,N_17442,N_17436);
and U17938 (N_17938,N_17143,N_17208);
nor U17939 (N_17939,N_17329,N_17214);
and U17940 (N_17940,N_17254,N_17369);
nand U17941 (N_17941,N_17279,N_17361);
and U17942 (N_17942,N_17434,N_17299);
or U17943 (N_17943,N_17454,N_17047);
nand U17944 (N_17944,N_17244,N_17114);
nor U17945 (N_17945,N_17099,N_17153);
nand U17946 (N_17946,N_17056,N_17179);
or U17947 (N_17947,N_17299,N_17125);
and U17948 (N_17948,N_17213,N_17027);
nand U17949 (N_17949,N_17216,N_17487);
or U17950 (N_17950,N_17363,N_17475);
nor U17951 (N_17951,N_17020,N_17184);
xor U17952 (N_17952,N_17235,N_17491);
or U17953 (N_17953,N_17074,N_17371);
or U17954 (N_17954,N_17498,N_17337);
or U17955 (N_17955,N_17044,N_17060);
and U17956 (N_17956,N_17499,N_17113);
and U17957 (N_17957,N_17251,N_17130);
and U17958 (N_17958,N_17175,N_17376);
or U17959 (N_17959,N_17047,N_17437);
nand U17960 (N_17960,N_17286,N_17067);
or U17961 (N_17961,N_17434,N_17247);
nor U17962 (N_17962,N_17302,N_17112);
or U17963 (N_17963,N_17454,N_17304);
or U17964 (N_17964,N_17018,N_17168);
or U17965 (N_17965,N_17402,N_17237);
nand U17966 (N_17966,N_17294,N_17199);
nor U17967 (N_17967,N_17017,N_17039);
and U17968 (N_17968,N_17336,N_17263);
nand U17969 (N_17969,N_17013,N_17316);
and U17970 (N_17970,N_17448,N_17447);
and U17971 (N_17971,N_17124,N_17122);
nor U17972 (N_17972,N_17296,N_17104);
and U17973 (N_17973,N_17370,N_17018);
nand U17974 (N_17974,N_17430,N_17147);
or U17975 (N_17975,N_17244,N_17364);
nand U17976 (N_17976,N_17009,N_17085);
nor U17977 (N_17977,N_17377,N_17358);
or U17978 (N_17978,N_17265,N_17391);
nor U17979 (N_17979,N_17052,N_17332);
nor U17980 (N_17980,N_17131,N_17281);
and U17981 (N_17981,N_17051,N_17044);
or U17982 (N_17982,N_17453,N_17400);
nand U17983 (N_17983,N_17151,N_17010);
or U17984 (N_17984,N_17400,N_17461);
and U17985 (N_17985,N_17408,N_17073);
or U17986 (N_17986,N_17398,N_17459);
nor U17987 (N_17987,N_17450,N_17023);
nor U17988 (N_17988,N_17132,N_17008);
nor U17989 (N_17989,N_17278,N_17354);
nand U17990 (N_17990,N_17133,N_17284);
and U17991 (N_17991,N_17445,N_17285);
nand U17992 (N_17992,N_17001,N_17075);
or U17993 (N_17993,N_17169,N_17207);
nor U17994 (N_17994,N_17093,N_17282);
or U17995 (N_17995,N_17386,N_17460);
nand U17996 (N_17996,N_17435,N_17443);
nand U17997 (N_17997,N_17039,N_17025);
and U17998 (N_17998,N_17483,N_17238);
or U17999 (N_17999,N_17484,N_17311);
or U18000 (N_18000,N_17743,N_17775);
nand U18001 (N_18001,N_17521,N_17547);
and U18002 (N_18002,N_17638,N_17873);
or U18003 (N_18003,N_17677,N_17757);
xor U18004 (N_18004,N_17527,N_17700);
and U18005 (N_18005,N_17805,N_17748);
nor U18006 (N_18006,N_17566,N_17745);
nor U18007 (N_18007,N_17500,N_17612);
or U18008 (N_18008,N_17905,N_17884);
nand U18009 (N_18009,N_17675,N_17698);
or U18010 (N_18010,N_17518,N_17906);
and U18011 (N_18011,N_17846,N_17550);
or U18012 (N_18012,N_17785,N_17519);
or U18013 (N_18013,N_17690,N_17574);
and U18014 (N_18014,N_17955,N_17716);
nor U18015 (N_18015,N_17866,N_17615);
or U18016 (N_18016,N_17871,N_17933);
or U18017 (N_18017,N_17856,N_17589);
and U18018 (N_18018,N_17825,N_17986);
nand U18019 (N_18019,N_17629,N_17980);
nor U18020 (N_18020,N_17751,N_17625);
or U18021 (N_18021,N_17947,N_17898);
and U18022 (N_18022,N_17809,N_17767);
and U18023 (N_18023,N_17647,N_17790);
nor U18024 (N_18024,N_17822,N_17702);
and U18025 (N_18025,N_17922,N_17842);
or U18026 (N_18026,N_17882,N_17573);
nand U18027 (N_18027,N_17931,N_17605);
nand U18028 (N_18028,N_17758,N_17673);
or U18029 (N_18029,N_17859,N_17685);
nor U18030 (N_18030,N_17771,N_17926);
or U18031 (N_18031,N_17534,N_17900);
or U18032 (N_18032,N_17735,N_17620);
nor U18033 (N_18033,N_17631,N_17575);
and U18034 (N_18034,N_17614,N_17928);
nor U18035 (N_18035,N_17979,N_17542);
nand U18036 (N_18036,N_17881,N_17599);
or U18037 (N_18037,N_17803,N_17813);
and U18038 (N_18038,N_17641,N_17650);
nand U18039 (N_18039,N_17711,N_17594);
or U18040 (N_18040,N_17619,N_17522);
and U18041 (N_18041,N_17988,N_17997);
nor U18042 (N_18042,N_17621,N_17543);
or U18043 (N_18043,N_17808,N_17652);
and U18044 (N_18044,N_17953,N_17705);
nand U18045 (N_18045,N_17667,N_17991);
and U18046 (N_18046,N_17733,N_17932);
nor U18047 (N_18047,N_17731,N_17781);
nand U18048 (N_18048,N_17925,N_17897);
nand U18049 (N_18049,N_17516,N_17965);
nand U18050 (N_18050,N_17510,N_17919);
nand U18051 (N_18051,N_17972,N_17760);
nand U18052 (N_18052,N_17970,N_17869);
nor U18053 (N_18053,N_17969,N_17513);
and U18054 (N_18054,N_17585,N_17904);
nor U18055 (N_18055,N_17936,N_17861);
nor U18056 (N_18056,N_17949,N_17727);
nand U18057 (N_18057,N_17603,N_17989);
nand U18058 (N_18058,N_17964,N_17666);
and U18059 (N_18059,N_17664,N_17627);
or U18060 (N_18060,N_17816,N_17982);
or U18061 (N_18061,N_17699,N_17613);
or U18062 (N_18062,N_17744,N_17867);
or U18063 (N_18063,N_17967,N_17577);
and U18064 (N_18064,N_17604,N_17895);
nand U18065 (N_18065,N_17927,N_17820);
or U18066 (N_18066,N_17801,N_17845);
or U18067 (N_18067,N_17773,N_17930);
xor U18068 (N_18068,N_17517,N_17857);
nand U18069 (N_18069,N_17501,N_17635);
nor U18070 (N_18070,N_17568,N_17862);
nand U18071 (N_18071,N_17506,N_17824);
nor U18072 (N_18072,N_17688,N_17976);
or U18073 (N_18073,N_17946,N_17984);
or U18074 (N_18074,N_17537,N_17794);
and U18075 (N_18075,N_17870,N_17659);
or U18076 (N_18076,N_17956,N_17572);
nor U18077 (N_18077,N_17876,N_17592);
nand U18078 (N_18078,N_17784,N_17749);
nor U18079 (N_18079,N_17832,N_17747);
and U18080 (N_18080,N_17941,N_17774);
or U18081 (N_18081,N_17549,N_17670);
or U18082 (N_18082,N_17732,N_17863);
or U18083 (N_18083,N_17907,N_17893);
and U18084 (N_18084,N_17657,N_17724);
or U18085 (N_18085,N_17512,N_17601);
nor U18086 (N_18086,N_17783,N_17720);
nand U18087 (N_18087,N_17581,N_17660);
nand U18088 (N_18088,N_17722,N_17583);
and U18089 (N_18089,N_17737,N_17899);
or U18090 (N_18090,N_17539,N_17559);
and U18091 (N_18091,N_17715,N_17918);
or U18092 (N_18092,N_17600,N_17750);
and U18093 (N_18093,N_17562,N_17954);
nand U18094 (N_18094,N_17942,N_17709);
nand U18095 (N_18095,N_17695,N_17879);
and U18096 (N_18096,N_17786,N_17766);
nor U18097 (N_18097,N_17944,N_17890);
nor U18098 (N_18098,N_17836,N_17548);
nand U18099 (N_18099,N_17913,N_17741);
nor U18100 (N_18100,N_17502,N_17520);
nor U18101 (N_18101,N_17530,N_17514);
and U18102 (N_18102,N_17811,N_17754);
nor U18103 (N_18103,N_17579,N_17691);
nand U18104 (N_18104,N_17687,N_17838);
or U18105 (N_18105,N_17992,N_17847);
nand U18106 (N_18106,N_17830,N_17819);
nor U18107 (N_18107,N_17778,N_17633);
nand U18108 (N_18108,N_17681,N_17987);
nor U18109 (N_18109,N_17901,N_17787);
nor U18110 (N_18110,N_17602,N_17843);
nor U18111 (N_18111,N_17523,N_17763);
nand U18112 (N_18112,N_17655,N_17597);
nand U18113 (N_18113,N_17776,N_17834);
and U18114 (N_18114,N_17511,N_17804);
nand U18115 (N_18115,N_17990,N_17628);
nor U18116 (N_18116,N_17833,N_17759);
or U18117 (N_18117,N_17772,N_17903);
nor U18118 (N_18118,N_17515,N_17817);
nand U18119 (N_18119,N_17563,N_17639);
nor U18120 (N_18120,N_17792,N_17995);
nor U18121 (N_18121,N_17590,N_17915);
or U18122 (N_18122,N_17938,N_17793);
or U18123 (N_18123,N_17841,N_17536);
or U18124 (N_18124,N_17999,N_17694);
nand U18125 (N_18125,N_17689,N_17962);
and U18126 (N_18126,N_17526,N_17560);
nand U18127 (N_18127,N_17648,N_17739);
or U18128 (N_18128,N_17762,N_17826);
nand U18129 (N_18129,N_17827,N_17570);
nand U18130 (N_18130,N_17780,N_17571);
nor U18131 (N_18131,N_17883,N_17552);
or U18132 (N_18132,N_17975,N_17917);
nand U18133 (N_18133,N_17889,N_17504);
nand U18134 (N_18134,N_17935,N_17524);
and U18135 (N_18135,N_17914,N_17634);
nor U18136 (N_18136,N_17654,N_17551);
or U18137 (N_18137,N_17706,N_17582);
nor U18138 (N_18138,N_17503,N_17789);
and U18139 (N_18139,N_17959,N_17874);
and U18140 (N_18140,N_17981,N_17740);
or U18141 (N_18141,N_17908,N_17978);
and U18142 (N_18142,N_17966,N_17920);
and U18143 (N_18143,N_17544,N_17802);
and U18144 (N_18144,N_17676,N_17977);
nor U18145 (N_18145,N_17593,N_17616);
or U18146 (N_18146,N_17996,N_17645);
nand U18147 (N_18147,N_17578,N_17823);
nor U18148 (N_18148,N_17864,N_17814);
nand U18149 (N_18149,N_17952,N_17661);
nor U18150 (N_18150,N_17929,N_17880);
nor U18151 (N_18151,N_17642,N_17858);
nand U18152 (N_18152,N_17958,N_17726);
or U18153 (N_18153,N_17692,N_17561);
nor U18154 (N_18154,N_17665,N_17878);
nand U18155 (N_18155,N_17565,N_17556);
and U18156 (N_18156,N_17658,N_17831);
and U18157 (N_18157,N_17939,N_17607);
nor U18158 (N_18158,N_17753,N_17788);
or U18159 (N_18159,N_17569,N_17674);
nor U18160 (N_18160,N_17974,N_17531);
nand U18161 (N_18161,N_17892,N_17678);
or U18162 (N_18162,N_17668,N_17679);
or U18163 (N_18163,N_17968,N_17818);
nand U18164 (N_18164,N_17948,N_17921);
and U18165 (N_18165,N_17580,N_17940);
or U18166 (N_18166,N_17528,N_17855);
and U18167 (N_18167,N_17896,N_17606);
and U18168 (N_18168,N_17672,N_17937);
nand U18169 (N_18169,N_17505,N_17640);
or U18170 (N_18170,N_17718,N_17971);
nand U18171 (N_18171,N_17957,N_17755);
or U18172 (N_18172,N_17800,N_17555);
nor U18173 (N_18173,N_17799,N_17909);
nor U18174 (N_18174,N_17782,N_17529);
nor U18175 (N_18175,N_17951,N_17742);
and U18176 (N_18176,N_17721,N_17894);
or U18177 (N_18177,N_17916,N_17837);
nand U18178 (N_18178,N_17910,N_17624);
nor U18179 (N_18179,N_17777,N_17696);
and U18180 (N_18180,N_17545,N_17872);
nand U18181 (N_18181,N_17911,N_17587);
or U18182 (N_18182,N_17507,N_17643);
nor U18183 (N_18183,N_17626,N_17752);
nand U18184 (N_18184,N_17769,N_17934);
or U18185 (N_18185,N_17710,N_17714);
or U18186 (N_18186,N_17888,N_17853);
nor U18187 (N_18187,N_17779,N_17798);
and U18188 (N_18188,N_17584,N_17712);
and U18189 (N_18189,N_17564,N_17595);
nor U18190 (N_18190,N_17983,N_17756);
nor U18191 (N_18191,N_17963,N_17553);
nor U18192 (N_18192,N_17795,N_17651);
nor U18193 (N_18193,N_17994,N_17993);
or U18194 (N_18194,N_17588,N_17693);
or U18195 (N_18195,N_17596,N_17684);
or U18196 (N_18196,N_17796,N_17950);
nor U18197 (N_18197,N_17868,N_17567);
and U18198 (N_18198,N_17812,N_17765);
and U18199 (N_18199,N_17623,N_17703);
nor U18200 (N_18200,N_17973,N_17761);
nand U18201 (N_18201,N_17828,N_17707);
nor U18202 (N_18202,N_17865,N_17807);
or U18203 (N_18203,N_17886,N_17509);
nor U18204 (N_18204,N_17558,N_17637);
or U18205 (N_18205,N_17821,N_17704);
and U18206 (N_18206,N_17618,N_17686);
nor U18207 (N_18207,N_17554,N_17508);
xor U18208 (N_18208,N_17546,N_17630);
and U18209 (N_18209,N_17960,N_17860);
nor U18210 (N_18210,N_17924,N_17653);
nand U18211 (N_18211,N_17998,N_17611);
and U18212 (N_18212,N_17636,N_17851);
and U18213 (N_18213,N_17840,N_17746);
nand U18214 (N_18214,N_17540,N_17810);
and U18215 (N_18215,N_17912,N_17701);
nor U18216 (N_18216,N_17945,N_17610);
or U18217 (N_18217,N_17656,N_17525);
nor U18218 (N_18218,N_17644,N_17854);
and U18219 (N_18219,N_17533,N_17849);
nand U18220 (N_18220,N_17680,N_17697);
and U18221 (N_18221,N_17738,N_17791);
and U18222 (N_18222,N_17535,N_17961);
and U18223 (N_18223,N_17815,N_17850);
nand U18224 (N_18224,N_17891,N_17887);
or U18225 (N_18225,N_17729,N_17797);
nor U18226 (N_18226,N_17844,N_17591);
and U18227 (N_18227,N_17770,N_17806);
or U18228 (N_18228,N_17829,N_17835);
nor U18229 (N_18229,N_17839,N_17541);
nand U18230 (N_18230,N_17708,N_17730);
nand U18231 (N_18231,N_17877,N_17622);
or U18232 (N_18232,N_17725,N_17734);
or U18233 (N_18233,N_17609,N_17683);
nand U18234 (N_18234,N_17649,N_17713);
nand U18235 (N_18235,N_17923,N_17717);
nor U18236 (N_18236,N_17682,N_17586);
and U18237 (N_18237,N_17617,N_17669);
or U18238 (N_18238,N_17557,N_17608);
nor U18239 (N_18239,N_17663,N_17723);
or U18240 (N_18240,N_17848,N_17885);
or U18241 (N_18241,N_17943,N_17671);
or U18242 (N_18242,N_17719,N_17875);
nand U18243 (N_18243,N_17576,N_17985);
or U18244 (N_18244,N_17902,N_17538);
and U18245 (N_18245,N_17662,N_17598);
nand U18246 (N_18246,N_17728,N_17736);
nand U18247 (N_18247,N_17768,N_17646);
nor U18248 (N_18248,N_17632,N_17852);
or U18249 (N_18249,N_17532,N_17764);
nand U18250 (N_18250,N_17508,N_17828);
or U18251 (N_18251,N_17936,N_17515);
nand U18252 (N_18252,N_17683,N_17948);
and U18253 (N_18253,N_17894,N_17773);
xor U18254 (N_18254,N_17819,N_17684);
and U18255 (N_18255,N_17917,N_17825);
or U18256 (N_18256,N_17956,N_17626);
nor U18257 (N_18257,N_17538,N_17659);
nor U18258 (N_18258,N_17527,N_17539);
or U18259 (N_18259,N_17716,N_17873);
nand U18260 (N_18260,N_17659,N_17841);
nand U18261 (N_18261,N_17997,N_17758);
nand U18262 (N_18262,N_17875,N_17935);
and U18263 (N_18263,N_17585,N_17706);
nor U18264 (N_18264,N_17853,N_17844);
nor U18265 (N_18265,N_17758,N_17830);
nor U18266 (N_18266,N_17559,N_17791);
nand U18267 (N_18267,N_17630,N_17700);
nor U18268 (N_18268,N_17929,N_17963);
nand U18269 (N_18269,N_17861,N_17681);
and U18270 (N_18270,N_17578,N_17752);
and U18271 (N_18271,N_17724,N_17654);
nor U18272 (N_18272,N_17664,N_17618);
and U18273 (N_18273,N_17521,N_17934);
nor U18274 (N_18274,N_17750,N_17989);
or U18275 (N_18275,N_17713,N_17757);
nor U18276 (N_18276,N_17629,N_17762);
and U18277 (N_18277,N_17640,N_17741);
nand U18278 (N_18278,N_17876,N_17706);
or U18279 (N_18279,N_17899,N_17787);
nand U18280 (N_18280,N_17546,N_17945);
nand U18281 (N_18281,N_17735,N_17716);
nand U18282 (N_18282,N_17647,N_17872);
nor U18283 (N_18283,N_17832,N_17868);
nor U18284 (N_18284,N_17980,N_17640);
and U18285 (N_18285,N_17870,N_17752);
and U18286 (N_18286,N_17743,N_17624);
and U18287 (N_18287,N_17733,N_17769);
nand U18288 (N_18288,N_17522,N_17590);
nand U18289 (N_18289,N_17676,N_17518);
nand U18290 (N_18290,N_17815,N_17646);
and U18291 (N_18291,N_17566,N_17729);
nand U18292 (N_18292,N_17640,N_17800);
or U18293 (N_18293,N_17641,N_17881);
and U18294 (N_18294,N_17978,N_17907);
nand U18295 (N_18295,N_17589,N_17605);
nand U18296 (N_18296,N_17541,N_17726);
nand U18297 (N_18297,N_17815,N_17950);
nor U18298 (N_18298,N_17595,N_17869);
nor U18299 (N_18299,N_17732,N_17606);
nor U18300 (N_18300,N_17533,N_17693);
xor U18301 (N_18301,N_17686,N_17811);
nor U18302 (N_18302,N_17940,N_17973);
and U18303 (N_18303,N_17777,N_17571);
nand U18304 (N_18304,N_17960,N_17791);
xnor U18305 (N_18305,N_17705,N_17981);
and U18306 (N_18306,N_17843,N_17943);
or U18307 (N_18307,N_17585,N_17966);
and U18308 (N_18308,N_17960,N_17862);
nand U18309 (N_18309,N_17861,N_17807);
nor U18310 (N_18310,N_17740,N_17760);
nor U18311 (N_18311,N_17746,N_17702);
or U18312 (N_18312,N_17831,N_17680);
and U18313 (N_18313,N_17518,N_17993);
xor U18314 (N_18314,N_17770,N_17909);
nor U18315 (N_18315,N_17771,N_17795);
nand U18316 (N_18316,N_17842,N_17994);
or U18317 (N_18317,N_17846,N_17583);
nand U18318 (N_18318,N_17520,N_17892);
nand U18319 (N_18319,N_17799,N_17540);
nor U18320 (N_18320,N_17930,N_17714);
nor U18321 (N_18321,N_17677,N_17832);
nand U18322 (N_18322,N_17679,N_17508);
and U18323 (N_18323,N_17870,N_17826);
and U18324 (N_18324,N_17977,N_17913);
or U18325 (N_18325,N_17681,N_17625);
nor U18326 (N_18326,N_17592,N_17934);
nor U18327 (N_18327,N_17766,N_17908);
or U18328 (N_18328,N_17757,N_17587);
or U18329 (N_18329,N_17861,N_17887);
and U18330 (N_18330,N_17647,N_17624);
nand U18331 (N_18331,N_17612,N_17576);
and U18332 (N_18332,N_17786,N_17624);
nor U18333 (N_18333,N_17680,N_17578);
or U18334 (N_18334,N_17506,N_17819);
nand U18335 (N_18335,N_17780,N_17981);
xor U18336 (N_18336,N_17861,N_17656);
nor U18337 (N_18337,N_17611,N_17509);
or U18338 (N_18338,N_17525,N_17719);
nor U18339 (N_18339,N_17661,N_17637);
nand U18340 (N_18340,N_17604,N_17994);
nand U18341 (N_18341,N_17787,N_17685);
and U18342 (N_18342,N_17792,N_17867);
nor U18343 (N_18343,N_17683,N_17719);
or U18344 (N_18344,N_17736,N_17531);
and U18345 (N_18345,N_17977,N_17635);
or U18346 (N_18346,N_17927,N_17511);
and U18347 (N_18347,N_17912,N_17592);
nor U18348 (N_18348,N_17858,N_17557);
and U18349 (N_18349,N_17755,N_17557);
nor U18350 (N_18350,N_17654,N_17696);
and U18351 (N_18351,N_17698,N_17778);
nor U18352 (N_18352,N_17628,N_17730);
nor U18353 (N_18353,N_17617,N_17503);
nand U18354 (N_18354,N_17928,N_17816);
or U18355 (N_18355,N_17868,N_17797);
nor U18356 (N_18356,N_17770,N_17546);
and U18357 (N_18357,N_17690,N_17851);
nor U18358 (N_18358,N_17552,N_17769);
nor U18359 (N_18359,N_17673,N_17685);
or U18360 (N_18360,N_17926,N_17721);
nor U18361 (N_18361,N_17983,N_17804);
nor U18362 (N_18362,N_17662,N_17555);
nand U18363 (N_18363,N_17790,N_17697);
or U18364 (N_18364,N_17807,N_17750);
or U18365 (N_18365,N_17715,N_17567);
nor U18366 (N_18366,N_17953,N_17819);
nand U18367 (N_18367,N_17864,N_17563);
nand U18368 (N_18368,N_17909,N_17835);
nand U18369 (N_18369,N_17799,N_17884);
nor U18370 (N_18370,N_17916,N_17770);
and U18371 (N_18371,N_17908,N_17882);
nand U18372 (N_18372,N_17506,N_17751);
or U18373 (N_18373,N_17970,N_17630);
nor U18374 (N_18374,N_17967,N_17936);
nand U18375 (N_18375,N_17557,N_17741);
nor U18376 (N_18376,N_17577,N_17726);
nor U18377 (N_18377,N_17850,N_17784);
nand U18378 (N_18378,N_17556,N_17524);
nor U18379 (N_18379,N_17833,N_17687);
or U18380 (N_18380,N_17557,N_17891);
or U18381 (N_18381,N_17671,N_17639);
xnor U18382 (N_18382,N_17571,N_17696);
and U18383 (N_18383,N_17678,N_17960);
xnor U18384 (N_18384,N_17787,N_17890);
and U18385 (N_18385,N_17558,N_17679);
and U18386 (N_18386,N_17512,N_17640);
nand U18387 (N_18387,N_17906,N_17677);
nor U18388 (N_18388,N_17711,N_17927);
nor U18389 (N_18389,N_17771,N_17950);
nand U18390 (N_18390,N_17570,N_17839);
nor U18391 (N_18391,N_17839,N_17574);
and U18392 (N_18392,N_17652,N_17642);
or U18393 (N_18393,N_17562,N_17684);
or U18394 (N_18394,N_17530,N_17913);
or U18395 (N_18395,N_17850,N_17721);
and U18396 (N_18396,N_17914,N_17909);
and U18397 (N_18397,N_17618,N_17953);
and U18398 (N_18398,N_17820,N_17771);
or U18399 (N_18399,N_17697,N_17597);
nand U18400 (N_18400,N_17658,N_17940);
or U18401 (N_18401,N_17602,N_17694);
or U18402 (N_18402,N_17547,N_17688);
nand U18403 (N_18403,N_17984,N_17596);
nor U18404 (N_18404,N_17748,N_17854);
or U18405 (N_18405,N_17874,N_17750);
and U18406 (N_18406,N_17858,N_17606);
and U18407 (N_18407,N_17592,N_17514);
nand U18408 (N_18408,N_17866,N_17916);
and U18409 (N_18409,N_17791,N_17804);
and U18410 (N_18410,N_17953,N_17990);
or U18411 (N_18411,N_17598,N_17538);
nand U18412 (N_18412,N_17639,N_17617);
nand U18413 (N_18413,N_17629,N_17806);
or U18414 (N_18414,N_17930,N_17994);
and U18415 (N_18415,N_17943,N_17700);
and U18416 (N_18416,N_17786,N_17539);
nand U18417 (N_18417,N_17841,N_17535);
or U18418 (N_18418,N_17901,N_17781);
nor U18419 (N_18419,N_17661,N_17795);
nor U18420 (N_18420,N_17665,N_17998);
or U18421 (N_18421,N_17935,N_17880);
nor U18422 (N_18422,N_17517,N_17837);
nand U18423 (N_18423,N_17620,N_17708);
or U18424 (N_18424,N_17715,N_17619);
and U18425 (N_18425,N_17889,N_17572);
nor U18426 (N_18426,N_17865,N_17526);
and U18427 (N_18427,N_17590,N_17794);
or U18428 (N_18428,N_17519,N_17685);
and U18429 (N_18429,N_17856,N_17692);
or U18430 (N_18430,N_17970,N_17996);
or U18431 (N_18431,N_17853,N_17514);
nand U18432 (N_18432,N_17783,N_17679);
or U18433 (N_18433,N_17581,N_17548);
and U18434 (N_18434,N_17593,N_17940);
or U18435 (N_18435,N_17843,N_17858);
and U18436 (N_18436,N_17504,N_17907);
or U18437 (N_18437,N_17774,N_17746);
or U18438 (N_18438,N_17753,N_17963);
nand U18439 (N_18439,N_17683,N_17512);
and U18440 (N_18440,N_17585,N_17718);
nor U18441 (N_18441,N_17676,N_17891);
nand U18442 (N_18442,N_17551,N_17685);
nand U18443 (N_18443,N_17842,N_17921);
nand U18444 (N_18444,N_17843,N_17741);
nor U18445 (N_18445,N_17743,N_17607);
nor U18446 (N_18446,N_17642,N_17830);
nand U18447 (N_18447,N_17892,N_17506);
or U18448 (N_18448,N_17921,N_17750);
nor U18449 (N_18449,N_17559,N_17757);
nand U18450 (N_18450,N_17725,N_17583);
nor U18451 (N_18451,N_17980,N_17793);
or U18452 (N_18452,N_17925,N_17789);
or U18453 (N_18453,N_17930,N_17711);
and U18454 (N_18454,N_17844,N_17947);
or U18455 (N_18455,N_17524,N_17960);
and U18456 (N_18456,N_17863,N_17600);
or U18457 (N_18457,N_17546,N_17569);
and U18458 (N_18458,N_17995,N_17647);
and U18459 (N_18459,N_17527,N_17634);
and U18460 (N_18460,N_17951,N_17588);
nand U18461 (N_18461,N_17667,N_17569);
and U18462 (N_18462,N_17744,N_17559);
nor U18463 (N_18463,N_17979,N_17564);
nor U18464 (N_18464,N_17862,N_17781);
nor U18465 (N_18465,N_17645,N_17817);
nor U18466 (N_18466,N_17504,N_17521);
nand U18467 (N_18467,N_17690,N_17810);
nor U18468 (N_18468,N_17622,N_17957);
and U18469 (N_18469,N_17883,N_17841);
nand U18470 (N_18470,N_17605,N_17882);
or U18471 (N_18471,N_17915,N_17816);
or U18472 (N_18472,N_17557,N_17764);
and U18473 (N_18473,N_17763,N_17637);
or U18474 (N_18474,N_17737,N_17963);
nand U18475 (N_18475,N_17714,N_17750);
nand U18476 (N_18476,N_17545,N_17798);
and U18477 (N_18477,N_17554,N_17852);
or U18478 (N_18478,N_17588,N_17776);
nor U18479 (N_18479,N_17772,N_17954);
or U18480 (N_18480,N_17692,N_17923);
and U18481 (N_18481,N_17942,N_17722);
nand U18482 (N_18482,N_17907,N_17595);
or U18483 (N_18483,N_17656,N_17766);
nand U18484 (N_18484,N_17996,N_17579);
nor U18485 (N_18485,N_17740,N_17952);
nor U18486 (N_18486,N_17715,N_17653);
or U18487 (N_18487,N_17541,N_17963);
or U18488 (N_18488,N_17941,N_17853);
or U18489 (N_18489,N_17751,N_17727);
nand U18490 (N_18490,N_17755,N_17659);
nor U18491 (N_18491,N_17549,N_17970);
and U18492 (N_18492,N_17892,N_17675);
and U18493 (N_18493,N_17857,N_17555);
nor U18494 (N_18494,N_17889,N_17653);
nand U18495 (N_18495,N_17889,N_17575);
or U18496 (N_18496,N_17548,N_17681);
or U18497 (N_18497,N_17847,N_17522);
and U18498 (N_18498,N_17969,N_17989);
nor U18499 (N_18499,N_17723,N_17871);
nor U18500 (N_18500,N_18237,N_18051);
or U18501 (N_18501,N_18132,N_18014);
and U18502 (N_18502,N_18311,N_18407);
nand U18503 (N_18503,N_18251,N_18425);
nand U18504 (N_18504,N_18163,N_18182);
and U18505 (N_18505,N_18245,N_18455);
or U18506 (N_18506,N_18027,N_18316);
nor U18507 (N_18507,N_18491,N_18437);
nand U18508 (N_18508,N_18441,N_18410);
or U18509 (N_18509,N_18204,N_18208);
or U18510 (N_18510,N_18092,N_18254);
nor U18511 (N_18511,N_18498,N_18247);
nand U18512 (N_18512,N_18057,N_18406);
and U18513 (N_18513,N_18065,N_18048);
nand U18514 (N_18514,N_18099,N_18398);
or U18515 (N_18515,N_18438,N_18330);
nand U18516 (N_18516,N_18055,N_18058);
or U18517 (N_18517,N_18395,N_18078);
nor U18518 (N_18518,N_18201,N_18120);
nand U18519 (N_18519,N_18459,N_18453);
nor U18520 (N_18520,N_18292,N_18326);
and U18521 (N_18521,N_18177,N_18412);
nand U18522 (N_18522,N_18362,N_18135);
and U18523 (N_18523,N_18273,N_18130);
nor U18524 (N_18524,N_18107,N_18216);
and U18525 (N_18525,N_18198,N_18018);
or U18526 (N_18526,N_18408,N_18206);
nor U18527 (N_18527,N_18463,N_18084);
nor U18528 (N_18528,N_18187,N_18282);
and U18529 (N_18529,N_18169,N_18286);
nand U18530 (N_18530,N_18172,N_18059);
nand U18531 (N_18531,N_18225,N_18307);
nand U18532 (N_18532,N_18195,N_18497);
nor U18533 (N_18533,N_18464,N_18222);
or U18534 (N_18534,N_18287,N_18006);
nor U18535 (N_18535,N_18147,N_18250);
nor U18536 (N_18536,N_18343,N_18233);
nor U18537 (N_18537,N_18476,N_18019);
and U18538 (N_18538,N_18365,N_18496);
or U18539 (N_18539,N_18461,N_18442);
or U18540 (N_18540,N_18089,N_18348);
nor U18541 (N_18541,N_18414,N_18114);
and U18542 (N_18542,N_18475,N_18429);
or U18543 (N_18543,N_18054,N_18259);
nand U18544 (N_18544,N_18255,N_18210);
nand U18545 (N_18545,N_18199,N_18258);
nor U18546 (N_18546,N_18062,N_18073);
or U18547 (N_18547,N_18028,N_18495);
or U18548 (N_18548,N_18241,N_18377);
nand U18549 (N_18549,N_18191,N_18007);
or U18550 (N_18550,N_18074,N_18445);
or U18551 (N_18551,N_18189,N_18378);
and U18552 (N_18552,N_18372,N_18448);
and U18553 (N_18553,N_18327,N_18040);
or U18554 (N_18554,N_18338,N_18068);
and U18555 (N_18555,N_18389,N_18413);
and U18556 (N_18556,N_18149,N_18269);
nand U18557 (N_18557,N_18175,N_18226);
and U18558 (N_18558,N_18129,N_18390);
nor U18559 (N_18559,N_18318,N_18275);
nand U18560 (N_18560,N_18298,N_18309);
or U18561 (N_18561,N_18447,N_18080);
or U18562 (N_18562,N_18053,N_18482);
nor U18563 (N_18563,N_18271,N_18391);
nand U18564 (N_18564,N_18203,N_18202);
or U18565 (N_18565,N_18076,N_18218);
nor U18566 (N_18566,N_18388,N_18263);
and U18567 (N_18567,N_18399,N_18394);
nand U18568 (N_18568,N_18095,N_18050);
and U18569 (N_18569,N_18243,N_18017);
or U18570 (N_18570,N_18492,N_18402);
nand U18571 (N_18571,N_18479,N_18490);
nor U18572 (N_18572,N_18368,N_18001);
and U18573 (N_18573,N_18321,N_18088);
nand U18574 (N_18574,N_18457,N_18026);
nand U18575 (N_18575,N_18002,N_18416);
nor U18576 (N_18576,N_18284,N_18151);
or U18577 (N_18577,N_18443,N_18152);
nor U18578 (N_18578,N_18252,N_18133);
nor U18579 (N_18579,N_18436,N_18109);
or U18580 (N_18580,N_18117,N_18168);
nand U18581 (N_18581,N_18484,N_18323);
nor U18582 (N_18582,N_18383,N_18462);
and U18583 (N_18583,N_18353,N_18184);
or U18584 (N_18584,N_18229,N_18033);
or U18585 (N_18585,N_18194,N_18385);
nor U18586 (N_18586,N_18418,N_18417);
and U18587 (N_18587,N_18320,N_18483);
or U18588 (N_18588,N_18473,N_18344);
and U18589 (N_18589,N_18106,N_18003);
or U18590 (N_18590,N_18232,N_18127);
and U18591 (N_18591,N_18224,N_18192);
nand U18592 (N_18592,N_18242,N_18270);
or U18593 (N_18593,N_18043,N_18119);
nor U18594 (N_18594,N_18113,N_18214);
and U18595 (N_18595,N_18023,N_18397);
nand U18596 (N_18596,N_18261,N_18101);
or U18597 (N_18597,N_18052,N_18086);
or U18598 (N_18598,N_18238,N_18487);
nand U18599 (N_18599,N_18347,N_18422);
nand U18600 (N_18600,N_18349,N_18474);
and U18601 (N_18601,N_18393,N_18249);
or U18602 (N_18602,N_18016,N_18167);
nor U18603 (N_18603,N_18010,N_18031);
nand U18604 (N_18604,N_18341,N_18087);
nor U18605 (N_18605,N_18278,N_18209);
nor U18606 (N_18606,N_18221,N_18339);
nand U18607 (N_18607,N_18403,N_18193);
and U18608 (N_18608,N_18317,N_18156);
or U18609 (N_18609,N_18302,N_18319);
or U18610 (N_18610,N_18162,N_18379);
nor U18611 (N_18611,N_18313,N_18337);
or U18612 (N_18612,N_18144,N_18158);
nor U18613 (N_18613,N_18426,N_18432);
nand U18614 (N_18614,N_18098,N_18046);
nand U18615 (N_18615,N_18430,N_18069);
and U18616 (N_18616,N_18246,N_18472);
or U18617 (N_18617,N_18021,N_18289);
nand U18618 (N_18618,N_18427,N_18067);
and U18619 (N_18619,N_18424,N_18469);
xor U18620 (N_18620,N_18035,N_18082);
and U18621 (N_18621,N_18387,N_18126);
and U18622 (N_18622,N_18439,N_18124);
and U18623 (N_18623,N_18421,N_18244);
nand U18624 (N_18624,N_18083,N_18093);
nand U18625 (N_18625,N_18139,N_18205);
and U18626 (N_18626,N_18303,N_18234);
and U18627 (N_18627,N_18036,N_18111);
or U18628 (N_18628,N_18297,N_18037);
or U18629 (N_18629,N_18489,N_18174);
and U18630 (N_18630,N_18071,N_18200);
nor U18631 (N_18631,N_18161,N_18364);
and U18632 (N_18632,N_18142,N_18308);
nor U18633 (N_18633,N_18154,N_18000);
and U18634 (N_18634,N_18304,N_18435);
nand U18635 (N_18635,N_18207,N_18150);
and U18636 (N_18636,N_18056,N_18440);
or U18637 (N_18637,N_18405,N_18470);
nand U18638 (N_18638,N_18256,N_18186);
or U18639 (N_18639,N_18257,N_18009);
xor U18640 (N_18640,N_18110,N_18179);
nor U18641 (N_18641,N_18239,N_18166);
and U18642 (N_18642,N_18108,N_18356);
or U18643 (N_18643,N_18228,N_18456);
nand U18644 (N_18644,N_18183,N_18091);
nor U18645 (N_18645,N_18293,N_18220);
and U18646 (N_18646,N_18012,N_18291);
or U18647 (N_18647,N_18454,N_18382);
nor U18648 (N_18648,N_18159,N_18478);
and U18649 (N_18649,N_18351,N_18411);
nand U18650 (N_18650,N_18369,N_18038);
and U18651 (N_18651,N_18346,N_18419);
and U18652 (N_18652,N_18141,N_18451);
nor U18653 (N_18653,N_18165,N_18452);
nand U18654 (N_18654,N_18140,N_18359);
or U18655 (N_18655,N_18458,N_18336);
and U18656 (N_18656,N_18283,N_18115);
and U18657 (N_18657,N_18375,N_18279);
or U18658 (N_18658,N_18400,N_18294);
and U18659 (N_18659,N_18248,N_18094);
nand U18660 (N_18660,N_18466,N_18404);
nor U18661 (N_18661,N_18075,N_18471);
nand U18662 (N_18662,N_18380,N_18328);
nor U18663 (N_18663,N_18285,N_18295);
and U18664 (N_18664,N_18240,N_18164);
and U18665 (N_18665,N_18125,N_18301);
nor U18666 (N_18666,N_18288,N_18434);
nand U18667 (N_18667,N_18123,N_18034);
nand U18668 (N_18668,N_18486,N_18180);
xor U18669 (N_18669,N_18181,N_18314);
and U18670 (N_18670,N_18116,N_18290);
or U18671 (N_18671,N_18153,N_18047);
nand U18672 (N_18672,N_18370,N_18433);
nand U18673 (N_18673,N_18299,N_18219);
or U18674 (N_18674,N_18102,N_18020);
or U18675 (N_18675,N_18444,N_18468);
nor U18676 (N_18676,N_18061,N_18333);
and U18677 (N_18677,N_18386,N_18100);
nor U18678 (N_18678,N_18431,N_18305);
nor U18679 (N_18679,N_18231,N_18262);
or U18680 (N_18680,N_18090,N_18396);
or U18681 (N_18681,N_18460,N_18121);
or U18682 (N_18682,N_18276,N_18188);
nor U18683 (N_18683,N_18401,N_18494);
nor U18684 (N_18684,N_18296,N_18310);
and U18685 (N_18685,N_18260,N_18097);
and U18686 (N_18686,N_18267,N_18428);
nand U18687 (N_18687,N_18392,N_18358);
nand U18688 (N_18688,N_18281,N_18064);
nand U18689 (N_18689,N_18485,N_18420);
and U18690 (N_18690,N_18081,N_18024);
nand U18691 (N_18691,N_18331,N_18063);
and U18692 (N_18692,N_18143,N_18213);
nor U18693 (N_18693,N_18384,N_18361);
and U18694 (N_18694,N_18367,N_18423);
nand U18695 (N_18695,N_18060,N_18176);
and U18696 (N_18696,N_18446,N_18079);
nor U18697 (N_18697,N_18042,N_18355);
nor U18698 (N_18698,N_18335,N_18465);
and U18699 (N_18699,N_18415,N_18145);
nor U18700 (N_18700,N_18322,N_18312);
nor U18701 (N_18701,N_18467,N_18105);
or U18702 (N_18702,N_18072,N_18373);
and U18703 (N_18703,N_18266,N_18357);
nand U18704 (N_18704,N_18077,N_18274);
nor U18705 (N_18705,N_18196,N_18134);
or U18706 (N_18706,N_18315,N_18155);
or U18707 (N_18707,N_18157,N_18374);
nand U18708 (N_18708,N_18146,N_18025);
or U18709 (N_18709,N_18136,N_18215);
nor U18710 (N_18710,N_18211,N_18170);
or U18711 (N_18711,N_18280,N_18268);
nor U18712 (N_18712,N_18197,N_18371);
nor U18713 (N_18713,N_18178,N_18324);
or U18714 (N_18714,N_18131,N_18223);
nor U18715 (N_18715,N_18148,N_18477);
and U18716 (N_18716,N_18481,N_18488);
and U18717 (N_18717,N_18230,N_18352);
and U18718 (N_18718,N_18070,N_18300);
or U18719 (N_18719,N_18044,N_18029);
or U18720 (N_18720,N_18015,N_18039);
and U18721 (N_18721,N_18272,N_18409);
nand U18722 (N_18722,N_18340,N_18171);
and U18723 (N_18723,N_18066,N_18118);
or U18724 (N_18724,N_18185,N_18306);
and U18725 (N_18725,N_18360,N_18325);
and U18726 (N_18726,N_18480,N_18013);
nand U18727 (N_18727,N_18264,N_18137);
nor U18728 (N_18728,N_18190,N_18045);
and U18729 (N_18729,N_18253,N_18104);
and U18730 (N_18730,N_18332,N_18499);
nor U18731 (N_18731,N_18008,N_18493);
nor U18732 (N_18732,N_18096,N_18212);
nor U18733 (N_18733,N_18032,N_18265);
and U18734 (N_18734,N_18329,N_18030);
nand U18735 (N_18735,N_18049,N_18450);
nor U18736 (N_18736,N_18004,N_18138);
or U18737 (N_18737,N_18128,N_18217);
nor U18738 (N_18738,N_18235,N_18112);
nand U18739 (N_18739,N_18173,N_18376);
and U18740 (N_18740,N_18122,N_18277);
and U18741 (N_18741,N_18085,N_18366);
nand U18742 (N_18742,N_18381,N_18350);
nor U18743 (N_18743,N_18345,N_18005);
nor U18744 (N_18744,N_18449,N_18041);
nor U18745 (N_18745,N_18227,N_18236);
nor U18746 (N_18746,N_18160,N_18363);
or U18747 (N_18747,N_18022,N_18342);
nor U18748 (N_18748,N_18011,N_18103);
xnor U18749 (N_18749,N_18354,N_18334);
nand U18750 (N_18750,N_18087,N_18054);
nor U18751 (N_18751,N_18206,N_18444);
or U18752 (N_18752,N_18022,N_18123);
nor U18753 (N_18753,N_18173,N_18056);
nor U18754 (N_18754,N_18224,N_18184);
and U18755 (N_18755,N_18363,N_18058);
nand U18756 (N_18756,N_18291,N_18013);
nand U18757 (N_18757,N_18029,N_18430);
or U18758 (N_18758,N_18040,N_18003);
or U18759 (N_18759,N_18004,N_18134);
or U18760 (N_18760,N_18180,N_18244);
nor U18761 (N_18761,N_18097,N_18150);
and U18762 (N_18762,N_18171,N_18229);
nand U18763 (N_18763,N_18461,N_18335);
and U18764 (N_18764,N_18113,N_18061);
nand U18765 (N_18765,N_18050,N_18462);
and U18766 (N_18766,N_18111,N_18034);
and U18767 (N_18767,N_18302,N_18488);
nor U18768 (N_18768,N_18095,N_18107);
nor U18769 (N_18769,N_18152,N_18383);
nor U18770 (N_18770,N_18419,N_18107);
nand U18771 (N_18771,N_18347,N_18372);
nand U18772 (N_18772,N_18378,N_18381);
and U18773 (N_18773,N_18436,N_18246);
or U18774 (N_18774,N_18314,N_18131);
or U18775 (N_18775,N_18470,N_18210);
or U18776 (N_18776,N_18296,N_18242);
xor U18777 (N_18777,N_18298,N_18337);
and U18778 (N_18778,N_18422,N_18367);
nand U18779 (N_18779,N_18452,N_18083);
and U18780 (N_18780,N_18189,N_18358);
nor U18781 (N_18781,N_18412,N_18435);
or U18782 (N_18782,N_18209,N_18235);
nand U18783 (N_18783,N_18067,N_18353);
nand U18784 (N_18784,N_18190,N_18206);
or U18785 (N_18785,N_18296,N_18161);
nand U18786 (N_18786,N_18076,N_18048);
or U18787 (N_18787,N_18459,N_18373);
and U18788 (N_18788,N_18122,N_18162);
and U18789 (N_18789,N_18074,N_18313);
nor U18790 (N_18790,N_18299,N_18443);
nor U18791 (N_18791,N_18475,N_18233);
nand U18792 (N_18792,N_18426,N_18133);
or U18793 (N_18793,N_18207,N_18049);
and U18794 (N_18794,N_18274,N_18168);
nand U18795 (N_18795,N_18359,N_18434);
nor U18796 (N_18796,N_18328,N_18413);
nand U18797 (N_18797,N_18221,N_18172);
and U18798 (N_18798,N_18263,N_18393);
or U18799 (N_18799,N_18326,N_18358);
or U18800 (N_18800,N_18092,N_18104);
and U18801 (N_18801,N_18177,N_18339);
nor U18802 (N_18802,N_18324,N_18213);
nor U18803 (N_18803,N_18341,N_18027);
and U18804 (N_18804,N_18167,N_18036);
nand U18805 (N_18805,N_18388,N_18081);
or U18806 (N_18806,N_18194,N_18478);
and U18807 (N_18807,N_18410,N_18285);
or U18808 (N_18808,N_18015,N_18103);
or U18809 (N_18809,N_18460,N_18410);
and U18810 (N_18810,N_18345,N_18031);
nor U18811 (N_18811,N_18148,N_18211);
or U18812 (N_18812,N_18301,N_18199);
nand U18813 (N_18813,N_18273,N_18279);
nor U18814 (N_18814,N_18244,N_18474);
nand U18815 (N_18815,N_18142,N_18035);
nand U18816 (N_18816,N_18427,N_18095);
and U18817 (N_18817,N_18199,N_18082);
and U18818 (N_18818,N_18126,N_18401);
and U18819 (N_18819,N_18469,N_18328);
or U18820 (N_18820,N_18074,N_18480);
nor U18821 (N_18821,N_18386,N_18429);
and U18822 (N_18822,N_18333,N_18122);
nor U18823 (N_18823,N_18153,N_18181);
and U18824 (N_18824,N_18065,N_18431);
nor U18825 (N_18825,N_18411,N_18014);
and U18826 (N_18826,N_18194,N_18263);
and U18827 (N_18827,N_18074,N_18136);
nor U18828 (N_18828,N_18490,N_18208);
nor U18829 (N_18829,N_18003,N_18404);
or U18830 (N_18830,N_18187,N_18418);
nand U18831 (N_18831,N_18154,N_18133);
nor U18832 (N_18832,N_18040,N_18344);
nand U18833 (N_18833,N_18113,N_18330);
and U18834 (N_18834,N_18064,N_18243);
nand U18835 (N_18835,N_18057,N_18229);
nor U18836 (N_18836,N_18291,N_18033);
nand U18837 (N_18837,N_18498,N_18046);
or U18838 (N_18838,N_18033,N_18230);
xnor U18839 (N_18839,N_18485,N_18043);
and U18840 (N_18840,N_18471,N_18008);
and U18841 (N_18841,N_18140,N_18279);
or U18842 (N_18842,N_18330,N_18048);
nor U18843 (N_18843,N_18082,N_18209);
and U18844 (N_18844,N_18341,N_18090);
nor U18845 (N_18845,N_18358,N_18280);
nor U18846 (N_18846,N_18231,N_18086);
nor U18847 (N_18847,N_18469,N_18249);
nor U18848 (N_18848,N_18228,N_18081);
or U18849 (N_18849,N_18208,N_18292);
nor U18850 (N_18850,N_18072,N_18153);
nand U18851 (N_18851,N_18045,N_18153);
or U18852 (N_18852,N_18450,N_18361);
nor U18853 (N_18853,N_18457,N_18475);
nand U18854 (N_18854,N_18226,N_18423);
and U18855 (N_18855,N_18141,N_18136);
nand U18856 (N_18856,N_18487,N_18208);
and U18857 (N_18857,N_18271,N_18083);
nor U18858 (N_18858,N_18334,N_18381);
nand U18859 (N_18859,N_18368,N_18182);
nor U18860 (N_18860,N_18367,N_18494);
and U18861 (N_18861,N_18016,N_18472);
nor U18862 (N_18862,N_18465,N_18341);
or U18863 (N_18863,N_18161,N_18368);
nor U18864 (N_18864,N_18255,N_18356);
or U18865 (N_18865,N_18428,N_18482);
or U18866 (N_18866,N_18039,N_18193);
nor U18867 (N_18867,N_18260,N_18283);
nand U18868 (N_18868,N_18020,N_18246);
nand U18869 (N_18869,N_18309,N_18394);
nand U18870 (N_18870,N_18274,N_18130);
nor U18871 (N_18871,N_18410,N_18060);
nor U18872 (N_18872,N_18280,N_18092);
or U18873 (N_18873,N_18121,N_18049);
and U18874 (N_18874,N_18110,N_18255);
or U18875 (N_18875,N_18495,N_18490);
or U18876 (N_18876,N_18050,N_18382);
nor U18877 (N_18877,N_18489,N_18261);
or U18878 (N_18878,N_18420,N_18349);
nor U18879 (N_18879,N_18341,N_18227);
and U18880 (N_18880,N_18136,N_18383);
nand U18881 (N_18881,N_18013,N_18046);
or U18882 (N_18882,N_18285,N_18044);
nand U18883 (N_18883,N_18442,N_18020);
or U18884 (N_18884,N_18101,N_18117);
nand U18885 (N_18885,N_18352,N_18129);
nand U18886 (N_18886,N_18218,N_18350);
nand U18887 (N_18887,N_18467,N_18336);
and U18888 (N_18888,N_18410,N_18288);
or U18889 (N_18889,N_18399,N_18347);
nand U18890 (N_18890,N_18200,N_18486);
and U18891 (N_18891,N_18349,N_18158);
nand U18892 (N_18892,N_18472,N_18336);
nand U18893 (N_18893,N_18029,N_18138);
or U18894 (N_18894,N_18001,N_18401);
and U18895 (N_18895,N_18336,N_18137);
nand U18896 (N_18896,N_18267,N_18408);
nor U18897 (N_18897,N_18132,N_18354);
and U18898 (N_18898,N_18296,N_18046);
nand U18899 (N_18899,N_18316,N_18489);
or U18900 (N_18900,N_18441,N_18276);
or U18901 (N_18901,N_18143,N_18057);
nor U18902 (N_18902,N_18438,N_18180);
and U18903 (N_18903,N_18335,N_18407);
or U18904 (N_18904,N_18113,N_18249);
or U18905 (N_18905,N_18114,N_18237);
nand U18906 (N_18906,N_18016,N_18161);
and U18907 (N_18907,N_18376,N_18223);
nor U18908 (N_18908,N_18410,N_18491);
nor U18909 (N_18909,N_18465,N_18163);
or U18910 (N_18910,N_18126,N_18375);
or U18911 (N_18911,N_18001,N_18260);
or U18912 (N_18912,N_18036,N_18070);
nand U18913 (N_18913,N_18275,N_18289);
or U18914 (N_18914,N_18326,N_18327);
and U18915 (N_18915,N_18094,N_18329);
nor U18916 (N_18916,N_18436,N_18301);
nand U18917 (N_18917,N_18067,N_18362);
nor U18918 (N_18918,N_18485,N_18151);
and U18919 (N_18919,N_18113,N_18079);
nand U18920 (N_18920,N_18391,N_18198);
and U18921 (N_18921,N_18027,N_18268);
nor U18922 (N_18922,N_18396,N_18229);
or U18923 (N_18923,N_18005,N_18373);
nor U18924 (N_18924,N_18315,N_18355);
or U18925 (N_18925,N_18011,N_18222);
nand U18926 (N_18926,N_18423,N_18305);
nand U18927 (N_18927,N_18099,N_18399);
nand U18928 (N_18928,N_18010,N_18197);
nand U18929 (N_18929,N_18223,N_18452);
and U18930 (N_18930,N_18451,N_18167);
nor U18931 (N_18931,N_18337,N_18429);
nand U18932 (N_18932,N_18009,N_18449);
nor U18933 (N_18933,N_18297,N_18058);
nand U18934 (N_18934,N_18012,N_18103);
and U18935 (N_18935,N_18269,N_18134);
or U18936 (N_18936,N_18342,N_18042);
nand U18937 (N_18937,N_18071,N_18427);
or U18938 (N_18938,N_18218,N_18017);
or U18939 (N_18939,N_18350,N_18137);
or U18940 (N_18940,N_18241,N_18162);
nand U18941 (N_18941,N_18174,N_18344);
or U18942 (N_18942,N_18183,N_18177);
nand U18943 (N_18943,N_18283,N_18424);
or U18944 (N_18944,N_18279,N_18492);
or U18945 (N_18945,N_18162,N_18385);
nor U18946 (N_18946,N_18029,N_18283);
nand U18947 (N_18947,N_18001,N_18147);
and U18948 (N_18948,N_18400,N_18173);
nand U18949 (N_18949,N_18195,N_18361);
or U18950 (N_18950,N_18415,N_18162);
nor U18951 (N_18951,N_18191,N_18396);
or U18952 (N_18952,N_18457,N_18255);
nor U18953 (N_18953,N_18178,N_18118);
nand U18954 (N_18954,N_18422,N_18437);
and U18955 (N_18955,N_18224,N_18118);
nand U18956 (N_18956,N_18267,N_18406);
nor U18957 (N_18957,N_18021,N_18367);
or U18958 (N_18958,N_18030,N_18414);
nand U18959 (N_18959,N_18100,N_18486);
and U18960 (N_18960,N_18416,N_18482);
nor U18961 (N_18961,N_18464,N_18350);
xnor U18962 (N_18962,N_18024,N_18221);
or U18963 (N_18963,N_18217,N_18371);
nand U18964 (N_18964,N_18161,N_18427);
and U18965 (N_18965,N_18265,N_18122);
or U18966 (N_18966,N_18268,N_18067);
or U18967 (N_18967,N_18275,N_18081);
nor U18968 (N_18968,N_18261,N_18072);
or U18969 (N_18969,N_18109,N_18132);
and U18970 (N_18970,N_18461,N_18073);
nand U18971 (N_18971,N_18323,N_18012);
and U18972 (N_18972,N_18229,N_18197);
nor U18973 (N_18973,N_18294,N_18158);
or U18974 (N_18974,N_18004,N_18265);
and U18975 (N_18975,N_18124,N_18448);
nor U18976 (N_18976,N_18411,N_18179);
xor U18977 (N_18977,N_18490,N_18029);
nor U18978 (N_18978,N_18083,N_18037);
nand U18979 (N_18979,N_18360,N_18090);
nand U18980 (N_18980,N_18223,N_18144);
and U18981 (N_18981,N_18291,N_18116);
or U18982 (N_18982,N_18260,N_18341);
or U18983 (N_18983,N_18436,N_18404);
and U18984 (N_18984,N_18478,N_18022);
and U18985 (N_18985,N_18453,N_18432);
nand U18986 (N_18986,N_18010,N_18009);
nand U18987 (N_18987,N_18025,N_18296);
or U18988 (N_18988,N_18320,N_18440);
or U18989 (N_18989,N_18403,N_18166);
and U18990 (N_18990,N_18110,N_18385);
or U18991 (N_18991,N_18405,N_18309);
nor U18992 (N_18992,N_18288,N_18394);
nand U18993 (N_18993,N_18468,N_18378);
and U18994 (N_18994,N_18212,N_18379);
nand U18995 (N_18995,N_18037,N_18286);
nor U18996 (N_18996,N_18212,N_18062);
nand U18997 (N_18997,N_18275,N_18460);
or U18998 (N_18998,N_18360,N_18475);
and U18999 (N_18999,N_18017,N_18317);
nand U19000 (N_19000,N_18837,N_18741);
or U19001 (N_19001,N_18593,N_18824);
nand U19002 (N_19002,N_18768,N_18610);
nor U19003 (N_19003,N_18985,N_18885);
nor U19004 (N_19004,N_18980,N_18952);
or U19005 (N_19005,N_18806,N_18523);
nor U19006 (N_19006,N_18779,N_18875);
or U19007 (N_19007,N_18692,N_18799);
nand U19008 (N_19008,N_18962,N_18902);
nand U19009 (N_19009,N_18889,N_18819);
nor U19010 (N_19010,N_18918,N_18625);
or U19011 (N_19011,N_18677,N_18746);
nand U19012 (N_19012,N_18512,N_18560);
and U19013 (N_19013,N_18568,N_18800);
and U19014 (N_19014,N_18955,N_18898);
and U19015 (N_19015,N_18706,N_18878);
and U19016 (N_19016,N_18825,N_18522);
nand U19017 (N_19017,N_18872,N_18859);
or U19018 (N_19018,N_18906,N_18785);
and U19019 (N_19019,N_18589,N_18650);
and U19020 (N_19020,N_18782,N_18506);
and U19021 (N_19021,N_18660,N_18618);
nand U19022 (N_19022,N_18971,N_18763);
nor U19023 (N_19023,N_18626,N_18826);
nor U19024 (N_19024,N_18754,N_18731);
nand U19025 (N_19025,N_18551,N_18659);
and U19026 (N_19026,N_18707,N_18877);
nand U19027 (N_19027,N_18930,N_18944);
and U19028 (N_19028,N_18655,N_18682);
and U19029 (N_19029,N_18748,N_18908);
or U19030 (N_19030,N_18718,N_18844);
nor U19031 (N_19031,N_18616,N_18515);
nor U19032 (N_19032,N_18619,N_18788);
nand U19033 (N_19033,N_18776,N_18901);
nand U19034 (N_19034,N_18835,N_18862);
and U19035 (N_19035,N_18828,N_18654);
nand U19036 (N_19036,N_18674,N_18578);
and U19037 (N_19037,N_18967,N_18668);
nand U19038 (N_19038,N_18595,N_18511);
and U19039 (N_19039,N_18897,N_18698);
nor U19040 (N_19040,N_18851,N_18533);
and U19041 (N_19041,N_18501,N_18950);
and U19042 (N_19042,N_18689,N_18599);
or U19043 (N_19043,N_18998,N_18888);
or U19044 (N_19044,N_18993,N_18608);
and U19045 (N_19045,N_18657,N_18986);
nor U19046 (N_19046,N_18874,N_18700);
and U19047 (N_19047,N_18678,N_18594);
nand U19048 (N_19048,N_18588,N_18663);
nor U19049 (N_19049,N_18792,N_18848);
or U19050 (N_19050,N_18736,N_18892);
and U19051 (N_19051,N_18548,N_18696);
or U19052 (N_19052,N_18658,N_18643);
and U19053 (N_19053,N_18507,N_18920);
nor U19054 (N_19054,N_18517,N_18852);
or U19055 (N_19055,N_18840,N_18894);
and U19056 (N_19056,N_18518,N_18752);
or U19057 (N_19057,N_18639,N_18559);
and U19058 (N_19058,N_18742,N_18747);
and U19059 (N_19059,N_18795,N_18831);
nand U19060 (N_19060,N_18635,N_18703);
nor U19061 (N_19061,N_18645,N_18863);
nand U19062 (N_19062,N_18673,N_18529);
or U19063 (N_19063,N_18600,N_18603);
or U19064 (N_19064,N_18953,N_18652);
nor U19065 (N_19065,N_18966,N_18999);
or U19066 (N_19066,N_18509,N_18605);
nand U19067 (N_19067,N_18900,N_18526);
and U19068 (N_19068,N_18803,N_18520);
or U19069 (N_19069,N_18869,N_18991);
nand U19070 (N_19070,N_18676,N_18644);
nand U19071 (N_19071,N_18646,N_18536);
nand U19072 (N_19072,N_18883,N_18500);
nand U19073 (N_19073,N_18917,N_18726);
nand U19074 (N_19074,N_18807,N_18813);
nor U19075 (N_19075,N_18601,N_18974);
or U19076 (N_19076,N_18850,N_18777);
nor U19077 (N_19077,N_18789,N_18633);
and U19078 (N_19078,N_18946,N_18717);
nand U19079 (N_19079,N_18879,N_18954);
nor U19080 (N_19080,N_18973,N_18784);
nor U19081 (N_19081,N_18948,N_18994);
nand U19082 (N_19082,N_18691,N_18925);
nor U19083 (N_19083,N_18503,N_18729);
nand U19084 (N_19084,N_18539,N_18627);
and U19085 (N_19085,N_18933,N_18727);
nor U19086 (N_19086,N_18725,N_18555);
or U19087 (N_19087,N_18535,N_18912);
or U19088 (N_19088,N_18904,N_18730);
and U19089 (N_19089,N_18921,N_18550);
and U19090 (N_19090,N_18662,N_18783);
nor U19091 (N_19091,N_18801,N_18505);
and U19092 (N_19092,N_18915,N_18680);
or U19093 (N_19093,N_18567,N_18965);
and U19094 (N_19094,N_18981,N_18577);
and U19095 (N_19095,N_18956,N_18584);
nand U19096 (N_19096,N_18556,N_18797);
and U19097 (N_19097,N_18716,N_18670);
nor U19098 (N_19098,N_18563,N_18988);
nand U19099 (N_19099,N_18821,N_18721);
nand U19100 (N_19100,N_18934,N_18990);
or U19101 (N_19101,N_18531,N_18870);
nand U19102 (N_19102,N_18834,N_18695);
nor U19103 (N_19103,N_18764,N_18972);
nor U19104 (N_19104,N_18951,N_18534);
or U19105 (N_19105,N_18771,N_18665);
nor U19106 (N_19106,N_18832,N_18775);
nand U19107 (N_19107,N_18949,N_18566);
nor U19108 (N_19108,N_18936,N_18621);
nor U19109 (N_19109,N_18823,N_18611);
nor U19110 (N_19110,N_18569,N_18984);
nand U19111 (N_19111,N_18576,N_18694);
and U19112 (N_19112,N_18675,N_18932);
and U19113 (N_19113,N_18562,N_18739);
nor U19114 (N_19114,N_18620,N_18581);
or U19115 (N_19115,N_18854,N_18519);
and U19116 (N_19116,N_18609,N_18772);
or U19117 (N_19117,N_18672,N_18697);
and U19118 (N_19118,N_18637,N_18818);
and U19119 (N_19119,N_18558,N_18614);
or U19120 (N_19120,N_18532,N_18570);
nor U19121 (N_19121,N_18749,N_18711);
and U19122 (N_19122,N_18745,N_18853);
or U19123 (N_19123,N_18709,N_18669);
and U19124 (N_19124,N_18798,N_18910);
and U19125 (N_19125,N_18929,N_18762);
and U19126 (N_19126,N_18592,N_18649);
and U19127 (N_19127,N_18805,N_18615);
nand U19128 (N_19128,N_18767,N_18829);
nor U19129 (N_19129,N_18597,N_18671);
nand U19130 (N_19130,N_18634,N_18638);
and U19131 (N_19131,N_18759,N_18893);
nor U19132 (N_19132,N_18540,N_18722);
and U19133 (N_19133,N_18681,N_18564);
and U19134 (N_19134,N_18849,N_18876);
nor U19135 (N_19135,N_18856,N_18873);
nor U19136 (N_19136,N_18867,N_18773);
and U19137 (N_19137,N_18565,N_18541);
nor U19138 (N_19138,N_18891,N_18780);
nand U19139 (N_19139,N_18791,N_18508);
nor U19140 (N_19140,N_18648,N_18911);
and U19141 (N_19141,N_18757,N_18743);
or U19142 (N_19142,N_18820,N_18702);
and U19143 (N_19143,N_18774,N_18604);
and U19144 (N_19144,N_18552,N_18733);
nand U19145 (N_19145,N_18723,N_18842);
or U19146 (N_19146,N_18941,N_18781);
or U19147 (N_19147,N_18896,N_18712);
and U19148 (N_19148,N_18557,N_18661);
or U19149 (N_19149,N_18710,N_18542);
nand U19150 (N_19150,N_18909,N_18907);
and U19151 (N_19151,N_18547,N_18579);
nor U19152 (N_19152,N_18786,N_18963);
nor U19153 (N_19153,N_18744,N_18945);
nand U19154 (N_19154,N_18886,N_18613);
or U19155 (N_19155,N_18684,N_18631);
or U19156 (N_19156,N_18755,N_18530);
and U19157 (N_19157,N_18513,N_18868);
nor U19158 (N_19158,N_18760,N_18811);
nor U19159 (N_19159,N_18571,N_18651);
or U19160 (N_19160,N_18528,N_18705);
nor U19161 (N_19161,N_18628,N_18935);
nor U19162 (N_19162,N_18516,N_18766);
and U19163 (N_19163,N_18502,N_18838);
and U19164 (N_19164,N_18793,N_18575);
nor U19165 (N_19165,N_18719,N_18815);
or U19166 (N_19166,N_18860,N_18734);
or U19167 (N_19167,N_18514,N_18942);
nand U19168 (N_19168,N_18688,N_18855);
xnor U19169 (N_19169,N_18622,N_18940);
nand U19170 (N_19170,N_18997,N_18939);
or U19171 (N_19171,N_18943,N_18538);
nand U19172 (N_19172,N_18927,N_18740);
or U19173 (N_19173,N_18713,N_18687);
and U19174 (N_19174,N_18959,N_18561);
nor U19175 (N_19175,N_18960,N_18794);
nor U19176 (N_19176,N_18602,N_18970);
and U19177 (N_19177,N_18871,N_18735);
and U19178 (N_19178,N_18632,N_18732);
and U19179 (N_19179,N_18667,N_18903);
nand U19180 (N_19180,N_18653,N_18841);
or U19181 (N_19181,N_18814,N_18865);
nor U19182 (N_19182,N_18715,N_18937);
nand U19183 (N_19183,N_18699,N_18720);
or U19184 (N_19184,N_18510,N_18881);
or U19185 (N_19185,N_18574,N_18996);
or U19186 (N_19186,N_18708,N_18630);
nand U19187 (N_19187,N_18938,N_18612);
and U19188 (N_19188,N_18679,N_18714);
or U19189 (N_19189,N_18922,N_18812);
or U19190 (N_19190,N_18968,N_18787);
and U19191 (N_19191,N_18958,N_18525);
and U19192 (N_19192,N_18836,N_18761);
nor U19193 (N_19193,N_18884,N_18847);
or U19194 (N_19194,N_18987,N_18690);
nor U19195 (N_19195,N_18737,N_18923);
nor U19196 (N_19196,N_18899,N_18586);
or U19197 (N_19197,N_18753,N_18802);
nor U19198 (N_19198,N_18890,N_18913);
nand U19199 (N_19199,N_18804,N_18857);
or U19200 (N_19200,N_18641,N_18977);
nand U19201 (N_19201,N_18724,N_18607);
and U19202 (N_19202,N_18833,N_18827);
and U19203 (N_19203,N_18765,N_18664);
nand U19204 (N_19204,N_18979,N_18553);
nor U19205 (N_19205,N_18957,N_18978);
or U19206 (N_19206,N_18926,N_18524);
nand U19207 (N_19207,N_18549,N_18982);
nand U19208 (N_19208,N_18598,N_18527);
or U19209 (N_19209,N_18861,N_18629);
nand U19210 (N_19210,N_18931,N_18636);
nand U19211 (N_19211,N_18537,N_18544);
and U19212 (N_19212,N_18858,N_18769);
nand U19213 (N_19213,N_18573,N_18642);
xor U19214 (N_19214,N_18983,N_18961);
nor U19215 (N_19215,N_18572,N_18623);
or U19216 (N_19216,N_18882,N_18656);
and U19217 (N_19217,N_18686,N_18704);
nand U19218 (N_19218,N_18590,N_18947);
and U19219 (N_19219,N_18790,N_18624);
nor U19220 (N_19220,N_18816,N_18756);
and U19221 (N_19221,N_18866,N_18845);
nand U19222 (N_19222,N_18864,N_18683);
or U19223 (N_19223,N_18685,N_18969);
or U19224 (N_19224,N_18647,N_18606);
nand U19225 (N_19225,N_18617,N_18596);
and U19226 (N_19226,N_18914,N_18543);
or U19227 (N_19227,N_18905,N_18810);
nor U19228 (N_19228,N_18701,N_18995);
nor U19229 (N_19229,N_18770,N_18846);
nand U19230 (N_19230,N_18554,N_18591);
and U19231 (N_19231,N_18546,N_18976);
and U19232 (N_19232,N_18693,N_18587);
nand U19233 (N_19233,N_18640,N_18817);
nand U19234 (N_19234,N_18989,N_18796);
nor U19235 (N_19235,N_18887,N_18808);
and U19236 (N_19236,N_18880,N_18822);
nand U19237 (N_19237,N_18521,N_18964);
nor U19238 (N_19238,N_18585,N_18928);
nand U19239 (N_19239,N_18582,N_18738);
nand U19240 (N_19240,N_18839,N_18751);
and U19241 (N_19241,N_18583,N_18545);
nand U19242 (N_19242,N_18843,N_18580);
nor U19243 (N_19243,N_18830,N_18750);
and U19244 (N_19244,N_18504,N_18916);
nand U19245 (N_19245,N_18728,N_18758);
or U19246 (N_19246,N_18895,N_18992);
nand U19247 (N_19247,N_18975,N_18924);
or U19248 (N_19248,N_18919,N_18666);
nor U19249 (N_19249,N_18778,N_18809);
nand U19250 (N_19250,N_18750,N_18573);
nand U19251 (N_19251,N_18815,N_18936);
nand U19252 (N_19252,N_18697,N_18743);
or U19253 (N_19253,N_18715,N_18941);
nor U19254 (N_19254,N_18669,N_18694);
nor U19255 (N_19255,N_18998,N_18982);
nor U19256 (N_19256,N_18605,N_18975);
nand U19257 (N_19257,N_18522,N_18818);
or U19258 (N_19258,N_18892,N_18867);
nor U19259 (N_19259,N_18550,N_18696);
and U19260 (N_19260,N_18589,N_18696);
and U19261 (N_19261,N_18942,N_18579);
or U19262 (N_19262,N_18542,N_18649);
nor U19263 (N_19263,N_18629,N_18806);
nor U19264 (N_19264,N_18779,N_18673);
nand U19265 (N_19265,N_18820,N_18794);
nor U19266 (N_19266,N_18795,N_18754);
and U19267 (N_19267,N_18616,N_18567);
or U19268 (N_19268,N_18605,N_18690);
and U19269 (N_19269,N_18747,N_18513);
nand U19270 (N_19270,N_18728,N_18801);
and U19271 (N_19271,N_18626,N_18859);
or U19272 (N_19272,N_18629,N_18976);
and U19273 (N_19273,N_18500,N_18748);
and U19274 (N_19274,N_18715,N_18988);
or U19275 (N_19275,N_18628,N_18978);
nor U19276 (N_19276,N_18916,N_18590);
or U19277 (N_19277,N_18794,N_18562);
nand U19278 (N_19278,N_18815,N_18766);
nand U19279 (N_19279,N_18853,N_18957);
and U19280 (N_19280,N_18509,N_18982);
nand U19281 (N_19281,N_18870,N_18656);
or U19282 (N_19282,N_18887,N_18782);
nand U19283 (N_19283,N_18942,N_18886);
or U19284 (N_19284,N_18896,N_18790);
nor U19285 (N_19285,N_18840,N_18794);
or U19286 (N_19286,N_18907,N_18866);
and U19287 (N_19287,N_18885,N_18698);
and U19288 (N_19288,N_18997,N_18602);
nor U19289 (N_19289,N_18578,N_18623);
nor U19290 (N_19290,N_18816,N_18598);
and U19291 (N_19291,N_18886,N_18808);
nand U19292 (N_19292,N_18656,N_18680);
nor U19293 (N_19293,N_18553,N_18703);
nand U19294 (N_19294,N_18679,N_18525);
and U19295 (N_19295,N_18847,N_18976);
and U19296 (N_19296,N_18563,N_18667);
nor U19297 (N_19297,N_18864,N_18657);
nand U19298 (N_19298,N_18825,N_18778);
and U19299 (N_19299,N_18557,N_18703);
and U19300 (N_19300,N_18735,N_18878);
or U19301 (N_19301,N_18947,N_18555);
and U19302 (N_19302,N_18725,N_18661);
nand U19303 (N_19303,N_18725,N_18592);
nor U19304 (N_19304,N_18707,N_18760);
nor U19305 (N_19305,N_18982,N_18686);
nand U19306 (N_19306,N_18913,N_18807);
nand U19307 (N_19307,N_18762,N_18866);
nor U19308 (N_19308,N_18923,N_18604);
or U19309 (N_19309,N_18552,N_18526);
xor U19310 (N_19310,N_18613,N_18753);
and U19311 (N_19311,N_18606,N_18652);
or U19312 (N_19312,N_18835,N_18698);
nor U19313 (N_19313,N_18544,N_18509);
or U19314 (N_19314,N_18618,N_18824);
and U19315 (N_19315,N_18754,N_18593);
nand U19316 (N_19316,N_18660,N_18762);
xor U19317 (N_19317,N_18514,N_18818);
nor U19318 (N_19318,N_18858,N_18608);
and U19319 (N_19319,N_18615,N_18870);
nor U19320 (N_19320,N_18975,N_18529);
nor U19321 (N_19321,N_18640,N_18720);
nand U19322 (N_19322,N_18648,N_18925);
nor U19323 (N_19323,N_18906,N_18952);
or U19324 (N_19324,N_18622,N_18883);
nor U19325 (N_19325,N_18886,N_18911);
or U19326 (N_19326,N_18587,N_18766);
or U19327 (N_19327,N_18870,N_18970);
nand U19328 (N_19328,N_18738,N_18956);
and U19329 (N_19329,N_18665,N_18838);
nand U19330 (N_19330,N_18920,N_18547);
or U19331 (N_19331,N_18877,N_18632);
or U19332 (N_19332,N_18872,N_18605);
nand U19333 (N_19333,N_18549,N_18706);
nor U19334 (N_19334,N_18581,N_18653);
nor U19335 (N_19335,N_18897,N_18564);
and U19336 (N_19336,N_18860,N_18924);
nor U19337 (N_19337,N_18756,N_18586);
nor U19338 (N_19338,N_18863,N_18935);
nor U19339 (N_19339,N_18587,N_18785);
and U19340 (N_19340,N_18948,N_18810);
or U19341 (N_19341,N_18608,N_18701);
nand U19342 (N_19342,N_18505,N_18770);
nor U19343 (N_19343,N_18767,N_18866);
or U19344 (N_19344,N_18662,N_18848);
nor U19345 (N_19345,N_18960,N_18764);
nand U19346 (N_19346,N_18925,N_18708);
nand U19347 (N_19347,N_18905,N_18504);
nor U19348 (N_19348,N_18855,N_18860);
nand U19349 (N_19349,N_18544,N_18999);
nor U19350 (N_19350,N_18987,N_18600);
nor U19351 (N_19351,N_18807,N_18758);
or U19352 (N_19352,N_18516,N_18638);
or U19353 (N_19353,N_18894,N_18834);
and U19354 (N_19354,N_18563,N_18782);
nor U19355 (N_19355,N_18609,N_18935);
and U19356 (N_19356,N_18635,N_18653);
or U19357 (N_19357,N_18773,N_18624);
nand U19358 (N_19358,N_18908,N_18872);
and U19359 (N_19359,N_18708,N_18818);
nand U19360 (N_19360,N_18586,N_18975);
nand U19361 (N_19361,N_18937,N_18706);
xnor U19362 (N_19362,N_18658,N_18976);
nand U19363 (N_19363,N_18611,N_18899);
nor U19364 (N_19364,N_18611,N_18561);
and U19365 (N_19365,N_18545,N_18700);
or U19366 (N_19366,N_18964,N_18998);
nor U19367 (N_19367,N_18585,N_18973);
nor U19368 (N_19368,N_18698,N_18872);
nand U19369 (N_19369,N_18638,N_18580);
nand U19370 (N_19370,N_18883,N_18954);
and U19371 (N_19371,N_18949,N_18587);
nor U19372 (N_19372,N_18973,N_18940);
nor U19373 (N_19373,N_18504,N_18908);
nor U19374 (N_19374,N_18658,N_18959);
or U19375 (N_19375,N_18751,N_18976);
or U19376 (N_19376,N_18571,N_18508);
nor U19377 (N_19377,N_18521,N_18992);
or U19378 (N_19378,N_18740,N_18921);
nand U19379 (N_19379,N_18873,N_18902);
nor U19380 (N_19380,N_18943,N_18523);
nand U19381 (N_19381,N_18940,N_18627);
and U19382 (N_19382,N_18684,N_18660);
or U19383 (N_19383,N_18577,N_18629);
nand U19384 (N_19384,N_18742,N_18736);
nand U19385 (N_19385,N_18522,N_18504);
nand U19386 (N_19386,N_18902,N_18679);
and U19387 (N_19387,N_18777,N_18731);
and U19388 (N_19388,N_18761,N_18772);
or U19389 (N_19389,N_18574,N_18609);
and U19390 (N_19390,N_18922,N_18880);
nor U19391 (N_19391,N_18705,N_18887);
nor U19392 (N_19392,N_18791,N_18606);
nor U19393 (N_19393,N_18931,N_18587);
nor U19394 (N_19394,N_18501,N_18629);
or U19395 (N_19395,N_18991,N_18768);
nor U19396 (N_19396,N_18714,N_18988);
and U19397 (N_19397,N_18738,N_18860);
nand U19398 (N_19398,N_18745,N_18657);
or U19399 (N_19399,N_18976,N_18720);
and U19400 (N_19400,N_18738,N_18880);
or U19401 (N_19401,N_18862,N_18564);
nand U19402 (N_19402,N_18868,N_18947);
nor U19403 (N_19403,N_18703,N_18632);
nor U19404 (N_19404,N_18881,N_18755);
nand U19405 (N_19405,N_18521,N_18666);
nor U19406 (N_19406,N_18977,N_18994);
or U19407 (N_19407,N_18854,N_18627);
nand U19408 (N_19408,N_18543,N_18659);
or U19409 (N_19409,N_18945,N_18502);
nand U19410 (N_19410,N_18634,N_18981);
or U19411 (N_19411,N_18923,N_18516);
xnor U19412 (N_19412,N_18617,N_18857);
or U19413 (N_19413,N_18890,N_18500);
nor U19414 (N_19414,N_18993,N_18525);
nand U19415 (N_19415,N_18562,N_18812);
nand U19416 (N_19416,N_18777,N_18970);
nor U19417 (N_19417,N_18650,N_18510);
nor U19418 (N_19418,N_18615,N_18741);
and U19419 (N_19419,N_18841,N_18502);
nor U19420 (N_19420,N_18945,N_18875);
and U19421 (N_19421,N_18912,N_18711);
and U19422 (N_19422,N_18874,N_18866);
and U19423 (N_19423,N_18896,N_18584);
nand U19424 (N_19424,N_18557,N_18970);
nand U19425 (N_19425,N_18757,N_18656);
or U19426 (N_19426,N_18840,N_18855);
nand U19427 (N_19427,N_18779,N_18954);
nand U19428 (N_19428,N_18887,N_18687);
and U19429 (N_19429,N_18667,N_18940);
or U19430 (N_19430,N_18666,N_18938);
nor U19431 (N_19431,N_18681,N_18934);
nand U19432 (N_19432,N_18908,N_18554);
nor U19433 (N_19433,N_18521,N_18888);
nor U19434 (N_19434,N_18608,N_18759);
or U19435 (N_19435,N_18934,N_18861);
and U19436 (N_19436,N_18804,N_18991);
nand U19437 (N_19437,N_18734,N_18926);
or U19438 (N_19438,N_18939,N_18728);
nand U19439 (N_19439,N_18513,N_18849);
nor U19440 (N_19440,N_18713,N_18810);
nor U19441 (N_19441,N_18803,N_18804);
or U19442 (N_19442,N_18825,N_18794);
nor U19443 (N_19443,N_18570,N_18908);
nor U19444 (N_19444,N_18636,N_18938);
nor U19445 (N_19445,N_18993,N_18598);
nor U19446 (N_19446,N_18994,N_18574);
and U19447 (N_19447,N_18738,N_18516);
or U19448 (N_19448,N_18769,N_18591);
or U19449 (N_19449,N_18962,N_18630);
nor U19450 (N_19450,N_18775,N_18774);
nand U19451 (N_19451,N_18947,N_18886);
and U19452 (N_19452,N_18790,N_18591);
and U19453 (N_19453,N_18607,N_18572);
or U19454 (N_19454,N_18832,N_18890);
nor U19455 (N_19455,N_18647,N_18899);
nor U19456 (N_19456,N_18650,N_18579);
and U19457 (N_19457,N_18572,N_18554);
nand U19458 (N_19458,N_18571,N_18533);
nand U19459 (N_19459,N_18543,N_18921);
nor U19460 (N_19460,N_18539,N_18745);
and U19461 (N_19461,N_18887,N_18682);
and U19462 (N_19462,N_18704,N_18743);
and U19463 (N_19463,N_18889,N_18771);
and U19464 (N_19464,N_18755,N_18611);
nor U19465 (N_19465,N_18958,N_18774);
nor U19466 (N_19466,N_18511,N_18577);
or U19467 (N_19467,N_18596,N_18972);
or U19468 (N_19468,N_18602,N_18914);
or U19469 (N_19469,N_18650,N_18776);
nor U19470 (N_19470,N_18798,N_18616);
or U19471 (N_19471,N_18795,N_18950);
nand U19472 (N_19472,N_18748,N_18879);
nand U19473 (N_19473,N_18805,N_18656);
nor U19474 (N_19474,N_18557,N_18629);
and U19475 (N_19475,N_18843,N_18533);
nand U19476 (N_19476,N_18792,N_18717);
nor U19477 (N_19477,N_18847,N_18556);
and U19478 (N_19478,N_18735,N_18812);
and U19479 (N_19479,N_18510,N_18515);
nand U19480 (N_19480,N_18575,N_18523);
nor U19481 (N_19481,N_18800,N_18910);
and U19482 (N_19482,N_18684,N_18625);
nand U19483 (N_19483,N_18563,N_18949);
nor U19484 (N_19484,N_18857,N_18551);
nor U19485 (N_19485,N_18656,N_18537);
nor U19486 (N_19486,N_18736,N_18739);
and U19487 (N_19487,N_18973,N_18689);
nor U19488 (N_19488,N_18546,N_18924);
or U19489 (N_19489,N_18922,N_18902);
nor U19490 (N_19490,N_18831,N_18739);
and U19491 (N_19491,N_18540,N_18766);
xnor U19492 (N_19492,N_18592,N_18682);
or U19493 (N_19493,N_18799,N_18632);
nand U19494 (N_19494,N_18853,N_18935);
nor U19495 (N_19495,N_18924,N_18931);
nand U19496 (N_19496,N_18623,N_18978);
nor U19497 (N_19497,N_18912,N_18956);
and U19498 (N_19498,N_18570,N_18747);
nor U19499 (N_19499,N_18713,N_18997);
or U19500 (N_19500,N_19001,N_19318);
nor U19501 (N_19501,N_19340,N_19078);
and U19502 (N_19502,N_19122,N_19240);
nand U19503 (N_19503,N_19155,N_19499);
or U19504 (N_19504,N_19422,N_19171);
and U19505 (N_19505,N_19326,N_19428);
nor U19506 (N_19506,N_19012,N_19113);
and U19507 (N_19507,N_19485,N_19408);
nor U19508 (N_19508,N_19441,N_19072);
nor U19509 (N_19509,N_19332,N_19263);
nor U19510 (N_19510,N_19009,N_19299);
and U19511 (N_19511,N_19343,N_19261);
nand U19512 (N_19512,N_19472,N_19459);
nor U19513 (N_19513,N_19149,N_19243);
and U19514 (N_19514,N_19123,N_19145);
nor U19515 (N_19515,N_19363,N_19384);
nand U19516 (N_19516,N_19455,N_19147);
nand U19517 (N_19517,N_19169,N_19436);
nor U19518 (N_19518,N_19304,N_19370);
nor U19519 (N_19519,N_19496,N_19062);
nand U19520 (N_19520,N_19355,N_19467);
nor U19521 (N_19521,N_19423,N_19295);
and U19522 (N_19522,N_19392,N_19082);
or U19523 (N_19523,N_19196,N_19110);
nand U19524 (N_19524,N_19206,N_19470);
and U19525 (N_19525,N_19069,N_19247);
nor U19526 (N_19526,N_19347,N_19089);
and U19527 (N_19527,N_19404,N_19151);
and U19528 (N_19528,N_19382,N_19088);
nand U19529 (N_19529,N_19164,N_19456);
and U19530 (N_19530,N_19195,N_19121);
nand U19531 (N_19531,N_19081,N_19060);
nand U19532 (N_19532,N_19492,N_19100);
nor U19533 (N_19533,N_19204,N_19481);
or U19534 (N_19534,N_19271,N_19024);
and U19535 (N_19535,N_19098,N_19115);
and U19536 (N_19536,N_19041,N_19112);
and U19537 (N_19537,N_19337,N_19039);
nor U19538 (N_19538,N_19443,N_19365);
nand U19539 (N_19539,N_19053,N_19253);
or U19540 (N_19540,N_19323,N_19330);
or U19541 (N_19541,N_19292,N_19190);
nor U19542 (N_19542,N_19236,N_19478);
or U19543 (N_19543,N_19182,N_19463);
nor U19544 (N_19544,N_19006,N_19083);
and U19545 (N_19545,N_19358,N_19313);
nor U19546 (N_19546,N_19157,N_19135);
nor U19547 (N_19547,N_19168,N_19440);
and U19548 (N_19548,N_19437,N_19460);
nand U19549 (N_19549,N_19439,N_19005);
nor U19550 (N_19550,N_19224,N_19497);
nor U19551 (N_19551,N_19327,N_19461);
and U19552 (N_19552,N_19391,N_19425);
nor U19553 (N_19553,N_19093,N_19156);
nor U19554 (N_19554,N_19143,N_19040);
or U19555 (N_19555,N_19430,N_19360);
nand U19556 (N_19556,N_19378,N_19312);
or U19557 (N_19557,N_19294,N_19427);
and U19558 (N_19558,N_19033,N_19176);
nor U19559 (N_19559,N_19124,N_19361);
or U19560 (N_19560,N_19488,N_19424);
or U19561 (N_19561,N_19191,N_19230);
nand U19562 (N_19562,N_19092,N_19364);
nand U19563 (N_19563,N_19338,N_19202);
nand U19564 (N_19564,N_19008,N_19002);
nand U19565 (N_19565,N_19153,N_19162);
nor U19566 (N_19566,N_19346,N_19303);
nand U19567 (N_19567,N_19289,N_19244);
nor U19568 (N_19568,N_19293,N_19200);
nor U19569 (N_19569,N_19042,N_19207);
and U19570 (N_19570,N_19057,N_19410);
and U19571 (N_19571,N_19442,N_19117);
nor U19572 (N_19572,N_19381,N_19141);
and U19573 (N_19573,N_19302,N_19016);
nor U19574 (N_19574,N_19187,N_19220);
and U19575 (N_19575,N_19268,N_19179);
nor U19576 (N_19576,N_19477,N_19239);
and U19577 (N_19577,N_19109,N_19248);
or U19578 (N_19578,N_19366,N_19315);
nor U19579 (N_19579,N_19394,N_19102);
nor U19580 (N_19580,N_19257,N_19129);
or U19581 (N_19581,N_19125,N_19379);
or U19582 (N_19582,N_19090,N_19446);
and U19583 (N_19583,N_19061,N_19166);
nand U19584 (N_19584,N_19105,N_19297);
or U19585 (N_19585,N_19415,N_19007);
nand U19586 (N_19586,N_19344,N_19291);
nor U19587 (N_19587,N_19262,N_19199);
nor U19588 (N_19588,N_19493,N_19300);
nor U19589 (N_19589,N_19174,N_19405);
nor U19590 (N_19590,N_19298,N_19094);
nor U19591 (N_19591,N_19375,N_19377);
or U19592 (N_19592,N_19480,N_19177);
nor U19593 (N_19593,N_19142,N_19211);
nor U19594 (N_19594,N_19227,N_19023);
and U19595 (N_19595,N_19296,N_19071);
nor U19596 (N_19596,N_19101,N_19235);
nand U19597 (N_19597,N_19362,N_19158);
or U19598 (N_19598,N_19019,N_19498);
nand U19599 (N_19599,N_19465,N_19342);
nor U19600 (N_19600,N_19272,N_19486);
nand U19601 (N_19601,N_19278,N_19281);
nand U19602 (N_19602,N_19201,N_19473);
and U19603 (N_19603,N_19047,N_19409);
nand U19604 (N_19604,N_19325,N_19310);
nand U19605 (N_19605,N_19468,N_19390);
nand U19606 (N_19606,N_19046,N_19170);
nor U19607 (N_19607,N_19445,N_19106);
and U19608 (N_19608,N_19031,N_19130);
and U19609 (N_19609,N_19104,N_19412);
nor U19610 (N_19610,N_19311,N_19221);
nor U19611 (N_19611,N_19017,N_19354);
or U19612 (N_19612,N_19067,N_19189);
nand U19613 (N_19613,N_19120,N_19103);
nor U19614 (N_19614,N_19079,N_19035);
and U19615 (N_19615,N_19249,N_19055);
and U19616 (N_19616,N_19475,N_19048);
and U19617 (N_19617,N_19334,N_19225);
and U19618 (N_19618,N_19237,N_19218);
nand U19619 (N_19619,N_19353,N_19396);
or U19620 (N_19620,N_19414,N_19373);
nand U19621 (N_19621,N_19215,N_19161);
or U19622 (N_19622,N_19265,N_19194);
or U19623 (N_19623,N_19228,N_19466);
and U19624 (N_19624,N_19350,N_19116);
and U19625 (N_19625,N_19021,N_19146);
nand U19626 (N_19626,N_19438,N_19469);
nor U19627 (N_19627,N_19181,N_19188);
nand U19628 (N_19628,N_19417,N_19231);
nor U19629 (N_19629,N_19399,N_19301);
nand U19630 (N_19630,N_19011,N_19385);
and U19631 (N_19631,N_19096,N_19139);
nor U19632 (N_19632,N_19052,N_19288);
nand U19633 (N_19633,N_19434,N_19027);
or U19634 (N_19634,N_19341,N_19322);
nor U19635 (N_19635,N_19000,N_19420);
nand U19636 (N_19636,N_19004,N_19336);
nand U19637 (N_19637,N_19026,N_19095);
or U19638 (N_19638,N_19321,N_19285);
and U19639 (N_19639,N_19260,N_19119);
nand U19640 (N_19640,N_19256,N_19279);
and U19641 (N_19641,N_19213,N_19449);
nor U19642 (N_19642,N_19163,N_19407);
and U19643 (N_19643,N_19320,N_19359);
and U19644 (N_19644,N_19212,N_19474);
and U19645 (N_19645,N_19136,N_19074);
nor U19646 (N_19646,N_19172,N_19209);
nand U19647 (N_19647,N_19028,N_19056);
and U19648 (N_19648,N_19490,N_19015);
and U19649 (N_19649,N_19203,N_19229);
or U19650 (N_19650,N_19085,N_19383);
nand U19651 (N_19651,N_19406,N_19097);
or U19652 (N_19652,N_19058,N_19210);
nand U19653 (N_19653,N_19454,N_19232);
or U19654 (N_19654,N_19077,N_19051);
nor U19655 (N_19655,N_19064,N_19482);
nor U19656 (N_19656,N_19114,N_19352);
and U19657 (N_19657,N_19198,N_19144);
nand U19658 (N_19658,N_19270,N_19214);
and U19659 (N_19659,N_19154,N_19403);
nand U19660 (N_19660,N_19025,N_19371);
nand U19661 (N_19661,N_19043,N_19429);
and U19662 (N_19662,N_19380,N_19118);
nand U19663 (N_19663,N_19167,N_19111);
nor U19664 (N_19664,N_19108,N_19258);
and U19665 (N_19665,N_19367,N_19233);
nand U19666 (N_19666,N_19329,N_19433);
and U19667 (N_19667,N_19222,N_19137);
and U19668 (N_19668,N_19476,N_19173);
or U19669 (N_19669,N_19387,N_19165);
and U19670 (N_19670,N_19284,N_19416);
or U19671 (N_19671,N_19063,N_19448);
and U19672 (N_19672,N_19277,N_19208);
or U19673 (N_19673,N_19418,N_19070);
nand U19674 (N_19674,N_19290,N_19132);
xnor U19675 (N_19675,N_19357,N_19251);
and U19676 (N_19676,N_19014,N_19241);
and U19677 (N_19677,N_19266,N_19388);
xnor U19678 (N_19678,N_19250,N_19489);
nand U19679 (N_19679,N_19020,N_19273);
nor U19680 (N_19680,N_19216,N_19259);
nand U19681 (N_19681,N_19086,N_19398);
or U19682 (N_19682,N_19462,N_19032);
or U19683 (N_19683,N_19345,N_19226);
or U19684 (N_19684,N_19305,N_19234);
or U19685 (N_19685,N_19107,N_19030);
and U19686 (N_19686,N_19049,N_19450);
nand U19687 (N_19687,N_19252,N_19317);
and U19688 (N_19688,N_19324,N_19044);
nor U19689 (N_19689,N_19283,N_19186);
and U19690 (N_19690,N_19495,N_19010);
or U19691 (N_19691,N_19319,N_19457);
nand U19692 (N_19692,N_19453,N_19374);
nand U19693 (N_19693,N_19134,N_19307);
nor U19694 (N_19694,N_19084,N_19185);
nor U19695 (N_19695,N_19421,N_19286);
nand U19696 (N_19696,N_19494,N_19076);
nand U19697 (N_19697,N_19451,N_19065);
and U19698 (N_19698,N_19148,N_19356);
or U19699 (N_19699,N_19389,N_19219);
nor U19700 (N_19700,N_19160,N_19386);
or U19701 (N_19701,N_19184,N_19059);
and U19702 (N_19702,N_19217,N_19029);
and U19703 (N_19703,N_19128,N_19397);
nand U19704 (N_19704,N_19447,N_19126);
nand U19705 (N_19705,N_19099,N_19133);
and U19706 (N_19706,N_19037,N_19335);
nor U19707 (N_19707,N_19393,N_19054);
and U19708 (N_19708,N_19238,N_19282);
nand U19709 (N_19709,N_19314,N_19431);
nor U19710 (N_19710,N_19287,N_19087);
nor U19711 (N_19711,N_19245,N_19242);
and U19712 (N_19712,N_19068,N_19045);
or U19713 (N_19713,N_19483,N_19308);
or U19714 (N_19714,N_19197,N_19432);
and U19715 (N_19715,N_19036,N_19034);
or U19716 (N_19716,N_19400,N_19152);
and U19717 (N_19717,N_19276,N_19066);
or U19718 (N_19718,N_19444,N_19178);
or U19719 (N_19719,N_19419,N_19267);
nor U19720 (N_19720,N_19376,N_19280);
or U19721 (N_19721,N_19269,N_19018);
nor U19722 (N_19722,N_19264,N_19351);
nand U19723 (N_19723,N_19331,N_19401);
nand U19724 (N_19724,N_19491,N_19193);
or U19725 (N_19725,N_19038,N_19205);
nand U19726 (N_19726,N_19254,N_19150);
nand U19727 (N_19727,N_19487,N_19091);
or U19728 (N_19728,N_19435,N_19131);
and U19729 (N_19729,N_19411,N_19073);
or U19730 (N_19730,N_19013,N_19138);
nand U19731 (N_19731,N_19180,N_19316);
nand U19732 (N_19732,N_19309,N_19413);
nor U19733 (N_19733,N_19471,N_19349);
nor U19734 (N_19734,N_19368,N_19140);
or U19735 (N_19735,N_19479,N_19050);
nand U19736 (N_19736,N_19484,N_19369);
nand U19737 (N_19737,N_19255,N_19075);
or U19738 (N_19738,N_19333,N_19080);
nand U19739 (N_19739,N_19372,N_19274);
nand U19740 (N_19740,N_19306,N_19452);
or U19741 (N_19741,N_19328,N_19402);
or U19742 (N_19742,N_19395,N_19183);
and U19743 (N_19743,N_19275,N_19175);
nor U19744 (N_19744,N_19022,N_19339);
xor U19745 (N_19745,N_19464,N_19003);
nor U19746 (N_19746,N_19192,N_19127);
and U19747 (N_19747,N_19159,N_19348);
nand U19748 (N_19748,N_19426,N_19246);
nand U19749 (N_19749,N_19223,N_19458);
and U19750 (N_19750,N_19264,N_19468);
and U19751 (N_19751,N_19073,N_19023);
nor U19752 (N_19752,N_19357,N_19171);
nand U19753 (N_19753,N_19144,N_19086);
and U19754 (N_19754,N_19216,N_19184);
nor U19755 (N_19755,N_19168,N_19042);
and U19756 (N_19756,N_19069,N_19055);
nor U19757 (N_19757,N_19147,N_19328);
nand U19758 (N_19758,N_19228,N_19292);
nor U19759 (N_19759,N_19174,N_19181);
or U19760 (N_19760,N_19010,N_19106);
and U19761 (N_19761,N_19047,N_19019);
and U19762 (N_19762,N_19336,N_19233);
and U19763 (N_19763,N_19155,N_19308);
nand U19764 (N_19764,N_19121,N_19224);
nor U19765 (N_19765,N_19475,N_19338);
nand U19766 (N_19766,N_19369,N_19334);
or U19767 (N_19767,N_19065,N_19091);
or U19768 (N_19768,N_19338,N_19411);
or U19769 (N_19769,N_19146,N_19469);
or U19770 (N_19770,N_19275,N_19334);
nand U19771 (N_19771,N_19337,N_19281);
nor U19772 (N_19772,N_19300,N_19360);
nand U19773 (N_19773,N_19484,N_19100);
nand U19774 (N_19774,N_19458,N_19252);
or U19775 (N_19775,N_19164,N_19044);
or U19776 (N_19776,N_19125,N_19342);
nand U19777 (N_19777,N_19164,N_19184);
nand U19778 (N_19778,N_19389,N_19180);
nor U19779 (N_19779,N_19046,N_19197);
or U19780 (N_19780,N_19045,N_19054);
or U19781 (N_19781,N_19130,N_19185);
or U19782 (N_19782,N_19433,N_19174);
or U19783 (N_19783,N_19052,N_19081);
nand U19784 (N_19784,N_19371,N_19078);
nand U19785 (N_19785,N_19090,N_19461);
nand U19786 (N_19786,N_19125,N_19404);
nor U19787 (N_19787,N_19159,N_19464);
and U19788 (N_19788,N_19028,N_19061);
nand U19789 (N_19789,N_19291,N_19424);
or U19790 (N_19790,N_19331,N_19154);
nand U19791 (N_19791,N_19141,N_19015);
or U19792 (N_19792,N_19005,N_19474);
nand U19793 (N_19793,N_19010,N_19490);
nand U19794 (N_19794,N_19080,N_19068);
or U19795 (N_19795,N_19068,N_19490);
or U19796 (N_19796,N_19054,N_19275);
nand U19797 (N_19797,N_19227,N_19476);
nor U19798 (N_19798,N_19108,N_19219);
nand U19799 (N_19799,N_19308,N_19040);
and U19800 (N_19800,N_19225,N_19248);
or U19801 (N_19801,N_19362,N_19471);
nand U19802 (N_19802,N_19472,N_19046);
and U19803 (N_19803,N_19052,N_19478);
nand U19804 (N_19804,N_19184,N_19395);
nor U19805 (N_19805,N_19207,N_19144);
nand U19806 (N_19806,N_19492,N_19457);
and U19807 (N_19807,N_19404,N_19261);
nand U19808 (N_19808,N_19331,N_19162);
and U19809 (N_19809,N_19254,N_19483);
nand U19810 (N_19810,N_19301,N_19188);
or U19811 (N_19811,N_19386,N_19437);
nand U19812 (N_19812,N_19444,N_19184);
nand U19813 (N_19813,N_19458,N_19140);
nor U19814 (N_19814,N_19357,N_19039);
xor U19815 (N_19815,N_19064,N_19422);
nand U19816 (N_19816,N_19094,N_19115);
or U19817 (N_19817,N_19452,N_19498);
and U19818 (N_19818,N_19072,N_19292);
and U19819 (N_19819,N_19308,N_19290);
nand U19820 (N_19820,N_19017,N_19232);
nor U19821 (N_19821,N_19298,N_19301);
nor U19822 (N_19822,N_19435,N_19434);
or U19823 (N_19823,N_19174,N_19301);
or U19824 (N_19824,N_19346,N_19425);
nand U19825 (N_19825,N_19488,N_19099);
nand U19826 (N_19826,N_19296,N_19144);
or U19827 (N_19827,N_19226,N_19079);
nand U19828 (N_19828,N_19484,N_19129);
and U19829 (N_19829,N_19234,N_19037);
nor U19830 (N_19830,N_19106,N_19416);
or U19831 (N_19831,N_19481,N_19090);
and U19832 (N_19832,N_19460,N_19449);
nand U19833 (N_19833,N_19069,N_19495);
nand U19834 (N_19834,N_19034,N_19272);
nand U19835 (N_19835,N_19460,N_19203);
and U19836 (N_19836,N_19361,N_19255);
xnor U19837 (N_19837,N_19286,N_19156);
nor U19838 (N_19838,N_19231,N_19153);
nor U19839 (N_19839,N_19217,N_19038);
nor U19840 (N_19840,N_19283,N_19488);
or U19841 (N_19841,N_19074,N_19309);
nor U19842 (N_19842,N_19473,N_19485);
nand U19843 (N_19843,N_19432,N_19113);
and U19844 (N_19844,N_19315,N_19436);
nor U19845 (N_19845,N_19033,N_19495);
nand U19846 (N_19846,N_19063,N_19383);
nor U19847 (N_19847,N_19077,N_19429);
or U19848 (N_19848,N_19054,N_19038);
nor U19849 (N_19849,N_19060,N_19121);
or U19850 (N_19850,N_19056,N_19246);
and U19851 (N_19851,N_19391,N_19280);
nor U19852 (N_19852,N_19060,N_19043);
nand U19853 (N_19853,N_19348,N_19424);
nand U19854 (N_19854,N_19129,N_19415);
or U19855 (N_19855,N_19109,N_19163);
and U19856 (N_19856,N_19018,N_19453);
or U19857 (N_19857,N_19077,N_19176);
nor U19858 (N_19858,N_19038,N_19391);
or U19859 (N_19859,N_19001,N_19310);
nor U19860 (N_19860,N_19119,N_19308);
nor U19861 (N_19861,N_19214,N_19153);
or U19862 (N_19862,N_19238,N_19443);
and U19863 (N_19863,N_19090,N_19436);
and U19864 (N_19864,N_19483,N_19111);
nor U19865 (N_19865,N_19125,N_19217);
and U19866 (N_19866,N_19362,N_19387);
nand U19867 (N_19867,N_19036,N_19408);
nor U19868 (N_19868,N_19051,N_19388);
nand U19869 (N_19869,N_19061,N_19169);
and U19870 (N_19870,N_19413,N_19350);
or U19871 (N_19871,N_19150,N_19018);
nor U19872 (N_19872,N_19243,N_19008);
nand U19873 (N_19873,N_19155,N_19059);
nor U19874 (N_19874,N_19338,N_19469);
or U19875 (N_19875,N_19360,N_19357);
nor U19876 (N_19876,N_19237,N_19096);
nor U19877 (N_19877,N_19045,N_19299);
nand U19878 (N_19878,N_19012,N_19451);
or U19879 (N_19879,N_19080,N_19048);
nor U19880 (N_19880,N_19233,N_19105);
or U19881 (N_19881,N_19273,N_19108);
or U19882 (N_19882,N_19142,N_19441);
nor U19883 (N_19883,N_19293,N_19322);
or U19884 (N_19884,N_19282,N_19144);
nor U19885 (N_19885,N_19083,N_19213);
or U19886 (N_19886,N_19094,N_19027);
and U19887 (N_19887,N_19066,N_19196);
and U19888 (N_19888,N_19227,N_19243);
and U19889 (N_19889,N_19011,N_19207);
or U19890 (N_19890,N_19366,N_19311);
nor U19891 (N_19891,N_19205,N_19443);
nand U19892 (N_19892,N_19100,N_19454);
nand U19893 (N_19893,N_19181,N_19082);
nand U19894 (N_19894,N_19195,N_19392);
nor U19895 (N_19895,N_19165,N_19119);
nor U19896 (N_19896,N_19259,N_19055);
nand U19897 (N_19897,N_19047,N_19146);
nand U19898 (N_19898,N_19102,N_19411);
nand U19899 (N_19899,N_19383,N_19053);
xor U19900 (N_19900,N_19464,N_19022);
nor U19901 (N_19901,N_19344,N_19085);
or U19902 (N_19902,N_19194,N_19042);
nand U19903 (N_19903,N_19148,N_19436);
nand U19904 (N_19904,N_19035,N_19285);
or U19905 (N_19905,N_19308,N_19170);
and U19906 (N_19906,N_19124,N_19313);
nand U19907 (N_19907,N_19258,N_19187);
nand U19908 (N_19908,N_19126,N_19037);
nor U19909 (N_19909,N_19324,N_19396);
and U19910 (N_19910,N_19103,N_19435);
and U19911 (N_19911,N_19191,N_19138);
or U19912 (N_19912,N_19471,N_19273);
or U19913 (N_19913,N_19379,N_19335);
and U19914 (N_19914,N_19285,N_19100);
nor U19915 (N_19915,N_19063,N_19409);
nand U19916 (N_19916,N_19069,N_19134);
nor U19917 (N_19917,N_19092,N_19122);
or U19918 (N_19918,N_19353,N_19000);
and U19919 (N_19919,N_19208,N_19176);
and U19920 (N_19920,N_19208,N_19464);
and U19921 (N_19921,N_19235,N_19146);
nand U19922 (N_19922,N_19386,N_19492);
or U19923 (N_19923,N_19493,N_19104);
or U19924 (N_19924,N_19192,N_19396);
and U19925 (N_19925,N_19062,N_19371);
nand U19926 (N_19926,N_19294,N_19131);
and U19927 (N_19927,N_19344,N_19202);
nor U19928 (N_19928,N_19292,N_19253);
and U19929 (N_19929,N_19337,N_19245);
and U19930 (N_19930,N_19386,N_19220);
nor U19931 (N_19931,N_19139,N_19259);
or U19932 (N_19932,N_19305,N_19200);
or U19933 (N_19933,N_19252,N_19384);
or U19934 (N_19934,N_19369,N_19088);
nand U19935 (N_19935,N_19287,N_19414);
nand U19936 (N_19936,N_19158,N_19356);
or U19937 (N_19937,N_19113,N_19034);
nand U19938 (N_19938,N_19335,N_19084);
and U19939 (N_19939,N_19049,N_19128);
nand U19940 (N_19940,N_19212,N_19179);
nand U19941 (N_19941,N_19275,N_19480);
and U19942 (N_19942,N_19358,N_19376);
and U19943 (N_19943,N_19012,N_19029);
or U19944 (N_19944,N_19423,N_19057);
nor U19945 (N_19945,N_19075,N_19489);
nand U19946 (N_19946,N_19024,N_19286);
nor U19947 (N_19947,N_19110,N_19416);
nand U19948 (N_19948,N_19191,N_19283);
nor U19949 (N_19949,N_19027,N_19038);
xor U19950 (N_19950,N_19493,N_19340);
nand U19951 (N_19951,N_19362,N_19041);
nor U19952 (N_19952,N_19023,N_19486);
and U19953 (N_19953,N_19276,N_19121);
nor U19954 (N_19954,N_19455,N_19069);
and U19955 (N_19955,N_19207,N_19021);
and U19956 (N_19956,N_19417,N_19463);
nand U19957 (N_19957,N_19199,N_19446);
and U19958 (N_19958,N_19296,N_19318);
nand U19959 (N_19959,N_19464,N_19201);
nand U19960 (N_19960,N_19457,N_19072);
nor U19961 (N_19961,N_19472,N_19157);
or U19962 (N_19962,N_19055,N_19324);
or U19963 (N_19963,N_19347,N_19122);
nand U19964 (N_19964,N_19282,N_19124);
nor U19965 (N_19965,N_19423,N_19317);
nand U19966 (N_19966,N_19060,N_19271);
nor U19967 (N_19967,N_19124,N_19109);
and U19968 (N_19968,N_19039,N_19292);
or U19969 (N_19969,N_19319,N_19490);
nor U19970 (N_19970,N_19058,N_19372);
or U19971 (N_19971,N_19353,N_19099);
and U19972 (N_19972,N_19229,N_19351);
nor U19973 (N_19973,N_19041,N_19129);
nor U19974 (N_19974,N_19247,N_19304);
and U19975 (N_19975,N_19260,N_19355);
nand U19976 (N_19976,N_19452,N_19433);
or U19977 (N_19977,N_19255,N_19347);
nand U19978 (N_19978,N_19053,N_19027);
or U19979 (N_19979,N_19276,N_19383);
and U19980 (N_19980,N_19123,N_19128);
nor U19981 (N_19981,N_19033,N_19283);
nor U19982 (N_19982,N_19146,N_19428);
and U19983 (N_19983,N_19329,N_19201);
nor U19984 (N_19984,N_19193,N_19489);
nand U19985 (N_19985,N_19409,N_19405);
nor U19986 (N_19986,N_19391,N_19051);
or U19987 (N_19987,N_19156,N_19426);
nand U19988 (N_19988,N_19292,N_19466);
nand U19989 (N_19989,N_19485,N_19048);
nand U19990 (N_19990,N_19287,N_19388);
nor U19991 (N_19991,N_19120,N_19034);
and U19992 (N_19992,N_19234,N_19173);
nor U19993 (N_19993,N_19224,N_19399);
nand U19994 (N_19994,N_19369,N_19329);
nor U19995 (N_19995,N_19411,N_19311);
nor U19996 (N_19996,N_19032,N_19033);
or U19997 (N_19997,N_19226,N_19158);
nand U19998 (N_19998,N_19490,N_19057);
or U19999 (N_19999,N_19024,N_19263);
or UO_0 (O_0,N_19905,N_19775);
nor UO_1 (O_1,N_19908,N_19979);
or UO_2 (O_2,N_19831,N_19797);
and UO_3 (O_3,N_19944,N_19836);
or UO_4 (O_4,N_19880,N_19695);
and UO_5 (O_5,N_19582,N_19902);
nand UO_6 (O_6,N_19869,N_19606);
nor UO_7 (O_7,N_19983,N_19516);
or UO_8 (O_8,N_19533,N_19593);
nand UO_9 (O_9,N_19631,N_19649);
or UO_10 (O_10,N_19567,N_19921);
nand UO_11 (O_11,N_19827,N_19923);
nand UO_12 (O_12,N_19885,N_19657);
and UO_13 (O_13,N_19772,N_19559);
and UO_14 (O_14,N_19914,N_19592);
and UO_15 (O_15,N_19726,N_19652);
nand UO_16 (O_16,N_19656,N_19971);
and UO_17 (O_17,N_19874,N_19724);
nor UO_18 (O_18,N_19688,N_19760);
or UO_19 (O_19,N_19798,N_19694);
nand UO_20 (O_20,N_19612,N_19574);
nand UO_21 (O_21,N_19632,N_19852);
nor UO_22 (O_22,N_19994,N_19997);
nand UO_23 (O_23,N_19583,N_19960);
nor UO_24 (O_24,N_19662,N_19986);
nor UO_25 (O_25,N_19515,N_19881);
or UO_26 (O_26,N_19517,N_19759);
and UO_27 (O_27,N_19858,N_19868);
and UO_28 (O_28,N_19890,N_19973);
nand UO_29 (O_29,N_19672,N_19528);
nor UO_30 (O_30,N_19544,N_19581);
nand UO_31 (O_31,N_19505,N_19791);
nand UO_32 (O_32,N_19703,N_19549);
nor UO_33 (O_33,N_19901,N_19660);
nor UO_34 (O_34,N_19906,N_19721);
or UO_35 (O_35,N_19771,N_19774);
or UO_36 (O_36,N_19783,N_19830);
nor UO_37 (O_37,N_19933,N_19638);
and UO_38 (O_38,N_19879,N_19807);
or UO_39 (O_39,N_19961,N_19982);
nor UO_40 (O_40,N_19750,N_19706);
nor UO_41 (O_41,N_19822,N_19806);
nor UO_42 (O_42,N_19598,N_19835);
nor UO_43 (O_43,N_19898,N_19911);
nand UO_44 (O_44,N_19635,N_19571);
or UO_45 (O_45,N_19794,N_19641);
nand UO_46 (O_46,N_19870,N_19915);
nand UO_47 (O_47,N_19620,N_19848);
and UO_48 (O_48,N_19539,N_19556);
or UO_49 (O_49,N_19940,N_19990);
nand UO_50 (O_50,N_19579,N_19773);
or UO_51 (O_51,N_19931,N_19745);
nand UO_52 (O_52,N_19817,N_19823);
nand UO_53 (O_53,N_19749,N_19934);
and UO_54 (O_54,N_19849,N_19551);
nand UO_55 (O_55,N_19670,N_19865);
and UO_56 (O_56,N_19954,N_19946);
nor UO_57 (O_57,N_19648,N_19838);
or UO_58 (O_58,N_19613,N_19536);
and UO_59 (O_59,N_19634,N_19628);
nor UO_60 (O_60,N_19607,N_19938);
xor UO_61 (O_61,N_19702,N_19991);
nor UO_62 (O_62,N_19969,N_19562);
or UO_63 (O_63,N_19913,N_19941);
and UO_64 (O_64,N_19585,N_19644);
or UO_65 (O_65,N_19734,N_19981);
nor UO_66 (O_66,N_19597,N_19844);
and UO_67 (O_67,N_19968,N_19900);
and UO_68 (O_68,N_19919,N_19978);
or UO_69 (O_69,N_19603,N_19553);
nand UO_70 (O_70,N_19594,N_19936);
nor UO_71 (O_71,N_19777,N_19565);
nand UO_72 (O_72,N_19639,N_19974);
or UO_73 (O_73,N_19625,N_19570);
nor UO_74 (O_74,N_19821,N_19850);
or UO_75 (O_75,N_19698,N_19563);
nand UO_76 (O_76,N_19996,N_19928);
and UO_77 (O_77,N_19526,N_19650);
nor UO_78 (O_78,N_19564,N_19867);
and UO_79 (O_79,N_19897,N_19595);
xnor UO_80 (O_80,N_19792,N_19600);
nand UO_81 (O_81,N_19682,N_19531);
or UO_82 (O_82,N_19808,N_19939);
nor UO_83 (O_83,N_19891,N_19521);
nor UO_84 (O_84,N_19882,N_19601);
or UO_85 (O_85,N_19833,N_19910);
nor UO_86 (O_86,N_19679,N_19520);
nand UO_87 (O_87,N_19976,N_19876);
nand UO_88 (O_88,N_19655,N_19989);
nand UO_89 (O_89,N_19930,N_19788);
or UO_90 (O_90,N_19937,N_19610);
nor UO_91 (O_91,N_19999,N_19691);
and UO_92 (O_92,N_19664,N_19751);
or UO_93 (O_93,N_19731,N_19646);
nor UO_94 (O_94,N_19853,N_19545);
or UO_95 (O_95,N_19741,N_19569);
nor UO_96 (O_96,N_19675,N_19727);
nor UO_97 (O_97,N_19503,N_19918);
and UO_98 (O_98,N_19681,N_19965);
nand UO_99 (O_99,N_19604,N_19651);
nor UO_100 (O_100,N_19627,N_19894);
nor UO_101 (O_101,N_19711,N_19926);
or UO_102 (O_102,N_19828,N_19889);
or UO_103 (O_103,N_19769,N_19952);
and UO_104 (O_104,N_19715,N_19815);
and UO_105 (O_105,N_19927,N_19744);
and UO_106 (O_106,N_19614,N_19813);
or UO_107 (O_107,N_19532,N_19980);
or UO_108 (O_108,N_19924,N_19862);
or UO_109 (O_109,N_19733,N_19696);
and UO_110 (O_110,N_19818,N_19514);
nand UO_111 (O_111,N_19780,N_19878);
nand UO_112 (O_112,N_19693,N_19617);
or UO_113 (O_113,N_19587,N_19500);
nand UO_114 (O_114,N_19762,N_19608);
nand UO_115 (O_115,N_19998,N_19800);
nor UO_116 (O_116,N_19804,N_19642);
and UO_117 (O_117,N_19895,N_19524);
nor UO_118 (O_118,N_19713,N_19697);
nor UO_119 (O_119,N_19511,N_19609);
or UO_120 (O_120,N_19837,N_19955);
or UO_121 (O_121,N_19640,N_19964);
and UO_122 (O_122,N_19674,N_19892);
nor UO_123 (O_123,N_19737,N_19596);
or UO_124 (O_124,N_19963,N_19554);
and UO_125 (O_125,N_19787,N_19666);
nor UO_126 (O_126,N_19805,N_19790);
or UO_127 (O_127,N_19728,N_19912);
or UO_128 (O_128,N_19720,N_19739);
nand UO_129 (O_129,N_19586,N_19678);
nand UO_130 (O_130,N_19856,N_19685);
and UO_131 (O_131,N_19776,N_19538);
nor UO_132 (O_132,N_19757,N_19943);
nand UO_133 (O_133,N_19863,N_19584);
or UO_134 (O_134,N_19802,N_19875);
and UO_135 (O_135,N_19784,N_19920);
nor UO_136 (O_136,N_19888,N_19717);
or UO_137 (O_137,N_19967,N_19993);
nor UO_138 (O_138,N_19883,N_19873);
nor UO_139 (O_139,N_19846,N_19618);
nor UO_140 (O_140,N_19667,N_19866);
nand UO_141 (O_141,N_19832,N_19576);
nand UO_142 (O_142,N_19899,N_19506);
nor UO_143 (O_143,N_19537,N_19718);
nand UO_144 (O_144,N_19507,N_19962);
or UO_145 (O_145,N_19884,N_19530);
nor UO_146 (O_146,N_19752,N_19854);
xor UO_147 (O_147,N_19985,N_19522);
or UO_148 (O_148,N_19768,N_19743);
nand UO_149 (O_149,N_19577,N_19972);
and UO_150 (O_150,N_19732,N_19810);
or UO_151 (O_151,N_19557,N_19599);
nand UO_152 (O_152,N_19909,N_19668);
or UO_153 (O_153,N_19578,N_19723);
and UO_154 (O_154,N_19619,N_19840);
nor UO_155 (O_155,N_19621,N_19636);
nor UO_156 (O_156,N_19987,N_19527);
and UO_157 (O_157,N_19623,N_19633);
and UO_158 (O_158,N_19630,N_19548);
or UO_159 (O_159,N_19730,N_19842);
nor UO_160 (O_160,N_19786,N_19781);
nand UO_161 (O_161,N_19575,N_19859);
and UO_162 (O_162,N_19966,N_19782);
or UO_163 (O_163,N_19949,N_19669);
nand UO_164 (O_164,N_19887,N_19673);
nor UO_165 (O_165,N_19701,N_19801);
or UO_166 (O_166,N_19676,N_19796);
nand UO_167 (O_167,N_19712,N_19543);
nand UO_168 (O_168,N_19550,N_19951);
and UO_169 (O_169,N_19716,N_19518);
nand UO_170 (O_170,N_19851,N_19977);
nor UO_171 (O_171,N_19922,N_19795);
or UO_172 (O_172,N_19568,N_19573);
nand UO_173 (O_173,N_19742,N_19552);
nor UO_174 (O_174,N_19812,N_19611);
nor UO_175 (O_175,N_19546,N_19659);
nand UO_176 (O_176,N_19907,N_19513);
or UO_177 (O_177,N_19975,N_19722);
or UO_178 (O_178,N_19756,N_19626);
nor UO_179 (O_179,N_19605,N_19841);
nand UO_180 (O_180,N_19629,N_19956);
nor UO_181 (O_181,N_19917,N_19705);
nor UO_182 (O_182,N_19534,N_19942);
nor UO_183 (O_183,N_19845,N_19714);
nor UO_184 (O_184,N_19764,N_19680);
xnor UO_185 (O_185,N_19708,N_19510);
and UO_186 (O_186,N_19725,N_19803);
or UO_187 (O_187,N_19529,N_19541);
nor UO_188 (O_188,N_19825,N_19658);
and UO_189 (O_189,N_19809,N_19893);
and UO_190 (O_190,N_19872,N_19671);
and UO_191 (O_191,N_19778,N_19643);
nand UO_192 (O_192,N_19519,N_19896);
and UO_193 (O_193,N_19948,N_19677);
nand UO_194 (O_194,N_19589,N_19709);
or UO_195 (O_195,N_19653,N_19735);
or UO_196 (O_196,N_19847,N_19616);
or UO_197 (O_197,N_19591,N_19523);
nor UO_198 (O_198,N_19729,N_19748);
and UO_199 (O_199,N_19588,N_19740);
and UO_200 (O_200,N_19689,N_19645);
and UO_201 (O_201,N_19829,N_19699);
nor UO_202 (O_202,N_19566,N_19779);
and UO_203 (O_203,N_19861,N_19710);
or UO_204 (O_204,N_19590,N_19560);
and UO_205 (O_205,N_19504,N_19819);
nor UO_206 (O_206,N_19864,N_19558);
and UO_207 (O_207,N_19785,N_19793);
and UO_208 (O_208,N_19502,N_19647);
nand UO_209 (O_209,N_19970,N_19811);
nor UO_210 (O_210,N_19663,N_19857);
nand UO_211 (O_211,N_19755,N_19707);
or UO_212 (O_212,N_19860,N_19959);
or UO_213 (O_213,N_19988,N_19665);
xor UO_214 (O_214,N_19816,N_19525);
nor UO_215 (O_215,N_19947,N_19766);
and UO_216 (O_216,N_19501,N_19767);
nor UO_217 (O_217,N_19763,N_19738);
and UO_218 (O_218,N_19834,N_19615);
nand UO_219 (O_219,N_19684,N_19542);
or UO_220 (O_220,N_19984,N_19916);
or UO_221 (O_221,N_19704,N_19687);
nor UO_222 (O_222,N_19690,N_19929);
nor UO_223 (O_223,N_19508,N_19746);
nor UO_224 (O_224,N_19839,N_19904);
nor UO_225 (O_225,N_19903,N_19602);
nor UO_226 (O_226,N_19761,N_19719);
nor UO_227 (O_227,N_19950,N_19572);
nand UO_228 (O_228,N_19753,N_19789);
nand UO_229 (O_229,N_19561,N_19624);
nor UO_230 (O_230,N_19692,N_19871);
nand UO_231 (O_231,N_19995,N_19540);
nand UO_232 (O_232,N_19637,N_19953);
nor UO_233 (O_233,N_19935,N_19799);
or UO_234 (O_234,N_19855,N_19958);
or UO_235 (O_235,N_19945,N_19820);
and UO_236 (O_236,N_19555,N_19843);
and UO_237 (O_237,N_19765,N_19877);
nand UO_238 (O_238,N_19770,N_19826);
and UO_239 (O_239,N_19509,N_19824);
nand UO_240 (O_240,N_19547,N_19686);
and UO_241 (O_241,N_19754,N_19512);
nand UO_242 (O_242,N_19932,N_19992);
and UO_243 (O_243,N_19683,N_19814);
or UO_244 (O_244,N_19654,N_19747);
nand UO_245 (O_245,N_19580,N_19535);
nand UO_246 (O_246,N_19886,N_19758);
nand UO_247 (O_247,N_19661,N_19622);
nand UO_248 (O_248,N_19700,N_19957);
nand UO_249 (O_249,N_19925,N_19736);
nand UO_250 (O_250,N_19745,N_19832);
nor UO_251 (O_251,N_19877,N_19673);
nor UO_252 (O_252,N_19902,N_19815);
or UO_253 (O_253,N_19569,N_19926);
or UO_254 (O_254,N_19872,N_19708);
and UO_255 (O_255,N_19686,N_19892);
nand UO_256 (O_256,N_19745,N_19557);
and UO_257 (O_257,N_19878,N_19699);
or UO_258 (O_258,N_19531,N_19528);
and UO_259 (O_259,N_19747,N_19717);
or UO_260 (O_260,N_19593,N_19766);
or UO_261 (O_261,N_19535,N_19934);
nand UO_262 (O_262,N_19618,N_19525);
nor UO_263 (O_263,N_19880,N_19706);
nand UO_264 (O_264,N_19685,N_19602);
nor UO_265 (O_265,N_19923,N_19955);
or UO_266 (O_266,N_19615,N_19919);
and UO_267 (O_267,N_19912,N_19609);
and UO_268 (O_268,N_19803,N_19844);
nand UO_269 (O_269,N_19664,N_19633);
and UO_270 (O_270,N_19978,N_19682);
nand UO_271 (O_271,N_19506,N_19608);
or UO_272 (O_272,N_19714,N_19567);
nor UO_273 (O_273,N_19795,N_19827);
or UO_274 (O_274,N_19616,N_19811);
or UO_275 (O_275,N_19648,N_19802);
nor UO_276 (O_276,N_19928,N_19873);
nor UO_277 (O_277,N_19641,N_19976);
nor UO_278 (O_278,N_19837,N_19566);
and UO_279 (O_279,N_19848,N_19699);
nor UO_280 (O_280,N_19800,N_19549);
or UO_281 (O_281,N_19598,N_19850);
nand UO_282 (O_282,N_19879,N_19626);
or UO_283 (O_283,N_19575,N_19844);
nor UO_284 (O_284,N_19904,N_19878);
or UO_285 (O_285,N_19623,N_19859);
nor UO_286 (O_286,N_19870,N_19956);
and UO_287 (O_287,N_19665,N_19506);
and UO_288 (O_288,N_19772,N_19633);
nand UO_289 (O_289,N_19936,N_19828);
and UO_290 (O_290,N_19524,N_19810);
and UO_291 (O_291,N_19611,N_19757);
nand UO_292 (O_292,N_19646,N_19927);
nand UO_293 (O_293,N_19667,N_19530);
nor UO_294 (O_294,N_19937,N_19591);
nor UO_295 (O_295,N_19700,N_19863);
nor UO_296 (O_296,N_19595,N_19622);
and UO_297 (O_297,N_19750,N_19798);
nor UO_298 (O_298,N_19584,N_19793);
nor UO_299 (O_299,N_19504,N_19943);
or UO_300 (O_300,N_19607,N_19895);
nand UO_301 (O_301,N_19695,N_19863);
nand UO_302 (O_302,N_19882,N_19815);
and UO_303 (O_303,N_19818,N_19930);
or UO_304 (O_304,N_19708,N_19831);
or UO_305 (O_305,N_19622,N_19587);
nor UO_306 (O_306,N_19734,N_19920);
nor UO_307 (O_307,N_19727,N_19682);
and UO_308 (O_308,N_19996,N_19975);
or UO_309 (O_309,N_19542,N_19838);
nor UO_310 (O_310,N_19993,N_19728);
nor UO_311 (O_311,N_19929,N_19954);
and UO_312 (O_312,N_19720,N_19575);
and UO_313 (O_313,N_19884,N_19595);
or UO_314 (O_314,N_19961,N_19803);
and UO_315 (O_315,N_19698,N_19938);
nor UO_316 (O_316,N_19895,N_19835);
or UO_317 (O_317,N_19726,N_19731);
nand UO_318 (O_318,N_19845,N_19533);
and UO_319 (O_319,N_19719,N_19619);
nand UO_320 (O_320,N_19611,N_19887);
nand UO_321 (O_321,N_19677,N_19659);
nor UO_322 (O_322,N_19557,N_19762);
or UO_323 (O_323,N_19721,N_19641);
xnor UO_324 (O_324,N_19787,N_19892);
nor UO_325 (O_325,N_19589,N_19710);
or UO_326 (O_326,N_19735,N_19748);
nor UO_327 (O_327,N_19518,N_19782);
or UO_328 (O_328,N_19628,N_19973);
and UO_329 (O_329,N_19834,N_19942);
nor UO_330 (O_330,N_19690,N_19535);
nand UO_331 (O_331,N_19835,N_19886);
nor UO_332 (O_332,N_19541,N_19663);
or UO_333 (O_333,N_19912,N_19561);
and UO_334 (O_334,N_19807,N_19570);
and UO_335 (O_335,N_19712,N_19736);
xor UO_336 (O_336,N_19690,N_19661);
or UO_337 (O_337,N_19978,N_19642);
nor UO_338 (O_338,N_19653,N_19654);
or UO_339 (O_339,N_19667,N_19918);
nand UO_340 (O_340,N_19671,N_19606);
or UO_341 (O_341,N_19530,N_19974);
nand UO_342 (O_342,N_19960,N_19531);
nor UO_343 (O_343,N_19864,N_19640);
and UO_344 (O_344,N_19513,N_19611);
nand UO_345 (O_345,N_19817,N_19831);
and UO_346 (O_346,N_19901,N_19543);
or UO_347 (O_347,N_19641,N_19595);
and UO_348 (O_348,N_19637,N_19845);
nor UO_349 (O_349,N_19850,N_19589);
and UO_350 (O_350,N_19742,N_19981);
or UO_351 (O_351,N_19637,N_19904);
or UO_352 (O_352,N_19506,N_19618);
nand UO_353 (O_353,N_19944,N_19562);
or UO_354 (O_354,N_19567,N_19975);
nor UO_355 (O_355,N_19624,N_19957);
or UO_356 (O_356,N_19685,N_19596);
and UO_357 (O_357,N_19769,N_19937);
and UO_358 (O_358,N_19760,N_19996);
and UO_359 (O_359,N_19874,N_19737);
or UO_360 (O_360,N_19866,N_19560);
nor UO_361 (O_361,N_19672,N_19765);
and UO_362 (O_362,N_19875,N_19525);
and UO_363 (O_363,N_19873,N_19878);
and UO_364 (O_364,N_19872,N_19580);
nand UO_365 (O_365,N_19689,N_19623);
nor UO_366 (O_366,N_19896,N_19637);
or UO_367 (O_367,N_19732,N_19885);
nor UO_368 (O_368,N_19804,N_19987);
nor UO_369 (O_369,N_19973,N_19583);
nand UO_370 (O_370,N_19775,N_19866);
nand UO_371 (O_371,N_19614,N_19611);
nor UO_372 (O_372,N_19940,N_19710);
or UO_373 (O_373,N_19755,N_19819);
and UO_374 (O_374,N_19730,N_19921);
or UO_375 (O_375,N_19977,N_19984);
nand UO_376 (O_376,N_19713,N_19902);
or UO_377 (O_377,N_19759,N_19718);
and UO_378 (O_378,N_19936,N_19768);
nand UO_379 (O_379,N_19936,N_19813);
and UO_380 (O_380,N_19551,N_19872);
nand UO_381 (O_381,N_19623,N_19991);
nand UO_382 (O_382,N_19733,N_19545);
xnor UO_383 (O_383,N_19999,N_19573);
nand UO_384 (O_384,N_19936,N_19656);
and UO_385 (O_385,N_19876,N_19777);
nor UO_386 (O_386,N_19653,N_19793);
nand UO_387 (O_387,N_19563,N_19723);
nor UO_388 (O_388,N_19810,N_19911);
and UO_389 (O_389,N_19979,N_19718);
or UO_390 (O_390,N_19925,N_19755);
and UO_391 (O_391,N_19876,N_19826);
or UO_392 (O_392,N_19698,N_19557);
and UO_393 (O_393,N_19896,N_19975);
nand UO_394 (O_394,N_19881,N_19806);
or UO_395 (O_395,N_19810,N_19811);
and UO_396 (O_396,N_19845,N_19874);
nand UO_397 (O_397,N_19598,N_19587);
nor UO_398 (O_398,N_19778,N_19975);
or UO_399 (O_399,N_19773,N_19567);
or UO_400 (O_400,N_19778,N_19583);
and UO_401 (O_401,N_19516,N_19894);
nor UO_402 (O_402,N_19720,N_19886);
nor UO_403 (O_403,N_19531,N_19673);
nand UO_404 (O_404,N_19816,N_19960);
or UO_405 (O_405,N_19611,N_19553);
nor UO_406 (O_406,N_19996,N_19796);
nor UO_407 (O_407,N_19709,N_19566);
nor UO_408 (O_408,N_19772,N_19604);
nand UO_409 (O_409,N_19842,N_19761);
and UO_410 (O_410,N_19977,N_19784);
nor UO_411 (O_411,N_19909,N_19795);
nand UO_412 (O_412,N_19593,N_19804);
nand UO_413 (O_413,N_19584,N_19575);
or UO_414 (O_414,N_19728,N_19533);
nor UO_415 (O_415,N_19989,N_19525);
or UO_416 (O_416,N_19936,N_19806);
and UO_417 (O_417,N_19616,N_19537);
nand UO_418 (O_418,N_19524,N_19887);
nand UO_419 (O_419,N_19509,N_19829);
and UO_420 (O_420,N_19910,N_19544);
nor UO_421 (O_421,N_19626,N_19646);
nor UO_422 (O_422,N_19668,N_19774);
nor UO_423 (O_423,N_19860,N_19790);
or UO_424 (O_424,N_19704,N_19620);
nor UO_425 (O_425,N_19899,N_19613);
nand UO_426 (O_426,N_19704,N_19595);
or UO_427 (O_427,N_19990,N_19616);
nand UO_428 (O_428,N_19638,N_19932);
nand UO_429 (O_429,N_19556,N_19618);
nor UO_430 (O_430,N_19838,N_19813);
nand UO_431 (O_431,N_19729,N_19596);
nand UO_432 (O_432,N_19732,N_19505);
or UO_433 (O_433,N_19674,N_19690);
and UO_434 (O_434,N_19886,N_19794);
nor UO_435 (O_435,N_19778,N_19941);
and UO_436 (O_436,N_19567,N_19663);
and UO_437 (O_437,N_19728,N_19654);
nand UO_438 (O_438,N_19521,N_19804);
or UO_439 (O_439,N_19800,N_19792);
nor UO_440 (O_440,N_19811,N_19974);
nor UO_441 (O_441,N_19879,N_19844);
and UO_442 (O_442,N_19550,N_19646);
and UO_443 (O_443,N_19864,N_19614);
and UO_444 (O_444,N_19662,N_19963);
nand UO_445 (O_445,N_19962,N_19580);
nand UO_446 (O_446,N_19608,N_19872);
nand UO_447 (O_447,N_19898,N_19799);
and UO_448 (O_448,N_19996,N_19902);
and UO_449 (O_449,N_19830,N_19858);
nor UO_450 (O_450,N_19984,N_19773);
and UO_451 (O_451,N_19978,N_19660);
or UO_452 (O_452,N_19591,N_19826);
nand UO_453 (O_453,N_19592,N_19679);
and UO_454 (O_454,N_19835,N_19720);
and UO_455 (O_455,N_19834,N_19921);
and UO_456 (O_456,N_19583,N_19500);
nand UO_457 (O_457,N_19653,N_19611);
or UO_458 (O_458,N_19662,N_19722);
or UO_459 (O_459,N_19776,N_19850);
or UO_460 (O_460,N_19934,N_19678);
or UO_461 (O_461,N_19841,N_19961);
or UO_462 (O_462,N_19956,N_19758);
and UO_463 (O_463,N_19534,N_19963);
and UO_464 (O_464,N_19530,N_19622);
nor UO_465 (O_465,N_19625,N_19891);
or UO_466 (O_466,N_19997,N_19538);
nor UO_467 (O_467,N_19756,N_19636);
and UO_468 (O_468,N_19651,N_19657);
and UO_469 (O_469,N_19613,N_19677);
and UO_470 (O_470,N_19884,N_19674);
and UO_471 (O_471,N_19987,N_19832);
or UO_472 (O_472,N_19989,N_19617);
or UO_473 (O_473,N_19765,N_19778);
or UO_474 (O_474,N_19662,N_19867);
nand UO_475 (O_475,N_19507,N_19702);
nand UO_476 (O_476,N_19940,N_19591);
and UO_477 (O_477,N_19803,N_19812);
nand UO_478 (O_478,N_19833,N_19703);
and UO_479 (O_479,N_19841,N_19615);
or UO_480 (O_480,N_19517,N_19977);
nor UO_481 (O_481,N_19544,N_19909);
nand UO_482 (O_482,N_19961,N_19744);
or UO_483 (O_483,N_19804,N_19793);
nand UO_484 (O_484,N_19881,N_19868);
nor UO_485 (O_485,N_19827,N_19617);
nand UO_486 (O_486,N_19750,N_19640);
and UO_487 (O_487,N_19646,N_19705);
or UO_488 (O_488,N_19643,N_19937);
and UO_489 (O_489,N_19981,N_19948);
nor UO_490 (O_490,N_19518,N_19656);
xor UO_491 (O_491,N_19823,N_19838);
or UO_492 (O_492,N_19652,N_19776);
nor UO_493 (O_493,N_19571,N_19560);
and UO_494 (O_494,N_19599,N_19613);
and UO_495 (O_495,N_19888,N_19981);
or UO_496 (O_496,N_19517,N_19762);
and UO_497 (O_497,N_19740,N_19931);
nor UO_498 (O_498,N_19653,N_19780);
nand UO_499 (O_499,N_19678,N_19849);
or UO_500 (O_500,N_19829,N_19611);
and UO_501 (O_501,N_19845,N_19871);
or UO_502 (O_502,N_19741,N_19675);
and UO_503 (O_503,N_19875,N_19536);
xor UO_504 (O_504,N_19968,N_19561);
and UO_505 (O_505,N_19843,N_19802);
or UO_506 (O_506,N_19987,N_19972);
nor UO_507 (O_507,N_19861,N_19957);
nor UO_508 (O_508,N_19704,N_19880);
and UO_509 (O_509,N_19741,N_19853);
and UO_510 (O_510,N_19590,N_19818);
or UO_511 (O_511,N_19841,N_19589);
or UO_512 (O_512,N_19789,N_19780);
or UO_513 (O_513,N_19671,N_19764);
or UO_514 (O_514,N_19595,N_19527);
nor UO_515 (O_515,N_19554,N_19760);
nand UO_516 (O_516,N_19566,N_19972);
and UO_517 (O_517,N_19655,N_19690);
nor UO_518 (O_518,N_19935,N_19859);
and UO_519 (O_519,N_19949,N_19807);
nand UO_520 (O_520,N_19908,N_19821);
and UO_521 (O_521,N_19547,N_19609);
and UO_522 (O_522,N_19681,N_19809);
and UO_523 (O_523,N_19546,N_19893);
and UO_524 (O_524,N_19594,N_19678);
or UO_525 (O_525,N_19783,N_19742);
or UO_526 (O_526,N_19937,N_19790);
and UO_527 (O_527,N_19765,N_19871);
xor UO_528 (O_528,N_19852,N_19978);
or UO_529 (O_529,N_19844,N_19951);
nand UO_530 (O_530,N_19965,N_19769);
nand UO_531 (O_531,N_19998,N_19602);
nor UO_532 (O_532,N_19724,N_19706);
nand UO_533 (O_533,N_19828,N_19862);
nand UO_534 (O_534,N_19544,N_19528);
nand UO_535 (O_535,N_19963,N_19944);
and UO_536 (O_536,N_19729,N_19740);
nand UO_537 (O_537,N_19707,N_19963);
nor UO_538 (O_538,N_19925,N_19852);
nand UO_539 (O_539,N_19631,N_19887);
and UO_540 (O_540,N_19939,N_19695);
nand UO_541 (O_541,N_19999,N_19805);
or UO_542 (O_542,N_19519,N_19818);
or UO_543 (O_543,N_19690,N_19557);
nor UO_544 (O_544,N_19790,N_19895);
or UO_545 (O_545,N_19532,N_19664);
nand UO_546 (O_546,N_19840,N_19775);
and UO_547 (O_547,N_19562,N_19719);
nor UO_548 (O_548,N_19922,N_19618);
nand UO_549 (O_549,N_19755,N_19520);
nor UO_550 (O_550,N_19770,N_19868);
nor UO_551 (O_551,N_19955,N_19851);
nand UO_552 (O_552,N_19764,N_19995);
nand UO_553 (O_553,N_19767,N_19693);
nand UO_554 (O_554,N_19810,N_19909);
nand UO_555 (O_555,N_19983,N_19727);
or UO_556 (O_556,N_19792,N_19509);
or UO_557 (O_557,N_19581,N_19538);
nor UO_558 (O_558,N_19706,N_19510);
nand UO_559 (O_559,N_19914,N_19681);
or UO_560 (O_560,N_19845,N_19582);
and UO_561 (O_561,N_19742,N_19739);
nand UO_562 (O_562,N_19621,N_19684);
nor UO_563 (O_563,N_19949,N_19511);
and UO_564 (O_564,N_19593,N_19601);
or UO_565 (O_565,N_19612,N_19779);
nor UO_566 (O_566,N_19911,N_19998);
or UO_567 (O_567,N_19663,N_19796);
nand UO_568 (O_568,N_19540,N_19954);
nor UO_569 (O_569,N_19610,N_19896);
and UO_570 (O_570,N_19634,N_19850);
or UO_571 (O_571,N_19559,N_19871);
and UO_572 (O_572,N_19706,N_19624);
and UO_573 (O_573,N_19684,N_19941);
or UO_574 (O_574,N_19898,N_19847);
nand UO_575 (O_575,N_19900,N_19923);
and UO_576 (O_576,N_19965,N_19533);
nor UO_577 (O_577,N_19844,N_19829);
and UO_578 (O_578,N_19930,N_19505);
nand UO_579 (O_579,N_19771,N_19616);
nand UO_580 (O_580,N_19811,N_19635);
and UO_581 (O_581,N_19582,N_19644);
or UO_582 (O_582,N_19559,N_19784);
nor UO_583 (O_583,N_19599,N_19945);
nor UO_584 (O_584,N_19808,N_19829);
nor UO_585 (O_585,N_19695,N_19889);
nand UO_586 (O_586,N_19807,N_19709);
and UO_587 (O_587,N_19600,N_19695);
or UO_588 (O_588,N_19601,N_19739);
nand UO_589 (O_589,N_19521,N_19564);
or UO_590 (O_590,N_19571,N_19942);
or UO_591 (O_591,N_19620,N_19808);
nand UO_592 (O_592,N_19640,N_19606);
or UO_593 (O_593,N_19780,N_19921);
and UO_594 (O_594,N_19898,N_19641);
nand UO_595 (O_595,N_19545,N_19512);
nor UO_596 (O_596,N_19783,N_19632);
or UO_597 (O_597,N_19994,N_19814);
and UO_598 (O_598,N_19620,N_19778);
or UO_599 (O_599,N_19753,N_19846);
and UO_600 (O_600,N_19849,N_19730);
nand UO_601 (O_601,N_19649,N_19939);
or UO_602 (O_602,N_19503,N_19921);
nor UO_603 (O_603,N_19906,N_19739);
or UO_604 (O_604,N_19854,N_19767);
nand UO_605 (O_605,N_19667,N_19814);
xnor UO_606 (O_606,N_19758,N_19939);
nand UO_607 (O_607,N_19517,N_19826);
and UO_608 (O_608,N_19840,N_19979);
nand UO_609 (O_609,N_19588,N_19710);
nor UO_610 (O_610,N_19966,N_19704);
nand UO_611 (O_611,N_19851,N_19633);
and UO_612 (O_612,N_19874,N_19706);
and UO_613 (O_613,N_19925,N_19689);
nand UO_614 (O_614,N_19859,N_19547);
or UO_615 (O_615,N_19808,N_19784);
and UO_616 (O_616,N_19799,N_19971);
or UO_617 (O_617,N_19870,N_19561);
and UO_618 (O_618,N_19715,N_19928);
or UO_619 (O_619,N_19793,N_19991);
and UO_620 (O_620,N_19850,N_19965);
nand UO_621 (O_621,N_19643,N_19646);
and UO_622 (O_622,N_19571,N_19995);
and UO_623 (O_623,N_19747,N_19787);
and UO_624 (O_624,N_19661,N_19907);
and UO_625 (O_625,N_19622,N_19869);
nor UO_626 (O_626,N_19974,N_19966);
and UO_627 (O_627,N_19981,N_19717);
or UO_628 (O_628,N_19535,N_19847);
or UO_629 (O_629,N_19848,N_19657);
and UO_630 (O_630,N_19595,N_19911);
nand UO_631 (O_631,N_19560,N_19777);
or UO_632 (O_632,N_19943,N_19780);
or UO_633 (O_633,N_19842,N_19746);
nand UO_634 (O_634,N_19800,N_19686);
nor UO_635 (O_635,N_19585,N_19717);
nand UO_636 (O_636,N_19587,N_19823);
and UO_637 (O_637,N_19833,N_19541);
nand UO_638 (O_638,N_19976,N_19902);
or UO_639 (O_639,N_19819,N_19824);
or UO_640 (O_640,N_19519,N_19764);
or UO_641 (O_641,N_19955,N_19904);
and UO_642 (O_642,N_19869,N_19589);
nand UO_643 (O_643,N_19683,N_19551);
nand UO_644 (O_644,N_19993,N_19630);
and UO_645 (O_645,N_19717,N_19999);
nand UO_646 (O_646,N_19718,N_19800);
nor UO_647 (O_647,N_19625,N_19552);
nor UO_648 (O_648,N_19943,N_19844);
and UO_649 (O_649,N_19602,N_19607);
nor UO_650 (O_650,N_19647,N_19906);
nor UO_651 (O_651,N_19641,N_19684);
or UO_652 (O_652,N_19661,N_19659);
or UO_653 (O_653,N_19543,N_19618);
nor UO_654 (O_654,N_19559,N_19825);
or UO_655 (O_655,N_19672,N_19539);
nor UO_656 (O_656,N_19529,N_19727);
or UO_657 (O_657,N_19601,N_19791);
nand UO_658 (O_658,N_19698,N_19954);
nand UO_659 (O_659,N_19700,N_19557);
and UO_660 (O_660,N_19516,N_19753);
nor UO_661 (O_661,N_19553,N_19849);
nor UO_662 (O_662,N_19714,N_19685);
and UO_663 (O_663,N_19615,N_19866);
nand UO_664 (O_664,N_19586,N_19676);
or UO_665 (O_665,N_19508,N_19842);
nand UO_666 (O_666,N_19586,N_19519);
nor UO_667 (O_667,N_19908,N_19589);
and UO_668 (O_668,N_19719,N_19657);
or UO_669 (O_669,N_19527,N_19661);
or UO_670 (O_670,N_19540,N_19589);
nand UO_671 (O_671,N_19581,N_19662);
nand UO_672 (O_672,N_19736,N_19678);
or UO_673 (O_673,N_19709,N_19763);
nor UO_674 (O_674,N_19562,N_19902);
and UO_675 (O_675,N_19725,N_19916);
nor UO_676 (O_676,N_19995,N_19601);
and UO_677 (O_677,N_19542,N_19736);
nand UO_678 (O_678,N_19604,N_19975);
or UO_679 (O_679,N_19822,N_19730);
or UO_680 (O_680,N_19540,N_19712);
or UO_681 (O_681,N_19935,N_19972);
and UO_682 (O_682,N_19815,N_19692);
nand UO_683 (O_683,N_19781,N_19609);
nand UO_684 (O_684,N_19816,N_19544);
nand UO_685 (O_685,N_19729,N_19997);
nand UO_686 (O_686,N_19671,N_19506);
or UO_687 (O_687,N_19869,N_19569);
nor UO_688 (O_688,N_19548,N_19576);
or UO_689 (O_689,N_19529,N_19548);
nor UO_690 (O_690,N_19783,N_19514);
nor UO_691 (O_691,N_19595,N_19721);
or UO_692 (O_692,N_19687,N_19717);
nand UO_693 (O_693,N_19793,N_19822);
nand UO_694 (O_694,N_19901,N_19646);
nor UO_695 (O_695,N_19777,N_19598);
nor UO_696 (O_696,N_19992,N_19929);
nand UO_697 (O_697,N_19898,N_19553);
nor UO_698 (O_698,N_19590,N_19982);
and UO_699 (O_699,N_19951,N_19721);
nor UO_700 (O_700,N_19899,N_19771);
nand UO_701 (O_701,N_19575,N_19749);
or UO_702 (O_702,N_19697,N_19602);
nand UO_703 (O_703,N_19556,N_19666);
nand UO_704 (O_704,N_19785,N_19556);
nor UO_705 (O_705,N_19677,N_19671);
and UO_706 (O_706,N_19632,N_19562);
and UO_707 (O_707,N_19873,N_19793);
nor UO_708 (O_708,N_19539,N_19749);
and UO_709 (O_709,N_19729,N_19672);
nand UO_710 (O_710,N_19682,N_19721);
xor UO_711 (O_711,N_19986,N_19858);
or UO_712 (O_712,N_19755,N_19853);
nor UO_713 (O_713,N_19772,N_19928);
nor UO_714 (O_714,N_19717,N_19718);
or UO_715 (O_715,N_19980,N_19930);
nand UO_716 (O_716,N_19746,N_19982);
nor UO_717 (O_717,N_19553,N_19688);
nor UO_718 (O_718,N_19702,N_19820);
and UO_719 (O_719,N_19889,N_19905);
and UO_720 (O_720,N_19905,N_19559);
or UO_721 (O_721,N_19578,N_19877);
nor UO_722 (O_722,N_19855,N_19960);
nor UO_723 (O_723,N_19533,N_19704);
or UO_724 (O_724,N_19596,N_19543);
or UO_725 (O_725,N_19682,N_19800);
nand UO_726 (O_726,N_19800,N_19855);
and UO_727 (O_727,N_19777,N_19747);
and UO_728 (O_728,N_19756,N_19779);
nand UO_729 (O_729,N_19794,N_19700);
nor UO_730 (O_730,N_19861,N_19506);
nand UO_731 (O_731,N_19966,N_19764);
or UO_732 (O_732,N_19565,N_19912);
or UO_733 (O_733,N_19964,N_19559);
or UO_734 (O_734,N_19545,N_19522);
xnor UO_735 (O_735,N_19762,N_19505);
or UO_736 (O_736,N_19857,N_19513);
or UO_737 (O_737,N_19643,N_19909);
or UO_738 (O_738,N_19639,N_19617);
nor UO_739 (O_739,N_19939,N_19887);
nand UO_740 (O_740,N_19602,N_19582);
nor UO_741 (O_741,N_19791,N_19953);
nor UO_742 (O_742,N_19616,N_19784);
or UO_743 (O_743,N_19602,N_19614);
nor UO_744 (O_744,N_19618,N_19969);
nor UO_745 (O_745,N_19951,N_19881);
nand UO_746 (O_746,N_19762,N_19860);
or UO_747 (O_747,N_19875,N_19786);
or UO_748 (O_748,N_19542,N_19931);
and UO_749 (O_749,N_19515,N_19507);
or UO_750 (O_750,N_19671,N_19844);
nand UO_751 (O_751,N_19870,N_19797);
and UO_752 (O_752,N_19737,N_19916);
nand UO_753 (O_753,N_19855,N_19726);
nor UO_754 (O_754,N_19649,N_19633);
or UO_755 (O_755,N_19861,N_19842);
nand UO_756 (O_756,N_19776,N_19557);
nor UO_757 (O_757,N_19835,N_19551);
nand UO_758 (O_758,N_19616,N_19799);
nor UO_759 (O_759,N_19977,N_19767);
and UO_760 (O_760,N_19519,N_19668);
and UO_761 (O_761,N_19889,N_19677);
nand UO_762 (O_762,N_19511,N_19578);
nand UO_763 (O_763,N_19546,N_19959);
nor UO_764 (O_764,N_19838,N_19923);
nor UO_765 (O_765,N_19617,N_19893);
and UO_766 (O_766,N_19750,N_19673);
or UO_767 (O_767,N_19703,N_19901);
nor UO_768 (O_768,N_19686,N_19581);
or UO_769 (O_769,N_19771,N_19748);
and UO_770 (O_770,N_19948,N_19564);
nand UO_771 (O_771,N_19516,N_19860);
and UO_772 (O_772,N_19582,N_19726);
and UO_773 (O_773,N_19738,N_19789);
nor UO_774 (O_774,N_19660,N_19891);
nand UO_775 (O_775,N_19862,N_19978);
nor UO_776 (O_776,N_19659,N_19982);
nand UO_777 (O_777,N_19802,N_19571);
and UO_778 (O_778,N_19670,N_19809);
nand UO_779 (O_779,N_19859,N_19646);
or UO_780 (O_780,N_19601,N_19948);
and UO_781 (O_781,N_19994,N_19586);
and UO_782 (O_782,N_19500,N_19925);
nand UO_783 (O_783,N_19897,N_19967);
or UO_784 (O_784,N_19780,N_19742);
nor UO_785 (O_785,N_19736,N_19670);
nor UO_786 (O_786,N_19858,N_19813);
nand UO_787 (O_787,N_19664,N_19827);
nor UO_788 (O_788,N_19732,N_19867);
or UO_789 (O_789,N_19694,N_19687);
or UO_790 (O_790,N_19519,N_19939);
nor UO_791 (O_791,N_19573,N_19889);
nor UO_792 (O_792,N_19926,N_19923);
or UO_793 (O_793,N_19657,N_19773);
nand UO_794 (O_794,N_19671,N_19769);
nor UO_795 (O_795,N_19555,N_19554);
nor UO_796 (O_796,N_19866,N_19781);
or UO_797 (O_797,N_19975,N_19641);
and UO_798 (O_798,N_19735,N_19824);
or UO_799 (O_799,N_19981,N_19774);
and UO_800 (O_800,N_19976,N_19892);
and UO_801 (O_801,N_19784,N_19504);
and UO_802 (O_802,N_19683,N_19605);
nand UO_803 (O_803,N_19870,N_19791);
nor UO_804 (O_804,N_19765,N_19716);
and UO_805 (O_805,N_19993,N_19877);
nor UO_806 (O_806,N_19597,N_19767);
nor UO_807 (O_807,N_19577,N_19766);
or UO_808 (O_808,N_19873,N_19606);
and UO_809 (O_809,N_19641,N_19835);
and UO_810 (O_810,N_19673,N_19600);
and UO_811 (O_811,N_19867,N_19902);
nand UO_812 (O_812,N_19855,N_19887);
nand UO_813 (O_813,N_19884,N_19897);
or UO_814 (O_814,N_19609,N_19554);
and UO_815 (O_815,N_19867,N_19901);
nand UO_816 (O_816,N_19953,N_19738);
and UO_817 (O_817,N_19831,N_19643);
and UO_818 (O_818,N_19818,N_19651);
and UO_819 (O_819,N_19875,N_19542);
or UO_820 (O_820,N_19791,N_19542);
or UO_821 (O_821,N_19866,N_19503);
and UO_822 (O_822,N_19900,N_19589);
nor UO_823 (O_823,N_19949,N_19568);
nor UO_824 (O_824,N_19519,N_19921);
nand UO_825 (O_825,N_19807,N_19971);
nor UO_826 (O_826,N_19774,N_19697);
or UO_827 (O_827,N_19881,N_19807);
and UO_828 (O_828,N_19860,N_19742);
nand UO_829 (O_829,N_19870,N_19722);
nand UO_830 (O_830,N_19595,N_19535);
nand UO_831 (O_831,N_19970,N_19559);
nand UO_832 (O_832,N_19782,N_19916);
and UO_833 (O_833,N_19815,N_19568);
or UO_834 (O_834,N_19639,N_19527);
nor UO_835 (O_835,N_19791,N_19683);
and UO_836 (O_836,N_19879,N_19596);
and UO_837 (O_837,N_19522,N_19898);
nor UO_838 (O_838,N_19792,N_19840);
nand UO_839 (O_839,N_19811,N_19873);
xor UO_840 (O_840,N_19742,N_19812);
or UO_841 (O_841,N_19655,N_19761);
or UO_842 (O_842,N_19727,N_19505);
or UO_843 (O_843,N_19571,N_19607);
nor UO_844 (O_844,N_19903,N_19872);
and UO_845 (O_845,N_19732,N_19628);
nor UO_846 (O_846,N_19960,N_19780);
or UO_847 (O_847,N_19720,N_19642);
nor UO_848 (O_848,N_19865,N_19974);
nor UO_849 (O_849,N_19509,N_19692);
and UO_850 (O_850,N_19802,N_19702);
and UO_851 (O_851,N_19571,N_19864);
or UO_852 (O_852,N_19614,N_19588);
nand UO_853 (O_853,N_19823,N_19578);
or UO_854 (O_854,N_19755,N_19941);
nand UO_855 (O_855,N_19623,N_19584);
and UO_856 (O_856,N_19896,N_19744);
or UO_857 (O_857,N_19836,N_19872);
or UO_858 (O_858,N_19931,N_19801);
nand UO_859 (O_859,N_19810,N_19863);
and UO_860 (O_860,N_19604,N_19836);
and UO_861 (O_861,N_19509,N_19550);
and UO_862 (O_862,N_19981,N_19579);
or UO_863 (O_863,N_19520,N_19933);
and UO_864 (O_864,N_19571,N_19504);
or UO_865 (O_865,N_19711,N_19989);
nor UO_866 (O_866,N_19685,N_19946);
or UO_867 (O_867,N_19721,N_19800);
and UO_868 (O_868,N_19668,N_19900);
nand UO_869 (O_869,N_19734,N_19889);
nor UO_870 (O_870,N_19922,N_19927);
or UO_871 (O_871,N_19695,N_19675);
or UO_872 (O_872,N_19548,N_19675);
nand UO_873 (O_873,N_19598,N_19732);
nor UO_874 (O_874,N_19693,N_19982);
and UO_875 (O_875,N_19738,N_19620);
and UO_876 (O_876,N_19919,N_19893);
nand UO_877 (O_877,N_19779,N_19958);
nor UO_878 (O_878,N_19785,N_19987);
nand UO_879 (O_879,N_19923,N_19839);
nor UO_880 (O_880,N_19635,N_19995);
or UO_881 (O_881,N_19788,N_19781);
nand UO_882 (O_882,N_19637,N_19625);
and UO_883 (O_883,N_19827,N_19531);
or UO_884 (O_884,N_19864,N_19996);
and UO_885 (O_885,N_19614,N_19545);
nor UO_886 (O_886,N_19812,N_19784);
nand UO_887 (O_887,N_19981,N_19512);
nor UO_888 (O_888,N_19601,N_19781);
nor UO_889 (O_889,N_19835,N_19980);
and UO_890 (O_890,N_19517,N_19664);
nand UO_891 (O_891,N_19754,N_19979);
nand UO_892 (O_892,N_19765,N_19605);
nand UO_893 (O_893,N_19691,N_19885);
xor UO_894 (O_894,N_19845,N_19515);
and UO_895 (O_895,N_19800,N_19713);
nor UO_896 (O_896,N_19581,N_19909);
xnor UO_897 (O_897,N_19934,N_19521);
or UO_898 (O_898,N_19953,N_19990);
or UO_899 (O_899,N_19627,N_19563);
nor UO_900 (O_900,N_19861,N_19865);
nand UO_901 (O_901,N_19646,N_19592);
nand UO_902 (O_902,N_19579,N_19940);
nand UO_903 (O_903,N_19759,N_19779);
nand UO_904 (O_904,N_19960,N_19763);
nand UO_905 (O_905,N_19910,N_19881);
or UO_906 (O_906,N_19625,N_19897);
and UO_907 (O_907,N_19857,N_19728);
nand UO_908 (O_908,N_19555,N_19619);
nand UO_909 (O_909,N_19865,N_19989);
and UO_910 (O_910,N_19565,N_19979);
nand UO_911 (O_911,N_19644,N_19941);
and UO_912 (O_912,N_19683,N_19648);
and UO_913 (O_913,N_19601,N_19520);
or UO_914 (O_914,N_19862,N_19592);
nand UO_915 (O_915,N_19615,N_19585);
and UO_916 (O_916,N_19843,N_19943);
nand UO_917 (O_917,N_19938,N_19999);
nor UO_918 (O_918,N_19522,N_19798);
nand UO_919 (O_919,N_19945,N_19649);
and UO_920 (O_920,N_19668,N_19508);
nand UO_921 (O_921,N_19750,N_19765);
and UO_922 (O_922,N_19519,N_19958);
and UO_923 (O_923,N_19984,N_19978);
or UO_924 (O_924,N_19627,N_19782);
nand UO_925 (O_925,N_19762,N_19908);
nor UO_926 (O_926,N_19820,N_19785);
and UO_927 (O_927,N_19516,N_19680);
and UO_928 (O_928,N_19778,N_19798);
and UO_929 (O_929,N_19751,N_19841);
nor UO_930 (O_930,N_19727,N_19763);
nand UO_931 (O_931,N_19918,N_19739);
or UO_932 (O_932,N_19922,N_19635);
nand UO_933 (O_933,N_19618,N_19694);
nand UO_934 (O_934,N_19829,N_19503);
and UO_935 (O_935,N_19829,N_19890);
and UO_936 (O_936,N_19640,N_19678);
nor UO_937 (O_937,N_19684,N_19531);
or UO_938 (O_938,N_19544,N_19993);
nor UO_939 (O_939,N_19747,N_19557);
and UO_940 (O_940,N_19605,N_19587);
and UO_941 (O_941,N_19789,N_19552);
nand UO_942 (O_942,N_19714,N_19690);
and UO_943 (O_943,N_19995,N_19688);
nor UO_944 (O_944,N_19534,N_19624);
nor UO_945 (O_945,N_19860,N_19870);
and UO_946 (O_946,N_19626,N_19743);
xnor UO_947 (O_947,N_19956,N_19672);
and UO_948 (O_948,N_19901,N_19796);
nor UO_949 (O_949,N_19515,N_19764);
nor UO_950 (O_950,N_19744,N_19656);
and UO_951 (O_951,N_19991,N_19553);
nand UO_952 (O_952,N_19869,N_19715);
nand UO_953 (O_953,N_19670,N_19536);
or UO_954 (O_954,N_19726,N_19994);
nand UO_955 (O_955,N_19663,N_19545);
nand UO_956 (O_956,N_19677,N_19966);
nand UO_957 (O_957,N_19857,N_19946);
and UO_958 (O_958,N_19766,N_19820);
nand UO_959 (O_959,N_19747,N_19968);
nor UO_960 (O_960,N_19733,N_19689);
nor UO_961 (O_961,N_19564,N_19528);
and UO_962 (O_962,N_19932,N_19843);
nor UO_963 (O_963,N_19799,N_19882);
nand UO_964 (O_964,N_19501,N_19543);
or UO_965 (O_965,N_19677,N_19515);
and UO_966 (O_966,N_19854,N_19739);
or UO_967 (O_967,N_19515,N_19918);
or UO_968 (O_968,N_19816,N_19584);
or UO_969 (O_969,N_19777,N_19595);
nor UO_970 (O_970,N_19553,N_19759);
nand UO_971 (O_971,N_19975,N_19617);
xor UO_972 (O_972,N_19808,N_19597);
or UO_973 (O_973,N_19509,N_19675);
nor UO_974 (O_974,N_19969,N_19801);
and UO_975 (O_975,N_19618,N_19779);
or UO_976 (O_976,N_19926,N_19909);
and UO_977 (O_977,N_19769,N_19859);
nand UO_978 (O_978,N_19693,N_19624);
and UO_979 (O_979,N_19669,N_19618);
nor UO_980 (O_980,N_19805,N_19998);
or UO_981 (O_981,N_19800,N_19719);
or UO_982 (O_982,N_19882,N_19871);
nand UO_983 (O_983,N_19700,N_19518);
nand UO_984 (O_984,N_19906,N_19693);
or UO_985 (O_985,N_19612,N_19753);
nand UO_986 (O_986,N_19801,N_19843);
nand UO_987 (O_987,N_19769,N_19685);
or UO_988 (O_988,N_19852,N_19699);
nand UO_989 (O_989,N_19749,N_19950);
or UO_990 (O_990,N_19789,N_19510);
nor UO_991 (O_991,N_19853,N_19815);
or UO_992 (O_992,N_19847,N_19892);
nand UO_993 (O_993,N_19540,N_19965);
or UO_994 (O_994,N_19807,N_19672);
and UO_995 (O_995,N_19502,N_19661);
nor UO_996 (O_996,N_19748,N_19709);
and UO_997 (O_997,N_19988,N_19693);
and UO_998 (O_998,N_19828,N_19782);
and UO_999 (O_999,N_19899,N_19759);
nand UO_1000 (O_1000,N_19790,N_19955);
nor UO_1001 (O_1001,N_19989,N_19584);
nand UO_1002 (O_1002,N_19936,N_19870);
nand UO_1003 (O_1003,N_19506,N_19932);
nand UO_1004 (O_1004,N_19749,N_19597);
nand UO_1005 (O_1005,N_19793,N_19583);
and UO_1006 (O_1006,N_19770,N_19880);
nor UO_1007 (O_1007,N_19593,N_19746);
nor UO_1008 (O_1008,N_19842,N_19822);
and UO_1009 (O_1009,N_19774,N_19929);
xnor UO_1010 (O_1010,N_19526,N_19868);
nand UO_1011 (O_1011,N_19571,N_19634);
or UO_1012 (O_1012,N_19741,N_19565);
or UO_1013 (O_1013,N_19899,N_19894);
and UO_1014 (O_1014,N_19964,N_19990);
nor UO_1015 (O_1015,N_19824,N_19981);
or UO_1016 (O_1016,N_19969,N_19569);
or UO_1017 (O_1017,N_19700,N_19582);
nor UO_1018 (O_1018,N_19534,N_19925);
xnor UO_1019 (O_1019,N_19572,N_19672);
and UO_1020 (O_1020,N_19721,N_19652);
or UO_1021 (O_1021,N_19869,N_19603);
nor UO_1022 (O_1022,N_19602,N_19675);
or UO_1023 (O_1023,N_19641,N_19604);
or UO_1024 (O_1024,N_19647,N_19634);
nor UO_1025 (O_1025,N_19600,N_19955);
or UO_1026 (O_1026,N_19569,N_19799);
and UO_1027 (O_1027,N_19791,N_19980);
and UO_1028 (O_1028,N_19546,N_19698);
nand UO_1029 (O_1029,N_19951,N_19811);
nor UO_1030 (O_1030,N_19644,N_19861);
or UO_1031 (O_1031,N_19664,N_19630);
xor UO_1032 (O_1032,N_19667,N_19788);
and UO_1033 (O_1033,N_19503,N_19959);
and UO_1034 (O_1034,N_19540,N_19662);
and UO_1035 (O_1035,N_19660,N_19841);
and UO_1036 (O_1036,N_19787,N_19742);
nor UO_1037 (O_1037,N_19662,N_19538);
nand UO_1038 (O_1038,N_19862,N_19747);
or UO_1039 (O_1039,N_19785,N_19851);
or UO_1040 (O_1040,N_19872,N_19575);
nand UO_1041 (O_1041,N_19957,N_19608);
nand UO_1042 (O_1042,N_19665,N_19813);
or UO_1043 (O_1043,N_19884,N_19698);
xor UO_1044 (O_1044,N_19951,N_19916);
nor UO_1045 (O_1045,N_19513,N_19961);
or UO_1046 (O_1046,N_19752,N_19822);
and UO_1047 (O_1047,N_19796,N_19596);
nand UO_1048 (O_1048,N_19655,N_19671);
or UO_1049 (O_1049,N_19695,N_19561);
and UO_1050 (O_1050,N_19969,N_19671);
or UO_1051 (O_1051,N_19513,N_19770);
nor UO_1052 (O_1052,N_19573,N_19846);
and UO_1053 (O_1053,N_19924,N_19666);
nand UO_1054 (O_1054,N_19874,N_19888);
or UO_1055 (O_1055,N_19728,N_19851);
nor UO_1056 (O_1056,N_19514,N_19959);
xnor UO_1057 (O_1057,N_19680,N_19953);
nand UO_1058 (O_1058,N_19518,N_19729);
nor UO_1059 (O_1059,N_19906,N_19713);
nand UO_1060 (O_1060,N_19832,N_19547);
nand UO_1061 (O_1061,N_19910,N_19859);
and UO_1062 (O_1062,N_19586,N_19863);
or UO_1063 (O_1063,N_19585,N_19721);
and UO_1064 (O_1064,N_19662,N_19852);
and UO_1065 (O_1065,N_19641,N_19671);
or UO_1066 (O_1066,N_19657,N_19560);
or UO_1067 (O_1067,N_19709,N_19796);
nand UO_1068 (O_1068,N_19631,N_19623);
nand UO_1069 (O_1069,N_19776,N_19825);
xnor UO_1070 (O_1070,N_19967,N_19922);
nor UO_1071 (O_1071,N_19978,N_19956);
and UO_1072 (O_1072,N_19507,N_19837);
and UO_1073 (O_1073,N_19847,N_19991);
or UO_1074 (O_1074,N_19630,N_19720);
or UO_1075 (O_1075,N_19645,N_19641);
or UO_1076 (O_1076,N_19826,N_19910);
nor UO_1077 (O_1077,N_19559,N_19854);
and UO_1078 (O_1078,N_19794,N_19774);
nand UO_1079 (O_1079,N_19996,N_19852);
nand UO_1080 (O_1080,N_19994,N_19977);
nor UO_1081 (O_1081,N_19644,N_19586);
or UO_1082 (O_1082,N_19942,N_19542);
and UO_1083 (O_1083,N_19879,N_19861);
nand UO_1084 (O_1084,N_19645,N_19909);
nand UO_1085 (O_1085,N_19782,N_19970);
nand UO_1086 (O_1086,N_19556,N_19737);
nor UO_1087 (O_1087,N_19782,N_19842);
nor UO_1088 (O_1088,N_19736,N_19738);
and UO_1089 (O_1089,N_19740,N_19517);
nand UO_1090 (O_1090,N_19977,N_19844);
or UO_1091 (O_1091,N_19886,N_19619);
or UO_1092 (O_1092,N_19858,N_19637);
or UO_1093 (O_1093,N_19684,N_19897);
and UO_1094 (O_1094,N_19941,N_19788);
or UO_1095 (O_1095,N_19770,N_19515);
or UO_1096 (O_1096,N_19574,N_19851);
nor UO_1097 (O_1097,N_19698,N_19810);
nand UO_1098 (O_1098,N_19742,N_19990);
nor UO_1099 (O_1099,N_19975,N_19678);
or UO_1100 (O_1100,N_19698,N_19603);
and UO_1101 (O_1101,N_19607,N_19968);
and UO_1102 (O_1102,N_19875,N_19883);
nand UO_1103 (O_1103,N_19821,N_19635);
and UO_1104 (O_1104,N_19643,N_19980);
nor UO_1105 (O_1105,N_19846,N_19843);
nor UO_1106 (O_1106,N_19712,N_19747);
nand UO_1107 (O_1107,N_19906,N_19585);
or UO_1108 (O_1108,N_19951,N_19958);
or UO_1109 (O_1109,N_19977,N_19765);
or UO_1110 (O_1110,N_19805,N_19690);
xor UO_1111 (O_1111,N_19632,N_19854);
nor UO_1112 (O_1112,N_19996,N_19889);
nor UO_1113 (O_1113,N_19638,N_19642);
and UO_1114 (O_1114,N_19924,N_19510);
and UO_1115 (O_1115,N_19574,N_19980);
and UO_1116 (O_1116,N_19661,N_19882);
nor UO_1117 (O_1117,N_19804,N_19871);
and UO_1118 (O_1118,N_19655,N_19823);
and UO_1119 (O_1119,N_19639,N_19985);
nor UO_1120 (O_1120,N_19793,N_19759);
and UO_1121 (O_1121,N_19581,N_19582);
or UO_1122 (O_1122,N_19637,N_19704);
or UO_1123 (O_1123,N_19900,N_19669);
nand UO_1124 (O_1124,N_19782,N_19836);
nor UO_1125 (O_1125,N_19647,N_19787);
nand UO_1126 (O_1126,N_19818,N_19831);
or UO_1127 (O_1127,N_19941,N_19577);
nand UO_1128 (O_1128,N_19669,N_19604);
nor UO_1129 (O_1129,N_19948,N_19990);
and UO_1130 (O_1130,N_19767,N_19885);
or UO_1131 (O_1131,N_19957,N_19591);
nand UO_1132 (O_1132,N_19992,N_19517);
nor UO_1133 (O_1133,N_19556,N_19608);
and UO_1134 (O_1134,N_19524,N_19601);
or UO_1135 (O_1135,N_19985,N_19717);
and UO_1136 (O_1136,N_19709,N_19701);
nand UO_1137 (O_1137,N_19677,N_19917);
nand UO_1138 (O_1138,N_19520,N_19848);
and UO_1139 (O_1139,N_19608,N_19947);
or UO_1140 (O_1140,N_19507,N_19926);
nand UO_1141 (O_1141,N_19788,N_19915);
nand UO_1142 (O_1142,N_19909,N_19570);
or UO_1143 (O_1143,N_19528,N_19754);
nand UO_1144 (O_1144,N_19671,N_19539);
nor UO_1145 (O_1145,N_19720,N_19898);
nor UO_1146 (O_1146,N_19820,N_19594);
or UO_1147 (O_1147,N_19631,N_19856);
and UO_1148 (O_1148,N_19512,N_19573);
and UO_1149 (O_1149,N_19679,N_19628);
nor UO_1150 (O_1150,N_19900,N_19852);
or UO_1151 (O_1151,N_19860,N_19631);
xor UO_1152 (O_1152,N_19785,N_19776);
and UO_1153 (O_1153,N_19986,N_19827);
nor UO_1154 (O_1154,N_19913,N_19946);
and UO_1155 (O_1155,N_19729,N_19870);
nor UO_1156 (O_1156,N_19859,N_19722);
nand UO_1157 (O_1157,N_19807,N_19713);
nand UO_1158 (O_1158,N_19529,N_19692);
and UO_1159 (O_1159,N_19698,N_19500);
nand UO_1160 (O_1160,N_19840,N_19816);
and UO_1161 (O_1161,N_19501,N_19526);
nor UO_1162 (O_1162,N_19699,N_19612);
or UO_1163 (O_1163,N_19529,N_19795);
and UO_1164 (O_1164,N_19976,N_19616);
and UO_1165 (O_1165,N_19845,N_19620);
or UO_1166 (O_1166,N_19819,N_19562);
and UO_1167 (O_1167,N_19999,N_19534);
or UO_1168 (O_1168,N_19999,N_19623);
and UO_1169 (O_1169,N_19877,N_19873);
and UO_1170 (O_1170,N_19948,N_19684);
nor UO_1171 (O_1171,N_19614,N_19838);
and UO_1172 (O_1172,N_19567,N_19808);
nand UO_1173 (O_1173,N_19802,N_19983);
or UO_1174 (O_1174,N_19971,N_19763);
nand UO_1175 (O_1175,N_19790,N_19907);
or UO_1176 (O_1176,N_19533,N_19560);
nand UO_1177 (O_1177,N_19784,N_19900);
nand UO_1178 (O_1178,N_19550,N_19960);
and UO_1179 (O_1179,N_19824,N_19592);
or UO_1180 (O_1180,N_19666,N_19535);
nor UO_1181 (O_1181,N_19709,N_19872);
nor UO_1182 (O_1182,N_19936,N_19856);
nand UO_1183 (O_1183,N_19950,N_19893);
and UO_1184 (O_1184,N_19538,N_19825);
nand UO_1185 (O_1185,N_19582,N_19783);
or UO_1186 (O_1186,N_19953,N_19814);
xnor UO_1187 (O_1187,N_19600,N_19710);
nand UO_1188 (O_1188,N_19816,N_19731);
and UO_1189 (O_1189,N_19621,N_19557);
and UO_1190 (O_1190,N_19744,N_19536);
nor UO_1191 (O_1191,N_19964,N_19575);
nor UO_1192 (O_1192,N_19984,N_19625);
nand UO_1193 (O_1193,N_19608,N_19675);
nor UO_1194 (O_1194,N_19689,N_19840);
nor UO_1195 (O_1195,N_19784,N_19758);
and UO_1196 (O_1196,N_19745,N_19894);
nand UO_1197 (O_1197,N_19540,N_19795);
nand UO_1198 (O_1198,N_19731,N_19990);
nand UO_1199 (O_1199,N_19545,N_19555);
nor UO_1200 (O_1200,N_19731,N_19670);
nand UO_1201 (O_1201,N_19700,N_19604);
or UO_1202 (O_1202,N_19744,N_19693);
nand UO_1203 (O_1203,N_19621,N_19967);
or UO_1204 (O_1204,N_19816,N_19841);
or UO_1205 (O_1205,N_19824,N_19601);
and UO_1206 (O_1206,N_19525,N_19927);
and UO_1207 (O_1207,N_19801,N_19828);
or UO_1208 (O_1208,N_19869,N_19988);
nor UO_1209 (O_1209,N_19841,N_19696);
and UO_1210 (O_1210,N_19894,N_19764);
and UO_1211 (O_1211,N_19509,N_19798);
or UO_1212 (O_1212,N_19873,N_19580);
nor UO_1213 (O_1213,N_19865,N_19901);
nand UO_1214 (O_1214,N_19741,N_19554);
and UO_1215 (O_1215,N_19554,N_19531);
nand UO_1216 (O_1216,N_19600,N_19566);
and UO_1217 (O_1217,N_19588,N_19758);
nor UO_1218 (O_1218,N_19741,N_19713);
or UO_1219 (O_1219,N_19779,N_19800);
or UO_1220 (O_1220,N_19831,N_19763);
and UO_1221 (O_1221,N_19696,N_19948);
and UO_1222 (O_1222,N_19637,N_19684);
nand UO_1223 (O_1223,N_19797,N_19538);
and UO_1224 (O_1224,N_19568,N_19813);
or UO_1225 (O_1225,N_19957,N_19982);
and UO_1226 (O_1226,N_19501,N_19995);
nand UO_1227 (O_1227,N_19560,N_19861);
or UO_1228 (O_1228,N_19990,N_19913);
or UO_1229 (O_1229,N_19522,N_19650);
nor UO_1230 (O_1230,N_19649,N_19895);
nand UO_1231 (O_1231,N_19796,N_19941);
or UO_1232 (O_1232,N_19729,N_19837);
nand UO_1233 (O_1233,N_19795,N_19576);
nand UO_1234 (O_1234,N_19585,N_19669);
nor UO_1235 (O_1235,N_19699,N_19807);
nor UO_1236 (O_1236,N_19569,N_19976);
nor UO_1237 (O_1237,N_19617,N_19612);
nand UO_1238 (O_1238,N_19897,N_19724);
and UO_1239 (O_1239,N_19835,N_19832);
or UO_1240 (O_1240,N_19795,N_19881);
nand UO_1241 (O_1241,N_19950,N_19606);
or UO_1242 (O_1242,N_19991,N_19714);
nand UO_1243 (O_1243,N_19859,N_19731);
nor UO_1244 (O_1244,N_19584,N_19565);
nor UO_1245 (O_1245,N_19764,N_19511);
nand UO_1246 (O_1246,N_19663,N_19695);
nor UO_1247 (O_1247,N_19974,N_19888);
nand UO_1248 (O_1248,N_19571,N_19889);
nand UO_1249 (O_1249,N_19656,N_19553);
and UO_1250 (O_1250,N_19726,N_19644);
nor UO_1251 (O_1251,N_19560,N_19691);
nor UO_1252 (O_1252,N_19601,N_19834);
or UO_1253 (O_1253,N_19838,N_19618);
xor UO_1254 (O_1254,N_19817,N_19920);
nor UO_1255 (O_1255,N_19686,N_19691);
and UO_1256 (O_1256,N_19620,N_19837);
or UO_1257 (O_1257,N_19556,N_19949);
or UO_1258 (O_1258,N_19846,N_19895);
nand UO_1259 (O_1259,N_19965,N_19557);
nand UO_1260 (O_1260,N_19962,N_19863);
and UO_1261 (O_1261,N_19648,N_19769);
and UO_1262 (O_1262,N_19666,N_19730);
or UO_1263 (O_1263,N_19566,N_19678);
nor UO_1264 (O_1264,N_19877,N_19964);
or UO_1265 (O_1265,N_19564,N_19763);
nor UO_1266 (O_1266,N_19600,N_19698);
and UO_1267 (O_1267,N_19931,N_19993);
and UO_1268 (O_1268,N_19541,N_19603);
nand UO_1269 (O_1269,N_19792,N_19926);
or UO_1270 (O_1270,N_19678,N_19584);
and UO_1271 (O_1271,N_19684,N_19646);
nor UO_1272 (O_1272,N_19668,N_19615);
nand UO_1273 (O_1273,N_19850,N_19814);
nor UO_1274 (O_1274,N_19578,N_19722);
nor UO_1275 (O_1275,N_19664,N_19665);
nand UO_1276 (O_1276,N_19890,N_19743);
nor UO_1277 (O_1277,N_19897,N_19851);
nand UO_1278 (O_1278,N_19730,N_19785);
and UO_1279 (O_1279,N_19978,N_19586);
nor UO_1280 (O_1280,N_19850,N_19856);
or UO_1281 (O_1281,N_19821,N_19952);
and UO_1282 (O_1282,N_19637,N_19875);
nor UO_1283 (O_1283,N_19954,N_19938);
and UO_1284 (O_1284,N_19942,N_19882);
nand UO_1285 (O_1285,N_19522,N_19983);
and UO_1286 (O_1286,N_19885,N_19785);
or UO_1287 (O_1287,N_19950,N_19551);
or UO_1288 (O_1288,N_19706,N_19546);
nand UO_1289 (O_1289,N_19523,N_19816);
nor UO_1290 (O_1290,N_19783,N_19987);
or UO_1291 (O_1291,N_19601,N_19827);
or UO_1292 (O_1292,N_19720,N_19757);
or UO_1293 (O_1293,N_19966,N_19862);
nor UO_1294 (O_1294,N_19604,N_19849);
or UO_1295 (O_1295,N_19967,N_19550);
or UO_1296 (O_1296,N_19770,N_19755);
nor UO_1297 (O_1297,N_19730,N_19904);
xor UO_1298 (O_1298,N_19603,N_19743);
and UO_1299 (O_1299,N_19640,N_19643);
or UO_1300 (O_1300,N_19559,N_19725);
or UO_1301 (O_1301,N_19959,N_19867);
and UO_1302 (O_1302,N_19649,N_19853);
or UO_1303 (O_1303,N_19832,N_19803);
nor UO_1304 (O_1304,N_19721,N_19597);
and UO_1305 (O_1305,N_19955,N_19897);
and UO_1306 (O_1306,N_19874,N_19980);
nor UO_1307 (O_1307,N_19808,N_19850);
and UO_1308 (O_1308,N_19749,N_19941);
nand UO_1309 (O_1309,N_19673,N_19870);
nand UO_1310 (O_1310,N_19729,N_19968);
xor UO_1311 (O_1311,N_19716,N_19998);
nor UO_1312 (O_1312,N_19856,N_19829);
and UO_1313 (O_1313,N_19896,N_19673);
nand UO_1314 (O_1314,N_19837,N_19686);
or UO_1315 (O_1315,N_19996,N_19729);
nand UO_1316 (O_1316,N_19894,N_19771);
or UO_1317 (O_1317,N_19932,N_19603);
nand UO_1318 (O_1318,N_19994,N_19549);
or UO_1319 (O_1319,N_19926,N_19743);
and UO_1320 (O_1320,N_19959,N_19536);
or UO_1321 (O_1321,N_19864,N_19709);
or UO_1322 (O_1322,N_19824,N_19792);
and UO_1323 (O_1323,N_19581,N_19683);
and UO_1324 (O_1324,N_19774,N_19521);
nor UO_1325 (O_1325,N_19635,N_19816);
nor UO_1326 (O_1326,N_19586,N_19708);
nor UO_1327 (O_1327,N_19580,N_19987);
or UO_1328 (O_1328,N_19575,N_19614);
and UO_1329 (O_1329,N_19900,N_19876);
and UO_1330 (O_1330,N_19975,N_19652);
or UO_1331 (O_1331,N_19822,N_19955);
nor UO_1332 (O_1332,N_19641,N_19937);
nand UO_1333 (O_1333,N_19609,N_19939);
nand UO_1334 (O_1334,N_19901,N_19872);
and UO_1335 (O_1335,N_19645,N_19642);
or UO_1336 (O_1336,N_19758,N_19966);
nor UO_1337 (O_1337,N_19920,N_19716);
and UO_1338 (O_1338,N_19507,N_19874);
and UO_1339 (O_1339,N_19792,N_19514);
or UO_1340 (O_1340,N_19541,N_19639);
or UO_1341 (O_1341,N_19502,N_19852);
or UO_1342 (O_1342,N_19598,N_19986);
and UO_1343 (O_1343,N_19614,N_19737);
and UO_1344 (O_1344,N_19590,N_19878);
nor UO_1345 (O_1345,N_19721,N_19820);
nor UO_1346 (O_1346,N_19557,N_19514);
nor UO_1347 (O_1347,N_19744,N_19646);
nand UO_1348 (O_1348,N_19613,N_19914);
and UO_1349 (O_1349,N_19616,N_19829);
nand UO_1350 (O_1350,N_19577,N_19758);
nand UO_1351 (O_1351,N_19849,N_19723);
or UO_1352 (O_1352,N_19964,N_19744);
nor UO_1353 (O_1353,N_19728,N_19918);
and UO_1354 (O_1354,N_19674,N_19732);
xnor UO_1355 (O_1355,N_19598,N_19922);
or UO_1356 (O_1356,N_19688,N_19921);
or UO_1357 (O_1357,N_19501,N_19828);
or UO_1358 (O_1358,N_19915,N_19705);
and UO_1359 (O_1359,N_19784,N_19571);
or UO_1360 (O_1360,N_19788,N_19533);
or UO_1361 (O_1361,N_19688,N_19773);
nand UO_1362 (O_1362,N_19537,N_19950);
and UO_1363 (O_1363,N_19910,N_19754);
nand UO_1364 (O_1364,N_19900,N_19826);
or UO_1365 (O_1365,N_19735,N_19988);
nor UO_1366 (O_1366,N_19865,N_19645);
and UO_1367 (O_1367,N_19505,N_19734);
or UO_1368 (O_1368,N_19972,N_19841);
and UO_1369 (O_1369,N_19842,N_19871);
and UO_1370 (O_1370,N_19934,N_19974);
nor UO_1371 (O_1371,N_19977,N_19741);
and UO_1372 (O_1372,N_19828,N_19511);
nor UO_1373 (O_1373,N_19591,N_19533);
nand UO_1374 (O_1374,N_19736,N_19563);
and UO_1375 (O_1375,N_19925,N_19709);
or UO_1376 (O_1376,N_19712,N_19719);
nand UO_1377 (O_1377,N_19780,N_19563);
nand UO_1378 (O_1378,N_19882,N_19804);
or UO_1379 (O_1379,N_19536,N_19914);
or UO_1380 (O_1380,N_19938,N_19553);
or UO_1381 (O_1381,N_19597,N_19608);
and UO_1382 (O_1382,N_19973,N_19925);
nor UO_1383 (O_1383,N_19833,N_19594);
nand UO_1384 (O_1384,N_19540,N_19501);
nand UO_1385 (O_1385,N_19954,N_19795);
and UO_1386 (O_1386,N_19816,N_19709);
and UO_1387 (O_1387,N_19622,N_19652);
or UO_1388 (O_1388,N_19713,N_19953);
or UO_1389 (O_1389,N_19940,N_19946);
nor UO_1390 (O_1390,N_19502,N_19941);
or UO_1391 (O_1391,N_19906,N_19640);
and UO_1392 (O_1392,N_19972,N_19850);
and UO_1393 (O_1393,N_19660,N_19667);
nor UO_1394 (O_1394,N_19755,N_19996);
nor UO_1395 (O_1395,N_19574,N_19828);
and UO_1396 (O_1396,N_19681,N_19892);
or UO_1397 (O_1397,N_19794,N_19630);
and UO_1398 (O_1398,N_19811,N_19968);
nand UO_1399 (O_1399,N_19648,N_19698);
nor UO_1400 (O_1400,N_19984,N_19592);
nor UO_1401 (O_1401,N_19838,N_19801);
nor UO_1402 (O_1402,N_19884,N_19833);
or UO_1403 (O_1403,N_19674,N_19665);
nor UO_1404 (O_1404,N_19776,N_19510);
nand UO_1405 (O_1405,N_19890,N_19798);
nor UO_1406 (O_1406,N_19939,N_19803);
and UO_1407 (O_1407,N_19612,N_19830);
nand UO_1408 (O_1408,N_19653,N_19686);
and UO_1409 (O_1409,N_19926,N_19704);
and UO_1410 (O_1410,N_19707,N_19851);
nand UO_1411 (O_1411,N_19889,N_19599);
nor UO_1412 (O_1412,N_19891,N_19509);
or UO_1413 (O_1413,N_19670,N_19874);
nand UO_1414 (O_1414,N_19883,N_19747);
nor UO_1415 (O_1415,N_19703,N_19734);
nor UO_1416 (O_1416,N_19760,N_19602);
nor UO_1417 (O_1417,N_19917,N_19701);
and UO_1418 (O_1418,N_19830,N_19736);
nand UO_1419 (O_1419,N_19568,N_19933);
or UO_1420 (O_1420,N_19502,N_19561);
and UO_1421 (O_1421,N_19599,N_19684);
nor UO_1422 (O_1422,N_19951,N_19988);
and UO_1423 (O_1423,N_19507,N_19799);
nor UO_1424 (O_1424,N_19559,N_19909);
nor UO_1425 (O_1425,N_19984,N_19712);
nor UO_1426 (O_1426,N_19894,N_19855);
or UO_1427 (O_1427,N_19786,N_19843);
and UO_1428 (O_1428,N_19883,N_19782);
nor UO_1429 (O_1429,N_19686,N_19596);
or UO_1430 (O_1430,N_19764,N_19779);
nor UO_1431 (O_1431,N_19774,N_19916);
and UO_1432 (O_1432,N_19793,N_19967);
and UO_1433 (O_1433,N_19913,N_19956);
and UO_1434 (O_1434,N_19863,N_19741);
and UO_1435 (O_1435,N_19524,N_19517);
nand UO_1436 (O_1436,N_19636,N_19917);
or UO_1437 (O_1437,N_19643,N_19570);
or UO_1438 (O_1438,N_19984,N_19919);
nor UO_1439 (O_1439,N_19916,N_19501);
or UO_1440 (O_1440,N_19619,N_19512);
nand UO_1441 (O_1441,N_19799,N_19572);
and UO_1442 (O_1442,N_19819,N_19936);
and UO_1443 (O_1443,N_19685,N_19762);
or UO_1444 (O_1444,N_19884,N_19721);
nand UO_1445 (O_1445,N_19717,N_19650);
and UO_1446 (O_1446,N_19780,N_19905);
nor UO_1447 (O_1447,N_19504,N_19723);
or UO_1448 (O_1448,N_19652,N_19936);
nor UO_1449 (O_1449,N_19861,N_19828);
xnor UO_1450 (O_1450,N_19745,N_19972);
nor UO_1451 (O_1451,N_19554,N_19643);
nor UO_1452 (O_1452,N_19904,N_19897);
nor UO_1453 (O_1453,N_19560,N_19908);
or UO_1454 (O_1454,N_19501,N_19718);
nand UO_1455 (O_1455,N_19722,N_19972);
or UO_1456 (O_1456,N_19560,N_19589);
nand UO_1457 (O_1457,N_19975,N_19912);
nor UO_1458 (O_1458,N_19833,N_19526);
or UO_1459 (O_1459,N_19642,N_19963);
or UO_1460 (O_1460,N_19985,N_19939);
or UO_1461 (O_1461,N_19585,N_19782);
or UO_1462 (O_1462,N_19562,N_19583);
and UO_1463 (O_1463,N_19637,N_19538);
nor UO_1464 (O_1464,N_19617,N_19507);
nand UO_1465 (O_1465,N_19950,N_19817);
nand UO_1466 (O_1466,N_19620,N_19669);
nor UO_1467 (O_1467,N_19549,N_19936);
or UO_1468 (O_1468,N_19994,N_19649);
nand UO_1469 (O_1469,N_19625,N_19555);
nand UO_1470 (O_1470,N_19738,N_19931);
nor UO_1471 (O_1471,N_19695,N_19543);
nor UO_1472 (O_1472,N_19919,N_19983);
nand UO_1473 (O_1473,N_19829,N_19787);
nand UO_1474 (O_1474,N_19994,N_19656);
and UO_1475 (O_1475,N_19668,N_19995);
nand UO_1476 (O_1476,N_19889,N_19973);
and UO_1477 (O_1477,N_19612,N_19773);
nor UO_1478 (O_1478,N_19883,N_19725);
nand UO_1479 (O_1479,N_19639,N_19748);
nor UO_1480 (O_1480,N_19503,N_19993);
and UO_1481 (O_1481,N_19804,N_19737);
nor UO_1482 (O_1482,N_19780,N_19815);
and UO_1483 (O_1483,N_19651,N_19772);
or UO_1484 (O_1484,N_19610,N_19591);
nand UO_1485 (O_1485,N_19588,N_19870);
and UO_1486 (O_1486,N_19803,N_19670);
or UO_1487 (O_1487,N_19559,N_19845);
and UO_1488 (O_1488,N_19726,N_19587);
nand UO_1489 (O_1489,N_19888,N_19690);
or UO_1490 (O_1490,N_19796,N_19773);
nor UO_1491 (O_1491,N_19868,N_19589);
and UO_1492 (O_1492,N_19955,N_19573);
and UO_1493 (O_1493,N_19971,N_19813);
nand UO_1494 (O_1494,N_19942,N_19986);
nor UO_1495 (O_1495,N_19730,N_19701);
and UO_1496 (O_1496,N_19634,N_19616);
nor UO_1497 (O_1497,N_19859,N_19993);
nand UO_1498 (O_1498,N_19749,N_19734);
nand UO_1499 (O_1499,N_19596,N_19827);
nor UO_1500 (O_1500,N_19766,N_19967);
or UO_1501 (O_1501,N_19855,N_19554);
nor UO_1502 (O_1502,N_19508,N_19715);
and UO_1503 (O_1503,N_19787,N_19957);
and UO_1504 (O_1504,N_19898,N_19559);
nor UO_1505 (O_1505,N_19731,N_19937);
or UO_1506 (O_1506,N_19844,N_19510);
or UO_1507 (O_1507,N_19849,N_19779);
and UO_1508 (O_1508,N_19565,N_19758);
nand UO_1509 (O_1509,N_19935,N_19744);
or UO_1510 (O_1510,N_19570,N_19569);
or UO_1511 (O_1511,N_19675,N_19842);
xor UO_1512 (O_1512,N_19886,N_19915);
nor UO_1513 (O_1513,N_19853,N_19687);
or UO_1514 (O_1514,N_19955,N_19745);
or UO_1515 (O_1515,N_19687,N_19772);
or UO_1516 (O_1516,N_19818,N_19559);
or UO_1517 (O_1517,N_19873,N_19716);
and UO_1518 (O_1518,N_19593,N_19975);
nor UO_1519 (O_1519,N_19624,N_19505);
nor UO_1520 (O_1520,N_19574,N_19698);
nand UO_1521 (O_1521,N_19694,N_19529);
nand UO_1522 (O_1522,N_19677,N_19551);
and UO_1523 (O_1523,N_19743,N_19826);
and UO_1524 (O_1524,N_19636,N_19995);
or UO_1525 (O_1525,N_19851,N_19668);
and UO_1526 (O_1526,N_19686,N_19865);
nand UO_1527 (O_1527,N_19939,N_19790);
nor UO_1528 (O_1528,N_19854,N_19725);
xnor UO_1529 (O_1529,N_19679,N_19798);
nor UO_1530 (O_1530,N_19785,N_19794);
nand UO_1531 (O_1531,N_19675,N_19860);
and UO_1532 (O_1532,N_19908,N_19790);
nor UO_1533 (O_1533,N_19630,N_19982);
nand UO_1534 (O_1534,N_19556,N_19711);
nor UO_1535 (O_1535,N_19635,N_19987);
and UO_1536 (O_1536,N_19828,N_19983);
nor UO_1537 (O_1537,N_19627,N_19872);
or UO_1538 (O_1538,N_19621,N_19572);
nor UO_1539 (O_1539,N_19611,N_19506);
or UO_1540 (O_1540,N_19810,N_19716);
and UO_1541 (O_1541,N_19726,N_19650);
or UO_1542 (O_1542,N_19650,N_19926);
nor UO_1543 (O_1543,N_19695,N_19654);
nor UO_1544 (O_1544,N_19888,N_19622);
or UO_1545 (O_1545,N_19926,N_19757);
and UO_1546 (O_1546,N_19853,N_19771);
or UO_1547 (O_1547,N_19623,N_19572);
nand UO_1548 (O_1548,N_19503,N_19566);
and UO_1549 (O_1549,N_19850,N_19679);
and UO_1550 (O_1550,N_19556,N_19512);
nor UO_1551 (O_1551,N_19724,N_19591);
or UO_1552 (O_1552,N_19609,N_19944);
and UO_1553 (O_1553,N_19661,N_19707);
nor UO_1554 (O_1554,N_19854,N_19791);
nor UO_1555 (O_1555,N_19604,N_19805);
and UO_1556 (O_1556,N_19572,N_19592);
and UO_1557 (O_1557,N_19823,N_19839);
or UO_1558 (O_1558,N_19729,N_19784);
nor UO_1559 (O_1559,N_19979,N_19916);
and UO_1560 (O_1560,N_19945,N_19724);
and UO_1561 (O_1561,N_19603,N_19524);
nand UO_1562 (O_1562,N_19619,N_19502);
nor UO_1563 (O_1563,N_19540,N_19996);
nand UO_1564 (O_1564,N_19831,N_19682);
and UO_1565 (O_1565,N_19527,N_19799);
nand UO_1566 (O_1566,N_19905,N_19633);
nand UO_1567 (O_1567,N_19557,N_19641);
and UO_1568 (O_1568,N_19787,N_19539);
or UO_1569 (O_1569,N_19635,N_19532);
or UO_1570 (O_1570,N_19566,N_19865);
and UO_1571 (O_1571,N_19697,N_19763);
or UO_1572 (O_1572,N_19982,N_19984);
and UO_1573 (O_1573,N_19766,N_19801);
nor UO_1574 (O_1574,N_19978,N_19980);
or UO_1575 (O_1575,N_19720,N_19729);
nor UO_1576 (O_1576,N_19763,N_19821);
nand UO_1577 (O_1577,N_19899,N_19781);
or UO_1578 (O_1578,N_19920,N_19887);
nor UO_1579 (O_1579,N_19905,N_19669);
or UO_1580 (O_1580,N_19831,N_19760);
nor UO_1581 (O_1581,N_19532,N_19758);
nor UO_1582 (O_1582,N_19913,N_19934);
nor UO_1583 (O_1583,N_19613,N_19578);
nor UO_1584 (O_1584,N_19816,N_19639);
and UO_1585 (O_1585,N_19725,N_19855);
nand UO_1586 (O_1586,N_19848,N_19542);
or UO_1587 (O_1587,N_19953,N_19579);
nand UO_1588 (O_1588,N_19956,N_19664);
nor UO_1589 (O_1589,N_19605,N_19675);
nand UO_1590 (O_1590,N_19826,N_19623);
nor UO_1591 (O_1591,N_19663,N_19531);
nand UO_1592 (O_1592,N_19924,N_19635);
nor UO_1593 (O_1593,N_19594,N_19861);
and UO_1594 (O_1594,N_19792,N_19788);
nand UO_1595 (O_1595,N_19729,N_19761);
or UO_1596 (O_1596,N_19645,N_19854);
and UO_1597 (O_1597,N_19597,N_19928);
and UO_1598 (O_1598,N_19866,N_19783);
nand UO_1599 (O_1599,N_19971,N_19854);
and UO_1600 (O_1600,N_19826,N_19864);
nand UO_1601 (O_1601,N_19648,N_19536);
or UO_1602 (O_1602,N_19735,N_19644);
and UO_1603 (O_1603,N_19916,N_19726);
and UO_1604 (O_1604,N_19641,N_19771);
and UO_1605 (O_1605,N_19966,N_19719);
or UO_1606 (O_1606,N_19948,N_19539);
nor UO_1607 (O_1607,N_19668,N_19704);
or UO_1608 (O_1608,N_19777,N_19690);
or UO_1609 (O_1609,N_19743,N_19930);
or UO_1610 (O_1610,N_19593,N_19541);
xnor UO_1611 (O_1611,N_19716,N_19861);
xnor UO_1612 (O_1612,N_19819,N_19500);
xor UO_1613 (O_1613,N_19817,N_19549);
and UO_1614 (O_1614,N_19548,N_19855);
nor UO_1615 (O_1615,N_19519,N_19923);
and UO_1616 (O_1616,N_19877,N_19941);
nand UO_1617 (O_1617,N_19508,N_19987);
nor UO_1618 (O_1618,N_19970,N_19541);
and UO_1619 (O_1619,N_19735,N_19537);
nand UO_1620 (O_1620,N_19953,N_19777);
and UO_1621 (O_1621,N_19765,N_19913);
and UO_1622 (O_1622,N_19859,N_19533);
nand UO_1623 (O_1623,N_19978,N_19623);
and UO_1624 (O_1624,N_19719,N_19673);
and UO_1625 (O_1625,N_19639,N_19728);
and UO_1626 (O_1626,N_19557,N_19815);
nor UO_1627 (O_1627,N_19878,N_19644);
nand UO_1628 (O_1628,N_19927,N_19670);
or UO_1629 (O_1629,N_19579,N_19848);
or UO_1630 (O_1630,N_19608,N_19986);
and UO_1631 (O_1631,N_19633,N_19921);
and UO_1632 (O_1632,N_19652,N_19709);
nand UO_1633 (O_1633,N_19609,N_19882);
or UO_1634 (O_1634,N_19790,N_19995);
nand UO_1635 (O_1635,N_19900,N_19514);
nor UO_1636 (O_1636,N_19974,N_19672);
and UO_1637 (O_1637,N_19766,N_19920);
nor UO_1638 (O_1638,N_19672,N_19766);
and UO_1639 (O_1639,N_19842,N_19739);
and UO_1640 (O_1640,N_19752,N_19916);
and UO_1641 (O_1641,N_19701,N_19583);
or UO_1642 (O_1642,N_19963,N_19672);
or UO_1643 (O_1643,N_19752,N_19664);
or UO_1644 (O_1644,N_19933,N_19993);
nand UO_1645 (O_1645,N_19535,N_19890);
or UO_1646 (O_1646,N_19990,N_19792);
or UO_1647 (O_1647,N_19986,N_19585);
nor UO_1648 (O_1648,N_19745,N_19661);
or UO_1649 (O_1649,N_19659,N_19897);
or UO_1650 (O_1650,N_19580,N_19961);
nor UO_1651 (O_1651,N_19643,N_19620);
nand UO_1652 (O_1652,N_19521,N_19689);
or UO_1653 (O_1653,N_19629,N_19662);
and UO_1654 (O_1654,N_19804,N_19699);
nor UO_1655 (O_1655,N_19526,N_19654);
nor UO_1656 (O_1656,N_19933,N_19909);
or UO_1657 (O_1657,N_19893,N_19970);
and UO_1658 (O_1658,N_19750,N_19566);
or UO_1659 (O_1659,N_19872,N_19819);
or UO_1660 (O_1660,N_19923,N_19936);
nor UO_1661 (O_1661,N_19509,N_19568);
nor UO_1662 (O_1662,N_19661,N_19649);
nor UO_1663 (O_1663,N_19533,N_19857);
xor UO_1664 (O_1664,N_19842,N_19911);
nand UO_1665 (O_1665,N_19624,N_19546);
nor UO_1666 (O_1666,N_19975,N_19561);
nand UO_1667 (O_1667,N_19991,N_19927);
and UO_1668 (O_1668,N_19507,N_19875);
and UO_1669 (O_1669,N_19721,N_19632);
nand UO_1670 (O_1670,N_19606,N_19747);
and UO_1671 (O_1671,N_19962,N_19749);
nor UO_1672 (O_1672,N_19859,N_19883);
nand UO_1673 (O_1673,N_19800,N_19628);
and UO_1674 (O_1674,N_19849,N_19696);
nor UO_1675 (O_1675,N_19553,N_19713);
and UO_1676 (O_1676,N_19681,N_19986);
nor UO_1677 (O_1677,N_19829,N_19763);
nor UO_1678 (O_1678,N_19595,N_19829);
nand UO_1679 (O_1679,N_19771,N_19570);
or UO_1680 (O_1680,N_19819,N_19952);
xnor UO_1681 (O_1681,N_19578,N_19576);
or UO_1682 (O_1682,N_19802,N_19545);
and UO_1683 (O_1683,N_19701,N_19710);
and UO_1684 (O_1684,N_19842,N_19929);
nand UO_1685 (O_1685,N_19842,N_19775);
and UO_1686 (O_1686,N_19882,N_19976);
nor UO_1687 (O_1687,N_19954,N_19737);
and UO_1688 (O_1688,N_19890,N_19939);
or UO_1689 (O_1689,N_19813,N_19703);
or UO_1690 (O_1690,N_19828,N_19723);
or UO_1691 (O_1691,N_19976,N_19526);
nor UO_1692 (O_1692,N_19563,N_19781);
nor UO_1693 (O_1693,N_19909,N_19745);
nor UO_1694 (O_1694,N_19718,N_19875);
nor UO_1695 (O_1695,N_19607,N_19758);
nand UO_1696 (O_1696,N_19636,N_19909);
or UO_1697 (O_1697,N_19769,N_19635);
and UO_1698 (O_1698,N_19616,N_19879);
and UO_1699 (O_1699,N_19720,N_19698);
nand UO_1700 (O_1700,N_19524,N_19673);
nand UO_1701 (O_1701,N_19742,N_19734);
nand UO_1702 (O_1702,N_19592,N_19622);
or UO_1703 (O_1703,N_19933,N_19805);
nand UO_1704 (O_1704,N_19642,N_19610);
nand UO_1705 (O_1705,N_19958,N_19914);
nand UO_1706 (O_1706,N_19701,N_19620);
nand UO_1707 (O_1707,N_19786,N_19681);
and UO_1708 (O_1708,N_19731,N_19522);
or UO_1709 (O_1709,N_19768,N_19905);
nor UO_1710 (O_1710,N_19524,N_19994);
nor UO_1711 (O_1711,N_19619,N_19988);
xnor UO_1712 (O_1712,N_19826,N_19993);
and UO_1713 (O_1713,N_19640,N_19644);
nor UO_1714 (O_1714,N_19658,N_19989);
nand UO_1715 (O_1715,N_19642,N_19749);
and UO_1716 (O_1716,N_19918,N_19862);
nand UO_1717 (O_1717,N_19843,N_19834);
nor UO_1718 (O_1718,N_19903,N_19905);
or UO_1719 (O_1719,N_19539,N_19605);
and UO_1720 (O_1720,N_19797,N_19933);
and UO_1721 (O_1721,N_19585,N_19727);
nor UO_1722 (O_1722,N_19785,N_19596);
xor UO_1723 (O_1723,N_19610,N_19828);
nand UO_1724 (O_1724,N_19896,N_19790);
or UO_1725 (O_1725,N_19954,N_19680);
nor UO_1726 (O_1726,N_19774,N_19784);
and UO_1727 (O_1727,N_19693,N_19761);
or UO_1728 (O_1728,N_19674,N_19963);
nand UO_1729 (O_1729,N_19575,N_19689);
and UO_1730 (O_1730,N_19663,N_19737);
nor UO_1731 (O_1731,N_19988,N_19736);
nor UO_1732 (O_1732,N_19507,N_19637);
nor UO_1733 (O_1733,N_19912,N_19562);
nand UO_1734 (O_1734,N_19869,N_19530);
and UO_1735 (O_1735,N_19713,N_19748);
and UO_1736 (O_1736,N_19995,N_19899);
nor UO_1737 (O_1737,N_19893,N_19901);
and UO_1738 (O_1738,N_19640,N_19627);
or UO_1739 (O_1739,N_19912,N_19626);
nor UO_1740 (O_1740,N_19504,N_19716);
or UO_1741 (O_1741,N_19514,N_19591);
nand UO_1742 (O_1742,N_19550,N_19806);
nor UO_1743 (O_1743,N_19592,N_19992);
and UO_1744 (O_1744,N_19889,N_19906);
nor UO_1745 (O_1745,N_19556,N_19693);
and UO_1746 (O_1746,N_19695,N_19530);
and UO_1747 (O_1747,N_19572,N_19707);
nand UO_1748 (O_1748,N_19547,N_19669);
nand UO_1749 (O_1749,N_19726,N_19803);
nand UO_1750 (O_1750,N_19624,N_19520);
and UO_1751 (O_1751,N_19500,N_19831);
and UO_1752 (O_1752,N_19779,N_19515);
and UO_1753 (O_1753,N_19612,N_19994);
or UO_1754 (O_1754,N_19768,N_19815);
nand UO_1755 (O_1755,N_19921,N_19738);
or UO_1756 (O_1756,N_19607,N_19852);
and UO_1757 (O_1757,N_19713,N_19575);
and UO_1758 (O_1758,N_19930,N_19831);
nor UO_1759 (O_1759,N_19736,N_19731);
and UO_1760 (O_1760,N_19956,N_19999);
nor UO_1761 (O_1761,N_19528,N_19774);
or UO_1762 (O_1762,N_19604,N_19568);
or UO_1763 (O_1763,N_19802,N_19646);
nand UO_1764 (O_1764,N_19823,N_19925);
nand UO_1765 (O_1765,N_19975,N_19964);
or UO_1766 (O_1766,N_19527,N_19725);
nand UO_1767 (O_1767,N_19732,N_19965);
and UO_1768 (O_1768,N_19657,N_19888);
nor UO_1769 (O_1769,N_19971,N_19538);
nor UO_1770 (O_1770,N_19971,N_19633);
or UO_1771 (O_1771,N_19507,N_19555);
nand UO_1772 (O_1772,N_19591,N_19605);
or UO_1773 (O_1773,N_19572,N_19546);
and UO_1774 (O_1774,N_19724,N_19771);
and UO_1775 (O_1775,N_19874,N_19953);
nand UO_1776 (O_1776,N_19550,N_19741);
nand UO_1777 (O_1777,N_19617,N_19868);
and UO_1778 (O_1778,N_19573,N_19746);
nand UO_1779 (O_1779,N_19536,N_19842);
nand UO_1780 (O_1780,N_19907,N_19583);
nor UO_1781 (O_1781,N_19572,N_19910);
nand UO_1782 (O_1782,N_19818,N_19602);
nor UO_1783 (O_1783,N_19551,N_19634);
and UO_1784 (O_1784,N_19543,N_19876);
and UO_1785 (O_1785,N_19620,N_19563);
and UO_1786 (O_1786,N_19714,N_19676);
or UO_1787 (O_1787,N_19702,N_19776);
or UO_1788 (O_1788,N_19718,N_19555);
nand UO_1789 (O_1789,N_19811,N_19760);
and UO_1790 (O_1790,N_19552,N_19800);
nand UO_1791 (O_1791,N_19668,N_19864);
or UO_1792 (O_1792,N_19934,N_19876);
nor UO_1793 (O_1793,N_19563,N_19921);
and UO_1794 (O_1794,N_19848,N_19847);
nor UO_1795 (O_1795,N_19931,N_19880);
nand UO_1796 (O_1796,N_19514,N_19655);
and UO_1797 (O_1797,N_19671,N_19636);
nand UO_1798 (O_1798,N_19838,N_19870);
or UO_1799 (O_1799,N_19858,N_19906);
nor UO_1800 (O_1800,N_19550,N_19564);
nand UO_1801 (O_1801,N_19750,N_19829);
or UO_1802 (O_1802,N_19781,N_19653);
nand UO_1803 (O_1803,N_19709,N_19746);
nand UO_1804 (O_1804,N_19721,N_19758);
or UO_1805 (O_1805,N_19710,N_19879);
nand UO_1806 (O_1806,N_19846,N_19662);
nand UO_1807 (O_1807,N_19802,N_19744);
and UO_1808 (O_1808,N_19964,N_19732);
or UO_1809 (O_1809,N_19909,N_19538);
and UO_1810 (O_1810,N_19513,N_19968);
nand UO_1811 (O_1811,N_19858,N_19886);
nand UO_1812 (O_1812,N_19733,N_19935);
nor UO_1813 (O_1813,N_19538,N_19740);
xnor UO_1814 (O_1814,N_19802,N_19642);
or UO_1815 (O_1815,N_19706,N_19700);
nand UO_1816 (O_1816,N_19719,N_19650);
and UO_1817 (O_1817,N_19947,N_19829);
or UO_1818 (O_1818,N_19527,N_19803);
nand UO_1819 (O_1819,N_19775,N_19530);
and UO_1820 (O_1820,N_19535,N_19528);
nand UO_1821 (O_1821,N_19518,N_19554);
or UO_1822 (O_1822,N_19818,N_19713);
nor UO_1823 (O_1823,N_19996,N_19913);
nor UO_1824 (O_1824,N_19756,N_19623);
nand UO_1825 (O_1825,N_19751,N_19593);
nand UO_1826 (O_1826,N_19768,N_19670);
nand UO_1827 (O_1827,N_19883,N_19962);
and UO_1828 (O_1828,N_19802,N_19757);
and UO_1829 (O_1829,N_19639,N_19646);
nor UO_1830 (O_1830,N_19775,N_19731);
nand UO_1831 (O_1831,N_19695,N_19909);
or UO_1832 (O_1832,N_19980,N_19959);
nor UO_1833 (O_1833,N_19613,N_19520);
or UO_1834 (O_1834,N_19812,N_19671);
nand UO_1835 (O_1835,N_19827,N_19808);
or UO_1836 (O_1836,N_19657,N_19512);
or UO_1837 (O_1837,N_19955,N_19821);
xor UO_1838 (O_1838,N_19890,N_19536);
and UO_1839 (O_1839,N_19553,N_19506);
nor UO_1840 (O_1840,N_19580,N_19829);
and UO_1841 (O_1841,N_19669,N_19568);
nor UO_1842 (O_1842,N_19545,N_19513);
or UO_1843 (O_1843,N_19955,N_19594);
nor UO_1844 (O_1844,N_19937,N_19509);
or UO_1845 (O_1845,N_19961,N_19523);
nor UO_1846 (O_1846,N_19881,N_19909);
nor UO_1847 (O_1847,N_19613,N_19564);
nor UO_1848 (O_1848,N_19860,N_19593);
or UO_1849 (O_1849,N_19809,N_19901);
nand UO_1850 (O_1850,N_19793,N_19974);
nor UO_1851 (O_1851,N_19762,N_19554);
and UO_1852 (O_1852,N_19806,N_19913);
xor UO_1853 (O_1853,N_19782,N_19508);
or UO_1854 (O_1854,N_19694,N_19951);
nand UO_1855 (O_1855,N_19700,N_19630);
and UO_1856 (O_1856,N_19566,N_19629);
nor UO_1857 (O_1857,N_19779,N_19930);
nand UO_1858 (O_1858,N_19684,N_19803);
and UO_1859 (O_1859,N_19504,N_19581);
nor UO_1860 (O_1860,N_19660,N_19676);
and UO_1861 (O_1861,N_19907,N_19506);
nor UO_1862 (O_1862,N_19930,N_19561);
nor UO_1863 (O_1863,N_19649,N_19796);
xor UO_1864 (O_1864,N_19750,N_19736);
nor UO_1865 (O_1865,N_19753,N_19686);
nand UO_1866 (O_1866,N_19779,N_19875);
and UO_1867 (O_1867,N_19565,N_19740);
and UO_1868 (O_1868,N_19830,N_19557);
and UO_1869 (O_1869,N_19654,N_19858);
nand UO_1870 (O_1870,N_19613,N_19618);
nor UO_1871 (O_1871,N_19576,N_19981);
or UO_1872 (O_1872,N_19519,N_19842);
and UO_1873 (O_1873,N_19680,N_19525);
and UO_1874 (O_1874,N_19677,N_19571);
and UO_1875 (O_1875,N_19646,N_19959);
and UO_1876 (O_1876,N_19758,N_19608);
and UO_1877 (O_1877,N_19508,N_19697);
or UO_1878 (O_1878,N_19878,N_19997);
and UO_1879 (O_1879,N_19664,N_19586);
and UO_1880 (O_1880,N_19806,N_19888);
nand UO_1881 (O_1881,N_19840,N_19507);
and UO_1882 (O_1882,N_19995,N_19938);
or UO_1883 (O_1883,N_19577,N_19528);
nor UO_1884 (O_1884,N_19769,N_19892);
or UO_1885 (O_1885,N_19754,N_19545);
and UO_1886 (O_1886,N_19849,N_19989);
or UO_1887 (O_1887,N_19571,N_19981);
or UO_1888 (O_1888,N_19691,N_19692);
nand UO_1889 (O_1889,N_19820,N_19897);
nand UO_1890 (O_1890,N_19831,N_19704);
or UO_1891 (O_1891,N_19916,N_19971);
nor UO_1892 (O_1892,N_19755,N_19923);
nand UO_1893 (O_1893,N_19531,N_19653);
nand UO_1894 (O_1894,N_19772,N_19964);
and UO_1895 (O_1895,N_19688,N_19967);
nand UO_1896 (O_1896,N_19838,N_19844);
and UO_1897 (O_1897,N_19958,N_19788);
nor UO_1898 (O_1898,N_19920,N_19722);
nand UO_1899 (O_1899,N_19940,N_19666);
nor UO_1900 (O_1900,N_19747,N_19731);
nand UO_1901 (O_1901,N_19729,N_19603);
or UO_1902 (O_1902,N_19755,N_19709);
nand UO_1903 (O_1903,N_19579,N_19897);
or UO_1904 (O_1904,N_19618,N_19921);
or UO_1905 (O_1905,N_19604,N_19821);
nor UO_1906 (O_1906,N_19547,N_19922);
nor UO_1907 (O_1907,N_19895,N_19600);
nor UO_1908 (O_1908,N_19701,N_19742);
and UO_1909 (O_1909,N_19825,N_19690);
nor UO_1910 (O_1910,N_19545,N_19964);
or UO_1911 (O_1911,N_19835,N_19587);
nand UO_1912 (O_1912,N_19782,N_19677);
nand UO_1913 (O_1913,N_19650,N_19834);
nor UO_1914 (O_1914,N_19883,N_19716);
and UO_1915 (O_1915,N_19648,N_19575);
nor UO_1916 (O_1916,N_19926,N_19584);
or UO_1917 (O_1917,N_19662,N_19691);
nand UO_1918 (O_1918,N_19675,N_19577);
nor UO_1919 (O_1919,N_19711,N_19515);
or UO_1920 (O_1920,N_19572,N_19747);
xnor UO_1921 (O_1921,N_19971,N_19563);
and UO_1922 (O_1922,N_19596,N_19604);
nor UO_1923 (O_1923,N_19853,N_19671);
and UO_1924 (O_1924,N_19563,N_19891);
nand UO_1925 (O_1925,N_19870,N_19747);
nor UO_1926 (O_1926,N_19826,N_19843);
and UO_1927 (O_1927,N_19921,N_19901);
nor UO_1928 (O_1928,N_19501,N_19713);
nor UO_1929 (O_1929,N_19742,N_19984);
or UO_1930 (O_1930,N_19834,N_19876);
nor UO_1931 (O_1931,N_19512,N_19884);
nand UO_1932 (O_1932,N_19918,N_19816);
nor UO_1933 (O_1933,N_19508,N_19705);
nand UO_1934 (O_1934,N_19711,N_19682);
or UO_1935 (O_1935,N_19720,N_19962);
nand UO_1936 (O_1936,N_19702,N_19571);
nor UO_1937 (O_1937,N_19633,N_19770);
nand UO_1938 (O_1938,N_19984,N_19650);
and UO_1939 (O_1939,N_19763,N_19760);
or UO_1940 (O_1940,N_19546,N_19700);
nand UO_1941 (O_1941,N_19874,N_19565);
nand UO_1942 (O_1942,N_19965,N_19976);
and UO_1943 (O_1943,N_19918,N_19588);
nor UO_1944 (O_1944,N_19852,N_19636);
and UO_1945 (O_1945,N_19779,N_19938);
and UO_1946 (O_1946,N_19672,N_19675);
and UO_1947 (O_1947,N_19663,N_19834);
or UO_1948 (O_1948,N_19923,N_19580);
nand UO_1949 (O_1949,N_19600,N_19941);
and UO_1950 (O_1950,N_19551,N_19597);
and UO_1951 (O_1951,N_19580,N_19784);
and UO_1952 (O_1952,N_19741,N_19636);
xnor UO_1953 (O_1953,N_19703,N_19655);
nand UO_1954 (O_1954,N_19713,N_19793);
nor UO_1955 (O_1955,N_19853,N_19586);
and UO_1956 (O_1956,N_19912,N_19748);
and UO_1957 (O_1957,N_19710,N_19640);
and UO_1958 (O_1958,N_19871,N_19747);
nor UO_1959 (O_1959,N_19612,N_19952);
nand UO_1960 (O_1960,N_19768,N_19841);
or UO_1961 (O_1961,N_19561,N_19823);
or UO_1962 (O_1962,N_19794,N_19973);
nor UO_1963 (O_1963,N_19795,N_19663);
and UO_1964 (O_1964,N_19829,N_19828);
or UO_1965 (O_1965,N_19649,N_19846);
or UO_1966 (O_1966,N_19740,N_19929);
and UO_1967 (O_1967,N_19500,N_19604);
and UO_1968 (O_1968,N_19684,N_19519);
nor UO_1969 (O_1969,N_19511,N_19717);
or UO_1970 (O_1970,N_19651,N_19521);
nand UO_1971 (O_1971,N_19814,N_19992);
nand UO_1972 (O_1972,N_19800,N_19807);
or UO_1973 (O_1973,N_19770,N_19747);
nand UO_1974 (O_1974,N_19758,N_19704);
nand UO_1975 (O_1975,N_19683,N_19550);
nor UO_1976 (O_1976,N_19650,N_19676);
or UO_1977 (O_1977,N_19551,N_19807);
or UO_1978 (O_1978,N_19687,N_19840);
nor UO_1979 (O_1979,N_19566,N_19506);
and UO_1980 (O_1980,N_19888,N_19818);
or UO_1981 (O_1981,N_19928,N_19553);
nand UO_1982 (O_1982,N_19724,N_19720);
nand UO_1983 (O_1983,N_19910,N_19899);
nand UO_1984 (O_1984,N_19761,N_19918);
nor UO_1985 (O_1985,N_19970,N_19581);
nor UO_1986 (O_1986,N_19624,N_19814);
nor UO_1987 (O_1987,N_19513,N_19565);
nand UO_1988 (O_1988,N_19643,N_19813);
and UO_1989 (O_1989,N_19537,N_19782);
nor UO_1990 (O_1990,N_19782,N_19887);
nand UO_1991 (O_1991,N_19904,N_19505);
nand UO_1992 (O_1992,N_19841,N_19622);
or UO_1993 (O_1993,N_19675,N_19829);
and UO_1994 (O_1994,N_19596,N_19602);
or UO_1995 (O_1995,N_19971,N_19603);
nand UO_1996 (O_1996,N_19597,N_19942);
or UO_1997 (O_1997,N_19917,N_19515);
nand UO_1998 (O_1998,N_19704,N_19787);
nand UO_1999 (O_1999,N_19967,N_19537);
and UO_2000 (O_2000,N_19887,N_19729);
and UO_2001 (O_2001,N_19737,N_19574);
nand UO_2002 (O_2002,N_19520,N_19799);
and UO_2003 (O_2003,N_19691,N_19796);
nand UO_2004 (O_2004,N_19569,N_19927);
nand UO_2005 (O_2005,N_19831,N_19895);
nor UO_2006 (O_2006,N_19926,N_19867);
and UO_2007 (O_2007,N_19869,N_19691);
or UO_2008 (O_2008,N_19910,N_19612);
nand UO_2009 (O_2009,N_19592,N_19763);
nand UO_2010 (O_2010,N_19888,N_19979);
nor UO_2011 (O_2011,N_19603,N_19595);
and UO_2012 (O_2012,N_19661,N_19654);
and UO_2013 (O_2013,N_19609,N_19689);
nor UO_2014 (O_2014,N_19784,N_19870);
nor UO_2015 (O_2015,N_19788,N_19815);
or UO_2016 (O_2016,N_19853,N_19698);
or UO_2017 (O_2017,N_19843,N_19893);
nor UO_2018 (O_2018,N_19969,N_19551);
nor UO_2019 (O_2019,N_19757,N_19570);
nand UO_2020 (O_2020,N_19780,N_19889);
nand UO_2021 (O_2021,N_19994,N_19709);
or UO_2022 (O_2022,N_19857,N_19818);
or UO_2023 (O_2023,N_19586,N_19595);
and UO_2024 (O_2024,N_19753,N_19603);
nor UO_2025 (O_2025,N_19630,N_19695);
nor UO_2026 (O_2026,N_19975,N_19646);
nand UO_2027 (O_2027,N_19953,N_19686);
nor UO_2028 (O_2028,N_19665,N_19843);
xnor UO_2029 (O_2029,N_19516,N_19793);
nand UO_2030 (O_2030,N_19555,N_19674);
and UO_2031 (O_2031,N_19954,N_19700);
nor UO_2032 (O_2032,N_19944,N_19641);
nor UO_2033 (O_2033,N_19923,N_19595);
and UO_2034 (O_2034,N_19972,N_19673);
or UO_2035 (O_2035,N_19653,N_19752);
and UO_2036 (O_2036,N_19850,N_19673);
or UO_2037 (O_2037,N_19866,N_19804);
or UO_2038 (O_2038,N_19852,N_19844);
nand UO_2039 (O_2039,N_19645,N_19729);
or UO_2040 (O_2040,N_19573,N_19558);
nor UO_2041 (O_2041,N_19922,N_19673);
or UO_2042 (O_2042,N_19570,N_19796);
nor UO_2043 (O_2043,N_19620,N_19852);
nor UO_2044 (O_2044,N_19525,N_19918);
nor UO_2045 (O_2045,N_19505,N_19764);
and UO_2046 (O_2046,N_19885,N_19706);
nor UO_2047 (O_2047,N_19651,N_19980);
and UO_2048 (O_2048,N_19721,N_19789);
nand UO_2049 (O_2049,N_19930,N_19623);
or UO_2050 (O_2050,N_19758,N_19720);
nor UO_2051 (O_2051,N_19596,N_19500);
nor UO_2052 (O_2052,N_19981,N_19831);
nand UO_2053 (O_2053,N_19882,N_19974);
or UO_2054 (O_2054,N_19568,N_19797);
or UO_2055 (O_2055,N_19733,N_19849);
or UO_2056 (O_2056,N_19587,N_19624);
nand UO_2057 (O_2057,N_19731,N_19620);
or UO_2058 (O_2058,N_19722,N_19833);
and UO_2059 (O_2059,N_19928,N_19650);
nand UO_2060 (O_2060,N_19512,N_19883);
and UO_2061 (O_2061,N_19831,N_19993);
or UO_2062 (O_2062,N_19856,N_19701);
nand UO_2063 (O_2063,N_19674,N_19747);
nand UO_2064 (O_2064,N_19864,N_19782);
or UO_2065 (O_2065,N_19765,N_19806);
nand UO_2066 (O_2066,N_19978,N_19608);
nor UO_2067 (O_2067,N_19791,N_19572);
and UO_2068 (O_2068,N_19825,N_19959);
or UO_2069 (O_2069,N_19682,N_19597);
nor UO_2070 (O_2070,N_19834,N_19904);
or UO_2071 (O_2071,N_19994,N_19580);
nor UO_2072 (O_2072,N_19990,N_19727);
nor UO_2073 (O_2073,N_19618,N_19929);
or UO_2074 (O_2074,N_19550,N_19837);
nor UO_2075 (O_2075,N_19944,N_19751);
nor UO_2076 (O_2076,N_19661,N_19533);
nand UO_2077 (O_2077,N_19510,N_19537);
nand UO_2078 (O_2078,N_19686,N_19631);
or UO_2079 (O_2079,N_19903,N_19735);
and UO_2080 (O_2080,N_19823,N_19989);
nor UO_2081 (O_2081,N_19870,N_19692);
nor UO_2082 (O_2082,N_19961,N_19970);
nand UO_2083 (O_2083,N_19959,N_19793);
nand UO_2084 (O_2084,N_19699,N_19680);
or UO_2085 (O_2085,N_19701,N_19809);
and UO_2086 (O_2086,N_19698,N_19814);
and UO_2087 (O_2087,N_19967,N_19819);
and UO_2088 (O_2088,N_19631,N_19690);
and UO_2089 (O_2089,N_19524,N_19862);
nand UO_2090 (O_2090,N_19685,N_19823);
or UO_2091 (O_2091,N_19884,N_19611);
and UO_2092 (O_2092,N_19972,N_19834);
nand UO_2093 (O_2093,N_19580,N_19759);
and UO_2094 (O_2094,N_19867,N_19737);
nor UO_2095 (O_2095,N_19640,N_19842);
nor UO_2096 (O_2096,N_19769,N_19586);
or UO_2097 (O_2097,N_19977,N_19914);
nand UO_2098 (O_2098,N_19980,N_19768);
nor UO_2099 (O_2099,N_19910,N_19831);
and UO_2100 (O_2100,N_19860,N_19689);
or UO_2101 (O_2101,N_19828,N_19564);
or UO_2102 (O_2102,N_19798,N_19511);
nand UO_2103 (O_2103,N_19651,N_19946);
nand UO_2104 (O_2104,N_19987,N_19912);
and UO_2105 (O_2105,N_19903,N_19514);
or UO_2106 (O_2106,N_19892,N_19948);
nand UO_2107 (O_2107,N_19594,N_19928);
nand UO_2108 (O_2108,N_19574,N_19586);
nor UO_2109 (O_2109,N_19677,N_19757);
nand UO_2110 (O_2110,N_19526,N_19559);
nor UO_2111 (O_2111,N_19930,N_19861);
or UO_2112 (O_2112,N_19674,N_19677);
nor UO_2113 (O_2113,N_19829,N_19838);
nor UO_2114 (O_2114,N_19834,N_19661);
nor UO_2115 (O_2115,N_19587,N_19504);
nor UO_2116 (O_2116,N_19668,N_19724);
nor UO_2117 (O_2117,N_19676,N_19576);
and UO_2118 (O_2118,N_19929,N_19525);
nor UO_2119 (O_2119,N_19822,N_19935);
and UO_2120 (O_2120,N_19789,N_19629);
and UO_2121 (O_2121,N_19774,N_19522);
nand UO_2122 (O_2122,N_19882,N_19633);
and UO_2123 (O_2123,N_19701,N_19723);
nand UO_2124 (O_2124,N_19726,N_19962);
and UO_2125 (O_2125,N_19550,N_19830);
nor UO_2126 (O_2126,N_19785,N_19991);
nand UO_2127 (O_2127,N_19676,N_19953);
nand UO_2128 (O_2128,N_19817,N_19591);
or UO_2129 (O_2129,N_19649,N_19754);
and UO_2130 (O_2130,N_19526,N_19638);
or UO_2131 (O_2131,N_19548,N_19535);
or UO_2132 (O_2132,N_19780,N_19664);
nand UO_2133 (O_2133,N_19749,N_19669);
nor UO_2134 (O_2134,N_19918,N_19544);
and UO_2135 (O_2135,N_19684,N_19787);
nor UO_2136 (O_2136,N_19633,N_19854);
nor UO_2137 (O_2137,N_19861,N_19926);
nand UO_2138 (O_2138,N_19618,N_19913);
nand UO_2139 (O_2139,N_19547,N_19600);
and UO_2140 (O_2140,N_19993,N_19815);
or UO_2141 (O_2141,N_19746,N_19843);
or UO_2142 (O_2142,N_19709,N_19721);
and UO_2143 (O_2143,N_19694,N_19693);
and UO_2144 (O_2144,N_19700,N_19712);
and UO_2145 (O_2145,N_19607,N_19850);
and UO_2146 (O_2146,N_19748,N_19618);
or UO_2147 (O_2147,N_19985,N_19710);
nor UO_2148 (O_2148,N_19559,N_19750);
or UO_2149 (O_2149,N_19759,N_19849);
nor UO_2150 (O_2150,N_19661,N_19874);
nor UO_2151 (O_2151,N_19537,N_19775);
nor UO_2152 (O_2152,N_19582,N_19829);
or UO_2153 (O_2153,N_19550,N_19500);
and UO_2154 (O_2154,N_19952,N_19953);
nand UO_2155 (O_2155,N_19506,N_19559);
and UO_2156 (O_2156,N_19772,N_19856);
nor UO_2157 (O_2157,N_19953,N_19685);
nand UO_2158 (O_2158,N_19782,N_19982);
and UO_2159 (O_2159,N_19987,N_19764);
or UO_2160 (O_2160,N_19560,N_19999);
nor UO_2161 (O_2161,N_19992,N_19883);
and UO_2162 (O_2162,N_19512,N_19636);
or UO_2163 (O_2163,N_19936,N_19687);
or UO_2164 (O_2164,N_19562,N_19828);
or UO_2165 (O_2165,N_19640,N_19650);
or UO_2166 (O_2166,N_19528,N_19709);
or UO_2167 (O_2167,N_19558,N_19956);
nor UO_2168 (O_2168,N_19938,N_19692);
xnor UO_2169 (O_2169,N_19620,N_19860);
nor UO_2170 (O_2170,N_19763,N_19601);
nand UO_2171 (O_2171,N_19704,N_19898);
nand UO_2172 (O_2172,N_19990,N_19623);
and UO_2173 (O_2173,N_19823,N_19802);
nor UO_2174 (O_2174,N_19995,N_19742);
nand UO_2175 (O_2175,N_19820,N_19748);
nor UO_2176 (O_2176,N_19908,N_19805);
and UO_2177 (O_2177,N_19875,N_19767);
and UO_2178 (O_2178,N_19632,N_19708);
nand UO_2179 (O_2179,N_19572,N_19646);
xor UO_2180 (O_2180,N_19525,N_19591);
and UO_2181 (O_2181,N_19907,N_19918);
nand UO_2182 (O_2182,N_19777,N_19731);
and UO_2183 (O_2183,N_19706,N_19731);
or UO_2184 (O_2184,N_19520,N_19981);
or UO_2185 (O_2185,N_19810,N_19930);
or UO_2186 (O_2186,N_19821,N_19987);
and UO_2187 (O_2187,N_19925,N_19945);
nand UO_2188 (O_2188,N_19510,N_19927);
and UO_2189 (O_2189,N_19651,N_19693);
nand UO_2190 (O_2190,N_19614,N_19606);
or UO_2191 (O_2191,N_19512,N_19537);
nand UO_2192 (O_2192,N_19967,N_19957);
and UO_2193 (O_2193,N_19742,N_19925);
or UO_2194 (O_2194,N_19798,N_19721);
nand UO_2195 (O_2195,N_19504,N_19572);
nand UO_2196 (O_2196,N_19833,N_19839);
or UO_2197 (O_2197,N_19659,N_19657);
or UO_2198 (O_2198,N_19723,N_19958);
or UO_2199 (O_2199,N_19535,N_19776);
nand UO_2200 (O_2200,N_19689,N_19909);
or UO_2201 (O_2201,N_19658,N_19848);
nor UO_2202 (O_2202,N_19584,N_19638);
nor UO_2203 (O_2203,N_19634,N_19703);
or UO_2204 (O_2204,N_19536,N_19561);
or UO_2205 (O_2205,N_19683,N_19714);
nor UO_2206 (O_2206,N_19701,N_19924);
nor UO_2207 (O_2207,N_19545,N_19631);
or UO_2208 (O_2208,N_19661,N_19508);
and UO_2209 (O_2209,N_19652,N_19855);
nor UO_2210 (O_2210,N_19513,N_19828);
xnor UO_2211 (O_2211,N_19737,N_19561);
and UO_2212 (O_2212,N_19667,N_19617);
nor UO_2213 (O_2213,N_19845,N_19945);
or UO_2214 (O_2214,N_19650,N_19550);
or UO_2215 (O_2215,N_19679,N_19970);
and UO_2216 (O_2216,N_19549,N_19894);
or UO_2217 (O_2217,N_19886,N_19653);
nand UO_2218 (O_2218,N_19987,N_19743);
or UO_2219 (O_2219,N_19534,N_19617);
or UO_2220 (O_2220,N_19709,N_19704);
and UO_2221 (O_2221,N_19893,N_19657);
or UO_2222 (O_2222,N_19668,N_19876);
nor UO_2223 (O_2223,N_19587,N_19758);
or UO_2224 (O_2224,N_19539,N_19508);
and UO_2225 (O_2225,N_19940,N_19796);
and UO_2226 (O_2226,N_19784,N_19684);
nor UO_2227 (O_2227,N_19796,N_19536);
or UO_2228 (O_2228,N_19636,N_19595);
nand UO_2229 (O_2229,N_19889,N_19675);
nand UO_2230 (O_2230,N_19690,N_19604);
nor UO_2231 (O_2231,N_19714,N_19565);
nand UO_2232 (O_2232,N_19577,N_19740);
and UO_2233 (O_2233,N_19748,N_19672);
or UO_2234 (O_2234,N_19788,N_19769);
and UO_2235 (O_2235,N_19953,N_19745);
or UO_2236 (O_2236,N_19826,N_19643);
and UO_2237 (O_2237,N_19727,N_19773);
and UO_2238 (O_2238,N_19654,N_19638);
and UO_2239 (O_2239,N_19720,N_19812);
nor UO_2240 (O_2240,N_19517,N_19594);
nor UO_2241 (O_2241,N_19559,N_19959);
nand UO_2242 (O_2242,N_19569,N_19895);
or UO_2243 (O_2243,N_19939,N_19946);
xor UO_2244 (O_2244,N_19886,N_19818);
and UO_2245 (O_2245,N_19731,N_19551);
and UO_2246 (O_2246,N_19535,N_19806);
nor UO_2247 (O_2247,N_19832,N_19528);
nor UO_2248 (O_2248,N_19609,N_19896);
and UO_2249 (O_2249,N_19788,N_19976);
and UO_2250 (O_2250,N_19815,N_19667);
nand UO_2251 (O_2251,N_19939,N_19811);
nand UO_2252 (O_2252,N_19508,N_19578);
and UO_2253 (O_2253,N_19528,N_19839);
nor UO_2254 (O_2254,N_19726,N_19673);
or UO_2255 (O_2255,N_19799,N_19604);
or UO_2256 (O_2256,N_19544,N_19559);
and UO_2257 (O_2257,N_19646,N_19574);
or UO_2258 (O_2258,N_19666,N_19550);
and UO_2259 (O_2259,N_19790,N_19756);
and UO_2260 (O_2260,N_19883,N_19774);
nand UO_2261 (O_2261,N_19918,N_19639);
nand UO_2262 (O_2262,N_19737,N_19504);
or UO_2263 (O_2263,N_19809,N_19870);
or UO_2264 (O_2264,N_19991,N_19728);
and UO_2265 (O_2265,N_19841,N_19748);
and UO_2266 (O_2266,N_19782,N_19880);
nand UO_2267 (O_2267,N_19866,N_19634);
and UO_2268 (O_2268,N_19738,N_19781);
nand UO_2269 (O_2269,N_19964,N_19992);
or UO_2270 (O_2270,N_19718,N_19935);
and UO_2271 (O_2271,N_19734,N_19598);
nor UO_2272 (O_2272,N_19765,N_19885);
nand UO_2273 (O_2273,N_19788,N_19506);
and UO_2274 (O_2274,N_19603,N_19903);
nor UO_2275 (O_2275,N_19992,N_19723);
nand UO_2276 (O_2276,N_19812,N_19651);
and UO_2277 (O_2277,N_19962,N_19660);
and UO_2278 (O_2278,N_19603,N_19983);
or UO_2279 (O_2279,N_19723,N_19608);
nand UO_2280 (O_2280,N_19868,N_19979);
nor UO_2281 (O_2281,N_19760,N_19748);
nand UO_2282 (O_2282,N_19860,N_19850);
or UO_2283 (O_2283,N_19792,N_19737);
and UO_2284 (O_2284,N_19647,N_19533);
nand UO_2285 (O_2285,N_19786,N_19872);
nand UO_2286 (O_2286,N_19553,N_19536);
nor UO_2287 (O_2287,N_19666,N_19605);
or UO_2288 (O_2288,N_19504,N_19926);
or UO_2289 (O_2289,N_19962,N_19815);
nor UO_2290 (O_2290,N_19794,N_19784);
nand UO_2291 (O_2291,N_19553,N_19758);
xor UO_2292 (O_2292,N_19822,N_19536);
and UO_2293 (O_2293,N_19530,N_19644);
nor UO_2294 (O_2294,N_19549,N_19664);
nand UO_2295 (O_2295,N_19826,N_19685);
and UO_2296 (O_2296,N_19908,N_19947);
nor UO_2297 (O_2297,N_19573,N_19732);
nand UO_2298 (O_2298,N_19743,N_19590);
nor UO_2299 (O_2299,N_19999,N_19765);
or UO_2300 (O_2300,N_19740,N_19920);
or UO_2301 (O_2301,N_19734,N_19942);
or UO_2302 (O_2302,N_19735,N_19742);
nor UO_2303 (O_2303,N_19596,N_19553);
and UO_2304 (O_2304,N_19504,N_19789);
and UO_2305 (O_2305,N_19909,N_19526);
nor UO_2306 (O_2306,N_19936,N_19684);
nor UO_2307 (O_2307,N_19922,N_19964);
or UO_2308 (O_2308,N_19869,N_19638);
nand UO_2309 (O_2309,N_19929,N_19837);
and UO_2310 (O_2310,N_19981,N_19959);
or UO_2311 (O_2311,N_19785,N_19619);
nand UO_2312 (O_2312,N_19792,N_19721);
or UO_2313 (O_2313,N_19951,N_19835);
and UO_2314 (O_2314,N_19653,N_19840);
nor UO_2315 (O_2315,N_19760,N_19536);
and UO_2316 (O_2316,N_19633,N_19619);
and UO_2317 (O_2317,N_19926,N_19651);
and UO_2318 (O_2318,N_19658,N_19838);
or UO_2319 (O_2319,N_19812,N_19512);
or UO_2320 (O_2320,N_19535,N_19780);
nor UO_2321 (O_2321,N_19551,N_19726);
or UO_2322 (O_2322,N_19711,N_19799);
or UO_2323 (O_2323,N_19748,N_19664);
and UO_2324 (O_2324,N_19795,N_19781);
or UO_2325 (O_2325,N_19992,N_19969);
nand UO_2326 (O_2326,N_19742,N_19623);
or UO_2327 (O_2327,N_19774,N_19621);
or UO_2328 (O_2328,N_19591,N_19854);
and UO_2329 (O_2329,N_19603,N_19647);
or UO_2330 (O_2330,N_19685,N_19516);
nand UO_2331 (O_2331,N_19655,N_19829);
nor UO_2332 (O_2332,N_19696,N_19974);
nor UO_2333 (O_2333,N_19913,N_19673);
or UO_2334 (O_2334,N_19982,N_19992);
nand UO_2335 (O_2335,N_19767,N_19880);
and UO_2336 (O_2336,N_19684,N_19793);
or UO_2337 (O_2337,N_19532,N_19997);
and UO_2338 (O_2338,N_19614,N_19678);
nand UO_2339 (O_2339,N_19825,N_19541);
nor UO_2340 (O_2340,N_19667,N_19824);
and UO_2341 (O_2341,N_19930,N_19782);
or UO_2342 (O_2342,N_19914,N_19744);
xnor UO_2343 (O_2343,N_19622,N_19671);
nor UO_2344 (O_2344,N_19900,N_19989);
or UO_2345 (O_2345,N_19810,N_19785);
and UO_2346 (O_2346,N_19883,N_19890);
and UO_2347 (O_2347,N_19828,N_19580);
and UO_2348 (O_2348,N_19571,N_19737);
nor UO_2349 (O_2349,N_19695,N_19830);
and UO_2350 (O_2350,N_19931,N_19823);
or UO_2351 (O_2351,N_19622,N_19624);
and UO_2352 (O_2352,N_19523,N_19660);
or UO_2353 (O_2353,N_19651,N_19594);
nand UO_2354 (O_2354,N_19684,N_19517);
nor UO_2355 (O_2355,N_19534,N_19695);
and UO_2356 (O_2356,N_19729,N_19574);
nand UO_2357 (O_2357,N_19609,N_19746);
nand UO_2358 (O_2358,N_19890,N_19929);
nor UO_2359 (O_2359,N_19848,N_19842);
and UO_2360 (O_2360,N_19523,N_19904);
and UO_2361 (O_2361,N_19522,N_19726);
and UO_2362 (O_2362,N_19774,N_19567);
nand UO_2363 (O_2363,N_19610,N_19501);
and UO_2364 (O_2364,N_19731,N_19720);
nand UO_2365 (O_2365,N_19606,N_19778);
and UO_2366 (O_2366,N_19533,N_19836);
or UO_2367 (O_2367,N_19875,N_19917);
nand UO_2368 (O_2368,N_19985,N_19983);
and UO_2369 (O_2369,N_19516,N_19556);
and UO_2370 (O_2370,N_19855,N_19573);
or UO_2371 (O_2371,N_19731,N_19657);
nor UO_2372 (O_2372,N_19658,N_19667);
nand UO_2373 (O_2373,N_19650,N_19985);
and UO_2374 (O_2374,N_19676,N_19987);
nand UO_2375 (O_2375,N_19975,N_19647);
and UO_2376 (O_2376,N_19744,N_19794);
and UO_2377 (O_2377,N_19598,N_19533);
nor UO_2378 (O_2378,N_19525,N_19977);
and UO_2379 (O_2379,N_19993,N_19997);
and UO_2380 (O_2380,N_19644,N_19594);
and UO_2381 (O_2381,N_19559,N_19860);
or UO_2382 (O_2382,N_19898,N_19617);
nor UO_2383 (O_2383,N_19530,N_19503);
nor UO_2384 (O_2384,N_19814,N_19535);
and UO_2385 (O_2385,N_19684,N_19536);
nor UO_2386 (O_2386,N_19669,N_19849);
or UO_2387 (O_2387,N_19663,N_19758);
and UO_2388 (O_2388,N_19838,N_19925);
and UO_2389 (O_2389,N_19903,N_19564);
nand UO_2390 (O_2390,N_19855,N_19552);
nand UO_2391 (O_2391,N_19900,N_19994);
nand UO_2392 (O_2392,N_19955,N_19587);
and UO_2393 (O_2393,N_19900,N_19574);
nand UO_2394 (O_2394,N_19811,N_19546);
nor UO_2395 (O_2395,N_19553,N_19845);
nor UO_2396 (O_2396,N_19992,N_19798);
and UO_2397 (O_2397,N_19765,N_19801);
nand UO_2398 (O_2398,N_19737,N_19704);
or UO_2399 (O_2399,N_19542,N_19505);
nor UO_2400 (O_2400,N_19604,N_19730);
or UO_2401 (O_2401,N_19571,N_19606);
and UO_2402 (O_2402,N_19663,N_19890);
or UO_2403 (O_2403,N_19830,N_19649);
nor UO_2404 (O_2404,N_19568,N_19614);
and UO_2405 (O_2405,N_19932,N_19618);
nor UO_2406 (O_2406,N_19525,N_19900);
nand UO_2407 (O_2407,N_19945,N_19544);
nor UO_2408 (O_2408,N_19530,N_19924);
nand UO_2409 (O_2409,N_19647,N_19804);
or UO_2410 (O_2410,N_19781,N_19689);
nor UO_2411 (O_2411,N_19712,N_19974);
nand UO_2412 (O_2412,N_19839,N_19960);
nor UO_2413 (O_2413,N_19794,N_19949);
nor UO_2414 (O_2414,N_19851,N_19501);
or UO_2415 (O_2415,N_19834,N_19822);
or UO_2416 (O_2416,N_19880,N_19571);
or UO_2417 (O_2417,N_19605,N_19711);
nor UO_2418 (O_2418,N_19522,N_19826);
nand UO_2419 (O_2419,N_19634,N_19742);
and UO_2420 (O_2420,N_19907,N_19950);
and UO_2421 (O_2421,N_19520,N_19541);
nor UO_2422 (O_2422,N_19951,N_19923);
nor UO_2423 (O_2423,N_19606,N_19655);
or UO_2424 (O_2424,N_19936,N_19691);
nor UO_2425 (O_2425,N_19675,N_19996);
nand UO_2426 (O_2426,N_19936,N_19524);
xnor UO_2427 (O_2427,N_19523,N_19938);
and UO_2428 (O_2428,N_19838,N_19628);
and UO_2429 (O_2429,N_19769,N_19904);
nand UO_2430 (O_2430,N_19709,N_19580);
nor UO_2431 (O_2431,N_19814,N_19712);
nand UO_2432 (O_2432,N_19832,N_19740);
nand UO_2433 (O_2433,N_19816,N_19576);
and UO_2434 (O_2434,N_19854,N_19894);
or UO_2435 (O_2435,N_19782,N_19621);
nor UO_2436 (O_2436,N_19893,N_19685);
nand UO_2437 (O_2437,N_19593,N_19689);
nand UO_2438 (O_2438,N_19704,N_19561);
or UO_2439 (O_2439,N_19776,N_19903);
nor UO_2440 (O_2440,N_19932,N_19891);
and UO_2441 (O_2441,N_19604,N_19756);
nand UO_2442 (O_2442,N_19788,N_19650);
or UO_2443 (O_2443,N_19505,N_19932);
nor UO_2444 (O_2444,N_19792,N_19520);
nand UO_2445 (O_2445,N_19646,N_19712);
nor UO_2446 (O_2446,N_19802,N_19919);
and UO_2447 (O_2447,N_19644,N_19702);
and UO_2448 (O_2448,N_19895,N_19969);
nand UO_2449 (O_2449,N_19671,N_19752);
or UO_2450 (O_2450,N_19833,N_19602);
nor UO_2451 (O_2451,N_19578,N_19625);
nand UO_2452 (O_2452,N_19749,N_19622);
nand UO_2453 (O_2453,N_19620,N_19830);
or UO_2454 (O_2454,N_19685,N_19654);
and UO_2455 (O_2455,N_19982,N_19616);
and UO_2456 (O_2456,N_19723,N_19517);
nand UO_2457 (O_2457,N_19919,N_19805);
and UO_2458 (O_2458,N_19899,N_19792);
nor UO_2459 (O_2459,N_19693,N_19976);
nor UO_2460 (O_2460,N_19700,N_19605);
or UO_2461 (O_2461,N_19794,N_19887);
nor UO_2462 (O_2462,N_19743,N_19585);
and UO_2463 (O_2463,N_19988,N_19582);
nand UO_2464 (O_2464,N_19972,N_19971);
or UO_2465 (O_2465,N_19922,N_19634);
or UO_2466 (O_2466,N_19524,N_19657);
and UO_2467 (O_2467,N_19714,N_19527);
or UO_2468 (O_2468,N_19699,N_19633);
and UO_2469 (O_2469,N_19919,N_19663);
nor UO_2470 (O_2470,N_19590,N_19562);
and UO_2471 (O_2471,N_19839,N_19959);
nor UO_2472 (O_2472,N_19830,N_19925);
or UO_2473 (O_2473,N_19967,N_19577);
or UO_2474 (O_2474,N_19510,N_19555);
or UO_2475 (O_2475,N_19564,N_19701);
nand UO_2476 (O_2476,N_19646,N_19885);
and UO_2477 (O_2477,N_19929,N_19800);
nand UO_2478 (O_2478,N_19558,N_19905);
and UO_2479 (O_2479,N_19886,N_19956);
nand UO_2480 (O_2480,N_19628,N_19678);
or UO_2481 (O_2481,N_19958,N_19546);
nand UO_2482 (O_2482,N_19773,N_19701);
nand UO_2483 (O_2483,N_19734,N_19611);
or UO_2484 (O_2484,N_19743,N_19822);
and UO_2485 (O_2485,N_19590,N_19516);
nor UO_2486 (O_2486,N_19924,N_19636);
nor UO_2487 (O_2487,N_19966,N_19877);
nand UO_2488 (O_2488,N_19644,N_19855);
nor UO_2489 (O_2489,N_19537,N_19875);
or UO_2490 (O_2490,N_19715,N_19824);
and UO_2491 (O_2491,N_19851,N_19619);
and UO_2492 (O_2492,N_19861,N_19724);
nand UO_2493 (O_2493,N_19724,N_19554);
or UO_2494 (O_2494,N_19903,N_19937);
or UO_2495 (O_2495,N_19831,N_19995);
or UO_2496 (O_2496,N_19654,N_19935);
nand UO_2497 (O_2497,N_19655,N_19554);
nand UO_2498 (O_2498,N_19653,N_19900);
or UO_2499 (O_2499,N_19639,N_19923);
endmodule