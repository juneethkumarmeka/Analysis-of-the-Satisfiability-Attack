module basic_5000_50000_5000_100_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_731,In_4620);
or U1 (N_1,In_2641,In_2340);
or U2 (N_2,In_1245,In_4260);
or U3 (N_3,In_4799,In_290);
and U4 (N_4,In_2350,In_4793);
nand U5 (N_5,In_592,In_4494);
and U6 (N_6,In_3069,In_4445);
nor U7 (N_7,In_765,In_3297);
xor U8 (N_8,In_3369,In_581);
or U9 (N_9,In_4004,In_3557);
xor U10 (N_10,In_104,In_4606);
and U11 (N_11,In_4283,In_1054);
nand U12 (N_12,In_3517,In_4390);
xor U13 (N_13,In_1661,In_1573);
and U14 (N_14,In_3026,In_1780);
xor U15 (N_15,In_4427,In_2649);
xnor U16 (N_16,In_1428,In_1451);
nor U17 (N_17,In_2258,In_4495);
and U18 (N_18,In_3308,In_1420);
xnor U19 (N_19,In_469,In_3251);
or U20 (N_20,In_1691,In_3351);
and U21 (N_21,In_435,In_445);
and U22 (N_22,In_1898,In_1916);
or U23 (N_23,In_4994,In_3003);
xor U24 (N_24,In_4790,In_798);
nor U25 (N_25,In_3712,In_2661);
xnor U26 (N_26,In_3994,In_430);
xnor U27 (N_27,In_4281,In_2458);
xnor U28 (N_28,In_498,In_478);
nor U29 (N_29,In_800,In_194);
and U30 (N_30,In_1777,In_420);
xnor U31 (N_31,In_3671,In_4855);
nor U32 (N_32,In_1453,In_2611);
or U33 (N_33,In_4212,In_2363);
xor U34 (N_34,In_1045,In_4282);
xor U35 (N_35,In_2370,In_2738);
nand U36 (N_36,In_1183,In_1943);
xnor U37 (N_37,In_1776,In_449);
nor U38 (N_38,In_3818,In_4755);
or U39 (N_39,In_3909,In_2797);
and U40 (N_40,In_1019,In_145);
or U41 (N_41,In_990,In_4277);
nor U42 (N_42,In_3244,In_801);
nor U43 (N_43,In_3809,In_551);
xnor U44 (N_44,In_3408,In_4584);
and U45 (N_45,In_3017,In_4866);
and U46 (N_46,In_1624,In_3625);
or U47 (N_47,In_1538,In_2352);
nor U48 (N_48,In_2506,In_2076);
xor U49 (N_49,In_3180,In_540);
or U50 (N_50,In_1031,In_804);
nor U51 (N_51,In_233,In_2986);
or U52 (N_52,In_2440,In_3225);
xor U53 (N_53,In_2090,In_4334);
or U54 (N_54,In_1528,In_1440);
or U55 (N_55,In_2201,In_1036);
nor U56 (N_56,In_4108,In_319);
and U57 (N_57,In_681,In_3572);
nand U58 (N_58,In_3025,In_1846);
nand U59 (N_59,In_2502,In_41);
xor U60 (N_60,In_4264,In_944);
xor U61 (N_61,In_2106,In_4347);
nor U62 (N_62,In_96,In_4090);
and U63 (N_63,In_1973,In_617);
and U64 (N_64,In_379,In_958);
nand U65 (N_65,In_2803,In_4549);
or U66 (N_66,In_1713,In_1734);
and U67 (N_67,In_156,In_3460);
and U68 (N_68,In_3159,In_1864);
or U69 (N_69,In_2313,In_3824);
xor U70 (N_70,In_2407,In_1417);
nand U71 (N_71,In_499,In_2992);
nor U72 (N_72,In_2279,In_3758);
or U73 (N_73,In_682,In_719);
or U74 (N_74,In_336,In_3558);
nor U75 (N_75,In_3386,In_4517);
nor U76 (N_76,In_1291,In_2474);
or U77 (N_77,In_458,In_4024);
or U78 (N_78,In_1845,In_3704);
nor U79 (N_79,In_133,In_4422);
or U80 (N_80,In_246,In_1379);
or U81 (N_81,In_1458,In_1304);
nand U82 (N_82,In_3998,In_2442);
or U83 (N_83,In_454,In_4993);
nand U84 (N_84,In_1210,In_4527);
nand U85 (N_85,In_170,In_4167);
and U86 (N_86,In_1491,In_1415);
nand U87 (N_87,In_4311,In_63);
and U88 (N_88,In_2063,In_3525);
nor U89 (N_89,In_512,In_1231);
nor U90 (N_90,In_2037,In_1197);
or U91 (N_91,In_314,In_1191);
xnor U92 (N_92,In_2403,In_3198);
and U93 (N_93,In_2957,In_2745);
nor U94 (N_94,In_3237,In_1771);
xor U95 (N_95,In_1312,In_2102);
nand U96 (N_96,In_2118,In_2445);
nor U97 (N_97,In_875,In_425);
nor U98 (N_98,In_2470,In_3102);
xor U99 (N_99,In_3469,In_4098);
and U100 (N_100,In_8,In_3637);
nor U101 (N_101,In_4101,In_4275);
nor U102 (N_102,In_4752,In_2364);
nand U103 (N_103,In_4384,In_3729);
xor U104 (N_104,In_1341,In_966);
nand U105 (N_105,In_1619,In_189);
or U106 (N_106,In_4178,In_4516);
nor U107 (N_107,In_271,In_2113);
xor U108 (N_108,In_1112,In_120);
and U109 (N_109,In_548,In_3732);
or U110 (N_110,In_2507,In_2938);
and U111 (N_111,In_2375,In_1370);
nand U112 (N_112,In_4883,In_1232);
nand U113 (N_113,In_1480,In_963);
or U114 (N_114,In_2717,In_1295);
nand U115 (N_115,In_4986,In_2761);
xor U116 (N_116,In_3040,In_1686);
and U117 (N_117,In_1648,In_4915);
or U118 (N_118,In_821,In_3510);
nand U119 (N_119,In_2225,In_4195);
nand U120 (N_120,In_2633,In_3784);
or U121 (N_121,In_310,In_1882);
xnor U122 (N_122,In_4204,In_2389);
xnor U123 (N_123,In_1052,In_556);
or U124 (N_124,In_3427,In_1187);
xnor U125 (N_125,In_4289,In_3163);
and U126 (N_126,In_3654,In_2110);
nor U127 (N_127,In_1710,In_3128);
xor U128 (N_128,In_619,In_4411);
nor U129 (N_129,In_1283,In_4571);
and U130 (N_130,In_1336,In_470);
and U131 (N_131,In_2744,In_1506);
and U132 (N_132,In_4135,In_3344);
nand U133 (N_133,In_642,In_1023);
xor U134 (N_134,In_3433,In_1501);
or U135 (N_135,In_2792,In_4647);
and U136 (N_136,In_3452,In_4969);
xnor U137 (N_137,In_659,In_3161);
nand U138 (N_138,In_4019,In_1723);
nand U139 (N_139,In_1028,In_2590);
nor U140 (N_140,In_2381,In_3752);
nor U141 (N_141,In_2259,In_345);
xor U142 (N_142,In_2295,In_224);
nor U143 (N_143,In_2368,In_4632);
nor U144 (N_144,In_1891,In_2007);
and U145 (N_145,In_2194,In_2322);
xor U146 (N_146,In_3630,In_1721);
and U147 (N_147,In_4326,In_2701);
nor U148 (N_148,In_2487,In_3717);
and U149 (N_149,In_25,In_4707);
and U150 (N_150,In_2480,In_3219);
or U151 (N_151,In_1027,In_3530);
nand U152 (N_152,In_2786,In_1152);
nor U153 (N_153,In_4984,In_1629);
and U154 (N_154,In_1168,In_4722);
or U155 (N_155,In_1137,In_1783);
and U156 (N_156,In_3489,In_455);
or U157 (N_157,In_3772,In_2139);
xnor U158 (N_158,In_555,In_1014);
nand U159 (N_159,In_3294,In_3734);
or U160 (N_160,In_466,In_616);
and U161 (N_161,In_4745,In_44);
xor U162 (N_162,In_1806,In_213);
xnor U163 (N_163,In_1055,In_4600);
nand U164 (N_164,In_1349,In_2134);
nor U165 (N_165,In_1466,In_1794);
or U166 (N_166,In_2847,In_2149);
nor U167 (N_167,In_706,In_2568);
xor U168 (N_168,In_601,In_927);
or U169 (N_169,In_1472,In_221);
nand U170 (N_170,In_3569,In_3259);
or U171 (N_171,In_2861,In_1994);
and U172 (N_172,In_2299,In_741);
xor U173 (N_173,In_3399,In_1442);
nor U174 (N_174,In_3691,In_2962);
nor U175 (N_175,In_885,In_3721);
and U176 (N_176,In_1211,In_4359);
and U177 (N_177,In_173,In_951);
nor U178 (N_178,In_3971,In_2123);
and U179 (N_179,In_3126,In_4845);
xor U180 (N_180,In_190,In_1171);
nand U181 (N_181,In_1563,In_4618);
and U182 (N_182,In_1526,In_123);
or U183 (N_183,In_1524,In_2539);
xnor U184 (N_184,In_1522,In_978);
and U185 (N_185,In_3580,In_366);
nor U186 (N_186,In_198,In_2509);
or U187 (N_187,In_4579,In_3747);
nand U188 (N_188,In_1747,In_2260);
xor U189 (N_189,In_2970,In_607);
xor U190 (N_190,In_37,In_4307);
xnor U191 (N_191,In_4300,In_1952);
or U192 (N_192,In_3154,In_3289);
xnor U193 (N_193,In_4923,In_2273);
nor U194 (N_194,In_1577,In_31);
xnor U195 (N_195,In_479,In_2443);
xor U196 (N_196,In_3547,In_1178);
nor U197 (N_197,In_2604,In_2706);
nor U198 (N_198,In_1966,In_2203);
and U199 (N_199,In_3107,In_3820);
nand U200 (N_200,In_4137,In_4528);
nand U201 (N_201,In_3829,In_4370);
xnor U202 (N_202,In_768,In_273);
nor U203 (N_203,In_4627,In_3903);
xnor U204 (N_204,In_2163,In_3761);
nor U205 (N_205,In_2573,In_1658);
nor U206 (N_206,In_486,In_47);
nor U207 (N_207,In_3118,In_3108);
or U208 (N_208,In_799,In_250);
xnor U209 (N_209,In_4198,In_2151);
and U210 (N_210,In_612,In_4244);
and U211 (N_211,In_3078,In_3071);
nor U212 (N_212,In_3479,In_2642);
or U213 (N_213,In_1227,In_1249);
or U214 (N_214,In_1585,In_4132);
nor U215 (N_215,In_1987,In_4727);
and U216 (N_216,In_2012,In_3008);
or U217 (N_217,In_4960,In_1770);
nor U218 (N_218,In_152,In_441);
and U219 (N_219,In_1354,In_679);
xnor U220 (N_220,In_934,In_3813);
nor U221 (N_221,In_1956,In_418);
nand U222 (N_222,In_1463,In_2082);
nor U223 (N_223,In_2892,In_2186);
nand U224 (N_224,In_209,In_2955);
nor U225 (N_225,In_4830,In_1058);
nor U226 (N_226,In_1678,In_265);
xor U227 (N_227,In_4958,In_4286);
nand U228 (N_228,In_1228,In_2070);
xnor U229 (N_229,In_2348,In_253);
or U230 (N_230,In_694,In_2906);
or U231 (N_231,In_3565,In_3168);
or U232 (N_232,In_2692,In_1605);
and U233 (N_233,In_4064,In_3715);
xor U234 (N_234,In_4572,In_3674);
and U235 (N_235,In_3816,In_3948);
and U236 (N_236,In_4942,In_2434);
xor U237 (N_237,In_1155,In_4176);
xnor U238 (N_238,In_4642,In_447);
nand U239 (N_239,In_892,In_3002);
nor U240 (N_240,In_2668,In_4483);
and U241 (N_241,In_4497,In_3092);
or U242 (N_242,In_4710,In_1841);
nand U243 (N_243,In_3410,In_4512);
and U244 (N_244,In_810,In_773);
nor U245 (N_245,In_4654,In_2265);
xnor U246 (N_246,In_4846,In_1300);
nand U247 (N_247,In_4777,In_1495);
xor U248 (N_248,In_2280,In_1346);
and U249 (N_249,In_1512,In_627);
nor U250 (N_250,In_3009,In_620);
xor U251 (N_251,In_2612,In_2831);
nor U252 (N_252,In_1550,In_1999);
nand U253 (N_253,In_4189,In_3528);
nor U254 (N_254,In_2083,In_3497);
nor U255 (N_255,In_1953,In_4577);
nand U256 (N_256,In_2215,In_2321);
nor U257 (N_257,In_3760,In_1792);
and U258 (N_258,In_1715,In_1906);
or U259 (N_259,In_1900,In_4037);
and U260 (N_260,In_3390,In_30);
nand U261 (N_261,In_1860,In_4059);
xor U262 (N_262,In_3051,In_3810);
nand U263 (N_263,In_89,In_4086);
xnor U264 (N_264,In_1494,In_1797);
and U265 (N_265,In_2137,In_457);
nand U266 (N_266,In_4522,In_4876);
nand U267 (N_267,In_400,In_1631);
xor U268 (N_268,In_3561,In_3937);
nand U269 (N_269,In_1209,In_439);
nor U270 (N_270,In_2428,In_3455);
xnor U271 (N_271,In_355,In_2989);
and U272 (N_272,In_1340,In_4215);
xnor U273 (N_273,In_4809,In_2143);
nor U274 (N_274,In_354,In_2415);
and U275 (N_275,In_4330,In_2292);
nand U276 (N_276,In_4989,In_1358);
nor U277 (N_277,In_2593,In_3582);
or U278 (N_278,In_2629,In_2705);
xor U279 (N_279,In_2610,In_1339);
nor U280 (N_280,In_4025,In_1077);
xor U281 (N_281,In_1143,In_2896);
nand U282 (N_282,In_1912,In_4997);
nor U283 (N_283,In_3970,In_3856);
nor U284 (N_284,In_2773,In_2859);
or U285 (N_285,In_2990,In_29);
nand U286 (N_286,In_3210,In_4256);
nor U287 (N_287,In_3104,In_4821);
nand U288 (N_288,In_2079,In_4559);
xnor U289 (N_289,In_3591,In_1212);
xor U290 (N_290,In_1311,In_4806);
nand U291 (N_291,In_2144,In_3177);
nor U292 (N_292,In_4336,In_2067);
and U293 (N_293,In_2730,In_2553);
xor U294 (N_294,In_59,In_4177);
and U295 (N_295,In_2595,In_1041);
and U296 (N_296,In_4742,In_3267);
and U297 (N_297,In_1018,In_264);
xor U298 (N_298,In_2704,In_4922);
nor U299 (N_299,In_3743,In_3944);
nor U300 (N_300,In_916,In_4708);
nor U301 (N_301,In_4121,In_753);
or U302 (N_302,In_3663,In_3043);
or U303 (N_303,In_570,In_2103);
xor U304 (N_304,In_1596,In_1892);
nand U305 (N_305,In_3894,In_378);
nand U306 (N_306,In_3788,In_4931);
nand U307 (N_307,In_3187,In_4099);
nor U308 (N_308,In_1922,In_2010);
or U309 (N_309,In_1421,In_4791);
nand U310 (N_310,In_4812,In_4168);
xor U311 (N_311,In_4760,In_1432);
and U312 (N_312,In_1962,In_1328);
and U313 (N_313,In_2058,In_868);
nand U314 (N_314,In_384,In_901);
xor U315 (N_315,In_117,In_4697);
or U316 (N_316,In_3919,In_318);
and U317 (N_317,In_1760,In_4951);
or U318 (N_318,In_4506,In_3955);
xor U319 (N_319,In_401,In_4623);
nor U320 (N_320,In_4419,In_1518);
and U321 (N_321,In_3320,In_2623);
nand U322 (N_322,In_3859,In_2882);
xnor U323 (N_323,In_1481,In_889);
or U324 (N_324,In_3462,In_1646);
nor U325 (N_325,In_1179,In_1293);
nand U326 (N_326,In_4655,In_1343);
or U327 (N_327,In_1630,In_3453);
xor U328 (N_328,In_1695,In_72);
and U329 (N_329,In_881,In_234);
or U330 (N_330,In_137,In_614);
nand U331 (N_331,In_4119,In_1753);
or U332 (N_332,In_2444,In_1218);
or U333 (N_333,In_60,In_3030);
xnor U334 (N_334,In_1887,In_181);
nor U335 (N_335,In_2331,In_3623);
nand U336 (N_336,In_3819,In_1359);
or U337 (N_337,In_1690,In_3035);
xor U338 (N_338,In_2314,In_188);
or U339 (N_339,In_4925,In_1119);
nor U340 (N_340,In_2587,In_2323);
nand U341 (N_341,In_576,In_4630);
or U342 (N_342,In_3905,In_1562);
xor U343 (N_343,In_1870,In_2810);
xor U344 (N_344,In_2531,In_4114);
and U345 (N_345,In_703,In_1683);
and U346 (N_346,In_2647,In_1233);
xor U347 (N_347,In_594,In_146);
or U348 (N_348,In_444,In_2920);
and U349 (N_349,In_3087,In_4263);
or U350 (N_350,In_3765,In_1787);
or U351 (N_351,In_3551,In_907);
nor U352 (N_352,In_3740,In_3349);
nor U353 (N_353,In_90,In_184);
nand U354 (N_354,In_1822,In_3151);
xnor U355 (N_355,In_1410,In_1221);
nor U356 (N_356,In_1539,In_3476);
xor U357 (N_357,In_787,In_3302);
nand U358 (N_358,In_3535,In_3534);
or U359 (N_359,In_4852,In_1065);
nor U360 (N_360,In_2697,In_1645);
xor U361 (N_361,In_1251,In_2833);
nand U362 (N_362,In_58,In_3616);
nor U363 (N_363,In_1722,In_1148);
nand U364 (N_364,In_2140,In_1486);
or U365 (N_365,In_1542,In_776);
xnor U366 (N_366,In_1335,In_2011);
nand U367 (N_367,In_4992,In_4658);
and U368 (N_368,In_2249,In_1280);
or U369 (N_369,In_948,In_1190);
and U370 (N_370,In_2605,In_1059);
nand U371 (N_371,In_4629,In_81);
or U372 (N_372,In_1225,In_3389);
xor U373 (N_373,In_3720,In_4148);
or U374 (N_374,In_95,In_4956);
nand U375 (N_375,In_1772,In_4619);
or U376 (N_376,In_3848,In_920);
xor U377 (N_377,In_1653,In_3148);
or U378 (N_378,In_2173,In_3121);
nand U379 (N_379,In_791,In_1213);
and U380 (N_380,In_1735,In_2659);
xor U381 (N_381,In_3446,In_4673);
xnor U382 (N_382,In_895,In_2491);
xnor U383 (N_383,In_4371,In_2236);
nand U384 (N_384,In_501,In_3306);
and U385 (N_385,In_4804,In_942);
xor U386 (N_386,In_3963,In_2358);
xnor U387 (N_387,In_2196,In_482);
and U388 (N_388,In_3432,In_3062);
xnor U389 (N_389,In_392,In_4128);
xnor U390 (N_390,In_1174,In_274);
nor U391 (N_391,In_3340,In_827);
xor U392 (N_392,In_3862,In_4570);
nor U393 (N_393,In_1593,In_4161);
or U394 (N_394,In_403,In_4000);
xor U395 (N_395,In_1220,In_1934);
nor U396 (N_396,In_1600,In_4479);
xor U397 (N_397,In_1356,In_353);
nor U398 (N_398,In_2963,In_4557);
and U399 (N_399,In_3256,In_1732);
nand U400 (N_400,In_4605,In_4920);
nor U401 (N_401,In_3714,In_3444);
nor U402 (N_402,In_671,In_3366);
xor U403 (N_403,In_3440,In_3004);
nand U404 (N_404,In_4917,In_4196);
and U405 (N_405,In_835,In_1242);
and U406 (N_406,In_279,In_537);
or U407 (N_407,In_487,In_1007);
nand U408 (N_408,In_4872,In_4899);
or U409 (N_409,In_292,In_3579);
nor U410 (N_410,In_4368,In_3425);
or U411 (N_411,In_4007,In_1826);
or U412 (N_412,In_2680,In_1241);
or U413 (N_413,In_180,In_846);
nand U414 (N_414,In_1151,In_3304);
xor U415 (N_415,In_2429,In_4814);
and U416 (N_416,In_2126,In_4954);
nand U417 (N_417,In_849,In_2816);
nand U418 (N_418,In_38,In_1849);
and U419 (N_419,In_3207,In_774);
xnor U420 (N_420,In_4729,In_1673);
nand U421 (N_421,In_3238,In_4301);
or U422 (N_422,In_2270,In_3860);
nor U423 (N_423,In_4157,In_1337);
xnor U424 (N_424,In_3834,In_3336);
or U425 (N_425,In_2663,In_3795);
nor U426 (N_426,In_2820,In_2278);
or U427 (N_427,In_3613,In_4662);
nand U428 (N_428,In_483,In_1660);
and U429 (N_429,In_4335,In_866);
and U430 (N_430,In_1157,In_1871);
and U431 (N_431,In_2529,In_1546);
nand U432 (N_432,In_107,In_1382);
or U433 (N_433,In_2341,In_4272);
or U434 (N_434,In_448,In_1561);
or U435 (N_435,In_643,In_1261);
nand U436 (N_436,In_4405,In_3928);
and U437 (N_437,In_3893,In_1099);
xnor U438 (N_438,In_969,In_3622);
nand U439 (N_439,In_4711,In_2987);
or U440 (N_440,In_3814,In_3968);
xnor U441 (N_441,In_4279,In_4604);
nor U442 (N_442,In_2922,In_4893);
or U443 (N_443,In_3539,In_1172);
nand U444 (N_444,In_2361,In_3603);
nand U445 (N_445,In_3388,In_3023);
nor U446 (N_446,In_3633,In_1011);
nor U447 (N_447,In_2893,In_2868);
or U448 (N_448,In_2806,In_3072);
or U449 (N_449,In_102,In_1778);
and U450 (N_450,In_1047,In_4660);
nor U451 (N_451,In_2956,In_4728);
nand U452 (N_452,In_2679,In_4221);
or U453 (N_453,In_33,In_3578);
and U454 (N_454,In_3507,In_3318);
and U455 (N_455,In_4808,In_4113);
nand U456 (N_456,In_1983,In_4996);
nor U457 (N_457,In_707,In_1034);
and U458 (N_458,In_4743,In_3034);
and U459 (N_459,In_85,In_993);
and U460 (N_460,In_4753,In_3438);
nand U461 (N_461,In_1586,In_4910);
nor U462 (N_462,In_4226,In_22);
nor U463 (N_463,In_1613,In_1423);
and U464 (N_464,In_1061,In_943);
nor U465 (N_465,In_4952,In_2645);
and U466 (N_466,In_2253,In_532);
nor U467 (N_467,In_422,In_771);
nand U468 (N_468,In_3398,In_3404);
and U469 (N_469,In_1560,In_3934);
xnor U470 (N_470,In_4703,In_4525);
nor U471 (N_471,In_4935,In_4180);
or U472 (N_472,In_3989,In_4249);
nor U473 (N_473,In_3686,In_2296);
and U474 (N_474,In_4612,In_908);
or U475 (N_475,In_1493,In_3012);
nand U476 (N_476,In_609,In_4932);
xnor U477 (N_477,In_3212,In_2085);
nand U478 (N_478,In_3684,In_1124);
nand U479 (N_479,In_3261,In_186);
xnor U480 (N_480,In_2535,In_4237);
xnor U481 (N_481,In_3531,In_3755);
nand U482 (N_482,In_2513,In_1067);
nand U483 (N_483,In_4832,In_481);
and U484 (N_484,In_2580,In_3575);
xnor U485 (N_485,In_1136,In_1590);
nand U486 (N_486,In_1529,In_2698);
nand U487 (N_487,In_4122,In_135);
nand U488 (N_488,In_756,In_3962);
nand U489 (N_489,In_1044,In_1610);
nor U490 (N_490,In_4415,In_3335);
nand U491 (N_491,In_717,In_2823);
xor U492 (N_492,In_1635,In_495);
nor U493 (N_493,In_3595,In_4058);
xnor U494 (N_494,In_269,In_3113);
xor U495 (N_495,In_3277,In_1122);
nand U496 (N_496,In_1940,In_1697);
and U497 (N_497,In_3123,In_4949);
xnor U498 (N_498,In_4229,In_196);
and U499 (N_499,In_1547,In_4937);
xor U500 (N_500,In_2684,In_1073);
and U501 (N_501,In_3013,In_4125);
xnor U502 (N_502,In_557,N_495);
nand U503 (N_503,In_1872,In_4719);
and U504 (N_504,In_20,In_2822);
and U505 (N_505,In_10,In_2282);
and U506 (N_506,N_426,In_2227);
nor U507 (N_507,In_3769,In_4267);
nand U508 (N_508,In_1075,In_4201);
nor U509 (N_509,In_2667,In_786);
and U510 (N_510,In_3101,N_242);
nand U511 (N_511,In_3536,In_788);
or U512 (N_512,In_3594,In_4568);
xnor U513 (N_513,In_3888,In_1255);
and U514 (N_514,N_391,In_3844);
xnor U515 (N_515,In_3932,In_1671);
nor U516 (N_516,In_1615,In_4181);
nand U517 (N_517,In_764,N_71);
or U518 (N_518,N_223,In_1830);
nor U519 (N_519,In_3434,In_4414);
nor U520 (N_520,In_1572,In_3659);
and U521 (N_521,In_4453,N_345);
xor U522 (N_522,In_4199,N_256);
and U523 (N_523,In_2943,In_428);
xnor U524 (N_524,In_2515,In_591);
xnor U525 (N_525,In_1319,In_3458);
nor U526 (N_526,In_1009,In_844);
nand U527 (N_527,In_3983,In_3640);
and U528 (N_528,In_4325,In_3950);
and U529 (N_529,In_4535,In_4903);
or U530 (N_530,In_3491,In_1127);
and U531 (N_531,In_3858,In_1567);
xnor U532 (N_532,N_474,In_4720);
xnor U533 (N_533,In_2914,In_4555);
nand U534 (N_534,In_3726,N_166);
or U535 (N_535,In_204,In_1755);
and U536 (N_536,N_456,In_4353);
xor U537 (N_537,In_2223,In_3111);
or U538 (N_538,In_1521,N_141);
nor U539 (N_539,N_3,In_1957);
or U540 (N_540,In_516,In_283);
nor U541 (N_541,In_1394,In_3906);
xor U542 (N_542,In_3857,In_174);
xor U543 (N_543,N_179,In_4117);
or U544 (N_544,In_1094,In_3706);
nand U545 (N_545,In_1165,In_4761);
and U546 (N_546,In_4145,In_3874);
nor U547 (N_547,In_931,In_3549);
nand U548 (N_548,In_1926,N_350);
nand U549 (N_549,In_562,In_4164);
or U550 (N_550,In_636,In_1488);
xnor U551 (N_551,In_2499,In_4228);
and U552 (N_552,In_2241,N_151);
nand U553 (N_553,In_2141,In_590);
and U554 (N_554,In_3631,In_4182);
xor U555 (N_555,In_2116,In_489);
and U556 (N_556,N_23,In_2808);
or U557 (N_557,In_1048,In_3406);
and U558 (N_558,In_670,In_2152);
and U559 (N_559,In_2516,In_1523);
or U560 (N_560,In_3585,In_4828);
nor U561 (N_561,In_1651,In_2627);
xnor U562 (N_562,In_4840,In_2237);
or U563 (N_563,In_3355,N_306);
nand U564 (N_564,In_3619,In_127);
nand U565 (N_565,In_573,In_4941);
xor U566 (N_566,N_486,In_2939);
or U567 (N_567,In_4550,N_340);
xor U568 (N_568,In_2760,In_1030);
and U569 (N_569,In_3952,In_4787);
or U570 (N_570,In_4686,In_1142);
or U571 (N_571,In_2660,In_4853);
or U572 (N_572,In_4048,In_2231);
or U573 (N_573,In_3502,In_2589);
nor U574 (N_574,In_2763,In_795);
xnor U575 (N_575,In_1729,In_86);
or U576 (N_576,In_1807,In_4343);
and U577 (N_577,In_4913,In_3307);
xor U578 (N_578,In_3204,N_484);
and U579 (N_579,In_2383,In_3922);
or U580 (N_580,In_4185,In_2162);
nor U581 (N_581,In_3799,N_312);
nor U582 (N_582,In_3339,In_1718);
nor U583 (N_583,N_30,In_3951);
nor U584 (N_584,In_1996,In_3429);
nand U585 (N_585,In_3374,In_3094);
xnor U586 (N_586,In_1855,In_53);
xor U587 (N_587,In_1568,In_1654);
or U588 (N_588,N_387,In_1267);
nand U589 (N_589,In_130,In_1371);
and U590 (N_590,In_1198,In_2379);
nor U591 (N_591,In_1626,N_244);
and U592 (N_592,In_1049,In_2357);
nor U593 (N_593,In_744,In_1080);
xnor U594 (N_594,In_2427,N_294);
and U595 (N_595,In_3213,In_697);
nand U596 (N_596,In_2023,In_4675);
nand U597 (N_597,In_2827,In_4316);
nand U598 (N_598,In_505,N_475);
xor U599 (N_599,In_1680,In_2872);
or U600 (N_600,In_716,In_4026);
nor U601 (N_601,In_3276,In_3786);
nor U602 (N_602,In_2088,In_2302);
nor U603 (N_603,N_75,In_3378);
xnor U604 (N_604,N_487,In_2136);
xor U605 (N_605,In_4582,In_62);
and U606 (N_606,In_3883,In_3195);
or U607 (N_607,In_3960,In_1400);
nand U608 (N_608,In_4597,In_2669);
nor U609 (N_609,In_3007,In_4592);
xor U610 (N_610,In_2671,In_100);
xor U611 (N_611,In_3678,In_730);
or U612 (N_612,In_1991,In_442);
nor U613 (N_613,In_830,In_4039);
or U614 (N_614,N_451,In_3878);
and U615 (N_615,In_4640,In_4936);
xor U616 (N_616,In_3537,In_2133);
or U617 (N_617,In_1696,In_2096);
nor U618 (N_618,In_3300,In_2053);
and U619 (N_619,In_2874,In_2080);
nand U620 (N_620,In_3485,In_2554);
nand U621 (N_621,In_4569,In_1514);
and U622 (N_622,In_2543,In_1789);
and U623 (N_623,In_3606,In_1470);
nor U624 (N_624,In_1821,In_3647);
and U625 (N_625,N_217,In_3559);
xor U626 (N_626,In_2422,In_608);
and U627 (N_627,In_2749,In_1373);
and U628 (N_628,In_2880,In_2873);
and U629 (N_629,In_1464,In_1297);
xnor U630 (N_630,In_1079,In_2387);
xor U631 (N_631,N_397,In_21);
and U632 (N_632,In_2332,In_2670);
nand U633 (N_633,N_485,In_1985);
and U634 (N_634,In_50,In_408);
or U635 (N_635,N_300,In_4447);
and U636 (N_636,N_349,In_4639);
or U637 (N_637,In_2431,In_2490);
nand U638 (N_638,N_342,In_51);
or U639 (N_639,In_550,N_260);
and U640 (N_640,In_1497,In_777);
nor U641 (N_641,In_4778,In_349);
nand U642 (N_642,In_282,In_4624);
or U643 (N_643,In_251,In_1469);
xnor U644 (N_644,N_432,In_3509);
nor U645 (N_645,In_92,In_2864);
nand U646 (N_646,In_4152,In_1450);
nor U647 (N_647,In_962,In_3642);
or U648 (N_648,In_1214,In_4398);
xor U649 (N_649,In_4046,In_926);
and U650 (N_650,In_3312,In_3315);
or U651 (N_651,N_73,N_59);
nor U652 (N_652,In_1634,In_1436);
xnor U653 (N_653,N_493,In_2312);
or U654 (N_654,In_1189,In_3405);
nor U655 (N_655,In_2805,In_2902);
or U656 (N_656,In_3738,In_4222);
nand U657 (N_657,In_1076,N_227);
xor U658 (N_658,In_1802,In_411);
or U659 (N_659,In_4481,In_4551);
xor U660 (N_660,In_2104,In_199);
nor U661 (N_661,In_2787,N_282);
nand U662 (N_662,In_4469,In_3419);
nand U663 (N_663,In_3070,In_3666);
nand U664 (N_664,In_2742,In_49);
and U665 (N_665,In_1445,In_3975);
and U666 (N_666,In_3665,In_3278);
or U667 (N_667,In_633,In_3992);
and U668 (N_668,In_2954,In_1914);
and U669 (N_669,In_3941,In_4027);
nor U670 (N_670,In_2599,In_2598);
nand U671 (N_671,In_4467,In_824);
xor U672 (N_672,In_4354,In_2210);
and U673 (N_673,In_3227,In_845);
nand U674 (N_674,In_1633,N_215);
and U675 (N_675,In_1642,In_453);
nor U676 (N_676,N_24,In_1668);
nor U677 (N_677,In_884,In_1711);
xnor U678 (N_678,In_3424,In_4504);
or U679 (N_679,In_419,In_1186);
nand U680 (N_680,In_940,In_4147);
nand U681 (N_681,In_348,N_467);
nor U682 (N_682,In_3988,N_434);
nand U683 (N_683,In_363,In_1460);
xor U684 (N_684,In_1963,In_3454);
and U685 (N_685,In_2617,In_3759);
and U686 (N_686,In_2586,In_2522);
nor U687 (N_687,In_638,In_4439);
nand U688 (N_688,In_3202,In_3608);
or U689 (N_689,N_332,In_202);
or U690 (N_690,In_329,In_3915);
xnor U691 (N_691,In_247,In_568);
xor U692 (N_692,In_4734,In_970);
nand U693 (N_693,In_586,In_243);
and U694 (N_694,In_2775,In_2496);
or U695 (N_695,In_3965,In_2433);
or U696 (N_696,In_4385,In_4259);
and U697 (N_697,N_238,In_4564);
nor U698 (N_698,In_1150,In_3725);
nand U699 (N_699,In_3334,In_4669);
nor U700 (N_700,In_3626,In_1948);
or U701 (N_701,In_16,In_521);
nor U702 (N_702,In_953,In_4127);
or U703 (N_703,In_3898,In_4313);
nand U704 (N_704,In_1727,N_408);
xnor U705 (N_705,In_1093,In_2951);
or U706 (N_706,In_825,In_2737);
or U707 (N_707,In_834,N_313);
xnor U708 (N_708,In_2266,In_1618);
and U709 (N_709,In_4558,In_3242);
nand U710 (N_710,In_930,In_1589);
nor U711 (N_711,In_291,In_3296);
nor U712 (N_712,In_1230,In_412);
or U713 (N_713,In_3492,In_1184);
nor U714 (N_714,In_2243,In_175);
nor U715 (N_715,In_3041,N_357);
xnor U716 (N_716,In_686,In_3567);
and U717 (N_717,In_3744,In_249);
nor U718 (N_718,In_4010,In_1443);
nand U719 (N_719,In_4268,In_4888);
or U720 (N_720,N_130,In_3215);
nor U721 (N_721,In_806,N_352);
and U722 (N_722,N_374,In_2983);
or U723 (N_723,In_630,In_2965);
and U724 (N_724,In_3478,In_1247);
xor U725 (N_725,In_4451,N_386);
xnor U726 (N_726,In_2703,In_141);
or U727 (N_727,In_3781,In_748);
xnor U728 (N_728,In_4056,In_1986);
nand U729 (N_729,In_1674,N_52);
or U730 (N_730,In_3269,In_1487);
nand U731 (N_731,In_4902,In_3086);
nand U732 (N_732,In_959,In_150);
nor U733 (N_733,In_4914,In_2439);
nand U734 (N_734,In_3196,In_3787);
nor U735 (N_735,In_3605,In_3807);
nand U736 (N_736,In_2547,In_3806);
nand U737 (N_737,In_3855,In_3682);
nor U738 (N_738,In_1046,In_2028);
nor U739 (N_739,In_4638,In_4713);
nand U740 (N_740,In_2320,In_2437);
nor U741 (N_741,N_424,In_4403);
nand U742 (N_742,N_189,In_3480);
nor U743 (N_743,In_1395,In_3867);
xnor U744 (N_744,In_4789,In_887);
nor U745 (N_745,In_4982,N_385);
or U746 (N_746,In_2384,In_2460);
nand U747 (N_747,In_4187,In_4854);
xor U748 (N_748,In_3966,In_2014);
nor U749 (N_749,In_514,N_65);
nand U750 (N_750,In_4169,In_2246);
nor U751 (N_751,In_3423,In_421);
nor U752 (N_752,In_4104,In_1035);
nor U753 (N_753,In_2767,In_66);
nor U754 (N_754,In_995,In_3607);
nor U755 (N_755,In_272,In_1505);
nand U756 (N_756,In_1176,In_1402);
or U757 (N_757,In_2917,In_3628);
and U758 (N_758,In_4008,In_2129);
or U759 (N_759,In_2863,In_3171);
and U760 (N_760,In_4015,In_2532);
nand U761 (N_761,N_347,In_4700);
nand U762 (N_762,In_4454,In_1202);
nand U763 (N_763,In_3545,In_4002);
nand U764 (N_764,In_4455,In_2417);
or U765 (N_765,In_1820,In_1072);
or U766 (N_766,In_4863,In_270);
nand U767 (N_767,In_2638,In_1632);
nand U768 (N_768,In_365,In_3343);
nor U769 (N_769,In_1757,In_1516);
and U770 (N_770,N_239,In_2412);
nor U771 (N_771,In_2190,N_417);
nand U772 (N_772,In_4085,In_3835);
or U773 (N_773,In_1706,In_2526);
or U774 (N_774,In_2182,In_4794);
xor U775 (N_775,In_4593,In_2108);
xnor U776 (N_776,In_303,In_64);
or U777 (N_777,In_3050,In_3014);
xor U778 (N_778,In_814,In_289);
or U779 (N_779,In_779,In_2945);
nor U780 (N_780,In_220,In_1154);
nor U781 (N_781,In_2318,N_112);
nand U782 (N_782,In_2559,In_1852);
nand U783 (N_783,In_2362,In_1286);
or U784 (N_784,In_2338,In_3938);
nand U785 (N_785,In_3586,N_336);
xor U786 (N_786,In_4440,N_490);
and U787 (N_787,In_4733,In_1954);
or U788 (N_788,In_1576,In_3907);
nor U789 (N_789,In_3887,In_1367);
nand U790 (N_790,In_2432,In_496);
nand U791 (N_791,In_1207,N_222);
and U792 (N_792,In_1925,In_3328);
or U793 (N_793,In_98,In_1088);
nor U794 (N_794,In_140,In_1268);
nor U795 (N_795,N_409,In_4251);
or U796 (N_796,In_1108,In_2921);
nor U797 (N_797,In_1303,In_4220);
nor U798 (N_798,In_3015,In_280);
or U799 (N_799,In_702,In_3493);
and U800 (N_800,In_2397,In_2334);
xor U801 (N_801,In_1945,In_361);
or U802 (N_802,In_2187,In_2753);
nor U803 (N_803,In_2727,In_2105);
nor U804 (N_804,In_1431,In_820);
nand U805 (N_805,In_2838,In_649);
or U806 (N_806,In_1978,N_462);
xor U807 (N_807,In_1140,In_1750);
xnor U808 (N_808,In_1074,In_4988);
or U809 (N_809,In_905,In_3570);
nor U810 (N_810,In_4670,In_4363);
or U811 (N_811,In_1050,N_93);
nand U812 (N_812,In_1100,In_3046);
xor U813 (N_813,In_2138,In_1639);
and U814 (N_814,In_3785,In_3233);
xnor U815 (N_815,In_3387,In_3789);
nand U816 (N_816,In_4524,In_4337);
nor U817 (N_817,In_3341,In_124);
nand U818 (N_818,In_4587,In_4140);
xnor U819 (N_819,In_2206,In_1650);
nand U820 (N_820,In_1259,In_1203);
nand U821 (N_821,In_1,In_42);
nor U822 (N_822,In_3815,N_303);
or U823 (N_823,In_3282,In_3719);
xor U824 (N_824,In_1182,In_157);
xor U825 (N_825,In_3653,In_560);
xnor U826 (N_826,In_4921,In_1726);
nor U827 (N_827,N_278,In_4068);
nor U828 (N_828,In_2324,In_337);
nor U829 (N_829,In_4520,In_772);
and U830 (N_830,In_2124,In_1938);
nand U831 (N_831,In_183,In_1201);
and U832 (N_832,In_4744,N_271);
nor U833 (N_833,In_1164,N_246);
nor U834 (N_834,In_3100,In_4172);
or U835 (N_835,In_1502,In_1950);
nor U836 (N_836,N_181,In_976);
or U837 (N_837,In_1038,In_3687);
or U838 (N_838,In_2839,In_2707);
xor U839 (N_839,In_4241,In_2414);
nor U840 (N_840,In_1663,In_464);
and U841 (N_841,In_3381,In_2240);
xnor U842 (N_842,In_1180,In_4437);
or U843 (N_843,In_1138,In_3439);
nand U844 (N_844,In_893,In_1452);
xnor U845 (N_845,In_239,In_212);
nand U846 (N_846,In_2248,In_2915);
nor U847 (N_847,In_4306,In_1944);
and U848 (N_848,N_115,In_472);
and U849 (N_849,In_4069,In_2488);
and U850 (N_850,In_626,In_1156);
nand U851 (N_851,In_1917,In_3403);
nand U852 (N_852,N_68,N_472);
nand U853 (N_853,In_2303,In_1873);
nand U854 (N_854,In_1327,N_245);
or U855 (N_855,N_279,In_2032);
nor U856 (N_856,In_1398,In_4491);
and U857 (N_857,In_4158,N_168);
xor U858 (N_858,In_3754,In_4092);
nor U859 (N_859,In_4238,In_4036);
nor U860 (N_860,In_295,N_310);
or U861 (N_861,In_1265,In_2218);
or U862 (N_862,In_2166,In_1482);
nand U863 (N_863,In_1118,In_4699);
xnor U864 (N_864,In_727,In_4933);
or U865 (N_865,In_503,In_3853);
and U866 (N_866,N_445,In_278);
xor U867 (N_867,In_2029,In_2075);
nand U868 (N_868,In_2211,In_4716);
or U869 (N_869,In_164,In_2495);
xor U870 (N_870,In_4433,In_1575);
xor U871 (N_871,In_2555,N_4);
and U872 (N_872,In_2216,In_3749);
xor U873 (N_873,In_4561,In_2674);
or U874 (N_874,In_3037,In_3953);
and U875 (N_875,In_2446,In_3472);
and U876 (N_876,N_96,N_262);
or U877 (N_877,In_4088,In_604);
xnor U878 (N_878,In_3413,N_492);
nor U879 (N_879,In_2183,In_898);
nand U880 (N_880,In_1854,In_153);
nor U881 (N_881,In_2789,N_182);
and U882 (N_882,In_4436,In_1693);
or U883 (N_883,In_967,In_74);
or U884 (N_884,In_778,In_599);
nand U885 (N_885,In_2024,In_4502);
or U886 (N_886,In_394,N_66);
nor U887 (N_887,In_4252,In_4317);
and U888 (N_888,In_669,In_4702);
and U889 (N_889,In_2448,In_525);
xor U890 (N_890,N_89,In_3876);
or U891 (N_891,In_3257,In_477);
and U892 (N_892,In_2172,In_1439);
or U893 (N_893,In_504,In_2171);
and U894 (N_894,In_1385,In_1989);
xnor U895 (N_895,In_2018,In_3317);
nand U896 (N_896,In_2766,In_2702);
xor U897 (N_897,In_4858,In_1559);
xnor U898 (N_898,In_4545,In_3332);
and U899 (N_899,In_2074,In_3152);
and U900 (N_900,In_3345,N_145);
or U901 (N_901,In_3409,In_1116);
nand U902 (N_902,In_4782,In_4166);
nor U903 (N_903,In_3979,In_4802);
or U904 (N_904,In_522,In_119);
xor U905 (N_905,N_101,In_3393);
or U906 (N_906,In_2916,In_321);
nor U907 (N_907,In_2325,In_2998);
nor U908 (N_908,N_202,In_1017);
nand U909 (N_909,In_4531,In_2114);
nor U910 (N_910,In_2854,In_2783);
nor U911 (N_911,In_40,In_2117);
nand U912 (N_912,In_1459,In_1306);
or U913 (N_913,In_2923,In_575);
nand U914 (N_914,In_3564,In_3822);
nand U915 (N_915,In_2814,In_925);
xnor U916 (N_916,N_309,In_3634);
or U917 (N_917,In_4418,In_735);
xnor U918 (N_918,In_1288,In_1130);
or U919 (N_919,In_3698,In_4050);
nand U920 (N_920,In_4972,In_2927);
nor U921 (N_921,In_4747,In_3442);
or U922 (N_922,In_3911,In_4153);
or U923 (N_923,In_2855,In_4065);
nor U924 (N_924,N_436,N_285);
xor U925 (N_925,In_0,In_3353);
nand U926 (N_926,In_3969,In_4851);
xor U927 (N_927,In_4839,In_4850);
nor U928 (N_928,In_2301,In_2051);
nand U929 (N_929,In_4273,In_4870);
nand U930 (N_930,In_3803,In_3513);
nand U931 (N_931,In_46,In_1535);
nor U932 (N_932,In_759,N_118);
nor U933 (N_933,In_1270,In_2457);
xnor U934 (N_934,In_1687,In_922);
nor U935 (N_935,In_4590,N_191);
or U936 (N_936,In_661,In_3756);
or U937 (N_937,In_3203,In_914);
nand U938 (N_938,In_3839,In_3521);
nand U939 (N_939,In_1796,In_2949);
nand U940 (N_940,In_1941,In_4739);
xnor U941 (N_941,In_2952,In_3930);
or U942 (N_942,In_1347,In_4519);
and U943 (N_943,N_94,In_4562);
and U944 (N_944,In_933,In_3872);
nor U945 (N_945,In_4146,In_3120);
nor U946 (N_946,In_238,In_4342);
or U947 (N_947,In_1160,In_4781);
xnor U948 (N_948,In_2656,In_623);
and U949 (N_949,N_164,In_1062);
nand U950 (N_950,In_1918,In_1549);
nand U951 (N_951,In_4573,In_2512);
or U952 (N_952,In_4738,In_1976);
or U953 (N_953,In_2993,In_3266);
xnor U954 (N_954,N_290,In_195);
or U955 (N_955,In_4442,In_4095);
nand U956 (N_956,In_1566,In_985);
nand U957 (N_957,In_4603,N_393);
nand U958 (N_958,In_4779,In_3599);
or U959 (N_959,In_2356,In_775);
or U960 (N_960,In_4235,In_1819);
nor U961 (N_961,In_2049,N_479);
nor U962 (N_962,In_4424,In_4081);
nand U963 (N_963,In_1909,In_4514);
and U964 (N_964,In_1897,In_2648);
and U965 (N_965,In_2089,In_3902);
nor U966 (N_966,In_4349,In_24);
nor U967 (N_967,In_558,N_116);
xnor U968 (N_968,In_4400,In_2652);
or U969 (N_969,In_4186,N_471);
xor U970 (N_970,In_1256,In_2988);
xor U971 (N_971,In_2360,N_401);
nor U972 (N_972,In_1798,In_2452);
nand U973 (N_973,In_4302,In_2693);
or U974 (N_974,In_4123,In_2888);
nand U975 (N_975,In_1840,In_2628);
or U976 (N_976,In_4541,In_2365);
nor U977 (N_977,In_4692,In_2748);
or U978 (N_978,In_4677,In_4962);
nand U979 (N_979,In_603,In_2399);
xor U980 (N_980,In_2944,N_140);
nand U981 (N_981,In_1611,In_4309);
nor U982 (N_982,N_488,In_9);
nor U983 (N_983,In_4314,In_3904);
xor U984 (N_984,In_2653,In_1544);
or U985 (N_985,N_446,N_341);
nand U986 (N_986,In_3986,In_3149);
nand U987 (N_987,In_1805,In_4084);
or U988 (N_988,N_25,In_3552);
nand U989 (N_989,In_1756,In_2681);
or U990 (N_990,In_4072,In_709);
nor U991 (N_991,N_252,In_4881);
and U992 (N_992,In_4413,In_1363);
nor U993 (N_993,In_1708,In_3379);
and U994 (N_994,In_3508,In_3656);
nand U995 (N_995,In_3556,N_284);
xnor U996 (N_996,In_2287,In_839);
nand U997 (N_997,In_3075,In_2276);
and U998 (N_998,In_4886,N_33);
nand U999 (N_999,In_1977,In_2345);
nand U1000 (N_1000,In_2907,N_649);
and U1001 (N_1001,N_715,N_193);
nor U1002 (N_1002,In_4224,In_3518);
or U1003 (N_1003,In_256,In_2235);
and U1004 (N_1004,In_4822,In_4857);
xor U1005 (N_1005,In_3383,In_2678);
xnor U1006 (N_1006,In_177,N_125);
xor U1007 (N_1007,In_3873,N_692);
xor U1008 (N_1008,In_1426,N_8);
xor U1009 (N_1009,In_1369,In_645);
and U1010 (N_1010,In_3563,In_4718);
xor U1011 (N_1011,In_4526,In_4995);
or U1012 (N_1012,In_2145,In_3745);
nor U1013 (N_1013,N_305,In_1342);
or U1014 (N_1014,In_2826,In_1013);
nand U1015 (N_1015,N_927,In_4539);
nand U1016 (N_1016,N_185,In_3246);
nand U1017 (N_1017,In_1838,In_3958);
xnor U1018 (N_1018,In_785,In_2420);
xor U1019 (N_1019,In_4537,In_1556);
nor U1020 (N_1020,N_95,N_824);
nor U1021 (N_1021,In_4484,In_577);
and U1022 (N_1022,N_581,In_2071);
or U1023 (N_1023,In_1097,In_3139);
or U1024 (N_1024,In_4978,N_734);
and U1025 (N_1025,In_4230,In_2722);
xnor U1026 (N_1026,In_4575,In_1086);
nand U1027 (N_1027,In_1500,In_3058);
nor U1028 (N_1028,In_1537,In_3548);
and U1029 (N_1029,In_4308,N_578);
and U1030 (N_1030,In_1874,In_399);
or U1031 (N_1031,In_1159,In_1345);
xnor U1032 (N_1032,In_2003,In_57);
xor U1033 (N_1033,In_1479,N_536);
xnor U1034 (N_1034,N_835,In_1217);
nand U1035 (N_1035,N_293,N_85);
nor U1036 (N_1036,In_2942,N_162);
or U1037 (N_1037,In_2618,In_2167);
nand U1038 (N_1038,N_532,In_4383);
nand U1039 (N_1039,N_861,In_1541);
and U1040 (N_1040,In_4750,In_242);
nor U1041 (N_1041,In_3006,In_3167);
xnor U1042 (N_1042,N_876,In_1578);
and U1043 (N_1043,N_769,In_2207);
and U1044 (N_1044,In_121,In_356);
nand U1045 (N_1045,N_620,In_561);
or U1046 (N_1046,In_3270,In_1754);
nand U1047 (N_1047,In_3032,In_4255);
or U1048 (N_1048,In_2461,In_97);
and U1049 (N_1049,In_4908,N_206);
nand U1050 (N_1050,N_803,N_520);
or U1051 (N_1051,In_856,In_511);
or U1052 (N_1052,N_392,In_1548);
or U1053 (N_1053,In_3338,In_2683);
xor U1054 (N_1054,In_3602,In_2482);
and U1055 (N_1055,In_1877,In_364);
nor U1056 (N_1056,N_188,In_3074);
nand U1057 (N_1057,N_40,In_1832);
nand U1058 (N_1058,In_3923,In_4163);
xor U1059 (N_1059,In_767,In_1621);
or U1060 (N_1060,In_1597,In_1329);
and U1061 (N_1061,N_200,In_4396);
and U1062 (N_1062,In_3779,N_758);
xor U1063 (N_1063,In_171,In_999);
nand U1064 (N_1064,In_3775,In_4482);
and U1065 (N_1065,N_287,N_833);
nor U1066 (N_1066,In_4834,In_2563);
nor U1067 (N_1067,In_3864,In_2247);
nand U1068 (N_1068,In_287,In_924);
nand U1069 (N_1069,In_1955,In_2751);
nor U1070 (N_1070,In_2695,N_353);
nor U1071 (N_1071,N_954,In_1517);
or U1072 (N_1072,In_4175,In_2408);
or U1073 (N_1073,N_134,In_3077);
nor U1074 (N_1074,In_3990,In_2250);
nand U1075 (N_1075,In_929,In_3064);
and U1076 (N_1076,In_3800,In_1484);
nand U1077 (N_1077,In_4819,N_776);
nand U1078 (N_1078,In_4380,N_525);
and U1079 (N_1079,N_449,In_308);
and U1080 (N_1080,In_4576,N_518);
nor U1081 (N_1081,In_236,In_3279);
nand U1082 (N_1082,N_967,N_562);
nor U1083 (N_1083,In_2588,In_847);
or U1084 (N_1084,In_1764,In_2541);
nor U1085 (N_1085,In_3363,In_2665);
nor U1086 (N_1086,N_988,N_883);
and U1087 (N_1087,In_1582,In_2731);
xnor U1088 (N_1088,N_204,In_3620);
nor U1089 (N_1089,In_4684,In_1919);
nor U1090 (N_1090,In_4503,In_4274);
or U1091 (N_1091,In_4310,N_892);
and U1092 (N_1092,In_475,In_4665);
and U1093 (N_1093,In_872,N_730);
and U1094 (N_1094,In_333,In_1274);
nor U1095 (N_1095,In_1786,In_1998);
or U1096 (N_1096,N_782,In_3197);
nor U1097 (N_1097,In_397,In_4835);
and U1098 (N_1098,In_2081,In_4805);
nor U1099 (N_1099,In_3140,In_1939);
nand U1100 (N_1100,N_973,In_1098);
or U1101 (N_1101,In_436,In_569);
nand U1102 (N_1102,N_302,N_13);
and U1103 (N_1103,In_1216,In_1808);
or U1104 (N_1104,In_3206,In_4731);
nor U1105 (N_1105,In_1425,In_3222);
or U1106 (N_1106,In_3757,In_1644);
xor U1107 (N_1107,In_416,In_4878);
or U1108 (N_1108,In_1029,In_2176);
nor U1109 (N_1109,In_572,In_4818);
nand U1110 (N_1110,In_936,In_4801);
nand U1111 (N_1111,In_2536,N_104);
and U1112 (N_1112,N_573,In_3931);
nor U1113 (N_1113,In_409,In_549);
and U1114 (N_1114,In_2747,In_360);
nand U1115 (N_1115,In_201,In_909);
nand U1116 (N_1116,In_1701,In_1837);
and U1117 (N_1117,N_497,In_3741);
or U1118 (N_1118,In_1923,N_653);
or U1119 (N_1119,In_4348,In_387);
xnor U1120 (N_1120,In_600,In_3352);
xor U1121 (N_1121,In_1403,In_4462);
nor U1122 (N_1122,N_477,In_4685);
xor U1123 (N_1123,In_2002,In_1121);
and U1124 (N_1124,In_2382,In_1990);
and U1125 (N_1125,N_567,In_4295);
or U1126 (N_1126,In_2711,In_3373);
nand U1127 (N_1127,N_795,In_3218);
nor U1128 (N_1128,In_2031,In_4206);
nand U1129 (N_1129,In_688,In_4011);
nand U1130 (N_1130,N_798,In_2277);
and U1131 (N_1131,In_2958,In_3977);
nor U1132 (N_1132,N_241,In_4841);
xor U1133 (N_1133,In_877,In_1579);
xor U1134 (N_1134,In_2550,In_4197);
nor U1135 (N_1135,In_4416,In_766);
xor U1136 (N_1136,In_832,In_4094);
xor U1137 (N_1137,In_377,N_339);
xnor U1138 (N_1138,N_872,In_2475);
xnor U1139 (N_1139,In_3964,In_677);
nor U1140 (N_1140,N_491,In_760);
or U1141 (N_1141,In_3401,In_4381);
and U1142 (N_1142,N_219,N_742);
xnor U1143 (N_1143,In_3303,In_3957);
nand U1144 (N_1144,N_931,In_1509);
nand U1145 (N_1145,N_346,In_3524);
nand U1146 (N_1146,In_2904,In_2758);
nand U1147 (N_1147,In_3411,In_3199);
nand U1148 (N_1148,In_4776,In_4783);
nor U1149 (N_1149,In_4659,N_503);
xnor U1150 (N_1150,In_4130,In_3885);
and U1151 (N_1151,In_1475,In_2643);
nand U1152 (N_1152,In_2040,N_688);
and U1153 (N_1153,In_3481,N_368);
nor U1154 (N_1154,In_2019,In_2009);
nand U1155 (N_1155,N_127,In_3562);
and U1156 (N_1156,N_388,In_2878);
nand U1157 (N_1157,In_3224,In_4633);
xnor U1158 (N_1158,In_1282,In_1814);
and U1159 (N_1159,In_4929,In_3326);
or U1160 (N_1160,In_4820,In_1738);
nor U1161 (N_1161,N_534,In_1773);
and U1162 (N_1162,In_3746,In_971);
nor U1163 (N_1163,In_3943,In_3596);
xor U1164 (N_1164,In_818,In_4192);
nand U1165 (N_1165,In_3193,In_618);
nand U1166 (N_1166,In_1932,In_4324);
xnor U1167 (N_1167,In_648,In_3936);
xnor U1168 (N_1168,N_42,In_3420);
nand U1169 (N_1169,N_43,N_155);
xor U1170 (N_1170,In_3748,In_3090);
xnor U1171 (N_1171,In_125,In_2204);
nand U1172 (N_1172,In_2777,N_898);
xnor U1173 (N_1173,In_3415,In_2158);
and U1174 (N_1174,In_3701,N_713);
or U1175 (N_1175,In_1260,In_1237);
and U1176 (N_1176,N_187,In_1188);
or U1177 (N_1177,In_598,In_1889);
nor U1178 (N_1178,N_631,In_1441);
or U1179 (N_1179,In_4351,In_4456);
and U1180 (N_1180,In_1307,In_4296);
and U1181 (N_1181,In_1931,In_517);
xnor U1182 (N_1182,N_466,In_4786);
xor U1183 (N_1183,In_4772,In_3778);
xnor U1184 (N_1184,N_270,In_2466);
and U1185 (N_1185,N_156,In_232);
nand U1186 (N_1186,In_1647,In_4402);
nand U1187 (N_1187,In_4667,In_2597);
and U1188 (N_1188,N_660,In_4831);
nand U1189 (N_1189,In_1829,In_737);
nor U1190 (N_1190,In_4165,In_1271);
nand U1191 (N_1191,In_2718,In_1318);
nor U1192 (N_1192,In_2602,N_367);
or U1193 (N_1193,In_3287,In_327);
and U1194 (N_1194,In_2575,In_2632);
or U1195 (N_1195,In_3459,In_4443);
nor U1196 (N_1196,In_749,In_4118);
or U1197 (N_1197,In_4200,N_113);
nor U1198 (N_1198,In_2840,In_474);
xnor U1199 (N_1199,In_2972,In_4290);
nand U1200 (N_1200,In_4625,In_4214);
nand U1201 (N_1201,In_4216,In_3005);
nand U1202 (N_1202,In_757,In_4966);
nand U1203 (N_1203,N_757,In_426);
or U1204 (N_1204,In_2997,In_2848);
and U1205 (N_1205,In_2614,In_3053);
or U1206 (N_1206,In_4111,In_2682);
xnor U1207 (N_1207,In_4672,In_1862);
and U1208 (N_1208,In_374,In_1389);
nor U1209 (N_1209,N_325,N_987);
or U1210 (N_1210,In_1238,In_2298);
nand U1211 (N_1211,In_2057,In_4930);
or U1212 (N_1212,In_1250,In_3185);
nor U1213 (N_1213,In_3700,In_2780);
nor U1214 (N_1214,In_4970,In_4862);
nand U1215 (N_1215,N_907,N_781);
xor U1216 (N_1216,In_1057,In_1377);
and U1217 (N_1217,In_1290,In_3716);
nor U1218 (N_1218,In_4939,In_4412);
nor U1219 (N_1219,N_739,In_3044);
or U1220 (N_1220,In_1467,In_1924);
xnor U1221 (N_1221,In_4131,N_224);
nor U1222 (N_1222,In_1478,N_79);
xor U1223 (N_1223,In_148,N_568);
and U1224 (N_1224,In_743,In_2054);
xnor U1225 (N_1225,N_383,In_952);
or U1226 (N_1226,In_1357,In_3496);
nand U1227 (N_1227,In_259,N_546);
or U1228 (N_1228,N_825,In_1392);
and U1229 (N_1229,In_851,In_4554);
nor U1230 (N_1230,In_4057,N_827);
or U1231 (N_1231,N_674,In_1114);
and U1232 (N_1232,In_812,In_4243);
and U1233 (N_1233,In_977,In_4284);
nand U1234 (N_1234,In_1641,In_4885);
nand U1235 (N_1235,In_750,N_274);
nand U1236 (N_1236,N_828,In_207);
nand U1237 (N_1237,In_2562,In_2520);
xor U1238 (N_1238,In_1815,In_1433);
nor U1239 (N_1239,In_1682,In_56);
nor U1240 (N_1240,In_1571,In_4919);
or U1241 (N_1241,In_3846,In_729);
or U1242 (N_1242,In_813,In_665);
nand U1243 (N_1243,In_4293,N_259);
nor U1244 (N_1244,In_3029,In_1699);
nor U1245 (N_1245,In_4464,In_1606);
nor U1246 (N_1246,In_1637,N_494);
and U1247 (N_1247,In_105,In_4097);
nand U1248 (N_1248,N_530,N_921);
nor U1249 (N_1249,In_2100,In_3650);
and U1250 (N_1250,In_4950,N_558);
xor U1251 (N_1251,In_692,In_2879);
or U1252 (N_1252,In_3201,In_3782);
nand U1253 (N_1253,In_3473,In_3949);
or U1254 (N_1254,In_3059,In_3614);
and U1255 (N_1255,In_2128,In_2026);
nor U1256 (N_1256,In_65,N_315);
nor U1257 (N_1257,In_2087,In_3529);
nand U1258 (N_1258,N_802,In_3801);
and U1259 (N_1259,In_1042,In_2281);
nor U1260 (N_1260,N_86,In_2999);
and U1261 (N_1261,In_4179,In_4758);
xor U1262 (N_1262,In_1253,In_2824);
xnor U1263 (N_1263,N_153,In_781);
or U1264 (N_1264,In_4061,In_1595);
nor U1265 (N_1265,In_2662,In_1703);
or U1266 (N_1266,N_110,N_192);
nand U1267 (N_1267,In_968,In_6);
nand U1268 (N_1268,In_2416,In_210);
nor U1269 (N_1269,In_494,In_4848);
and U1270 (N_1270,In_4588,In_214);
nand U1271 (N_1271,In_1333,N_559);
nand U1272 (N_1272,In_2154,N_109);
or U1273 (N_1273,N_787,In_4967);
nor U1274 (N_1274,In_3877,In_2768);
nor U1275 (N_1275,N_76,In_4948);
xor U1276 (N_1276,In_3156,In_2592);
and U1277 (N_1277,In_1625,In_4615);
nor U1278 (N_1278,N_460,In_429);
nand U1279 (N_1279,In_2869,In_1608);
nor U1280 (N_1280,In_4110,N_976);
and U1281 (N_1281,In_446,N_31);
xnor U1282 (N_1282,In_4246,N_762);
or U1283 (N_1283,N_10,In_733);
xor U1284 (N_1284,In_3119,In_584);
xnor U1285 (N_1285,In_987,In_1455);
xnor U1286 (N_1286,N_866,N_571);
xor U1287 (N_1287,N_612,In_4709);
nor U1288 (N_1288,N_785,In_939);
nor U1289 (N_1289,In_1847,In_696);
nor U1290 (N_1290,In_3054,In_217);
or U1291 (N_1291,In_3361,N_16);
nor U1292 (N_1292,In_1315,N_505);
nor U1293 (N_1293,N_380,N_799);
or U1294 (N_1294,In_1332,In_858);
and U1295 (N_1295,In_4435,In_2369);
nor U1296 (N_1296,In_3713,N_815);
and U1297 (N_1297,In_3066,In_27);
nor U1298 (N_1298,In_3290,In_4100);
nor U1299 (N_1299,In_3096,N_980);
nor U1300 (N_1300,N_400,In_1551);
nor U1301 (N_1301,In_2041,N_459);
nand U1302 (N_1302,In_582,In_4565);
or U1303 (N_1303,N_512,In_463);
nand U1304 (N_1304,In_1884,In_4102);
and U1305 (N_1305,In_330,In_1907);
xnor U1306 (N_1306,N_237,N_557);
xor U1307 (N_1307,In_1006,In_973);
or U1308 (N_1308,In_12,In_5);
or U1309 (N_1309,In_1483,In_1204);
or U1310 (N_1310,In_3370,In_3112);
nor U1311 (N_1311,In_663,In_1285);
nor U1312 (N_1312,N_502,N_129);
and U1313 (N_1313,In_4231,N_122);
xor U1314 (N_1314,In_4388,N_510);
and U1315 (N_1315,In_4879,In_4312);
or U1316 (N_1316,In_979,In_4142);
or U1317 (N_1317,In_84,In_178);
or U1318 (N_1318,In_637,In_4190);
nand U1319 (N_1319,In_3929,In_624);
nand U1320 (N_1320,N_634,In_3309);
or U1321 (N_1321,In_932,In_4622);
xnor U1322 (N_1322,In_32,In_4394);
xor U1323 (N_1323,In_2269,In_2481);
and U1324 (N_1324,In_2616,In_2367);
nor U1325 (N_1325,In_1904,In_3675);
or U1326 (N_1326,In_1935,In_3790);
nand U1327 (N_1327,In_998,In_4695);
nor U1328 (N_1328,In_739,N_569);
xnor U1329 (N_1329,In_398,In_3868);
xor U1330 (N_1330,In_689,In_2091);
xnor U1331 (N_1331,In_4796,In_4894);
xnor U1332 (N_1332,In_1813,In_4943);
nor U1333 (N_1333,In_1263,In_2036);
or U1334 (N_1334,N_190,In_2146);
and U1335 (N_1335,In_211,N_21);
nand U1336 (N_1336,In_4430,In_2006);
xor U1337 (N_1337,In_4001,In_2947);
xor U1338 (N_1338,In_3639,In_2570);
or U1339 (N_1339,In_3648,In_4493);
or U1340 (N_1340,In_2566,In_1324);
nor U1341 (N_1341,In_497,N_720);
xor U1342 (N_1342,In_129,In_4947);
or U1343 (N_1343,In_1790,In_2453);
nand U1344 (N_1344,In_3681,In_1831);
nor U1345 (N_1345,In_3866,N_207);
xnor U1346 (N_1346,In_1795,In_4628);
and U1347 (N_1347,In_2918,In_2465);
nand U1348 (N_1348,In_4511,In_2581);
and U1349 (N_1349,N_0,In_3079);
nand U1350 (N_1350,In_1883,In_192);
or U1351 (N_1351,In_3875,In_1564);
or U1352 (N_1352,In_1676,In_988);
or U1353 (N_1353,N_695,In_2251);
or U1354 (N_1354,In_1273,In_535);
nor U1355 (N_1355,N_627,In_3490);
nand U1356 (N_1356,In_4397,In_4082);
or U1357 (N_1357,In_3841,In_465);
nand U1358 (N_1358,In_1053,In_2901);
or U1359 (N_1359,In_3311,In_566);
nand U1360 (N_1360,N_233,In_625);
nor U1361 (N_1361,In_680,In_2615);
nand U1362 (N_1362,N_675,N_407);
nand U1363 (N_1363,In_2905,In_595);
and U1364 (N_1364,In_320,N_788);
or U1365 (N_1365,N_899,N_12);
and U1366 (N_1366,N_248,In_1863);
and U1367 (N_1367,In_3391,N_968);
or U1368 (N_1368,N_60,N_133);
nand U1369 (N_1369,In_2055,In_528);
or U1370 (N_1370,In_393,In_1742);
or U1371 (N_1371,In_4792,N_994);
nand U1372 (N_1372,In_2409,In_3350);
nor U1373 (N_1373,In_1144,In_3621);
xor U1374 (N_1374,In_294,In_2725);
and U1375 (N_1375,N_329,In_3465);
or U1376 (N_1376,In_2690,In_1964);
nor U1377 (N_1377,In_4070,In_4864);
nor U1378 (N_1378,In_3974,In_2094);
xor U1379 (N_1379,N_470,In_3135);
nor U1380 (N_1380,In_904,In_1396);
nor U1381 (N_1381,N_576,In_4450);
and U1382 (N_1382,In_1454,In_1087);
xor U1383 (N_1383,In_4965,In_2001);
nand U1384 (N_1384,In_910,In_2583);
and U1385 (N_1385,In_2086,In_3323);
nand U1386 (N_1386,In_507,N_359);
xnor U1387 (N_1387,In_1401,In_4813);
nand U1388 (N_1388,In_1037,In_2242);
and U1389 (N_1389,In_1570,In_2464);
xor U1390 (N_1390,In_485,In_2043);
or U1391 (N_1391,In_4827,N_705);
nand U1392 (N_1392,N_639,N_513);
nand U1393 (N_1393,N_990,In_1881);
or U1394 (N_1394,N_778,In_4704);
nand U1395 (N_1395,In_792,N_657);
xnor U1396 (N_1396,N_652,In_471);
xnor U1397 (N_1397,In_989,In_3627);
nand U1398 (N_1398,In_819,N_69);
xnor U1399 (N_1399,In_3239,In_945);
and U1400 (N_1400,In_4171,In_226);
nor U1401 (N_1401,In_3487,In_870);
or U1402 (N_1402,In_1302,In_628);
nor U1403 (N_1403,N_186,In_1323);
or U1404 (N_1404,In_3593,In_2219);
or U1405 (N_1405,In_980,In_2625);
or U1406 (N_1406,In_3209,In_1393);
and U1407 (N_1407,In_149,In_2672);
xnor U1408 (N_1408,In_2666,In_1961);
or U1409 (N_1409,In_3028,In_2447);
or U1410 (N_1410,In_3226,In_427);
and U1411 (N_1411,In_3060,In_3783);
nand U1412 (N_1412,In_3610,In_3661);
or U1413 (N_1413,In_2107,In_2980);
xor U1414 (N_1414,In_1404,In_2378);
nand U1415 (N_1415,In_3486,In_2849);
or U1416 (N_1416,N_738,N_521);
nand U1417 (N_1417,In_132,In_3768);
and U1418 (N_1418,In_4961,In_2209);
xor U1419 (N_1419,N_670,N_759);
nand U1420 (N_1420,In_4924,In_2065);
xor U1421 (N_1421,In_3400,In_3475);
or U1422 (N_1422,In_4139,In_19);
nor U1423 (N_1423,In_678,In_3836);
nor U1424 (N_1424,In_3519,In_1744);
or U1425 (N_1425,In_3057,In_2720);
xor U1426 (N_1426,N_131,N_535);
and U1427 (N_1427,In_3116,In_1135);
and U1428 (N_1428,In_4595,In_1702);
or U1429 (N_1429,In_3145,In_2489);
or U1430 (N_1430,In_1946,N_707);
nand U1431 (N_1431,In_4749,N_996);
or U1432 (N_1432,N_137,N_819);
xnor U1433 (N_1433,In_567,In_1292);
xnor U1434 (N_1434,In_4617,In_3501);
nand U1435 (N_1435,In_1043,In_4159);
nor U1436 (N_1436,In_4877,In_1096);
nor U1437 (N_1437,In_4780,N_914);
nand U1438 (N_1438,In_34,In_524);
nand U1439 (N_1439,In_277,N_682);
and U1440 (N_1440,In_1993,N_381);
and U1441 (N_1441,In_4022,N_724);
and U1442 (N_1442,In_4507,N_362);
nor U1443 (N_1443,In_1848,N_937);
and U1444 (N_1444,In_4458,In_1942);
xnor U1445 (N_1445,In_4679,In_2867);
or U1446 (N_1446,In_4896,In_3430);
xor U1447 (N_1447,N_854,N_526);
xor U1448 (N_1448,In_4884,In_2467);
nor U1449 (N_1449,In_2101,N_375);
or U1450 (N_1450,In_3376,In_554);
and U1451 (N_1451,In_2402,In_4486);
and U1452 (N_1452,In_3292,N_948);
or U1453 (N_1453,In_3649,N_845);
nor U1454 (N_1454,In_4979,In_1139);
nor U1455 (N_1455,In_2812,In_2286);
and U1456 (N_1456,In_2577,In_919);
and U1457 (N_1457,N_697,In_2342);
and U1458 (N_1458,N_596,N_638);
nand U1459 (N_1459,In_2772,In_1269);
and U1460 (N_1460,N_38,In_3737);
xnor U1461 (N_1461,In_67,In_4106);
nand U1462 (N_1462,In_2423,In_1173);
nand U1463 (N_1463,N_264,N_884);
nand U1464 (N_1464,In_3024,N_791);
or U1465 (N_1465,In_2455,In_2050);
or U1466 (N_1466,In_36,N_851);
and U1467 (N_1467,N_458,In_4544);
and U1468 (N_1468,In_2354,In_2729);
or U1469 (N_1469,In_2835,In_2304);
nand U1470 (N_1470,In_1959,N_46);
xor U1471 (N_1471,In_3155,In_4807);
xor U1472 (N_1472,In_2039,In_2712);
or U1473 (N_1473,In_298,In_4266);
xnor U1474 (N_1474,N_696,In_4523);
nand U1475 (N_1475,In_3048,In_3697);
xor U1476 (N_1476,In_2540,In_1811);
nand U1477 (N_1477,In_4901,In_4116);
and U1478 (N_1478,In_3677,In_4270);
and U1479 (N_1479,In_921,In_4234);
nand U1480 (N_1480,In_983,In_515);
or U1481 (N_1481,N_149,N_810);
nand U1482 (N_1482,In_1622,In_2967);
nand U1483 (N_1483,N_746,N_677);
nand U1484 (N_1484,In_1447,In_718);
nand U1485 (N_1485,N_555,In_3055);
or U1486 (N_1486,N_56,In_3298);
xnor U1487 (N_1487,N_425,In_4346);
nor U1488 (N_1488,In_1492,N_600);
xnor U1489 (N_1489,In_4060,In_339);
nor U1490 (N_1490,In_865,In_2584);
and U1491 (N_1491,In_2494,N_553);
xnor U1492 (N_1492,In_3397,N_36);
nand U1493 (N_1493,In_144,N_906);
and U1494 (N_1494,N_993,N_814);
nor U1495 (N_1495,In_2121,In_2991);
nand U1496 (N_1496,In_2932,In_3618);
or U1497 (N_1497,In_2476,In_2946);
nor U1498 (N_1498,N_7,In_3364);
nand U1499 (N_1499,In_3688,In_2908);
and U1500 (N_1500,In_3597,In_1158);
xnor U1501 (N_1501,In_2436,N_1246);
xnor U1502 (N_1502,In_4991,In_1468);
nor U1503 (N_1503,In_1126,In_4193);
nor U1504 (N_1504,N_1133,In_1405);
and U1505 (N_1505,In_1128,In_3443);
or U1506 (N_1506,In_2845,In_4645);
and U1507 (N_1507,In_351,In_1022);
nor U1508 (N_1508,In_3708,In_3445);
nor U1509 (N_1509,In_720,In_4631);
and U1510 (N_1510,N_1330,N_1098);
nor U1511 (N_1511,In_1448,In_1352);
nand U1512 (N_1512,In_2619,In_3211);
or U1513 (N_1513,In_510,N_1020);
nor U1514 (N_1514,In_4223,In_78);
xor U1515 (N_1515,In_1381,In_3849);
and U1516 (N_1516,In_1519,In_1219);
nor U1517 (N_1517,In_842,N_862);
nand U1518 (N_1518,N_889,N_942);
nor U1519 (N_1519,In_4320,In_2156);
nand U1520 (N_1520,In_1812,In_913);
or U1521 (N_1521,N_941,In_2289);
and U1522 (N_1522,N_2,N_905);
xor U1523 (N_1523,N_1427,N_194);
nor U1524 (N_1524,In_2048,In_2858);
xnor U1525 (N_1525,N_587,In_4990);
nor U1526 (N_1526,In_1473,N_415);
or U1527 (N_1527,In_4953,In_946);
nand U1528 (N_1528,In_3416,In_1951);
or U1529 (N_1529,In_1588,In_3474);
and U1530 (N_1530,In_704,N_318);
nand U1531 (N_1531,N_146,N_998);
and U1532 (N_1532,In_3186,In_4401);
and U1533 (N_1533,N_496,N_1001);
and U1534 (N_1534,In_4080,In_4150);
xnor U1535 (N_1535,In_2525,N_176);
nand U1536 (N_1536,N_965,In_4465);
or U1537 (N_1537,In_685,In_1659);
and U1538 (N_1538,In_206,N_1352);
or U1539 (N_1539,In_3601,In_4183);
or U1540 (N_1540,N_611,N_384);
xnor U1541 (N_1541,In_4712,In_3166);
or U1542 (N_1542,In_644,In_698);
or U1543 (N_1543,N_763,In_2911);
nand U1544 (N_1544,N_676,N_626);
or U1545 (N_1545,In_4417,In_2337);
or U1546 (N_1546,N_641,In_80);
and U1547 (N_1547,N_135,In_4678);
xor U1548 (N_1548,N_882,In_2097);
nor U1549 (N_1549,In_752,In_2222);
nand U1550 (N_1550,In_4262,In_1609);
and U1551 (N_1551,In_803,In_3313);
or U1552 (N_1552,In_4358,In_2971);
nand U1553 (N_1553,In_2811,In_2027);
xor U1554 (N_1554,N_1419,N_891);
nand U1555 (N_1555,In_2275,N_565);
xor U1556 (N_1556,In_915,In_1762);
and U1557 (N_1557,In_3375,In_1670);
and U1558 (N_1558,In_4566,In_4063);
or U1559 (N_1559,In_4344,In_1397);
nor U1560 (N_1560,In_1584,N_750);
and U1561 (N_1561,In_1272,In_822);
nor U1562 (N_1562,In_3843,In_306);
or U1563 (N_1563,In_3056,In_1457);
nand U1564 (N_1564,In_4895,In_4898);
nand U1565 (N_1565,N_673,In_3542);
or U1566 (N_1566,In_4425,In_2862);
nand U1567 (N_1567,In_229,N_1088);
or U1568 (N_1568,In_547,In_3676);
nor U1569 (N_1569,In_650,In_3020);
or U1570 (N_1570,In_2719,In_176);
nand U1571 (N_1571,In_1824,In_4563);
and U1572 (N_1572,N_1402,N_575);
and U1573 (N_1573,In_3512,In_837);
nand U1574 (N_1574,In_4079,In_1915);
nand U1575 (N_1575,N_794,In_3577);
or U1576 (N_1576,In_894,In_2413);
and U1577 (N_1577,N_989,In_654);
or U1578 (N_1578,N_838,In_874);
or U1579 (N_1579,N_1117,N_454);
or U1580 (N_1580,In_4746,In_2685);
and U1581 (N_1581,N_860,In_1301);
or U1582 (N_1582,In_2919,In_1390);
and U1583 (N_1583,N_689,N_1432);
nor U1584 (N_1584,In_2400,In_2851);
or U1585 (N_1585,In_438,N_473);
or U1586 (N_1586,In_782,In_3372);
xnor U1587 (N_1587,In_1666,N_171);
xor U1588 (N_1588,N_197,In_2511);
xor U1589 (N_1589,N_178,In_4596);
nor U1590 (N_1590,In_579,In_2925);
nor U1591 (N_1591,N_1264,In_1365);
nor U1592 (N_1592,N_647,In_3097);
or U1593 (N_1593,In_2462,In_3538);
nor U1594 (N_1594,In_4042,In_3357);
or U1595 (N_1595,N_1200,In_2825);
nand U1596 (N_1596,In_4297,In_4247);
nor U1597 (N_1597,In_519,In_231);
or U1598 (N_1598,In_4648,N_962);
xor U1599 (N_1599,In_2799,In_3083);
nand U1600 (N_1600,In_459,N_509);
xnor U1601 (N_1601,In_2644,In_960);
xor U1602 (N_1602,In_673,In_4741);
or U1603 (N_1603,N_1313,In_1257);
nor U1604 (N_1604,In_4420,N_1182);
and U1605 (N_1605,In_1223,In_3428);
nand U1606 (N_1606,In_2708,N_430);
or U1607 (N_1607,N_212,N_395);
and U1608 (N_1608,In_863,In_235);
or U1609 (N_1609,In_169,N_91);
nand U1610 (N_1610,In_3160,N_665);
nor U1611 (N_1611,In_268,In_1685);
and U1612 (N_1612,In_3764,In_1540);
nand U1613 (N_1613,In_961,In_867);
or U1614 (N_1614,In_1842,N_1170);
xor U1615 (N_1615,In_158,In_1001);
nand U1616 (N_1616,N_205,N_527);
or U1617 (N_1617,N_253,In_1236);
or U1618 (N_1618,In_4093,In_2646);
and U1619 (N_1619,N_982,In_109);
or U1620 (N_1620,In_541,N_1120);
and U1621 (N_1621,In_1461,N_726);
nand U1622 (N_1622,N_945,N_1066);
nor U1623 (N_1623,In_2142,In_769);
and U1624 (N_1624,N_98,N_108);
nand U1625 (N_1625,In_2578,In_1199);
nor U1626 (N_1626,In_1129,In_1206);
or U1627 (N_1627,N_554,In_200);
or U1628 (N_1628,N_429,In_1344);
or U1629 (N_1629,In_3348,In_4585);
nor U1630 (N_1630,N_196,N_266);
and U1631 (N_1631,N_1413,In_3724);
and U1632 (N_1632,In_708,N_628);
nor U1633 (N_1633,In_4052,In_928);
and U1634 (N_1634,In_4843,In_2734);
xnor U1635 (N_1635,In_4374,N_210);
and U1636 (N_1636,N_1174,In_1779);
and U1637 (N_1637,In_161,In_3329);
or U1638 (N_1638,In_4449,In_4421);
or U1639 (N_1639,In_539,In_3886);
xnor U1640 (N_1640,In_371,In_4666);
and U1641 (N_1641,N_842,In_414);
xor U1642 (N_1642,N_365,N_103);
or U1643 (N_1643,N_541,N_917);
nor U1644 (N_1644,In_2900,In_1309);
and U1645 (N_1645,In_2774,N_121);
xor U1646 (N_1646,In_1002,In_2634);
nor U1647 (N_1647,In_2759,N_280);
xor U1648 (N_1648,N_594,In_4798);
and U1649 (N_1649,N_1282,In_1091);
and U1650 (N_1650,In_2372,In_2636);
and U1651 (N_1651,N_265,In_1021);
and U1652 (N_1652,In_2800,N_956);
xor U1653 (N_1653,In_4946,N_900);
or U1654 (N_1654,N_1058,N_894);
nand U1655 (N_1655,In_869,In_1733);
and U1656 (N_1656,In_4041,N_1480);
xor U1657 (N_1657,In_262,In_4715);
and U1658 (N_1658,N_1354,N_1263);
or U1659 (N_1659,In_879,N_1141);
nor U1660 (N_1660,In_4556,N_297);
xor U1661 (N_1661,In_1262,N_1081);
or U1662 (N_1662,N_1321,In_2542);
or U1663 (N_1663,In_4706,In_4698);
and U1664 (N_1664,N_1028,N_1010);
and U1665 (N_1665,N_786,In_2315);
and U1666 (N_1666,N_714,In_343);
xnor U1667 (N_1667,In_903,In_4696);
xnor U1668 (N_1668,In_1192,In_4735);
xnor U1669 (N_1669,In_4912,N_1166);
or U1670 (N_1670,N_1342,In_1419);
and U1671 (N_1671,In_899,In_1543);
or U1672 (N_1672,In_2343,N_659);
nor U1673 (N_1673,In_701,In_1025);
or U1674 (N_1674,N_1431,In_114);
nor U1675 (N_1675,In_3482,In_975);
nor U1676 (N_1676,In_3973,N_1059);
nor U1677 (N_1677,In_635,N_5);
nor U1678 (N_1678,In_2960,In_2519);
nor U1679 (N_1679,N_154,In_2016);
or U1680 (N_1680,N_1255,In_2004);
xor U1681 (N_1681,In_3367,In_1147);
or U1682 (N_1682,In_1728,In_4770);
xnor U1683 (N_1683,In_4428,In_4073);
nor U1684 (N_1684,In_3660,N_128);
xnor U1685 (N_1685,N_1159,In_1875);
and U1686 (N_1686,In_2694,N_544);
and U1687 (N_1687,N_963,In_882);
nor U1688 (N_1688,In_1880,In_1095);
nor U1689 (N_1689,In_2866,N_1488);
nor U1690 (N_1690,In_4291,In_1766);
nand U1691 (N_1691,In_4838,N_1485);
xor U1692 (N_1692,In_2484,N_855);
nand U1693 (N_1693,N_548,In_1296);
xnor U1694 (N_1694,N_1325,In_2733);
nand U1695 (N_1695,N_935,In_508);
xor U1696 (N_1696,N_944,In_4078);
nor U1697 (N_1697,In_1244,In_4498);
nand U1698 (N_1698,In_1316,N_439);
and U1699 (N_1699,In_3515,In_4553);
xnor U1700 (N_1700,In_159,In_3284);
nor U1701 (N_1701,N_1498,In_2995);
xor U1702 (N_1702,In_880,In_691);
or U1703 (N_1703,In_2099,In_745);
nand U1704 (N_1704,In_4829,In_742);
nor U1705 (N_1705,In_651,In_3467);
nand U1706 (N_1706,N_1324,N_1481);
or U1707 (N_1707,In_1008,In_193);
and U1708 (N_1708,In_664,N_865);
nor U1709 (N_1709,In_790,In_3581);
and U1710 (N_1710,N_1031,N_1228);
nor U1711 (N_1711,In_2676,In_26);
nor U1712 (N_1712,N_773,In_4856);
or U1713 (N_1713,N_625,In_1070);
or U1714 (N_1714,N_610,In_693);
and U1715 (N_1715,In_3285,In_2651);
nor U1716 (N_1716,In_476,In_4028);
or U1717 (N_1717,In_493,In_2836);
xnor U1718 (N_1718,In_2966,N_1172);
nor U1719 (N_1719,In_4548,N_1111);
nor U1720 (N_1720,N_1099,N_875);
or U1721 (N_1721,In_3016,N_1415);
and U1722 (N_1722,In_3234,N_609);
or U1723 (N_1723,In_4248,N_580);
and U1724 (N_1724,In_2655,N_1288);
or U1725 (N_1725,In_2046,N_1305);
nor U1726 (N_1726,In_3337,In_3999);
xnor U1727 (N_1727,In_3750,In_3587);
or U1728 (N_1728,In_836,In_2451);
xnor U1729 (N_1729,In_1170,In_1513);
nor U1730 (N_1730,N_584,In_2969);
nand U1731 (N_1731,In_3612,In_388);
xnor U1732 (N_1732,N_6,N_99);
and U1733 (N_1733,N_1425,In_2870);
xnor U1734 (N_1734,In_3314,In_3652);
xnor U1735 (N_1735,N_1048,In_4998);
and U1736 (N_1736,In_3771,In_2244);
or U1737 (N_1737,In_3667,N_1251);
and U1738 (N_1738,N_167,In_4032);
xor U1739 (N_1739,In_1879,In_1090);
and U1740 (N_1740,In_2159,N_744);
and U1741 (N_1741,N_1138,In_4610);
nor U1742 (N_1742,N_722,In_854);
nand U1743 (N_1743,In_3791,In_1132);
xor U1744 (N_1744,In_2109,In_1843);
xor U1745 (N_1745,N_1337,In_3103);
and U1746 (N_1746,N_1094,N_1323);
xor U1747 (N_1747,In_3162,In_520);
or U1748 (N_1748,N_1140,In_3972);
nand U1749 (N_1749,N_234,In_1499);
nor U1750 (N_1750,In_3085,In_3553);
xor U1751 (N_1751,N_1336,N_1343);
or U1752 (N_1752,N_686,In_372);
xnor U1753 (N_1753,In_2635,In_4188);
nand U1754 (N_1754,In_4859,In_1320);
and U1755 (N_1755,In_2545,In_1992);
and U1756 (N_1756,In_2374,In_1679);
and U1757 (N_1757,In_4534,N_1);
xor U1758 (N_1758,N_483,In_2268);
nor U1759 (N_1759,In_3689,N_373);
and U1760 (N_1760,In_4641,In_3208);
nand U1761 (N_1761,In_3360,In_917);
and U1762 (N_1762,In_4377,N_933);
and U1763 (N_1763,N_298,In_4294);
xor U1764 (N_1764,N_410,In_2200);
xnor U1765 (N_1765,In_335,In_2127);
xor U1766 (N_1766,In_4771,N_1450);
or U1767 (N_1767,In_3900,In_593);
xor U1768 (N_1768,N_1089,In_225);
nand U1769 (N_1769,In_2518,N_396);
xor U1770 (N_1770,N_524,In_2832);
or U1771 (N_1771,In_3464,In_4530);
and U1772 (N_1772,In_2131,In_2887);
nand U1773 (N_1773,In_4034,In_1299);
nand U1774 (N_1774,N_1334,In_4250);
nor U1775 (N_1775,In_4963,N_804);
nor U1776 (N_1776,In_1851,N_874);
or U1777 (N_1777,In_154,N_1420);
or U1778 (N_1778,In_1827,N_597);
or U1779 (N_1779,In_4446,In_313);
nand U1780 (N_1780,In_3505,In_136);
and U1781 (N_1781,In_2226,In_2386);
xor U1782 (N_1782,In_122,In_2856);
or U1783 (N_1783,In_3047,In_2622);
and U1784 (N_1784,N_1077,N_1389);
nand U1785 (N_1785,In_3723,In_565);
nand U1786 (N_1786,N_45,In_1740);
or U1787 (N_1787,N_923,N_1491);
and U1788 (N_1788,In_3200,In_2224);
and U1789 (N_1789,In_4513,In_3477);
xor U1790 (N_1790,N_511,In_531);
xnor U1791 (N_1791,In_2964,N_543);
xor U1792 (N_1792,In_2373,In_2894);
nor U1793 (N_1793,N_857,In_886);
or U1794 (N_1794,N_1212,N_1142);
nand U1795 (N_1795,In_1947,In_1767);
and U1796 (N_1796,In_4389,N_770);
and U1797 (N_1797,In_3122,In_2293);
xnor U1798 (N_1798,N_1436,In_4408);
or U1799 (N_1799,N_143,N_1079);
or U1800 (N_1800,In_305,N_593);
xor U1801 (N_1801,N_537,In_809);
xor U1802 (N_1802,In_2621,N_480);
nor U1803 (N_1803,In_2197,In_340);
and U1804 (N_1804,In_385,In_1162);
nor U1805 (N_1805,In_4693,In_3191);
or U1806 (N_1806,N_161,In_2060);
or U1807 (N_1807,In_4410,In_4889);
nand U1808 (N_1808,N_247,N_447);
xnor U1809 (N_1809,N_228,In_3089);
nand U1810 (N_1810,In_2229,In_4897);
and U1811 (N_1811,N_372,N_1092);
nor U1812 (N_1812,N_661,N_55);
or U1813 (N_1813,N_1146,In_2351);
or U1814 (N_1814,In_2169,N_403);
and U1815 (N_1815,In_2807,In_155);
and U1816 (N_1816,N_901,In_4269);
xnor U1817 (N_1817,In_1558,N_1414);
and U1818 (N_1818,In_1010,In_2174);
nor U1819 (N_1819,N_438,In_3805);
nand U1820 (N_1820,In_855,In_163);
xnor U1821 (N_1821,In_2059,In_1930);
and U1822 (N_1822,In_93,N_841);
nor U1823 (N_1823,In_695,N_1440);
xor U1824 (N_1824,In_2654,In_352);
nand U1825 (N_1825,In_4880,In_1321);
and U1826 (N_1826,In_833,In_3272);
xor U1827 (N_1827,In_574,In_1525);
and U1828 (N_1828,In_1774,N_1000);
and U1829 (N_1829,In_2936,In_4957);
nand U1830 (N_1830,In_1859,N_687);
nor U1831 (N_1831,In_3080,N_809);
or U1832 (N_1832,In_1655,In_2177);
nand U1833 (N_1833,N_528,In_3651);
or U1834 (N_1834,In_168,N_1297);
nand U1835 (N_1835,N_806,In_4053);
and U1836 (N_1836,N_856,In_2316);
and U1837 (N_1837,In_2005,In_43);
and U1838 (N_1838,N_117,In_2813);
or U1839 (N_1839,In_1195,In_4687);
xor U1840 (N_1840,In_1465,In_4155);
nand U1841 (N_1841,N_893,N_1071);
or U1842 (N_1842,In_2020,N_919);
nor U1843 (N_1843,N_198,In_1868);
xnor U1844 (N_1844,In_1391,N_1009);
xor U1845 (N_1845,In_1591,In_3371);
xor U1846 (N_1846,In_2609,In_3321);
nand U1847 (N_1847,In_2834,In_4141);
and U1848 (N_1848,In_4489,In_3001);
and U1849 (N_1849,N_737,In_2288);
nand U1850 (N_1850,N_668,In_4160);
xnor U1851 (N_1851,In_1799,In_4151);
and U1852 (N_1852,In_2485,In_4810);
nand U1853 (N_1853,In_1716,N_643);
nor U1854 (N_1854,In_1462,N_371);
xor U1855 (N_1855,N_422,In_4271);
nor U1856 (N_1856,In_3996,N_1421);
nor U1857 (N_1857,N_1219,In_3220);
nor U1858 (N_1858,N_335,N_820);
xor U1859 (N_1859,In_2620,In_1731);
nor U1860 (N_1860,In_754,In_4940);
xor U1861 (N_1861,In_2735,In_2530);
nand U1862 (N_1862,N_455,In_134);
nand U1863 (N_1863,N_1497,In_2933);
or U1864 (N_1864,In_3901,N_971);
or U1865 (N_1865,In_4476,In_3942);
or U1866 (N_1866,In_1496,In_3718);
nand U1867 (N_1867,In_344,In_4510);
or U1868 (N_1868,In_653,In_4350);
nand U1869 (N_1869,N_723,N_1201);
xnor U1870 (N_1870,N_1441,In_3946);
xnor U1871 (N_1871,In_3347,In_3624);
and U1872 (N_1872,In_2715,In_3441);
or U1873 (N_1873,In_1704,In_1026);
nand U1874 (N_1874,N_864,N_598);
and U1875 (N_1875,N_896,N_1476);
and U1876 (N_1876,In_1921,N_760);
and U1877 (N_1877,N_736,In_203);
xor U1878 (N_1878,N_1315,N_107);
or U1879 (N_1879,In_3412,In_1899);
or U1880 (N_1880,N_319,In_2976);
nor U1881 (N_1881,In_1743,N_1284);
and U1882 (N_1882,N_1404,N_732);
nand U1883 (N_1883,In_1408,In_4811);
xor U1884 (N_1884,In_4257,N_717);
nand U1885 (N_1885,In_1981,In_2157);
nand U1886 (N_1886,In_3840,N_1203);
nand U1887 (N_1887,In_2503,In_3727);
xnor U1888 (N_1888,In_1793,In_3899);
nor U1889 (N_1889,N_17,In_1657);
or U1890 (N_1890,In_1387,In_4657);
nor U1891 (N_1891,N_1380,N_476);
and U1892 (N_1892,N_801,N_666);
and U1893 (N_1893,In_3330,In_2815);
nand U1894 (N_1894,In_2713,N_873);
or U1895 (N_1895,In_2883,In_4217);
or U1896 (N_1896,In_165,In_1380);
and U1897 (N_1897,In_3184,In_2898);
or U1898 (N_1898,In_2477,N_1273);
or U1899 (N_1899,In_3742,In_2533);
nor U1900 (N_1900,In_1888,In_2709);
xor U1901 (N_1901,N_150,In_529);
and U1902 (N_1902,In_71,In_4691);
nand U1903 (N_1903,In_3908,N_27);
or U1904 (N_1904,In_4369,N_811);
and U1905 (N_1905,In_4668,N_563);
and U1906 (N_1906,In_2073,In_1627);
and U1907 (N_1907,In_4356,N_269);
xor U1908 (N_1908,In_241,In_2022);
nor U1909 (N_1909,N_1293,In_3692);
and U1910 (N_1910,In_3138,In_4826);
nor U1911 (N_1911,N_740,In_341);
xnor U1912 (N_1912,N_550,In_4646);
xor U1913 (N_1913,In_3735,N_834);
nand U1914 (N_1914,In_2,In_1598);
nand U1915 (N_1915,In_3346,In_2508);
nor U1916 (N_1916,In_2062,N_120);
nor U1917 (N_1917,In_3774,In_2624);
xnor U1918 (N_1918,N_1266,N_482);
nand U1919 (N_1919,N_1112,In_3382);
nor U1920 (N_1920,N_276,N_1412);
nor U1921 (N_1921,In_4533,In_3812);
or U1922 (N_1922,In_986,In_3828);
nor U1923 (N_1923,In_88,In_3414);
nand U1924 (N_1924,N_817,In_1980);
and U1925 (N_1925,In_4487,In_4361);
and U1926 (N_1926,N_18,In_237);
nand U1927 (N_1927,N_416,In_1374);
xnor U1928 (N_1928,In_941,N_1261);
xor U1929 (N_1929,In_2192,In_3137);
nand U1930 (N_1930,In_2339,N_1472);
and U1931 (N_1931,In_4748,In_1652);
xnor U1932 (N_1932,In_2425,In_309);
or U1933 (N_1933,In_1737,N_694);
nand U1934 (N_1934,In_3174,In_2264);
or U1935 (N_1935,N_203,N_1135);
nor U1936 (N_1936,In_4663,In_4636);
and U1937 (N_1937,N_41,In_684);
nand U1938 (N_1938,In_2045,In_166);
and U1939 (N_1939,N_531,In_1604);
and U1940 (N_1940,N_428,N_1461);
xnor U1941 (N_1941,In_2765,N_624);
or U1942 (N_1942,N_1143,In_2935);
nand U1943 (N_1943,In_2430,N_1169);
and U1944 (N_1944,In_2501,In_1933);
nor U1945 (N_1945,In_1833,In_2228);
or U1946 (N_1946,In_2877,In_338);
xor U1947 (N_1947,In_861,In_4103);
and U1948 (N_1948,In_4681,In_2410);
or U1949 (N_1949,In_1520,In_1617);
and U1950 (N_1950,In_3730,In_3500);
and U1951 (N_1951,In_3954,In_334);
and U1952 (N_1952,In_2626,N_1162);
nand U1953 (N_1953,N_616,In_3780);
and U1954 (N_1954,N_379,N_1333);
xor U1955 (N_1955,N_1335,In_2978);
xor U1956 (N_1956,N_1150,N_586);
or U1957 (N_1957,In_2426,In_784);
or U1958 (N_1958,In_1350,N_63);
nor U1959 (N_1959,N_1344,N_26);
or U1960 (N_1960,In_182,N_1483);
or U1961 (N_1961,In_4496,In_390);
or U1962 (N_1962,In_4460,In_3739);
and U1963 (N_1963,N_1178,In_383);
nor U1964 (N_1964,In_3881,In_2929);
nand U1965 (N_1965,N_1473,In_1131);
or U1966 (N_1966,In_3042,N_1306);
nor U1967 (N_1967,In_1856,N_1435);
or U1968 (N_1968,N_478,In_1056);
xor U1969 (N_1969,In_2327,In_91);
xor U1970 (N_1970,N_909,In_3484);
or U1971 (N_1971,N_9,In_3598);
nor U1972 (N_1972,In_3098,N_77);
and U1973 (N_1973,In_4112,In_1688);
xnor U1974 (N_1974,N_1381,In_2521);
nor U1975 (N_1975,N_405,In_4836);
xnor U1976 (N_1976,N_830,N_589);
nand U1977 (N_1977,In_1853,In_1175);
or U1978 (N_1978,N_1177,N_1399);
xnor U1979 (N_1979,In_4372,N_254);
and U1980 (N_1980,In_3889,In_3010);
or U1981 (N_1981,In_2353,In_2571);
and U1982 (N_1982,In_2700,N_421);
nand U1983 (N_1983,In_1226,In_2377);
xor U1984 (N_1984,N_1267,N_406);
and U1985 (N_1985,In_167,N_1453);
nor U1986 (N_1986,In_4705,In_1003);
xnor U1987 (N_1987,In_3920,N_49);
nand U1988 (N_1988,In_4466,In_1317);
nand U1989 (N_1989,N_582,In_1834);
xnor U1990 (N_1990,In_2785,In_1665);
xor U1991 (N_1991,In_1113,N_1218);
nor U1992 (N_1992,N_499,N_881);
and U1993 (N_1993,In_1066,In_4299);
and U1994 (N_1994,In_3105,In_1970);
nor U1995 (N_1995,In_1599,In_4378);
xor U1996 (N_1996,In_2781,In_4134);
nand U1997 (N_1997,N_818,In_3384);
or U1998 (N_1998,In_1368,In_2996);
or U1999 (N_1999,In_4253,In_3673);
nand U2000 (N_2000,In_2757,In_1308);
or U2001 (N_2001,N_602,N_1965);
and U2002 (N_2002,In_2546,In_3223);
xor U2003 (N_2003,In_381,In_2329);
xor U2004 (N_2004,In_3084,In_1749);
xor U2005 (N_2005,In_3158,In_4355);
nor U2006 (N_2006,N_1318,In_83);
or U2007 (N_2007,In_2212,N_1350);
or U2008 (N_2008,N_334,In_4338);
xor U2009 (N_2009,In_4366,In_2860);
and U2010 (N_2010,In_2245,In_683);
nand U2011 (N_2011,N_1585,N_1184);
and U2012 (N_2012,N_230,In_4944);
nand U2013 (N_2013,In_2013,In_4452);
xnor U2014 (N_2014,N_1706,N_376);
nand U2015 (N_2015,In_667,N_1652);
nor U2016 (N_2016,In_3327,In_4823);
xor U2017 (N_2017,N_614,In_713);
xor U2018 (N_2018,N_850,N_216);
xnor U2019 (N_2019,N_1696,In_3693);
and U2020 (N_2020,In_2366,N_943);
and U2021 (N_2021,N_251,N_1395);
and U2022 (N_2022,N_1980,In_3777);
or U2023 (N_2023,In_2214,In_862);
or U2024 (N_2024,N_1160,N_807);
nand U2025 (N_2025,N_1806,In_4934);
xor U2026 (N_2026,In_2596,In_4367);
nor U2027 (N_2027,In_1361,In_1839);
xnor U2028 (N_2028,N_1836,N_1231);
nand U2029 (N_2029,In_2818,N_1644);
or U2030 (N_2030,In_2077,N_1582);
nor U2031 (N_2031,In_3664,N_19);
and U2032 (N_2032,In_3188,In_738);
or U2033 (N_2033,In_2650,N_1349);
nand U2034 (N_2034,N_1737,In_3879);
or U2035 (N_2035,In_4844,N_678);
nand U2036 (N_2036,In_2688,N_1383);
nand U2037 (N_2037,In_128,In_1508);
nor U2038 (N_2038,N_1416,In_2283);
and U2039 (N_2039,In_1515,In_2940);
and U2040 (N_2040,In_3629,In_4003);
or U2041 (N_2041,In_597,N_886);
xor U2042 (N_2042,In_3600,N_1669);
nand U2043 (N_2043,N_1125,N_1877);
or U2044 (N_2044,In_2220,In_1890);
nor U2045 (N_2045,In_4357,N_1490);
and U2046 (N_2046,In_722,In_758);
nand U2047 (N_2047,N_1546,In_3959);
nor U2048 (N_2048,In_2189,In_1110);
nor U2049 (N_2049,In_492,N_1942);
and U2050 (N_2050,In_3926,N_1827);
nand U2051 (N_2051,In_3093,N_1191);
xor U2052 (N_2052,N_1428,N_1698);
or U2053 (N_2053,In_3258,N_1408);
nand U2054 (N_2054,N_867,N_983);
and U2055 (N_2055,N_613,N_1770);
and U2056 (N_2056,N_1357,In_4927);
nand U2057 (N_2057,N_1748,N_1258);
or U2058 (N_2058,In_546,N_1959);
and U2059 (N_2059,In_3571,In_723);
xnor U2060 (N_2060,N_1889,In_293);
and U2061 (N_2061,In_3831,In_2608);
or U2062 (N_2062,In_3142,N_1275);
nor U2063 (N_2063,In_407,In_3141);
or U2064 (N_2064,N_1848,In_3504);
or U2065 (N_2065,In_1662,In_4438);
xnor U2066 (N_2066,In_2903,In_3690);
or U2067 (N_2067,In_3655,N_1502);
xnor U2068 (N_2068,N_1062,N_1767);
and U2069 (N_2069,In_1039,N_1039);
and U2070 (N_2070,In_70,In_2388);
nor U2071 (N_2071,N_1478,N_1403);
or U2072 (N_2072,N_1785,In_747);
nor U2073 (N_2073,In_3421,N_1976);
or U2074 (N_2074,In_4723,In_3680);
and U2075 (N_2075,In_3129,In_589);
or U2076 (N_2076,In_3021,N_62);
and U2077 (N_2077,In_1435,N_1804);
nand U2078 (N_2078,In_1069,In_687);
nor U2079 (N_2079,In_4345,N_636);
nor U2080 (N_2080,In_4105,In_4607);
nand U2081 (N_2081,N_1008,In_1785);
xnor U2082 (N_2082,N_1677,In_4304);
xnor U2083 (N_2083,In_3178,In_3031);
and U2084 (N_2084,In_578,In_3773);
nor U2085 (N_2085,N_812,N_1155);
xor U2086 (N_2086,In_4754,In_2637);
and U2087 (N_2087,N_1660,N_1881);
nand U2088 (N_2088,In_4473,N_566);
and U2089 (N_2089,In_1051,In_1607);
and U2090 (N_2090,N_1875,N_699);
xnor U2091 (N_2091,In_3792,In_1612);
and U2092 (N_2092,N_170,In_4194);
nor U2093 (N_2093,N_796,N_608);
nand U2094 (N_2094,N_765,N_296);
and U2095 (N_2095,In_1681,In_1406);
and U2096 (N_2096,In_373,In_1330);
nor U2097 (N_2097,In_3243,In_2305);
and U2098 (N_2098,In_1338,In_2017);
or U2099 (N_2099,N_1443,N_1810);
xnor U2100 (N_2100,N_1890,N_831);
nand U2101 (N_2101,In_245,N_1750);
nor U2102 (N_2102,In_545,In_2132);
xnor U2103 (N_2103,In_2613,N_1691);
nor U2104 (N_2104,In_982,N_1656);
or U2105 (N_2105,N_813,N_1659);
xor U2106 (N_2106,In_1725,N_1126);
and U2107 (N_2107,N_654,In_563);
or U2108 (N_2108,In_1684,In_3216);
nor U2109 (N_2109,N_123,In_2411);
or U2110 (N_2110,N_999,N_1361);
and U2111 (N_2111,N_1674,In_4278);
nor U2112 (N_2112,In_3817,N_1590);
or U2113 (N_2113,N_1635,In_3165);
nand U2114 (N_2114,In_2396,N_1041);
xnor U2115 (N_2115,In_502,N_1320);
and U2116 (N_2116,N_1382,In_4054);
xnor U2117 (N_2117,N_1463,N_1701);
nand U2118 (N_2118,In_68,N_779);
and U2119 (N_2119,In_2779,N_583);
nand U2120 (N_2120,N_1518,In_3368);
or U2121 (N_2121,In_2317,N_1681);
xnor U2122 (N_2122,In_4406,In_1982);
nor U2123 (N_2123,N_1236,N_1665);
or U2124 (N_2124,N_1196,In_2191);
and U2125 (N_2125,In_1133,In_1967);
nor U2126 (N_2126,In_935,In_4051);
xor U2127 (N_2127,In_2344,In_359);
nand U2128 (N_2128,In_2424,N_1295);
or U2129 (N_2129,N_549,N_1931);
or U2130 (N_2130,In_1979,N_78);
and U2131 (N_2131,In_2178,N_1688);
or U2132 (N_2132,N_916,In_2724);
nor U2133 (N_2133,In_2852,N_1739);
and U2134 (N_2134,In_3073,In_1929);
nand U2135 (N_2135,N_1601,In_629);
and U2136 (N_2136,N_1575,In_4521);
nor U2137 (N_2137,In_1224,In_3550);
or U2138 (N_2138,In_4261,In_950);
and U2139 (N_2139,In_3657,In_571);
and U2140 (N_2140,In_4423,In_2035);
and U2141 (N_2141,N_1554,N_1646);
or U2142 (N_2142,In_431,In_4774);
xor U2143 (N_2143,N_961,In_2330);
xnor U2144 (N_2144,N_1553,In_1234);
and U2145 (N_2145,N_949,N_617);
or U2146 (N_2146,N_789,N_839);
and U2147 (N_2147,In_2600,N_1479);
nor U2148 (N_2148,N_1016,In_230);
nor U2149 (N_2149,In_1769,N_747);
nor U2150 (N_2150,In_2291,In_4767);
nand U2151 (N_2151,N_1406,N_1558);
nor U2152 (N_2152,In_77,In_375);
nor U2153 (N_2153,N_1904,In_2881);
or U2154 (N_2154,In_1181,In_674);
and U2155 (N_2155,N_756,N_930);
or U2156 (N_2156,In_3770,N_1061);
or U2157 (N_2157,In_4909,N_805);
nor U2158 (N_2158,N_1626,N_1386);
nor U2159 (N_2159,N_547,In_712);
nor U2160 (N_2160,In_4784,N_1523);
and U2161 (N_2161,In_4067,In_3431);
nor U2162 (N_2162,In_631,N_1327);
and U2163 (N_2163,In_3260,N_1276);
or U2164 (N_2164,N_836,N_1532);
xnor U2165 (N_2165,N_764,In_11);
and U2166 (N_2166,In_4472,N_1825);
or U2167 (N_2167,N_1708,In_3604);
or U2168 (N_2168,In_4096,N_1823);
xor U2169 (N_2169,In_4030,In_138);
or U2170 (N_2170,In_2769,In_831);
nand U2171 (N_2171,N_1918,In_1628);
nor U2172 (N_2172,In_4674,In_3838);
nand U2173 (N_2173,In_1675,N_1715);
and U2174 (N_2174,N_1882,N_1080);
nor U2175 (N_2175,In_4865,N_1482);
nand U2176 (N_2176,N_1913,In_1314);
xor U2177 (N_2177,N_1407,N_1452);
or U2178 (N_2178,N_1630,In_2125);
and U2179 (N_2179,In_248,N_1969);
and U2180 (N_2180,In_2579,N_1740);
or U2181 (N_2181,N_327,N_142);
nand U2182 (N_2182,In_996,N_1168);
and U2183 (N_2183,N_1190,N_1851);
xor U2184 (N_2184,In_1015,In_4842);
and U2185 (N_2185,In_4701,In_4945);
or U2186 (N_2186,N_74,In_2658);
nor U2187 (N_2187,In_326,N_32);
and U2188 (N_2188,In_3217,In_3248);
nor U2189 (N_2189,N_1824,In_2934);
or U2190 (N_2190,N_1619,In_1229);
or U2191 (N_2191,In_4926,In_3365);
or U2192 (N_2192,In_4129,In_805);
nand U2193 (N_2193,N_175,N_1572);
nor U2194 (N_2194,In_162,In_4552);
nor U2195 (N_2195,In_2752,N_754);
nor U2196 (N_2196,N_1250,N_1923);
nand U2197 (N_2197,N_1738,N_1879);
nand U2198 (N_2198,N_1455,N_323);
nor U2199 (N_2199,In_1413,N_701);
nand U2200 (N_2200,In_4480,In_2391);
nor U2201 (N_2201,In_324,N_136);
xnor U2202 (N_2202,N_1650,In_1972);
or U2203 (N_2203,N_1963,N_240);
xnor U2204 (N_2204,In_3978,In_2728);
xor U2205 (N_2205,N_1202,In_2716);
nand U2206 (N_2206,In_2721,N_1087);
xnor U2207 (N_2207,N_87,N_800);
nor U2208 (N_2208,In_3262,In_734);
and U2209 (N_2209,In_4202,In_4717);
nor U2210 (N_2210,In_602,In_240);
or U2211 (N_2211,N_1322,N_1730);
or U2212 (N_2212,N_1903,In_4205);
nor U2213 (N_2213,N_1137,In_4386);
and U2214 (N_2214,In_2890,N_1581);
nor U2215 (N_2215,In_108,In_3837);
nor U2216 (N_2216,In_4574,In_3283);
nor U2217 (N_2217,N_1616,In_3728);
and U2218 (N_2218,N_314,N_1710);
nor U2219 (N_2219,In_3589,In_588);
nand U2220 (N_2220,N_220,N_1916);
nor U2221 (N_2221,N_1181,N_1759);
or U2222 (N_2222,In_634,N_1339);
or U2223 (N_2223,In_860,N_1373);
nand U2224 (N_2224,N_1232,In_4508);
xnor U2225 (N_2225,In_538,N_1880);
xor U2226 (N_2226,In_252,In_3981);
or U2227 (N_2227,In_1758,N_904);
nand U2228 (N_2228,In_761,N_774);
and U2229 (N_2229,N_853,N_1624);
nand U2230 (N_2230,In_1936,N_1265);
or U2231 (N_2231,In_3264,N_1854);
nor U2232 (N_2232,N_1636,In_3609);
and U2233 (N_2233,In_2926,In_3984);
and U2234 (N_2234,N_1743,In_639);
or U2235 (N_2235,N_1514,N_1884);
or U2236 (N_2236,N_1217,In_1386);
nor U2237 (N_2237,N_1818,In_2056);
nand U2238 (N_2238,N_1257,In_2030);
nor U2239 (N_2239,N_378,In_518);
nand U2240 (N_2240,N_928,In_2493);
or U2241 (N_2241,In_4207,In_1905);
xor U2242 (N_2242,N_870,N_1151);
or U2243 (N_2243,In_3192,In_2828);
xor U2244 (N_2244,N_465,N_1521);
or U2245 (N_2245,In_1664,In_4694);
nand U2246 (N_2246,N_437,N_1438);
and U2247 (N_2247,In_2181,In_2309);
xor U2248 (N_2248,N_947,In_2047);
nand U2249 (N_2249,In_2930,In_3022);
xor U2250 (N_2250,In_4432,In_3130);
nor U2251 (N_2251,In_2147,N_1362);
nand U2252 (N_2252,In_796,N_1298);
or U2253 (N_2253,In_3288,N_1180);
nand U2254 (N_2254,N_516,N_1358);
xor U2255 (N_2255,In_4532,In_1937);
or U2256 (N_2256,N_1781,N_1912);
xnor U2257 (N_2257,In_1788,N_749);
and U2258 (N_2258,In_1169,N_389);
or U2259 (N_2259,N_158,In_583);
nor U2260 (N_2260,In_3358,In_2548);
and U2261 (N_2261,N_321,In_4768);
xor U2262 (N_2262,N_741,N_1887);
nor U2263 (N_2263,N_1456,N_523);
nor U2264 (N_2264,N_1686,In_4258);
nand U2265 (N_2265,In_2238,In_3980);
xor U2266 (N_2266,In_3291,N_671);
nor U2267 (N_2267,In_1298,In_3114);
nor U2268 (N_2268,In_2438,N_1653);
or U2269 (N_2269,In_632,In_4239);
nor U2270 (N_2270,In_611,N_1899);
and U2271 (N_2271,In_676,In_1700);
nand U2272 (N_2272,N_100,In_3240);
xor U2273 (N_2273,In_4580,In_2941);
xnor U2274 (N_2274,In_1490,N_1447);
xnor U2275 (N_2275,In_2319,In_2841);
nand U2276 (N_2276,In_4076,In_2853);
nor U2277 (N_2277,N_539,In_2505);
nand U2278 (N_2278,N_289,N_1173);
or U2279 (N_2279,In_1372,In_3435);
nand U2280 (N_2280,N_684,N_958);
xnor U2281 (N_2281,In_802,In_2092);
nand U2282 (N_2282,N_1049,In_3136);
or U2283 (N_2283,In_587,N_1775);
and U2284 (N_2284,In_4882,In_376);
nor U2285 (N_2285,In_4976,N_1939);
nand U2286 (N_2286,In_3038,In_467);
xor U2287 (N_2287,N_1494,In_4376);
and U2288 (N_2288,In_1958,In_1414);
and U2289 (N_2289,In_423,In_1781);
nor U2290 (N_2290,N_1798,N_1697);
or U2291 (N_2291,N_1869,N_433);
nand U2292 (N_2292,N_718,N_173);
nand U2293 (N_2293,N_1017,N_1346);
nor U2294 (N_2294,N_1290,In_4515);
and U2295 (N_2295,N_1136,In_4529);
nand U2296 (N_2296,N_977,In_3205);
and U2297 (N_2297,In_142,In_4341);
and U2298 (N_2298,N_1026,In_1616);
xnor U2299 (N_2299,In_4184,In_3751);
xor U2300 (N_2300,In_2000,In_2804);
and U2301 (N_2301,N_1394,N_144);
and U2302 (N_2302,N_311,In_2112);
or U2303 (N_2303,In_3532,In_3275);
and U2304 (N_2304,N_985,In_4075);
and U2305 (N_2305,In_255,In_1334);
nand U2306 (N_2306,N_1347,N_1766);
nand U2307 (N_2307,In_115,In_2161);
and U2308 (N_2308,N_630,N_1405);
nand U2309 (N_2309,N_1746,In_1287);
xnor U2310 (N_2310,In_3027,In_3705);
or U2311 (N_2311,In_2468,N_1375);
xor U2312 (N_2312,In_3457,In_3925);
nand U2313 (N_2313,In_4683,In_4721);
xor U2314 (N_2314,In_450,In_2762);
nand U2315 (N_2315,In_4975,In_1071);
nand U2316 (N_2316,N_1083,In_947);
nor U2317 (N_2317,In_3214,N_1384);
or U2318 (N_2318,N_1458,In_2537);
or U2319 (N_2319,N_646,In_2790);
or U2320 (N_2320,N_1941,N_1620);
xnor U2321 (N_2321,In_3991,In_957);
nor U2322 (N_2322,N_1519,N_1005);
nor U2323 (N_2323,N_1496,N_229);
nor U2324 (N_2324,N_1911,N_1807);
or U2325 (N_2325,N_1296,N_1769);
nand U2326 (N_2326,In_4318,In_3494);
or U2327 (N_2327,In_3850,In_14);
xor U2328 (N_2328,In_1741,In_2441);
nand U2329 (N_2329,N_1424,N_533);
or U2330 (N_2330,N_366,N_844);
nor U2331 (N_2331,In_1885,In_4873);
xnor U2332 (N_2332,N_637,In_380);
and U2333 (N_2333,N_361,N_887);
and U2334 (N_2334,In_1867,In_1325);
nor U2335 (N_2335,In_2549,In_552);
and U2336 (N_2336,N_316,In_3333);
or U2337 (N_2337,N_920,N_1524);
xor U2338 (N_2338,N_1666,N_1615);
nand U2339 (N_2339,N_382,N_1351);
nor U2340 (N_2340,N_1477,N_221);
nand U2341 (N_2341,In_2631,In_3331);
or U2342 (N_2342,In_2601,In_3967);
xnor U2343 (N_2343,In_4591,N_1771);
and U2344 (N_2344,N_1580,N_1702);
and U2345 (N_2345,N_1309,In_2754);
or U2346 (N_2346,In_389,In_3733);
or U2347 (N_2347,N_605,In_2756);
or U2348 (N_2348,N_291,N_570);
nor U2349 (N_2349,N_1703,N_1679);
or U2350 (N_2350,In_4764,In_3061);
or U2351 (N_2351,In_4492,In_3890);
and U2352 (N_2352,N_1509,In_1636);
and U2353 (N_2353,N_1091,In_4887);
nand U2354 (N_2354,N_975,In_1997);
nand U2355 (N_2355,In_1313,N_721);
nand U2356 (N_2356,N_679,In_1153);
nand U2357 (N_2357,N_1093,In_3449);
nand U2358 (N_2358,In_906,In_523);
and U2359 (N_2359,N_959,N_771);
nand U2360 (N_2360,In_1284,In_1456);
nor U2361 (N_2361,In_1709,In_1902);
nor U2362 (N_2362,N_114,In_3456);
xnor U2363 (N_2363,In_2740,In_2392);
nand U2364 (N_2364,N_1856,In_4399);
or U2365 (N_2365,N_1067,N_1158);
nand U2366 (N_2366,In_3736,N_1789);
xor U2367 (N_2367,N_1409,N_879);
xnor U2368 (N_2368,In_2837,N_420);
or U2369 (N_2369,In_2865,N_88);
nand U2370 (N_2370,In_2675,N_871);
nand U2371 (N_2371,N_1589,In_4635);
nor U2372 (N_2372,In_4977,In_2985);
or U2373 (N_2373,N_1920,In_3418);
or U2374 (N_2374,In_2454,In_3450);
nand U2375 (N_2375,N_1778,N_1095);
xnor U2376 (N_2376,In_2582,N_984);
and U2377 (N_2377,In_4463,N_1611);
or U2378 (N_2378,In_596,N_1813);
xnor U2379 (N_2379,N_1946,N_1499);
nor U2380 (N_2380,In_1430,In_1289);
and U2381 (N_2381,N_72,In_4156);
nor U2382 (N_2382,N_1057,In_3796);
nand U2383 (N_2383,N_1014,N_1462);
xnor U2384 (N_2384,N_431,In_4426);
nand U2385 (N_2385,In_23,In_1082);
nand U2386 (N_2386,In_3914,In_4211);
nor U2387 (N_2387,N_1139,N_1247);
nand U2388 (N_2388,N_1894,In_331);
or U2389 (N_2389,N_1986,In_3254);
or U2390 (N_2390,In_2385,In_111);
and U2391 (N_2391,N_1101,In_1016);
or U2392 (N_2392,In_3039,In_1751);
xnor U2393 (N_2393,In_4501,In_3235);
or U2394 (N_2394,N_702,In_4490);
nand U2395 (N_2395,In_2418,In_4091);
nand U2396 (N_2396,In_972,N_1467);
nand U2397 (N_2397,In_3709,In_770);
nor U2398 (N_2398,N_1253,N_1426);
nand U2399 (N_2399,In_2961,In_4485);
and U2400 (N_2400,N_1515,In_460);
nand U2401 (N_2401,N_82,In_1040);
nor U2402 (N_2402,In_94,In_4362);
nand U2403 (N_2403,In_1115,N_1045);
nor U2404 (N_2404,N_826,N_231);
and U2405 (N_2405,In_859,N_991);
and U2406 (N_2406,In_3695,In_4732);
nor U2407 (N_2407,In_1266,In_4170);
and U2408 (N_2408,In_3324,In_358);
nor U2409 (N_2409,N_356,N_1951);
and U2410 (N_2410,In_1085,N_35);
or U2411 (N_2411,N_579,N_1516);
nor U2412 (N_2412,In_3150,N_138);
or U2413 (N_2413,N_1300,In_3830);
and U2414 (N_2414,In_1109,In_2230);
and U2415 (N_2415,In_2572,N_1925);
xnor U2416 (N_2416,N_1501,In_4968);
and U2417 (N_2417,N_832,N_1304);
or U2418 (N_2418,N_925,In_2755);
and U2419 (N_2419,N_1225,N_263);
xor U2420 (N_2420,In_2284,N_704);
nand U2421 (N_2421,In_1736,In_2311);
nand U2422 (N_2422,In_3823,N_1459);
and U2423 (N_2423,N_1221,In_4955);
nor U2424 (N_2424,N_1627,In_2042);
and U2425 (N_2425,N_938,In_1857);
xnor U2426 (N_2426,N_767,In_1974);
nand U2427 (N_2427,In_991,N_1861);
nand U2428 (N_2428,In_1120,In_3945);
nor U2429 (N_2429,N_922,In_112);
and U2430 (N_2430,In_151,N_506);
or U2431 (N_2431,N_1832,In_2500);
or U2432 (N_2432,In_286,In_4614);
xor U2433 (N_2433,N_1910,N_1299);
nor U2434 (N_2434,In_3,In_369);
xor U2435 (N_2435,In_613,N_1280);
nor U2436 (N_2436,In_1276,In_559);
nor U2437 (N_2437,In_4448,N_1747);
xor U2438 (N_2438,In_4680,In_2135);
xnor U2439 (N_2439,In_2677,In_1968);
nor U2440 (N_2440,In_4203,N_992);
xor U2441 (N_2441,N_1038,In_147);
xnor U2442 (N_2442,N_1664,In_1920);
and U2443 (N_2443,In_2347,In_3566);
nor U2444 (N_2444,In_1449,In_1724);
or U2445 (N_2445,N_1973,N_1368);
xnor U2446 (N_2446,N_326,In_1531);
xnor U2447 (N_2447,N_1042,N_1374);
nor U2448 (N_2448,N_1983,In_1105);
and U2449 (N_2449,In_726,In_3131);
or U2450 (N_2450,In_1878,N_1100);
nor U2451 (N_2451,In_1587,N_1123);
nor U2452 (N_2452,In_205,In_4087);
nand U2453 (N_2453,In_2564,In_2398);
or U2454 (N_2454,In_533,N_272);
nor U2455 (N_2455,In_4488,In_3672);
and U2456 (N_2456,In_2743,N_1994);
or U2457 (N_2457,N_1507,In_4288);
nand U2458 (N_2458,In_3776,In_1020);
or U2459 (N_2459,In_4847,N_635);
nor U2460 (N_2460,In_2687,N_1849);
or U2461 (N_2461,In_2842,N_418);
and U2462 (N_2462,N_1090,N_1718);
and U2463 (N_2463,N_299,N_1752);
xor U2464 (N_2464,N_572,N_880);
nand U2465 (N_2465,In_2084,In_143);
nand U2466 (N_2466,In_4149,In_1103);
xor U2467 (N_2467,N_1471,In_1489);
and U2468 (N_2468,N_1118,N_1517);
nor U2469 (N_2469,N_1915,In_3422);
or U2470 (N_2470,N_1513,In_284);
and U2471 (N_2471,N_1922,In_1278);
nand U2472 (N_2472,N_1905,In_3463);
nand U2473 (N_2473,N_184,In_4974);
and U2474 (N_2474,N_148,N_226);
and U2475 (N_2475,In_1791,N_1329);
nor U2476 (N_2476,N_1993,In_424);
nor U2477 (N_2477,N_1549,N_348);
xnor U2478 (N_2478,N_208,N_507);
xor U2479 (N_2479,In_721,In_2290);
xor U2480 (N_2480,In_2686,In_2796);
or U2481 (N_2481,In_2710,N_1044);
xnor U2482 (N_2482,In_811,In_4751);
xor U2483 (N_2483,In_3033,N_355);
nand U2484 (N_2484,In_4005,N_1147);
xor U2485 (N_2485,N_1596,N_498);
and U2486 (N_2486,In_3821,In_3895);
nor U2487 (N_2487,In_4,In_4904);
nor U2488 (N_2488,N_1237,In_871);
xnor U2489 (N_2489,N_929,In_2809);
nor U2490 (N_2490,In_76,In_2982);
nand U2491 (N_2491,In_4763,In_2795);
xnor U2492 (N_2492,In_506,In_2052);
and U2493 (N_2493,In_829,N_1663);
and U2494 (N_2494,In_3833,In_1886);
nand U2495 (N_2495,In_3851,N_890);
nand U2496 (N_2496,In_13,In_4328);
and U2497 (N_2497,N_165,N_1536);
or U2498 (N_2498,N_1864,N_1153);
nor U2499 (N_2499,N_1113,N_619);
and U2500 (N_2500,N_1676,In_4518);
nor U2501 (N_2501,In_3426,N_1640);
xnor U2502 (N_2502,N_2200,N_1895);
or U2503 (N_2503,N_607,N_751);
nand U2504 (N_2504,In_725,In_3115);
or U2505 (N_2505,In_740,In_4392);
or U2506 (N_2506,N_1629,N_1933);
nor U2507 (N_2507,N_2392,In_139);
and U2508 (N_2508,In_564,In_876);
nand U2509 (N_2509,In_2726,N_1948);
nand U2510 (N_2510,N_441,N_1085);
or U2511 (N_2511,In_4816,N_1945);
and U2512 (N_2512,In_1532,N_2403);
nor U2513 (N_2513,In_55,N_1115);
nor U2514 (N_2514,In_2691,In_3470);
xor U2515 (N_2515,In_4474,N_2358);
and U2516 (N_2516,N_1032,N_1732);
xnor U2517 (N_2517,In_4303,N_1543);
nor U2518 (N_2518,In_2297,In_307);
nand U2519 (N_2519,N_1874,In_3133);
nand U2520 (N_2520,In_1803,N_2110);
nor U2521 (N_2521,N_1811,In_828);
nand U2522 (N_2522,In_1081,N_1522);
nor U2523 (N_2523,N_2378,In_1835);
xor U2524 (N_2524,N_2149,N_132);
and U2525 (N_2525,In_3143,N_2404);
nand U2526 (N_2526,In_2723,In_1064);
or U2527 (N_2527,In_323,N_2319);
nand U2528 (N_2528,N_2480,In_1378);
nand U2529 (N_2529,In_1024,In_1275);
and U2530 (N_2530,In_4409,In_755);
nand U2531 (N_2531,In_1580,In_281);
nor U2532 (N_2532,N_816,N_1648);
nand U2533 (N_2533,In_3520,In_666);
xnor U2534 (N_2534,N_1504,N_2076);
or U2535 (N_2535,In_3342,In_1163);
or U2536 (N_2536,N_1410,In_553);
and U2537 (N_2537,N_2112,N_1858);
or U2538 (N_2538,In_2830,In_1705);
nand U2539 (N_2539,N_1259,N_2376);
nand U2540 (N_2540,N_1128,N_599);
and U2541 (N_2541,In_7,In_2267);
and U2542 (N_2542,N_2073,In_2233);
and U2543 (N_2543,N_595,In_1574);
xor U2544 (N_2544,In_2534,N_1921);
nand U2545 (N_2545,In_4973,N_1613);
nand U2546 (N_2546,N_2005,N_2287);
or U2547 (N_2547,N_517,In_1601);
nand U2548 (N_2548,N_1949,N_292);
nor U2549 (N_2549,In_1910,N_1570);
nor U2550 (N_2550,N_249,In_3483);
nor U2551 (N_2551,In_1825,In_4232);
or U2552 (N_2552,N_1274,In_2168);
nor U2553 (N_2553,N_236,N_939);
or U2554 (N_2554,N_1249,In_4586);
or U2555 (N_2555,N_139,N_2062);
nor U2556 (N_2556,N_1387,N_2482);
xnor U2557 (N_2557,In_2336,N_1909);
or U2558 (N_2558,N_1979,N_1487);
or U2559 (N_2559,In_1583,In_3169);
or U2560 (N_2560,In_4689,N_1776);
nand U2561 (N_2561,N_2194,In_1557);
or U2562 (N_2562,N_2387,N_147);
and U2563 (N_2563,In_126,N_2447);
and U2564 (N_2564,In_4637,In_4688);
nand U2565 (N_2565,N_1363,In_288);
nor U2566 (N_2566,N_808,In_2066);
nand U2567 (N_2567,In_2478,In_509);
and U2568 (N_2568,N_1577,N_394);
nand U2569 (N_2569,In_3638,In_4817);
or U2570 (N_2570,N_2428,N_2228);
and U2571 (N_2571,N_2310,In_434);
nor U2572 (N_2572,N_545,N_2486);
nor U2573 (N_2573,N_2126,In_4598);
or U2574 (N_2574,In_3286,N_2033);
nand U2575 (N_2575,In_3516,In_3913);
xnor U2576 (N_2576,N_2008,N_2271);
xnor U2577 (N_2577,N_2182,N_1056);
nand U2578 (N_2578,In_4626,N_159);
xor U2579 (N_2579,N_1685,N_2165);
or U2580 (N_2580,N_58,N_1134);
nor U2581 (N_2581,N_1567,N_753);
xnor U2582 (N_2582,In_2784,N_1814);
and U2583 (N_2583,N_822,In_3245);
and U2584 (N_2584,In_3271,N_14);
nor U2585 (N_2585,N_2125,N_2253);
xnor U2586 (N_2586,In_728,In_312);
xnor U2587 (N_2587,In_3767,N_1418);
nor U2588 (N_2588,N_1256,N_2069);
nor U2589 (N_2589,N_2240,In_807);
or U2590 (N_2590,N_1565,In_902);
xnor U2591 (N_2591,N_452,N_2470);
nand U2592 (N_2592,In_652,In_3377);
nand U2593 (N_2593,N_604,N_1484);
xor U2594 (N_2594,N_1353,N_2103);
or U2595 (N_2595,In_4726,In_3190);
xor U2596 (N_2596,N_1960,N_1185);
xor U2597 (N_2597,In_3280,In_3884);
or U2598 (N_2598,N_1209,In_2994);
nor U2599 (N_2599,N_1645,N_2262);
nor U2600 (N_2600,In_4120,N_615);
xor U2601 (N_2601,N_1855,N_423);
xnor U2602 (N_2602,N_1011,N_2329);
nand U2603 (N_2603,In_2346,N_1693);
or U2604 (N_2604,In_3526,In_1208);
nand U2605 (N_2605,N_20,N_2321);
nor U2606 (N_2606,In_2165,N_564);
xnor U2607 (N_2607,In_99,N_783);
nand U2608 (N_2608,N_1720,N_2421);
nand U2609 (N_2609,In_580,N_81);
nor U2610 (N_2610,N_2229,N_911);
xnor U2611 (N_2611,N_2087,In_1896);
nand U2612 (N_2612,N_213,N_727);
or U2613 (N_2613,In_2008,N_320);
nand U2614 (N_2614,In_4321,In_4382);
nand U2615 (N_2615,N_1243,N_2440);
nand U2616 (N_2616,N_1835,N_852);
xnor U2617 (N_2617,In_3274,N_2356);
nor U2618 (N_2618,N_2151,N_243);
or U2619 (N_2619,N_2435,N_969);
nand U2620 (N_2620,N_2374,In_3802);
nand U2621 (N_2621,N_1244,N_1857);
nor U2622 (N_2622,N_1262,In_2390);
nor U2623 (N_2623,In_1089,In_4560);
or U2624 (N_2624,N_1366,In_2959);
and U2625 (N_2625,In_3273,In_300);
nand U2626 (N_2626,N_1872,N_337);
and U2627 (N_2627,N_1199,In_3897);
or U2628 (N_2628,In_3869,N_2266);
nand U2629 (N_2629,In_4124,N_2295);
xnor U2630 (N_2630,N_2085,In_4040);
nand U2631 (N_2631,N_2070,In_4323);
nand U2632 (N_2632,N_1935,N_1116);
nor U2633 (N_2633,N_1828,N_1628);
and U2634 (N_2634,N_2192,N_1027);
or U2635 (N_2635,N_2108,In_4756);
nor U2636 (N_2636,N_51,In_332);
xnor U2637 (N_2637,N_1893,N_1655);
nand U2638 (N_2638,N_275,N_22);
and U2639 (N_2639,N_1540,N_1223);
nor U2640 (N_2640,N_2298,N_1878);
nand U2641 (N_2641,N_1021,In_2376);
nor U2642 (N_2642,In_2696,N_2397);
or U2643 (N_2643,In_794,In_2913);
or U2644 (N_2644,In_410,N_1271);
nand U2645 (N_2645,N_1595,In_3144);
xnor U2646 (N_2646,N_1968,In_4653);
nor U2647 (N_2647,N_2361,N_1850);
nor U2648 (N_2648,N_1668,N_1186);
or U2649 (N_2649,N_2464,In_2843);
and U2650 (N_2650,N_995,N_1932);
nor U2651 (N_2651,In_2394,N_655);
and U2652 (N_2652,N_2124,N_333);
nor U2653 (N_2653,In_2234,In_266);
and U2654 (N_2654,N_2036,In_3385);
and U2655 (N_2655,N_37,In_2393);
nor U2656 (N_2656,N_2299,In_4536);
or U2657 (N_2657,N_1392,In_3592);
or U2658 (N_2658,N_1962,In_4045);
and U2659 (N_2659,In_2072,N_90);
and U2660 (N_2660,In_4825,N_1505);
nor U2661 (N_2661,N_1534,N_2483);
nor U2662 (N_2662,In_3832,In_1412);
or U2663 (N_2663,N_1721,In_2252);
nand U2664 (N_2664,N_1029,In_2736);
or U2665 (N_2665,N_2465,N_2267);
xnor U2666 (N_2666,In_1712,N_1562);
nand U2667 (N_2667,In_873,In_640);
or U2668 (N_2668,In_4319,N_1050);
and U2669 (N_2669,In_3495,In_4505);
nor U2670 (N_2670,N_2268,In_3863);
and U2671 (N_2671,In_2170,In_4589);
and U2672 (N_2672,In_2068,N_180);
xnor U2673 (N_2673,N_2457,N_1588);
xnor U2674 (N_2674,In_2044,In_4077);
and U2675 (N_2675,N_304,In_2471);
xnor U2676 (N_2676,N_1820,N_2128);
nor U2677 (N_2677,N_1446,N_1977);
nand U2678 (N_2678,In_1429,N_1982);
and U2679 (N_2679,In_838,N_2446);
xnor U2680 (N_2680,In_2119,N_1830);
xor U2681 (N_2681,N_1222,In_2953);
or U2682 (N_2682,N_1326,N_719);
and U2683 (N_2683,In_1894,N_257);
or U2684 (N_2684,N_2383,N_552);
nor U2685 (N_2685,N_2285,N_2414);
xnor U2686 (N_2686,N_2123,N_1310);
or U2687 (N_2687,N_1970,In_2912);
xnor U2688 (N_2688,N_710,N_2187);
or U2689 (N_2689,In_1533,N_2216);
nor U2690 (N_2690,N_2381,In_690);
and U2691 (N_2691,N_1176,In_2981);
nand U2692 (N_2692,N_2060,In_1193);
and U2693 (N_2693,In_3574,In_850);
nor U2694 (N_2694,In_4905,N_859);
or U2695 (N_2695,In_3170,In_4287);
xor U2696 (N_2696,In_896,N_2065);
and U2697 (N_2697,N_2203,In_3106);
or U2698 (N_2698,In_2776,In_4333);
and U2699 (N_2699,In_4062,In_3554);
nor U2700 (N_2700,In_3865,N_1400);
nand U2701 (N_2701,In_923,In_3699);
xor U2702 (N_2702,N_1082,N_1316);
or U2703 (N_2703,N_1002,N_940);
or U2704 (N_2704,N_1379,In_2950);
and U2705 (N_2705,In_4682,N_1608);
xnor U2706 (N_2706,In_4609,In_3947);
xor U2707 (N_2707,In_3052,N_324);
and U2708 (N_2708,N_2016,N_2167);
or U2709 (N_2709,In_3325,N_2490);
xnor U2710 (N_2710,In_3395,In_2180);
or U2711 (N_2711,N_1314,N_1610);
and U2712 (N_2712,In_3175,N_981);
and U2713 (N_2713,N_2232,In_3543);
xor U2714 (N_2714,In_1005,In_2771);
nand U2715 (N_2715,N_1245,In_75);
nor U2716 (N_2716,N_2372,N_1966);
nor U2717 (N_2717,In_2435,In_2984);
and U2718 (N_2718,N_1684,In_4634);
or U2719 (N_2719,In_2310,In_18);
nor U2720 (N_2720,N_974,N_2154);
or U2721 (N_2721,N_283,In_1707);
xor U2722 (N_2722,N_1312,N_1385);
nand U2723 (N_2723,N_1833,In_2449);
or U2724 (N_2724,In_4457,In_2817);
xor U2725 (N_2725,In_2202,N_2422);
or U2726 (N_2726,N_1755,N_2233);
and U2727 (N_2727,N_2202,N_2044);
and U2728 (N_2728,In_350,In_843);
nor U2729 (N_2729,In_1638,N_97);
nand U2730 (N_2730,N_1157,N_731);
xor U2731 (N_2731,In_4671,N_1815);
and U2732 (N_2732,N_1633,N_463);
xor U2733 (N_2733,In_4762,In_4173);
nor U2734 (N_2734,In_2802,N_1705);
and U2735 (N_2735,N_934,In_1698);
xnor U2736 (N_2736,In_1869,In_4690);
nor U2737 (N_2737,In_2185,N_399);
and U2738 (N_2738,In_4867,In_4006);
xnor U2739 (N_2739,N_2145,In_3711);
or U2740 (N_2740,N_53,In_984);
or U2741 (N_2741,In_3164,In_4133);
nand U2742 (N_2742,N_2393,N_2015);
xor U2743 (N_2743,In_227,In_3845);
xnor U2744 (N_2744,In_2565,N_2385);
nand U2745 (N_2745,N_2411,In_823);
xor U2746 (N_2746,N_1862,N_2037);
nor U2747 (N_2747,N_2014,N_1741);
or U2748 (N_2748,In_2473,In_1033);
nor U2749 (N_2749,In_4837,In_4581);
xnor U2750 (N_2750,In_4017,In_3091);
or U2751 (N_2751,In_1196,N_2109);
xnor U2752 (N_2752,N_912,In_2148);
xnor U2753 (N_2753,In_276,N_1901);
and U2754 (N_2754,In_1913,N_1023);
and U2755 (N_2755,N_1108,N_2283);
nor U2756 (N_2756,N_1469,In_3268);
xnor U2757 (N_2757,N_2019,In_451);
xor U2758 (N_2758,In_1782,In_3132);
xnor U2759 (N_2759,N_1533,In_897);
and U2760 (N_2760,N_469,In_1383);
and U2761 (N_2761,In_4332,In_4391);
and U2762 (N_2762,N_1900,In_1640);
or U2763 (N_2763,N_590,N_1930);
nor U2764 (N_2764,N_1999,In_4233);
or U2765 (N_2765,In_4611,N_1070);
xnor U2766 (N_2766,N_28,In_1101);
xor U2767 (N_2767,In_3956,N_1242);
or U2768 (N_2768,In_275,N_1754);
or U2769 (N_2769,In_2524,N_268);
xnor U2770 (N_2770,N_2003,N_2223);
and U2771 (N_2771,In_3685,N_632);
nor U2772 (N_2772,N_1204,N_2067);
and U2773 (N_2773,In_1246,In_3499);
or U2774 (N_2774,N_1187,N_2193);
nand U2775 (N_2775,N_761,In_4861);
or U2776 (N_2776,In_2569,N_2484);
xor U2777 (N_2777,In_3632,N_1530);
nor U2778 (N_2778,N_267,N_1579);
and U2779 (N_2779,In_4971,In_2794);
nand U2780 (N_2780,In_3910,N_1390);
nor U2781 (N_2781,N_1682,N_1544);
or U2782 (N_2782,N_2280,N_2261);
nor U2783 (N_2783,In_1984,In_1643);
nand U2784 (N_2784,N_177,In_1222);
nand U2785 (N_2785,N_1958,In_4785);
or U2786 (N_2786,In_2450,N_2157);
nor U2787 (N_2787,N_2188,N_1605);
or U2788 (N_2788,In_4379,In_3095);
or U2789 (N_2789,In_955,N_1583);
nor U2790 (N_2790,N_797,In_2188);
nand U2791 (N_2791,N_1551,In_2405);
or U2792 (N_2792,In_3451,In_362);
nor U2793 (N_2793,In_1552,In_1866);
nand U2794 (N_2794,N_2418,N_706);
nor U2795 (N_2795,N_2477,In_1901);
or U2796 (N_2796,In_1068,N_1216);
nand U2797 (N_2797,N_667,N_1433);
nor U2798 (N_2798,In_3762,N_1726);
nand U2799 (N_2799,N_1670,N_1625);
nand U2800 (N_2800,N_1763,N_1121);
nand U2801 (N_2801,In_710,N_328);
or U2802 (N_2802,In_4434,N_2024);
or U2803 (N_2803,In_118,N_1792);
and U2804 (N_2804,In_2514,N_1638);
nand U2805 (N_2805,N_1226,In_2699);
nand U2806 (N_2806,In_1281,N_1198);
xor U2807 (N_2807,In_48,In_3916);
and U2808 (N_2808,N_1842,N_126);
nor U2809 (N_2809,N_1692,In_3546);
nand U2810 (N_2810,N_2454,N_2330);
nor U2811 (N_2811,N_1578,N_1512);
or U2812 (N_2812,N_1793,In_4643);
and U2813 (N_2813,In_473,In_3088);
xnor U2814 (N_2814,N_1791,N_1055);
nor U2815 (N_2815,N_1106,N_2495);
or U2816 (N_2816,N_1808,In_1667);
and U2817 (N_2817,N_1097,In_3359);
xnor U2818 (N_2818,In_1995,In_1083);
or U2819 (N_2819,In_368,In_2567);
nor U2820 (N_2820,In_367,N_680);
nand U2821 (N_2821,In_4737,In_655);
nor U2822 (N_2822,N_2023,In_382);
nand U2823 (N_2823,In_2895,N_1840);
and U2824 (N_2824,N_1012,N_54);
and U2825 (N_2825,In_2419,In_3798);
or U2826 (N_2826,N_1278,In_3703);
nor U2827 (N_2827,N_358,N_1675);
or U2828 (N_2828,N_1831,In_2349);
and U2829 (N_2829,N_2166,In_3019);
or U2830 (N_2830,In_2150,In_1692);
xnor U2831 (N_2831,In_480,N_1838);
or U2832 (N_2832,N_2496,In_4339);
and U2833 (N_2833,In_780,N_29);
nand U2834 (N_2834,In_2974,N_2175);
or U2835 (N_2835,In_1279,In_3766);
nand U2836 (N_2836,N_1317,In_3099);
xor U2837 (N_2837,In_3076,N_2173);
nor U2838 (N_2838,N_2029,N_1809);
xnor U2839 (N_2839,In_4245,N_1319);
nand U2840 (N_2840,In_61,N_1657);
or U2841 (N_2841,N_106,In_1388);
or U2842 (N_2842,N_1984,N_2102);
and U2843 (N_2843,N_2026,In_4714);
and U2844 (N_2844,N_2423,N_2021);
or U2845 (N_2845,In_1422,In_3997);
or U2846 (N_2846,N_1800,N_2155);
xnor U2847 (N_2847,N_1768,N_295);
nand U2848 (N_2848,N_1024,N_11);
and U2849 (N_2849,In_3173,N_2066);
nor U2850 (N_2850,N_2186,N_2391);
nor U2851 (N_2851,In_815,N_2335);
xor U2852 (N_2852,In_1305,In_3847);
nand U2853 (N_2853,N_1537,In_3696);
nand U2854 (N_2854,In_4305,N_1690);
and U2855 (N_2855,In_4292,In_432);
and U2856 (N_2856,In_215,N_1972);
and U2857 (N_2857,N_1950,N_1064);
nor U2858 (N_2858,In_4327,N_1762);
or U2859 (N_2859,N_712,N_2050);
or U2860 (N_2860,N_2409,N_2281);
nand U2861 (N_2861,N_1821,N_1529);
xor U2862 (N_2862,In_3045,N_1926);
or U2863 (N_2863,In_2421,N_2000);
nand U2864 (N_2864,N_2022,In_900);
or U2865 (N_2865,In_322,In_3065);
nor U2866 (N_2866,N_1179,N_2147);
nor U2867 (N_2867,In_2164,In_3231);
nor U2868 (N_2868,N_2315,N_2270);
and U2869 (N_2869,In_4769,In_1817);
and U2870 (N_2870,N_1673,N_1367);
and U2871 (N_2871,In_3448,In_4999);
nand U2872 (N_2872,In_3880,In_2801);
nand U2873 (N_2873,In_4393,In_3935);
nand U2874 (N_2874,In_2033,N_1454);
xor U2875 (N_2875,In_4538,N_1761);
nor U2876 (N_2876,In_3396,In_4583);
nand U2877 (N_2877,N_1541,In_4322);
xnor U2878 (N_2878,N_2251,N_1015);
nor U2879 (N_2879,In_1554,N_606);
xor U2880 (N_2880,In_2078,In_3731);
and U2881 (N_2881,N_2220,N_1448);
and U2882 (N_2882,N_846,In_3182);
nor U2883 (N_2883,N_681,N_1928);
nor U2884 (N_2884,N_878,N_823);
nand U2885 (N_2885,N_92,In_2850);
xor U2886 (N_2886,N_2027,In_918);
nand U2887 (N_2887,In_1614,N_858);
nor U2888 (N_2888,In_1809,N_1704);
nand U2889 (N_2889,N_1078,N_2197);
and U2890 (N_2890,N_2325,In_4475);
nor U2891 (N_2891,N_913,N_2237);
or U2892 (N_2892,In_2294,In_484);
or U2893 (N_2893,In_2254,N_2412);
xnor U2894 (N_2894,N_2056,In_3305);
and U2895 (N_2895,N_1211,N_664);
or U2896 (N_2896,N_398,N_1722);
nor U2897 (N_2897,N_2399,In_763);
xnor U2898 (N_2898,In_3514,In_1248);
and U2899 (N_2899,N_2088,In_3993);
nand U2900 (N_2900,N_277,In_3861);
nor U2901 (N_2901,In_530,N_61);
or U2902 (N_2902,In_3917,N_895);
nand U2903 (N_2903,N_2068,In_3870);
nand U2904 (N_2904,In_106,In_1106);
nand U2905 (N_2905,N_752,In_2657);
or U2906 (N_2906,N_1034,N_2278);
or U2907 (N_2907,In_3533,N_322);
nand U2908 (N_2908,N_2456,N_2386);
nor U2909 (N_2909,In_4331,In_4298);
nor U2910 (N_2910,In_1800,N_780);
nand U2911 (N_2911,N_1341,N_468);
xnor U2912 (N_2912,N_1643,N_1084);
xnor U2913 (N_2913,N_2394,N_2401);
nor U2914 (N_2914,In_3117,In_2239);
and U2915 (N_2915,In_1205,In_1861);
nand U2916 (N_2916,N_2035,In_4875);
and U2917 (N_2917,N_1268,N_307);
or U2918 (N_2918,N_644,N_2277);
or U2919 (N_2919,N_2263,In_711);
and U2920 (N_2920,In_4227,In_500);
and U2921 (N_2921,In_848,In_4014);
nor U2922 (N_2922,N_1991,N_2196);
or U2923 (N_2923,N_2142,In_317);
or U2924 (N_2924,N_2293,N_211);
or U2925 (N_2925,N_2450,N_1154);
nand U2926 (N_2926,N_1780,In_3299);
nand U2927 (N_2927,In_3179,N_2028);
nor U2928 (N_2928,In_3668,N_2105);
or U2929 (N_2929,N_1765,In_938);
and U2930 (N_2930,N_1707,N_691);
and U2931 (N_2931,N_1873,In_1656);
or U2932 (N_2932,In_3127,In_4892);
or U2933 (N_2933,In_2510,N_2095);
xnor U2934 (N_2934,N_1345,N_1215);
nand U2935 (N_2935,N_1552,In_2937);
nor U2936 (N_2936,N_1460,In_3232);
nand U2937 (N_2937,In_1407,In_2770);
nor U2938 (N_2938,N_2320,N_2297);
nand U2939 (N_2939,In_1971,N_1285);
xor U2940 (N_2940,In_3617,In_3265);
and U2941 (N_2941,N_1074,N_2489);
nand U2942 (N_2942,N_1661,N_152);
xnor U2943 (N_2943,N_519,In_116);
nor U2944 (N_2944,In_4724,In_101);
or U2945 (N_2945,In_258,In_1850);
nand U2946 (N_2946,In_3710,N_1526);
or U2947 (N_2947,In_3541,N_1165);
xnor U2948 (N_2948,In_736,N_2282);
and U2949 (N_2949,N_1022,N_1545);
nor U2950 (N_2950,In_3540,N_629);
or U2951 (N_2951,In_4013,In_3573);
or U2952 (N_2952,N_897,N_2221);
nor U2953 (N_2953,N_1593,N_1525);
or U2954 (N_2954,N_2180,N_2213);
nand U2955 (N_2955,In_4208,In_2528);
xor U2956 (N_2956,N_2474,N_1528);
nand U2957 (N_2957,N_2499,N_683);
nand U2958 (N_2958,N_1883,In_2523);
nand U2959 (N_2959,N_978,N_1124);
xnor U2960 (N_2960,N_501,In_4621);
or U2961 (N_2961,N_2244,In_2456);
and U2962 (N_2962,In_223,In_1322);
and U2963 (N_2963,N_1283,In_2931);
nor U2964 (N_2964,N_2207,In_2857);
or U2965 (N_2965,In_513,In_1102);
xnor U2966 (N_2966,In_949,N_1784);
or U2967 (N_2967,N_932,N_1205);
xnor U2968 (N_2968,In_2221,N_669);
and U2969 (N_2969,In_4174,In_1504);
and U2970 (N_2970,N_1531,N_1556);
or U2971 (N_2971,In_4644,In_4803);
nor U2972 (N_2972,N_2048,In_4599);
xnor U2973 (N_2973,In_2395,In_732);
and U2974 (N_2974,N_522,N_1649);
xor U2975 (N_2975,N_1745,In_2897);
xnor U2976 (N_2976,N_1075,N_708);
nand U2977 (N_2977,N_2306,N_1886);
nor U2978 (N_2978,N_1206,N_1742);
and U2979 (N_2979,N_1289,N_2079);
nand U2980 (N_2980,In_3940,N_1195);
nor U2981 (N_2981,In_2193,In_4191);
or U2982 (N_2982,In_2198,In_4540);
or U2983 (N_2983,In_1366,In_4016);
and U2984 (N_2984,N_1749,N_1105);
or U2985 (N_2985,N_2336,In_4815);
xnor U2986 (N_2986,N_622,In_1485);
and U2987 (N_2987,In_2844,N_2437);
nand U2988 (N_2988,N_2059,In_1536);
nand U2989 (N_2989,N_119,N_1149);
xnor U2990 (N_2990,In_2130,N_2260);
and U2991 (N_2991,N_1622,In_3110);
or U2992 (N_2992,N_2045,N_1119);
nand U2993 (N_2993,N_2494,N_1538);
or U2994 (N_2994,In_1761,In_3961);
and U2995 (N_2995,N_848,In_402);
and U2996 (N_2996,In_4265,N_1129);
nand U2997 (N_2997,In_4676,N_1758);
or U2998 (N_2998,In_4578,In_2517);
xnor U2999 (N_2999,N_1422,In_1752);
and U3000 (N_3000,In_2486,N_1355);
xor U3001 (N_3001,In_1592,In_4759);
and U3002 (N_3002,In_1107,N_2398);
or U3003 (N_3003,N_1470,In_4213);
or U3004 (N_3004,In_857,N_837);
nand U3005 (N_3005,N_2864,N_1060);
nand U3006 (N_3006,N_2098,N_514);
and U3007 (N_3007,N_733,In_1928);
nand U3008 (N_3008,N_2309,N_2375);
and U3009 (N_3009,N_1311,N_183);
xor U3010 (N_3010,N_1826,N_489);
or U3011 (N_3011,In_3281,N_2672);
nand U3012 (N_3012,N_551,N_2168);
nor U3013 (N_3013,N_1906,N_2684);
or U3014 (N_3014,N_2322,In_1768);
nand U3015 (N_3015,N_2350,N_2296);
or U3016 (N_3016,N_370,In_218);
or U3017 (N_3017,N_2535,N_1975);
nor U3018 (N_3018,In_301,N_2812);
nand U3019 (N_3019,N_1360,N_775);
and U3020 (N_3020,N_2370,N_2837);
nand U3021 (N_3021,In_615,N_1573);
or U3022 (N_3022,N_709,In_1893);
nor U3023 (N_3023,N_1846,N_1837);
and U3024 (N_3024,In_2798,N_2866);
xnor U3025 (N_3025,In_964,N_2549);
nand U3026 (N_3026,N_2658,N_2692);
or U3027 (N_3027,N_1724,N_2835);
and U3028 (N_3028,N_1511,N_2243);
nand U3029 (N_3029,N_2536,N_2011);
nor U3030 (N_3030,N_2983,N_2257);
xor U3031 (N_3031,N_903,In_3933);
nor U3032 (N_3032,In_2308,In_2928);
or U3033 (N_3033,N_1576,N_1822);
or U3034 (N_3034,In_817,N_2586);
xnor U3035 (N_3035,In_1032,In_342);
xnor U3036 (N_3036,N_1812,In_1254);
or U3037 (N_3037,N_235,N_1520);
or U3038 (N_3038,N_2764,N_2051);
xnor U3039 (N_3039,In_4138,N_1208);
and U3040 (N_3040,N_2762,In_413);
and U3041 (N_3041,N_1104,N_450);
nor U3042 (N_3042,In_1969,N_2791);
xor U3043 (N_3043,N_2651,N_2500);
xor U3044 (N_3044,N_2531,In_4089);
nor U3045 (N_3045,N_2670,N_344);
xnor U3046 (N_3046,N_2212,In_1865);
xnor U3047 (N_3047,In_404,N_2575);
xnor U3048 (N_3048,N_2521,In_3437);
xor U3049 (N_3049,In_3825,N_2734);
or U3050 (N_3050,N_2057,N_2150);
and U3051 (N_3051,N_2827,N_2727);
xnor U3052 (N_3052,N_1388,N_1797);
or U3053 (N_3053,N_1302,In_3380);
or U3054 (N_3054,In_1200,In_4649);
nand U3055 (N_3055,N_2130,In_1004);
or U3056 (N_3056,In_1775,N_2195);
or U3057 (N_3057,In_2492,N_102);
xnor U3058 (N_3058,N_1566,N_1816);
or U3059 (N_3059,N_44,N_2425);
nand U3060 (N_3060,N_2810,N_2615);
or U3061 (N_3061,N_1637,N_2384);
or U3062 (N_3062,In_3082,N_2915);
nor U3063 (N_3063,N_1127,N_2120);
nor U3064 (N_3064,N_2099,N_2780);
nor U3065 (N_3065,In_3255,In_3263);
nor U3066 (N_3066,In_853,In_191);
or U3067 (N_3067,N_2638,In_890);
or U3068 (N_3068,N_1439,In_3250);
nand U3069 (N_3069,N_1235,N_2815);
and U3070 (N_3070,In_4959,N_2255);
xnor U3071 (N_3071,N_2679,N_2713);
or U3072 (N_3072,N_2921,N_2994);
nand U3073 (N_3073,N_2341,N_2181);
or U3074 (N_3074,N_1717,N_2807);
nor U3075 (N_3075,In_3658,N_2612);
or U3076 (N_3076,N_1885,In_2973);
xor U3077 (N_3077,In_3247,In_4340);
nor U3078 (N_3078,In_4797,In_296);
nor U3079 (N_3079,In_2406,N_2134);
or U3080 (N_3080,N_57,N_2596);
and U3081 (N_3081,In_1384,N_2633);
and U3082 (N_3082,In_2576,In_3322);
or U3083 (N_3083,N_561,In_1565);
or U3084 (N_3084,N_2113,N_2153);
xor U3085 (N_3085,N_2510,N_2595);
or U3086 (N_3086,N_1871,N_354);
and U3087 (N_3087,N_1919,N_1025);
xnor U3088 (N_3088,N_515,In_3230);
nor U3089 (N_3089,N_2647,In_1476);
nand U3090 (N_3090,N_650,N_2390);
nand U3091 (N_3091,N_2639,In_2271);
and U3092 (N_3092,N_2303,N_1073);
and U3093 (N_3093,N_2289,N_1891);
nor U3094 (N_3094,In_2217,N_2567);
or U3095 (N_3095,N_1639,In_3183);
xor U3096 (N_3096,In_4499,In_3471);
xor U3097 (N_3097,N_926,In_2479);
nor U3098 (N_3098,In_1471,N_1043);
xor U3099 (N_3099,In_912,N_2380);
and U3100 (N_3100,In_395,N_2569);
nand U3101 (N_3101,N_1727,In_1988);
xor U3102 (N_3102,N_2581,In_1623);
nand U3103 (N_3103,N_2851,In_1759);
nor U3104 (N_3104,In_3871,In_4020);
nor U3105 (N_3105,N_2184,In_610);
and U3106 (N_3106,In_2556,In_2263);
and U3107 (N_3107,In_714,In_888);
xnor U3108 (N_3108,N_877,N_2211);
xor U3109 (N_3109,In_724,In_3172);
or U3110 (N_3110,In_79,In_1063);
and U3111 (N_3111,N_2395,N_157);
xor U3112 (N_3112,N_2580,N_2745);
or U3113 (N_3113,N_2442,N_725);
and U3114 (N_3114,N_2417,In_4043);
and U3115 (N_3115,In_1060,In_4373);
nand U3116 (N_3116,In_2285,N_2118);
nor U3117 (N_3117,N_2230,N_2973);
or U3118 (N_3118,N_2231,N_2883);
nand U3119 (N_3119,N_199,In_1828);
xor U3120 (N_3120,In_841,N_2614);
nor U3121 (N_3121,N_2577,N_2975);
xor U3122 (N_3122,In_622,In_3892);
and U3123 (N_3123,N_2603,N_1756);
nand U3124 (N_3124,N_2726,In_4352);
and U3125 (N_3125,N_2879,In_4509);
nand U3126 (N_3126,N_957,N_2845);
xnor U3127 (N_3127,N_2782,In_4471);
xnor U3128 (N_3128,In_660,N_2463);
and U3129 (N_3129,N_2174,N_2628);
or U3130 (N_3130,In_2673,N_2821);
nor U3131 (N_3131,In_406,N_2101);
nor U3132 (N_3132,N_1054,N_2605);
nor U3133 (N_3133,N_2313,N_1474);
and U3134 (N_3134,N_1606,N_1867);
xnor U3135 (N_3135,N_2671,N_172);
nand U3136 (N_3136,In_1240,N_2140);
nand U3137 (N_3137,In_852,In_2274);
xnor U3138 (N_3138,N_2792,N_2055);
or U3139 (N_3139,In_3793,N_1254);
or U3140 (N_3140,N_2591,N_2985);
or U3141 (N_3141,N_2317,N_910);
or U3142 (N_3142,N_651,In_1434);
xnor U3143 (N_3143,N_2860,In_4038);
nand U3144 (N_3144,In_2778,N_2597);
or U3145 (N_3145,N_1978,N_2141);
xnor U3146 (N_3146,In_646,N_2508);
xnor U3147 (N_3147,N_2579,N_2433);
or U3148 (N_3148,In_433,N_648);
xor U3149 (N_3149,N_1985,In_1765);
and U3150 (N_3150,N_728,N_1294);
and U3151 (N_3151,N_1753,In_662);
nand U3152 (N_3152,N_2136,N_2646);
nor U3153 (N_3153,In_542,N_70);
and U3154 (N_3154,In_2061,N_951);
and U3155 (N_3155,In_244,N_1007);
xor U3156 (N_3156,N_2530,In_2261);
and U3157 (N_3157,N_2968,In_1530);
nor U3158 (N_3158,In_4736,N_2757);
or U3159 (N_3159,N_1796,N_2371);
nor U3160 (N_3160,N_793,In_2741);
nand U3161 (N_3161,In_2184,N_2804);
nand U3162 (N_3162,N_2898,N_1944);
xor U3163 (N_3163,N_2522,N_2645);
xnor U3164 (N_3164,N_2709,N_1102);
nand U3165 (N_3165,N_2678,N_790);
or U3166 (N_3166,In_261,In_3468);
or U3167 (N_3167,N_1757,N_574);
xor U3168 (N_3168,In_937,N_2675);
or U3169 (N_3169,In_534,In_3301);
and U3170 (N_3170,In_3644,N_2171);
nor U3171 (N_3171,In_2603,In_840);
and U3172 (N_3172,N_2424,In_1092);
nor U3173 (N_3173,In_715,N_2980);
nand U3174 (N_3174,In_2871,N_2674);
nand U3175 (N_3175,In_1908,In_4071);
nor U3176 (N_3176,N_2458,In_3827);
nand U3177 (N_3177,In_1527,N_1971);
or U3178 (N_3178,N_2627,N_2498);
nand U3179 (N_3179,In_4387,N_868);
xor U3180 (N_3180,N_2349,In_2093);
or U3181 (N_3181,N_2419,N_2504);
or U3182 (N_3182,In_4594,N_2957);
and U3183 (N_3183,N_2725,In_3417);
nand U3184 (N_3184,In_437,In_1555);
nor U3185 (N_3185,N_849,In_417);
and U3186 (N_3186,N_1035,N_1794);
or U3187 (N_3187,N_2867,In_370);
or U3188 (N_3188,N_1687,In_3722);
or U3189 (N_3189,N_2776,N_2618);
xor U3190 (N_3190,In_2213,In_1511);
and U3191 (N_3191,In_2639,N_2448);
nand U3192 (N_3192,N_2524,In_656);
nand U3193 (N_3193,N_1144,N_2763);
nand U3194 (N_3194,N_2491,In_826);
or U3195 (N_3195,N_2426,N_1019);
xor U3196 (N_3196,N_2626,In_4083);
or U3197 (N_3197,In_187,N_1961);
nor U3198 (N_3198,N_2509,N_2998);
xnor U3199 (N_3199,N_2723,In_73);
nor U3200 (N_3200,N_2922,N_698);
and U3201 (N_3201,N_2018,N_2354);
and U3202 (N_3202,In_2199,In_3447);
and U3203 (N_3203,N_1356,N_2528);
nor U3204 (N_3204,In_4407,In_997);
xnor U3205 (N_3205,In_1375,N_2342);
nor U3206 (N_3206,N_2686,In_657);
and U3207 (N_3207,N_1711,In_1720);
or U3208 (N_3208,N_2304,N_2224);
nand U3209 (N_3209,In_3241,N_1952);
nor U3210 (N_3210,N_1725,N_2565);
or U3211 (N_3211,In_4225,N_2460);
xnor U3212 (N_3212,In_956,N_1260);
and U3213 (N_3213,N_2129,N_48);
nand U3214 (N_3214,N_1500,N_685);
or U3215 (N_3215,N_1647,N_2570);
xnor U3216 (N_3216,In_3461,N_2363);
and U3217 (N_3217,N_2669,N_2198);
nor U3218 (N_3218,In_1146,N_1731);
xnor U3219 (N_3219,N_1503,N_308);
nand U3220 (N_3220,N_1229,N_404);
or U3221 (N_3221,In_1818,N_1004);
or U3222 (N_3222,N_2654,N_2075);
and U3223 (N_3223,In_1161,N_2160);
xor U3224 (N_3224,N_2944,In_3036);
nor U3225 (N_3225,In_1510,N_1843);
nor U3226 (N_3226,N_2388,In_2750);
nor U3227 (N_3227,N_2331,N_1506);
nand U3228 (N_3228,N_1908,In_1409);
nand U3229 (N_3229,N_2061,In_1876);
xnor U3230 (N_3230,N_955,N_2755);
or U3231 (N_3231,In_3584,N_2945);
nor U3232 (N_3232,In_3252,In_2328);
xnor U3233 (N_3233,N_2752,In_4468);
or U3234 (N_3234,In_185,N_1779);
and U3235 (N_3235,N_448,In_4143);
and U3236 (N_3236,In_2560,N_1654);
xor U3237 (N_3237,N_658,In_2630);
xor U3238 (N_3238,In_2714,N_2806);
nand U3239 (N_3239,N_2765,N_2553);
or U3240 (N_3240,N_2751,In_1858);
or U3241 (N_3241,N_50,In_2069);
nor U3242 (N_3242,N_656,In_4983);
and U3243 (N_3243,N_2637,N_2012);
xor U3244 (N_3244,N_2481,N_2183);
nor U3245 (N_3245,N_946,In_2205);
and U3246 (N_3246,In_2788,N_2487);
or U3247 (N_3247,N_538,N_2852);
nand U3248 (N_3248,In_3194,N_1451);
and U3249 (N_3249,N_1829,N_1847);
nand U3250 (N_3250,N_1307,In_2640);
xnor U3251 (N_3251,In_311,N_2933);
or U3252 (N_3252,N_1131,N_2001);
or U3253 (N_3253,N_1281,N_2226);
and U3254 (N_3254,In_2483,In_4023);
and U3255 (N_3255,N_2235,N_2238);
or U3256 (N_3256,N_2185,N_1764);
and U3257 (N_3257,N_1365,N_936);
xor U3258 (N_3258,N_2288,In_647);
nand U3259 (N_3259,N_2373,N_2929);
xnor U3260 (N_3260,N_2659,N_1286);
or U3261 (N_3261,N_2119,N_2636);
and U3262 (N_3262,N_2609,In_878);
xor U3263 (N_3263,N_1489,N_621);
and U3264 (N_3264,N_1086,In_3249);
nand U3265 (N_3265,N_2415,In_285);
and U3266 (N_3266,N_2932,N_2039);
or U3267 (N_3267,In_789,In_3176);
nor U3268 (N_3268,N_1240,In_4136);
and U3269 (N_3269,N_442,In_3511);
or U3270 (N_3270,N_1391,In_4031);
nor U3271 (N_3271,N_1076,In_4874);
and U3272 (N_3272,N_1866,N_2931);
xor U3273 (N_3273,N_2988,N_2996);
and U3274 (N_3274,N_2885,N_2090);
nor U3275 (N_3275,N_1238,N_2660);
nand U3276 (N_3276,N_1370,N_2164);
nand U3277 (N_3277,N_2908,N_2537);
nand U3278 (N_3278,In_3560,N_2733);
xor U3279 (N_3279,In_208,In_4431);
nor U3280 (N_3280,In_2552,N_1069);
nor U3281 (N_3281,N_1037,N_1156);
xor U3282 (N_3282,N_1642,N_1550);
and U3283 (N_3283,N_2492,N_2209);
nor U3284 (N_3284,N_2546,In_2819);
or U3285 (N_3285,N_1651,N_2416);
or U3286 (N_3286,N_2708,N_2700);
xnor U3287 (N_3287,N_2767,N_1539);
and U3288 (N_3288,In_4869,N_2308);
nor U3289 (N_3289,N_1917,N_2786);
and U3290 (N_3290,N_453,N_2813);
and U3291 (N_3291,In_4543,In_4911);
xor U3292 (N_3292,N_2870,In_3852);
nor U3293 (N_3293,In_864,N_2959);
nor U3294 (N_3294,In_1123,In_1823);
nor U3295 (N_3295,N_1592,N_2972);
nor U3296 (N_3296,N_2252,In_2821);
nand U3297 (N_3297,In_3645,N_2302);
and U3298 (N_3298,N_1863,N_821);
and U3299 (N_3299,N_1587,N_663);
xor U3300 (N_3300,N_2248,N_1109);
and U3301 (N_3301,N_2444,In_1474);
or U3302 (N_3302,N_1773,In_2255);
nand U3303 (N_3303,N_2720,N_1603);
or U3304 (N_3304,In_4900,In_3753);
xor U3305 (N_3305,In_4218,In_4651);
and U3306 (N_3306,In_4365,N_1658);
xnor U3307 (N_3307,N_2839,N_2892);
nor U3308 (N_3308,In_4602,N_2617);
and U3309 (N_3309,In_219,N_2602);
nor U3310 (N_3310,N_2139,In_1117);
xor U3311 (N_3311,N_1723,N_2990);
xor U3312 (N_3312,In_1975,In_1362);
and U3313 (N_3313,N_2405,N_1401);
nor U3314 (N_3314,N_2759,N_1466);
nand U3315 (N_3315,N_281,N_2402);
and U3316 (N_3316,In_315,N_2882);
xnor U3317 (N_3317,N_1694,In_2968);
or U3318 (N_3318,N_1892,In_793);
nor U3319 (N_3319,In_1185,N_1192);
and U3320 (N_3320,N_2683,N_2621);
nor U3321 (N_3321,N_2247,N_2236);
nor U3322 (N_3322,In_3918,In_4868);
nand U3323 (N_3323,N_1535,In_2095);
xnor U3324 (N_3324,N_2642,In_4656);
nor U3325 (N_3325,In_2256,N_964);
xor U3326 (N_3326,N_1068,N_1801);
xnor U3327 (N_3327,N_1040,N_2503);
nand U3328 (N_3328,N_2445,In_4144);
nor U3329 (N_3329,In_3011,N_1995);
or U3330 (N_3330,N_2993,N_174);
nor U3331 (N_3331,N_2178,N_2995);
nand U3332 (N_3332,N_2563,N_2013);
xor U3333 (N_3333,N_2662,N_2004);
xor U3334 (N_3334,N_952,N_2133);
nor U3335 (N_3335,N_2300,In_4981);
or U3336 (N_3336,In_1149,In_2307);
and U3337 (N_3337,N_2078,N_2828);
nand U3338 (N_3338,N_2469,In_3882);
xor U3339 (N_3339,N_1667,In_69);
xnor U3340 (N_3340,In_808,N_124);
xnor U3341 (N_3341,N_2156,N_402);
nor U3342 (N_3342,N_2808,N_351);
xnor U3343 (N_3343,N_2227,N_2587);
and U3344 (N_3344,In_4240,N_2657);
nor U3345 (N_3345,In_3181,N_1047);
nand U3346 (N_3346,N_1689,N_2697);
or U3347 (N_3347,N_2511,N_2523);
nor U3348 (N_3348,In_4795,In_2179);
nor U3349 (N_3349,N_1964,N_2054);
and U3350 (N_3350,In_2160,N_1210);
xor U3351 (N_3351,N_2847,In_1243);
or U3352 (N_3352,In_1719,N_2665);
or U3353 (N_3353,N_2451,N_1332);
nand U3354 (N_3354,In_254,N_2034);
xor U3355 (N_3355,In_2064,N_2775);
nand U3356 (N_3356,In_4478,N_2046);
nor U3357 (N_3357,In_4938,N_2688);
xnor U3358 (N_3358,N_2176,In_1569);
nand U3359 (N_3359,In_2115,N_1683);
or U3360 (N_3360,In_4066,N_2094);
nor U3361 (N_3361,N_748,N_2246);
and U3362 (N_3362,N_2290,N_1790);
and U3363 (N_3363,N_711,N_2953);
or U3364 (N_3364,N_2739,N_1834);
and U3365 (N_3365,In_1294,N_2740);
or U3366 (N_3366,In_751,N_1729);
xor U3367 (N_3367,N_1230,In_2504);
xor U3368 (N_3368,N_2115,N_2844);
and U3369 (N_3369,In_1730,In_585);
xnor U3370 (N_3370,N_2877,N_2601);
and U3371 (N_3371,N_2473,N_588);
xor U3372 (N_3372,N_1870,N_716);
and U3373 (N_3373,N_1152,In_2793);
nor U3374 (N_3374,In_1689,N_2091);
nor U3375 (N_3375,N_1751,N_508);
nand U3376 (N_3376,N_105,N_2007);
nor U3377 (N_3377,N_1559,N_2365);
and U3378 (N_3378,In_2355,In_4444);
or U3379 (N_3379,In_2746,N_2934);
xor U3380 (N_3380,In_3891,N_2505);
nor U3381 (N_3381,In_3896,N_2161);
nand U3382 (N_3382,N_672,In_2782);
xnor U3383 (N_3383,N_2942,N_1859);
nor U3384 (N_3384,In_536,N_2009);
and U3385 (N_3385,N_1695,In_4375);
or U3386 (N_3386,N_2360,N_792);
nand U3387 (N_3387,N_2848,In_1911);
nand U3388 (N_3388,N_2986,N_2919);
and U3389 (N_3389,N_918,N_1634);
or U3390 (N_3390,N_1030,In_2899);
and U3391 (N_3391,N_2872,N_1929);
nor U3392 (N_3392,N_2170,In_3068);
nand U3393 (N_3393,N_1234,N_2191);
nor U3394 (N_3394,N_1444,In_1620);
xnor U3395 (N_3395,N_1167,N_255);
and U3396 (N_3396,N_2053,N_2598);
nor U3397 (N_3397,In_347,In_658);
nand U3398 (N_3398,N_2876,N_2543);
xnor U3399 (N_3399,N_2805,N_2210);
xor U3400 (N_3400,N_2557,N_1599);
and U3401 (N_3401,N_924,In_3125);
nor U3402 (N_3402,In_3134,N_2080);
and U3403 (N_3403,N_1988,In_3912);
and U3404 (N_3404,N_2121,N_1876);
and U3405 (N_3405,N_2097,N_2548);
or U3406 (N_3406,In_2975,N_377);
xnor U3407 (N_3407,N_1560,N_2620);
xnor U3408 (N_3408,In_2371,N_1700);
or U3409 (N_3409,N_1103,N_1183);
and U3410 (N_3410,N_1348,N_2241);
or U3411 (N_3411,In_4276,N_2920);
nor U3412 (N_3412,N_1292,N_412);
nand U3413 (N_3413,N_1868,N_1734);
or U3414 (N_3414,In_2333,In_4542);
and U3415 (N_3415,In_1399,N_2869);
and U3416 (N_3416,N_2958,N_2894);
nor U3417 (N_3417,N_2897,N_1548);
nand U3418 (N_3418,N_2352,In_4871);
nor U3419 (N_3419,In_3643,N_2578);
and U3420 (N_3420,N_2083,N_2798);
or U3421 (N_3421,N_2208,N_2781);
xor U3422 (N_3422,N_1671,N_2369);
and U3423 (N_3423,N_2006,N_444);
or U3424 (N_3424,N_2348,N_591);
nor U3425 (N_3425,In_4029,In_4725);
nor U3426 (N_3426,N_601,N_1175);
nand U3427 (N_3427,N_829,N_2607);
nand U3428 (N_3428,N_2472,N_1013);
xor U3429 (N_3429,N_2696,In_2015);
nor U3430 (N_3430,N_2588,N_2766);
xor U3431 (N_3431,N_364,In_2380);
and U3432 (N_3432,In_3356,N_1786);
nand U3433 (N_3433,N_2324,N_2179);
or U3434 (N_3434,In_2300,N_2410);
or U3435 (N_3435,N_413,In_4461);
and U3436 (N_3436,In_891,N_330);
or U3437 (N_3437,N_2093,In_816);
nor U3438 (N_3438,In_2924,N_2842);
nand U3439 (N_3439,In_4360,In_216);
and U3440 (N_3440,In_4035,N_2868);
or U3441 (N_3441,N_163,In_954);
and U3442 (N_3442,N_84,N_2721);
nand U3443 (N_3443,N_369,In_4860);
nor U3444 (N_3444,N_2400,N_1586);
nor U3445 (N_3445,N_2682,N_1122);
or U3446 (N_3446,N_2924,In_4021);
and U3447 (N_3447,N_2653,N_363);
or U3448 (N_3448,N_2131,In_4916);
and U3449 (N_3449,In_3670,N_540);
nor U3450 (N_3450,N_1331,N_201);
nor U3451 (N_3451,In_1804,N_2438);
nand U3452 (N_3452,N_273,N_2641);
or U3453 (N_3453,N_2152,N_2629);
and U3454 (N_3454,N_1046,In_4773);
xor U3455 (N_3455,N_1712,In_3253);
xor U3456 (N_3456,In_1331,N_1591);
nor U3457 (N_3457,N_645,In_1364);
nor U3458 (N_3458,In_1649,N_2971);
or U3459 (N_3459,N_2803,N_2071);
and U3460 (N_3460,N_2312,N_1464);
nor U3461 (N_3461,N_1065,N_2576);
nand U3462 (N_3462,N_1774,In_4980);
nand U3463 (N_3463,In_2664,In_440);
and U3464 (N_3464,N_2930,N_2514);
and U3465 (N_3465,N_1398,N_2092);
nand U3466 (N_3466,N_2701,N_2327);
or U3467 (N_3467,N_950,N_2162);
nor U3468 (N_3468,N_2925,In_2034);
nand U3469 (N_3469,In_1418,N_2918);
nand U3470 (N_3470,N_2611,In_260);
xnor U3471 (N_3471,N_1547,In_3310);
nand U3472 (N_3472,In_2527,In_2764);
xnor U3473 (N_3473,N_2783,N_2789);
nand U3474 (N_3474,In_172,N_2239);
nor U3475 (N_3475,N_1308,N_2538);
and U3476 (N_3476,N_1641,In_4154);
or U3477 (N_3477,N_2286,N_577);
nor U3478 (N_3478,In_1810,N_2096);
nand U3479 (N_3479,N_2541,N_2711);
nor U3480 (N_3480,N_2562,In_1411);
or U3481 (N_3481,In_1603,N_2461);
xnor U3482 (N_3482,N_1937,N_2455);
or U3483 (N_3483,N_2199,In_2574);
nand U3484 (N_3484,N_461,N_1998);
nor U3485 (N_3485,N_2917,In_490);
nand U3486 (N_3486,In_1903,In_3811);
xnor U3487 (N_3487,In_4018,N_343);
xor U3488 (N_3488,N_2476,N_1291);
and U3489 (N_3489,N_504,In_1927);
nand U3490 (N_3490,In_415,In_3854);
xor U3491 (N_3491,N_1338,N_2038);
xnor U3492 (N_3492,N_39,N_2856);
nor U3493 (N_3493,In_1602,N_2506);
xor U3494 (N_3494,In_3146,N_2900);
nand U3495 (N_3495,N_2952,In_4661);
or U3496 (N_3496,N_2163,N_2488);
nor U3497 (N_3497,N_2825,N_1003);
or U3498 (N_3498,In_4107,N_2938);
or U3499 (N_3499,N_1369,N_2564);
nor U3500 (N_3500,N_3452,N_457);
xor U3501 (N_3501,N_3300,In_2038);
xor U3502 (N_3502,N_2946,N_411);
or U3503 (N_3503,In_1348,In_1258);
nand U3504 (N_3504,N_3347,N_2064);
xnor U3505 (N_3505,N_2613,N_3226);
nor U3506 (N_3506,N_2955,N_2853);
xor U3507 (N_3507,N_3149,N_3138);
and U3508 (N_3508,N_3121,N_1888);
and U3509 (N_3509,N_2214,N_3040);
nor U3510 (N_3510,N_2533,N_2143);
nand U3511 (N_3511,N_2784,N_2795);
and U3512 (N_3512,N_2222,N_2468);
xor U3513 (N_3513,N_3013,N_3042);
xnor U3514 (N_3514,N_3081,In_4126);
nand U3515 (N_3515,N_2794,In_3362);
nand U3516 (N_3516,N_3242,N_3409);
or U3517 (N_3517,N_3389,In_1437);
and U3518 (N_3518,N_3312,In_2885);
nor U3519 (N_3519,N_2824,In_1111);
nor U3520 (N_3520,In_3976,N_3302);
xor U3521 (N_3521,N_2190,N_3303);
nand U3522 (N_3522,N_1772,N_2761);
xnor U3523 (N_3523,In_2732,N_2030);
and U3524 (N_3524,In_3544,N_2608);
xor U3525 (N_3525,N_3442,In_4664);
xnor U3526 (N_3526,N_3498,N_3399);
nand U3527 (N_3527,N_3211,N_1631);
nor U3528 (N_3528,N_2351,In_462);
xor U3529 (N_3529,In_54,In_3804);
and U3530 (N_3530,N_2706,In_4766);
and U3531 (N_3531,N_2225,N_1956);
or U3532 (N_3532,N_1445,N_662);
and U3533 (N_3533,N_1233,N_3499);
and U3534 (N_3534,N_3333,N_2217);
and U3535 (N_3535,N_3043,N_2107);
xnor U3536 (N_3536,N_2259,N_3461);
xnor U3537 (N_3537,In_3763,N_2049);
or U3538 (N_3538,N_2816,N_1555);
xor U3539 (N_3539,N_3497,In_3236);
nor U3540 (N_3540,N_3207,N_2729);
and U3541 (N_3541,N_3221,N_2002);
and U3542 (N_3542,N_863,N_2127);
nand U3543 (N_3543,N_3202,N_3344);
nand U3544 (N_3544,In_3568,In_1545);
nor U3545 (N_3545,N_3425,N_700);
xnor U3546 (N_3546,N_768,In_3063);
nor U3547 (N_3547,N_1269,In_2232);
or U3548 (N_3548,N_640,In_304);
xnor U3549 (N_3549,In_672,N_3083);
and U3550 (N_3550,N_3435,N_3018);
nand U3551 (N_3551,N_3245,N_1372);
nor U3552 (N_3552,N_693,In_1594);
or U3553 (N_3553,N_3387,In_3826);
nor U3554 (N_3554,N_3392,N_3210);
nor U3555 (N_3555,N_2630,N_3342);
nor U3556 (N_3556,N_3106,In_1784);
xor U3557 (N_3557,N_2873,N_2497);
nand U3558 (N_3558,N_3220,In_1444);
nor U3559 (N_3559,N_3160,N_2625);
nor U3560 (N_3560,N_1248,N_3129);
nor U3561 (N_3561,N_2744,N_3096);
nor U3562 (N_3562,In_197,N_2074);
and U3563 (N_3563,N_2471,N_3477);
nand U3564 (N_3564,N_3156,N_2820);
nor U3565 (N_3565,N_2981,N_2017);
and U3566 (N_3566,N_3429,N_1006);
xor U3567 (N_3567,N_3223,In_4650);
nand U3568 (N_3568,N_2632,N_3157);
xnor U3569 (N_3569,N_2772,N_2616);
and U3570 (N_3570,In_2889,N_618);
and U3571 (N_3571,N_3430,N_3325);
and U3572 (N_3572,In_2558,N_1063);
nand U3573 (N_3573,In_222,N_1148);
xnor U3574 (N_3574,In_1355,N_2718);
nor U3575 (N_3575,N_2406,N_1598);
xnor U3576 (N_3576,In_3498,N_3424);
or U3577 (N_3577,N_3092,In_3921);
nor U3578 (N_3578,N_3068,N_1241);
and U3579 (N_3579,N_2279,N_2785);
xor U3580 (N_3580,N_443,N_3175);
or U3581 (N_3581,N_3168,N_3099);
nor U3582 (N_3582,N_556,N_3427);
or U3583 (N_3583,In_4315,N_258);
xnor U3584 (N_3584,N_3123,N_1990);
and U3585 (N_3585,N_3196,N_3098);
xor U3586 (N_3586,In_4757,N_2631);
nor U3587 (N_3587,In_2551,N_3402);
or U3588 (N_3588,N_3236,N_3276);
nor U3589 (N_3589,In_4209,N_3114);
and U3590 (N_3590,N_3381,N_3416);
and U3591 (N_3591,N_2756,N_2396);
or U3592 (N_3592,In_2469,N_3215);
nor U3593 (N_3593,N_3462,N_1787);
xor U3594 (N_3594,In_2120,N_3239);
and U3595 (N_3595,N_3067,N_2106);
and U3596 (N_3596,N_1364,In_103);
and U3597 (N_3597,N_3496,N_2969);
or U3598 (N_3598,N_3272,N_2362);
and U3599 (N_3599,N_2838,In_3590);
nor U3600 (N_3600,N_2997,N_2089);
xor U3601 (N_3601,In_974,N_3310);
nand U3602 (N_3602,N_1220,N_3295);
or U3603 (N_3603,N_3252,N_2606);
or U3604 (N_3604,N_1272,N_2871);
nor U3605 (N_3605,In_4115,N_2800);
and U3606 (N_3606,In_110,N_703);
nand U3607 (N_3607,In_4395,In_4546);
nand U3608 (N_3608,N_2687,N_3415);
xor U3609 (N_3609,N_2771,N_3326);
xnor U3610 (N_3610,N_2717,In_1669);
nor U3611 (N_3611,In_641,N_3063);
nand U3612 (N_3612,N_2773,In_4254);
and U3613 (N_3613,N_2935,N_3120);
nor U3614 (N_3614,In_994,N_2843);
and U3615 (N_3615,N_2977,N_2552);
nor U3616 (N_3616,N_1744,N_3036);
and U3617 (N_3617,In_3662,N_3084);
xnor U3618 (N_3618,N_2874,N_3493);
or U3619 (N_3619,N_2832,N_1396);
nand U3620 (N_3620,In_17,N_888);
nand U3621 (N_3621,N_3187,In_160);
xor U3622 (N_3622,N_3137,N_3027);
and U3623 (N_3623,N_3074,In_1534);
nand U3624 (N_3624,N_1795,In_2876);
xor U3625 (N_3625,In_4907,N_2063);
xnor U3626 (N_3626,In_1714,In_346);
and U3627 (N_3627,N_3154,N_2507);
nand U3628 (N_3628,In_2948,N_3048);
nand U3629 (N_3629,N_3471,N_3087);
xnor U3630 (N_3630,N_3185,In_2557);
nor U3631 (N_3631,N_1161,N_2831);
nand U3632 (N_3632,N_3369,N_3472);
nor U3633 (N_3633,N_3173,N_2501);
or U3634 (N_3634,N_3396,N_3118);
xnor U3635 (N_3635,In_1581,N_301);
or U3636 (N_3636,N_3062,N_2545);
xor U3637 (N_3637,N_2950,N_3230);
nand U3638 (N_3638,N_1860,In_28);
and U3639 (N_3639,N_2663,N_3391);
nand U3640 (N_3640,N_2357,N_3296);
or U3641 (N_3641,N_2941,N_1417);
and U3642 (N_3642,In_461,N_2132);
or U3643 (N_3643,N_3025,N_3204);
or U3644 (N_3644,N_3274,N_3193);
nor U3645 (N_3645,N_1981,In_3488);
nor U3646 (N_3646,In_443,N_3290);
xnor U3647 (N_3647,In_3924,N_3308);
xnor U3648 (N_3648,In_1252,N_3127);
nand U3649 (N_3649,N_3380,N_2961);
nand U3650 (N_3650,In_3394,N_3393);
nor U3651 (N_3651,N_743,N_2690);
and U3652 (N_3652,N_2951,N_3004);
nor U3653 (N_3653,N_2540,N_3282);
xnor U3654 (N_3654,N_2420,N_3201);
nor U3655 (N_3655,N_2189,In_3646);
or U3656 (N_3656,N_3216,N_1561);
xnor U3657 (N_3657,N_3489,N_2964);
xnor U3658 (N_3658,N_2809,N_2436);
nand U3659 (N_3659,N_3332,N_1527);
and U3660 (N_3660,N_2940,N_3263);
nor U3661 (N_3661,N_1051,N_3377);
nor U3662 (N_3662,N_3261,N_3008);
nor U3663 (N_3663,N_3420,N_3269);
xor U3664 (N_3664,N_3135,N_2573);
nor U3665 (N_3665,N_3119,N_2716);
and U3666 (N_3666,N_2084,N_2693);
xor U3667 (N_3667,N_3468,N_1359);
or U3668 (N_3668,In_2025,N_3029);
and U3669 (N_3669,N_1680,N_3264);
xnor U3670 (N_3670,N_2355,N_2584);
xnor U3671 (N_3671,In_113,N_3304);
nor U3672 (N_3672,N_3438,In_405);
or U3673 (N_3673,N_3246,N_111);
xnor U3674 (N_3674,N_2862,In_1503);
nor U3675 (N_3675,In_3049,N_2272);
xnor U3676 (N_3676,N_1110,In_911);
xnor U3677 (N_3677,N_1719,N_1145);
or U3678 (N_3678,N_2790,N_2555);
and U3679 (N_3679,In_3018,N_1714);
nand U3680 (N_3680,In_2098,N_2551);
nand U3681 (N_3681,In_468,N_3315);
nand U3682 (N_3682,In_2829,N_3355);
and U3683 (N_3683,N_2215,N_1279);
xor U3684 (N_3684,N_1597,N_2466);
nor U3685 (N_3685,N_3335,N_3161);
or U3686 (N_3686,N_2041,N_2880);
nand U3687 (N_3687,N_1839,N_3426);
xnor U3688 (N_3688,N_3233,In_2561);
nand U3689 (N_3689,N_2703,N_755);
xor U3690 (N_3690,N_2714,N_2520);
nor U3691 (N_3691,N_1584,In_2498);
or U3692 (N_3692,N_3324,N_3108);
nand U3693 (N_3693,N_2754,In_527);
and U3694 (N_3694,N_1713,N_1442);
nand U3695 (N_3695,N_3058,N_2624);
nor U3696 (N_3696,N_261,N_2314);
or U3697 (N_3697,N_2778,N_1803);
or U3698 (N_3698,N_3217,In_4074);
and U3699 (N_3699,In_2153,N_3132);
xor U3700 (N_3700,N_2966,N_2082);
or U3701 (N_3701,N_3488,N_3423);
nor U3702 (N_3702,In_1895,N_3117);
or U3703 (N_3703,N_3197,In_297);
and U3704 (N_3704,N_2366,N_3400);
and U3705 (N_3705,N_1457,N_2705);
nor U3706 (N_3706,N_3495,In_1125);
nor U3707 (N_3707,N_2273,In_3522);
and U3708 (N_3708,N_2429,N_3406);
nor U3709 (N_3709,N_1493,N_3080);
and U3710 (N_3710,In_1134,N_3401);
or U3711 (N_3711,N_2982,N_2865);
nor U3712 (N_3712,N_3268,N_2710);
nand U3713 (N_3713,N_1107,N_3449);
and U3714 (N_3714,N_2218,In_2195);
nor U3715 (N_3715,N_3163,N_3445);
nand U3716 (N_3716,N_2250,N_585);
xor U3717 (N_3717,N_3294,N_2592);
or U3718 (N_3718,N_2600,N_3234);
nor U3719 (N_3719,N_2452,N_2478);
xor U3720 (N_3720,In_4162,N_218);
nor U3721 (N_3721,In_3939,N_2594);
xor U3722 (N_3722,In_2257,N_2730);
nor U3723 (N_3723,N_1036,N_2724);
xnor U3724 (N_3724,N_2956,N_3078);
nor U3725 (N_3725,N_3021,N_2158);
nand U3726 (N_3726,N_2284,N_3407);
and U3727 (N_3727,In_3669,N_1974);
nand U3728 (N_3728,N_1475,N_2863);
nor U3729 (N_3729,In_3794,In_2262);
xnor U3730 (N_3730,N_3384,N_2746);
xor U3731 (N_3731,N_3146,N_2699);
xnor U3732 (N_3732,N_3309,In_3583);
nor U3733 (N_3733,N_2787,N_1897);
nand U3734 (N_3734,In_3229,N_3247);
xor U3735 (N_3735,N_2854,N_2912);
nor U3736 (N_3736,N_2389,N_3020);
xor U3737 (N_3737,N_3237,N_3102);
xor U3738 (N_3738,N_2031,N_2137);
or U3739 (N_3739,N_633,N_3260);
nand U3740 (N_3740,In_2607,N_2572);
nor U3741 (N_3741,In_1739,N_3066);
xnor U3742 (N_3742,In_2594,N_3208);
xor U3743 (N_3743,In_4849,N_3050);
nand U3744 (N_3744,In_4890,N_3041);
nand U3745 (N_3745,N_3411,N_3136);
and U3746 (N_3746,In_3402,N_1171);
xnor U3747 (N_3747,N_2737,N_2561);
xor U3748 (N_3748,N_2834,N_1938);
or U3749 (N_3749,N_3443,N_2467);
nor U3750 (N_3750,N_2441,N_2256);
nor U3751 (N_3751,In_797,In_3354);
or U3752 (N_3752,In_4652,N_1802);
nor U3753 (N_3753,N_3113,N_1270);
or U3754 (N_3754,In_2021,In_3228);
xor U3755 (N_3755,N_2462,In_3124);
nand U3756 (N_3756,N_3035,N_1574);
and U3757 (N_3757,N_3006,In_1427);
and U3758 (N_3758,In_1104,N_2547);
nor U3759 (N_3759,In_3436,N_3244);
nand U3760 (N_3760,N_2796,N_390);
nor U3761 (N_3761,N_2840,N_2475);
nor U3762 (N_3762,N_2571,N_2811);
nand U3763 (N_3763,N_1845,N_3176);
nor U3764 (N_3764,N_915,N_3280);
or U3765 (N_3765,In_1416,In_456);
xnor U3766 (N_3766,N_3318,In_2884);
nor U3767 (N_3767,In_1215,N_2965);
or U3768 (N_3768,N_1328,N_3364);
or U3769 (N_3769,N_2819,In_1746);
and U3770 (N_3770,In_316,In_883);
xnor U3771 (N_3771,N_3459,In_1672);
nand U3772 (N_3772,N_2719,N_2989);
or U3773 (N_3773,In_82,N_1495);
xor U3774 (N_3774,N_3142,N_3356);
nor U3775 (N_3775,N_3386,In_4280);
nand U3776 (N_3776,In_179,N_3271);
or U3777 (N_3777,N_2172,N_2443);
xnor U3778 (N_3778,N_1736,N_3436);
nor U3779 (N_3779,N_3378,N_3405);
or U3780 (N_3780,In_783,N_3052);
and U3781 (N_3781,N_3343,In_3503);
nor U3782 (N_3782,In_2272,N_2738);
or U3783 (N_3783,N_1287,N_3334);
or U3784 (N_3784,N_160,In_1477);
nor U3785 (N_3785,In_700,N_3016);
and U3786 (N_3786,In_3189,N_2344);
xor U3787 (N_3787,N_1569,N_1617);
nand U3788 (N_3788,N_3352,In_1424);
or U3789 (N_3789,N_745,In_2544);
or U3790 (N_3790,N_3316,In_396);
and U3791 (N_3791,N_1934,In_267);
xnor U3792 (N_3792,N_2430,N_1853);
nand U3793 (N_3793,N_2513,In_4219);
nand U3794 (N_3794,N_735,N_1411);
or U3795 (N_3795,In_4459,N_3177);
and U3796 (N_3796,N_1777,N_3055);
xnor U3797 (N_3797,N_1709,In_2979);
nand U3798 (N_3798,N_3394,N_2408);
and U3799 (N_3799,N_3228,N_623);
nor U3800 (N_3800,N_34,N_3075);
or U3801 (N_3801,In_2891,N_3241);
nand U3802 (N_3802,N_3198,N_3174);
and U3803 (N_3803,N_2704,N_3227);
and U3804 (N_3804,N_3284,N_1492);
and U3805 (N_3805,N_2529,N_1898);
nor U3806 (N_3806,In_1000,N_3181);
xor U3807 (N_3807,N_2799,N_2987);
or U3808 (N_3808,N_2889,N_1277);
nor U3809 (N_3809,N_3141,N_2316);
nor U3810 (N_3810,N_3336,N_500);
xor U3811 (N_3811,N_3253,N_3285);
nand U3812 (N_3812,N_1940,N_1733);
xnor U3813 (N_3813,N_3147,In_3842);
or U3814 (N_3814,In_1801,N_2685);
or U3815 (N_3815,N_3487,N_1943);
nand U3816 (N_3816,In_52,N_3270);
xnor U3817 (N_3817,In_3392,N_288);
xor U3818 (N_3818,In_4730,N_885);
or U3819 (N_3819,In_3982,In_3611);
xnor U3820 (N_3820,In_3694,N_840);
xnor U3821 (N_3821,N_1987,In_4985);
nand U3822 (N_3822,N_2689,N_3434);
nand U3823 (N_3823,N_3069,N_2432);
nand U3824 (N_3824,In_4049,N_2590);
nand U3825 (N_3825,N_1429,N_2691);
and U3826 (N_3826,In_3506,N_2991);
or U3827 (N_3827,N_1423,N_3238);
and U3828 (N_3828,In_488,N_3143);
xor U3829 (N_3829,N_3022,N_3034);
xnor U3830 (N_3830,N_2407,In_3987);
nand U3831 (N_3831,In_1360,N_3115);
or U3832 (N_3832,N_3028,N_729);
nand U3833 (N_3833,N_1371,N_3446);
nand U3834 (N_3834,N_481,N_3456);
and U3835 (N_3835,N_1018,N_1612);
xor U3836 (N_3836,N_1716,In_746);
nand U3837 (N_3837,N_1955,N_214);
xor U3838 (N_3838,N_3414,N_3417);
or U3839 (N_3839,N_2622,N_2916);
nand U3840 (N_3840,N_2205,N_3444);
and U3841 (N_3841,N_1376,N_3323);
and U3842 (N_3842,N_3385,In_1694);
nand U3843 (N_3843,N_3003,N_3093);
or U3844 (N_3844,N_2769,N_3278);
nor U3845 (N_3845,In_4987,N_979);
xor U3846 (N_3846,N_338,N_3045);
nand U3847 (N_3847,N_2875,N_2116);
nand U3848 (N_3848,N_3205,In_4765);
xor U3849 (N_3849,N_2788,In_299);
or U3850 (N_3850,N_3189,N_2453);
nand U3851 (N_3851,N_419,In_3641);
nand U3852 (N_3852,N_3365,In_1353);
nor U3853 (N_3853,N_3116,N_3071);
nand U3854 (N_3854,N_209,In_1326);
and U3855 (N_3855,N_3124,N_2913);
nor U3856 (N_3856,In_4800,N_3422);
or U3857 (N_3857,N_1799,In_4964);
nor U3858 (N_3858,N_2903,N_2275);
nor U3859 (N_3859,N_2855,In_1141);
xnor U3860 (N_3860,N_3015,N_3251);
xnor U3861 (N_3861,In_3067,N_1805);
and U3862 (N_3862,N_2242,N_1164);
xnor U3863 (N_3863,N_2566,In_2910);
xnor U3864 (N_3864,N_414,N_1953);
nand U3865 (N_3865,N_2338,N_1377);
or U3866 (N_3866,N_3413,N_2413);
xnor U3867 (N_3867,N_3460,N_1163);
xnor U3868 (N_3868,In_2739,N_2861);
nor U3869 (N_3869,N_2104,N_2517);
nand U3870 (N_3870,N_2206,N_2887);
nand U3871 (N_3871,N_3257,N_2294);
and U3872 (N_3872,N_3301,N_2568);
xnor U3873 (N_3873,N_3383,In_4470);
nor U3874 (N_3874,N_2904,N_2656);
nand U3875 (N_3875,N_2736,In_2472);
nor U3876 (N_3876,N_2542,N_3109);
nand U3877 (N_3877,N_2434,N_843);
nor U3878 (N_3878,In_3221,N_2667);
xnor U3879 (N_3879,N_2159,N_3457);
xor U3880 (N_3880,N_2249,In_3588);
and U3881 (N_3881,N_2144,In_2463);
nand U3882 (N_3882,N_3397,N_2258);
or U3883 (N_3883,N_3345,N_1947);
nand U3884 (N_3884,In_2977,N_3464);
or U3885 (N_3885,N_2676,N_2850);
and U3886 (N_3886,In_2909,N_2245);
nor U3887 (N_3887,N_1907,N_225);
nor U3888 (N_3888,N_3321,N_3293);
and U3889 (N_3889,N_2345,N_3180);
xor U3890 (N_3890,N_2891,N_1841);
xnor U3891 (N_3891,N_2292,In_4236);
nor U3892 (N_3892,In_1264,N_2943);
and U3893 (N_3893,N_3103,N_3485);
xor U3894 (N_3894,N_15,N_2367);
xnor U3895 (N_3895,N_2728,N_3395);
xor U3896 (N_3896,N_3473,N_2818);
nor U3897 (N_3897,In_3081,N_2556);
nand U3898 (N_3898,N_3349,N_2939);
xor U3899 (N_3899,In_39,N_3100);
and U3900 (N_3900,N_3060,N_3277);
nand U3901 (N_3901,N_2502,N_2439);
and U3902 (N_3902,N_3319,N_3011);
xor U3903 (N_3903,N_3484,N_2753);
nand U3904 (N_3904,N_3299,In_491);
or U3905 (N_3905,N_1563,N_2914);
nand U3906 (N_3906,N_3267,N_2936);
or U3907 (N_3907,N_2516,N_2643);
nand U3908 (N_3908,In_4477,In_2585);
xnor U3909 (N_3909,N_972,N_3059);
or U3910 (N_3910,In_2111,N_3089);
and U3911 (N_3911,N_1449,N_2814);
nand U3912 (N_3912,N_3017,In_1177);
or U3913 (N_3913,In_4429,In_4833);
and U3914 (N_3914,In_2791,N_2774);
or U3915 (N_3915,N_3104,N_3101);
and U3916 (N_3916,N_2648,In_1960);
nor U3917 (N_3917,N_1967,In_3808);
nand U3918 (N_3918,N_777,N_2593);
nor U3919 (N_3919,N_3331,N_1465);
or U3920 (N_3920,N_3085,N_3486);
and U3921 (N_3921,N_953,N_3072);
nor U3922 (N_3922,N_2077,In_3636);
or U3923 (N_3923,N_1301,N_3038);
or U3924 (N_3924,N_2750,N_2695);
xnor U3925 (N_3925,In_981,N_1997);
nor U3926 (N_3926,N_2911,In_1438);
xnor U3927 (N_3927,N_3064,N_3195);
or U3928 (N_3928,N_1865,N_1957);
nand U3929 (N_3929,N_902,N_1130);
nor U3930 (N_3930,N_3130,N_2905);
nand U3931 (N_3931,N_3398,N_3191);
and U3932 (N_3932,N_3000,N_3418);
nor U3933 (N_3933,N_2770,In_543);
or U3934 (N_3934,In_2401,N_3128);
nand U3935 (N_3935,N_64,In_1717);
or U3936 (N_3936,N_542,N_2359);
nor U3937 (N_3937,N_2893,In_386);
nor U3938 (N_3938,N_3079,N_3030);
or U3939 (N_3939,N_1468,N_2544);
and U3940 (N_3940,N_2878,N_2910);
nor U3941 (N_3941,N_3338,N_3353);
and U3942 (N_3942,N_2527,In_1844);
or U3943 (N_3943,In_4109,In_2122);
or U3944 (N_3944,N_2680,N_3357);
or U3945 (N_3945,N_3474,N_1252);
xnor U3946 (N_3946,N_2301,N_3390);
or U3947 (N_3947,N_2826,N_3095);
nand U3948 (N_3948,N_2760,In_1965);
nand U3949 (N_3949,N_2427,N_2604);
nor U3950 (N_3950,N_2635,In_4242);
nor U3951 (N_3951,N_3458,N_3432);
or U3952 (N_3952,In_263,In_2326);
and U3953 (N_3953,In_3153,N_3266);
nand U3954 (N_3954,In_1553,N_2122);
or U3955 (N_3955,N_2201,N_3286);
nor U3956 (N_3956,N_2949,N_3351);
nand U3957 (N_3957,N_1224,N_2583);
nand U3958 (N_3958,In_3527,N_3186);
nand U3959 (N_3959,N_3240,N_2318);
or U3960 (N_3960,N_1621,N_3077);
nor U3961 (N_3961,N_3306,N_2574);
nand U3962 (N_3962,N_3363,N_2640);
xor U3963 (N_3963,N_2901,In_2359);
and U3964 (N_3964,N_3155,N_3322);
nand U3965 (N_3965,N_3148,N_1896);
and U3966 (N_3966,N_83,N_3371);
and U3967 (N_3967,N_3480,N_2610);
nor U3968 (N_3968,In_1376,N_3009);
or U3969 (N_3969,N_1052,N_1508);
and U3970 (N_3970,N_2849,N_3051);
and U3971 (N_3971,N_2377,N_2732);
or U3972 (N_3972,In_228,In_1836);
or U3973 (N_3973,N_3454,In_2497);
and U3974 (N_3974,N_3231,N_2560);
or U3975 (N_3975,N_3151,N_3479);
nor U3976 (N_3976,In_1078,N_3007);
xnor U3977 (N_3977,N_1678,N_2974);
xnor U3978 (N_3978,N_1817,N_3491);
nand U3979 (N_3979,N_2138,In_1310);
and U3980 (N_3980,N_2081,N_3107);
and U3981 (N_3981,N_1632,N_2830);
and U3982 (N_3982,N_3232,N_3481);
or U3983 (N_3983,In_4616,N_3256);
nor U3984 (N_3984,In_4441,N_2382);
xnor U3985 (N_3985,N_3291,N_3337);
and U3986 (N_3986,N_464,N_1996);
nand U3987 (N_3987,N_2978,N_2265);
xor U3988 (N_3988,N_3061,N_2534);
nand U3989 (N_3989,N_3475,N_2111);
and U3990 (N_3990,N_1510,N_3346);
nor U3991 (N_3991,N_3388,N_1672);
nand U3992 (N_3992,N_3213,N_2379);
xnor U3993 (N_3993,N_2923,N_2902);
xor U3994 (N_3994,N_2694,N_2731);
or U3995 (N_3995,N_2020,In_2886);
nand U3996 (N_3996,In_302,N_317);
and U3997 (N_3997,N_2927,N_3329);
or U3998 (N_3998,N_2777,N_2550);
xnor U3999 (N_3999,N_3297,N_2768);
xnor U4000 (N_4000,N_3817,In_1084);
or U4001 (N_4001,N_3659,N_1033);
nor U4002 (N_4002,N_3724,N_3552);
and U4003 (N_4003,N_3235,N_3670);
and U4004 (N_4004,In_2591,N_3262);
nand U4005 (N_4005,N_2823,N_3421);
nor U4006 (N_4006,N_3584,N_3412);
xnor U4007 (N_4007,N_3854,In_3147);
and U4008 (N_4008,N_3005,N_3134);
xor U4009 (N_4009,In_4404,N_3769);
nand U4010 (N_4010,N_3797,N_3654);
or U4011 (N_4011,In_2846,N_2291);
and U4012 (N_4012,N_3718,N_3706);
nand U4013 (N_4013,N_3070,N_3634);
nand U4014 (N_4014,N_2364,N_3839);
or U4015 (N_4015,N_3523,N_3746);
and U4016 (N_4016,N_3957,N_3937);
xor U4017 (N_4017,N_3647,N_3538);
or U4018 (N_4018,N_3627,In_45);
xor U4019 (N_4019,N_3643,N_3997);
or U4020 (N_4020,In_3679,N_2712);
and U4021 (N_4021,N_3856,N_3713);
or U4022 (N_4022,N_1557,N_3806);
xnor U4023 (N_4023,N_3980,N_3861);
nor U4024 (N_4024,N_3556,N_2269);
and U4025 (N_4025,N_3049,N_3292);
and U4026 (N_4026,N_3790,N_3212);
xor U4027 (N_4027,N_2886,N_3599);
xor U4028 (N_4028,N_3681,In_3995);
nand U4029 (N_4029,N_3809,N_960);
nand U4030 (N_4030,N_3023,N_2307);
or U4031 (N_4031,N_3663,N_3638);
nor U4032 (N_4032,N_3249,N_3732);
or U4033 (N_4033,N_1193,N_3620);
nand U4034 (N_4034,In_1166,N_3852);
and U4035 (N_4035,N_2339,N_3695);
xnor U4036 (N_4036,N_784,N_3339);
or U4037 (N_4037,N_2333,N_3767);
nand U4038 (N_4038,N_1699,In_4740);
or U4039 (N_4039,N_3625,In_3635);
nor U4040 (N_4040,N_3152,N_3209);
and U4041 (N_4041,N_3086,N_3094);
nor U4042 (N_4042,N_195,In_3000);
and U4043 (N_4043,N_3841,N_3886);
xnor U4044 (N_4044,N_3974,N_3577);
nand U4045 (N_4045,N_3037,N_2264);
and U4046 (N_4046,N_3558,N_1819);
and U4047 (N_4047,N_3788,N_3637);
xor U4048 (N_4048,N_1239,N_3404);
xnor U4049 (N_4049,N_2890,N_3529);
nor U4050 (N_4050,N_3735,In_4012);
nand U4051 (N_4051,In_4567,N_2347);
xor U4052 (N_4052,N_3618,N_2722);
and U4053 (N_4053,N_3614,In_1498);
xnor U4054 (N_4054,N_3830,N_3860);
or U4055 (N_4055,N_3948,N_3988);
xnor U4056 (N_4056,N_3761,N_3571);
nand U4057 (N_4057,N_3636,N_3279);
nand U4058 (N_4058,N_3044,N_3952);
nor U4059 (N_4059,N_3891,N_3676);
xor U4060 (N_4060,N_3824,N_3705);
nand U4061 (N_4061,N_2254,N_3557);
and U4062 (N_4062,N_2906,N_2884);
xnor U4063 (N_4063,N_3684,N_3725);
xor U4064 (N_4064,N_3573,N_1053);
nand U4065 (N_4065,N_3626,N_3702);
xnor U4066 (N_4066,N_3379,N_3953);
or U4067 (N_4067,N_3799,N_232);
and U4068 (N_4068,N_3943,N_3375);
or U4069 (N_4069,N_3190,N_3900);
nand U4070 (N_4070,N_3553,N_908);
nand U4071 (N_4071,N_3991,N_2802);
nand U4072 (N_4072,N_3916,N_3590);
nor U4073 (N_4073,N_3540,N_2493);
or U4074 (N_4074,N_3574,N_3091);
nand U4075 (N_4075,N_2999,N_2963);
nor U4076 (N_4076,N_3470,N_603);
xnor U4077 (N_4077,N_3170,N_3924);
xnor U4078 (N_4078,N_3978,N_3831);
nor U4079 (N_4079,N_2962,N_3815);
and U4080 (N_4080,N_3609,N_3660);
xor U4081 (N_4081,N_1197,N_2960);
or U4082 (N_4082,N_3655,N_3619);
nor U4083 (N_4083,N_2276,N_3275);
nand U4084 (N_4084,N_3877,N_3907);
or U4085 (N_4085,N_3979,N_3728);
nand U4086 (N_4086,In_1507,N_3782);
or U4087 (N_4087,N_3621,N_3169);
nand U4088 (N_4088,N_3179,N_3845);
or U4089 (N_4089,N_3754,N_3740);
and U4090 (N_4090,N_3804,N_3938);
or U4091 (N_4091,N_2881,N_3358);
or U4092 (N_4092,N_3539,In_3295);
or U4093 (N_4093,In_4285,N_3184);
and U4094 (N_4094,N_2526,In_3985);
or U4095 (N_4095,N_3835,N_3823);
or U4096 (N_4096,N_3834,N_3367);
and U4097 (N_4097,N_2846,N_1852);
and U4098 (N_4098,N_3441,In_1816);
and U4099 (N_4099,N_3199,N_3640);
or U4100 (N_4100,N_3697,N_2274);
and U4101 (N_4101,N_3598,N_3776);
nor U4102 (N_4102,N_3903,N_3993);
xnor U4103 (N_4103,N_3930,N_3850);
and U4104 (N_4104,In_391,N_2743);
nand U4105 (N_4105,N_3842,N_3942);
or U4106 (N_4106,N_529,N_3921);
xnor U4107 (N_4107,N_3774,N_3905);
and U4108 (N_4108,N_3666,In_2175);
xor U4109 (N_4109,N_3884,N_3354);
xor U4110 (N_4110,N_3046,N_1303);
and U4111 (N_4111,N_3958,In_705);
xor U4112 (N_4112,N_3165,N_3816);
nor U4113 (N_4113,In_1239,N_3734);
nor U4114 (N_4114,N_2234,N_1927);
nor U4115 (N_4115,N_3500,N_1207);
nand U4116 (N_4116,N_3989,In_2606);
xnor U4117 (N_4117,N_3999,N_3675);
and U4118 (N_4118,N_3673,N_3596);
or U4119 (N_4119,N_2655,N_3910);
or U4120 (N_4120,N_3723,In_3707);
nand U4121 (N_4121,N_3088,N_3727);
nor U4122 (N_4122,N_3514,In_621);
xnor U4123 (N_4123,N_2305,N_3001);
xnor U4124 (N_4124,N_3455,N_3581);
and U4125 (N_4125,N_3631,N_2661);
nor U4126 (N_4126,N_3126,N_3887);
or U4127 (N_4127,N_3853,N_1989);
xor U4128 (N_4128,N_3987,N_3778);
xor U4129 (N_4129,N_2634,N_3273);
nand U4130 (N_4130,N_690,N_3469);
xor U4131 (N_4131,N_169,N_3671);
xnor U4132 (N_4132,N_3503,N_3373);
nor U4133 (N_4133,N_3182,N_3755);
or U4134 (N_4134,N_3701,N_3158);
or U4135 (N_4135,N_3642,N_3014);
xor U4136 (N_4136,N_3564,N_1604);
and U4137 (N_4137,In_4918,N_3328);
and U4138 (N_4138,N_3786,N_3977);
nor U4139 (N_4139,N_3635,N_3868);
or U4140 (N_4140,N_3433,N_3255);
nor U4141 (N_4141,N_3661,N_3898);
nand U4142 (N_4142,N_2148,N_3623);
nand U4143 (N_4143,N_3569,N_3054);
and U4144 (N_4144,N_3359,N_3463);
nand U4145 (N_4145,N_3606,N_3410);
xnor U4146 (N_4146,N_3646,N_3465);
or U4147 (N_4147,N_3690,N_3779);
or U4148 (N_4148,In_2306,N_3603);
nor U4149 (N_4149,N_3305,N_2539);
and U4150 (N_4150,N_3934,N_3720);
or U4151 (N_4151,N_3982,N_2532);
and U4152 (N_4152,N_2909,N_3314);
and U4153 (N_4153,N_2043,N_3530);
nor U4154 (N_4154,In_2459,N_1618);
and U4155 (N_4155,N_869,N_3832);
or U4156 (N_4156,N_2047,N_2485);
or U4157 (N_4157,N_2052,N_3327);
xor U4158 (N_4158,N_3644,In_3319);
xor U4159 (N_4159,N_3846,N_3795);
nor U4160 (N_4160,N_3829,N_3111);
nand U4161 (N_4161,N_1132,N_3857);
nand U4162 (N_4162,N_2328,N_3851);
nor U4163 (N_4163,N_3976,N_3990);
and U4164 (N_4164,N_2337,N_3229);
nand U4165 (N_4165,N_3885,N_3372);
nor U4166 (N_4166,N_3664,N_3704);
nand U4167 (N_4167,N_3909,In_4824);
and U4168 (N_4168,N_3750,N_3696);
or U4169 (N_4169,N_3531,N_3139);
nor U4170 (N_4170,N_3032,N_3737);
or U4171 (N_4171,N_2841,N_3753);
nor U4172 (N_4172,N_3825,N_3225);
and U4173 (N_4173,N_3768,N_3448);
nor U4174 (N_4174,N_3936,N_1072);
or U4175 (N_4175,N_3466,N_3546);
or U4176 (N_4176,N_2937,N_3519);
and U4177 (N_4177,N_3366,N_3652);
or U4178 (N_4178,N_3879,N_2010);
or U4179 (N_4179,In_4500,N_3726);
nor U4180 (N_4180,N_1340,In_3797);
xor U4181 (N_4181,N_3721,N_3781);
or U4182 (N_4182,N_3616,N_3419);
xnor U4183 (N_4183,In_3293,N_3019);
nand U4184 (N_4184,N_3447,N_2707);
nor U4185 (N_4185,N_3954,N_3320);
nor U4186 (N_4186,N_1954,N_3583);
nor U4187 (N_4187,N_3298,N_3712);
xor U4188 (N_4188,N_1607,N_3535);
or U4189 (N_4189,N_2512,N_3862);
or U4190 (N_4190,N_3742,N_1902);
nand U4191 (N_4191,N_1609,N_3747);
or U4192 (N_4192,N_3812,N_1600);
or U4193 (N_4193,In_2538,In_4329);
or U4194 (N_4194,N_3505,N_2353);
or U4195 (N_4195,N_3167,N_3528);
nand U4196 (N_4196,N_3065,N_1735);
nand U4197 (N_4197,In_3683,N_3789);
nand U4198 (N_4198,N_3586,N_3785);
nor U4199 (N_4199,N_3194,N_3951);
nand U4200 (N_4200,N_3729,N_3949);
or U4201 (N_4201,N_1783,In_3576);
nand U4202 (N_4202,N_3694,N_3875);
nor U4203 (N_4203,N_3855,N_3506);
xor U4204 (N_4204,N_1992,In_2689);
nand U4205 (N_4205,N_331,N_3513);
xor U4206 (N_4206,N_3922,N_2947);
or U4207 (N_4207,N_3250,N_3883);
nor U4208 (N_4208,In_3316,N_3504);
or U4209 (N_4209,N_3555,N_2858);
xnor U4210 (N_4210,N_3478,N_1788);
nand U4211 (N_4211,N_3764,N_2650);
or U4212 (N_4212,N_3521,N_3919);
or U4213 (N_4213,N_3870,N_250);
nand U4214 (N_4214,N_3524,N_3150);
nor U4215 (N_4215,In_4906,N_1568);
nand U4216 (N_4216,N_3844,In_4608);
nor U4217 (N_4217,N_1397,N_2836);
nor U4218 (N_4218,N_3218,N_3926);
or U4219 (N_4219,N_3683,N_3047);
nand U4220 (N_4220,N_3517,N_3657);
and U4221 (N_4221,N_1227,N_3986);
and U4222 (N_4222,N_3730,N_3490);
nor U4223 (N_4223,N_3752,N_3882);
xor U4224 (N_4224,N_2032,N_3617);
xor U4225 (N_4225,N_3341,N_3956);
xnor U4226 (N_4226,N_3733,N_3362);
nor U4227 (N_4227,N_3214,N_3933);
nand U4228 (N_4228,N_3669,N_3672);
xor U4229 (N_4229,N_3710,N_3711);
nor U4230 (N_4230,N_3689,N_3863);
and U4231 (N_4231,N_3840,N_3983);
nor U4232 (N_4232,N_3431,N_2332);
or U4233 (N_4233,N_3892,In_4547);
or U4234 (N_4234,N_3549,N_3607);
and U4235 (N_4235,N_3762,N_1214);
or U4236 (N_4236,N_2169,N_3827);
or U4237 (N_4237,N_3476,N_3902);
nand U4238 (N_4238,N_3962,N_3914);
xnor U4239 (N_4239,N_3222,N_3203);
or U4240 (N_4240,N_3807,N_1486);
or U4241 (N_4241,N_3656,N_3698);
nor U4242 (N_4242,N_1602,N_3076);
or U4243 (N_4243,N_3805,N_80);
or U4244 (N_4244,N_3801,N_1393);
nor U4245 (N_4245,In_1949,N_3699);
nor U4246 (N_4246,N_3533,N_3012);
nand U4247 (N_4247,N_2698,N_3551);
nand U4248 (N_4248,N_3439,N_286);
or U4249 (N_4249,N_3739,N_47);
and U4250 (N_4250,N_3794,N_3591);
or U4251 (N_4251,In_1145,N_3133);
and U4252 (N_4252,N_3867,N_3796);
xnor U4253 (N_4253,N_3678,In_328);
nand U4254 (N_4254,N_3527,N_3950);
nand U4255 (N_4255,N_3687,N_3594);
nor U4256 (N_4256,N_2559,N_3881);
nand U4257 (N_4257,N_2895,N_2954);
nand U4258 (N_4258,N_3512,N_3330);
or U4259 (N_4259,N_3945,N_1542);
nor U4260 (N_4260,In_2335,N_3450);
nor U4261 (N_4261,N_3348,N_2558);
and U4262 (N_4262,N_3518,N_3595);
nor U4263 (N_4263,In_4775,N_2623);
or U4264 (N_4264,N_2926,N_3878);
and U4265 (N_4265,N_3668,N_3716);
or U4266 (N_4266,N_3145,N_3243);
nor U4267 (N_4267,N_3685,In_1745);
nand U4268 (N_4268,N_3544,N_2859);
and U4269 (N_4269,N_3649,N_3639);
and U4270 (N_4270,In_131,N_3561);
xnor U4271 (N_4271,N_3917,N_3961);
and U4272 (N_4272,N_1914,N_3923);
xor U4273 (N_4273,N_3053,N_3947);
and U4274 (N_4274,N_3880,N_3893);
or U4275 (N_4275,N_2100,N_3927);
or U4276 (N_4276,N_592,In_4891);
or U4277 (N_4277,N_360,N_1437);
xor U4278 (N_4278,N_2177,N_3691);
xor U4279 (N_4279,N_3370,In_87);
or U4280 (N_4280,N_2976,N_3254);
nor U4281 (N_4281,N_3650,N_1434);
nor U4282 (N_4282,N_3492,N_3073);
nand U4283 (N_4283,In_668,N_3002);
or U4284 (N_4284,N_440,N_3188);
xor U4285 (N_4285,N_2040,N_3570);
or U4286 (N_4286,In_452,N_2644);
xor U4287 (N_4287,N_3865,N_2135);
nor U4288 (N_4288,N_1594,N_1924);
nor U4289 (N_4289,N_3876,N_3382);
and U4290 (N_4290,N_3939,N_3248);
xor U4291 (N_4291,N_3602,N_3822);
nor U4292 (N_4292,N_3925,N_3722);
and U4293 (N_4293,In_606,N_3708);
nand U4294 (N_4294,N_3566,N_3688);
and U4295 (N_4295,N_3995,N_2114);
or U4296 (N_4296,N_3994,N_2334);
xnor U4297 (N_4297,In_3702,N_3667);
nand U4298 (N_4298,N_3568,N_3901);
nor U4299 (N_4299,N_3206,N_3559);
nand U4300 (N_4300,N_2779,N_3580);
or U4301 (N_4301,N_2715,N_2589);
nand U4302 (N_4302,N_3759,N_3766);
nor U4303 (N_4303,N_3680,N_3913);
or U4304 (N_4304,N_435,N_3800);
nor U4305 (N_4305,N_2204,N_2346);
nand U4306 (N_4306,N_3615,N_2749);
or U4307 (N_4307,N_3935,N_2219);
or U4308 (N_4308,N_2758,N_3112);
nand U4309 (N_4309,N_3965,N_2599);
and U4310 (N_4310,N_3849,N_3259);
and U4311 (N_4311,N_3033,N_3542);
nor U4312 (N_4312,In_4210,N_3105);
nor U4313 (N_4313,N_2117,N_1782);
xnor U4314 (N_4314,In_4047,N_3946);
and U4315 (N_4315,N_3547,N_3818);
or U4316 (N_4316,N_3200,N_3918);
nand U4317 (N_4317,N_3763,N_3562);
or U4318 (N_4318,N_3964,In_4055);
nand U4319 (N_4319,N_2742,N_2582);
or U4320 (N_4320,N_2666,In_3927);
xnor U4321 (N_4321,N_3645,N_3792);
xnor U4322 (N_4322,N_3632,N_3097);
nand U4323 (N_4323,In_4364,N_3090);
nor U4324 (N_4324,In_1446,N_3920);
and U4325 (N_4325,In_1235,N_3604);
and U4326 (N_4326,N_560,N_3289);
or U4327 (N_4327,In_325,N_3915);
nand U4328 (N_4328,N_3453,In_526);
or U4329 (N_4329,N_2431,N_3871);
nand U4330 (N_4330,N_3904,N_1194);
or U4331 (N_4331,N_3541,In_1763);
xor U4332 (N_4332,N_3281,N_3745);
or U4333 (N_4333,In_3157,N_3311);
and U4334 (N_4334,N_3748,N_3658);
nor U4335 (N_4335,N_3931,N_2459);
xnor U4336 (N_4336,N_2677,N_2326);
and U4337 (N_4337,N_3811,In_605);
nand U4338 (N_4338,N_642,N_3554);
nor U4339 (N_4339,N_3437,N_2793);
and U4340 (N_4340,N_2735,In_992);
or U4341 (N_4341,N_2907,In_4613);
or U4342 (N_4342,N_3010,N_3821);
nor U4343 (N_4343,N_3848,N_3941);
nand U4344 (N_4344,N_3828,N_772);
nor U4345 (N_4345,N_3837,N_3802);
nand U4346 (N_4346,N_3743,N_3633);
xnor U4347 (N_4347,N_3888,N_1844);
and U4348 (N_4348,N_3313,N_3674);
or U4349 (N_4349,N_2928,N_3803);
or U4350 (N_4350,N_3808,N_3731);
or U4351 (N_4351,N_2817,N_3543);
or U4352 (N_4352,N_3972,N_2888);
nor U4353 (N_4353,N_2822,N_3361);
nor U4354 (N_4354,N_3287,N_3996);
xor U4355 (N_4355,In_15,N_2449);
xor U4356 (N_4356,N_2702,N_3350);
nor U4357 (N_4357,N_3928,N_2967);
xnor U4358 (N_4358,N_3403,N_3611);
xnor U4359 (N_4359,N_3219,N_1430);
nor U4360 (N_4360,N_2072,N_3525);
nand U4361 (N_4361,N_3593,In_357);
nor U4362 (N_4362,N_3516,N_3975);
nor U4363 (N_4363,N_3897,N_3575);
and U4364 (N_4364,N_3536,N_3864);
and U4365 (N_4365,N_2857,In_4788);
nand U4366 (N_4366,In_4009,N_2311);
nand U4367 (N_4367,N_3629,N_2025);
nand U4368 (N_4368,N_3707,N_3166);
nor U4369 (N_4369,N_3428,N_3682);
and U4370 (N_4370,N_3511,In_762);
nor U4371 (N_4371,N_3520,N_3510);
or U4372 (N_4372,N_3858,N_3944);
nand U4373 (N_4373,In_1194,N_3866);
nor U4374 (N_4374,N_1571,In_257);
xnor U4375 (N_4375,N_3494,N_427);
xor U4376 (N_4376,N_3317,N_3912);
and U4377 (N_4377,N_3224,N_3969);
or U4378 (N_4378,N_3600,N_3814);
and U4379 (N_4379,N_3813,N_3451);
xnor U4380 (N_4380,N_3700,In_2208);
xnor U4381 (N_4381,N_3653,N_3765);
or U4382 (N_4382,N_3057,In_675);
xor U4383 (N_4383,N_3744,N_2747);
nor U4384 (N_4384,N_3787,N_970);
xor U4385 (N_4385,N_1096,N_3613);
and U4386 (N_4386,N_3651,N_3578);
nor U4387 (N_4387,N_3783,N_3131);
xor U4388 (N_4388,N_3758,N_3959);
and U4389 (N_4389,N_1728,N_2058);
nand U4390 (N_4390,N_3507,N_2899);
or U4391 (N_4391,N_3874,N_2748);
xor U4392 (N_4392,N_3908,In_4601);
or U4393 (N_4393,N_2519,N_3171);
nand U4394 (N_4394,N_3932,N_3610);
and U4395 (N_4395,N_1188,In_1351);
nand U4396 (N_4396,N_3172,N_67);
nand U4397 (N_4397,In_2404,N_3374);
xnor U4398 (N_4398,N_3579,N_2992);
nand U4399 (N_4399,N_3039,N_3981);
nor U4400 (N_4400,N_3890,In_1748);
nor U4401 (N_4401,N_3648,N_3501);
xnor U4402 (N_4402,N_3714,N_3741);
xnor U4403 (N_4403,N_3548,N_766);
or U4404 (N_4404,N_3192,N_3592);
or U4405 (N_4405,N_3960,In_35);
and U4406 (N_4406,N_2649,N_3056);
and U4407 (N_4407,N_1614,N_3360);
and U4408 (N_4408,N_3894,N_3677);
and U4409 (N_4409,N_3288,N_3408);
and U4410 (N_4410,N_3971,N_2984);
and U4411 (N_4411,N_3307,N_2518);
or U4412 (N_4412,N_3265,N_3164);
xor U4413 (N_4413,N_3026,N_2979);
nand U4414 (N_4414,N_3777,N_3826);
and U4415 (N_4415,N_3911,N_3340);
xnor U4416 (N_4416,N_3376,N_966);
nand U4417 (N_4417,N_3770,N_2086);
or U4418 (N_4418,N_3899,N_3509);
xnor U4419 (N_4419,N_3153,N_2619);
nor U4420 (N_4420,N_3122,N_2801);
and U4421 (N_4421,N_2829,N_2554);
xor U4422 (N_4422,N_3873,N_3283);
or U4423 (N_4423,N_3565,N_3798);
and U4424 (N_4424,N_2970,N_3502);
and U4425 (N_4425,N_3601,N_3140);
nor U4426 (N_4426,N_3889,N_3833);
nand U4427 (N_4427,N_3587,N_997);
or U4428 (N_4428,N_3757,N_3693);
xor U4429 (N_4429,N_3628,N_3031);
xnor U4430 (N_4430,N_2340,N_3738);
nor U4431 (N_4431,N_2343,N_3968);
nor U4432 (N_4432,In_2155,N_3775);
xnor U4433 (N_4433,In_2875,N_3793);
xor U4434 (N_4434,N_3780,N_3082);
nor U4435 (N_4435,N_3482,N_3368);
nand U4436 (N_4436,N_3756,N_3872);
nor U4437 (N_4437,N_3709,N_3622);
nand U4438 (N_4438,N_2673,N_3869);
or U4439 (N_4439,N_3605,N_3970);
or U4440 (N_4440,N_3630,N_3483);
nand U4441 (N_4441,N_3522,N_3773);
xnor U4442 (N_4442,N_3749,N_3772);
nand U4443 (N_4443,N_2948,N_3896);
and U4444 (N_4444,In_3109,N_3537);
xnor U4445 (N_4445,N_3545,N_3563);
and U4446 (N_4446,N_3906,In_4044);
nor U4447 (N_4447,N_3771,N_3819);
nor U4448 (N_4448,N_3955,N_2681);
xnor U4449 (N_4449,N_3662,In_3615);
or U4450 (N_4450,N_847,N_3992);
or U4451 (N_4451,N_3585,N_3534);
nand U4452 (N_4452,N_3515,N_3966);
nand U4453 (N_4453,N_2479,In_4033);
and U4454 (N_4454,N_3589,N_3612);
nor U4455 (N_4455,N_3588,N_2515);
nor U4456 (N_4456,N_3838,N_2042);
or U4457 (N_4457,N_3719,N_3984);
xor U4458 (N_4458,N_1378,N_3608);
and U4459 (N_4459,N_3736,N_3895);
nor U4460 (N_4460,In_3523,In_3466);
nor U4461 (N_4461,In_4928,N_3560);
nor U4462 (N_4462,In_699,N_1662);
nor U4463 (N_4463,In_1277,N_3440);
nand U4464 (N_4464,N_3144,N_3973);
nor U4465 (N_4465,N_3110,N_3162);
xor U4466 (N_4466,N_1213,N_2525);
nand U4467 (N_4467,N_3679,N_3159);
nand U4468 (N_4468,N_3791,N_3760);
or U4469 (N_4469,N_3576,N_3985);
nor U4470 (N_4470,N_2797,N_986);
xnor U4471 (N_4471,N_3717,N_2585);
nand U4472 (N_4472,In_1012,N_3784);
nor U4473 (N_4473,N_3810,N_2323);
nor U4474 (N_4474,N_2896,N_3859);
nor U4475 (N_4475,N_3183,N_3582);
or U4476 (N_4476,N_3024,N_3597);
or U4477 (N_4477,In_3555,N_3641);
nor U4478 (N_4478,N_1760,In_3407);
xor U4479 (N_4479,N_1623,N_3692);
xor U4480 (N_4480,N_2833,N_3963);
xor U4481 (N_4481,N_3665,N_3929);
xor U4482 (N_4482,N_3508,N_3550);
nor U4483 (N_4483,N_3572,N_3715);
xor U4484 (N_4484,In_1677,N_3751);
or U4485 (N_4485,In_965,N_3258);
nor U4486 (N_4486,N_3843,N_2741);
and U4487 (N_4487,N_3467,N_3178);
and U4488 (N_4488,N_1189,N_3567);
or U4489 (N_4489,N_3820,N_3686);
nor U4490 (N_4490,N_3526,N_1936);
or U4491 (N_4491,N_3532,N_2668);
and U4492 (N_4492,N_2368,N_3847);
nor U4493 (N_4493,N_2146,N_1564);
nand U4494 (N_4494,In_544,N_2652);
or U4495 (N_4495,N_3836,N_1114);
nor U4496 (N_4496,N_3125,N_2664);
xnor U4497 (N_4497,N_3940,N_3998);
and U4498 (N_4498,N_3624,N_3967);
nor U4499 (N_4499,N_3703,In_1167);
nor U4500 (N_4500,N_4148,N_4146);
nor U4501 (N_4501,N_4153,N_4415);
xor U4502 (N_4502,N_4094,N_4380);
nor U4503 (N_4503,N_4149,N_4121);
nor U4504 (N_4504,N_4004,N_4416);
nor U4505 (N_4505,N_4308,N_4221);
or U4506 (N_4506,N_4155,N_4126);
nor U4507 (N_4507,N_4186,N_4250);
nand U4508 (N_4508,N_4453,N_4367);
and U4509 (N_4509,N_4434,N_4396);
and U4510 (N_4510,N_4257,N_4074);
nor U4511 (N_4511,N_4339,N_4409);
nor U4512 (N_4512,N_4400,N_4029);
or U4513 (N_4513,N_4129,N_4353);
or U4514 (N_4514,N_4338,N_4133);
nand U4515 (N_4515,N_4337,N_4097);
xor U4516 (N_4516,N_4328,N_4332);
and U4517 (N_4517,N_4152,N_4194);
or U4518 (N_4518,N_4203,N_4124);
nor U4519 (N_4519,N_4267,N_4058);
xnor U4520 (N_4520,N_4189,N_4408);
and U4521 (N_4521,N_4410,N_4006);
and U4522 (N_4522,N_4040,N_4031);
nand U4523 (N_4523,N_4011,N_4106);
nand U4524 (N_4524,N_4301,N_4002);
xor U4525 (N_4525,N_4278,N_4484);
nor U4526 (N_4526,N_4254,N_4212);
nand U4527 (N_4527,N_4333,N_4336);
nor U4528 (N_4528,N_4405,N_4024);
and U4529 (N_4529,N_4340,N_4314);
nor U4530 (N_4530,N_4205,N_4362);
and U4531 (N_4531,N_4447,N_4052);
nor U4532 (N_4532,N_4320,N_4306);
nand U4533 (N_4533,N_4023,N_4483);
or U4534 (N_4534,N_4335,N_4185);
nor U4535 (N_4535,N_4385,N_4169);
nand U4536 (N_4536,N_4035,N_4219);
xnor U4537 (N_4537,N_4007,N_4230);
nor U4538 (N_4538,N_4099,N_4240);
nand U4539 (N_4539,N_4251,N_4083);
nor U4540 (N_4540,N_4210,N_4113);
nand U4541 (N_4541,N_4281,N_4142);
nor U4542 (N_4542,N_4411,N_4261);
nand U4543 (N_4543,N_4160,N_4324);
nor U4544 (N_4544,N_4275,N_4310);
nor U4545 (N_4545,N_4218,N_4063);
and U4546 (N_4546,N_4119,N_4343);
or U4547 (N_4547,N_4444,N_4055);
xor U4548 (N_4548,N_4065,N_4036);
or U4549 (N_4549,N_4430,N_4199);
xnor U4550 (N_4550,N_4322,N_4132);
or U4551 (N_4551,N_4445,N_4319);
nand U4552 (N_4552,N_4228,N_4491);
and U4553 (N_4553,N_4192,N_4485);
and U4554 (N_4554,N_4443,N_4073);
and U4555 (N_4555,N_4118,N_4349);
nand U4556 (N_4556,N_4307,N_4276);
and U4557 (N_4557,N_4158,N_4469);
nand U4558 (N_4558,N_4436,N_4022);
or U4559 (N_4559,N_4026,N_4348);
and U4560 (N_4560,N_4499,N_4493);
xor U4561 (N_4561,N_4216,N_4127);
nand U4562 (N_4562,N_4034,N_4141);
and U4563 (N_4563,N_4432,N_4401);
and U4564 (N_4564,N_4008,N_4331);
and U4565 (N_4565,N_4012,N_4171);
or U4566 (N_4566,N_4048,N_4390);
nor U4567 (N_4567,N_4170,N_4180);
and U4568 (N_4568,N_4070,N_4242);
xnor U4569 (N_4569,N_4360,N_4435);
and U4570 (N_4570,N_4454,N_4027);
xnor U4571 (N_4571,N_4406,N_4449);
nor U4572 (N_4572,N_4093,N_4279);
xnor U4573 (N_4573,N_4128,N_4223);
and U4574 (N_4574,N_4222,N_4032);
or U4575 (N_4575,N_4477,N_4196);
nor U4576 (N_4576,N_4269,N_4176);
and U4577 (N_4577,N_4000,N_4259);
nor U4578 (N_4578,N_4235,N_4159);
xnor U4579 (N_4579,N_4120,N_4174);
nor U4580 (N_4580,N_4283,N_4496);
or U4581 (N_4581,N_4231,N_4418);
xor U4582 (N_4582,N_4164,N_4138);
and U4583 (N_4583,N_4371,N_4227);
nor U4584 (N_4584,N_4383,N_4042);
or U4585 (N_4585,N_4086,N_4249);
and U4586 (N_4586,N_4071,N_4238);
or U4587 (N_4587,N_4078,N_4393);
xor U4588 (N_4588,N_4253,N_4271);
or U4589 (N_4589,N_4107,N_4274);
nand U4590 (N_4590,N_4357,N_4209);
and U4591 (N_4591,N_4215,N_4030);
nand U4592 (N_4592,N_4388,N_4183);
or U4593 (N_4593,N_4207,N_4244);
xnor U4594 (N_4594,N_4190,N_4243);
or U4595 (N_4595,N_4072,N_4028);
nor U4596 (N_4596,N_4168,N_4470);
xor U4597 (N_4597,N_4304,N_4287);
and U4598 (N_4598,N_4366,N_4461);
nor U4599 (N_4599,N_4116,N_4224);
nand U4600 (N_4600,N_4193,N_4211);
xnor U4601 (N_4601,N_4397,N_4019);
or U4602 (N_4602,N_4200,N_4479);
or U4603 (N_4603,N_4497,N_4090);
and U4604 (N_4604,N_4345,N_4407);
and U4605 (N_4605,N_4466,N_4041);
xor U4606 (N_4606,N_4291,N_4297);
xor U4607 (N_4607,N_4392,N_4213);
and U4608 (N_4608,N_4321,N_4471);
or U4609 (N_4609,N_4260,N_4025);
xor U4610 (N_4610,N_4423,N_4226);
nand U4611 (N_4611,N_4361,N_4359);
xnor U4612 (N_4612,N_4056,N_4151);
xnor U4613 (N_4613,N_4354,N_4412);
nor U4614 (N_4614,N_4247,N_4472);
or U4615 (N_4615,N_4474,N_4080);
nand U4616 (N_4616,N_4378,N_4398);
xor U4617 (N_4617,N_4315,N_4125);
nand U4618 (N_4618,N_4085,N_4368);
nor U4619 (N_4619,N_4233,N_4273);
or U4620 (N_4620,N_4091,N_4143);
nor U4621 (N_4621,N_4144,N_4114);
xor U4622 (N_4622,N_4054,N_4266);
or U4623 (N_4623,N_4448,N_4350);
nand U4624 (N_4624,N_4404,N_4187);
nand U4625 (N_4625,N_4014,N_4232);
nor U4626 (N_4626,N_4123,N_4122);
or U4627 (N_4627,N_4309,N_4191);
or U4628 (N_4628,N_4162,N_4492);
xor U4629 (N_4629,N_4369,N_4330);
and U4630 (N_4630,N_4312,N_4137);
nor U4631 (N_4631,N_4179,N_4280);
or U4632 (N_4632,N_4437,N_4376);
nor U4633 (N_4633,N_4341,N_4358);
nor U4634 (N_4634,N_4234,N_4285);
or U4635 (N_4635,N_4387,N_4016);
and U4636 (N_4636,N_4302,N_4165);
xor U4637 (N_4637,N_4346,N_4157);
nand U4638 (N_4638,N_4413,N_4255);
and U4639 (N_4639,N_4206,N_4356);
and U4640 (N_4640,N_4342,N_4069);
nor U4641 (N_4641,N_4105,N_4136);
or U4642 (N_4642,N_4262,N_4323);
xnor U4643 (N_4643,N_4057,N_4264);
nor U4644 (N_4644,N_4303,N_4134);
nand U4645 (N_4645,N_4139,N_4429);
and U4646 (N_4646,N_4467,N_4096);
nor U4647 (N_4647,N_4239,N_4017);
nor U4648 (N_4648,N_4427,N_4382);
xnor U4649 (N_4649,N_4064,N_4386);
or U4650 (N_4650,N_4379,N_4372);
nor U4651 (N_4651,N_4225,N_4464);
xor U4652 (N_4652,N_4050,N_4311);
and U4653 (N_4653,N_4166,N_4298);
and U4654 (N_4654,N_4403,N_4288);
and U4655 (N_4655,N_4059,N_4475);
nand U4656 (N_4656,N_4229,N_4109);
nor U4657 (N_4657,N_4439,N_4334);
and U4658 (N_4658,N_4292,N_4173);
or U4659 (N_4659,N_4363,N_4049);
or U4660 (N_4660,N_4208,N_4010);
nand U4661 (N_4661,N_4177,N_4018);
xor U4662 (N_4662,N_4381,N_4374);
nand U4663 (N_4663,N_4414,N_4438);
or U4664 (N_4664,N_4329,N_4377);
or U4665 (N_4665,N_4178,N_4263);
xor U4666 (N_4666,N_4295,N_4450);
xor U4667 (N_4667,N_4364,N_4061);
xnor U4668 (N_4668,N_4115,N_4277);
xor U4669 (N_4669,N_4431,N_4220);
xor U4670 (N_4670,N_4417,N_4294);
nand U4671 (N_4671,N_4481,N_4075);
xor U4672 (N_4672,N_4021,N_4013);
xor U4673 (N_4673,N_4131,N_4110);
nor U4674 (N_4674,N_4441,N_4480);
nor U4675 (N_4675,N_4150,N_4424);
and U4676 (N_4676,N_4163,N_4087);
or U4677 (N_4677,N_4462,N_4370);
or U4678 (N_4678,N_4038,N_4425);
nor U4679 (N_4679,N_4486,N_4317);
nor U4680 (N_4680,N_4428,N_4316);
and U4681 (N_4681,N_4422,N_4318);
xor U4682 (N_4682,N_4446,N_4062);
nor U4683 (N_4683,N_4076,N_4252);
or U4684 (N_4684,N_4457,N_4296);
and U4685 (N_4685,N_4351,N_4204);
nand U4686 (N_4686,N_4299,N_4112);
and U4687 (N_4687,N_4037,N_4108);
nor U4688 (N_4688,N_4045,N_4419);
xor U4689 (N_4689,N_4198,N_4420);
xor U4690 (N_4690,N_4305,N_4195);
xnor U4691 (N_4691,N_4033,N_4039);
nor U4692 (N_4692,N_4172,N_4102);
nand U4693 (N_4693,N_4005,N_4344);
or U4694 (N_4694,N_4015,N_4167);
or U4695 (N_4695,N_4389,N_4103);
nor U4696 (N_4696,N_4082,N_4084);
nor U4697 (N_4697,N_4079,N_4313);
nand U4698 (N_4698,N_4433,N_4268);
or U4699 (N_4699,N_4043,N_4442);
xnor U4700 (N_4700,N_4066,N_4347);
nor U4701 (N_4701,N_4001,N_4044);
nor U4702 (N_4702,N_4421,N_4375);
xor U4703 (N_4703,N_4286,N_4482);
nand U4704 (N_4704,N_4478,N_4463);
and U4705 (N_4705,N_4245,N_4009);
or U4706 (N_4706,N_4460,N_4384);
nand U4707 (N_4707,N_4217,N_4327);
nand U4708 (N_4708,N_4117,N_4440);
and U4709 (N_4709,N_4100,N_4175);
nand U4710 (N_4710,N_4325,N_4104);
nand U4711 (N_4711,N_4077,N_4053);
nand U4712 (N_4712,N_4181,N_4282);
and U4713 (N_4713,N_4156,N_4111);
xnor U4714 (N_4714,N_4394,N_4051);
nand U4715 (N_4715,N_4258,N_4293);
nor U4716 (N_4716,N_4468,N_4246);
or U4717 (N_4717,N_4399,N_4237);
xnor U4718 (N_4718,N_4202,N_4373);
or U4719 (N_4719,N_4490,N_4265);
or U4720 (N_4720,N_4489,N_4060);
and U4721 (N_4721,N_4289,N_4426);
nor U4722 (N_4722,N_4459,N_4095);
nand U4723 (N_4723,N_4081,N_4270);
nor U4724 (N_4724,N_4452,N_4465);
and U4725 (N_4725,N_4130,N_4182);
and U4726 (N_4726,N_4476,N_4197);
nand U4727 (N_4727,N_4188,N_4272);
or U4728 (N_4728,N_4147,N_4236);
or U4729 (N_4729,N_4046,N_4488);
nor U4730 (N_4730,N_4456,N_4003);
nand U4731 (N_4731,N_4092,N_4101);
nand U4732 (N_4732,N_4326,N_4047);
or U4733 (N_4733,N_4241,N_4473);
and U4734 (N_4734,N_4161,N_4391);
nand U4735 (N_4735,N_4402,N_4395);
and U4736 (N_4736,N_4067,N_4284);
and U4737 (N_4737,N_4455,N_4089);
xnor U4738 (N_4738,N_4495,N_4201);
or U4739 (N_4739,N_4088,N_4256);
and U4740 (N_4740,N_4140,N_4135);
nand U4741 (N_4741,N_4214,N_4355);
nand U4742 (N_4742,N_4020,N_4098);
or U4743 (N_4743,N_4365,N_4184);
and U4744 (N_4744,N_4300,N_4352);
nor U4745 (N_4745,N_4290,N_4154);
and U4746 (N_4746,N_4498,N_4451);
or U4747 (N_4747,N_4458,N_4068);
and U4748 (N_4748,N_4145,N_4487);
nor U4749 (N_4749,N_4248,N_4494);
or U4750 (N_4750,N_4138,N_4276);
and U4751 (N_4751,N_4254,N_4015);
nor U4752 (N_4752,N_4395,N_4239);
and U4753 (N_4753,N_4073,N_4445);
xnor U4754 (N_4754,N_4068,N_4161);
and U4755 (N_4755,N_4479,N_4259);
or U4756 (N_4756,N_4270,N_4463);
xor U4757 (N_4757,N_4220,N_4308);
xor U4758 (N_4758,N_4295,N_4363);
xnor U4759 (N_4759,N_4182,N_4280);
or U4760 (N_4760,N_4400,N_4335);
xnor U4761 (N_4761,N_4185,N_4459);
nand U4762 (N_4762,N_4432,N_4291);
xnor U4763 (N_4763,N_4353,N_4424);
nor U4764 (N_4764,N_4495,N_4492);
xor U4765 (N_4765,N_4162,N_4357);
xor U4766 (N_4766,N_4280,N_4243);
and U4767 (N_4767,N_4480,N_4364);
and U4768 (N_4768,N_4065,N_4496);
nor U4769 (N_4769,N_4462,N_4309);
and U4770 (N_4770,N_4200,N_4426);
xnor U4771 (N_4771,N_4042,N_4149);
xor U4772 (N_4772,N_4371,N_4213);
nor U4773 (N_4773,N_4153,N_4015);
and U4774 (N_4774,N_4284,N_4495);
nor U4775 (N_4775,N_4435,N_4003);
xnor U4776 (N_4776,N_4019,N_4224);
nor U4777 (N_4777,N_4484,N_4063);
and U4778 (N_4778,N_4317,N_4151);
nor U4779 (N_4779,N_4481,N_4479);
or U4780 (N_4780,N_4356,N_4161);
xor U4781 (N_4781,N_4197,N_4360);
nor U4782 (N_4782,N_4459,N_4311);
and U4783 (N_4783,N_4212,N_4040);
nor U4784 (N_4784,N_4412,N_4145);
nand U4785 (N_4785,N_4420,N_4316);
or U4786 (N_4786,N_4003,N_4252);
nand U4787 (N_4787,N_4306,N_4383);
nand U4788 (N_4788,N_4007,N_4191);
nor U4789 (N_4789,N_4084,N_4224);
or U4790 (N_4790,N_4386,N_4050);
xor U4791 (N_4791,N_4011,N_4214);
nor U4792 (N_4792,N_4211,N_4295);
xnor U4793 (N_4793,N_4228,N_4129);
and U4794 (N_4794,N_4047,N_4400);
xnor U4795 (N_4795,N_4142,N_4185);
or U4796 (N_4796,N_4265,N_4246);
and U4797 (N_4797,N_4306,N_4124);
or U4798 (N_4798,N_4313,N_4233);
and U4799 (N_4799,N_4483,N_4379);
or U4800 (N_4800,N_4477,N_4230);
and U4801 (N_4801,N_4318,N_4325);
nand U4802 (N_4802,N_4035,N_4276);
xor U4803 (N_4803,N_4059,N_4251);
nor U4804 (N_4804,N_4470,N_4110);
and U4805 (N_4805,N_4497,N_4226);
nor U4806 (N_4806,N_4251,N_4493);
or U4807 (N_4807,N_4263,N_4210);
or U4808 (N_4808,N_4165,N_4169);
xor U4809 (N_4809,N_4178,N_4217);
or U4810 (N_4810,N_4313,N_4070);
or U4811 (N_4811,N_4314,N_4400);
nor U4812 (N_4812,N_4154,N_4024);
nor U4813 (N_4813,N_4490,N_4272);
or U4814 (N_4814,N_4136,N_4178);
nor U4815 (N_4815,N_4053,N_4342);
or U4816 (N_4816,N_4432,N_4314);
nor U4817 (N_4817,N_4200,N_4173);
or U4818 (N_4818,N_4137,N_4398);
or U4819 (N_4819,N_4204,N_4214);
and U4820 (N_4820,N_4060,N_4362);
and U4821 (N_4821,N_4269,N_4298);
and U4822 (N_4822,N_4456,N_4317);
nand U4823 (N_4823,N_4191,N_4258);
xnor U4824 (N_4824,N_4340,N_4033);
nor U4825 (N_4825,N_4052,N_4156);
nor U4826 (N_4826,N_4290,N_4036);
and U4827 (N_4827,N_4003,N_4486);
xnor U4828 (N_4828,N_4367,N_4090);
and U4829 (N_4829,N_4106,N_4424);
or U4830 (N_4830,N_4414,N_4154);
or U4831 (N_4831,N_4054,N_4411);
and U4832 (N_4832,N_4093,N_4355);
or U4833 (N_4833,N_4208,N_4321);
or U4834 (N_4834,N_4075,N_4229);
xnor U4835 (N_4835,N_4369,N_4074);
xnor U4836 (N_4836,N_4110,N_4200);
nand U4837 (N_4837,N_4313,N_4314);
nand U4838 (N_4838,N_4313,N_4251);
and U4839 (N_4839,N_4186,N_4033);
or U4840 (N_4840,N_4115,N_4290);
nor U4841 (N_4841,N_4227,N_4295);
and U4842 (N_4842,N_4469,N_4437);
nand U4843 (N_4843,N_4179,N_4323);
nor U4844 (N_4844,N_4311,N_4338);
and U4845 (N_4845,N_4249,N_4434);
or U4846 (N_4846,N_4130,N_4201);
xnor U4847 (N_4847,N_4338,N_4242);
or U4848 (N_4848,N_4144,N_4308);
or U4849 (N_4849,N_4382,N_4222);
nor U4850 (N_4850,N_4151,N_4227);
or U4851 (N_4851,N_4250,N_4404);
and U4852 (N_4852,N_4230,N_4322);
or U4853 (N_4853,N_4220,N_4172);
xnor U4854 (N_4854,N_4172,N_4026);
xor U4855 (N_4855,N_4368,N_4293);
nor U4856 (N_4856,N_4425,N_4344);
or U4857 (N_4857,N_4125,N_4110);
xnor U4858 (N_4858,N_4305,N_4438);
and U4859 (N_4859,N_4401,N_4498);
or U4860 (N_4860,N_4085,N_4076);
or U4861 (N_4861,N_4384,N_4145);
or U4862 (N_4862,N_4370,N_4298);
nor U4863 (N_4863,N_4057,N_4141);
or U4864 (N_4864,N_4028,N_4271);
and U4865 (N_4865,N_4009,N_4301);
nor U4866 (N_4866,N_4030,N_4296);
xor U4867 (N_4867,N_4408,N_4164);
xor U4868 (N_4868,N_4412,N_4079);
and U4869 (N_4869,N_4126,N_4203);
xnor U4870 (N_4870,N_4154,N_4377);
nor U4871 (N_4871,N_4497,N_4083);
nor U4872 (N_4872,N_4300,N_4016);
nor U4873 (N_4873,N_4326,N_4312);
and U4874 (N_4874,N_4282,N_4273);
nor U4875 (N_4875,N_4158,N_4057);
or U4876 (N_4876,N_4327,N_4381);
nor U4877 (N_4877,N_4471,N_4285);
xor U4878 (N_4878,N_4402,N_4283);
nand U4879 (N_4879,N_4266,N_4073);
nand U4880 (N_4880,N_4312,N_4029);
nor U4881 (N_4881,N_4339,N_4475);
and U4882 (N_4882,N_4236,N_4440);
nor U4883 (N_4883,N_4007,N_4068);
nor U4884 (N_4884,N_4116,N_4373);
nand U4885 (N_4885,N_4421,N_4343);
nand U4886 (N_4886,N_4418,N_4084);
or U4887 (N_4887,N_4169,N_4213);
nand U4888 (N_4888,N_4331,N_4173);
nand U4889 (N_4889,N_4017,N_4300);
and U4890 (N_4890,N_4400,N_4404);
xnor U4891 (N_4891,N_4159,N_4304);
nand U4892 (N_4892,N_4111,N_4340);
xnor U4893 (N_4893,N_4316,N_4355);
or U4894 (N_4894,N_4164,N_4041);
nand U4895 (N_4895,N_4234,N_4327);
or U4896 (N_4896,N_4117,N_4192);
and U4897 (N_4897,N_4054,N_4031);
nor U4898 (N_4898,N_4115,N_4177);
or U4899 (N_4899,N_4497,N_4115);
or U4900 (N_4900,N_4073,N_4414);
or U4901 (N_4901,N_4190,N_4313);
nand U4902 (N_4902,N_4192,N_4405);
nor U4903 (N_4903,N_4103,N_4185);
or U4904 (N_4904,N_4317,N_4397);
nor U4905 (N_4905,N_4020,N_4131);
nand U4906 (N_4906,N_4295,N_4366);
nand U4907 (N_4907,N_4150,N_4495);
and U4908 (N_4908,N_4072,N_4432);
and U4909 (N_4909,N_4164,N_4351);
nor U4910 (N_4910,N_4327,N_4093);
or U4911 (N_4911,N_4096,N_4243);
and U4912 (N_4912,N_4137,N_4052);
nand U4913 (N_4913,N_4193,N_4342);
nor U4914 (N_4914,N_4450,N_4153);
nand U4915 (N_4915,N_4400,N_4225);
nand U4916 (N_4916,N_4382,N_4447);
or U4917 (N_4917,N_4480,N_4240);
xor U4918 (N_4918,N_4148,N_4453);
and U4919 (N_4919,N_4354,N_4284);
and U4920 (N_4920,N_4176,N_4191);
and U4921 (N_4921,N_4020,N_4222);
or U4922 (N_4922,N_4395,N_4137);
nand U4923 (N_4923,N_4428,N_4251);
nand U4924 (N_4924,N_4058,N_4393);
xnor U4925 (N_4925,N_4404,N_4226);
and U4926 (N_4926,N_4161,N_4464);
or U4927 (N_4927,N_4269,N_4062);
xnor U4928 (N_4928,N_4318,N_4470);
and U4929 (N_4929,N_4216,N_4051);
nand U4930 (N_4930,N_4035,N_4205);
nand U4931 (N_4931,N_4465,N_4389);
nand U4932 (N_4932,N_4462,N_4372);
and U4933 (N_4933,N_4402,N_4432);
and U4934 (N_4934,N_4073,N_4267);
xor U4935 (N_4935,N_4310,N_4231);
nand U4936 (N_4936,N_4153,N_4250);
xnor U4937 (N_4937,N_4015,N_4126);
xor U4938 (N_4938,N_4432,N_4373);
or U4939 (N_4939,N_4120,N_4252);
xor U4940 (N_4940,N_4182,N_4043);
and U4941 (N_4941,N_4276,N_4111);
and U4942 (N_4942,N_4256,N_4089);
xnor U4943 (N_4943,N_4336,N_4279);
nand U4944 (N_4944,N_4173,N_4156);
nor U4945 (N_4945,N_4100,N_4074);
or U4946 (N_4946,N_4450,N_4315);
nand U4947 (N_4947,N_4467,N_4072);
xnor U4948 (N_4948,N_4255,N_4435);
xor U4949 (N_4949,N_4257,N_4318);
nor U4950 (N_4950,N_4078,N_4314);
nor U4951 (N_4951,N_4481,N_4089);
nor U4952 (N_4952,N_4033,N_4176);
or U4953 (N_4953,N_4428,N_4297);
or U4954 (N_4954,N_4393,N_4296);
or U4955 (N_4955,N_4346,N_4071);
and U4956 (N_4956,N_4338,N_4134);
nand U4957 (N_4957,N_4482,N_4272);
xnor U4958 (N_4958,N_4147,N_4030);
nand U4959 (N_4959,N_4135,N_4082);
nor U4960 (N_4960,N_4147,N_4305);
nand U4961 (N_4961,N_4453,N_4153);
and U4962 (N_4962,N_4323,N_4141);
xnor U4963 (N_4963,N_4326,N_4330);
nor U4964 (N_4964,N_4241,N_4045);
and U4965 (N_4965,N_4115,N_4175);
and U4966 (N_4966,N_4286,N_4489);
nand U4967 (N_4967,N_4193,N_4234);
xnor U4968 (N_4968,N_4086,N_4147);
nor U4969 (N_4969,N_4354,N_4199);
or U4970 (N_4970,N_4460,N_4305);
or U4971 (N_4971,N_4201,N_4433);
nor U4972 (N_4972,N_4128,N_4381);
or U4973 (N_4973,N_4134,N_4077);
or U4974 (N_4974,N_4334,N_4051);
or U4975 (N_4975,N_4487,N_4370);
xnor U4976 (N_4976,N_4299,N_4032);
nand U4977 (N_4977,N_4017,N_4366);
xnor U4978 (N_4978,N_4199,N_4260);
nand U4979 (N_4979,N_4425,N_4184);
nor U4980 (N_4980,N_4278,N_4384);
nor U4981 (N_4981,N_4141,N_4015);
nand U4982 (N_4982,N_4384,N_4473);
xnor U4983 (N_4983,N_4091,N_4407);
nor U4984 (N_4984,N_4119,N_4073);
xor U4985 (N_4985,N_4295,N_4038);
xor U4986 (N_4986,N_4396,N_4475);
nand U4987 (N_4987,N_4183,N_4224);
nand U4988 (N_4988,N_4387,N_4080);
and U4989 (N_4989,N_4403,N_4113);
and U4990 (N_4990,N_4337,N_4232);
nand U4991 (N_4991,N_4087,N_4288);
or U4992 (N_4992,N_4149,N_4376);
and U4993 (N_4993,N_4395,N_4136);
xnor U4994 (N_4994,N_4139,N_4220);
xnor U4995 (N_4995,N_4204,N_4252);
nor U4996 (N_4996,N_4492,N_4076);
xnor U4997 (N_4997,N_4483,N_4193);
or U4998 (N_4998,N_4264,N_4172);
nand U4999 (N_4999,N_4490,N_4372);
or U5000 (N_5000,N_4765,N_4644);
and U5001 (N_5001,N_4978,N_4965);
or U5002 (N_5002,N_4591,N_4666);
nand U5003 (N_5003,N_4987,N_4661);
nor U5004 (N_5004,N_4599,N_4992);
and U5005 (N_5005,N_4981,N_4731);
nor U5006 (N_5006,N_4605,N_4529);
xor U5007 (N_5007,N_4640,N_4871);
xnor U5008 (N_5008,N_4789,N_4680);
and U5009 (N_5009,N_4810,N_4937);
and U5010 (N_5010,N_4690,N_4757);
and U5011 (N_5011,N_4723,N_4638);
nand U5012 (N_5012,N_4933,N_4946);
xor U5013 (N_5013,N_4645,N_4555);
xor U5014 (N_5014,N_4578,N_4925);
or U5015 (N_5015,N_4939,N_4692);
nand U5016 (N_5016,N_4567,N_4956);
and U5017 (N_5017,N_4909,N_4568);
and U5018 (N_5018,N_4853,N_4504);
or U5019 (N_5019,N_4865,N_4516);
or U5020 (N_5020,N_4560,N_4803);
nor U5021 (N_5021,N_4614,N_4807);
and U5022 (N_5022,N_4960,N_4609);
nand U5023 (N_5023,N_4740,N_4646);
xnor U5024 (N_5024,N_4603,N_4955);
nand U5025 (N_5025,N_4747,N_4660);
or U5026 (N_5026,N_4930,N_4636);
xor U5027 (N_5027,N_4677,N_4791);
nor U5028 (N_5028,N_4624,N_4940);
xnor U5029 (N_5029,N_4786,N_4727);
and U5030 (N_5030,N_4556,N_4682);
nor U5031 (N_5031,N_4641,N_4653);
nand U5032 (N_5032,N_4708,N_4797);
and U5033 (N_5033,N_4669,N_4744);
or U5034 (N_5034,N_4924,N_4974);
xor U5035 (N_5035,N_4957,N_4967);
nor U5036 (N_5036,N_4724,N_4995);
nor U5037 (N_5037,N_4730,N_4877);
xor U5038 (N_5038,N_4679,N_4558);
and U5039 (N_5039,N_4662,N_4761);
or U5040 (N_5040,N_4628,N_4647);
nand U5041 (N_5041,N_4966,N_4561);
nor U5042 (N_5042,N_4598,N_4545);
nand U5043 (N_5043,N_4948,N_4855);
or U5044 (N_5044,N_4982,N_4663);
nor U5045 (N_5045,N_4549,N_4863);
nor U5046 (N_5046,N_4854,N_4837);
nor U5047 (N_5047,N_4776,N_4952);
nor U5048 (N_5048,N_4927,N_4918);
or U5049 (N_5049,N_4583,N_4587);
and U5050 (N_5050,N_4543,N_4577);
nor U5051 (N_5051,N_4541,N_4538);
nor U5052 (N_5052,N_4537,N_4702);
xor U5053 (N_5053,N_4683,N_4906);
xor U5054 (N_5054,N_4824,N_4772);
nor U5055 (N_5055,N_4840,N_4620);
xor U5056 (N_5056,N_4608,N_4938);
xor U5057 (N_5057,N_4973,N_4695);
nor U5058 (N_5058,N_4586,N_4681);
and U5059 (N_5059,N_4832,N_4963);
xor U5060 (N_5060,N_4774,N_4536);
or U5061 (N_5061,N_4922,N_4672);
nand U5062 (N_5062,N_4751,N_4901);
and U5063 (N_5063,N_4709,N_4998);
nand U5064 (N_5064,N_4573,N_4522);
or U5065 (N_5065,N_4878,N_4932);
xor U5066 (N_5066,N_4858,N_4814);
or U5067 (N_5067,N_4782,N_4563);
xor U5068 (N_5068,N_4670,N_4613);
nor U5069 (N_5069,N_4625,N_4900);
and U5070 (N_5070,N_4535,N_4989);
xor U5071 (N_5071,N_4781,N_4633);
nand U5072 (N_5072,N_4711,N_4615);
or U5073 (N_5073,N_4651,N_4719);
or U5074 (N_5074,N_4953,N_4991);
and U5075 (N_5075,N_4593,N_4886);
and U5076 (N_5076,N_4746,N_4984);
xnor U5077 (N_5077,N_4894,N_4528);
and U5078 (N_5078,N_4508,N_4923);
xnor U5079 (N_5079,N_4795,N_4699);
nand U5080 (N_5080,N_4584,N_4562);
nand U5081 (N_5081,N_4919,N_4518);
and U5082 (N_5082,N_4696,N_4818);
or U5083 (N_5083,N_4775,N_4539);
and U5084 (N_5084,N_4852,N_4610);
and U5085 (N_5085,N_4929,N_4616);
xor U5086 (N_5086,N_4836,N_4867);
nand U5087 (N_5087,N_4705,N_4510);
nand U5088 (N_5088,N_4862,N_4700);
nor U5089 (N_5089,N_4513,N_4790);
nand U5090 (N_5090,N_4896,N_4714);
nor U5091 (N_5091,N_4564,N_4770);
and U5092 (N_5092,N_4764,N_4606);
and U5093 (N_5093,N_4860,N_4734);
nor U5094 (N_5094,N_4949,N_4511);
or U5095 (N_5095,N_4888,N_4559);
and U5096 (N_5096,N_4920,N_4542);
xor U5097 (N_5097,N_4602,N_4684);
xnor U5098 (N_5098,N_4856,N_4649);
and U5099 (N_5099,N_4656,N_4617);
or U5100 (N_5100,N_4942,N_4905);
and U5101 (N_5101,N_4926,N_4566);
xor U5102 (N_5102,N_4823,N_4597);
or U5103 (N_5103,N_4801,N_4519);
nand U5104 (N_5104,N_4704,N_4728);
nor U5105 (N_5105,N_4509,N_4703);
nor U5106 (N_5106,N_4621,N_4735);
nor U5107 (N_5107,N_4745,N_4986);
xor U5108 (N_5108,N_4749,N_4688);
or U5109 (N_5109,N_4619,N_4706);
and U5110 (N_5110,N_4712,N_4581);
nor U5111 (N_5111,N_4773,N_4943);
or U5112 (N_5112,N_4928,N_4874);
and U5113 (N_5113,N_4595,N_4622);
and U5114 (N_5114,N_4864,N_4768);
nand U5115 (N_5115,N_4691,N_4841);
nand U5116 (N_5116,N_4742,N_4861);
nand U5117 (N_5117,N_4611,N_4784);
nor U5118 (N_5118,N_4780,N_4753);
xnor U5119 (N_5119,N_4676,N_4652);
nor U5120 (N_5120,N_4501,N_4524);
or U5121 (N_5121,N_4988,N_4554);
nor U5122 (N_5122,N_4994,N_4870);
nor U5123 (N_5123,N_4551,N_4792);
nand U5124 (N_5124,N_4859,N_4582);
or U5125 (N_5125,N_4725,N_4710);
or U5126 (N_5126,N_4758,N_4884);
and U5127 (N_5127,N_4574,N_4895);
xor U5128 (N_5128,N_4547,N_4872);
nand U5129 (N_5129,N_4767,N_4607);
nor U5130 (N_5130,N_4755,N_4612);
nand U5131 (N_5131,N_4983,N_4815);
or U5132 (N_5132,N_4912,N_4594);
and U5133 (N_5133,N_4893,N_4793);
xnor U5134 (N_5134,N_4847,N_4806);
xor U5135 (N_5135,N_4826,N_4629);
xor U5136 (N_5136,N_4866,N_4515);
or U5137 (N_5137,N_4630,N_4715);
nor U5138 (N_5138,N_4701,N_4512);
nor U5139 (N_5139,N_4947,N_4544);
and U5140 (N_5140,N_4674,N_4569);
nor U5141 (N_5141,N_4717,N_4739);
and U5142 (N_5142,N_4526,N_4546);
xor U5143 (N_5143,N_4600,N_4941);
and U5144 (N_5144,N_4527,N_4990);
or U5145 (N_5145,N_4736,N_4809);
xor U5146 (N_5146,N_4525,N_4950);
nand U5147 (N_5147,N_4520,N_4650);
nand U5148 (N_5148,N_4777,N_4979);
nor U5149 (N_5149,N_4752,N_4882);
nand U5150 (N_5150,N_4601,N_4604);
nand U5151 (N_5151,N_4985,N_4643);
and U5152 (N_5152,N_4980,N_4876);
nand U5153 (N_5153,N_4763,N_4565);
nand U5154 (N_5154,N_4552,N_4548);
nand U5155 (N_5155,N_4828,N_4964);
or U5156 (N_5156,N_4917,N_4514);
nand U5157 (N_5157,N_4783,N_4869);
nand U5158 (N_5158,N_4580,N_4890);
or U5159 (N_5159,N_4500,N_4835);
and U5160 (N_5160,N_4634,N_4766);
xnor U5161 (N_5161,N_4825,N_4642);
xor U5162 (N_5162,N_4913,N_4618);
or U5163 (N_5163,N_4553,N_4827);
or U5164 (N_5164,N_4687,N_4954);
and U5165 (N_5165,N_4903,N_4842);
nor U5166 (N_5166,N_4596,N_4756);
nor U5167 (N_5167,N_4698,N_4590);
nor U5168 (N_5168,N_4899,N_4589);
xnor U5169 (N_5169,N_4833,N_4718);
nor U5170 (N_5170,N_4993,N_4729);
xnor U5171 (N_5171,N_4737,N_4532);
nand U5172 (N_5172,N_4750,N_4667);
xor U5173 (N_5173,N_4887,N_4685);
xor U5174 (N_5174,N_4557,N_4851);
and U5175 (N_5175,N_4813,N_4523);
or U5176 (N_5176,N_4713,N_4811);
nand U5177 (N_5177,N_4738,N_4846);
nor U5178 (N_5178,N_4579,N_4592);
xor U5179 (N_5179,N_4880,N_4707);
xor U5180 (N_5180,N_4969,N_4779);
and U5181 (N_5181,N_4977,N_4533);
or U5182 (N_5182,N_4848,N_4671);
xnor U5183 (N_5183,N_4654,N_4778);
and U5184 (N_5184,N_4834,N_4530);
or U5185 (N_5185,N_4534,N_4639);
or U5186 (N_5186,N_4936,N_4694);
xnor U5187 (N_5187,N_4655,N_4915);
and U5188 (N_5188,N_4972,N_4817);
and U5189 (N_5189,N_4976,N_4794);
nand U5190 (N_5190,N_4892,N_4507);
xor U5191 (N_5191,N_4506,N_4959);
xor U5192 (N_5192,N_4697,N_4741);
or U5193 (N_5193,N_4802,N_4722);
or U5194 (N_5194,N_4831,N_4799);
nor U5195 (N_5195,N_4951,N_4898);
nand U5196 (N_5196,N_4921,N_4975);
xnor U5197 (N_5197,N_4748,N_4911);
nor U5198 (N_5198,N_4648,N_4829);
and U5199 (N_5199,N_4958,N_4816);
nand U5200 (N_5200,N_4889,N_4850);
nor U5201 (N_5201,N_4849,N_4726);
and U5202 (N_5202,N_4588,N_4521);
nor U5203 (N_5203,N_4904,N_4798);
xnor U5204 (N_5204,N_4805,N_4762);
nor U5205 (N_5205,N_4868,N_4785);
xor U5206 (N_5206,N_4968,N_4830);
or U5207 (N_5207,N_4686,N_4668);
nand U5208 (N_5208,N_4787,N_4821);
and U5209 (N_5209,N_4873,N_4673);
and U5210 (N_5210,N_4843,N_4931);
nand U5211 (N_5211,N_4907,N_4845);
or U5212 (N_5212,N_4550,N_4908);
nor U5213 (N_5213,N_4885,N_4945);
and U5214 (N_5214,N_4720,N_4693);
or U5215 (N_5215,N_4769,N_4505);
and U5216 (N_5216,N_4971,N_4659);
nor U5217 (N_5217,N_4732,N_4883);
or U5218 (N_5218,N_4996,N_4503);
xor U5219 (N_5219,N_4572,N_4743);
and U5220 (N_5220,N_4678,N_4822);
nand U5221 (N_5221,N_4914,N_4576);
nand U5222 (N_5222,N_4623,N_4771);
nand U5223 (N_5223,N_4879,N_4935);
nor U5224 (N_5224,N_4800,N_4733);
or U5225 (N_5225,N_4759,N_4716);
nor U5226 (N_5226,N_4962,N_4540);
xor U5227 (N_5227,N_4570,N_4897);
xor U5228 (N_5228,N_4585,N_4631);
nor U5229 (N_5229,N_4970,N_4754);
and U5230 (N_5230,N_4916,N_4961);
xnor U5231 (N_5231,N_4788,N_4531);
xor U5232 (N_5232,N_4502,N_4571);
or U5233 (N_5233,N_4635,N_4808);
and U5234 (N_5234,N_4675,N_4839);
xor U5235 (N_5235,N_4804,N_4627);
nor U5236 (N_5236,N_4997,N_4875);
or U5237 (N_5237,N_4796,N_4881);
or U5238 (N_5238,N_4820,N_4902);
and U5239 (N_5239,N_4999,N_4689);
or U5240 (N_5240,N_4934,N_4575);
xnor U5241 (N_5241,N_4819,N_4891);
and U5242 (N_5242,N_4760,N_4838);
and U5243 (N_5243,N_4857,N_4637);
nor U5244 (N_5244,N_4721,N_4910);
or U5245 (N_5245,N_4812,N_4844);
nor U5246 (N_5246,N_4944,N_4626);
nor U5247 (N_5247,N_4665,N_4657);
nor U5248 (N_5248,N_4517,N_4664);
or U5249 (N_5249,N_4658,N_4632);
nor U5250 (N_5250,N_4703,N_4571);
or U5251 (N_5251,N_4733,N_4702);
nand U5252 (N_5252,N_4636,N_4912);
nor U5253 (N_5253,N_4674,N_4716);
nand U5254 (N_5254,N_4769,N_4897);
and U5255 (N_5255,N_4504,N_4791);
nor U5256 (N_5256,N_4858,N_4988);
xnor U5257 (N_5257,N_4664,N_4699);
xnor U5258 (N_5258,N_4565,N_4736);
nand U5259 (N_5259,N_4663,N_4971);
xor U5260 (N_5260,N_4975,N_4826);
xor U5261 (N_5261,N_4814,N_4959);
nand U5262 (N_5262,N_4963,N_4957);
and U5263 (N_5263,N_4925,N_4948);
or U5264 (N_5264,N_4636,N_4666);
and U5265 (N_5265,N_4606,N_4851);
and U5266 (N_5266,N_4789,N_4556);
xor U5267 (N_5267,N_4530,N_4765);
nor U5268 (N_5268,N_4843,N_4748);
and U5269 (N_5269,N_4683,N_4944);
and U5270 (N_5270,N_4802,N_4647);
or U5271 (N_5271,N_4871,N_4701);
nor U5272 (N_5272,N_4653,N_4771);
nor U5273 (N_5273,N_4518,N_4861);
nand U5274 (N_5274,N_4594,N_4900);
xnor U5275 (N_5275,N_4980,N_4578);
nand U5276 (N_5276,N_4693,N_4821);
and U5277 (N_5277,N_4826,N_4696);
nand U5278 (N_5278,N_4728,N_4509);
and U5279 (N_5279,N_4908,N_4768);
and U5280 (N_5280,N_4965,N_4820);
nand U5281 (N_5281,N_4582,N_4643);
nor U5282 (N_5282,N_4983,N_4526);
xnor U5283 (N_5283,N_4982,N_4909);
nand U5284 (N_5284,N_4733,N_4849);
nor U5285 (N_5285,N_4835,N_4597);
nor U5286 (N_5286,N_4547,N_4765);
xnor U5287 (N_5287,N_4572,N_4713);
xor U5288 (N_5288,N_4980,N_4831);
and U5289 (N_5289,N_4564,N_4670);
xor U5290 (N_5290,N_4579,N_4654);
or U5291 (N_5291,N_4563,N_4933);
xnor U5292 (N_5292,N_4638,N_4959);
nand U5293 (N_5293,N_4953,N_4763);
xnor U5294 (N_5294,N_4766,N_4791);
or U5295 (N_5295,N_4925,N_4585);
nand U5296 (N_5296,N_4558,N_4563);
or U5297 (N_5297,N_4857,N_4676);
xnor U5298 (N_5298,N_4890,N_4797);
or U5299 (N_5299,N_4899,N_4582);
nand U5300 (N_5300,N_4894,N_4568);
nand U5301 (N_5301,N_4956,N_4676);
xnor U5302 (N_5302,N_4597,N_4975);
or U5303 (N_5303,N_4967,N_4588);
nor U5304 (N_5304,N_4515,N_4900);
and U5305 (N_5305,N_4524,N_4946);
nor U5306 (N_5306,N_4732,N_4995);
nand U5307 (N_5307,N_4795,N_4616);
nor U5308 (N_5308,N_4965,N_4504);
nor U5309 (N_5309,N_4606,N_4819);
and U5310 (N_5310,N_4966,N_4844);
nand U5311 (N_5311,N_4888,N_4564);
or U5312 (N_5312,N_4629,N_4660);
xor U5313 (N_5313,N_4959,N_4507);
and U5314 (N_5314,N_4987,N_4602);
nor U5315 (N_5315,N_4800,N_4515);
or U5316 (N_5316,N_4513,N_4931);
xnor U5317 (N_5317,N_4626,N_4813);
nand U5318 (N_5318,N_4850,N_4535);
nand U5319 (N_5319,N_4938,N_4962);
and U5320 (N_5320,N_4803,N_4913);
nor U5321 (N_5321,N_4516,N_4869);
xor U5322 (N_5322,N_4756,N_4722);
xnor U5323 (N_5323,N_4940,N_4792);
and U5324 (N_5324,N_4619,N_4829);
xnor U5325 (N_5325,N_4515,N_4813);
and U5326 (N_5326,N_4897,N_4501);
or U5327 (N_5327,N_4762,N_4502);
nand U5328 (N_5328,N_4878,N_4508);
nor U5329 (N_5329,N_4655,N_4995);
nand U5330 (N_5330,N_4784,N_4752);
or U5331 (N_5331,N_4597,N_4832);
or U5332 (N_5332,N_4840,N_4964);
or U5333 (N_5333,N_4867,N_4630);
nor U5334 (N_5334,N_4673,N_4758);
xor U5335 (N_5335,N_4992,N_4794);
and U5336 (N_5336,N_4917,N_4692);
or U5337 (N_5337,N_4535,N_4690);
nor U5338 (N_5338,N_4610,N_4845);
xor U5339 (N_5339,N_4958,N_4880);
or U5340 (N_5340,N_4926,N_4896);
or U5341 (N_5341,N_4647,N_4505);
nor U5342 (N_5342,N_4774,N_4569);
xor U5343 (N_5343,N_4647,N_4930);
xnor U5344 (N_5344,N_4959,N_4919);
nand U5345 (N_5345,N_4797,N_4509);
nor U5346 (N_5346,N_4873,N_4807);
and U5347 (N_5347,N_4819,N_4662);
nand U5348 (N_5348,N_4580,N_4754);
nand U5349 (N_5349,N_4889,N_4976);
xnor U5350 (N_5350,N_4601,N_4507);
nor U5351 (N_5351,N_4948,N_4504);
nor U5352 (N_5352,N_4988,N_4524);
or U5353 (N_5353,N_4939,N_4956);
xnor U5354 (N_5354,N_4844,N_4736);
and U5355 (N_5355,N_4807,N_4937);
nor U5356 (N_5356,N_4542,N_4687);
and U5357 (N_5357,N_4748,N_4542);
nand U5358 (N_5358,N_4782,N_4681);
xor U5359 (N_5359,N_4736,N_4766);
nor U5360 (N_5360,N_4892,N_4999);
or U5361 (N_5361,N_4556,N_4899);
or U5362 (N_5362,N_4720,N_4819);
and U5363 (N_5363,N_4521,N_4881);
nor U5364 (N_5364,N_4916,N_4882);
nor U5365 (N_5365,N_4836,N_4930);
or U5366 (N_5366,N_4738,N_4711);
nor U5367 (N_5367,N_4508,N_4983);
nor U5368 (N_5368,N_4633,N_4888);
nand U5369 (N_5369,N_4705,N_4660);
and U5370 (N_5370,N_4781,N_4661);
or U5371 (N_5371,N_4618,N_4500);
nand U5372 (N_5372,N_4545,N_4672);
or U5373 (N_5373,N_4939,N_4950);
xor U5374 (N_5374,N_4675,N_4913);
nor U5375 (N_5375,N_4608,N_4576);
or U5376 (N_5376,N_4770,N_4776);
xnor U5377 (N_5377,N_4564,N_4842);
and U5378 (N_5378,N_4593,N_4753);
nor U5379 (N_5379,N_4563,N_4923);
xnor U5380 (N_5380,N_4654,N_4651);
and U5381 (N_5381,N_4842,N_4868);
or U5382 (N_5382,N_4762,N_4773);
and U5383 (N_5383,N_4952,N_4894);
and U5384 (N_5384,N_4992,N_4873);
nand U5385 (N_5385,N_4864,N_4745);
xor U5386 (N_5386,N_4745,N_4575);
xnor U5387 (N_5387,N_4660,N_4924);
xnor U5388 (N_5388,N_4752,N_4782);
and U5389 (N_5389,N_4898,N_4753);
nor U5390 (N_5390,N_4654,N_4549);
nor U5391 (N_5391,N_4862,N_4852);
and U5392 (N_5392,N_4829,N_4536);
or U5393 (N_5393,N_4932,N_4742);
xor U5394 (N_5394,N_4820,N_4911);
nor U5395 (N_5395,N_4763,N_4785);
nor U5396 (N_5396,N_4557,N_4883);
xor U5397 (N_5397,N_4790,N_4818);
nand U5398 (N_5398,N_4847,N_4822);
or U5399 (N_5399,N_4849,N_4921);
nand U5400 (N_5400,N_4789,N_4766);
and U5401 (N_5401,N_4583,N_4731);
nor U5402 (N_5402,N_4898,N_4676);
and U5403 (N_5403,N_4624,N_4629);
xnor U5404 (N_5404,N_4652,N_4690);
or U5405 (N_5405,N_4513,N_4847);
or U5406 (N_5406,N_4668,N_4780);
and U5407 (N_5407,N_4723,N_4621);
nor U5408 (N_5408,N_4821,N_4620);
nand U5409 (N_5409,N_4561,N_4988);
xor U5410 (N_5410,N_4758,N_4712);
nand U5411 (N_5411,N_4832,N_4770);
or U5412 (N_5412,N_4997,N_4791);
xor U5413 (N_5413,N_4976,N_4691);
or U5414 (N_5414,N_4983,N_4893);
xor U5415 (N_5415,N_4890,N_4945);
and U5416 (N_5416,N_4540,N_4855);
nand U5417 (N_5417,N_4500,N_4504);
or U5418 (N_5418,N_4546,N_4724);
and U5419 (N_5419,N_4542,N_4901);
nand U5420 (N_5420,N_4899,N_4696);
xor U5421 (N_5421,N_4880,N_4950);
xor U5422 (N_5422,N_4715,N_4927);
nor U5423 (N_5423,N_4541,N_4572);
and U5424 (N_5424,N_4893,N_4833);
xor U5425 (N_5425,N_4655,N_4837);
or U5426 (N_5426,N_4938,N_4918);
nor U5427 (N_5427,N_4561,N_4581);
nor U5428 (N_5428,N_4542,N_4601);
or U5429 (N_5429,N_4733,N_4589);
or U5430 (N_5430,N_4857,N_4604);
and U5431 (N_5431,N_4917,N_4528);
xor U5432 (N_5432,N_4602,N_4934);
and U5433 (N_5433,N_4686,N_4824);
nand U5434 (N_5434,N_4570,N_4604);
and U5435 (N_5435,N_4723,N_4537);
xnor U5436 (N_5436,N_4593,N_4748);
or U5437 (N_5437,N_4687,N_4589);
nand U5438 (N_5438,N_4918,N_4599);
or U5439 (N_5439,N_4803,N_4723);
xor U5440 (N_5440,N_4681,N_4748);
nand U5441 (N_5441,N_4902,N_4762);
and U5442 (N_5442,N_4750,N_4870);
xnor U5443 (N_5443,N_4910,N_4507);
nor U5444 (N_5444,N_4565,N_4512);
nor U5445 (N_5445,N_4934,N_4576);
nand U5446 (N_5446,N_4655,N_4943);
xnor U5447 (N_5447,N_4805,N_4627);
or U5448 (N_5448,N_4771,N_4610);
or U5449 (N_5449,N_4561,N_4755);
and U5450 (N_5450,N_4928,N_4969);
xor U5451 (N_5451,N_4747,N_4811);
nand U5452 (N_5452,N_4992,N_4622);
and U5453 (N_5453,N_4696,N_4937);
xor U5454 (N_5454,N_4581,N_4902);
xnor U5455 (N_5455,N_4969,N_4813);
xor U5456 (N_5456,N_4922,N_4651);
or U5457 (N_5457,N_4587,N_4838);
or U5458 (N_5458,N_4637,N_4773);
xor U5459 (N_5459,N_4603,N_4662);
and U5460 (N_5460,N_4641,N_4793);
xnor U5461 (N_5461,N_4844,N_4525);
and U5462 (N_5462,N_4719,N_4712);
nand U5463 (N_5463,N_4848,N_4687);
or U5464 (N_5464,N_4846,N_4892);
or U5465 (N_5465,N_4964,N_4571);
nor U5466 (N_5466,N_4736,N_4968);
or U5467 (N_5467,N_4850,N_4823);
nand U5468 (N_5468,N_4509,N_4515);
and U5469 (N_5469,N_4502,N_4537);
nor U5470 (N_5470,N_4727,N_4749);
and U5471 (N_5471,N_4857,N_4910);
xnor U5472 (N_5472,N_4822,N_4680);
nand U5473 (N_5473,N_4847,N_4503);
nor U5474 (N_5474,N_4557,N_4705);
and U5475 (N_5475,N_4524,N_4829);
or U5476 (N_5476,N_4536,N_4660);
nor U5477 (N_5477,N_4781,N_4677);
and U5478 (N_5478,N_4904,N_4627);
nor U5479 (N_5479,N_4719,N_4855);
nor U5480 (N_5480,N_4709,N_4892);
nand U5481 (N_5481,N_4504,N_4773);
xnor U5482 (N_5482,N_4896,N_4786);
nand U5483 (N_5483,N_4526,N_4590);
and U5484 (N_5484,N_4541,N_4884);
xnor U5485 (N_5485,N_4510,N_4693);
or U5486 (N_5486,N_4683,N_4952);
xnor U5487 (N_5487,N_4680,N_4563);
or U5488 (N_5488,N_4636,N_4667);
and U5489 (N_5489,N_4890,N_4713);
nand U5490 (N_5490,N_4789,N_4977);
nor U5491 (N_5491,N_4781,N_4973);
and U5492 (N_5492,N_4673,N_4692);
xor U5493 (N_5493,N_4731,N_4834);
nand U5494 (N_5494,N_4943,N_4587);
and U5495 (N_5495,N_4635,N_4591);
and U5496 (N_5496,N_4960,N_4778);
and U5497 (N_5497,N_4563,N_4607);
and U5498 (N_5498,N_4940,N_4934);
and U5499 (N_5499,N_4705,N_4579);
xor U5500 (N_5500,N_5059,N_5319);
or U5501 (N_5501,N_5025,N_5027);
or U5502 (N_5502,N_5355,N_5109);
or U5503 (N_5503,N_5402,N_5279);
or U5504 (N_5504,N_5242,N_5167);
nand U5505 (N_5505,N_5299,N_5272);
xnor U5506 (N_5506,N_5403,N_5186);
nand U5507 (N_5507,N_5060,N_5257);
nor U5508 (N_5508,N_5039,N_5107);
nand U5509 (N_5509,N_5216,N_5359);
and U5510 (N_5510,N_5317,N_5238);
xnor U5511 (N_5511,N_5003,N_5363);
nor U5512 (N_5512,N_5233,N_5201);
xnor U5513 (N_5513,N_5061,N_5419);
or U5514 (N_5514,N_5204,N_5354);
or U5515 (N_5515,N_5410,N_5019);
xor U5516 (N_5516,N_5148,N_5118);
xnor U5517 (N_5517,N_5357,N_5176);
nand U5518 (N_5518,N_5123,N_5044);
nand U5519 (N_5519,N_5084,N_5318);
nand U5520 (N_5520,N_5348,N_5280);
and U5521 (N_5521,N_5466,N_5293);
xor U5522 (N_5522,N_5478,N_5273);
and U5523 (N_5523,N_5305,N_5188);
nand U5524 (N_5524,N_5296,N_5420);
and U5525 (N_5525,N_5268,N_5428);
nand U5526 (N_5526,N_5253,N_5200);
or U5527 (N_5527,N_5414,N_5141);
xnor U5528 (N_5528,N_5117,N_5142);
and U5529 (N_5529,N_5068,N_5065);
or U5530 (N_5530,N_5347,N_5119);
xnor U5531 (N_5531,N_5490,N_5367);
xnor U5532 (N_5532,N_5438,N_5275);
xor U5533 (N_5533,N_5245,N_5062);
xor U5534 (N_5534,N_5153,N_5447);
or U5535 (N_5535,N_5362,N_5313);
nor U5536 (N_5536,N_5470,N_5212);
and U5537 (N_5537,N_5405,N_5443);
and U5538 (N_5538,N_5106,N_5441);
xnor U5539 (N_5539,N_5444,N_5450);
xor U5540 (N_5540,N_5089,N_5194);
nor U5541 (N_5541,N_5217,N_5255);
nand U5542 (N_5542,N_5283,N_5129);
nand U5543 (N_5543,N_5240,N_5365);
xor U5544 (N_5544,N_5380,N_5012);
nand U5545 (N_5545,N_5295,N_5446);
or U5546 (N_5546,N_5404,N_5267);
xor U5547 (N_5547,N_5198,N_5050);
xor U5548 (N_5548,N_5031,N_5277);
nand U5549 (N_5549,N_5138,N_5047);
nand U5550 (N_5550,N_5029,N_5094);
or U5551 (N_5551,N_5152,N_5057);
xnor U5552 (N_5552,N_5067,N_5353);
nor U5553 (N_5553,N_5221,N_5322);
xnor U5554 (N_5554,N_5227,N_5392);
xor U5555 (N_5555,N_5485,N_5225);
nor U5556 (N_5556,N_5099,N_5092);
xor U5557 (N_5557,N_5040,N_5173);
nand U5558 (N_5558,N_5488,N_5177);
nand U5559 (N_5559,N_5157,N_5232);
xnor U5560 (N_5560,N_5372,N_5008);
nand U5561 (N_5561,N_5294,N_5151);
xor U5562 (N_5562,N_5306,N_5035);
and U5563 (N_5563,N_5407,N_5376);
xor U5564 (N_5564,N_5038,N_5475);
nand U5565 (N_5565,N_5287,N_5252);
xnor U5566 (N_5566,N_5487,N_5437);
nor U5567 (N_5567,N_5320,N_5187);
xnor U5568 (N_5568,N_5077,N_5066);
nor U5569 (N_5569,N_5457,N_5385);
nand U5570 (N_5570,N_5463,N_5199);
nand U5571 (N_5571,N_5076,N_5069);
nor U5572 (N_5572,N_5368,N_5132);
xnor U5573 (N_5573,N_5143,N_5183);
nor U5574 (N_5574,N_5274,N_5303);
nand U5575 (N_5575,N_5374,N_5366);
nand U5576 (N_5576,N_5344,N_5350);
nor U5577 (N_5577,N_5424,N_5166);
and U5578 (N_5578,N_5468,N_5458);
xnor U5579 (N_5579,N_5330,N_5467);
and U5580 (N_5580,N_5005,N_5435);
nor U5581 (N_5581,N_5377,N_5103);
nand U5582 (N_5582,N_5125,N_5228);
nand U5583 (N_5583,N_5430,N_5338);
nand U5584 (N_5584,N_5196,N_5498);
xnor U5585 (N_5585,N_5087,N_5102);
or U5586 (N_5586,N_5381,N_5191);
xnor U5587 (N_5587,N_5134,N_5053);
or U5588 (N_5588,N_5128,N_5323);
nor U5589 (N_5589,N_5270,N_5165);
or U5590 (N_5590,N_5332,N_5417);
and U5591 (N_5591,N_5496,N_5442);
nand U5592 (N_5592,N_5120,N_5286);
nand U5593 (N_5593,N_5250,N_5345);
and U5594 (N_5594,N_5006,N_5269);
and U5595 (N_5595,N_5218,N_5433);
nor U5596 (N_5596,N_5397,N_5371);
or U5597 (N_5597,N_5130,N_5247);
xor U5598 (N_5598,N_5013,N_5408);
nand U5599 (N_5599,N_5292,N_5454);
nor U5600 (N_5600,N_5336,N_5464);
and U5601 (N_5601,N_5179,N_5406);
nand U5602 (N_5602,N_5284,N_5133);
nand U5603 (N_5603,N_5030,N_5456);
or U5604 (N_5604,N_5346,N_5045);
xor U5605 (N_5605,N_5429,N_5079);
or U5606 (N_5606,N_5156,N_5291);
nor U5607 (N_5607,N_5214,N_5018);
or U5608 (N_5608,N_5314,N_5088);
and U5609 (N_5609,N_5481,N_5288);
xor U5610 (N_5610,N_5266,N_5328);
or U5611 (N_5611,N_5394,N_5469);
nor U5612 (N_5612,N_5144,N_5351);
xnor U5613 (N_5613,N_5489,N_5070);
and U5614 (N_5614,N_5097,N_5427);
and U5615 (N_5615,N_5448,N_5360);
and U5616 (N_5616,N_5304,N_5472);
nor U5617 (N_5617,N_5259,N_5459);
nor U5618 (N_5618,N_5004,N_5190);
xnor U5619 (N_5619,N_5172,N_5096);
nor U5620 (N_5620,N_5041,N_5244);
and U5621 (N_5621,N_5154,N_5193);
or U5622 (N_5622,N_5022,N_5391);
and U5623 (N_5623,N_5264,N_5393);
nor U5624 (N_5624,N_5285,N_5072);
nand U5625 (N_5625,N_5074,N_5499);
or U5626 (N_5626,N_5369,N_5197);
nor U5627 (N_5627,N_5021,N_5388);
or U5628 (N_5628,N_5423,N_5054);
xnor U5629 (N_5629,N_5418,N_5297);
nand U5630 (N_5630,N_5256,N_5220);
and U5631 (N_5631,N_5122,N_5398);
xor U5632 (N_5632,N_5055,N_5113);
or U5633 (N_5633,N_5073,N_5017);
nor U5634 (N_5634,N_5411,N_5479);
xnor U5635 (N_5635,N_5222,N_5215);
nor U5636 (N_5636,N_5101,N_5189);
xnor U5637 (N_5637,N_5327,N_5339);
and U5638 (N_5638,N_5278,N_5364);
nand U5639 (N_5639,N_5010,N_5175);
nor U5640 (N_5640,N_5178,N_5486);
or U5641 (N_5641,N_5093,N_5384);
nand U5642 (N_5642,N_5248,N_5237);
xor U5643 (N_5643,N_5356,N_5168);
nand U5644 (N_5644,N_5495,N_5263);
xor U5645 (N_5645,N_5136,N_5254);
and U5646 (N_5646,N_5145,N_5034);
and U5647 (N_5647,N_5281,N_5493);
xnor U5648 (N_5648,N_5048,N_5171);
and U5649 (N_5649,N_5321,N_5422);
or U5650 (N_5650,N_5375,N_5452);
and U5651 (N_5651,N_5207,N_5383);
nand U5652 (N_5652,N_5115,N_5108);
or U5653 (N_5653,N_5431,N_5265);
or U5654 (N_5654,N_5036,N_5230);
or U5655 (N_5655,N_5210,N_5181);
nand U5656 (N_5656,N_5311,N_5020);
xor U5657 (N_5657,N_5149,N_5140);
or U5658 (N_5658,N_5432,N_5195);
or U5659 (N_5659,N_5382,N_5016);
xnor U5660 (N_5660,N_5436,N_5460);
nand U5661 (N_5661,N_5396,N_5037);
and U5662 (N_5662,N_5370,N_5262);
and U5663 (N_5663,N_5483,N_5425);
nor U5664 (N_5664,N_5078,N_5324);
or U5665 (N_5665,N_5112,N_5023);
or U5666 (N_5666,N_5261,N_5399);
and U5667 (N_5667,N_5461,N_5491);
and U5668 (N_5668,N_5378,N_5223);
or U5669 (N_5669,N_5024,N_5104);
nor U5670 (N_5670,N_5276,N_5241);
nor U5671 (N_5671,N_5208,N_5159);
and U5672 (N_5672,N_5032,N_5180);
xnor U5673 (N_5673,N_5043,N_5471);
xnor U5674 (N_5674,N_5484,N_5494);
nand U5675 (N_5675,N_5413,N_5439);
nor U5676 (N_5676,N_5307,N_5211);
or U5677 (N_5677,N_5409,N_5352);
nor U5678 (N_5678,N_5046,N_5342);
nor U5679 (N_5679,N_5209,N_5063);
xor U5680 (N_5680,N_5337,N_5434);
and U5681 (N_5681,N_5095,N_5401);
and U5682 (N_5682,N_5476,N_5312);
xor U5683 (N_5683,N_5465,N_5110);
nor U5684 (N_5684,N_5492,N_5182);
nand U5685 (N_5685,N_5146,N_5135);
or U5686 (N_5686,N_5213,N_5289);
xnor U5687 (N_5687,N_5091,N_5086);
xnor U5688 (N_5688,N_5056,N_5049);
and U5689 (N_5689,N_5075,N_5474);
and U5690 (N_5690,N_5473,N_5235);
xnor U5691 (N_5691,N_5082,N_5373);
xor U5692 (N_5692,N_5111,N_5080);
and U5693 (N_5693,N_5386,N_5480);
nand U5694 (N_5694,N_5333,N_5329);
xor U5695 (N_5695,N_5000,N_5331);
nand U5696 (N_5696,N_5085,N_5137);
nand U5697 (N_5697,N_5349,N_5009);
or U5698 (N_5698,N_5202,N_5226);
xnor U5699 (N_5699,N_5335,N_5387);
xor U5700 (N_5700,N_5064,N_5011);
nor U5701 (N_5701,N_5033,N_5361);
nand U5702 (N_5702,N_5158,N_5246);
or U5703 (N_5703,N_5126,N_5440);
xor U5704 (N_5704,N_5083,N_5127);
and U5705 (N_5705,N_5234,N_5098);
and U5706 (N_5706,N_5379,N_5071);
nand U5707 (N_5707,N_5100,N_5162);
xor U5708 (N_5708,N_5358,N_5081);
nand U5709 (N_5709,N_5309,N_5150);
xor U5710 (N_5710,N_5497,N_5326);
nand U5711 (N_5711,N_5170,N_5028);
nand U5712 (N_5712,N_5205,N_5325);
and U5713 (N_5713,N_5026,N_5343);
nand U5714 (N_5714,N_5160,N_5139);
and U5715 (N_5715,N_5341,N_5105);
and U5716 (N_5716,N_5298,N_5300);
nand U5717 (N_5717,N_5051,N_5315);
and U5718 (N_5718,N_5426,N_5400);
xnor U5719 (N_5719,N_5453,N_5015);
nand U5720 (N_5720,N_5058,N_5114);
nand U5721 (N_5721,N_5206,N_5249);
or U5722 (N_5722,N_5412,N_5224);
xor U5723 (N_5723,N_5147,N_5121);
or U5724 (N_5724,N_5090,N_5395);
and U5725 (N_5725,N_5390,N_5302);
and U5726 (N_5726,N_5449,N_5231);
nor U5727 (N_5727,N_5184,N_5251);
or U5728 (N_5728,N_5389,N_5239);
nor U5729 (N_5729,N_5462,N_5316);
nand U5730 (N_5730,N_5334,N_5271);
and U5731 (N_5731,N_5236,N_5451);
or U5732 (N_5732,N_5174,N_5445);
and U5733 (N_5733,N_5164,N_5042);
or U5734 (N_5734,N_5124,N_5290);
or U5735 (N_5735,N_5282,N_5192);
and U5736 (N_5736,N_5421,N_5229);
and U5737 (N_5737,N_5415,N_5001);
nor U5738 (N_5738,N_5116,N_5155);
or U5739 (N_5739,N_5416,N_5052);
xor U5740 (N_5740,N_5477,N_5301);
xnor U5741 (N_5741,N_5455,N_5169);
or U5742 (N_5742,N_5002,N_5203);
nand U5743 (N_5743,N_5131,N_5258);
or U5744 (N_5744,N_5310,N_5260);
xor U5745 (N_5745,N_5482,N_5163);
or U5746 (N_5746,N_5007,N_5014);
xnor U5747 (N_5747,N_5340,N_5243);
or U5748 (N_5748,N_5161,N_5185);
and U5749 (N_5749,N_5219,N_5308);
and U5750 (N_5750,N_5033,N_5123);
nand U5751 (N_5751,N_5235,N_5435);
xnor U5752 (N_5752,N_5065,N_5135);
or U5753 (N_5753,N_5385,N_5278);
nand U5754 (N_5754,N_5082,N_5094);
nor U5755 (N_5755,N_5371,N_5047);
nor U5756 (N_5756,N_5044,N_5273);
nor U5757 (N_5757,N_5478,N_5142);
and U5758 (N_5758,N_5162,N_5169);
xnor U5759 (N_5759,N_5452,N_5303);
or U5760 (N_5760,N_5364,N_5061);
nor U5761 (N_5761,N_5135,N_5020);
nand U5762 (N_5762,N_5332,N_5274);
nand U5763 (N_5763,N_5484,N_5374);
and U5764 (N_5764,N_5426,N_5445);
nor U5765 (N_5765,N_5088,N_5396);
xor U5766 (N_5766,N_5456,N_5353);
xor U5767 (N_5767,N_5422,N_5416);
or U5768 (N_5768,N_5146,N_5116);
and U5769 (N_5769,N_5403,N_5311);
xnor U5770 (N_5770,N_5003,N_5433);
xnor U5771 (N_5771,N_5335,N_5285);
and U5772 (N_5772,N_5497,N_5147);
nor U5773 (N_5773,N_5423,N_5044);
nand U5774 (N_5774,N_5246,N_5368);
or U5775 (N_5775,N_5083,N_5080);
or U5776 (N_5776,N_5201,N_5203);
nor U5777 (N_5777,N_5226,N_5283);
nand U5778 (N_5778,N_5314,N_5398);
nand U5779 (N_5779,N_5292,N_5052);
xnor U5780 (N_5780,N_5254,N_5157);
nor U5781 (N_5781,N_5460,N_5476);
and U5782 (N_5782,N_5102,N_5376);
or U5783 (N_5783,N_5279,N_5206);
xor U5784 (N_5784,N_5379,N_5044);
or U5785 (N_5785,N_5488,N_5186);
or U5786 (N_5786,N_5449,N_5178);
nor U5787 (N_5787,N_5498,N_5375);
nor U5788 (N_5788,N_5260,N_5484);
xor U5789 (N_5789,N_5491,N_5380);
nand U5790 (N_5790,N_5407,N_5046);
and U5791 (N_5791,N_5394,N_5035);
xnor U5792 (N_5792,N_5213,N_5149);
nand U5793 (N_5793,N_5400,N_5245);
and U5794 (N_5794,N_5183,N_5291);
nand U5795 (N_5795,N_5473,N_5339);
xnor U5796 (N_5796,N_5406,N_5088);
xor U5797 (N_5797,N_5455,N_5116);
and U5798 (N_5798,N_5190,N_5238);
nand U5799 (N_5799,N_5463,N_5419);
nor U5800 (N_5800,N_5253,N_5157);
nor U5801 (N_5801,N_5271,N_5286);
and U5802 (N_5802,N_5138,N_5489);
xor U5803 (N_5803,N_5165,N_5116);
nand U5804 (N_5804,N_5369,N_5408);
or U5805 (N_5805,N_5261,N_5407);
xor U5806 (N_5806,N_5275,N_5258);
nor U5807 (N_5807,N_5045,N_5071);
and U5808 (N_5808,N_5076,N_5118);
and U5809 (N_5809,N_5061,N_5251);
nor U5810 (N_5810,N_5377,N_5039);
and U5811 (N_5811,N_5229,N_5277);
nor U5812 (N_5812,N_5347,N_5177);
xnor U5813 (N_5813,N_5267,N_5331);
or U5814 (N_5814,N_5436,N_5341);
nand U5815 (N_5815,N_5145,N_5427);
xor U5816 (N_5816,N_5048,N_5106);
nor U5817 (N_5817,N_5330,N_5260);
xnor U5818 (N_5818,N_5035,N_5110);
xor U5819 (N_5819,N_5023,N_5397);
nor U5820 (N_5820,N_5453,N_5382);
nor U5821 (N_5821,N_5379,N_5249);
nor U5822 (N_5822,N_5238,N_5203);
and U5823 (N_5823,N_5188,N_5327);
or U5824 (N_5824,N_5233,N_5354);
nor U5825 (N_5825,N_5333,N_5271);
xnor U5826 (N_5826,N_5154,N_5106);
xor U5827 (N_5827,N_5172,N_5019);
xor U5828 (N_5828,N_5042,N_5009);
and U5829 (N_5829,N_5338,N_5149);
xor U5830 (N_5830,N_5119,N_5129);
nor U5831 (N_5831,N_5122,N_5188);
and U5832 (N_5832,N_5451,N_5166);
xor U5833 (N_5833,N_5345,N_5356);
and U5834 (N_5834,N_5443,N_5073);
or U5835 (N_5835,N_5289,N_5121);
nand U5836 (N_5836,N_5485,N_5355);
xnor U5837 (N_5837,N_5418,N_5210);
nand U5838 (N_5838,N_5142,N_5139);
or U5839 (N_5839,N_5360,N_5073);
xnor U5840 (N_5840,N_5022,N_5296);
and U5841 (N_5841,N_5023,N_5448);
and U5842 (N_5842,N_5254,N_5116);
xor U5843 (N_5843,N_5312,N_5344);
nor U5844 (N_5844,N_5161,N_5029);
nand U5845 (N_5845,N_5018,N_5438);
and U5846 (N_5846,N_5145,N_5066);
or U5847 (N_5847,N_5498,N_5458);
nand U5848 (N_5848,N_5205,N_5028);
xor U5849 (N_5849,N_5338,N_5309);
xor U5850 (N_5850,N_5112,N_5240);
or U5851 (N_5851,N_5486,N_5044);
and U5852 (N_5852,N_5018,N_5228);
xnor U5853 (N_5853,N_5276,N_5321);
nor U5854 (N_5854,N_5482,N_5006);
xnor U5855 (N_5855,N_5256,N_5443);
and U5856 (N_5856,N_5230,N_5352);
and U5857 (N_5857,N_5444,N_5058);
and U5858 (N_5858,N_5447,N_5495);
and U5859 (N_5859,N_5188,N_5349);
nand U5860 (N_5860,N_5222,N_5244);
nor U5861 (N_5861,N_5027,N_5496);
nor U5862 (N_5862,N_5285,N_5010);
and U5863 (N_5863,N_5342,N_5034);
nor U5864 (N_5864,N_5232,N_5255);
or U5865 (N_5865,N_5434,N_5422);
nand U5866 (N_5866,N_5230,N_5062);
nand U5867 (N_5867,N_5349,N_5198);
xor U5868 (N_5868,N_5039,N_5465);
and U5869 (N_5869,N_5243,N_5426);
nand U5870 (N_5870,N_5121,N_5142);
and U5871 (N_5871,N_5183,N_5349);
and U5872 (N_5872,N_5139,N_5247);
or U5873 (N_5873,N_5067,N_5348);
nor U5874 (N_5874,N_5382,N_5164);
or U5875 (N_5875,N_5427,N_5484);
nor U5876 (N_5876,N_5077,N_5053);
or U5877 (N_5877,N_5055,N_5266);
or U5878 (N_5878,N_5089,N_5255);
and U5879 (N_5879,N_5384,N_5455);
and U5880 (N_5880,N_5491,N_5435);
nand U5881 (N_5881,N_5391,N_5190);
nand U5882 (N_5882,N_5259,N_5320);
nand U5883 (N_5883,N_5489,N_5139);
nor U5884 (N_5884,N_5498,N_5349);
or U5885 (N_5885,N_5406,N_5063);
and U5886 (N_5886,N_5258,N_5343);
xnor U5887 (N_5887,N_5311,N_5023);
or U5888 (N_5888,N_5329,N_5385);
or U5889 (N_5889,N_5479,N_5292);
and U5890 (N_5890,N_5437,N_5349);
nand U5891 (N_5891,N_5365,N_5065);
nand U5892 (N_5892,N_5302,N_5491);
and U5893 (N_5893,N_5451,N_5488);
nor U5894 (N_5894,N_5331,N_5112);
or U5895 (N_5895,N_5010,N_5404);
nor U5896 (N_5896,N_5310,N_5308);
and U5897 (N_5897,N_5171,N_5350);
nand U5898 (N_5898,N_5259,N_5262);
and U5899 (N_5899,N_5231,N_5024);
and U5900 (N_5900,N_5148,N_5489);
xnor U5901 (N_5901,N_5279,N_5168);
and U5902 (N_5902,N_5230,N_5279);
and U5903 (N_5903,N_5001,N_5418);
nor U5904 (N_5904,N_5482,N_5074);
and U5905 (N_5905,N_5028,N_5193);
nand U5906 (N_5906,N_5272,N_5045);
nand U5907 (N_5907,N_5352,N_5164);
or U5908 (N_5908,N_5378,N_5451);
xor U5909 (N_5909,N_5323,N_5152);
nand U5910 (N_5910,N_5024,N_5188);
or U5911 (N_5911,N_5299,N_5211);
nand U5912 (N_5912,N_5040,N_5284);
and U5913 (N_5913,N_5373,N_5476);
or U5914 (N_5914,N_5139,N_5452);
xor U5915 (N_5915,N_5074,N_5031);
and U5916 (N_5916,N_5284,N_5008);
nand U5917 (N_5917,N_5238,N_5143);
and U5918 (N_5918,N_5459,N_5209);
nor U5919 (N_5919,N_5216,N_5165);
or U5920 (N_5920,N_5146,N_5181);
or U5921 (N_5921,N_5159,N_5043);
nand U5922 (N_5922,N_5340,N_5270);
or U5923 (N_5923,N_5205,N_5419);
and U5924 (N_5924,N_5083,N_5348);
or U5925 (N_5925,N_5309,N_5448);
nor U5926 (N_5926,N_5223,N_5083);
xor U5927 (N_5927,N_5047,N_5064);
nand U5928 (N_5928,N_5143,N_5083);
or U5929 (N_5929,N_5417,N_5411);
or U5930 (N_5930,N_5354,N_5346);
or U5931 (N_5931,N_5389,N_5140);
nor U5932 (N_5932,N_5441,N_5112);
or U5933 (N_5933,N_5474,N_5122);
nand U5934 (N_5934,N_5112,N_5267);
xor U5935 (N_5935,N_5206,N_5412);
and U5936 (N_5936,N_5092,N_5100);
and U5937 (N_5937,N_5079,N_5284);
and U5938 (N_5938,N_5209,N_5480);
xor U5939 (N_5939,N_5390,N_5416);
xnor U5940 (N_5940,N_5274,N_5295);
nor U5941 (N_5941,N_5475,N_5110);
xnor U5942 (N_5942,N_5314,N_5306);
or U5943 (N_5943,N_5005,N_5303);
xor U5944 (N_5944,N_5075,N_5306);
xnor U5945 (N_5945,N_5106,N_5129);
xnor U5946 (N_5946,N_5381,N_5487);
and U5947 (N_5947,N_5302,N_5473);
and U5948 (N_5948,N_5230,N_5354);
and U5949 (N_5949,N_5174,N_5040);
and U5950 (N_5950,N_5360,N_5385);
nand U5951 (N_5951,N_5081,N_5182);
or U5952 (N_5952,N_5324,N_5224);
nor U5953 (N_5953,N_5217,N_5440);
or U5954 (N_5954,N_5251,N_5085);
xnor U5955 (N_5955,N_5149,N_5366);
and U5956 (N_5956,N_5405,N_5418);
xnor U5957 (N_5957,N_5498,N_5007);
nor U5958 (N_5958,N_5137,N_5195);
nor U5959 (N_5959,N_5111,N_5112);
nor U5960 (N_5960,N_5230,N_5276);
xnor U5961 (N_5961,N_5474,N_5257);
nand U5962 (N_5962,N_5108,N_5453);
and U5963 (N_5963,N_5424,N_5068);
and U5964 (N_5964,N_5450,N_5156);
nand U5965 (N_5965,N_5157,N_5240);
or U5966 (N_5966,N_5414,N_5473);
nor U5967 (N_5967,N_5226,N_5249);
or U5968 (N_5968,N_5354,N_5226);
xor U5969 (N_5969,N_5223,N_5474);
nand U5970 (N_5970,N_5096,N_5051);
or U5971 (N_5971,N_5469,N_5160);
xnor U5972 (N_5972,N_5155,N_5345);
and U5973 (N_5973,N_5015,N_5184);
nand U5974 (N_5974,N_5075,N_5225);
and U5975 (N_5975,N_5062,N_5077);
or U5976 (N_5976,N_5067,N_5144);
or U5977 (N_5977,N_5498,N_5074);
xnor U5978 (N_5978,N_5274,N_5306);
nor U5979 (N_5979,N_5419,N_5079);
nand U5980 (N_5980,N_5073,N_5345);
nor U5981 (N_5981,N_5123,N_5421);
xnor U5982 (N_5982,N_5195,N_5496);
xor U5983 (N_5983,N_5289,N_5149);
and U5984 (N_5984,N_5163,N_5275);
and U5985 (N_5985,N_5470,N_5414);
xnor U5986 (N_5986,N_5177,N_5305);
xor U5987 (N_5987,N_5324,N_5118);
xor U5988 (N_5988,N_5031,N_5166);
nor U5989 (N_5989,N_5387,N_5301);
and U5990 (N_5990,N_5018,N_5060);
or U5991 (N_5991,N_5263,N_5069);
and U5992 (N_5992,N_5163,N_5334);
or U5993 (N_5993,N_5486,N_5199);
xor U5994 (N_5994,N_5170,N_5307);
nor U5995 (N_5995,N_5338,N_5372);
or U5996 (N_5996,N_5300,N_5119);
nor U5997 (N_5997,N_5027,N_5029);
or U5998 (N_5998,N_5222,N_5066);
nor U5999 (N_5999,N_5054,N_5273);
nor U6000 (N_6000,N_5756,N_5765);
or U6001 (N_6001,N_5889,N_5785);
nor U6002 (N_6002,N_5755,N_5534);
and U6003 (N_6003,N_5973,N_5566);
nor U6004 (N_6004,N_5955,N_5517);
and U6005 (N_6005,N_5683,N_5853);
xor U6006 (N_6006,N_5526,N_5875);
xnor U6007 (N_6007,N_5748,N_5682);
nand U6008 (N_6008,N_5710,N_5726);
and U6009 (N_6009,N_5998,N_5565);
xor U6010 (N_6010,N_5822,N_5637);
nand U6011 (N_6011,N_5883,N_5549);
or U6012 (N_6012,N_5645,N_5747);
or U6013 (N_6013,N_5821,N_5545);
xnor U6014 (N_6014,N_5538,N_5692);
or U6015 (N_6015,N_5704,N_5974);
and U6016 (N_6016,N_5562,N_5542);
nand U6017 (N_6017,N_5612,N_5760);
xor U6018 (N_6018,N_5700,N_5994);
or U6019 (N_6019,N_5766,N_5687);
or U6020 (N_6020,N_5978,N_5712);
xor U6021 (N_6021,N_5598,N_5690);
and U6022 (N_6022,N_5739,N_5695);
or U6023 (N_6023,N_5908,N_5813);
nand U6024 (N_6024,N_5663,N_5897);
or U6025 (N_6025,N_5650,N_5820);
xor U6026 (N_6026,N_5922,N_5948);
or U6027 (N_6027,N_5595,N_5884);
and U6028 (N_6028,N_5548,N_5582);
xor U6029 (N_6029,N_5706,N_5810);
xnor U6030 (N_6030,N_5774,N_5699);
or U6031 (N_6031,N_5902,N_5641);
xor U6032 (N_6032,N_5653,N_5623);
xnor U6033 (N_6033,N_5796,N_5910);
or U6034 (N_6034,N_5749,N_5917);
nand U6035 (N_6035,N_5604,N_5950);
or U6036 (N_6036,N_5896,N_5934);
or U6037 (N_6037,N_5986,N_5969);
xnor U6038 (N_6038,N_5901,N_5512);
or U6039 (N_6039,N_5980,N_5725);
xor U6040 (N_6040,N_5947,N_5944);
xnor U6041 (N_6041,N_5721,N_5560);
nor U6042 (N_6042,N_5688,N_5793);
nand U6043 (N_6043,N_5581,N_5768);
or U6044 (N_6044,N_5823,N_5913);
and U6045 (N_6045,N_5867,N_5886);
xnor U6046 (N_6046,N_5697,N_5946);
xor U6047 (N_6047,N_5675,N_5972);
or U6048 (N_6048,N_5809,N_5784);
xor U6049 (N_6049,N_5824,N_5656);
and U6050 (N_6050,N_5628,N_5790);
and U6051 (N_6051,N_5574,N_5968);
nand U6052 (N_6052,N_5804,N_5826);
nand U6053 (N_6053,N_5646,N_5631);
nor U6054 (N_6054,N_5546,N_5516);
nand U6055 (N_6055,N_5981,N_5619);
or U6056 (N_6056,N_5964,N_5557);
nand U6057 (N_6057,N_5520,N_5838);
or U6058 (N_6058,N_5527,N_5530);
xnor U6059 (N_6059,N_5627,N_5539);
nor U6060 (N_6060,N_5958,N_5782);
nor U6061 (N_6061,N_5655,N_5939);
or U6062 (N_6062,N_5938,N_5664);
nand U6063 (N_6063,N_5554,N_5904);
xnor U6064 (N_6064,N_5919,N_5674);
and U6065 (N_6065,N_5639,N_5533);
or U6066 (N_6066,N_5965,N_5870);
and U6067 (N_6067,N_5898,N_5833);
or U6068 (N_6068,N_5957,N_5659);
nand U6069 (N_6069,N_5584,N_5605);
xnor U6070 (N_6070,N_5563,N_5709);
and U6071 (N_6071,N_5818,N_5911);
nor U6072 (N_6072,N_5795,N_5817);
nand U6073 (N_6073,N_5845,N_5960);
or U6074 (N_6074,N_5511,N_5803);
nand U6075 (N_6075,N_5601,N_5521);
nand U6076 (N_6076,N_5698,N_5703);
nor U6077 (N_6077,N_5841,N_5864);
nand U6078 (N_6078,N_5647,N_5618);
and U6079 (N_6079,N_5787,N_5761);
or U6080 (N_6080,N_5607,N_5869);
and U6081 (N_6081,N_5622,N_5816);
and U6082 (N_6082,N_5658,N_5661);
and U6083 (N_6083,N_5773,N_5966);
xnor U6084 (N_6084,N_5708,N_5814);
nand U6085 (N_6085,N_5762,N_5811);
and U6086 (N_6086,N_5844,N_5812);
nor U6087 (N_6087,N_5727,N_5942);
nand U6088 (N_6088,N_5776,N_5900);
or U6089 (N_6089,N_5862,N_5890);
nand U6090 (N_6090,N_5596,N_5586);
and U6091 (N_6091,N_5713,N_5736);
nor U6092 (N_6092,N_5610,N_5636);
and U6093 (N_6093,N_5854,N_5732);
xor U6094 (N_6094,N_5518,N_5594);
nor U6095 (N_6095,N_5903,N_5851);
or U6096 (N_6096,N_5840,N_5996);
or U6097 (N_6097,N_5734,N_5532);
nand U6098 (N_6098,N_5829,N_5731);
xor U6099 (N_6099,N_5681,N_5626);
nand U6100 (N_6100,N_5672,N_5745);
nand U6101 (N_6101,N_5744,N_5573);
and U6102 (N_6102,N_5614,N_5931);
nor U6103 (N_6103,N_5592,N_5694);
xnor U6104 (N_6104,N_5673,N_5691);
nand U6105 (N_6105,N_5769,N_5617);
and U6106 (N_6106,N_5531,N_5899);
and U6107 (N_6107,N_5717,N_5894);
xor U6108 (N_6108,N_5746,N_5997);
nor U6109 (N_6109,N_5609,N_5602);
nand U6110 (N_6110,N_5990,N_5551);
nor U6111 (N_6111,N_5666,N_5729);
xor U6112 (N_6112,N_5528,N_5797);
or U6113 (N_6113,N_5979,N_5536);
nor U6114 (N_6114,N_5615,N_5832);
and U6115 (N_6115,N_5544,N_5662);
and U6116 (N_6116,N_5550,N_5949);
and U6117 (N_6117,N_5852,N_5715);
nand U6118 (N_6118,N_5789,N_5735);
nor U6119 (N_6119,N_5847,N_5611);
nand U6120 (N_6120,N_5943,N_5783);
or U6121 (N_6121,N_5589,N_5597);
or U6122 (N_6122,N_5846,N_5501);
and U6123 (N_6123,N_5878,N_5881);
and U6124 (N_6124,N_5936,N_5696);
or U6125 (N_6125,N_5885,N_5963);
nor U6126 (N_6126,N_5874,N_5503);
and U6127 (N_6127,N_5956,N_5752);
xor U6128 (N_6128,N_5634,N_5750);
xnor U6129 (N_6129,N_5825,N_5740);
nor U6130 (N_6130,N_5665,N_5871);
or U6131 (N_6131,N_5933,N_5770);
or U6132 (N_6132,N_5831,N_5916);
and U6133 (N_6133,N_5859,N_5830);
nor U6134 (N_6134,N_5578,N_5952);
xnor U6135 (N_6135,N_5892,N_5794);
nor U6136 (N_6136,N_5834,N_5772);
xor U6137 (N_6137,N_5928,N_5590);
nor U6138 (N_6138,N_5802,N_5504);
xnor U6139 (N_6139,N_5808,N_5730);
nor U6140 (N_6140,N_5780,N_5537);
or U6141 (N_6141,N_5941,N_5977);
xor U6142 (N_6142,N_5678,N_5720);
xor U6143 (N_6143,N_5705,N_5579);
xor U6144 (N_6144,N_5571,N_5788);
xor U6145 (N_6145,N_5975,N_5751);
xnor U6146 (N_6146,N_5991,N_5724);
and U6147 (N_6147,N_5567,N_5680);
nor U6148 (N_6148,N_5951,N_5920);
xor U6149 (N_6149,N_5993,N_5856);
xor U6150 (N_6150,N_5588,N_5849);
nor U6151 (N_6151,N_5667,N_5879);
and U6152 (N_6152,N_5753,N_5985);
xor U6153 (N_6153,N_5801,N_5880);
and U6154 (N_6154,N_5988,N_5807);
nand U6155 (N_6155,N_5524,N_5621);
or U6156 (N_6156,N_5995,N_5525);
nand U6157 (N_6157,N_5791,N_5778);
xnor U6158 (N_6158,N_5953,N_5915);
and U6159 (N_6159,N_5926,N_5543);
nand U6160 (N_6160,N_5519,N_5987);
or U6161 (N_6161,N_5630,N_5918);
nor U6162 (N_6162,N_5570,N_5945);
and U6163 (N_6163,N_5764,N_5912);
nor U6164 (N_6164,N_5967,N_5932);
nand U6165 (N_6165,N_5670,N_5798);
xnor U6166 (N_6166,N_5800,N_5547);
nand U6167 (N_6167,N_5767,N_5771);
or U6168 (N_6168,N_5819,N_5921);
nand U6169 (N_6169,N_5669,N_5781);
nand U6170 (N_6170,N_5906,N_5895);
or U6171 (N_6171,N_5937,N_5608);
nor U6172 (N_6172,N_5775,N_5576);
or U6173 (N_6173,N_5792,N_5722);
xnor U6174 (N_6174,N_5686,N_5893);
xor U6175 (N_6175,N_5848,N_5599);
or U6176 (N_6176,N_5759,N_5603);
or U6177 (N_6177,N_5676,N_5552);
or U6178 (N_6178,N_5535,N_5679);
nor U6179 (N_6179,N_5643,N_5959);
and U6180 (N_6180,N_5907,N_5507);
or U6181 (N_6181,N_5587,N_5754);
nor U6182 (N_6182,N_5799,N_5559);
nor U6183 (N_6183,N_5909,N_5671);
and U6184 (N_6184,N_5860,N_5925);
or U6185 (N_6185,N_5914,N_5569);
and U6186 (N_6186,N_5591,N_5983);
and U6187 (N_6187,N_5858,N_5887);
or U6188 (N_6188,N_5649,N_5723);
or U6189 (N_6189,N_5758,N_5651);
xor U6190 (N_6190,N_5733,N_5842);
nor U6191 (N_6191,N_5868,N_5558);
and U6192 (N_6192,N_5509,N_5684);
and U6193 (N_6193,N_5583,N_5502);
and U6194 (N_6194,N_5961,N_5891);
nand U6195 (N_6195,N_5638,N_5500);
xor U6196 (N_6196,N_5989,N_5835);
xor U6197 (N_6197,N_5515,N_5743);
nor U6198 (N_6198,N_5970,N_5593);
xnor U6199 (N_6199,N_5625,N_5962);
and U6200 (N_6200,N_5866,N_5843);
and U6201 (N_6201,N_5872,N_5648);
or U6202 (N_6202,N_5992,N_5624);
xnor U6203 (N_6203,N_5742,N_5577);
and U6204 (N_6204,N_5652,N_5660);
and U6205 (N_6205,N_5836,N_5982);
nor U6206 (N_6206,N_5522,N_5865);
and U6207 (N_6207,N_5632,N_5633);
and U6208 (N_6208,N_5513,N_5640);
nand U6209 (N_6209,N_5716,N_5737);
nor U6210 (N_6210,N_5564,N_5923);
xor U6211 (N_6211,N_5523,N_5728);
nand U6212 (N_6212,N_5850,N_5620);
nand U6213 (N_6213,N_5572,N_5927);
and U6214 (N_6214,N_5935,N_5719);
and U6215 (N_6215,N_5877,N_5689);
xnor U6216 (N_6216,N_5606,N_5575);
or U6217 (N_6217,N_5616,N_5553);
or U6218 (N_6218,N_5924,N_5555);
and U6219 (N_6219,N_5757,N_5805);
xnor U6220 (N_6220,N_5685,N_5561);
nand U6221 (N_6221,N_5718,N_5613);
or U6222 (N_6222,N_5541,N_5929);
nand U6223 (N_6223,N_5635,N_5971);
xnor U6224 (N_6224,N_5815,N_5529);
nand U6225 (N_6225,N_5888,N_5828);
xnor U6226 (N_6226,N_5707,N_5693);
nor U6227 (N_6227,N_5806,N_5827);
and U6228 (N_6228,N_5642,N_5702);
nor U6229 (N_6229,N_5514,N_5657);
nand U6230 (N_6230,N_5763,N_5714);
xor U6231 (N_6231,N_5777,N_5580);
or U6232 (N_6232,N_5677,N_5940);
nor U6233 (N_6233,N_5568,N_5999);
nor U6234 (N_6234,N_5779,N_5855);
and U6235 (N_6235,N_5629,N_5861);
nor U6236 (N_6236,N_5837,N_5930);
and U6237 (N_6237,N_5644,N_5882);
nand U6238 (N_6238,N_5738,N_5508);
or U6239 (N_6239,N_5839,N_5540);
and U6240 (N_6240,N_5786,N_5863);
or U6241 (N_6241,N_5506,N_5505);
or U6242 (N_6242,N_5654,N_5741);
nor U6243 (N_6243,N_5510,N_5600);
or U6244 (N_6244,N_5585,N_5976);
nand U6245 (N_6245,N_5701,N_5668);
xnor U6246 (N_6246,N_5711,N_5954);
and U6247 (N_6247,N_5876,N_5556);
nand U6248 (N_6248,N_5984,N_5873);
or U6249 (N_6249,N_5857,N_5905);
nor U6250 (N_6250,N_5826,N_5783);
nand U6251 (N_6251,N_5973,N_5938);
and U6252 (N_6252,N_5527,N_5849);
and U6253 (N_6253,N_5603,N_5830);
nor U6254 (N_6254,N_5856,N_5534);
nand U6255 (N_6255,N_5944,N_5658);
or U6256 (N_6256,N_5893,N_5679);
nor U6257 (N_6257,N_5591,N_5692);
nand U6258 (N_6258,N_5736,N_5945);
xor U6259 (N_6259,N_5585,N_5556);
nand U6260 (N_6260,N_5646,N_5689);
nor U6261 (N_6261,N_5517,N_5619);
or U6262 (N_6262,N_5911,N_5922);
and U6263 (N_6263,N_5610,N_5945);
or U6264 (N_6264,N_5900,N_5746);
nand U6265 (N_6265,N_5663,N_5592);
and U6266 (N_6266,N_5938,N_5552);
nor U6267 (N_6267,N_5753,N_5863);
nand U6268 (N_6268,N_5924,N_5548);
or U6269 (N_6269,N_5618,N_5695);
and U6270 (N_6270,N_5541,N_5522);
nand U6271 (N_6271,N_5958,N_5956);
nor U6272 (N_6272,N_5623,N_5739);
nor U6273 (N_6273,N_5852,N_5789);
xor U6274 (N_6274,N_5562,N_5771);
and U6275 (N_6275,N_5740,N_5714);
or U6276 (N_6276,N_5839,N_5714);
or U6277 (N_6277,N_5526,N_5705);
or U6278 (N_6278,N_5959,N_5565);
or U6279 (N_6279,N_5878,N_5715);
nand U6280 (N_6280,N_5652,N_5537);
xor U6281 (N_6281,N_5844,N_5807);
or U6282 (N_6282,N_5623,N_5920);
nor U6283 (N_6283,N_5501,N_5701);
and U6284 (N_6284,N_5952,N_5800);
xor U6285 (N_6285,N_5934,N_5673);
or U6286 (N_6286,N_5930,N_5976);
xnor U6287 (N_6287,N_5762,N_5832);
xor U6288 (N_6288,N_5543,N_5751);
nand U6289 (N_6289,N_5613,N_5738);
nor U6290 (N_6290,N_5708,N_5659);
xnor U6291 (N_6291,N_5887,N_5651);
or U6292 (N_6292,N_5759,N_5645);
or U6293 (N_6293,N_5674,N_5878);
and U6294 (N_6294,N_5709,N_5622);
and U6295 (N_6295,N_5695,N_5843);
or U6296 (N_6296,N_5569,N_5959);
nor U6297 (N_6297,N_5747,N_5756);
or U6298 (N_6298,N_5716,N_5724);
or U6299 (N_6299,N_5973,N_5559);
xor U6300 (N_6300,N_5562,N_5882);
or U6301 (N_6301,N_5723,N_5745);
xor U6302 (N_6302,N_5664,N_5844);
or U6303 (N_6303,N_5669,N_5625);
and U6304 (N_6304,N_5843,N_5949);
nor U6305 (N_6305,N_5856,N_5587);
nand U6306 (N_6306,N_5796,N_5807);
xor U6307 (N_6307,N_5707,N_5588);
or U6308 (N_6308,N_5887,N_5523);
or U6309 (N_6309,N_5741,N_5536);
nor U6310 (N_6310,N_5938,N_5940);
nand U6311 (N_6311,N_5847,N_5718);
or U6312 (N_6312,N_5992,N_5863);
or U6313 (N_6313,N_5580,N_5698);
nor U6314 (N_6314,N_5982,N_5790);
nand U6315 (N_6315,N_5751,N_5611);
nor U6316 (N_6316,N_5666,N_5898);
xnor U6317 (N_6317,N_5541,N_5706);
or U6318 (N_6318,N_5629,N_5668);
nor U6319 (N_6319,N_5870,N_5989);
and U6320 (N_6320,N_5974,N_5897);
nor U6321 (N_6321,N_5542,N_5972);
nor U6322 (N_6322,N_5858,N_5542);
nor U6323 (N_6323,N_5774,N_5966);
xnor U6324 (N_6324,N_5910,N_5772);
xor U6325 (N_6325,N_5726,N_5803);
or U6326 (N_6326,N_5743,N_5683);
or U6327 (N_6327,N_5523,N_5778);
or U6328 (N_6328,N_5764,N_5748);
xor U6329 (N_6329,N_5710,N_5745);
nand U6330 (N_6330,N_5846,N_5828);
and U6331 (N_6331,N_5553,N_5896);
nand U6332 (N_6332,N_5641,N_5785);
and U6333 (N_6333,N_5606,N_5503);
xnor U6334 (N_6334,N_5942,N_5808);
xor U6335 (N_6335,N_5677,N_5836);
xor U6336 (N_6336,N_5677,N_5982);
xnor U6337 (N_6337,N_5548,N_5675);
nand U6338 (N_6338,N_5946,N_5962);
nand U6339 (N_6339,N_5849,N_5973);
nand U6340 (N_6340,N_5621,N_5876);
or U6341 (N_6341,N_5579,N_5605);
and U6342 (N_6342,N_5985,N_5789);
or U6343 (N_6343,N_5655,N_5694);
xor U6344 (N_6344,N_5752,N_5973);
or U6345 (N_6345,N_5846,N_5579);
nor U6346 (N_6346,N_5703,N_5737);
nand U6347 (N_6347,N_5686,N_5782);
nand U6348 (N_6348,N_5874,N_5551);
nor U6349 (N_6349,N_5732,N_5899);
nor U6350 (N_6350,N_5645,N_5717);
or U6351 (N_6351,N_5945,N_5582);
nand U6352 (N_6352,N_5529,N_5628);
and U6353 (N_6353,N_5986,N_5698);
nor U6354 (N_6354,N_5807,N_5537);
or U6355 (N_6355,N_5654,N_5737);
or U6356 (N_6356,N_5613,N_5520);
or U6357 (N_6357,N_5618,N_5739);
and U6358 (N_6358,N_5873,N_5857);
xor U6359 (N_6359,N_5759,N_5523);
nand U6360 (N_6360,N_5718,N_5671);
nand U6361 (N_6361,N_5997,N_5813);
xnor U6362 (N_6362,N_5951,N_5675);
xor U6363 (N_6363,N_5602,N_5769);
xnor U6364 (N_6364,N_5809,N_5965);
xor U6365 (N_6365,N_5815,N_5510);
and U6366 (N_6366,N_5919,N_5775);
xor U6367 (N_6367,N_5946,N_5584);
nand U6368 (N_6368,N_5820,N_5668);
nand U6369 (N_6369,N_5648,N_5656);
and U6370 (N_6370,N_5572,N_5719);
or U6371 (N_6371,N_5805,N_5957);
xnor U6372 (N_6372,N_5767,N_5986);
xnor U6373 (N_6373,N_5684,N_5843);
nand U6374 (N_6374,N_5821,N_5897);
nand U6375 (N_6375,N_5870,N_5945);
and U6376 (N_6376,N_5723,N_5786);
nor U6377 (N_6377,N_5930,N_5910);
and U6378 (N_6378,N_5772,N_5532);
nand U6379 (N_6379,N_5773,N_5793);
nor U6380 (N_6380,N_5969,N_5938);
or U6381 (N_6381,N_5599,N_5832);
nand U6382 (N_6382,N_5995,N_5868);
and U6383 (N_6383,N_5851,N_5702);
and U6384 (N_6384,N_5715,N_5931);
or U6385 (N_6385,N_5824,N_5567);
nand U6386 (N_6386,N_5842,N_5573);
or U6387 (N_6387,N_5936,N_5630);
or U6388 (N_6388,N_5859,N_5883);
and U6389 (N_6389,N_5678,N_5883);
nand U6390 (N_6390,N_5546,N_5686);
or U6391 (N_6391,N_5555,N_5677);
and U6392 (N_6392,N_5949,N_5678);
nand U6393 (N_6393,N_5813,N_5807);
nand U6394 (N_6394,N_5756,N_5567);
or U6395 (N_6395,N_5858,N_5917);
nor U6396 (N_6396,N_5868,N_5997);
or U6397 (N_6397,N_5702,N_5582);
xor U6398 (N_6398,N_5711,N_5864);
xnor U6399 (N_6399,N_5619,N_5720);
and U6400 (N_6400,N_5873,N_5921);
nor U6401 (N_6401,N_5698,N_5828);
xnor U6402 (N_6402,N_5900,N_5829);
xnor U6403 (N_6403,N_5776,N_5632);
xnor U6404 (N_6404,N_5873,N_5859);
nand U6405 (N_6405,N_5679,N_5799);
xnor U6406 (N_6406,N_5610,N_5774);
nor U6407 (N_6407,N_5756,N_5988);
xor U6408 (N_6408,N_5825,N_5804);
nand U6409 (N_6409,N_5993,N_5763);
nor U6410 (N_6410,N_5918,N_5749);
and U6411 (N_6411,N_5742,N_5999);
nand U6412 (N_6412,N_5765,N_5506);
or U6413 (N_6413,N_5789,N_5794);
nand U6414 (N_6414,N_5775,N_5798);
nor U6415 (N_6415,N_5644,N_5833);
nand U6416 (N_6416,N_5954,N_5732);
nor U6417 (N_6417,N_5891,N_5672);
nor U6418 (N_6418,N_5811,N_5934);
nor U6419 (N_6419,N_5782,N_5623);
and U6420 (N_6420,N_5520,N_5880);
nor U6421 (N_6421,N_5773,N_5948);
nand U6422 (N_6422,N_5770,N_5664);
xnor U6423 (N_6423,N_5550,N_5517);
nand U6424 (N_6424,N_5508,N_5990);
nand U6425 (N_6425,N_5636,N_5917);
nand U6426 (N_6426,N_5814,N_5731);
nand U6427 (N_6427,N_5907,N_5606);
nand U6428 (N_6428,N_5906,N_5989);
nand U6429 (N_6429,N_5649,N_5977);
and U6430 (N_6430,N_5776,N_5856);
nor U6431 (N_6431,N_5712,N_5552);
xnor U6432 (N_6432,N_5874,N_5889);
nor U6433 (N_6433,N_5923,N_5980);
nor U6434 (N_6434,N_5648,N_5911);
or U6435 (N_6435,N_5824,N_5955);
and U6436 (N_6436,N_5889,N_5910);
xnor U6437 (N_6437,N_5697,N_5614);
and U6438 (N_6438,N_5790,N_5871);
and U6439 (N_6439,N_5545,N_5919);
and U6440 (N_6440,N_5749,N_5751);
nand U6441 (N_6441,N_5784,N_5762);
and U6442 (N_6442,N_5895,N_5847);
xor U6443 (N_6443,N_5883,N_5944);
xor U6444 (N_6444,N_5780,N_5768);
and U6445 (N_6445,N_5966,N_5675);
or U6446 (N_6446,N_5630,N_5664);
xor U6447 (N_6447,N_5615,N_5960);
nor U6448 (N_6448,N_5756,N_5694);
nand U6449 (N_6449,N_5946,N_5680);
nand U6450 (N_6450,N_5940,N_5660);
nor U6451 (N_6451,N_5603,N_5961);
and U6452 (N_6452,N_5766,N_5550);
or U6453 (N_6453,N_5500,N_5926);
nand U6454 (N_6454,N_5686,N_5587);
nand U6455 (N_6455,N_5917,N_5593);
and U6456 (N_6456,N_5804,N_5675);
and U6457 (N_6457,N_5765,N_5923);
or U6458 (N_6458,N_5741,N_5899);
nand U6459 (N_6459,N_5854,N_5662);
and U6460 (N_6460,N_5928,N_5569);
nor U6461 (N_6461,N_5552,N_5948);
xnor U6462 (N_6462,N_5819,N_5632);
xor U6463 (N_6463,N_5518,N_5804);
nand U6464 (N_6464,N_5759,N_5962);
xor U6465 (N_6465,N_5848,N_5592);
xor U6466 (N_6466,N_5802,N_5590);
and U6467 (N_6467,N_5548,N_5933);
xnor U6468 (N_6468,N_5529,N_5689);
nor U6469 (N_6469,N_5685,N_5777);
nor U6470 (N_6470,N_5573,N_5586);
or U6471 (N_6471,N_5580,N_5672);
nand U6472 (N_6472,N_5925,N_5523);
or U6473 (N_6473,N_5691,N_5588);
or U6474 (N_6474,N_5821,N_5911);
and U6475 (N_6475,N_5536,N_5594);
or U6476 (N_6476,N_5874,N_5653);
nor U6477 (N_6477,N_5982,N_5645);
xnor U6478 (N_6478,N_5922,N_5569);
and U6479 (N_6479,N_5956,N_5585);
xnor U6480 (N_6480,N_5829,N_5662);
and U6481 (N_6481,N_5780,N_5990);
or U6482 (N_6482,N_5564,N_5908);
and U6483 (N_6483,N_5623,N_5694);
xor U6484 (N_6484,N_5686,N_5851);
nor U6485 (N_6485,N_5615,N_5771);
or U6486 (N_6486,N_5516,N_5702);
xor U6487 (N_6487,N_5984,N_5654);
and U6488 (N_6488,N_5654,N_5661);
nand U6489 (N_6489,N_5605,N_5880);
nand U6490 (N_6490,N_5970,N_5886);
and U6491 (N_6491,N_5532,N_5783);
nand U6492 (N_6492,N_5897,N_5606);
or U6493 (N_6493,N_5724,N_5905);
or U6494 (N_6494,N_5786,N_5593);
xor U6495 (N_6495,N_5618,N_5875);
or U6496 (N_6496,N_5763,N_5896);
nor U6497 (N_6497,N_5816,N_5995);
nand U6498 (N_6498,N_5934,N_5788);
xnor U6499 (N_6499,N_5606,N_5926);
nor U6500 (N_6500,N_6330,N_6473);
or U6501 (N_6501,N_6421,N_6123);
nor U6502 (N_6502,N_6004,N_6024);
and U6503 (N_6503,N_6134,N_6069);
and U6504 (N_6504,N_6451,N_6106);
and U6505 (N_6505,N_6392,N_6308);
nand U6506 (N_6506,N_6447,N_6234);
nor U6507 (N_6507,N_6335,N_6213);
nor U6508 (N_6508,N_6083,N_6080);
nor U6509 (N_6509,N_6446,N_6386);
nand U6510 (N_6510,N_6283,N_6224);
or U6511 (N_6511,N_6315,N_6455);
and U6512 (N_6512,N_6485,N_6204);
and U6513 (N_6513,N_6270,N_6179);
xor U6514 (N_6514,N_6238,N_6305);
xnor U6515 (N_6515,N_6435,N_6404);
and U6516 (N_6516,N_6449,N_6073);
and U6517 (N_6517,N_6099,N_6381);
nor U6518 (N_6518,N_6103,N_6144);
nand U6519 (N_6519,N_6076,N_6332);
nor U6520 (N_6520,N_6138,N_6302);
or U6521 (N_6521,N_6383,N_6104);
and U6522 (N_6522,N_6297,N_6491);
xnor U6523 (N_6523,N_6460,N_6275);
or U6524 (N_6524,N_6107,N_6130);
or U6525 (N_6525,N_6109,N_6389);
and U6526 (N_6526,N_6272,N_6145);
nor U6527 (N_6527,N_6273,N_6118);
and U6528 (N_6528,N_6259,N_6405);
nand U6529 (N_6529,N_6163,N_6424);
xor U6530 (N_6530,N_6085,N_6427);
and U6531 (N_6531,N_6422,N_6431);
or U6532 (N_6532,N_6197,N_6229);
xnor U6533 (N_6533,N_6218,N_6369);
or U6534 (N_6534,N_6046,N_6125);
xor U6535 (N_6535,N_6260,N_6232);
nand U6536 (N_6536,N_6194,N_6137);
or U6537 (N_6537,N_6051,N_6286);
nand U6538 (N_6538,N_6129,N_6290);
nor U6539 (N_6539,N_6113,N_6139);
and U6540 (N_6540,N_6445,N_6100);
or U6541 (N_6541,N_6052,N_6434);
and U6542 (N_6542,N_6030,N_6044);
or U6543 (N_6543,N_6396,N_6461);
and U6544 (N_6544,N_6230,N_6146);
and U6545 (N_6545,N_6122,N_6184);
nand U6546 (N_6546,N_6457,N_6198);
nor U6547 (N_6547,N_6150,N_6350);
or U6548 (N_6548,N_6340,N_6394);
nand U6549 (N_6549,N_6426,N_6237);
nor U6550 (N_6550,N_6191,N_6147);
or U6551 (N_6551,N_6292,N_6212);
xnor U6552 (N_6552,N_6117,N_6410);
and U6553 (N_6553,N_6195,N_6497);
xnor U6554 (N_6554,N_6385,N_6050);
nand U6555 (N_6555,N_6187,N_6301);
nor U6556 (N_6556,N_6412,N_6274);
nor U6557 (N_6557,N_6235,N_6017);
and U6558 (N_6558,N_6417,N_6438);
nand U6559 (N_6559,N_6012,N_6231);
or U6560 (N_6560,N_6192,N_6020);
nor U6561 (N_6561,N_6151,N_6088);
and U6562 (N_6562,N_6217,N_6484);
nor U6563 (N_6563,N_6053,N_6200);
xnor U6564 (N_6564,N_6425,N_6007);
nand U6565 (N_6565,N_6078,N_6364);
nand U6566 (N_6566,N_6280,N_6486);
or U6567 (N_6567,N_6331,N_6271);
nor U6568 (N_6568,N_6241,N_6257);
or U6569 (N_6569,N_6016,N_6105);
xor U6570 (N_6570,N_6289,N_6097);
nand U6571 (N_6571,N_6495,N_6156);
xor U6572 (N_6572,N_6397,N_6077);
and U6573 (N_6573,N_6154,N_6023);
nor U6574 (N_6574,N_6346,N_6262);
xnor U6575 (N_6575,N_6468,N_6098);
and U6576 (N_6576,N_6066,N_6131);
xor U6577 (N_6577,N_6307,N_6482);
nand U6578 (N_6578,N_6295,N_6488);
and U6579 (N_6579,N_6027,N_6003);
nor U6580 (N_6580,N_6058,N_6035);
and U6581 (N_6581,N_6296,N_6313);
xnor U6582 (N_6582,N_6323,N_6005);
and U6583 (N_6583,N_6440,N_6176);
nor U6584 (N_6584,N_6048,N_6472);
or U6585 (N_6585,N_6177,N_6322);
or U6586 (N_6586,N_6032,N_6031);
and U6587 (N_6587,N_6496,N_6380);
or U6588 (N_6588,N_6463,N_6094);
nand U6589 (N_6589,N_6268,N_6084);
or U6590 (N_6590,N_6454,N_6357);
nor U6591 (N_6591,N_6402,N_6040);
and U6592 (N_6592,N_6306,N_6303);
nor U6593 (N_6593,N_6119,N_6116);
xor U6594 (N_6594,N_6294,N_6038);
nor U6595 (N_6595,N_6319,N_6183);
xor U6596 (N_6596,N_6328,N_6339);
nor U6597 (N_6597,N_6401,N_6281);
xnor U6598 (N_6598,N_6399,N_6493);
nand U6599 (N_6599,N_6370,N_6367);
or U6600 (N_6600,N_6376,N_6102);
nand U6601 (N_6601,N_6343,N_6341);
or U6602 (N_6602,N_6018,N_6382);
and U6603 (N_6603,N_6333,N_6403);
nand U6604 (N_6604,N_6208,N_6471);
or U6605 (N_6605,N_6450,N_6236);
nand U6606 (N_6606,N_6063,N_6459);
and U6607 (N_6607,N_6193,N_6247);
nor U6608 (N_6608,N_6026,N_6348);
and U6609 (N_6609,N_6390,N_6133);
xnor U6610 (N_6610,N_6143,N_6010);
and U6611 (N_6611,N_6407,N_6413);
xor U6612 (N_6612,N_6439,N_6135);
xnor U6613 (N_6613,N_6152,N_6190);
and U6614 (N_6614,N_6456,N_6054);
xor U6615 (N_6615,N_6068,N_6222);
xor U6616 (N_6616,N_6489,N_6014);
nand U6617 (N_6617,N_6310,N_6009);
or U6618 (N_6618,N_6042,N_6060);
or U6619 (N_6619,N_6279,N_6476);
or U6620 (N_6620,N_6324,N_6115);
nand U6621 (N_6621,N_6498,N_6266);
or U6622 (N_6622,N_6349,N_6096);
nand U6623 (N_6623,N_6362,N_6360);
or U6624 (N_6624,N_6141,N_6249);
xnor U6625 (N_6625,N_6062,N_6406);
nand U6626 (N_6626,N_6128,N_6374);
or U6627 (N_6627,N_6325,N_6359);
nand U6628 (N_6628,N_6379,N_6168);
or U6629 (N_6629,N_6164,N_6028);
or U6630 (N_6630,N_6065,N_6242);
or U6631 (N_6631,N_6481,N_6000);
nor U6632 (N_6632,N_6448,N_6186);
and U6633 (N_6633,N_6311,N_6226);
nand U6634 (N_6634,N_6127,N_6087);
or U6635 (N_6635,N_6391,N_6314);
xnor U6636 (N_6636,N_6162,N_6409);
and U6637 (N_6637,N_6452,N_6165);
and U6638 (N_6638,N_6312,N_6264);
nand U6639 (N_6639,N_6211,N_6377);
and U6640 (N_6640,N_6199,N_6181);
xnor U6641 (N_6641,N_6466,N_6365);
xnor U6642 (N_6642,N_6220,N_6006);
and U6643 (N_6643,N_6008,N_6255);
xnor U6644 (N_6644,N_6252,N_6371);
nand U6645 (N_6645,N_6470,N_6356);
nor U6646 (N_6646,N_6041,N_6161);
xor U6647 (N_6647,N_6172,N_6037);
xor U6648 (N_6648,N_6136,N_6246);
or U6649 (N_6649,N_6278,N_6221);
nor U6650 (N_6650,N_6479,N_6345);
xnor U6651 (N_6651,N_6091,N_6153);
and U6652 (N_6652,N_6132,N_6428);
xor U6653 (N_6653,N_6347,N_6329);
nor U6654 (N_6654,N_6423,N_6061);
nand U6655 (N_6655,N_6025,N_6254);
and U6656 (N_6656,N_6372,N_6419);
and U6657 (N_6657,N_6110,N_6291);
or U6658 (N_6658,N_6056,N_6180);
xor U6659 (N_6659,N_6499,N_6092);
and U6660 (N_6660,N_6298,N_6429);
and U6661 (N_6661,N_6079,N_6288);
nor U6662 (N_6662,N_6057,N_6142);
and U6663 (N_6663,N_6320,N_6090);
or U6664 (N_6664,N_6317,N_6022);
xor U6665 (N_6665,N_6011,N_6368);
nor U6666 (N_6666,N_6398,N_6318);
nor U6667 (N_6667,N_6039,N_6067);
nor U6668 (N_6668,N_6047,N_6189);
xor U6669 (N_6669,N_6064,N_6338);
or U6670 (N_6670,N_6355,N_6124);
or U6671 (N_6671,N_6477,N_6393);
and U6672 (N_6672,N_6443,N_6245);
or U6673 (N_6673,N_6304,N_6327);
nor U6674 (N_6674,N_6276,N_6469);
or U6675 (N_6675,N_6326,N_6244);
and U6676 (N_6676,N_6420,N_6384);
or U6677 (N_6677,N_6219,N_6111);
or U6678 (N_6678,N_6474,N_6086);
nor U6679 (N_6679,N_6081,N_6228);
and U6680 (N_6680,N_6001,N_6442);
nand U6681 (N_6681,N_6021,N_6361);
nor U6682 (N_6682,N_6201,N_6480);
nor U6683 (N_6683,N_6436,N_6101);
and U6684 (N_6684,N_6114,N_6336);
xnor U6685 (N_6685,N_6214,N_6248);
nor U6686 (N_6686,N_6240,N_6216);
nor U6687 (N_6687,N_6185,N_6112);
or U6688 (N_6688,N_6169,N_6159);
and U6689 (N_6689,N_6366,N_6160);
or U6690 (N_6690,N_6490,N_6344);
nand U6691 (N_6691,N_6203,N_6263);
nand U6692 (N_6692,N_6072,N_6167);
nor U6693 (N_6693,N_6227,N_6171);
and U6694 (N_6694,N_6174,N_6408);
and U6695 (N_6695,N_6074,N_6444);
nand U6696 (N_6696,N_6206,N_6082);
or U6697 (N_6697,N_6475,N_6277);
or U6698 (N_6698,N_6173,N_6055);
or U6699 (N_6699,N_6358,N_6209);
and U6700 (N_6700,N_6158,N_6019);
and U6701 (N_6701,N_6170,N_6353);
xnor U6702 (N_6702,N_6196,N_6478);
nand U6703 (N_6703,N_6071,N_6492);
and U6704 (N_6704,N_6182,N_6095);
and U6705 (N_6705,N_6418,N_6387);
nand U6706 (N_6706,N_6049,N_6239);
nand U6707 (N_6707,N_6126,N_6414);
nor U6708 (N_6708,N_6223,N_6175);
or U6709 (N_6709,N_6108,N_6494);
xor U6710 (N_6710,N_6258,N_6309);
and U6711 (N_6711,N_6155,N_6045);
nor U6712 (N_6712,N_6059,N_6433);
and U6713 (N_6713,N_6299,N_6215);
nand U6714 (N_6714,N_6437,N_6033);
or U6715 (N_6715,N_6002,N_6121);
nor U6716 (N_6716,N_6013,N_6029);
nor U6717 (N_6717,N_6070,N_6352);
nand U6718 (N_6718,N_6089,N_6034);
and U6719 (N_6719,N_6375,N_6373);
nand U6720 (N_6720,N_6351,N_6256);
and U6721 (N_6721,N_6411,N_6334);
xor U6722 (N_6722,N_6036,N_6300);
or U6723 (N_6723,N_6075,N_6120);
and U6724 (N_6724,N_6225,N_6464);
nand U6725 (N_6725,N_6467,N_6285);
nor U6726 (N_6726,N_6178,N_6316);
nand U6727 (N_6727,N_6205,N_6458);
nand U6728 (N_6728,N_6157,N_6282);
nand U6729 (N_6729,N_6416,N_6465);
nor U6730 (N_6730,N_6400,N_6462);
nand U6731 (N_6731,N_6483,N_6354);
nand U6732 (N_6732,N_6140,N_6149);
and U6733 (N_6733,N_6210,N_6337);
nor U6734 (N_6734,N_6243,N_6253);
xor U6735 (N_6735,N_6166,N_6202);
or U6736 (N_6736,N_6293,N_6342);
or U6737 (N_6737,N_6265,N_6321);
and U6738 (N_6738,N_6432,N_6233);
or U6739 (N_6739,N_6395,N_6388);
or U6740 (N_6740,N_6043,N_6430);
nand U6741 (N_6741,N_6378,N_6261);
and U6742 (N_6742,N_6251,N_6267);
xnor U6743 (N_6743,N_6015,N_6415);
and U6744 (N_6744,N_6441,N_6287);
xor U6745 (N_6745,N_6093,N_6188);
or U6746 (N_6746,N_6284,N_6250);
nand U6747 (N_6747,N_6148,N_6453);
xnor U6748 (N_6748,N_6207,N_6363);
xor U6749 (N_6749,N_6269,N_6487);
and U6750 (N_6750,N_6399,N_6381);
nor U6751 (N_6751,N_6354,N_6303);
nor U6752 (N_6752,N_6376,N_6189);
and U6753 (N_6753,N_6398,N_6196);
nand U6754 (N_6754,N_6489,N_6396);
xor U6755 (N_6755,N_6155,N_6054);
nand U6756 (N_6756,N_6073,N_6273);
nor U6757 (N_6757,N_6400,N_6346);
or U6758 (N_6758,N_6386,N_6489);
or U6759 (N_6759,N_6050,N_6397);
nor U6760 (N_6760,N_6287,N_6063);
nand U6761 (N_6761,N_6333,N_6125);
or U6762 (N_6762,N_6277,N_6032);
and U6763 (N_6763,N_6484,N_6304);
nor U6764 (N_6764,N_6486,N_6381);
xnor U6765 (N_6765,N_6321,N_6492);
and U6766 (N_6766,N_6272,N_6108);
or U6767 (N_6767,N_6382,N_6067);
nand U6768 (N_6768,N_6020,N_6256);
nand U6769 (N_6769,N_6056,N_6061);
and U6770 (N_6770,N_6204,N_6203);
or U6771 (N_6771,N_6074,N_6028);
and U6772 (N_6772,N_6319,N_6384);
and U6773 (N_6773,N_6345,N_6346);
xor U6774 (N_6774,N_6125,N_6241);
nor U6775 (N_6775,N_6133,N_6311);
xor U6776 (N_6776,N_6391,N_6311);
and U6777 (N_6777,N_6453,N_6014);
nand U6778 (N_6778,N_6012,N_6457);
and U6779 (N_6779,N_6323,N_6294);
xnor U6780 (N_6780,N_6071,N_6260);
xor U6781 (N_6781,N_6266,N_6465);
nor U6782 (N_6782,N_6013,N_6337);
xnor U6783 (N_6783,N_6188,N_6175);
nand U6784 (N_6784,N_6349,N_6412);
nor U6785 (N_6785,N_6158,N_6299);
and U6786 (N_6786,N_6243,N_6233);
nor U6787 (N_6787,N_6155,N_6201);
nand U6788 (N_6788,N_6449,N_6106);
or U6789 (N_6789,N_6035,N_6177);
nor U6790 (N_6790,N_6285,N_6213);
xor U6791 (N_6791,N_6011,N_6119);
xnor U6792 (N_6792,N_6487,N_6391);
or U6793 (N_6793,N_6492,N_6204);
xnor U6794 (N_6794,N_6117,N_6054);
or U6795 (N_6795,N_6081,N_6080);
nand U6796 (N_6796,N_6256,N_6466);
nor U6797 (N_6797,N_6273,N_6128);
nor U6798 (N_6798,N_6217,N_6004);
nand U6799 (N_6799,N_6221,N_6425);
or U6800 (N_6800,N_6062,N_6353);
nand U6801 (N_6801,N_6065,N_6081);
xnor U6802 (N_6802,N_6069,N_6461);
nand U6803 (N_6803,N_6104,N_6369);
and U6804 (N_6804,N_6063,N_6160);
nor U6805 (N_6805,N_6116,N_6423);
xor U6806 (N_6806,N_6132,N_6245);
and U6807 (N_6807,N_6418,N_6202);
or U6808 (N_6808,N_6131,N_6349);
nor U6809 (N_6809,N_6223,N_6338);
nand U6810 (N_6810,N_6435,N_6352);
or U6811 (N_6811,N_6200,N_6426);
and U6812 (N_6812,N_6199,N_6342);
and U6813 (N_6813,N_6116,N_6430);
xnor U6814 (N_6814,N_6464,N_6466);
xor U6815 (N_6815,N_6274,N_6262);
nor U6816 (N_6816,N_6341,N_6042);
and U6817 (N_6817,N_6223,N_6270);
nand U6818 (N_6818,N_6417,N_6182);
and U6819 (N_6819,N_6094,N_6160);
or U6820 (N_6820,N_6068,N_6459);
nor U6821 (N_6821,N_6111,N_6459);
or U6822 (N_6822,N_6108,N_6240);
and U6823 (N_6823,N_6485,N_6324);
nor U6824 (N_6824,N_6426,N_6026);
xnor U6825 (N_6825,N_6323,N_6090);
and U6826 (N_6826,N_6065,N_6040);
xnor U6827 (N_6827,N_6365,N_6046);
xnor U6828 (N_6828,N_6410,N_6046);
xnor U6829 (N_6829,N_6052,N_6114);
or U6830 (N_6830,N_6376,N_6202);
and U6831 (N_6831,N_6404,N_6050);
and U6832 (N_6832,N_6257,N_6183);
nand U6833 (N_6833,N_6050,N_6358);
nor U6834 (N_6834,N_6092,N_6084);
nand U6835 (N_6835,N_6217,N_6308);
nor U6836 (N_6836,N_6323,N_6377);
or U6837 (N_6837,N_6397,N_6123);
xnor U6838 (N_6838,N_6118,N_6284);
and U6839 (N_6839,N_6499,N_6201);
nand U6840 (N_6840,N_6095,N_6208);
xnor U6841 (N_6841,N_6325,N_6006);
nand U6842 (N_6842,N_6453,N_6196);
or U6843 (N_6843,N_6349,N_6193);
xnor U6844 (N_6844,N_6472,N_6133);
nand U6845 (N_6845,N_6125,N_6297);
xor U6846 (N_6846,N_6213,N_6297);
xor U6847 (N_6847,N_6499,N_6126);
xnor U6848 (N_6848,N_6326,N_6214);
nand U6849 (N_6849,N_6471,N_6206);
and U6850 (N_6850,N_6264,N_6362);
nand U6851 (N_6851,N_6103,N_6055);
nand U6852 (N_6852,N_6390,N_6155);
and U6853 (N_6853,N_6320,N_6001);
or U6854 (N_6854,N_6150,N_6322);
xor U6855 (N_6855,N_6099,N_6234);
nand U6856 (N_6856,N_6033,N_6172);
and U6857 (N_6857,N_6457,N_6070);
nand U6858 (N_6858,N_6052,N_6361);
xor U6859 (N_6859,N_6026,N_6159);
nor U6860 (N_6860,N_6379,N_6044);
xor U6861 (N_6861,N_6363,N_6211);
or U6862 (N_6862,N_6108,N_6154);
or U6863 (N_6863,N_6443,N_6098);
or U6864 (N_6864,N_6183,N_6132);
nor U6865 (N_6865,N_6282,N_6243);
nor U6866 (N_6866,N_6012,N_6046);
or U6867 (N_6867,N_6252,N_6388);
xnor U6868 (N_6868,N_6289,N_6291);
nor U6869 (N_6869,N_6090,N_6460);
or U6870 (N_6870,N_6131,N_6025);
or U6871 (N_6871,N_6296,N_6447);
or U6872 (N_6872,N_6312,N_6177);
nand U6873 (N_6873,N_6207,N_6221);
xor U6874 (N_6874,N_6154,N_6367);
or U6875 (N_6875,N_6052,N_6020);
xor U6876 (N_6876,N_6051,N_6418);
nand U6877 (N_6877,N_6466,N_6492);
or U6878 (N_6878,N_6115,N_6163);
xor U6879 (N_6879,N_6162,N_6298);
nor U6880 (N_6880,N_6246,N_6240);
and U6881 (N_6881,N_6392,N_6164);
and U6882 (N_6882,N_6154,N_6356);
nor U6883 (N_6883,N_6437,N_6120);
nor U6884 (N_6884,N_6417,N_6163);
and U6885 (N_6885,N_6185,N_6261);
nand U6886 (N_6886,N_6294,N_6037);
nand U6887 (N_6887,N_6012,N_6311);
nor U6888 (N_6888,N_6497,N_6322);
nor U6889 (N_6889,N_6488,N_6251);
or U6890 (N_6890,N_6138,N_6402);
nor U6891 (N_6891,N_6386,N_6205);
and U6892 (N_6892,N_6344,N_6117);
or U6893 (N_6893,N_6081,N_6001);
xnor U6894 (N_6894,N_6314,N_6201);
nor U6895 (N_6895,N_6388,N_6379);
nor U6896 (N_6896,N_6129,N_6187);
or U6897 (N_6897,N_6363,N_6176);
or U6898 (N_6898,N_6167,N_6239);
xor U6899 (N_6899,N_6085,N_6160);
nor U6900 (N_6900,N_6462,N_6454);
and U6901 (N_6901,N_6422,N_6011);
nand U6902 (N_6902,N_6321,N_6175);
or U6903 (N_6903,N_6430,N_6492);
xor U6904 (N_6904,N_6100,N_6498);
and U6905 (N_6905,N_6397,N_6168);
nor U6906 (N_6906,N_6285,N_6328);
xnor U6907 (N_6907,N_6226,N_6239);
or U6908 (N_6908,N_6337,N_6010);
or U6909 (N_6909,N_6231,N_6362);
nor U6910 (N_6910,N_6129,N_6364);
or U6911 (N_6911,N_6304,N_6085);
or U6912 (N_6912,N_6230,N_6088);
nand U6913 (N_6913,N_6162,N_6078);
and U6914 (N_6914,N_6300,N_6222);
nor U6915 (N_6915,N_6040,N_6080);
nor U6916 (N_6916,N_6044,N_6432);
nand U6917 (N_6917,N_6314,N_6340);
or U6918 (N_6918,N_6217,N_6485);
nor U6919 (N_6919,N_6012,N_6446);
nor U6920 (N_6920,N_6216,N_6183);
and U6921 (N_6921,N_6121,N_6297);
xor U6922 (N_6922,N_6411,N_6176);
nand U6923 (N_6923,N_6054,N_6104);
or U6924 (N_6924,N_6252,N_6240);
xor U6925 (N_6925,N_6206,N_6202);
nand U6926 (N_6926,N_6050,N_6261);
nand U6927 (N_6927,N_6101,N_6494);
or U6928 (N_6928,N_6012,N_6178);
nand U6929 (N_6929,N_6465,N_6485);
xor U6930 (N_6930,N_6128,N_6335);
xnor U6931 (N_6931,N_6129,N_6360);
xnor U6932 (N_6932,N_6226,N_6480);
and U6933 (N_6933,N_6091,N_6048);
xnor U6934 (N_6934,N_6174,N_6212);
nand U6935 (N_6935,N_6152,N_6038);
and U6936 (N_6936,N_6043,N_6435);
and U6937 (N_6937,N_6227,N_6161);
and U6938 (N_6938,N_6322,N_6248);
xor U6939 (N_6939,N_6103,N_6146);
and U6940 (N_6940,N_6264,N_6058);
nand U6941 (N_6941,N_6111,N_6262);
and U6942 (N_6942,N_6064,N_6344);
or U6943 (N_6943,N_6202,N_6110);
or U6944 (N_6944,N_6226,N_6326);
nor U6945 (N_6945,N_6162,N_6395);
nor U6946 (N_6946,N_6181,N_6167);
nor U6947 (N_6947,N_6286,N_6421);
or U6948 (N_6948,N_6089,N_6315);
xnor U6949 (N_6949,N_6211,N_6087);
xnor U6950 (N_6950,N_6267,N_6464);
nand U6951 (N_6951,N_6178,N_6164);
nor U6952 (N_6952,N_6252,N_6397);
and U6953 (N_6953,N_6401,N_6142);
xor U6954 (N_6954,N_6255,N_6427);
xnor U6955 (N_6955,N_6099,N_6093);
nand U6956 (N_6956,N_6121,N_6456);
or U6957 (N_6957,N_6376,N_6481);
and U6958 (N_6958,N_6175,N_6465);
and U6959 (N_6959,N_6059,N_6116);
xor U6960 (N_6960,N_6375,N_6318);
xor U6961 (N_6961,N_6437,N_6341);
and U6962 (N_6962,N_6420,N_6378);
nand U6963 (N_6963,N_6345,N_6018);
nor U6964 (N_6964,N_6409,N_6210);
xnor U6965 (N_6965,N_6023,N_6429);
and U6966 (N_6966,N_6296,N_6001);
or U6967 (N_6967,N_6037,N_6206);
nor U6968 (N_6968,N_6400,N_6369);
nor U6969 (N_6969,N_6267,N_6421);
nand U6970 (N_6970,N_6039,N_6049);
xor U6971 (N_6971,N_6142,N_6352);
nand U6972 (N_6972,N_6242,N_6481);
nor U6973 (N_6973,N_6289,N_6343);
and U6974 (N_6974,N_6202,N_6235);
nor U6975 (N_6975,N_6023,N_6455);
xor U6976 (N_6976,N_6230,N_6180);
and U6977 (N_6977,N_6396,N_6181);
or U6978 (N_6978,N_6226,N_6048);
nand U6979 (N_6979,N_6485,N_6032);
xor U6980 (N_6980,N_6335,N_6265);
or U6981 (N_6981,N_6015,N_6035);
or U6982 (N_6982,N_6237,N_6260);
xor U6983 (N_6983,N_6396,N_6313);
xor U6984 (N_6984,N_6309,N_6164);
nor U6985 (N_6985,N_6181,N_6265);
and U6986 (N_6986,N_6227,N_6023);
and U6987 (N_6987,N_6004,N_6022);
and U6988 (N_6988,N_6222,N_6257);
and U6989 (N_6989,N_6258,N_6052);
or U6990 (N_6990,N_6271,N_6499);
and U6991 (N_6991,N_6019,N_6401);
xor U6992 (N_6992,N_6323,N_6350);
and U6993 (N_6993,N_6166,N_6159);
or U6994 (N_6994,N_6223,N_6198);
and U6995 (N_6995,N_6181,N_6314);
xnor U6996 (N_6996,N_6096,N_6434);
nor U6997 (N_6997,N_6154,N_6168);
xor U6998 (N_6998,N_6388,N_6010);
and U6999 (N_6999,N_6472,N_6104);
and U7000 (N_7000,N_6644,N_6880);
nand U7001 (N_7001,N_6613,N_6507);
nor U7002 (N_7002,N_6844,N_6762);
or U7003 (N_7003,N_6637,N_6666);
or U7004 (N_7004,N_6500,N_6615);
nand U7005 (N_7005,N_6861,N_6651);
nand U7006 (N_7006,N_6915,N_6765);
or U7007 (N_7007,N_6771,N_6553);
and U7008 (N_7008,N_6531,N_6786);
or U7009 (N_7009,N_6751,N_6726);
nand U7010 (N_7010,N_6895,N_6526);
nand U7011 (N_7011,N_6974,N_6556);
nor U7012 (N_7012,N_6860,N_6816);
or U7013 (N_7013,N_6717,N_6777);
nand U7014 (N_7014,N_6910,N_6599);
nor U7015 (N_7015,N_6800,N_6977);
xnor U7016 (N_7016,N_6521,N_6967);
or U7017 (N_7017,N_6904,N_6769);
nand U7018 (N_7018,N_6929,N_6559);
xor U7019 (N_7019,N_6731,N_6601);
or U7020 (N_7020,N_6573,N_6900);
nand U7021 (N_7021,N_6891,N_6595);
nand U7022 (N_7022,N_6767,N_6505);
and U7023 (N_7023,N_6715,N_6571);
or U7024 (N_7024,N_6728,N_6886);
nor U7025 (N_7025,N_6652,N_6874);
xnor U7026 (N_7026,N_6923,N_6697);
nor U7027 (N_7027,N_6628,N_6789);
nor U7028 (N_7028,N_6858,N_6951);
xnor U7029 (N_7029,N_6940,N_6980);
nand U7030 (N_7030,N_6683,N_6945);
nor U7031 (N_7031,N_6782,N_6976);
nor U7032 (N_7032,N_6527,N_6864);
nand U7033 (N_7033,N_6987,N_6550);
nor U7034 (N_7034,N_6881,N_6828);
nand U7035 (N_7035,N_6722,N_6759);
or U7036 (N_7036,N_6854,N_6859);
and U7037 (N_7037,N_6956,N_6791);
nand U7038 (N_7038,N_6581,N_6862);
or U7039 (N_7039,N_6991,N_6914);
xnor U7040 (N_7040,N_6868,N_6947);
or U7041 (N_7041,N_6905,N_6834);
and U7042 (N_7042,N_6846,N_6654);
nor U7043 (N_7043,N_6582,N_6756);
nand U7044 (N_7044,N_6981,N_6889);
nand U7045 (N_7045,N_6774,N_6730);
and U7046 (N_7046,N_6803,N_6824);
and U7047 (N_7047,N_6810,N_6952);
and U7048 (N_7048,N_6622,N_6503);
xnor U7049 (N_7049,N_6733,N_6963);
nor U7050 (N_7050,N_6525,N_6982);
nor U7051 (N_7051,N_6566,N_6916);
and U7052 (N_7052,N_6607,N_6742);
nor U7053 (N_7053,N_6568,N_6872);
and U7054 (N_7054,N_6785,N_6994);
or U7055 (N_7055,N_6529,N_6937);
nor U7056 (N_7056,N_6631,N_6545);
nand U7057 (N_7057,N_6680,N_6734);
xor U7058 (N_7058,N_6646,N_6551);
nor U7059 (N_7059,N_6539,N_6931);
and U7060 (N_7060,N_6845,N_6993);
xor U7061 (N_7061,N_6924,N_6969);
or U7062 (N_7062,N_6564,N_6515);
or U7063 (N_7063,N_6784,N_6988);
xor U7064 (N_7064,N_6938,N_6509);
nor U7065 (N_7065,N_6533,N_6892);
nor U7066 (N_7066,N_6712,N_6577);
or U7067 (N_7067,N_6518,N_6598);
xor U7068 (N_7068,N_6962,N_6801);
or U7069 (N_7069,N_6692,N_6594);
nor U7070 (N_7070,N_6798,N_6708);
nor U7071 (N_7071,N_6537,N_6671);
or U7072 (N_7072,N_6657,N_6870);
xor U7073 (N_7073,N_6887,N_6829);
xor U7074 (N_7074,N_6656,N_6535);
nand U7075 (N_7075,N_6760,N_6688);
nand U7076 (N_7076,N_6627,N_6848);
xnor U7077 (N_7077,N_6971,N_6758);
or U7078 (N_7078,N_6517,N_6741);
or U7079 (N_7079,N_6635,N_6669);
and U7080 (N_7080,N_6705,N_6681);
xnor U7081 (N_7081,N_6569,N_6538);
or U7082 (N_7082,N_6778,N_6700);
or U7083 (N_7083,N_6841,N_6704);
xor U7084 (N_7084,N_6678,N_6839);
nor U7085 (N_7085,N_6580,N_6699);
and U7086 (N_7086,N_6735,N_6805);
and U7087 (N_7087,N_6833,N_6973);
nor U7088 (N_7088,N_6608,N_6794);
xnor U7089 (N_7089,N_6836,N_6561);
nand U7090 (N_7090,N_6847,N_6516);
nor U7091 (N_7091,N_6811,N_6621);
or U7092 (N_7092,N_6970,N_6686);
or U7093 (N_7093,N_6665,N_6941);
or U7094 (N_7094,N_6633,N_6992);
and U7095 (N_7095,N_6743,N_6783);
nand U7096 (N_7096,N_6546,N_6574);
nor U7097 (N_7097,N_6523,N_6832);
nand U7098 (N_7098,N_6648,N_6807);
nand U7099 (N_7099,N_6799,N_6512);
nand U7100 (N_7100,N_6694,N_6966);
nand U7101 (N_7101,N_6948,N_6701);
or U7102 (N_7102,N_6806,N_6558);
xnor U7103 (N_7103,N_6519,N_6884);
xor U7104 (N_7104,N_6689,N_6989);
nand U7105 (N_7105,N_6695,N_6894);
nand U7106 (N_7106,N_6592,N_6612);
and U7107 (N_7107,N_6618,N_6943);
nand U7108 (N_7108,N_6831,N_6685);
nand U7109 (N_7109,N_6640,N_6504);
and U7110 (N_7110,N_6912,N_6664);
or U7111 (N_7111,N_6953,N_6925);
or U7112 (N_7112,N_6714,N_6520);
and U7113 (N_7113,N_6885,N_6950);
nand U7114 (N_7114,N_6614,N_6918);
nand U7115 (N_7115,N_6638,N_6849);
xor U7116 (N_7116,N_6865,N_6590);
nor U7117 (N_7117,N_6548,N_6871);
and U7118 (N_7118,N_6957,N_6822);
or U7119 (N_7119,N_6761,N_6926);
nor U7120 (N_7120,N_6593,N_6619);
nor U7121 (N_7121,N_6532,N_6611);
or U7122 (N_7122,N_6610,N_6588);
nor U7123 (N_7123,N_6673,N_6522);
nor U7124 (N_7124,N_6932,N_6772);
nand U7125 (N_7125,N_6818,N_6634);
xor U7126 (N_7126,N_6825,N_6711);
xor U7127 (N_7127,N_6578,N_6764);
nand U7128 (N_7128,N_6837,N_6668);
or U7129 (N_7129,N_6720,N_6879);
nor U7130 (N_7130,N_6935,N_6755);
nand U7131 (N_7131,N_6746,N_6642);
or U7132 (N_7132,N_6819,N_6790);
and U7133 (N_7133,N_6721,N_6639);
xnor U7134 (N_7134,N_6620,N_6677);
nor U7135 (N_7135,N_6514,N_6934);
and U7136 (N_7136,N_6753,N_6852);
nand U7137 (N_7137,N_6792,N_6584);
xnor U7138 (N_7138,N_6534,N_6745);
and U7139 (N_7139,N_6661,N_6676);
nor U7140 (N_7140,N_6600,N_6687);
nand U7141 (N_7141,N_6587,N_6921);
or U7142 (N_7142,N_6867,N_6624);
and U7143 (N_7143,N_6552,N_6575);
and U7144 (N_7144,N_6773,N_6549);
nand U7145 (N_7145,N_6876,N_6530);
xor U7146 (N_7146,N_6675,N_6907);
nand U7147 (N_7147,N_6835,N_6986);
nor U7148 (N_7148,N_6682,N_6779);
and U7149 (N_7149,N_6738,N_6703);
nor U7150 (N_7150,N_6873,N_6606);
nor U7151 (N_7151,N_6897,N_6555);
nor U7152 (N_7152,N_6540,N_6911);
and U7153 (N_7153,N_6902,N_6576);
and U7154 (N_7154,N_6939,N_6890);
or U7155 (N_7155,N_6972,N_6709);
nand U7156 (N_7156,N_6729,N_6757);
and U7157 (N_7157,N_6579,N_6899);
xnor U7158 (N_7158,N_6853,N_6572);
and U7159 (N_7159,N_6723,N_6737);
and U7160 (N_7160,N_6842,N_6713);
and U7161 (N_7161,N_6616,N_6696);
nand U7162 (N_7162,N_6562,N_6649);
xor U7163 (N_7163,N_6547,N_6707);
or U7164 (N_7164,N_6903,N_6855);
nand U7165 (N_7165,N_6793,N_6716);
nand U7166 (N_7166,N_6510,N_6710);
xor U7167 (N_7167,N_6797,N_6843);
nand U7168 (N_7168,N_6597,N_6809);
nor U7169 (N_7169,N_6752,N_6693);
xor U7170 (N_7170,N_6630,N_6670);
or U7171 (N_7171,N_6511,N_6567);
nand U7172 (N_7172,N_6719,N_6602);
nand U7173 (N_7173,N_6660,N_6857);
xnor U7174 (N_7174,N_6754,N_6983);
nor U7175 (N_7175,N_6544,N_6732);
and U7176 (N_7176,N_6702,N_6998);
and U7177 (N_7177,N_6893,N_6999);
nand U7178 (N_7178,N_6698,N_6604);
xor U7179 (N_7179,N_6840,N_6820);
and U7180 (N_7180,N_6959,N_6508);
or U7181 (N_7181,N_6898,N_6570);
nor U7182 (N_7182,N_6827,N_6543);
nor U7183 (N_7183,N_6776,N_6913);
xnor U7184 (N_7184,N_6906,N_6869);
nor U7185 (N_7185,N_6796,N_6645);
or U7186 (N_7186,N_6740,N_6749);
nor U7187 (N_7187,N_6672,N_6863);
nand U7188 (N_7188,N_6659,N_6978);
xnor U7189 (N_7189,N_6933,N_6770);
nor U7190 (N_7190,N_6875,N_6922);
or U7191 (N_7191,N_6585,N_6795);
nor U7192 (N_7192,N_6690,N_6787);
nand U7193 (N_7193,N_6965,N_6985);
xnor U7194 (N_7194,N_6609,N_6821);
xnor U7195 (N_7195,N_6662,N_6815);
and U7196 (N_7196,N_6501,N_6856);
nor U7197 (N_7197,N_6586,N_6928);
xor U7198 (N_7198,N_6942,N_6882);
and U7199 (N_7199,N_6866,N_6768);
and U7200 (N_7200,N_6838,N_6725);
or U7201 (N_7201,N_6936,N_6917);
nand U7202 (N_7202,N_6927,N_6563);
and U7203 (N_7203,N_6812,N_6605);
nand U7204 (N_7204,N_6990,N_6896);
and U7205 (N_7205,N_6502,N_6641);
nand U7206 (N_7206,N_6650,N_6542);
nand U7207 (N_7207,N_6823,N_6850);
or U7208 (N_7208,N_6954,N_6766);
nand U7209 (N_7209,N_6817,N_6513);
nand U7210 (N_7210,N_6617,N_6653);
nor U7211 (N_7211,N_6663,N_6877);
nor U7212 (N_7212,N_6541,N_6920);
nand U7213 (N_7213,N_6591,N_6706);
or U7214 (N_7214,N_6826,N_6565);
and U7215 (N_7215,N_6739,N_6744);
and U7216 (N_7216,N_6629,N_6736);
xnor U7217 (N_7217,N_6727,N_6557);
xor U7218 (N_7218,N_6536,N_6908);
nand U7219 (N_7219,N_6747,N_6658);
nand U7220 (N_7220,N_6647,N_6997);
xor U7221 (N_7221,N_6830,N_6901);
xor U7222 (N_7222,N_6554,N_6775);
and U7223 (N_7223,N_6984,N_6560);
or U7224 (N_7224,N_6625,N_6748);
nand U7225 (N_7225,N_6968,N_6883);
and U7226 (N_7226,N_6691,N_6724);
and U7227 (N_7227,N_6909,N_6524);
or U7228 (N_7228,N_6679,N_6506);
or U7229 (N_7229,N_6655,N_6802);
or U7230 (N_7230,N_6949,N_6944);
nand U7231 (N_7231,N_6750,N_6788);
nand U7232 (N_7232,N_6946,N_6781);
nor U7233 (N_7233,N_6596,N_6979);
xor U7234 (N_7234,N_6964,N_6804);
nand U7235 (N_7235,N_6878,N_6995);
or U7236 (N_7236,N_6674,N_6960);
xnor U7237 (N_7237,N_6623,N_6583);
or U7238 (N_7238,N_6632,N_6961);
xor U7239 (N_7239,N_6958,N_6919);
xor U7240 (N_7240,N_6643,N_6780);
or U7241 (N_7241,N_6851,N_6888);
xnor U7242 (N_7242,N_6626,N_6996);
or U7243 (N_7243,N_6955,N_6528);
and U7244 (N_7244,N_6763,N_6718);
nand U7245 (N_7245,N_6636,N_6814);
xnor U7246 (N_7246,N_6813,N_6589);
xor U7247 (N_7247,N_6808,N_6603);
or U7248 (N_7248,N_6667,N_6975);
nand U7249 (N_7249,N_6930,N_6684);
nor U7250 (N_7250,N_6544,N_6537);
xnor U7251 (N_7251,N_6821,N_6990);
or U7252 (N_7252,N_6898,N_6777);
and U7253 (N_7253,N_6799,N_6888);
or U7254 (N_7254,N_6760,N_6785);
nor U7255 (N_7255,N_6611,N_6552);
and U7256 (N_7256,N_6932,N_6599);
nor U7257 (N_7257,N_6731,N_6685);
or U7258 (N_7258,N_6680,N_6884);
xor U7259 (N_7259,N_6526,N_6978);
xor U7260 (N_7260,N_6656,N_6642);
xor U7261 (N_7261,N_6846,N_6629);
xor U7262 (N_7262,N_6809,N_6855);
nand U7263 (N_7263,N_6864,N_6989);
nand U7264 (N_7264,N_6696,N_6906);
nand U7265 (N_7265,N_6818,N_6802);
xnor U7266 (N_7266,N_6757,N_6575);
nor U7267 (N_7267,N_6695,N_6602);
and U7268 (N_7268,N_6786,N_6710);
nand U7269 (N_7269,N_6916,N_6850);
nor U7270 (N_7270,N_6897,N_6858);
or U7271 (N_7271,N_6908,N_6659);
or U7272 (N_7272,N_6672,N_6587);
or U7273 (N_7273,N_6954,N_6581);
nand U7274 (N_7274,N_6725,N_6763);
or U7275 (N_7275,N_6631,N_6758);
nor U7276 (N_7276,N_6776,N_6722);
nor U7277 (N_7277,N_6957,N_6722);
and U7278 (N_7278,N_6629,N_6929);
and U7279 (N_7279,N_6932,N_6617);
and U7280 (N_7280,N_6614,N_6913);
nand U7281 (N_7281,N_6646,N_6739);
nor U7282 (N_7282,N_6677,N_6509);
or U7283 (N_7283,N_6557,N_6542);
and U7284 (N_7284,N_6872,N_6899);
nor U7285 (N_7285,N_6649,N_6956);
nor U7286 (N_7286,N_6634,N_6549);
or U7287 (N_7287,N_6569,N_6900);
nor U7288 (N_7288,N_6674,N_6842);
nand U7289 (N_7289,N_6505,N_6536);
xor U7290 (N_7290,N_6915,N_6888);
nand U7291 (N_7291,N_6650,N_6916);
nor U7292 (N_7292,N_6857,N_6598);
xor U7293 (N_7293,N_6645,N_6598);
or U7294 (N_7294,N_6513,N_6630);
xor U7295 (N_7295,N_6561,N_6978);
xnor U7296 (N_7296,N_6503,N_6998);
and U7297 (N_7297,N_6837,N_6956);
nor U7298 (N_7298,N_6759,N_6884);
nor U7299 (N_7299,N_6578,N_6601);
nor U7300 (N_7300,N_6531,N_6807);
or U7301 (N_7301,N_6777,N_6707);
or U7302 (N_7302,N_6504,N_6531);
nand U7303 (N_7303,N_6719,N_6752);
and U7304 (N_7304,N_6953,N_6681);
and U7305 (N_7305,N_6961,N_6590);
xor U7306 (N_7306,N_6806,N_6622);
nand U7307 (N_7307,N_6742,N_6563);
or U7308 (N_7308,N_6518,N_6769);
or U7309 (N_7309,N_6674,N_6791);
nand U7310 (N_7310,N_6720,N_6515);
nand U7311 (N_7311,N_6941,N_6787);
nand U7312 (N_7312,N_6507,N_6725);
xor U7313 (N_7313,N_6820,N_6899);
nand U7314 (N_7314,N_6714,N_6946);
nor U7315 (N_7315,N_6572,N_6966);
nand U7316 (N_7316,N_6854,N_6752);
and U7317 (N_7317,N_6939,N_6958);
or U7318 (N_7318,N_6686,N_6906);
or U7319 (N_7319,N_6684,N_6665);
xor U7320 (N_7320,N_6938,N_6518);
and U7321 (N_7321,N_6798,N_6677);
nand U7322 (N_7322,N_6742,N_6734);
or U7323 (N_7323,N_6757,N_6989);
xnor U7324 (N_7324,N_6766,N_6726);
and U7325 (N_7325,N_6841,N_6699);
nand U7326 (N_7326,N_6699,N_6977);
or U7327 (N_7327,N_6559,N_6863);
or U7328 (N_7328,N_6752,N_6840);
nor U7329 (N_7329,N_6791,N_6811);
and U7330 (N_7330,N_6766,N_6813);
nand U7331 (N_7331,N_6812,N_6869);
xnor U7332 (N_7332,N_6892,N_6827);
and U7333 (N_7333,N_6862,N_6847);
or U7334 (N_7334,N_6726,N_6597);
and U7335 (N_7335,N_6533,N_6557);
nand U7336 (N_7336,N_6820,N_6683);
or U7337 (N_7337,N_6571,N_6950);
or U7338 (N_7338,N_6820,N_6712);
or U7339 (N_7339,N_6983,N_6887);
xnor U7340 (N_7340,N_6677,N_6741);
xor U7341 (N_7341,N_6648,N_6751);
nor U7342 (N_7342,N_6623,N_6549);
and U7343 (N_7343,N_6604,N_6528);
nand U7344 (N_7344,N_6878,N_6682);
nand U7345 (N_7345,N_6904,N_6606);
and U7346 (N_7346,N_6911,N_6828);
nand U7347 (N_7347,N_6907,N_6659);
nor U7348 (N_7348,N_6535,N_6891);
xor U7349 (N_7349,N_6541,N_6586);
or U7350 (N_7350,N_6658,N_6950);
and U7351 (N_7351,N_6790,N_6970);
or U7352 (N_7352,N_6546,N_6825);
xnor U7353 (N_7353,N_6879,N_6643);
xnor U7354 (N_7354,N_6971,N_6754);
xor U7355 (N_7355,N_6940,N_6989);
xor U7356 (N_7356,N_6588,N_6875);
and U7357 (N_7357,N_6910,N_6629);
and U7358 (N_7358,N_6846,N_6792);
nand U7359 (N_7359,N_6698,N_6500);
or U7360 (N_7360,N_6806,N_6954);
nand U7361 (N_7361,N_6601,N_6510);
nand U7362 (N_7362,N_6556,N_6968);
and U7363 (N_7363,N_6971,N_6550);
nand U7364 (N_7364,N_6808,N_6538);
and U7365 (N_7365,N_6944,N_6963);
or U7366 (N_7366,N_6856,N_6874);
nor U7367 (N_7367,N_6524,N_6871);
nand U7368 (N_7368,N_6850,N_6645);
nand U7369 (N_7369,N_6771,N_6818);
nand U7370 (N_7370,N_6593,N_6597);
nor U7371 (N_7371,N_6862,N_6701);
or U7372 (N_7372,N_6729,N_6610);
or U7373 (N_7373,N_6970,N_6943);
nand U7374 (N_7374,N_6603,N_6771);
and U7375 (N_7375,N_6919,N_6852);
nor U7376 (N_7376,N_6825,N_6998);
or U7377 (N_7377,N_6836,N_6825);
xnor U7378 (N_7378,N_6818,N_6917);
xor U7379 (N_7379,N_6666,N_6663);
nand U7380 (N_7380,N_6622,N_6603);
or U7381 (N_7381,N_6791,N_6586);
xor U7382 (N_7382,N_6874,N_6825);
xor U7383 (N_7383,N_6783,N_6690);
nor U7384 (N_7384,N_6660,N_6959);
or U7385 (N_7385,N_6595,N_6983);
or U7386 (N_7386,N_6979,N_6915);
xor U7387 (N_7387,N_6634,N_6915);
or U7388 (N_7388,N_6588,N_6908);
and U7389 (N_7389,N_6691,N_6617);
nor U7390 (N_7390,N_6795,N_6810);
nand U7391 (N_7391,N_6965,N_6610);
or U7392 (N_7392,N_6870,N_6913);
xor U7393 (N_7393,N_6858,N_6838);
xor U7394 (N_7394,N_6837,N_6500);
or U7395 (N_7395,N_6963,N_6684);
nor U7396 (N_7396,N_6630,N_6991);
nor U7397 (N_7397,N_6971,N_6983);
nor U7398 (N_7398,N_6638,N_6799);
nand U7399 (N_7399,N_6632,N_6884);
xnor U7400 (N_7400,N_6794,N_6581);
xor U7401 (N_7401,N_6657,N_6960);
nand U7402 (N_7402,N_6766,N_6503);
or U7403 (N_7403,N_6708,N_6830);
or U7404 (N_7404,N_6979,N_6936);
and U7405 (N_7405,N_6879,N_6560);
nor U7406 (N_7406,N_6775,N_6532);
xor U7407 (N_7407,N_6628,N_6917);
nor U7408 (N_7408,N_6777,N_6738);
xnor U7409 (N_7409,N_6672,N_6510);
nor U7410 (N_7410,N_6549,N_6657);
nor U7411 (N_7411,N_6822,N_6813);
xor U7412 (N_7412,N_6942,N_6934);
nor U7413 (N_7413,N_6708,N_6605);
xor U7414 (N_7414,N_6825,N_6601);
xnor U7415 (N_7415,N_6746,N_6970);
or U7416 (N_7416,N_6821,N_6534);
or U7417 (N_7417,N_6599,N_6656);
nor U7418 (N_7418,N_6531,N_6507);
nand U7419 (N_7419,N_6944,N_6626);
and U7420 (N_7420,N_6540,N_6915);
nor U7421 (N_7421,N_6620,N_6796);
and U7422 (N_7422,N_6849,N_6574);
xor U7423 (N_7423,N_6717,N_6830);
nand U7424 (N_7424,N_6553,N_6759);
and U7425 (N_7425,N_6775,N_6829);
xnor U7426 (N_7426,N_6758,N_6764);
nand U7427 (N_7427,N_6509,N_6517);
and U7428 (N_7428,N_6861,N_6963);
and U7429 (N_7429,N_6536,N_6735);
xnor U7430 (N_7430,N_6565,N_6794);
nand U7431 (N_7431,N_6930,N_6848);
xor U7432 (N_7432,N_6787,N_6677);
nor U7433 (N_7433,N_6889,N_6784);
nand U7434 (N_7434,N_6518,N_6798);
nand U7435 (N_7435,N_6981,N_6735);
or U7436 (N_7436,N_6929,N_6617);
nand U7437 (N_7437,N_6717,N_6800);
nand U7438 (N_7438,N_6778,N_6962);
nand U7439 (N_7439,N_6652,N_6979);
or U7440 (N_7440,N_6528,N_6993);
nand U7441 (N_7441,N_6889,N_6702);
nor U7442 (N_7442,N_6806,N_6570);
or U7443 (N_7443,N_6737,N_6520);
and U7444 (N_7444,N_6723,N_6775);
or U7445 (N_7445,N_6749,N_6843);
nor U7446 (N_7446,N_6569,N_6665);
xnor U7447 (N_7447,N_6842,N_6535);
or U7448 (N_7448,N_6898,N_6969);
xnor U7449 (N_7449,N_6735,N_6639);
nand U7450 (N_7450,N_6581,N_6734);
or U7451 (N_7451,N_6820,N_6626);
xor U7452 (N_7452,N_6654,N_6533);
nand U7453 (N_7453,N_6586,N_6898);
xnor U7454 (N_7454,N_6512,N_6805);
nand U7455 (N_7455,N_6985,N_6983);
xnor U7456 (N_7456,N_6822,N_6582);
or U7457 (N_7457,N_6828,N_6708);
and U7458 (N_7458,N_6971,N_6647);
and U7459 (N_7459,N_6992,N_6586);
nand U7460 (N_7460,N_6598,N_6554);
or U7461 (N_7461,N_6560,N_6911);
or U7462 (N_7462,N_6726,N_6781);
nor U7463 (N_7463,N_6776,N_6620);
nor U7464 (N_7464,N_6667,N_6827);
nor U7465 (N_7465,N_6634,N_6676);
nand U7466 (N_7466,N_6868,N_6544);
and U7467 (N_7467,N_6915,N_6789);
nand U7468 (N_7468,N_6580,N_6533);
nor U7469 (N_7469,N_6781,N_6755);
nor U7470 (N_7470,N_6555,N_6539);
or U7471 (N_7471,N_6998,N_6956);
xnor U7472 (N_7472,N_6904,N_6842);
xor U7473 (N_7473,N_6819,N_6786);
nor U7474 (N_7474,N_6926,N_6583);
or U7475 (N_7475,N_6568,N_6803);
nand U7476 (N_7476,N_6796,N_6537);
xor U7477 (N_7477,N_6804,N_6706);
or U7478 (N_7478,N_6531,N_6675);
xnor U7479 (N_7479,N_6843,N_6693);
xnor U7480 (N_7480,N_6675,N_6772);
and U7481 (N_7481,N_6934,N_6927);
and U7482 (N_7482,N_6571,N_6553);
xnor U7483 (N_7483,N_6873,N_6710);
xor U7484 (N_7484,N_6965,N_6698);
nor U7485 (N_7485,N_6854,N_6509);
nor U7486 (N_7486,N_6682,N_6697);
xor U7487 (N_7487,N_6920,N_6970);
nand U7488 (N_7488,N_6875,N_6904);
and U7489 (N_7489,N_6545,N_6957);
xnor U7490 (N_7490,N_6771,N_6543);
xor U7491 (N_7491,N_6605,N_6730);
nand U7492 (N_7492,N_6760,N_6534);
nand U7493 (N_7493,N_6801,N_6679);
or U7494 (N_7494,N_6595,N_6674);
xor U7495 (N_7495,N_6822,N_6866);
nor U7496 (N_7496,N_6889,N_6831);
xor U7497 (N_7497,N_6944,N_6586);
nor U7498 (N_7498,N_6734,N_6960);
xor U7499 (N_7499,N_6536,N_6655);
xor U7500 (N_7500,N_7171,N_7216);
and U7501 (N_7501,N_7338,N_7007);
and U7502 (N_7502,N_7210,N_7089);
or U7503 (N_7503,N_7199,N_7107);
nor U7504 (N_7504,N_7293,N_7339);
nor U7505 (N_7505,N_7173,N_7077);
xnor U7506 (N_7506,N_7270,N_7308);
or U7507 (N_7507,N_7424,N_7140);
or U7508 (N_7508,N_7434,N_7301);
xor U7509 (N_7509,N_7200,N_7048);
and U7510 (N_7510,N_7175,N_7486);
nand U7511 (N_7511,N_7069,N_7119);
or U7512 (N_7512,N_7287,N_7294);
nand U7513 (N_7513,N_7458,N_7031);
and U7514 (N_7514,N_7192,N_7162);
and U7515 (N_7515,N_7215,N_7159);
and U7516 (N_7516,N_7321,N_7017);
or U7517 (N_7517,N_7496,N_7419);
xor U7518 (N_7518,N_7076,N_7320);
nand U7519 (N_7519,N_7278,N_7036);
xnor U7520 (N_7520,N_7473,N_7422);
or U7521 (N_7521,N_7435,N_7326);
nor U7522 (N_7522,N_7472,N_7292);
nand U7523 (N_7523,N_7023,N_7030);
and U7524 (N_7524,N_7291,N_7327);
nand U7525 (N_7525,N_7380,N_7393);
or U7526 (N_7526,N_7426,N_7351);
nor U7527 (N_7527,N_7300,N_7334);
or U7528 (N_7528,N_7405,N_7433);
nor U7529 (N_7529,N_7239,N_7184);
xnor U7530 (N_7530,N_7206,N_7428);
or U7531 (N_7531,N_7283,N_7260);
and U7532 (N_7532,N_7230,N_7440);
or U7533 (N_7533,N_7363,N_7147);
xnor U7534 (N_7534,N_7022,N_7432);
and U7535 (N_7535,N_7325,N_7382);
xor U7536 (N_7536,N_7404,N_7064);
and U7537 (N_7537,N_7138,N_7059);
nor U7538 (N_7538,N_7305,N_7438);
nor U7539 (N_7539,N_7085,N_7176);
or U7540 (N_7540,N_7224,N_7461);
nand U7541 (N_7541,N_7477,N_7005);
and U7542 (N_7542,N_7103,N_7227);
and U7543 (N_7543,N_7256,N_7333);
or U7544 (N_7544,N_7034,N_7324);
or U7545 (N_7545,N_7221,N_7483);
nor U7546 (N_7546,N_7011,N_7487);
xnor U7547 (N_7547,N_7371,N_7243);
nand U7548 (N_7548,N_7386,N_7248);
xnor U7549 (N_7549,N_7387,N_7273);
xor U7550 (N_7550,N_7266,N_7112);
and U7551 (N_7551,N_7302,N_7006);
nor U7552 (N_7552,N_7337,N_7254);
and U7553 (N_7553,N_7235,N_7049);
nor U7554 (N_7554,N_7368,N_7236);
or U7555 (N_7555,N_7106,N_7410);
and U7556 (N_7556,N_7413,N_7141);
xnor U7557 (N_7557,N_7484,N_7360);
and U7558 (N_7558,N_7051,N_7355);
and U7559 (N_7559,N_7272,N_7123);
and U7560 (N_7560,N_7403,N_7361);
nor U7561 (N_7561,N_7038,N_7412);
nand U7562 (N_7562,N_7460,N_7429);
or U7563 (N_7563,N_7309,N_7252);
nand U7564 (N_7564,N_7242,N_7479);
nor U7565 (N_7565,N_7449,N_7166);
nor U7566 (N_7566,N_7381,N_7280);
nand U7567 (N_7567,N_7485,N_7349);
nor U7568 (N_7568,N_7350,N_7116);
nor U7569 (N_7569,N_7060,N_7198);
and U7570 (N_7570,N_7401,N_7229);
nand U7571 (N_7571,N_7374,N_7190);
nor U7572 (N_7572,N_7331,N_7201);
xor U7573 (N_7573,N_7055,N_7269);
xnor U7574 (N_7574,N_7417,N_7398);
xnor U7575 (N_7575,N_7388,N_7154);
or U7576 (N_7576,N_7369,N_7411);
xnor U7577 (N_7577,N_7084,N_7120);
and U7578 (N_7578,N_7126,N_7491);
nand U7579 (N_7579,N_7421,N_7058);
xor U7580 (N_7580,N_7096,N_7376);
nor U7581 (N_7581,N_7191,N_7267);
nor U7582 (N_7582,N_7319,N_7020);
and U7583 (N_7583,N_7307,N_7197);
xnor U7584 (N_7584,N_7347,N_7204);
nor U7585 (N_7585,N_7218,N_7439);
xnor U7586 (N_7586,N_7183,N_7033);
xnor U7587 (N_7587,N_7013,N_7447);
and U7588 (N_7588,N_7169,N_7233);
xnor U7589 (N_7589,N_7246,N_7277);
and U7590 (N_7590,N_7443,N_7097);
nor U7591 (N_7591,N_7039,N_7346);
and U7592 (N_7592,N_7019,N_7232);
and U7593 (N_7593,N_7137,N_7041);
nor U7594 (N_7594,N_7214,N_7322);
nand U7595 (N_7595,N_7026,N_7481);
nand U7596 (N_7596,N_7099,N_7299);
nand U7597 (N_7597,N_7488,N_7075);
and U7598 (N_7598,N_7002,N_7179);
xor U7599 (N_7599,N_7185,N_7465);
and U7600 (N_7600,N_7336,N_7222);
or U7601 (N_7601,N_7394,N_7452);
nand U7602 (N_7602,N_7047,N_7152);
xor U7603 (N_7603,N_7091,N_7202);
nand U7604 (N_7604,N_7040,N_7430);
nand U7605 (N_7605,N_7037,N_7257);
nand U7606 (N_7606,N_7046,N_7455);
nand U7607 (N_7607,N_7415,N_7148);
and U7608 (N_7608,N_7027,N_7454);
xnor U7609 (N_7609,N_7332,N_7024);
or U7610 (N_7610,N_7219,N_7207);
or U7611 (N_7611,N_7328,N_7043);
nand U7612 (N_7612,N_7108,N_7220);
or U7613 (N_7613,N_7001,N_7493);
or U7614 (N_7614,N_7258,N_7470);
xnor U7615 (N_7615,N_7312,N_7110);
nand U7616 (N_7616,N_7193,N_7251);
and U7617 (N_7617,N_7244,N_7015);
nand U7618 (N_7618,N_7318,N_7478);
or U7619 (N_7619,N_7445,N_7181);
nor U7620 (N_7620,N_7453,N_7155);
or U7621 (N_7621,N_7276,N_7095);
or U7622 (N_7622,N_7052,N_7102);
and U7623 (N_7623,N_7090,N_7054);
and U7624 (N_7624,N_7344,N_7298);
xnor U7625 (N_7625,N_7436,N_7143);
and U7626 (N_7626,N_7245,N_7028);
nand U7627 (N_7627,N_7129,N_7228);
or U7628 (N_7628,N_7264,N_7286);
nand U7629 (N_7629,N_7446,N_7170);
nor U7630 (N_7630,N_7208,N_7342);
xnor U7631 (N_7631,N_7203,N_7340);
or U7632 (N_7632,N_7158,N_7035);
or U7633 (N_7633,N_7275,N_7092);
nand U7634 (N_7634,N_7008,N_7495);
nand U7635 (N_7635,N_7456,N_7250);
nor U7636 (N_7636,N_7464,N_7468);
nand U7637 (N_7637,N_7098,N_7128);
nor U7638 (N_7638,N_7385,N_7407);
or U7639 (N_7639,N_7157,N_7408);
nand U7640 (N_7640,N_7062,N_7330);
and U7641 (N_7641,N_7414,N_7010);
nor U7642 (N_7642,N_7187,N_7072);
nand U7643 (N_7643,N_7124,N_7442);
and U7644 (N_7644,N_7297,N_7127);
xnor U7645 (N_7645,N_7056,N_7014);
nor U7646 (N_7646,N_7271,N_7313);
nor U7647 (N_7647,N_7262,N_7114);
and U7648 (N_7648,N_7066,N_7253);
xnor U7649 (N_7649,N_7079,N_7012);
xnor U7650 (N_7650,N_7492,N_7153);
nor U7651 (N_7651,N_7150,N_7463);
nor U7652 (N_7652,N_7149,N_7316);
nand U7653 (N_7653,N_7373,N_7156);
xor U7654 (N_7654,N_7018,N_7145);
and U7655 (N_7655,N_7132,N_7000);
nor U7656 (N_7656,N_7306,N_7070);
nand U7657 (N_7657,N_7133,N_7209);
xor U7658 (N_7658,N_7282,N_7343);
nand U7659 (N_7659,N_7469,N_7462);
or U7660 (N_7660,N_7021,N_7101);
and U7661 (N_7661,N_7115,N_7279);
and U7662 (N_7662,N_7080,N_7451);
or U7663 (N_7663,N_7431,N_7480);
or U7664 (N_7664,N_7423,N_7418);
nor U7665 (N_7665,N_7094,N_7093);
and U7666 (N_7666,N_7378,N_7466);
and U7667 (N_7667,N_7081,N_7392);
or U7668 (N_7668,N_7188,N_7139);
and U7669 (N_7669,N_7310,N_7196);
nand U7670 (N_7670,N_7335,N_7240);
nand U7671 (N_7671,N_7044,N_7263);
nor U7672 (N_7672,N_7359,N_7444);
nand U7673 (N_7673,N_7100,N_7131);
nor U7674 (N_7674,N_7261,N_7061);
nand U7675 (N_7675,N_7195,N_7180);
nor U7676 (N_7676,N_7238,N_7074);
and U7677 (N_7677,N_7471,N_7255);
nand U7678 (N_7678,N_7078,N_7315);
and U7679 (N_7679,N_7177,N_7354);
nand U7680 (N_7680,N_7281,N_7174);
or U7681 (N_7681,N_7068,N_7163);
xnor U7682 (N_7682,N_7135,N_7009);
or U7683 (N_7683,N_7379,N_7314);
nand U7684 (N_7684,N_7004,N_7104);
xnor U7685 (N_7685,N_7105,N_7391);
nor U7686 (N_7686,N_7489,N_7358);
xor U7687 (N_7687,N_7241,N_7071);
and U7688 (N_7688,N_7402,N_7372);
nor U7689 (N_7689,N_7247,N_7390);
nand U7690 (N_7690,N_7289,N_7003);
nor U7691 (N_7691,N_7437,N_7370);
or U7692 (N_7692,N_7130,N_7144);
xnor U7693 (N_7693,N_7459,N_7409);
or U7694 (N_7694,N_7448,N_7259);
xnor U7695 (N_7695,N_7285,N_7063);
xnor U7696 (N_7696,N_7395,N_7383);
or U7697 (N_7697,N_7161,N_7441);
nand U7698 (N_7698,N_7189,N_7213);
and U7699 (N_7699,N_7311,N_7366);
xor U7700 (N_7700,N_7288,N_7226);
or U7701 (N_7701,N_7249,N_7353);
nor U7702 (N_7702,N_7474,N_7499);
or U7703 (N_7703,N_7268,N_7352);
nor U7704 (N_7704,N_7136,N_7290);
nand U7705 (N_7705,N_7025,N_7329);
and U7706 (N_7706,N_7475,N_7057);
xor U7707 (N_7707,N_7406,N_7323);
and U7708 (N_7708,N_7142,N_7032);
or U7709 (N_7709,N_7490,N_7303);
xnor U7710 (N_7710,N_7362,N_7476);
nand U7711 (N_7711,N_7164,N_7274);
nand U7712 (N_7712,N_7296,N_7497);
xnor U7713 (N_7713,N_7348,N_7400);
or U7714 (N_7714,N_7117,N_7045);
xnor U7715 (N_7715,N_7086,N_7420);
and U7716 (N_7716,N_7377,N_7029);
xor U7717 (N_7717,N_7494,N_7165);
nor U7718 (N_7718,N_7211,N_7087);
xor U7719 (N_7719,N_7168,N_7167);
xnor U7720 (N_7720,N_7178,N_7088);
and U7721 (N_7721,N_7225,N_7067);
nand U7722 (N_7722,N_7498,N_7304);
and U7723 (N_7723,N_7113,N_7364);
nor U7724 (N_7724,N_7425,N_7186);
or U7725 (N_7725,N_7125,N_7384);
or U7726 (N_7726,N_7151,N_7083);
nor U7727 (N_7727,N_7016,N_7237);
or U7728 (N_7728,N_7050,N_7217);
and U7729 (N_7729,N_7365,N_7284);
xnor U7730 (N_7730,N_7172,N_7345);
xor U7731 (N_7731,N_7053,N_7265);
and U7732 (N_7732,N_7427,N_7122);
or U7733 (N_7733,N_7416,N_7396);
nand U7734 (N_7734,N_7367,N_7205);
or U7735 (N_7735,N_7118,N_7356);
nor U7736 (N_7736,N_7467,N_7317);
xor U7737 (N_7737,N_7223,N_7357);
and U7738 (N_7738,N_7389,N_7194);
nand U7739 (N_7739,N_7134,N_7450);
nand U7740 (N_7740,N_7111,N_7065);
nor U7741 (N_7741,N_7182,N_7160);
nor U7742 (N_7742,N_7399,N_7121);
nor U7743 (N_7743,N_7082,N_7375);
xor U7744 (N_7744,N_7457,N_7146);
nor U7745 (N_7745,N_7212,N_7341);
or U7746 (N_7746,N_7042,N_7234);
nand U7747 (N_7747,N_7397,N_7482);
nor U7748 (N_7748,N_7295,N_7231);
or U7749 (N_7749,N_7109,N_7073);
xor U7750 (N_7750,N_7194,N_7254);
and U7751 (N_7751,N_7248,N_7258);
xnor U7752 (N_7752,N_7400,N_7281);
and U7753 (N_7753,N_7293,N_7370);
and U7754 (N_7754,N_7315,N_7125);
or U7755 (N_7755,N_7205,N_7141);
and U7756 (N_7756,N_7202,N_7339);
nor U7757 (N_7757,N_7081,N_7397);
or U7758 (N_7758,N_7114,N_7057);
xor U7759 (N_7759,N_7277,N_7197);
and U7760 (N_7760,N_7367,N_7081);
nor U7761 (N_7761,N_7155,N_7021);
nor U7762 (N_7762,N_7124,N_7128);
nor U7763 (N_7763,N_7359,N_7272);
nand U7764 (N_7764,N_7254,N_7448);
nand U7765 (N_7765,N_7270,N_7448);
nor U7766 (N_7766,N_7344,N_7072);
nor U7767 (N_7767,N_7238,N_7287);
nor U7768 (N_7768,N_7216,N_7358);
and U7769 (N_7769,N_7210,N_7147);
nand U7770 (N_7770,N_7232,N_7365);
and U7771 (N_7771,N_7243,N_7387);
xnor U7772 (N_7772,N_7030,N_7421);
nand U7773 (N_7773,N_7057,N_7312);
and U7774 (N_7774,N_7483,N_7067);
or U7775 (N_7775,N_7408,N_7306);
and U7776 (N_7776,N_7106,N_7284);
or U7777 (N_7777,N_7021,N_7358);
and U7778 (N_7778,N_7254,N_7474);
nand U7779 (N_7779,N_7112,N_7183);
or U7780 (N_7780,N_7256,N_7283);
or U7781 (N_7781,N_7463,N_7142);
or U7782 (N_7782,N_7223,N_7271);
nand U7783 (N_7783,N_7074,N_7291);
nand U7784 (N_7784,N_7008,N_7129);
nor U7785 (N_7785,N_7044,N_7347);
nand U7786 (N_7786,N_7092,N_7217);
xnor U7787 (N_7787,N_7419,N_7144);
nor U7788 (N_7788,N_7415,N_7376);
and U7789 (N_7789,N_7448,N_7029);
nor U7790 (N_7790,N_7402,N_7068);
xnor U7791 (N_7791,N_7420,N_7102);
or U7792 (N_7792,N_7371,N_7014);
nor U7793 (N_7793,N_7255,N_7468);
or U7794 (N_7794,N_7133,N_7061);
and U7795 (N_7795,N_7234,N_7033);
xor U7796 (N_7796,N_7101,N_7475);
and U7797 (N_7797,N_7296,N_7494);
and U7798 (N_7798,N_7408,N_7027);
xor U7799 (N_7799,N_7105,N_7310);
nand U7800 (N_7800,N_7409,N_7371);
nand U7801 (N_7801,N_7395,N_7485);
or U7802 (N_7802,N_7265,N_7481);
nor U7803 (N_7803,N_7142,N_7248);
or U7804 (N_7804,N_7009,N_7386);
xor U7805 (N_7805,N_7373,N_7392);
and U7806 (N_7806,N_7441,N_7098);
and U7807 (N_7807,N_7055,N_7235);
and U7808 (N_7808,N_7060,N_7112);
or U7809 (N_7809,N_7490,N_7210);
nor U7810 (N_7810,N_7318,N_7291);
and U7811 (N_7811,N_7338,N_7429);
xnor U7812 (N_7812,N_7186,N_7307);
or U7813 (N_7813,N_7227,N_7143);
or U7814 (N_7814,N_7469,N_7151);
xnor U7815 (N_7815,N_7014,N_7025);
or U7816 (N_7816,N_7487,N_7110);
nand U7817 (N_7817,N_7142,N_7268);
or U7818 (N_7818,N_7339,N_7058);
xor U7819 (N_7819,N_7116,N_7249);
or U7820 (N_7820,N_7406,N_7421);
or U7821 (N_7821,N_7496,N_7126);
nand U7822 (N_7822,N_7163,N_7388);
xor U7823 (N_7823,N_7203,N_7416);
and U7824 (N_7824,N_7062,N_7435);
xnor U7825 (N_7825,N_7283,N_7118);
and U7826 (N_7826,N_7136,N_7068);
and U7827 (N_7827,N_7010,N_7451);
and U7828 (N_7828,N_7297,N_7383);
nor U7829 (N_7829,N_7366,N_7217);
xnor U7830 (N_7830,N_7242,N_7430);
or U7831 (N_7831,N_7391,N_7189);
or U7832 (N_7832,N_7090,N_7473);
nand U7833 (N_7833,N_7123,N_7075);
and U7834 (N_7834,N_7475,N_7384);
nor U7835 (N_7835,N_7156,N_7102);
nand U7836 (N_7836,N_7106,N_7172);
and U7837 (N_7837,N_7490,N_7497);
xor U7838 (N_7838,N_7395,N_7075);
nand U7839 (N_7839,N_7467,N_7361);
nand U7840 (N_7840,N_7140,N_7366);
and U7841 (N_7841,N_7334,N_7143);
xnor U7842 (N_7842,N_7048,N_7039);
nand U7843 (N_7843,N_7221,N_7325);
nand U7844 (N_7844,N_7228,N_7067);
nor U7845 (N_7845,N_7230,N_7207);
xnor U7846 (N_7846,N_7406,N_7180);
and U7847 (N_7847,N_7323,N_7079);
xnor U7848 (N_7848,N_7010,N_7246);
nor U7849 (N_7849,N_7255,N_7473);
or U7850 (N_7850,N_7239,N_7408);
nor U7851 (N_7851,N_7267,N_7498);
nand U7852 (N_7852,N_7054,N_7093);
and U7853 (N_7853,N_7490,N_7153);
nor U7854 (N_7854,N_7486,N_7279);
xor U7855 (N_7855,N_7025,N_7175);
xor U7856 (N_7856,N_7006,N_7401);
and U7857 (N_7857,N_7040,N_7202);
and U7858 (N_7858,N_7036,N_7293);
nand U7859 (N_7859,N_7367,N_7287);
or U7860 (N_7860,N_7004,N_7484);
xor U7861 (N_7861,N_7014,N_7078);
or U7862 (N_7862,N_7261,N_7099);
nor U7863 (N_7863,N_7162,N_7002);
or U7864 (N_7864,N_7213,N_7046);
or U7865 (N_7865,N_7136,N_7001);
or U7866 (N_7866,N_7153,N_7484);
or U7867 (N_7867,N_7243,N_7372);
and U7868 (N_7868,N_7314,N_7466);
and U7869 (N_7869,N_7153,N_7489);
xor U7870 (N_7870,N_7436,N_7004);
xnor U7871 (N_7871,N_7347,N_7334);
or U7872 (N_7872,N_7396,N_7334);
xnor U7873 (N_7873,N_7315,N_7211);
nand U7874 (N_7874,N_7249,N_7437);
or U7875 (N_7875,N_7249,N_7454);
or U7876 (N_7876,N_7289,N_7119);
and U7877 (N_7877,N_7376,N_7139);
and U7878 (N_7878,N_7402,N_7239);
and U7879 (N_7879,N_7448,N_7372);
xnor U7880 (N_7880,N_7380,N_7345);
or U7881 (N_7881,N_7035,N_7180);
and U7882 (N_7882,N_7420,N_7052);
or U7883 (N_7883,N_7490,N_7187);
nor U7884 (N_7884,N_7341,N_7345);
or U7885 (N_7885,N_7189,N_7277);
xnor U7886 (N_7886,N_7174,N_7241);
or U7887 (N_7887,N_7146,N_7278);
and U7888 (N_7888,N_7367,N_7442);
nand U7889 (N_7889,N_7162,N_7016);
xor U7890 (N_7890,N_7356,N_7280);
nand U7891 (N_7891,N_7281,N_7444);
and U7892 (N_7892,N_7244,N_7434);
nand U7893 (N_7893,N_7413,N_7132);
xor U7894 (N_7894,N_7058,N_7369);
xnor U7895 (N_7895,N_7424,N_7030);
xor U7896 (N_7896,N_7444,N_7439);
or U7897 (N_7897,N_7494,N_7088);
and U7898 (N_7898,N_7438,N_7207);
or U7899 (N_7899,N_7417,N_7468);
nor U7900 (N_7900,N_7074,N_7213);
or U7901 (N_7901,N_7285,N_7211);
and U7902 (N_7902,N_7395,N_7000);
or U7903 (N_7903,N_7062,N_7468);
or U7904 (N_7904,N_7197,N_7407);
xnor U7905 (N_7905,N_7328,N_7275);
and U7906 (N_7906,N_7393,N_7331);
xnor U7907 (N_7907,N_7295,N_7135);
or U7908 (N_7908,N_7342,N_7439);
and U7909 (N_7909,N_7441,N_7111);
nor U7910 (N_7910,N_7193,N_7188);
or U7911 (N_7911,N_7311,N_7292);
and U7912 (N_7912,N_7436,N_7364);
nand U7913 (N_7913,N_7012,N_7085);
or U7914 (N_7914,N_7316,N_7158);
or U7915 (N_7915,N_7054,N_7466);
nor U7916 (N_7916,N_7179,N_7314);
nor U7917 (N_7917,N_7277,N_7403);
nand U7918 (N_7918,N_7482,N_7391);
or U7919 (N_7919,N_7208,N_7228);
and U7920 (N_7920,N_7299,N_7029);
xor U7921 (N_7921,N_7300,N_7412);
and U7922 (N_7922,N_7194,N_7441);
nor U7923 (N_7923,N_7195,N_7487);
or U7924 (N_7924,N_7402,N_7158);
nor U7925 (N_7925,N_7184,N_7236);
xnor U7926 (N_7926,N_7293,N_7067);
and U7927 (N_7927,N_7114,N_7468);
and U7928 (N_7928,N_7325,N_7050);
or U7929 (N_7929,N_7345,N_7370);
or U7930 (N_7930,N_7180,N_7040);
xor U7931 (N_7931,N_7300,N_7167);
xnor U7932 (N_7932,N_7332,N_7476);
nand U7933 (N_7933,N_7372,N_7489);
or U7934 (N_7934,N_7405,N_7057);
or U7935 (N_7935,N_7346,N_7415);
nor U7936 (N_7936,N_7055,N_7232);
xor U7937 (N_7937,N_7183,N_7255);
xnor U7938 (N_7938,N_7333,N_7056);
nor U7939 (N_7939,N_7299,N_7399);
or U7940 (N_7940,N_7083,N_7262);
or U7941 (N_7941,N_7220,N_7322);
xor U7942 (N_7942,N_7071,N_7370);
and U7943 (N_7943,N_7050,N_7135);
or U7944 (N_7944,N_7159,N_7354);
and U7945 (N_7945,N_7142,N_7051);
nand U7946 (N_7946,N_7273,N_7170);
xor U7947 (N_7947,N_7129,N_7070);
and U7948 (N_7948,N_7246,N_7327);
xor U7949 (N_7949,N_7422,N_7224);
xnor U7950 (N_7950,N_7128,N_7384);
xnor U7951 (N_7951,N_7268,N_7094);
nand U7952 (N_7952,N_7479,N_7395);
or U7953 (N_7953,N_7114,N_7340);
xor U7954 (N_7954,N_7182,N_7013);
nand U7955 (N_7955,N_7172,N_7157);
or U7956 (N_7956,N_7343,N_7441);
nand U7957 (N_7957,N_7352,N_7291);
nand U7958 (N_7958,N_7375,N_7113);
nand U7959 (N_7959,N_7262,N_7115);
nor U7960 (N_7960,N_7044,N_7199);
or U7961 (N_7961,N_7348,N_7095);
or U7962 (N_7962,N_7118,N_7420);
nand U7963 (N_7963,N_7231,N_7046);
nand U7964 (N_7964,N_7483,N_7090);
nand U7965 (N_7965,N_7235,N_7397);
nand U7966 (N_7966,N_7169,N_7153);
xor U7967 (N_7967,N_7467,N_7316);
nor U7968 (N_7968,N_7468,N_7192);
nand U7969 (N_7969,N_7203,N_7328);
and U7970 (N_7970,N_7140,N_7066);
and U7971 (N_7971,N_7321,N_7075);
or U7972 (N_7972,N_7385,N_7121);
or U7973 (N_7973,N_7332,N_7430);
nand U7974 (N_7974,N_7139,N_7337);
nor U7975 (N_7975,N_7475,N_7059);
or U7976 (N_7976,N_7273,N_7253);
xnor U7977 (N_7977,N_7352,N_7497);
nand U7978 (N_7978,N_7054,N_7186);
and U7979 (N_7979,N_7180,N_7462);
and U7980 (N_7980,N_7040,N_7361);
xnor U7981 (N_7981,N_7483,N_7025);
or U7982 (N_7982,N_7174,N_7317);
nand U7983 (N_7983,N_7186,N_7409);
nor U7984 (N_7984,N_7066,N_7008);
or U7985 (N_7985,N_7393,N_7091);
nor U7986 (N_7986,N_7088,N_7471);
and U7987 (N_7987,N_7254,N_7032);
xor U7988 (N_7988,N_7059,N_7062);
xnor U7989 (N_7989,N_7442,N_7425);
nor U7990 (N_7990,N_7086,N_7255);
and U7991 (N_7991,N_7327,N_7082);
or U7992 (N_7992,N_7206,N_7252);
nand U7993 (N_7993,N_7445,N_7104);
or U7994 (N_7994,N_7265,N_7344);
and U7995 (N_7995,N_7393,N_7031);
nor U7996 (N_7996,N_7400,N_7128);
or U7997 (N_7997,N_7100,N_7388);
nand U7998 (N_7998,N_7170,N_7464);
nor U7999 (N_7999,N_7199,N_7010);
nand U8000 (N_8000,N_7713,N_7577);
or U8001 (N_8001,N_7503,N_7761);
or U8002 (N_8002,N_7900,N_7770);
and U8003 (N_8003,N_7757,N_7815);
and U8004 (N_8004,N_7879,N_7665);
nor U8005 (N_8005,N_7931,N_7691);
xor U8006 (N_8006,N_7964,N_7942);
and U8007 (N_8007,N_7801,N_7715);
nand U8008 (N_8008,N_7819,N_7637);
nand U8009 (N_8009,N_7976,N_7929);
nor U8010 (N_8010,N_7889,N_7974);
xnor U8011 (N_8011,N_7887,N_7808);
xor U8012 (N_8012,N_7753,N_7543);
and U8013 (N_8013,N_7697,N_7988);
nand U8014 (N_8014,N_7528,N_7636);
nor U8015 (N_8015,N_7863,N_7935);
and U8016 (N_8016,N_7648,N_7828);
nand U8017 (N_8017,N_7594,N_7998);
nand U8018 (N_8018,N_7811,N_7807);
nor U8019 (N_8019,N_7597,N_7975);
or U8020 (N_8020,N_7512,N_7766);
nand U8021 (N_8021,N_7778,N_7871);
xor U8022 (N_8022,N_7690,N_7686);
nor U8023 (N_8023,N_7705,N_7995);
nor U8024 (N_8024,N_7752,N_7954);
nor U8025 (N_8025,N_7769,N_7525);
or U8026 (N_8026,N_7742,N_7728);
xnor U8027 (N_8027,N_7953,N_7551);
and U8028 (N_8028,N_7773,N_7714);
or U8029 (N_8029,N_7788,N_7751);
xnor U8030 (N_8030,N_7703,N_7673);
nand U8031 (N_8031,N_7780,N_7601);
nor U8032 (N_8032,N_7933,N_7843);
nor U8033 (N_8033,N_7687,N_7641);
or U8034 (N_8034,N_7764,N_7603);
nor U8035 (N_8035,N_7642,N_7620);
nor U8036 (N_8036,N_7559,N_7803);
nand U8037 (N_8037,N_7922,N_7930);
nand U8038 (N_8038,N_7650,N_7702);
nand U8039 (N_8039,N_7891,N_7746);
xnor U8040 (N_8040,N_7804,N_7578);
nand U8041 (N_8041,N_7692,N_7509);
nand U8042 (N_8042,N_7882,N_7548);
nor U8043 (N_8043,N_7963,N_7631);
and U8044 (N_8044,N_7500,N_7827);
xor U8045 (N_8045,N_7689,N_7937);
nor U8046 (N_8046,N_7730,N_7771);
nand U8047 (N_8047,N_7793,N_7888);
nand U8048 (N_8048,N_7736,N_7608);
nor U8049 (N_8049,N_7750,N_7949);
or U8050 (N_8050,N_7915,N_7894);
xnor U8051 (N_8051,N_7950,N_7600);
or U8052 (N_8052,N_7864,N_7607);
nand U8053 (N_8053,N_7540,N_7639);
nand U8054 (N_8054,N_7881,N_7716);
and U8055 (N_8055,N_7992,N_7623);
nand U8056 (N_8056,N_7850,N_7836);
nor U8057 (N_8057,N_7745,N_7831);
or U8058 (N_8058,N_7982,N_7837);
nand U8059 (N_8059,N_7779,N_7554);
nor U8060 (N_8060,N_7638,N_7524);
nor U8061 (N_8061,N_7602,N_7846);
or U8062 (N_8062,N_7535,N_7966);
and U8063 (N_8063,N_7901,N_7725);
xnor U8064 (N_8064,N_7852,N_7660);
nand U8065 (N_8065,N_7994,N_7531);
nor U8066 (N_8066,N_7786,N_7777);
nor U8067 (N_8067,N_7980,N_7977);
or U8068 (N_8068,N_7918,N_7979);
or U8069 (N_8069,N_7644,N_7719);
xnor U8070 (N_8070,N_7829,N_7563);
nor U8071 (N_8071,N_7762,N_7823);
or U8072 (N_8072,N_7606,N_7544);
nand U8073 (N_8073,N_7567,N_7549);
nand U8074 (N_8074,N_7885,N_7868);
or U8075 (N_8075,N_7957,N_7877);
xor U8076 (N_8076,N_7667,N_7883);
or U8077 (N_8077,N_7955,N_7855);
or U8078 (N_8078,N_7694,N_7721);
xor U8079 (N_8079,N_7537,N_7743);
nor U8080 (N_8080,N_7583,N_7903);
nand U8081 (N_8081,N_7755,N_7800);
nand U8082 (N_8082,N_7990,N_7926);
nand U8083 (N_8083,N_7890,N_7685);
and U8084 (N_8084,N_7521,N_7765);
nand U8085 (N_8085,N_7586,N_7802);
or U8086 (N_8086,N_7997,N_7860);
nor U8087 (N_8087,N_7612,N_7813);
nand U8088 (N_8088,N_7569,N_7566);
xnor U8089 (N_8089,N_7814,N_7904);
xnor U8090 (N_8090,N_7529,N_7984);
or U8091 (N_8091,N_7859,N_7733);
and U8092 (N_8092,N_7640,N_7884);
or U8093 (N_8093,N_7661,N_7940);
xnor U8094 (N_8094,N_7861,N_7727);
and U8095 (N_8095,N_7785,N_7710);
and U8096 (N_8096,N_7599,N_7739);
or U8097 (N_8097,N_7731,N_7522);
xnor U8098 (N_8098,N_7848,N_7987);
or U8099 (N_8099,N_7505,N_7649);
or U8100 (N_8100,N_7585,N_7670);
xnor U8101 (N_8101,N_7767,N_7820);
nor U8102 (N_8102,N_7527,N_7656);
nand U8103 (N_8103,N_7645,N_7632);
or U8104 (N_8104,N_7874,N_7886);
nor U8105 (N_8105,N_7999,N_7796);
nor U8106 (N_8106,N_7662,N_7504);
nor U8107 (N_8107,N_7619,N_7928);
and U8108 (N_8108,N_7655,N_7943);
xor U8109 (N_8109,N_7911,N_7948);
nor U8110 (N_8110,N_7916,N_7798);
nor U8111 (N_8111,N_7737,N_7782);
xnor U8112 (N_8112,N_7919,N_7774);
or U8113 (N_8113,N_7633,N_7643);
and U8114 (N_8114,N_7701,N_7658);
or U8115 (N_8115,N_7729,N_7553);
and U8116 (N_8116,N_7972,N_7838);
xor U8117 (N_8117,N_7546,N_7986);
or U8118 (N_8118,N_7910,N_7573);
or U8119 (N_8119,N_7945,N_7792);
or U8120 (N_8120,N_7595,N_7867);
nand U8121 (N_8121,N_7565,N_7625);
xor U8122 (N_8122,N_7653,N_7899);
xnor U8123 (N_8123,N_7628,N_7924);
and U8124 (N_8124,N_7555,N_7706);
nor U8125 (N_8125,N_7684,N_7865);
nor U8126 (N_8126,N_7854,N_7818);
nand U8127 (N_8127,N_7993,N_7572);
and U8128 (N_8128,N_7965,N_7672);
or U8129 (N_8129,N_7783,N_7609);
xor U8130 (N_8130,N_7962,N_7968);
and U8131 (N_8131,N_7634,N_7675);
and U8132 (N_8132,N_7647,N_7981);
or U8133 (N_8133,N_7556,N_7961);
or U8134 (N_8134,N_7781,N_7923);
and U8135 (N_8135,N_7635,N_7880);
or U8136 (N_8136,N_7519,N_7760);
xnor U8137 (N_8137,N_7614,N_7741);
nand U8138 (N_8138,N_7873,N_7932);
nand U8139 (N_8139,N_7724,N_7541);
or U8140 (N_8140,N_7946,N_7853);
and U8141 (N_8141,N_7822,N_7756);
xnor U8142 (N_8142,N_7613,N_7723);
xor U8143 (N_8143,N_7832,N_7775);
nor U8144 (N_8144,N_7616,N_7590);
nor U8145 (N_8145,N_7526,N_7789);
nand U8146 (N_8146,N_7562,N_7611);
xor U8147 (N_8147,N_7866,N_7768);
nor U8148 (N_8148,N_7669,N_7561);
nand U8149 (N_8149,N_7699,N_7615);
nand U8150 (N_8150,N_7817,N_7772);
nor U8151 (N_8151,N_7560,N_7671);
xnor U8152 (N_8152,N_7951,N_7726);
nand U8153 (N_8153,N_7794,N_7520);
nand U8154 (N_8154,N_7681,N_7914);
and U8155 (N_8155,N_7542,N_7787);
or U8156 (N_8156,N_7604,N_7576);
xor U8157 (N_8157,N_7844,N_7579);
or U8158 (N_8158,N_7591,N_7530);
or U8159 (N_8159,N_7805,N_7936);
and U8160 (N_8160,N_7759,N_7508);
nand U8161 (N_8161,N_7734,N_7841);
nand U8162 (N_8162,N_7797,N_7533);
xor U8163 (N_8163,N_7516,N_7917);
xor U8164 (N_8164,N_7709,N_7856);
nor U8165 (N_8165,N_7698,N_7664);
nor U8166 (N_8166,N_7680,N_7720);
and U8167 (N_8167,N_7676,N_7896);
and U8168 (N_8168,N_7996,N_7902);
or U8169 (N_8169,N_7791,N_7895);
xor U8170 (N_8170,N_7790,N_7857);
or U8171 (N_8171,N_7679,N_7517);
nor U8172 (N_8172,N_7682,N_7574);
xor U8173 (N_8173,N_7704,N_7515);
xnor U8174 (N_8174,N_7847,N_7589);
nand U8175 (N_8175,N_7826,N_7547);
and U8176 (N_8176,N_7906,N_7845);
nor U8177 (N_8177,N_7592,N_7905);
or U8178 (N_8178,N_7558,N_7744);
nor U8179 (N_8179,N_7907,N_7799);
xor U8180 (N_8180,N_7941,N_7913);
xnor U8181 (N_8181,N_7657,N_7510);
xor U8182 (N_8182,N_7564,N_7959);
nor U8183 (N_8183,N_7858,N_7707);
nor U8184 (N_8184,N_7912,N_7651);
nand U8185 (N_8185,N_7824,N_7587);
xnor U8186 (N_8186,N_7839,N_7830);
and U8187 (N_8187,N_7629,N_7552);
or U8188 (N_8188,N_7501,N_7627);
nor U8189 (N_8189,N_7652,N_7683);
xnor U8190 (N_8190,N_7763,N_7754);
nor U8191 (N_8191,N_7967,N_7654);
nand U8192 (N_8192,N_7518,N_7668);
and U8193 (N_8193,N_7983,N_7758);
xor U8194 (N_8194,N_7740,N_7575);
nor U8195 (N_8195,N_7735,N_7897);
and U8196 (N_8196,N_7545,N_7550);
nand U8197 (N_8197,N_7621,N_7598);
and U8198 (N_8198,N_7538,N_7626);
and U8199 (N_8199,N_7925,N_7816);
xor U8200 (N_8200,N_7666,N_7821);
nand U8201 (N_8201,N_7674,N_7718);
nor U8202 (N_8202,N_7747,N_7971);
or U8203 (N_8203,N_7956,N_7810);
or U8204 (N_8204,N_7610,N_7927);
or U8205 (N_8205,N_7938,N_7809);
or U8206 (N_8206,N_7878,N_7605);
nor U8207 (N_8207,N_7869,N_7557);
and U8208 (N_8208,N_7708,N_7700);
nor U8209 (N_8209,N_7534,N_7842);
or U8210 (N_8210,N_7696,N_7970);
and U8211 (N_8211,N_7588,N_7738);
nor U8212 (N_8212,N_7920,N_7834);
nor U8213 (N_8213,N_7712,N_7944);
nand U8214 (N_8214,N_7711,N_7502);
nand U8215 (N_8215,N_7571,N_7978);
xnor U8216 (N_8216,N_7893,N_7532);
or U8217 (N_8217,N_7622,N_7898);
nand U8218 (N_8218,N_7892,N_7677);
or U8219 (N_8219,N_7851,N_7678);
xnor U8220 (N_8220,N_7973,N_7939);
or U8221 (N_8221,N_7748,N_7833);
nor U8222 (N_8222,N_7875,N_7985);
xor U8223 (N_8223,N_7580,N_7513);
xnor U8224 (N_8224,N_7947,N_7776);
nand U8225 (N_8225,N_7618,N_7870);
or U8226 (N_8226,N_7536,N_7646);
or U8227 (N_8227,N_7630,N_7840);
xnor U8228 (N_8228,N_7795,N_7960);
and U8229 (N_8229,N_7593,N_7688);
xnor U8230 (N_8230,N_7806,N_7876);
xor U8231 (N_8231,N_7624,N_7717);
nor U8232 (N_8232,N_7825,N_7934);
xnor U8233 (N_8233,N_7921,N_7568);
xor U8234 (N_8234,N_7872,N_7969);
xnor U8235 (N_8235,N_7989,N_7581);
nand U8236 (N_8236,N_7659,N_7784);
and U8237 (N_8237,N_7695,N_7570);
or U8238 (N_8238,N_7835,N_7952);
nor U8239 (N_8239,N_7596,N_7582);
xor U8240 (N_8240,N_7511,N_7514);
or U8241 (N_8241,N_7849,N_7812);
and U8242 (N_8242,N_7749,N_7908);
and U8243 (N_8243,N_7722,N_7693);
or U8244 (N_8244,N_7862,N_7991);
xnor U8245 (N_8245,N_7539,N_7506);
and U8246 (N_8246,N_7663,N_7617);
or U8247 (N_8247,N_7909,N_7584);
nor U8248 (N_8248,N_7732,N_7958);
xnor U8249 (N_8249,N_7507,N_7523);
or U8250 (N_8250,N_7506,N_7807);
nand U8251 (N_8251,N_7976,N_7949);
or U8252 (N_8252,N_7777,N_7792);
nand U8253 (N_8253,N_7817,N_7647);
nand U8254 (N_8254,N_7998,N_7500);
and U8255 (N_8255,N_7739,N_7823);
nand U8256 (N_8256,N_7710,N_7755);
nor U8257 (N_8257,N_7529,N_7901);
nor U8258 (N_8258,N_7676,N_7741);
nor U8259 (N_8259,N_7845,N_7923);
nor U8260 (N_8260,N_7798,N_7930);
xnor U8261 (N_8261,N_7966,N_7560);
nor U8262 (N_8262,N_7697,N_7777);
nor U8263 (N_8263,N_7797,N_7815);
nor U8264 (N_8264,N_7653,N_7900);
xor U8265 (N_8265,N_7594,N_7727);
or U8266 (N_8266,N_7849,N_7630);
nor U8267 (N_8267,N_7813,N_7613);
or U8268 (N_8268,N_7822,N_7573);
xor U8269 (N_8269,N_7611,N_7586);
and U8270 (N_8270,N_7761,N_7597);
and U8271 (N_8271,N_7601,N_7954);
nand U8272 (N_8272,N_7927,N_7821);
nor U8273 (N_8273,N_7888,N_7557);
nor U8274 (N_8274,N_7517,N_7721);
and U8275 (N_8275,N_7999,N_7614);
nand U8276 (N_8276,N_7718,N_7890);
nor U8277 (N_8277,N_7824,N_7707);
or U8278 (N_8278,N_7994,N_7773);
or U8279 (N_8279,N_7838,N_7719);
xor U8280 (N_8280,N_7777,N_7599);
and U8281 (N_8281,N_7711,N_7569);
or U8282 (N_8282,N_7764,N_7991);
nand U8283 (N_8283,N_7978,N_7877);
nor U8284 (N_8284,N_7556,N_7953);
nor U8285 (N_8285,N_7802,N_7940);
or U8286 (N_8286,N_7824,N_7580);
or U8287 (N_8287,N_7783,N_7841);
nand U8288 (N_8288,N_7971,N_7604);
nor U8289 (N_8289,N_7865,N_7986);
xor U8290 (N_8290,N_7774,N_7736);
nor U8291 (N_8291,N_7756,N_7938);
nor U8292 (N_8292,N_7708,N_7692);
or U8293 (N_8293,N_7516,N_7794);
or U8294 (N_8294,N_7654,N_7959);
xor U8295 (N_8295,N_7510,N_7824);
xor U8296 (N_8296,N_7692,N_7646);
and U8297 (N_8297,N_7837,N_7518);
or U8298 (N_8298,N_7622,N_7605);
xor U8299 (N_8299,N_7654,N_7965);
xnor U8300 (N_8300,N_7708,N_7916);
nand U8301 (N_8301,N_7536,N_7915);
xor U8302 (N_8302,N_7583,N_7871);
and U8303 (N_8303,N_7658,N_7834);
and U8304 (N_8304,N_7749,N_7881);
and U8305 (N_8305,N_7905,N_7657);
and U8306 (N_8306,N_7680,N_7948);
nor U8307 (N_8307,N_7853,N_7691);
nor U8308 (N_8308,N_7954,N_7841);
nor U8309 (N_8309,N_7536,N_7659);
xnor U8310 (N_8310,N_7976,N_7894);
or U8311 (N_8311,N_7639,N_7514);
or U8312 (N_8312,N_7965,N_7777);
or U8313 (N_8313,N_7926,N_7505);
nand U8314 (N_8314,N_7773,N_7769);
xnor U8315 (N_8315,N_7946,N_7773);
or U8316 (N_8316,N_7607,N_7692);
or U8317 (N_8317,N_7639,N_7615);
nor U8318 (N_8318,N_7508,N_7611);
xor U8319 (N_8319,N_7864,N_7822);
xnor U8320 (N_8320,N_7697,N_7876);
or U8321 (N_8321,N_7918,N_7880);
or U8322 (N_8322,N_7868,N_7755);
xor U8323 (N_8323,N_7524,N_7641);
nand U8324 (N_8324,N_7982,N_7632);
or U8325 (N_8325,N_7964,N_7678);
xnor U8326 (N_8326,N_7612,N_7682);
or U8327 (N_8327,N_7708,N_7644);
xor U8328 (N_8328,N_7875,N_7808);
or U8329 (N_8329,N_7721,N_7593);
nor U8330 (N_8330,N_7873,N_7945);
and U8331 (N_8331,N_7765,N_7755);
or U8332 (N_8332,N_7762,N_7887);
nand U8333 (N_8333,N_7515,N_7532);
nand U8334 (N_8334,N_7534,N_7993);
xor U8335 (N_8335,N_7575,N_7701);
xnor U8336 (N_8336,N_7750,N_7747);
and U8337 (N_8337,N_7973,N_7976);
nor U8338 (N_8338,N_7629,N_7774);
and U8339 (N_8339,N_7688,N_7760);
or U8340 (N_8340,N_7567,N_7999);
nand U8341 (N_8341,N_7744,N_7807);
nand U8342 (N_8342,N_7990,N_7526);
nand U8343 (N_8343,N_7923,N_7980);
and U8344 (N_8344,N_7572,N_7856);
xor U8345 (N_8345,N_7702,N_7508);
and U8346 (N_8346,N_7768,N_7667);
xnor U8347 (N_8347,N_7825,N_7627);
nand U8348 (N_8348,N_7857,N_7842);
xor U8349 (N_8349,N_7731,N_7677);
and U8350 (N_8350,N_7715,N_7804);
nor U8351 (N_8351,N_7992,N_7837);
nand U8352 (N_8352,N_7902,N_7518);
nand U8353 (N_8353,N_7685,N_7767);
and U8354 (N_8354,N_7877,N_7583);
xor U8355 (N_8355,N_7803,N_7648);
or U8356 (N_8356,N_7990,N_7844);
nand U8357 (N_8357,N_7683,N_7635);
nor U8358 (N_8358,N_7836,N_7889);
or U8359 (N_8359,N_7526,N_7572);
xnor U8360 (N_8360,N_7685,N_7565);
xnor U8361 (N_8361,N_7586,N_7510);
nand U8362 (N_8362,N_7983,N_7548);
xnor U8363 (N_8363,N_7702,N_7843);
nand U8364 (N_8364,N_7643,N_7752);
and U8365 (N_8365,N_7598,N_7832);
nor U8366 (N_8366,N_7515,N_7765);
and U8367 (N_8367,N_7880,N_7738);
or U8368 (N_8368,N_7722,N_7841);
nand U8369 (N_8369,N_7674,N_7678);
or U8370 (N_8370,N_7933,N_7631);
nor U8371 (N_8371,N_7661,N_7511);
nor U8372 (N_8372,N_7837,N_7811);
nor U8373 (N_8373,N_7544,N_7663);
and U8374 (N_8374,N_7765,N_7842);
and U8375 (N_8375,N_7581,N_7771);
nand U8376 (N_8376,N_7765,N_7857);
xor U8377 (N_8377,N_7604,N_7743);
and U8378 (N_8378,N_7621,N_7919);
or U8379 (N_8379,N_7607,N_7941);
or U8380 (N_8380,N_7858,N_7940);
or U8381 (N_8381,N_7521,N_7661);
and U8382 (N_8382,N_7568,N_7504);
xor U8383 (N_8383,N_7985,N_7601);
and U8384 (N_8384,N_7516,N_7820);
or U8385 (N_8385,N_7500,N_7967);
and U8386 (N_8386,N_7535,N_7555);
and U8387 (N_8387,N_7829,N_7699);
and U8388 (N_8388,N_7839,N_7757);
xnor U8389 (N_8389,N_7951,N_7949);
or U8390 (N_8390,N_7518,N_7570);
xor U8391 (N_8391,N_7618,N_7880);
nor U8392 (N_8392,N_7848,N_7812);
nand U8393 (N_8393,N_7808,N_7535);
and U8394 (N_8394,N_7593,N_7507);
nor U8395 (N_8395,N_7699,N_7630);
nand U8396 (N_8396,N_7685,N_7668);
and U8397 (N_8397,N_7922,N_7803);
nor U8398 (N_8398,N_7946,N_7698);
or U8399 (N_8399,N_7821,N_7791);
and U8400 (N_8400,N_7771,N_7556);
nor U8401 (N_8401,N_7965,N_7529);
and U8402 (N_8402,N_7699,N_7597);
nand U8403 (N_8403,N_7679,N_7812);
and U8404 (N_8404,N_7969,N_7633);
nor U8405 (N_8405,N_7604,N_7867);
xnor U8406 (N_8406,N_7687,N_7892);
and U8407 (N_8407,N_7923,N_7952);
xnor U8408 (N_8408,N_7993,N_7846);
xor U8409 (N_8409,N_7545,N_7993);
nand U8410 (N_8410,N_7752,N_7930);
and U8411 (N_8411,N_7564,N_7743);
and U8412 (N_8412,N_7903,N_7598);
nor U8413 (N_8413,N_7684,N_7640);
nor U8414 (N_8414,N_7882,N_7738);
xnor U8415 (N_8415,N_7915,N_7895);
or U8416 (N_8416,N_7807,N_7621);
nand U8417 (N_8417,N_7611,N_7504);
nor U8418 (N_8418,N_7859,N_7564);
nand U8419 (N_8419,N_7701,N_7671);
nor U8420 (N_8420,N_7880,N_7957);
nor U8421 (N_8421,N_7825,N_7889);
nand U8422 (N_8422,N_7834,N_7629);
nand U8423 (N_8423,N_7784,N_7839);
or U8424 (N_8424,N_7793,N_7649);
xor U8425 (N_8425,N_7866,N_7650);
nand U8426 (N_8426,N_7704,N_7999);
and U8427 (N_8427,N_7991,N_7715);
nor U8428 (N_8428,N_7583,N_7705);
and U8429 (N_8429,N_7525,N_7929);
or U8430 (N_8430,N_7869,N_7725);
and U8431 (N_8431,N_7819,N_7941);
and U8432 (N_8432,N_7732,N_7946);
or U8433 (N_8433,N_7793,N_7733);
or U8434 (N_8434,N_7708,N_7929);
nor U8435 (N_8435,N_7513,N_7507);
and U8436 (N_8436,N_7793,N_7611);
or U8437 (N_8437,N_7681,N_7895);
nand U8438 (N_8438,N_7735,N_7583);
or U8439 (N_8439,N_7857,N_7990);
and U8440 (N_8440,N_7726,N_7979);
nand U8441 (N_8441,N_7833,N_7852);
nor U8442 (N_8442,N_7622,N_7927);
xor U8443 (N_8443,N_7962,N_7712);
or U8444 (N_8444,N_7545,N_7692);
nor U8445 (N_8445,N_7701,N_7509);
nand U8446 (N_8446,N_7969,N_7626);
nand U8447 (N_8447,N_7901,N_7641);
nand U8448 (N_8448,N_7735,N_7612);
and U8449 (N_8449,N_7808,N_7736);
nor U8450 (N_8450,N_7644,N_7863);
and U8451 (N_8451,N_7658,N_7692);
or U8452 (N_8452,N_7713,N_7632);
and U8453 (N_8453,N_7833,N_7985);
and U8454 (N_8454,N_7945,N_7852);
nand U8455 (N_8455,N_7693,N_7880);
or U8456 (N_8456,N_7681,N_7825);
and U8457 (N_8457,N_7988,N_7912);
or U8458 (N_8458,N_7746,N_7794);
nor U8459 (N_8459,N_7938,N_7632);
nand U8460 (N_8460,N_7715,N_7899);
nand U8461 (N_8461,N_7596,N_7854);
and U8462 (N_8462,N_7548,N_7788);
xnor U8463 (N_8463,N_7749,N_7833);
and U8464 (N_8464,N_7709,N_7922);
nand U8465 (N_8465,N_7672,N_7929);
or U8466 (N_8466,N_7766,N_7819);
and U8467 (N_8467,N_7856,N_7920);
and U8468 (N_8468,N_7898,N_7984);
xnor U8469 (N_8469,N_7704,N_7557);
xnor U8470 (N_8470,N_7647,N_7813);
or U8471 (N_8471,N_7660,N_7591);
or U8472 (N_8472,N_7873,N_7809);
nand U8473 (N_8473,N_7603,N_7912);
xnor U8474 (N_8474,N_7764,N_7750);
nor U8475 (N_8475,N_7841,N_7565);
or U8476 (N_8476,N_7906,N_7854);
and U8477 (N_8477,N_7644,N_7932);
or U8478 (N_8478,N_7509,N_7730);
or U8479 (N_8479,N_7879,N_7670);
nand U8480 (N_8480,N_7758,N_7936);
or U8481 (N_8481,N_7765,N_7875);
and U8482 (N_8482,N_7585,N_7870);
nor U8483 (N_8483,N_7972,N_7840);
and U8484 (N_8484,N_7924,N_7518);
nor U8485 (N_8485,N_7538,N_7733);
nand U8486 (N_8486,N_7645,N_7704);
and U8487 (N_8487,N_7645,N_7817);
and U8488 (N_8488,N_7661,N_7886);
nor U8489 (N_8489,N_7847,N_7595);
and U8490 (N_8490,N_7847,N_7982);
and U8491 (N_8491,N_7925,N_7815);
nor U8492 (N_8492,N_7735,N_7932);
xnor U8493 (N_8493,N_7746,N_7789);
nand U8494 (N_8494,N_7541,N_7887);
nor U8495 (N_8495,N_7912,N_7744);
nand U8496 (N_8496,N_7539,N_7782);
nand U8497 (N_8497,N_7579,N_7787);
xnor U8498 (N_8498,N_7863,N_7544);
xor U8499 (N_8499,N_7576,N_7952);
nor U8500 (N_8500,N_8212,N_8163);
and U8501 (N_8501,N_8433,N_8323);
nand U8502 (N_8502,N_8167,N_8075);
or U8503 (N_8503,N_8076,N_8297);
and U8504 (N_8504,N_8352,N_8121);
nor U8505 (N_8505,N_8048,N_8201);
nand U8506 (N_8506,N_8446,N_8105);
and U8507 (N_8507,N_8015,N_8128);
xor U8508 (N_8508,N_8218,N_8152);
and U8509 (N_8509,N_8235,N_8178);
nand U8510 (N_8510,N_8276,N_8210);
or U8511 (N_8511,N_8261,N_8228);
nor U8512 (N_8512,N_8329,N_8248);
nor U8513 (N_8513,N_8388,N_8209);
and U8514 (N_8514,N_8456,N_8394);
nor U8515 (N_8515,N_8362,N_8103);
xor U8516 (N_8516,N_8114,N_8101);
xnor U8517 (N_8517,N_8309,N_8030);
nor U8518 (N_8518,N_8018,N_8308);
xor U8519 (N_8519,N_8135,N_8390);
or U8520 (N_8520,N_8196,N_8255);
nand U8521 (N_8521,N_8017,N_8193);
and U8522 (N_8522,N_8392,N_8156);
and U8523 (N_8523,N_8066,N_8479);
nor U8524 (N_8524,N_8141,N_8002);
nor U8525 (N_8525,N_8377,N_8422);
xnor U8526 (N_8526,N_8151,N_8040);
or U8527 (N_8527,N_8189,N_8344);
nand U8528 (N_8528,N_8369,N_8359);
nand U8529 (N_8529,N_8117,N_8122);
and U8530 (N_8530,N_8085,N_8125);
nor U8531 (N_8531,N_8454,N_8476);
nor U8532 (N_8532,N_8160,N_8461);
or U8533 (N_8533,N_8036,N_8184);
nand U8534 (N_8534,N_8053,N_8473);
xor U8535 (N_8535,N_8245,N_8445);
nor U8536 (N_8536,N_8098,N_8090);
xnor U8537 (N_8537,N_8407,N_8269);
nor U8538 (N_8538,N_8343,N_8314);
xor U8539 (N_8539,N_8136,N_8350);
nand U8540 (N_8540,N_8417,N_8197);
or U8541 (N_8541,N_8188,N_8093);
nor U8542 (N_8542,N_8464,N_8325);
nand U8543 (N_8543,N_8347,N_8161);
nor U8544 (N_8544,N_8251,N_8234);
nor U8545 (N_8545,N_8299,N_8266);
xor U8546 (N_8546,N_8026,N_8318);
nor U8547 (N_8547,N_8247,N_8285);
or U8548 (N_8548,N_8070,N_8452);
or U8549 (N_8549,N_8181,N_8169);
xnor U8550 (N_8550,N_8466,N_8246);
nand U8551 (N_8551,N_8172,N_8435);
xor U8552 (N_8552,N_8219,N_8086);
and U8553 (N_8553,N_8284,N_8013);
and U8554 (N_8554,N_8168,N_8371);
nand U8555 (N_8555,N_8304,N_8496);
and U8556 (N_8556,N_8395,N_8425);
nand U8557 (N_8557,N_8370,N_8175);
nand U8558 (N_8558,N_8490,N_8354);
xnor U8559 (N_8559,N_8375,N_8112);
nand U8560 (N_8560,N_8233,N_8293);
or U8561 (N_8561,N_8379,N_8278);
nand U8562 (N_8562,N_8489,N_8328);
nand U8563 (N_8563,N_8191,N_8068);
xor U8564 (N_8564,N_8259,N_8029);
and U8565 (N_8565,N_8413,N_8404);
nor U8566 (N_8566,N_8094,N_8494);
or U8567 (N_8567,N_8250,N_8355);
nand U8568 (N_8568,N_8262,N_8241);
or U8569 (N_8569,N_8291,N_8001);
or U8570 (N_8570,N_8092,N_8202);
or U8571 (N_8571,N_8294,N_8238);
and U8572 (N_8572,N_8111,N_8436);
xor U8573 (N_8573,N_8140,N_8367);
or U8574 (N_8574,N_8383,N_8399);
nor U8575 (N_8575,N_8072,N_8418);
nor U8576 (N_8576,N_8408,N_8281);
and U8577 (N_8577,N_8062,N_8217);
and U8578 (N_8578,N_8470,N_8353);
and U8579 (N_8579,N_8173,N_8035);
xor U8580 (N_8580,N_8410,N_8481);
and U8581 (N_8581,N_8467,N_8236);
and U8582 (N_8582,N_8463,N_8084);
nor U8583 (N_8583,N_8215,N_8083);
and U8584 (N_8584,N_8447,N_8416);
and U8585 (N_8585,N_8147,N_8453);
nand U8586 (N_8586,N_8270,N_8120);
nor U8587 (N_8587,N_8483,N_8038);
and U8588 (N_8588,N_8044,N_8216);
nor U8589 (N_8589,N_8381,N_8356);
xor U8590 (N_8590,N_8346,N_8198);
nor U8591 (N_8591,N_8257,N_8031);
xor U8592 (N_8592,N_8214,N_8097);
nor U8593 (N_8593,N_8378,N_8115);
xnor U8594 (N_8594,N_8091,N_8339);
or U8595 (N_8595,N_8155,N_8012);
nor U8596 (N_8596,N_8372,N_8438);
xor U8597 (N_8597,N_8049,N_8337);
xor U8598 (N_8598,N_8348,N_8039);
nor U8599 (N_8599,N_8154,N_8272);
nor U8600 (N_8600,N_8492,N_8170);
nor U8601 (N_8601,N_8174,N_8267);
and U8602 (N_8602,N_8037,N_8386);
and U8603 (N_8603,N_8148,N_8171);
or U8604 (N_8604,N_8340,N_8341);
nor U8605 (N_8605,N_8254,N_8132);
nand U8606 (N_8606,N_8028,N_8055);
nand U8607 (N_8607,N_8471,N_8050);
or U8608 (N_8608,N_8474,N_8222);
xnor U8609 (N_8609,N_8402,N_8279);
and U8610 (N_8610,N_8162,N_8065);
xnor U8611 (N_8611,N_8130,N_8145);
or U8612 (N_8612,N_8441,N_8143);
nor U8613 (N_8613,N_8211,N_8127);
nor U8614 (N_8614,N_8139,N_8207);
or U8615 (N_8615,N_8421,N_8482);
nand U8616 (N_8616,N_8368,N_8208);
or U8617 (N_8617,N_8223,N_8336);
or U8618 (N_8618,N_8240,N_8296);
nor U8619 (N_8619,N_8468,N_8342);
and U8620 (N_8620,N_8321,N_8187);
xnor U8621 (N_8621,N_8007,N_8412);
xor U8622 (N_8622,N_8449,N_8498);
xor U8623 (N_8623,N_8003,N_8016);
xnor U8624 (N_8624,N_8290,N_8439);
nand U8625 (N_8625,N_8190,N_8424);
nand U8626 (N_8626,N_8491,N_8195);
or U8627 (N_8627,N_8054,N_8306);
nand U8628 (N_8628,N_8486,N_8063);
or U8629 (N_8629,N_8025,N_8082);
or U8630 (N_8630,N_8409,N_8067);
xor U8631 (N_8631,N_8319,N_8095);
and U8632 (N_8632,N_8009,N_8434);
nand U8633 (N_8633,N_8312,N_8074);
nor U8634 (N_8634,N_8249,N_8256);
nand U8635 (N_8635,N_8224,N_8387);
xnor U8636 (N_8636,N_8330,N_8406);
xor U8637 (N_8637,N_8391,N_8226);
nand U8638 (N_8638,N_8389,N_8046);
nor U8639 (N_8639,N_8363,N_8485);
xor U8640 (N_8640,N_8042,N_8420);
or U8641 (N_8641,N_8366,N_8004);
or U8642 (N_8642,N_8164,N_8428);
nand U8643 (N_8643,N_8260,N_8183);
and U8644 (N_8644,N_8385,N_8034);
nor U8645 (N_8645,N_8397,N_8374);
and U8646 (N_8646,N_8146,N_8008);
nand U8647 (N_8647,N_8089,N_8326);
and U8648 (N_8648,N_8430,N_8429);
xnor U8649 (N_8649,N_8024,N_8131);
or U8650 (N_8650,N_8165,N_8292);
nand U8651 (N_8651,N_8477,N_8316);
and U8652 (N_8652,N_8149,N_8398);
nand U8653 (N_8653,N_8403,N_8448);
or U8654 (N_8654,N_8286,N_8073);
xor U8655 (N_8655,N_8118,N_8088);
and U8656 (N_8656,N_8061,N_8019);
nor U8657 (N_8657,N_8023,N_8064);
xor U8658 (N_8658,N_8185,N_8079);
and U8659 (N_8659,N_8100,N_8032);
and U8660 (N_8660,N_8011,N_8153);
xnor U8661 (N_8661,N_8194,N_8123);
xor U8662 (N_8662,N_8493,N_8200);
and U8663 (N_8663,N_8205,N_8186);
xor U8664 (N_8664,N_8396,N_8334);
nand U8665 (N_8665,N_8440,N_8229);
or U8666 (N_8666,N_8313,N_8014);
or U8667 (N_8667,N_8225,N_8349);
nand U8668 (N_8668,N_8415,N_8443);
xnor U8669 (N_8669,N_8499,N_8041);
or U8670 (N_8670,N_8010,N_8232);
or U8671 (N_8671,N_8315,N_8231);
or U8672 (N_8672,N_8119,N_8124);
nand U8673 (N_8673,N_8472,N_8258);
nor U8674 (N_8674,N_8206,N_8033);
nand U8675 (N_8675,N_8203,N_8364);
nor U8676 (N_8676,N_8005,N_8332);
or U8677 (N_8677,N_8265,N_8077);
or U8678 (N_8678,N_8327,N_8204);
xnor U8679 (N_8679,N_8283,N_8144);
xnor U8680 (N_8680,N_8058,N_8027);
and U8681 (N_8681,N_8380,N_8134);
and U8682 (N_8682,N_8102,N_8271);
and U8683 (N_8683,N_8087,N_8045);
and U8684 (N_8684,N_8431,N_8335);
nand U8685 (N_8685,N_8444,N_8126);
nand U8686 (N_8686,N_8317,N_8192);
xnor U8687 (N_8687,N_8426,N_8282);
nand U8688 (N_8688,N_8052,N_8080);
nor U8689 (N_8689,N_8239,N_8405);
and U8690 (N_8690,N_8376,N_8137);
nor U8691 (N_8691,N_8459,N_8047);
or U8692 (N_8692,N_8277,N_8081);
nor U8693 (N_8693,N_8333,N_8107);
xor U8694 (N_8694,N_8138,N_8274);
xor U8695 (N_8695,N_8360,N_8020);
xor U8696 (N_8696,N_8303,N_8060);
xor U8697 (N_8697,N_8157,N_8495);
xnor U8698 (N_8698,N_8462,N_8237);
xor U8699 (N_8699,N_8227,N_8331);
or U8700 (N_8700,N_8320,N_8484);
nor U8701 (N_8701,N_8393,N_8338);
xnor U8702 (N_8702,N_8006,N_8051);
or U8703 (N_8703,N_8150,N_8469);
nor U8704 (N_8704,N_8022,N_8253);
nor U8705 (N_8705,N_8263,N_8182);
and U8706 (N_8706,N_8113,N_8307);
nand U8707 (N_8707,N_8458,N_8280);
xor U8708 (N_8708,N_8311,N_8180);
nor U8709 (N_8709,N_8043,N_8460);
and U8710 (N_8710,N_8159,N_8450);
and U8711 (N_8711,N_8289,N_8384);
or U8712 (N_8712,N_8302,N_8478);
and U8713 (N_8713,N_8457,N_8455);
nand U8714 (N_8714,N_8106,N_8268);
nor U8715 (N_8715,N_8305,N_8345);
nor U8716 (N_8716,N_8497,N_8221);
and U8717 (N_8717,N_8158,N_8351);
nor U8718 (N_8718,N_8488,N_8252);
nor U8719 (N_8719,N_8373,N_8109);
or U8720 (N_8720,N_8465,N_8166);
nand U8721 (N_8721,N_8365,N_8301);
xor U8722 (N_8722,N_8324,N_8116);
nor U8723 (N_8723,N_8475,N_8056);
or U8724 (N_8724,N_8419,N_8487);
nor U8725 (N_8725,N_8295,N_8361);
and U8726 (N_8726,N_8300,N_8199);
nand U8727 (N_8727,N_8059,N_8310);
nand U8728 (N_8728,N_8275,N_8401);
and U8729 (N_8729,N_8133,N_8110);
or U8730 (N_8730,N_8382,N_8273);
xor U8731 (N_8731,N_8078,N_8142);
and U8732 (N_8732,N_8176,N_8298);
and U8733 (N_8733,N_8179,N_8230);
and U8734 (N_8734,N_8432,N_8213);
nand U8735 (N_8735,N_8451,N_8000);
xor U8736 (N_8736,N_8414,N_8071);
xor U8737 (N_8737,N_8288,N_8322);
nor U8738 (N_8738,N_8021,N_8242);
or U8739 (N_8739,N_8244,N_8264);
nor U8740 (N_8740,N_8357,N_8243);
nand U8741 (N_8741,N_8427,N_8129);
or U8742 (N_8742,N_8442,N_8480);
and U8743 (N_8743,N_8057,N_8358);
nor U8744 (N_8744,N_8220,N_8104);
and U8745 (N_8745,N_8287,N_8437);
xnor U8746 (N_8746,N_8069,N_8096);
xor U8747 (N_8747,N_8108,N_8411);
nand U8748 (N_8748,N_8177,N_8423);
and U8749 (N_8749,N_8400,N_8099);
nand U8750 (N_8750,N_8302,N_8110);
or U8751 (N_8751,N_8364,N_8117);
nor U8752 (N_8752,N_8319,N_8433);
nand U8753 (N_8753,N_8289,N_8443);
and U8754 (N_8754,N_8147,N_8362);
nand U8755 (N_8755,N_8486,N_8286);
nor U8756 (N_8756,N_8170,N_8400);
xor U8757 (N_8757,N_8080,N_8299);
xnor U8758 (N_8758,N_8148,N_8313);
nand U8759 (N_8759,N_8266,N_8149);
or U8760 (N_8760,N_8263,N_8095);
xor U8761 (N_8761,N_8346,N_8039);
and U8762 (N_8762,N_8304,N_8228);
nor U8763 (N_8763,N_8330,N_8343);
and U8764 (N_8764,N_8026,N_8382);
or U8765 (N_8765,N_8158,N_8432);
and U8766 (N_8766,N_8171,N_8319);
and U8767 (N_8767,N_8350,N_8131);
nand U8768 (N_8768,N_8362,N_8046);
or U8769 (N_8769,N_8290,N_8386);
xnor U8770 (N_8770,N_8204,N_8114);
xor U8771 (N_8771,N_8484,N_8091);
nand U8772 (N_8772,N_8408,N_8378);
nand U8773 (N_8773,N_8208,N_8489);
and U8774 (N_8774,N_8393,N_8474);
and U8775 (N_8775,N_8357,N_8328);
and U8776 (N_8776,N_8189,N_8435);
nand U8777 (N_8777,N_8206,N_8013);
xnor U8778 (N_8778,N_8282,N_8460);
nand U8779 (N_8779,N_8211,N_8367);
and U8780 (N_8780,N_8070,N_8223);
nor U8781 (N_8781,N_8146,N_8245);
or U8782 (N_8782,N_8216,N_8090);
and U8783 (N_8783,N_8069,N_8103);
nand U8784 (N_8784,N_8130,N_8278);
nand U8785 (N_8785,N_8020,N_8437);
nand U8786 (N_8786,N_8311,N_8107);
or U8787 (N_8787,N_8184,N_8240);
and U8788 (N_8788,N_8079,N_8190);
and U8789 (N_8789,N_8115,N_8033);
and U8790 (N_8790,N_8385,N_8138);
nor U8791 (N_8791,N_8446,N_8428);
nand U8792 (N_8792,N_8497,N_8357);
nor U8793 (N_8793,N_8286,N_8299);
xor U8794 (N_8794,N_8136,N_8381);
or U8795 (N_8795,N_8164,N_8291);
nand U8796 (N_8796,N_8336,N_8019);
nor U8797 (N_8797,N_8327,N_8267);
nand U8798 (N_8798,N_8190,N_8421);
nand U8799 (N_8799,N_8181,N_8218);
xnor U8800 (N_8800,N_8378,N_8210);
nand U8801 (N_8801,N_8223,N_8250);
or U8802 (N_8802,N_8489,N_8102);
nor U8803 (N_8803,N_8299,N_8085);
and U8804 (N_8804,N_8099,N_8496);
nor U8805 (N_8805,N_8051,N_8304);
and U8806 (N_8806,N_8433,N_8082);
and U8807 (N_8807,N_8446,N_8168);
xnor U8808 (N_8808,N_8121,N_8278);
xnor U8809 (N_8809,N_8228,N_8193);
and U8810 (N_8810,N_8416,N_8070);
xor U8811 (N_8811,N_8125,N_8229);
and U8812 (N_8812,N_8021,N_8280);
and U8813 (N_8813,N_8051,N_8495);
or U8814 (N_8814,N_8194,N_8034);
xnor U8815 (N_8815,N_8105,N_8028);
nand U8816 (N_8816,N_8223,N_8387);
nor U8817 (N_8817,N_8223,N_8166);
and U8818 (N_8818,N_8008,N_8272);
nand U8819 (N_8819,N_8357,N_8414);
xnor U8820 (N_8820,N_8383,N_8056);
and U8821 (N_8821,N_8201,N_8361);
and U8822 (N_8822,N_8111,N_8161);
nand U8823 (N_8823,N_8460,N_8226);
and U8824 (N_8824,N_8138,N_8137);
or U8825 (N_8825,N_8112,N_8342);
xnor U8826 (N_8826,N_8147,N_8068);
and U8827 (N_8827,N_8152,N_8348);
or U8828 (N_8828,N_8480,N_8059);
nor U8829 (N_8829,N_8446,N_8229);
nand U8830 (N_8830,N_8227,N_8311);
xor U8831 (N_8831,N_8258,N_8316);
or U8832 (N_8832,N_8372,N_8385);
nor U8833 (N_8833,N_8075,N_8124);
and U8834 (N_8834,N_8133,N_8489);
nor U8835 (N_8835,N_8025,N_8453);
or U8836 (N_8836,N_8404,N_8172);
nor U8837 (N_8837,N_8305,N_8323);
and U8838 (N_8838,N_8417,N_8178);
nand U8839 (N_8839,N_8379,N_8243);
xnor U8840 (N_8840,N_8023,N_8291);
or U8841 (N_8841,N_8336,N_8390);
nand U8842 (N_8842,N_8247,N_8318);
nand U8843 (N_8843,N_8125,N_8249);
nand U8844 (N_8844,N_8049,N_8283);
nor U8845 (N_8845,N_8326,N_8016);
nand U8846 (N_8846,N_8192,N_8032);
xor U8847 (N_8847,N_8275,N_8496);
nand U8848 (N_8848,N_8149,N_8380);
and U8849 (N_8849,N_8498,N_8166);
xor U8850 (N_8850,N_8353,N_8173);
nand U8851 (N_8851,N_8195,N_8041);
or U8852 (N_8852,N_8197,N_8360);
nor U8853 (N_8853,N_8258,N_8168);
or U8854 (N_8854,N_8373,N_8497);
nor U8855 (N_8855,N_8148,N_8298);
and U8856 (N_8856,N_8424,N_8412);
xor U8857 (N_8857,N_8217,N_8201);
and U8858 (N_8858,N_8053,N_8166);
and U8859 (N_8859,N_8038,N_8118);
xnor U8860 (N_8860,N_8305,N_8382);
and U8861 (N_8861,N_8165,N_8384);
nand U8862 (N_8862,N_8032,N_8370);
nand U8863 (N_8863,N_8452,N_8016);
nor U8864 (N_8864,N_8019,N_8354);
and U8865 (N_8865,N_8484,N_8380);
or U8866 (N_8866,N_8300,N_8287);
nor U8867 (N_8867,N_8439,N_8057);
nor U8868 (N_8868,N_8126,N_8058);
and U8869 (N_8869,N_8000,N_8079);
nor U8870 (N_8870,N_8449,N_8171);
nor U8871 (N_8871,N_8138,N_8223);
or U8872 (N_8872,N_8032,N_8203);
nor U8873 (N_8873,N_8195,N_8135);
nand U8874 (N_8874,N_8224,N_8345);
or U8875 (N_8875,N_8221,N_8430);
nor U8876 (N_8876,N_8396,N_8464);
and U8877 (N_8877,N_8492,N_8015);
xnor U8878 (N_8878,N_8221,N_8350);
nor U8879 (N_8879,N_8198,N_8350);
and U8880 (N_8880,N_8138,N_8454);
nand U8881 (N_8881,N_8163,N_8162);
or U8882 (N_8882,N_8035,N_8021);
or U8883 (N_8883,N_8498,N_8248);
xnor U8884 (N_8884,N_8069,N_8368);
and U8885 (N_8885,N_8296,N_8291);
and U8886 (N_8886,N_8270,N_8283);
nand U8887 (N_8887,N_8091,N_8202);
or U8888 (N_8888,N_8332,N_8154);
and U8889 (N_8889,N_8380,N_8066);
nor U8890 (N_8890,N_8017,N_8327);
nand U8891 (N_8891,N_8062,N_8191);
or U8892 (N_8892,N_8054,N_8177);
and U8893 (N_8893,N_8285,N_8151);
or U8894 (N_8894,N_8333,N_8114);
nor U8895 (N_8895,N_8472,N_8295);
nor U8896 (N_8896,N_8014,N_8242);
nor U8897 (N_8897,N_8082,N_8171);
nand U8898 (N_8898,N_8459,N_8442);
nor U8899 (N_8899,N_8230,N_8327);
nor U8900 (N_8900,N_8436,N_8379);
and U8901 (N_8901,N_8100,N_8392);
or U8902 (N_8902,N_8169,N_8010);
or U8903 (N_8903,N_8242,N_8336);
xnor U8904 (N_8904,N_8227,N_8078);
xor U8905 (N_8905,N_8346,N_8008);
nand U8906 (N_8906,N_8144,N_8281);
or U8907 (N_8907,N_8309,N_8020);
xor U8908 (N_8908,N_8301,N_8038);
nand U8909 (N_8909,N_8400,N_8455);
and U8910 (N_8910,N_8462,N_8253);
and U8911 (N_8911,N_8487,N_8066);
xnor U8912 (N_8912,N_8456,N_8123);
or U8913 (N_8913,N_8490,N_8139);
nor U8914 (N_8914,N_8286,N_8245);
or U8915 (N_8915,N_8359,N_8059);
and U8916 (N_8916,N_8398,N_8221);
nand U8917 (N_8917,N_8442,N_8117);
or U8918 (N_8918,N_8424,N_8484);
nand U8919 (N_8919,N_8280,N_8302);
or U8920 (N_8920,N_8472,N_8437);
nor U8921 (N_8921,N_8359,N_8435);
xor U8922 (N_8922,N_8026,N_8022);
or U8923 (N_8923,N_8226,N_8484);
nand U8924 (N_8924,N_8216,N_8287);
xnor U8925 (N_8925,N_8367,N_8123);
nand U8926 (N_8926,N_8034,N_8420);
and U8927 (N_8927,N_8033,N_8132);
or U8928 (N_8928,N_8356,N_8385);
or U8929 (N_8929,N_8294,N_8020);
nor U8930 (N_8930,N_8177,N_8325);
and U8931 (N_8931,N_8162,N_8087);
and U8932 (N_8932,N_8382,N_8021);
nand U8933 (N_8933,N_8015,N_8314);
and U8934 (N_8934,N_8110,N_8006);
nor U8935 (N_8935,N_8491,N_8221);
and U8936 (N_8936,N_8076,N_8483);
nor U8937 (N_8937,N_8211,N_8488);
and U8938 (N_8938,N_8409,N_8390);
or U8939 (N_8939,N_8238,N_8061);
nand U8940 (N_8940,N_8116,N_8492);
and U8941 (N_8941,N_8066,N_8357);
nor U8942 (N_8942,N_8283,N_8323);
xnor U8943 (N_8943,N_8456,N_8056);
and U8944 (N_8944,N_8167,N_8355);
xnor U8945 (N_8945,N_8041,N_8464);
nand U8946 (N_8946,N_8473,N_8469);
or U8947 (N_8947,N_8277,N_8482);
and U8948 (N_8948,N_8172,N_8324);
nand U8949 (N_8949,N_8342,N_8196);
and U8950 (N_8950,N_8319,N_8265);
and U8951 (N_8951,N_8085,N_8383);
nor U8952 (N_8952,N_8014,N_8090);
nand U8953 (N_8953,N_8337,N_8109);
or U8954 (N_8954,N_8178,N_8281);
nand U8955 (N_8955,N_8489,N_8303);
nor U8956 (N_8956,N_8260,N_8044);
or U8957 (N_8957,N_8097,N_8034);
and U8958 (N_8958,N_8359,N_8283);
nor U8959 (N_8959,N_8194,N_8100);
nor U8960 (N_8960,N_8363,N_8251);
nand U8961 (N_8961,N_8244,N_8062);
nand U8962 (N_8962,N_8139,N_8331);
nor U8963 (N_8963,N_8428,N_8314);
and U8964 (N_8964,N_8352,N_8033);
or U8965 (N_8965,N_8400,N_8091);
and U8966 (N_8966,N_8244,N_8453);
or U8967 (N_8967,N_8412,N_8363);
nor U8968 (N_8968,N_8143,N_8386);
xnor U8969 (N_8969,N_8430,N_8305);
nor U8970 (N_8970,N_8493,N_8431);
xor U8971 (N_8971,N_8310,N_8222);
or U8972 (N_8972,N_8331,N_8475);
nor U8973 (N_8973,N_8335,N_8456);
nand U8974 (N_8974,N_8204,N_8124);
or U8975 (N_8975,N_8479,N_8296);
nor U8976 (N_8976,N_8412,N_8302);
nor U8977 (N_8977,N_8435,N_8461);
nand U8978 (N_8978,N_8090,N_8114);
or U8979 (N_8979,N_8255,N_8075);
xor U8980 (N_8980,N_8163,N_8211);
xnor U8981 (N_8981,N_8304,N_8300);
xor U8982 (N_8982,N_8327,N_8297);
nand U8983 (N_8983,N_8459,N_8044);
xor U8984 (N_8984,N_8363,N_8348);
xnor U8985 (N_8985,N_8017,N_8339);
nor U8986 (N_8986,N_8117,N_8428);
nor U8987 (N_8987,N_8304,N_8081);
nand U8988 (N_8988,N_8491,N_8159);
nor U8989 (N_8989,N_8268,N_8447);
nand U8990 (N_8990,N_8459,N_8251);
nand U8991 (N_8991,N_8037,N_8488);
or U8992 (N_8992,N_8477,N_8419);
or U8993 (N_8993,N_8095,N_8253);
nor U8994 (N_8994,N_8218,N_8185);
or U8995 (N_8995,N_8228,N_8022);
nor U8996 (N_8996,N_8234,N_8330);
or U8997 (N_8997,N_8150,N_8334);
or U8998 (N_8998,N_8155,N_8328);
xor U8999 (N_8999,N_8418,N_8121);
and U9000 (N_9000,N_8720,N_8793);
xor U9001 (N_9001,N_8846,N_8840);
xor U9002 (N_9002,N_8818,N_8817);
xor U9003 (N_9003,N_8651,N_8614);
xor U9004 (N_9004,N_8766,N_8969);
nand U9005 (N_9005,N_8533,N_8826);
and U9006 (N_9006,N_8900,N_8882);
and U9007 (N_9007,N_8868,N_8777);
and U9008 (N_9008,N_8652,N_8997);
nand U9009 (N_9009,N_8831,N_8770);
nand U9010 (N_9010,N_8843,N_8716);
or U9011 (N_9011,N_8906,N_8861);
nor U9012 (N_9012,N_8802,N_8837);
and U9013 (N_9013,N_8681,N_8984);
nand U9014 (N_9014,N_8623,N_8819);
and U9015 (N_9015,N_8690,N_8703);
nor U9016 (N_9016,N_8692,N_8705);
xor U9017 (N_9017,N_8803,N_8847);
and U9018 (N_9018,N_8822,N_8604);
nand U9019 (N_9019,N_8530,N_8591);
xnor U9020 (N_9020,N_8838,N_8568);
nor U9021 (N_9021,N_8794,N_8764);
nor U9022 (N_9022,N_8848,N_8684);
or U9023 (N_9023,N_8852,N_8780);
nand U9024 (N_9024,N_8582,N_8827);
and U9025 (N_9025,N_8999,N_8731);
nor U9026 (N_9026,N_8778,N_8760);
or U9027 (N_9027,N_8953,N_8636);
nand U9028 (N_9028,N_8736,N_8632);
and U9029 (N_9029,N_8695,N_8665);
nand U9030 (N_9030,N_8961,N_8552);
or U9031 (N_9031,N_8911,N_8729);
nand U9032 (N_9032,N_8896,N_8554);
nand U9033 (N_9033,N_8518,N_8643);
or U9034 (N_9034,N_8639,N_8740);
and U9035 (N_9035,N_8611,N_8721);
or U9036 (N_9036,N_8795,N_8768);
and U9037 (N_9037,N_8937,N_8546);
or U9038 (N_9038,N_8796,N_8556);
or U9039 (N_9039,N_8743,N_8815);
nand U9040 (N_9040,N_8842,N_8980);
xor U9041 (N_9041,N_8919,N_8517);
nand U9042 (N_9042,N_8691,N_8875);
nor U9043 (N_9043,N_8514,N_8516);
xnor U9044 (N_9044,N_8598,N_8547);
xnor U9045 (N_9045,N_8674,N_8976);
xor U9046 (N_9046,N_8507,N_8996);
nor U9047 (N_9047,N_8672,N_8987);
or U9048 (N_9048,N_8531,N_8801);
nor U9049 (N_9049,N_8913,N_8542);
nor U9050 (N_9050,N_8702,N_8677);
nor U9051 (N_9051,N_8759,N_8745);
xnor U9052 (N_9052,N_8733,N_8522);
or U9053 (N_9053,N_8773,N_8519);
xor U9054 (N_9054,N_8631,N_8946);
and U9055 (N_9055,N_8800,N_8851);
xor U9056 (N_9056,N_8626,N_8947);
xnor U9057 (N_9057,N_8503,N_8700);
nor U9058 (N_9058,N_8908,N_8888);
nor U9059 (N_9059,N_8874,N_8613);
and U9060 (N_9060,N_8675,N_8592);
or U9061 (N_9061,N_8862,N_8914);
and U9062 (N_9062,N_8741,N_8871);
and U9063 (N_9063,N_8685,N_8956);
nand U9064 (N_9064,N_8932,N_8960);
and U9065 (N_9065,N_8616,N_8910);
nor U9066 (N_9066,N_8983,N_8754);
or U9067 (N_9067,N_8739,N_8749);
and U9068 (N_9068,N_8918,N_8804);
and U9069 (N_9069,N_8710,N_8949);
and U9070 (N_9070,N_8979,N_8995);
nand U9071 (N_9071,N_8828,N_8967);
xor U9072 (N_9072,N_8808,N_8501);
and U9073 (N_9073,N_8574,N_8844);
or U9074 (N_9074,N_8915,N_8916);
nand U9075 (N_9075,N_8952,N_8939);
nand U9076 (N_9076,N_8634,N_8669);
xor U9077 (N_9077,N_8718,N_8571);
or U9078 (N_9078,N_8903,N_8789);
nand U9079 (N_9079,N_8673,N_8549);
xor U9080 (N_9080,N_8601,N_8894);
nor U9081 (N_9081,N_8873,N_8543);
xnor U9082 (N_9082,N_8859,N_8593);
or U9083 (N_9083,N_8708,N_8978);
and U9084 (N_9084,N_8779,N_8945);
and U9085 (N_9085,N_8781,N_8699);
and U9086 (N_9086,N_8661,N_8704);
nor U9087 (N_9087,N_8791,N_8620);
nor U9088 (N_9088,N_8858,N_8644);
or U9089 (N_9089,N_8816,N_8940);
and U9090 (N_9090,N_8562,N_8798);
nand U9091 (N_9091,N_8753,N_8608);
nor U9092 (N_9092,N_8662,N_8988);
nand U9093 (N_9093,N_8925,N_8658);
or U9094 (N_9094,N_8974,N_8893);
nor U9095 (N_9095,N_8876,N_8971);
nor U9096 (N_9096,N_8839,N_8878);
or U9097 (N_9097,N_8992,N_8510);
nand U9098 (N_9098,N_8646,N_8879);
nor U9099 (N_9099,N_8648,N_8590);
nor U9100 (N_9100,N_8688,N_8505);
xnor U9101 (N_9101,N_8551,N_8719);
nand U9102 (N_9102,N_8973,N_8724);
nor U9103 (N_9103,N_8727,N_8762);
xnor U9104 (N_9104,N_8653,N_8850);
or U9105 (N_9105,N_8742,N_8752);
and U9106 (N_9106,N_8560,N_8923);
and U9107 (N_9107,N_8845,N_8757);
nand U9108 (N_9108,N_8867,N_8748);
and U9109 (N_9109,N_8557,N_8735);
or U9110 (N_9110,N_8640,N_8587);
xnor U9111 (N_9111,N_8994,N_8563);
or U9112 (N_9112,N_8738,N_8583);
xor U9113 (N_9113,N_8659,N_8891);
xor U9114 (N_9114,N_8579,N_8811);
xor U9115 (N_9115,N_8954,N_8998);
and U9116 (N_9116,N_8670,N_8511);
nor U9117 (N_9117,N_8713,N_8657);
and U9118 (N_9118,N_8962,N_8892);
and U9119 (N_9119,N_8500,N_8717);
and U9120 (N_9120,N_8966,N_8540);
or U9121 (N_9121,N_8584,N_8792);
and U9122 (N_9122,N_8775,N_8865);
xnor U9123 (N_9123,N_8722,N_8991);
or U9124 (N_9124,N_8797,N_8609);
nor U9125 (N_9125,N_8606,N_8990);
nor U9126 (N_9126,N_8594,N_8890);
and U9127 (N_9127,N_8884,N_8809);
xor U9128 (N_9128,N_8854,N_8534);
xnor U9129 (N_9129,N_8870,N_8576);
nor U9130 (N_9130,N_8834,N_8504);
and U9131 (N_9131,N_8532,N_8641);
xnor U9132 (N_9132,N_8920,N_8943);
nand U9133 (N_9133,N_8885,N_8776);
nor U9134 (N_9134,N_8581,N_8881);
and U9135 (N_9135,N_8767,N_8678);
xnor U9136 (N_9136,N_8968,N_8849);
and U9137 (N_9137,N_8715,N_8734);
nand U9138 (N_9138,N_8539,N_8763);
and U9139 (N_9139,N_8508,N_8561);
and U9140 (N_9140,N_8972,N_8709);
xor U9141 (N_9141,N_8853,N_8820);
xor U9142 (N_9142,N_8625,N_8585);
nand U9143 (N_9143,N_8536,N_8898);
or U9144 (N_9144,N_8955,N_8570);
xnor U9145 (N_9145,N_8902,N_8559);
xnor U9146 (N_9146,N_8732,N_8696);
xor U9147 (N_9147,N_8989,N_8928);
and U9148 (N_9148,N_8981,N_8863);
nor U9149 (N_9149,N_8667,N_8635);
xnor U9150 (N_9150,N_8917,N_8941);
xnor U9151 (N_9151,N_8689,N_8664);
and U9152 (N_9152,N_8895,N_8676);
or U9153 (N_9153,N_8755,N_8694);
or U9154 (N_9154,N_8573,N_8602);
or U9155 (N_9155,N_8506,N_8771);
nand U9156 (N_9156,N_8693,N_8682);
nor U9157 (N_9157,N_8553,N_8805);
or U9158 (N_9158,N_8907,N_8600);
xor U9159 (N_9159,N_8619,N_8810);
nor U9160 (N_9160,N_8572,N_8899);
and U9161 (N_9161,N_8790,N_8872);
or U9162 (N_9162,N_8747,N_8813);
nor U9163 (N_9163,N_8605,N_8697);
nand U9164 (N_9164,N_8883,N_8597);
xnor U9165 (N_9165,N_8629,N_8577);
nor U9166 (N_9166,N_8575,N_8864);
xor U9167 (N_9167,N_8650,N_8723);
and U9168 (N_9168,N_8812,N_8783);
or U9169 (N_9169,N_8784,N_8525);
or U9170 (N_9170,N_8836,N_8886);
nor U9171 (N_9171,N_8714,N_8944);
nor U9172 (N_9172,N_8654,N_8904);
nor U9173 (N_9173,N_8832,N_8707);
nor U9174 (N_9174,N_8686,N_8958);
and U9175 (N_9175,N_8663,N_8567);
nand U9176 (N_9176,N_8746,N_8526);
and U9177 (N_9177,N_8564,N_8512);
xnor U9178 (N_9178,N_8578,N_8869);
or U9179 (N_9179,N_8965,N_8558);
or U9180 (N_9180,N_8628,N_8964);
nand U9181 (N_9181,N_8814,N_8829);
nor U9182 (N_9182,N_8683,N_8905);
and U9183 (N_9183,N_8698,N_8921);
and U9184 (N_9184,N_8857,N_8649);
nor U9185 (N_9185,N_8993,N_8712);
xor U9186 (N_9186,N_8589,N_8957);
and U9187 (N_9187,N_8774,N_8701);
and U9188 (N_9188,N_8982,N_8596);
nor U9189 (N_9189,N_8545,N_8786);
and U9190 (N_9190,N_8970,N_8825);
nor U9191 (N_9191,N_8521,N_8855);
nor U9192 (N_9192,N_8566,N_8889);
nand U9193 (N_9193,N_8887,N_8909);
nand U9194 (N_9194,N_8671,N_8824);
nand U9195 (N_9195,N_8821,N_8656);
nor U9196 (N_9196,N_8912,N_8985);
or U9197 (N_9197,N_8806,N_8856);
and U9198 (N_9198,N_8959,N_8535);
nand U9199 (N_9199,N_8926,N_8927);
nand U9200 (N_9200,N_8687,N_8627);
or U9201 (N_9201,N_8537,N_8901);
nor U9202 (N_9202,N_8924,N_8785);
xor U9203 (N_9203,N_8509,N_8833);
or U9204 (N_9204,N_8711,N_8638);
nor U9205 (N_9205,N_8835,N_8680);
or U9206 (N_9206,N_8929,N_8621);
or U9207 (N_9207,N_8725,N_8737);
xor U9208 (N_9208,N_8877,N_8615);
and U9209 (N_9209,N_8642,N_8569);
nor U9210 (N_9210,N_8951,N_8586);
or U9211 (N_9211,N_8544,N_8588);
or U9212 (N_9212,N_8538,N_8922);
nor U9213 (N_9213,N_8761,N_8950);
or U9214 (N_9214,N_8580,N_8618);
or U9215 (N_9215,N_8660,N_8942);
xor U9216 (N_9216,N_8935,N_8515);
xor U9217 (N_9217,N_8744,N_8948);
nand U9218 (N_9218,N_8529,N_8550);
xor U9219 (N_9219,N_8750,N_8617);
or U9220 (N_9220,N_8728,N_8624);
and U9221 (N_9221,N_8823,N_8751);
nor U9222 (N_9222,N_8930,N_8555);
or U9223 (N_9223,N_8612,N_8603);
and U9224 (N_9224,N_8758,N_8679);
nor U9225 (N_9225,N_8565,N_8655);
nand U9226 (N_9226,N_8807,N_8933);
nand U9227 (N_9227,N_8963,N_8938);
xor U9228 (N_9228,N_8880,N_8502);
xnor U9229 (N_9229,N_8787,N_8934);
and U9230 (N_9230,N_8513,N_8523);
or U9231 (N_9231,N_8541,N_8975);
nor U9232 (N_9232,N_8528,N_8645);
and U9233 (N_9233,N_8668,N_8772);
and U9234 (N_9234,N_8799,N_8548);
nand U9235 (N_9235,N_8730,N_8860);
xor U9236 (N_9236,N_8666,N_8520);
xnor U9237 (N_9237,N_8610,N_8841);
nor U9238 (N_9238,N_8765,N_8830);
nand U9239 (N_9239,N_8622,N_8599);
nor U9240 (N_9240,N_8524,N_8782);
or U9241 (N_9241,N_8706,N_8637);
xor U9242 (N_9242,N_8931,N_8607);
nor U9243 (N_9243,N_8897,N_8769);
or U9244 (N_9244,N_8595,N_8633);
or U9245 (N_9245,N_8936,N_8866);
or U9246 (N_9246,N_8986,N_8756);
xor U9247 (N_9247,N_8788,N_8726);
xor U9248 (N_9248,N_8647,N_8527);
and U9249 (N_9249,N_8630,N_8977);
nand U9250 (N_9250,N_8625,N_8688);
nand U9251 (N_9251,N_8754,N_8761);
nor U9252 (N_9252,N_8654,N_8746);
xnor U9253 (N_9253,N_8580,N_8726);
nor U9254 (N_9254,N_8534,N_8601);
and U9255 (N_9255,N_8634,N_8705);
nor U9256 (N_9256,N_8504,N_8968);
or U9257 (N_9257,N_8609,N_8863);
xnor U9258 (N_9258,N_8972,N_8594);
xnor U9259 (N_9259,N_8897,N_8878);
and U9260 (N_9260,N_8807,N_8592);
nor U9261 (N_9261,N_8527,N_8965);
nor U9262 (N_9262,N_8571,N_8781);
and U9263 (N_9263,N_8929,N_8546);
nor U9264 (N_9264,N_8820,N_8645);
or U9265 (N_9265,N_8571,N_8934);
xor U9266 (N_9266,N_8641,N_8716);
and U9267 (N_9267,N_8988,N_8555);
and U9268 (N_9268,N_8800,N_8938);
nor U9269 (N_9269,N_8758,N_8682);
or U9270 (N_9270,N_8588,N_8885);
xor U9271 (N_9271,N_8710,N_8836);
or U9272 (N_9272,N_8752,N_8773);
or U9273 (N_9273,N_8707,N_8734);
nor U9274 (N_9274,N_8597,N_8684);
nor U9275 (N_9275,N_8695,N_8514);
and U9276 (N_9276,N_8673,N_8741);
nor U9277 (N_9277,N_8971,N_8685);
and U9278 (N_9278,N_8994,N_8667);
and U9279 (N_9279,N_8809,N_8605);
and U9280 (N_9280,N_8875,N_8920);
nor U9281 (N_9281,N_8572,N_8871);
xor U9282 (N_9282,N_8614,N_8992);
or U9283 (N_9283,N_8566,N_8911);
xor U9284 (N_9284,N_8616,N_8885);
nand U9285 (N_9285,N_8848,N_8942);
and U9286 (N_9286,N_8800,N_8689);
nor U9287 (N_9287,N_8892,N_8903);
or U9288 (N_9288,N_8686,N_8874);
and U9289 (N_9289,N_8886,N_8864);
nor U9290 (N_9290,N_8632,N_8575);
nand U9291 (N_9291,N_8985,N_8676);
and U9292 (N_9292,N_8542,N_8975);
and U9293 (N_9293,N_8725,N_8546);
and U9294 (N_9294,N_8993,N_8794);
nand U9295 (N_9295,N_8865,N_8850);
xor U9296 (N_9296,N_8773,N_8961);
nand U9297 (N_9297,N_8808,N_8999);
or U9298 (N_9298,N_8586,N_8828);
and U9299 (N_9299,N_8812,N_8788);
nor U9300 (N_9300,N_8659,N_8877);
nand U9301 (N_9301,N_8602,N_8516);
nand U9302 (N_9302,N_8550,N_8518);
nand U9303 (N_9303,N_8736,N_8950);
nand U9304 (N_9304,N_8921,N_8753);
nand U9305 (N_9305,N_8827,N_8732);
nor U9306 (N_9306,N_8855,N_8918);
nor U9307 (N_9307,N_8596,N_8590);
nor U9308 (N_9308,N_8894,N_8678);
nand U9309 (N_9309,N_8697,N_8628);
and U9310 (N_9310,N_8743,N_8798);
nand U9311 (N_9311,N_8757,N_8514);
or U9312 (N_9312,N_8877,N_8699);
and U9313 (N_9313,N_8604,N_8743);
xor U9314 (N_9314,N_8543,N_8514);
nor U9315 (N_9315,N_8924,N_8933);
nor U9316 (N_9316,N_8992,N_8706);
nand U9317 (N_9317,N_8736,N_8791);
nor U9318 (N_9318,N_8600,N_8906);
nor U9319 (N_9319,N_8688,N_8554);
xor U9320 (N_9320,N_8840,N_8764);
and U9321 (N_9321,N_8714,N_8594);
xor U9322 (N_9322,N_8880,N_8809);
or U9323 (N_9323,N_8572,N_8914);
or U9324 (N_9324,N_8802,N_8785);
nor U9325 (N_9325,N_8922,N_8679);
nand U9326 (N_9326,N_8787,N_8960);
or U9327 (N_9327,N_8667,N_8650);
and U9328 (N_9328,N_8555,N_8923);
nor U9329 (N_9329,N_8932,N_8813);
and U9330 (N_9330,N_8580,N_8929);
xor U9331 (N_9331,N_8739,N_8762);
or U9332 (N_9332,N_8824,N_8999);
and U9333 (N_9333,N_8537,N_8918);
or U9334 (N_9334,N_8871,N_8710);
nor U9335 (N_9335,N_8831,N_8554);
nand U9336 (N_9336,N_8956,N_8613);
nand U9337 (N_9337,N_8787,N_8676);
xor U9338 (N_9338,N_8748,N_8700);
nor U9339 (N_9339,N_8961,N_8979);
xor U9340 (N_9340,N_8909,N_8705);
nand U9341 (N_9341,N_8530,N_8917);
or U9342 (N_9342,N_8913,N_8798);
nor U9343 (N_9343,N_8883,N_8615);
xor U9344 (N_9344,N_8850,N_8847);
and U9345 (N_9345,N_8756,N_8613);
and U9346 (N_9346,N_8739,N_8682);
or U9347 (N_9347,N_8905,N_8736);
and U9348 (N_9348,N_8749,N_8549);
and U9349 (N_9349,N_8742,N_8686);
or U9350 (N_9350,N_8993,N_8896);
nand U9351 (N_9351,N_8866,N_8585);
xor U9352 (N_9352,N_8504,N_8560);
or U9353 (N_9353,N_8754,N_8882);
or U9354 (N_9354,N_8621,N_8710);
xnor U9355 (N_9355,N_8917,N_8590);
nor U9356 (N_9356,N_8859,N_8892);
nor U9357 (N_9357,N_8787,N_8919);
xnor U9358 (N_9358,N_8708,N_8846);
xnor U9359 (N_9359,N_8730,N_8788);
or U9360 (N_9360,N_8593,N_8502);
nor U9361 (N_9361,N_8564,N_8946);
xor U9362 (N_9362,N_8550,N_8535);
nand U9363 (N_9363,N_8691,N_8548);
or U9364 (N_9364,N_8740,N_8730);
nand U9365 (N_9365,N_8804,N_8926);
or U9366 (N_9366,N_8797,N_8969);
nor U9367 (N_9367,N_8770,N_8718);
xor U9368 (N_9368,N_8684,N_8989);
xnor U9369 (N_9369,N_8669,N_8519);
nand U9370 (N_9370,N_8500,N_8877);
and U9371 (N_9371,N_8649,N_8620);
and U9372 (N_9372,N_8698,N_8704);
or U9373 (N_9373,N_8843,N_8872);
and U9374 (N_9374,N_8971,N_8589);
nand U9375 (N_9375,N_8803,N_8979);
nor U9376 (N_9376,N_8616,N_8990);
nand U9377 (N_9377,N_8575,N_8822);
nand U9378 (N_9378,N_8587,N_8816);
or U9379 (N_9379,N_8991,N_8961);
xor U9380 (N_9380,N_8972,N_8868);
or U9381 (N_9381,N_8786,N_8977);
xnor U9382 (N_9382,N_8732,N_8935);
nor U9383 (N_9383,N_8889,N_8934);
and U9384 (N_9384,N_8628,N_8645);
nor U9385 (N_9385,N_8712,N_8760);
and U9386 (N_9386,N_8727,N_8522);
and U9387 (N_9387,N_8821,N_8780);
xor U9388 (N_9388,N_8574,N_8521);
and U9389 (N_9389,N_8712,N_8571);
or U9390 (N_9390,N_8515,N_8810);
xor U9391 (N_9391,N_8738,N_8722);
or U9392 (N_9392,N_8829,N_8587);
or U9393 (N_9393,N_8616,N_8634);
xnor U9394 (N_9394,N_8892,N_8543);
xnor U9395 (N_9395,N_8682,N_8784);
or U9396 (N_9396,N_8849,N_8544);
nor U9397 (N_9397,N_8982,N_8760);
nand U9398 (N_9398,N_8938,N_8914);
nor U9399 (N_9399,N_8904,N_8836);
or U9400 (N_9400,N_8644,N_8650);
nor U9401 (N_9401,N_8731,N_8804);
xnor U9402 (N_9402,N_8824,N_8770);
nand U9403 (N_9403,N_8675,N_8720);
or U9404 (N_9404,N_8811,N_8814);
or U9405 (N_9405,N_8655,N_8576);
and U9406 (N_9406,N_8888,N_8645);
nand U9407 (N_9407,N_8524,N_8730);
nand U9408 (N_9408,N_8658,N_8794);
xor U9409 (N_9409,N_8790,N_8987);
xnor U9410 (N_9410,N_8941,N_8884);
and U9411 (N_9411,N_8874,N_8876);
and U9412 (N_9412,N_8659,N_8709);
nand U9413 (N_9413,N_8525,N_8549);
nor U9414 (N_9414,N_8747,N_8733);
and U9415 (N_9415,N_8837,N_8708);
nand U9416 (N_9416,N_8594,N_8848);
nor U9417 (N_9417,N_8900,N_8653);
xor U9418 (N_9418,N_8704,N_8869);
and U9419 (N_9419,N_8785,N_8554);
xor U9420 (N_9420,N_8651,N_8896);
nor U9421 (N_9421,N_8893,N_8611);
nor U9422 (N_9422,N_8878,N_8863);
or U9423 (N_9423,N_8851,N_8956);
nor U9424 (N_9424,N_8717,N_8748);
or U9425 (N_9425,N_8656,N_8797);
xor U9426 (N_9426,N_8971,N_8967);
and U9427 (N_9427,N_8805,N_8648);
nand U9428 (N_9428,N_8569,N_8906);
and U9429 (N_9429,N_8875,N_8672);
xor U9430 (N_9430,N_8607,N_8617);
nor U9431 (N_9431,N_8947,N_8826);
or U9432 (N_9432,N_8852,N_8739);
nand U9433 (N_9433,N_8903,N_8630);
and U9434 (N_9434,N_8911,N_8961);
nand U9435 (N_9435,N_8622,N_8839);
and U9436 (N_9436,N_8600,N_8872);
nand U9437 (N_9437,N_8958,N_8590);
xor U9438 (N_9438,N_8666,N_8824);
nor U9439 (N_9439,N_8761,N_8999);
nor U9440 (N_9440,N_8508,N_8819);
or U9441 (N_9441,N_8668,N_8940);
or U9442 (N_9442,N_8919,N_8976);
xor U9443 (N_9443,N_8623,N_8568);
nand U9444 (N_9444,N_8567,N_8929);
and U9445 (N_9445,N_8675,N_8986);
xnor U9446 (N_9446,N_8637,N_8713);
xor U9447 (N_9447,N_8594,N_8771);
xor U9448 (N_9448,N_8678,N_8668);
or U9449 (N_9449,N_8661,N_8827);
or U9450 (N_9450,N_8591,N_8876);
and U9451 (N_9451,N_8513,N_8964);
xor U9452 (N_9452,N_8768,N_8767);
nand U9453 (N_9453,N_8938,N_8602);
or U9454 (N_9454,N_8931,N_8949);
nor U9455 (N_9455,N_8691,N_8678);
nor U9456 (N_9456,N_8535,N_8588);
xnor U9457 (N_9457,N_8935,N_8842);
and U9458 (N_9458,N_8904,N_8869);
nand U9459 (N_9459,N_8643,N_8555);
xor U9460 (N_9460,N_8864,N_8882);
nor U9461 (N_9461,N_8516,N_8850);
nor U9462 (N_9462,N_8719,N_8965);
nor U9463 (N_9463,N_8680,N_8901);
nor U9464 (N_9464,N_8922,N_8891);
and U9465 (N_9465,N_8819,N_8998);
nor U9466 (N_9466,N_8520,N_8614);
or U9467 (N_9467,N_8626,N_8578);
nand U9468 (N_9468,N_8777,N_8733);
nand U9469 (N_9469,N_8871,N_8962);
and U9470 (N_9470,N_8501,N_8866);
nand U9471 (N_9471,N_8796,N_8763);
or U9472 (N_9472,N_8615,N_8681);
or U9473 (N_9473,N_8741,N_8592);
nor U9474 (N_9474,N_8545,N_8995);
xnor U9475 (N_9475,N_8768,N_8708);
xnor U9476 (N_9476,N_8652,N_8675);
or U9477 (N_9477,N_8618,N_8710);
nand U9478 (N_9478,N_8664,N_8718);
and U9479 (N_9479,N_8613,N_8867);
nand U9480 (N_9480,N_8658,N_8511);
or U9481 (N_9481,N_8624,N_8760);
nand U9482 (N_9482,N_8578,N_8799);
or U9483 (N_9483,N_8747,N_8728);
nand U9484 (N_9484,N_8880,N_8946);
nor U9485 (N_9485,N_8641,N_8823);
and U9486 (N_9486,N_8777,N_8523);
and U9487 (N_9487,N_8953,N_8509);
or U9488 (N_9488,N_8728,N_8957);
or U9489 (N_9489,N_8701,N_8572);
xor U9490 (N_9490,N_8826,N_8679);
nand U9491 (N_9491,N_8536,N_8595);
nor U9492 (N_9492,N_8820,N_8622);
or U9493 (N_9493,N_8896,N_8755);
nor U9494 (N_9494,N_8986,N_8596);
or U9495 (N_9495,N_8539,N_8796);
nor U9496 (N_9496,N_8802,N_8553);
nor U9497 (N_9497,N_8920,N_8819);
and U9498 (N_9498,N_8893,N_8664);
nand U9499 (N_9499,N_8798,N_8839);
or U9500 (N_9500,N_9404,N_9417);
nor U9501 (N_9501,N_9004,N_9012);
nand U9502 (N_9502,N_9364,N_9219);
nand U9503 (N_9503,N_9406,N_9422);
xor U9504 (N_9504,N_9427,N_9397);
and U9505 (N_9505,N_9450,N_9252);
or U9506 (N_9506,N_9069,N_9129);
xor U9507 (N_9507,N_9289,N_9437);
and U9508 (N_9508,N_9061,N_9368);
xnor U9509 (N_9509,N_9292,N_9043);
xnor U9510 (N_9510,N_9392,N_9466);
and U9511 (N_9511,N_9396,N_9463);
xor U9512 (N_9512,N_9309,N_9363);
nand U9513 (N_9513,N_9275,N_9373);
nor U9514 (N_9514,N_9193,N_9314);
nor U9515 (N_9515,N_9443,N_9105);
nor U9516 (N_9516,N_9197,N_9490);
xor U9517 (N_9517,N_9222,N_9032);
nand U9518 (N_9518,N_9305,N_9464);
nand U9519 (N_9519,N_9224,N_9018);
nor U9520 (N_9520,N_9452,N_9474);
nor U9521 (N_9521,N_9489,N_9117);
xor U9522 (N_9522,N_9050,N_9232);
xnor U9523 (N_9523,N_9174,N_9405);
nor U9524 (N_9524,N_9070,N_9107);
nand U9525 (N_9525,N_9272,N_9391);
or U9526 (N_9526,N_9451,N_9435);
xor U9527 (N_9527,N_9191,N_9058);
nand U9528 (N_9528,N_9449,N_9189);
xor U9529 (N_9529,N_9462,N_9277);
nand U9530 (N_9530,N_9166,N_9036);
or U9531 (N_9531,N_9425,N_9412);
and U9532 (N_9532,N_9182,N_9374);
and U9533 (N_9533,N_9125,N_9065);
or U9534 (N_9534,N_9134,N_9100);
nor U9535 (N_9535,N_9457,N_9481);
nor U9536 (N_9536,N_9256,N_9083);
or U9537 (N_9537,N_9271,N_9144);
or U9538 (N_9538,N_9328,N_9455);
and U9539 (N_9539,N_9122,N_9343);
nor U9540 (N_9540,N_9084,N_9044);
xor U9541 (N_9541,N_9110,N_9283);
xor U9542 (N_9542,N_9319,N_9133);
nand U9543 (N_9543,N_9408,N_9006);
nor U9544 (N_9544,N_9145,N_9411);
or U9545 (N_9545,N_9045,N_9211);
and U9546 (N_9546,N_9312,N_9048);
nand U9547 (N_9547,N_9354,N_9431);
and U9548 (N_9548,N_9262,N_9170);
xor U9549 (N_9549,N_9113,N_9313);
nand U9550 (N_9550,N_9241,N_9217);
nor U9551 (N_9551,N_9028,N_9395);
xnor U9552 (N_9552,N_9302,N_9274);
nor U9553 (N_9553,N_9239,N_9168);
xnor U9554 (N_9554,N_9049,N_9259);
or U9555 (N_9555,N_9321,N_9088);
and U9556 (N_9556,N_9495,N_9155);
and U9557 (N_9557,N_9024,N_9229);
or U9558 (N_9558,N_9162,N_9177);
or U9559 (N_9559,N_9441,N_9094);
nand U9560 (N_9560,N_9142,N_9424);
and U9561 (N_9561,N_9031,N_9114);
or U9562 (N_9562,N_9325,N_9423);
xnor U9563 (N_9563,N_9221,N_9086);
and U9564 (N_9564,N_9051,N_9152);
nor U9565 (N_9565,N_9357,N_9442);
xor U9566 (N_9566,N_9301,N_9027);
nor U9567 (N_9567,N_9019,N_9184);
xnor U9568 (N_9568,N_9258,N_9469);
nor U9569 (N_9569,N_9087,N_9073);
xnor U9570 (N_9570,N_9327,N_9478);
xnor U9571 (N_9571,N_9254,N_9208);
xor U9572 (N_9572,N_9226,N_9215);
xor U9573 (N_9573,N_9410,N_9293);
nor U9574 (N_9574,N_9351,N_9295);
and U9575 (N_9575,N_9360,N_9388);
or U9576 (N_9576,N_9488,N_9035);
or U9577 (N_9577,N_9244,N_9186);
or U9578 (N_9578,N_9336,N_9333);
or U9579 (N_9579,N_9160,N_9493);
or U9580 (N_9580,N_9276,N_9383);
nand U9581 (N_9581,N_9130,N_9334);
nor U9582 (N_9582,N_9230,N_9362);
or U9583 (N_9583,N_9118,N_9057);
nand U9584 (N_9584,N_9367,N_9338);
or U9585 (N_9585,N_9248,N_9220);
and U9586 (N_9586,N_9278,N_9267);
xnor U9587 (N_9587,N_9287,N_9445);
and U9588 (N_9588,N_9060,N_9151);
nor U9589 (N_9589,N_9456,N_9298);
xnor U9590 (N_9590,N_9382,N_9253);
nand U9591 (N_9591,N_9029,N_9461);
and U9592 (N_9592,N_9378,N_9156);
and U9593 (N_9593,N_9240,N_9420);
nand U9594 (N_9594,N_9340,N_9030);
or U9595 (N_9595,N_9085,N_9310);
or U9596 (N_9596,N_9096,N_9010);
xnor U9597 (N_9597,N_9480,N_9415);
and U9598 (N_9598,N_9007,N_9161);
xnor U9599 (N_9599,N_9263,N_9121);
and U9600 (N_9600,N_9470,N_9297);
xnor U9601 (N_9601,N_9243,N_9195);
xnor U9602 (N_9602,N_9013,N_9047);
nor U9603 (N_9603,N_9381,N_9273);
nand U9604 (N_9604,N_9475,N_9175);
and U9605 (N_9605,N_9074,N_9499);
xor U9606 (N_9606,N_9486,N_9089);
or U9607 (N_9607,N_9270,N_9201);
or U9608 (N_9608,N_9426,N_9136);
nor U9609 (N_9609,N_9320,N_9339);
and U9610 (N_9610,N_9235,N_9353);
or U9611 (N_9611,N_9356,N_9326);
nor U9612 (N_9612,N_9448,N_9337);
nor U9613 (N_9613,N_9202,N_9400);
or U9614 (N_9614,N_9076,N_9150);
and U9615 (N_9615,N_9147,N_9465);
or U9616 (N_9616,N_9119,N_9056);
xor U9617 (N_9617,N_9251,N_9139);
or U9618 (N_9618,N_9438,N_9279);
nor U9619 (N_9619,N_9228,N_9386);
or U9620 (N_9620,N_9370,N_9023);
nor U9621 (N_9621,N_9482,N_9346);
or U9622 (N_9622,N_9288,N_9454);
nor U9623 (N_9623,N_9436,N_9242);
nand U9624 (N_9624,N_9419,N_9233);
and U9625 (N_9625,N_9214,N_9433);
nand U9626 (N_9626,N_9483,N_9015);
and U9627 (N_9627,N_9323,N_9106);
and U9628 (N_9628,N_9471,N_9005);
and U9629 (N_9629,N_9183,N_9000);
or U9630 (N_9630,N_9429,N_9257);
or U9631 (N_9631,N_9385,N_9245);
or U9632 (N_9632,N_9380,N_9052);
nor U9633 (N_9633,N_9033,N_9393);
nand U9634 (N_9634,N_9223,N_9163);
or U9635 (N_9635,N_9308,N_9188);
and U9636 (N_9636,N_9141,N_9318);
xor U9637 (N_9637,N_9476,N_9154);
nand U9638 (N_9638,N_9020,N_9341);
xnor U9639 (N_9639,N_9081,N_9039);
xor U9640 (N_9640,N_9053,N_9042);
xnor U9641 (N_9641,N_9095,N_9112);
or U9642 (N_9642,N_9091,N_9284);
xor U9643 (N_9643,N_9187,N_9484);
xor U9644 (N_9644,N_9153,N_9205);
or U9645 (N_9645,N_9037,N_9440);
nand U9646 (N_9646,N_9067,N_9260);
nor U9647 (N_9647,N_9104,N_9428);
nand U9648 (N_9648,N_9082,N_9294);
nor U9649 (N_9649,N_9377,N_9280);
and U9650 (N_9650,N_9286,N_9255);
and U9651 (N_9651,N_9296,N_9331);
xnor U9652 (N_9652,N_9204,N_9250);
nor U9653 (N_9653,N_9485,N_9054);
or U9654 (N_9654,N_9164,N_9180);
or U9655 (N_9655,N_9332,N_9172);
and U9656 (N_9656,N_9398,N_9190);
nand U9657 (N_9657,N_9330,N_9498);
nand U9658 (N_9658,N_9358,N_9021);
nor U9659 (N_9659,N_9376,N_9306);
nor U9660 (N_9660,N_9290,N_9355);
nor U9661 (N_9661,N_9025,N_9022);
xor U9662 (N_9662,N_9079,N_9496);
xnor U9663 (N_9663,N_9098,N_9185);
and U9664 (N_9664,N_9046,N_9238);
nor U9665 (N_9665,N_9008,N_9348);
or U9666 (N_9666,N_9369,N_9102);
nand U9667 (N_9667,N_9101,N_9322);
or U9668 (N_9668,N_9432,N_9111);
or U9669 (N_9669,N_9418,N_9268);
or U9670 (N_9670,N_9361,N_9146);
nor U9671 (N_9671,N_9131,N_9207);
xnor U9672 (N_9672,N_9059,N_9090);
xnor U9673 (N_9673,N_9300,N_9324);
xor U9674 (N_9674,N_9209,N_9103);
nand U9675 (N_9675,N_9169,N_9062);
xnor U9676 (N_9676,N_9066,N_9158);
nand U9677 (N_9677,N_9194,N_9140);
or U9678 (N_9678,N_9307,N_9316);
and U9679 (N_9679,N_9116,N_9179);
nand U9680 (N_9680,N_9446,N_9165);
xnor U9681 (N_9681,N_9315,N_9199);
nand U9682 (N_9682,N_9213,N_9210);
nor U9683 (N_9683,N_9265,N_9206);
nor U9684 (N_9684,N_9421,N_9135);
nor U9685 (N_9685,N_9212,N_9345);
nand U9686 (N_9686,N_9472,N_9138);
nor U9687 (N_9687,N_9366,N_9123);
nand U9688 (N_9688,N_9402,N_9137);
or U9689 (N_9689,N_9040,N_9409);
xor U9690 (N_9690,N_9200,N_9414);
nand U9691 (N_9691,N_9269,N_9371);
nor U9692 (N_9692,N_9071,N_9093);
nor U9693 (N_9693,N_9120,N_9477);
nor U9694 (N_9694,N_9291,N_9092);
xnor U9695 (N_9695,N_9473,N_9157);
and U9696 (N_9696,N_9487,N_9080);
nor U9697 (N_9697,N_9299,N_9064);
nand U9698 (N_9698,N_9231,N_9178);
nand U9699 (N_9699,N_9261,N_9359);
nor U9700 (N_9700,N_9342,N_9394);
and U9701 (N_9701,N_9497,N_9001);
xor U9702 (N_9702,N_9109,N_9132);
or U9703 (N_9703,N_9365,N_9011);
xor U9704 (N_9704,N_9126,N_9491);
nand U9705 (N_9705,N_9492,N_9460);
nand U9706 (N_9706,N_9401,N_9329);
or U9707 (N_9707,N_9034,N_9143);
nand U9708 (N_9708,N_9003,N_9176);
nand U9709 (N_9709,N_9203,N_9017);
or U9710 (N_9710,N_9372,N_9072);
nand U9711 (N_9711,N_9458,N_9171);
nand U9712 (N_9712,N_9055,N_9068);
nor U9713 (N_9713,N_9075,N_9416);
or U9714 (N_9714,N_9249,N_9077);
nor U9715 (N_9715,N_9246,N_9108);
nand U9716 (N_9716,N_9281,N_9127);
nor U9717 (N_9717,N_9009,N_9403);
and U9718 (N_9718,N_9459,N_9379);
nand U9719 (N_9719,N_9434,N_9317);
xnor U9720 (N_9720,N_9303,N_9344);
or U9721 (N_9721,N_9399,N_9063);
and U9722 (N_9722,N_9349,N_9467);
nand U9723 (N_9723,N_9016,N_9198);
and U9724 (N_9724,N_9192,N_9430);
nor U9725 (N_9725,N_9468,N_9128);
xnor U9726 (N_9726,N_9375,N_9350);
nor U9727 (N_9727,N_9413,N_9439);
nand U9728 (N_9728,N_9264,N_9352);
or U9729 (N_9729,N_9247,N_9304);
nand U9730 (N_9730,N_9384,N_9196);
nor U9731 (N_9731,N_9026,N_9173);
and U9732 (N_9732,N_9218,N_9237);
nand U9733 (N_9733,N_9234,N_9447);
nor U9734 (N_9734,N_9014,N_9389);
xor U9735 (N_9735,N_9167,N_9002);
and U9736 (N_9736,N_9216,N_9311);
and U9737 (N_9737,N_9097,N_9124);
or U9738 (N_9738,N_9227,N_9078);
nand U9739 (N_9739,N_9494,N_9181);
xor U9740 (N_9740,N_9390,N_9453);
or U9741 (N_9741,N_9266,N_9159);
and U9742 (N_9742,N_9387,N_9407);
xnor U9743 (N_9743,N_9225,N_9285);
and U9744 (N_9744,N_9282,N_9347);
or U9745 (N_9745,N_9148,N_9444);
nor U9746 (N_9746,N_9479,N_9149);
nand U9747 (N_9747,N_9115,N_9041);
xor U9748 (N_9748,N_9038,N_9099);
and U9749 (N_9749,N_9335,N_9236);
and U9750 (N_9750,N_9282,N_9023);
nor U9751 (N_9751,N_9338,N_9053);
nor U9752 (N_9752,N_9054,N_9343);
xor U9753 (N_9753,N_9169,N_9254);
or U9754 (N_9754,N_9239,N_9146);
nor U9755 (N_9755,N_9004,N_9091);
or U9756 (N_9756,N_9271,N_9385);
or U9757 (N_9757,N_9313,N_9017);
and U9758 (N_9758,N_9230,N_9037);
nand U9759 (N_9759,N_9137,N_9429);
xor U9760 (N_9760,N_9333,N_9080);
nor U9761 (N_9761,N_9204,N_9017);
xnor U9762 (N_9762,N_9115,N_9418);
xnor U9763 (N_9763,N_9275,N_9060);
or U9764 (N_9764,N_9265,N_9101);
xnor U9765 (N_9765,N_9076,N_9255);
and U9766 (N_9766,N_9474,N_9424);
nand U9767 (N_9767,N_9390,N_9414);
nor U9768 (N_9768,N_9075,N_9258);
nor U9769 (N_9769,N_9174,N_9008);
nor U9770 (N_9770,N_9304,N_9186);
and U9771 (N_9771,N_9179,N_9068);
xor U9772 (N_9772,N_9012,N_9192);
and U9773 (N_9773,N_9309,N_9453);
and U9774 (N_9774,N_9219,N_9410);
nor U9775 (N_9775,N_9391,N_9197);
nand U9776 (N_9776,N_9056,N_9386);
nor U9777 (N_9777,N_9372,N_9463);
xor U9778 (N_9778,N_9243,N_9328);
nor U9779 (N_9779,N_9162,N_9246);
nor U9780 (N_9780,N_9088,N_9482);
nor U9781 (N_9781,N_9127,N_9464);
nand U9782 (N_9782,N_9491,N_9270);
xnor U9783 (N_9783,N_9197,N_9489);
and U9784 (N_9784,N_9377,N_9120);
or U9785 (N_9785,N_9301,N_9494);
nor U9786 (N_9786,N_9283,N_9049);
xnor U9787 (N_9787,N_9189,N_9017);
xnor U9788 (N_9788,N_9430,N_9123);
or U9789 (N_9789,N_9019,N_9390);
or U9790 (N_9790,N_9267,N_9167);
or U9791 (N_9791,N_9491,N_9297);
nor U9792 (N_9792,N_9129,N_9278);
nor U9793 (N_9793,N_9485,N_9497);
nor U9794 (N_9794,N_9445,N_9307);
and U9795 (N_9795,N_9283,N_9033);
and U9796 (N_9796,N_9053,N_9072);
and U9797 (N_9797,N_9305,N_9479);
and U9798 (N_9798,N_9157,N_9329);
xor U9799 (N_9799,N_9020,N_9485);
xnor U9800 (N_9800,N_9475,N_9264);
and U9801 (N_9801,N_9052,N_9021);
or U9802 (N_9802,N_9239,N_9357);
and U9803 (N_9803,N_9308,N_9439);
xnor U9804 (N_9804,N_9297,N_9159);
and U9805 (N_9805,N_9359,N_9035);
nor U9806 (N_9806,N_9032,N_9344);
or U9807 (N_9807,N_9457,N_9343);
xor U9808 (N_9808,N_9463,N_9072);
xnor U9809 (N_9809,N_9371,N_9442);
xor U9810 (N_9810,N_9424,N_9438);
nor U9811 (N_9811,N_9487,N_9185);
nand U9812 (N_9812,N_9200,N_9424);
nor U9813 (N_9813,N_9366,N_9373);
or U9814 (N_9814,N_9086,N_9387);
nand U9815 (N_9815,N_9408,N_9452);
or U9816 (N_9816,N_9493,N_9323);
xor U9817 (N_9817,N_9384,N_9012);
and U9818 (N_9818,N_9493,N_9437);
or U9819 (N_9819,N_9402,N_9384);
or U9820 (N_9820,N_9425,N_9413);
and U9821 (N_9821,N_9219,N_9207);
or U9822 (N_9822,N_9252,N_9394);
and U9823 (N_9823,N_9033,N_9057);
nor U9824 (N_9824,N_9062,N_9386);
and U9825 (N_9825,N_9280,N_9365);
nor U9826 (N_9826,N_9316,N_9448);
nor U9827 (N_9827,N_9351,N_9368);
xor U9828 (N_9828,N_9400,N_9451);
and U9829 (N_9829,N_9021,N_9057);
and U9830 (N_9830,N_9460,N_9040);
xnor U9831 (N_9831,N_9210,N_9350);
nor U9832 (N_9832,N_9209,N_9242);
or U9833 (N_9833,N_9495,N_9095);
or U9834 (N_9834,N_9319,N_9180);
nand U9835 (N_9835,N_9049,N_9173);
nand U9836 (N_9836,N_9478,N_9369);
or U9837 (N_9837,N_9052,N_9458);
xor U9838 (N_9838,N_9432,N_9112);
nor U9839 (N_9839,N_9069,N_9335);
xnor U9840 (N_9840,N_9241,N_9465);
xnor U9841 (N_9841,N_9144,N_9473);
and U9842 (N_9842,N_9305,N_9141);
or U9843 (N_9843,N_9472,N_9208);
or U9844 (N_9844,N_9092,N_9198);
xnor U9845 (N_9845,N_9153,N_9397);
nor U9846 (N_9846,N_9363,N_9416);
nor U9847 (N_9847,N_9495,N_9201);
xnor U9848 (N_9848,N_9385,N_9129);
or U9849 (N_9849,N_9370,N_9329);
nand U9850 (N_9850,N_9154,N_9152);
or U9851 (N_9851,N_9100,N_9444);
nand U9852 (N_9852,N_9181,N_9094);
xor U9853 (N_9853,N_9332,N_9257);
xor U9854 (N_9854,N_9450,N_9347);
nor U9855 (N_9855,N_9137,N_9225);
nor U9856 (N_9856,N_9021,N_9162);
xnor U9857 (N_9857,N_9088,N_9276);
or U9858 (N_9858,N_9425,N_9239);
nand U9859 (N_9859,N_9432,N_9199);
and U9860 (N_9860,N_9015,N_9485);
and U9861 (N_9861,N_9042,N_9440);
nand U9862 (N_9862,N_9160,N_9180);
and U9863 (N_9863,N_9485,N_9470);
xnor U9864 (N_9864,N_9407,N_9404);
nand U9865 (N_9865,N_9095,N_9146);
nor U9866 (N_9866,N_9064,N_9090);
and U9867 (N_9867,N_9142,N_9253);
or U9868 (N_9868,N_9442,N_9027);
and U9869 (N_9869,N_9219,N_9137);
nand U9870 (N_9870,N_9431,N_9014);
or U9871 (N_9871,N_9092,N_9040);
and U9872 (N_9872,N_9348,N_9470);
nand U9873 (N_9873,N_9025,N_9486);
nand U9874 (N_9874,N_9109,N_9328);
or U9875 (N_9875,N_9175,N_9213);
or U9876 (N_9876,N_9279,N_9387);
or U9877 (N_9877,N_9448,N_9048);
or U9878 (N_9878,N_9274,N_9413);
and U9879 (N_9879,N_9321,N_9202);
nand U9880 (N_9880,N_9134,N_9046);
and U9881 (N_9881,N_9494,N_9466);
nand U9882 (N_9882,N_9332,N_9247);
or U9883 (N_9883,N_9196,N_9037);
nor U9884 (N_9884,N_9011,N_9426);
or U9885 (N_9885,N_9348,N_9089);
nand U9886 (N_9886,N_9226,N_9200);
and U9887 (N_9887,N_9347,N_9072);
or U9888 (N_9888,N_9420,N_9096);
and U9889 (N_9889,N_9408,N_9474);
or U9890 (N_9890,N_9333,N_9259);
and U9891 (N_9891,N_9499,N_9322);
nand U9892 (N_9892,N_9249,N_9003);
and U9893 (N_9893,N_9454,N_9329);
or U9894 (N_9894,N_9166,N_9411);
and U9895 (N_9895,N_9047,N_9070);
and U9896 (N_9896,N_9446,N_9133);
nor U9897 (N_9897,N_9443,N_9021);
and U9898 (N_9898,N_9216,N_9387);
nand U9899 (N_9899,N_9257,N_9106);
and U9900 (N_9900,N_9342,N_9448);
and U9901 (N_9901,N_9475,N_9142);
nand U9902 (N_9902,N_9460,N_9269);
nand U9903 (N_9903,N_9454,N_9133);
nand U9904 (N_9904,N_9417,N_9435);
or U9905 (N_9905,N_9486,N_9261);
nor U9906 (N_9906,N_9224,N_9358);
nor U9907 (N_9907,N_9129,N_9032);
or U9908 (N_9908,N_9454,N_9433);
nand U9909 (N_9909,N_9144,N_9038);
xnor U9910 (N_9910,N_9336,N_9435);
and U9911 (N_9911,N_9181,N_9431);
nor U9912 (N_9912,N_9372,N_9257);
nor U9913 (N_9913,N_9031,N_9357);
nand U9914 (N_9914,N_9027,N_9139);
nor U9915 (N_9915,N_9472,N_9159);
nand U9916 (N_9916,N_9085,N_9306);
and U9917 (N_9917,N_9036,N_9097);
nand U9918 (N_9918,N_9188,N_9449);
nor U9919 (N_9919,N_9300,N_9468);
or U9920 (N_9920,N_9053,N_9404);
nor U9921 (N_9921,N_9363,N_9100);
nand U9922 (N_9922,N_9467,N_9354);
or U9923 (N_9923,N_9324,N_9342);
and U9924 (N_9924,N_9307,N_9174);
nand U9925 (N_9925,N_9247,N_9475);
xor U9926 (N_9926,N_9053,N_9496);
xor U9927 (N_9927,N_9204,N_9492);
nand U9928 (N_9928,N_9114,N_9301);
xor U9929 (N_9929,N_9247,N_9241);
xnor U9930 (N_9930,N_9048,N_9033);
xor U9931 (N_9931,N_9325,N_9335);
or U9932 (N_9932,N_9395,N_9352);
or U9933 (N_9933,N_9001,N_9084);
nor U9934 (N_9934,N_9217,N_9286);
and U9935 (N_9935,N_9043,N_9080);
xnor U9936 (N_9936,N_9206,N_9379);
nor U9937 (N_9937,N_9088,N_9278);
nor U9938 (N_9938,N_9361,N_9083);
nor U9939 (N_9939,N_9367,N_9176);
or U9940 (N_9940,N_9428,N_9297);
and U9941 (N_9941,N_9073,N_9212);
xor U9942 (N_9942,N_9028,N_9052);
nor U9943 (N_9943,N_9101,N_9362);
and U9944 (N_9944,N_9445,N_9497);
and U9945 (N_9945,N_9183,N_9445);
xor U9946 (N_9946,N_9486,N_9237);
or U9947 (N_9947,N_9367,N_9187);
and U9948 (N_9948,N_9384,N_9420);
xnor U9949 (N_9949,N_9058,N_9090);
nand U9950 (N_9950,N_9459,N_9377);
nand U9951 (N_9951,N_9321,N_9268);
and U9952 (N_9952,N_9086,N_9480);
or U9953 (N_9953,N_9432,N_9216);
nor U9954 (N_9954,N_9171,N_9075);
and U9955 (N_9955,N_9385,N_9098);
nand U9956 (N_9956,N_9336,N_9292);
nor U9957 (N_9957,N_9348,N_9314);
or U9958 (N_9958,N_9040,N_9158);
nor U9959 (N_9959,N_9356,N_9172);
xnor U9960 (N_9960,N_9333,N_9230);
nor U9961 (N_9961,N_9188,N_9143);
nand U9962 (N_9962,N_9243,N_9439);
or U9963 (N_9963,N_9447,N_9164);
or U9964 (N_9964,N_9219,N_9101);
xnor U9965 (N_9965,N_9463,N_9009);
nand U9966 (N_9966,N_9168,N_9408);
or U9967 (N_9967,N_9008,N_9043);
nand U9968 (N_9968,N_9449,N_9430);
nand U9969 (N_9969,N_9212,N_9215);
xor U9970 (N_9970,N_9020,N_9460);
xor U9971 (N_9971,N_9490,N_9210);
or U9972 (N_9972,N_9240,N_9499);
xnor U9973 (N_9973,N_9325,N_9042);
and U9974 (N_9974,N_9463,N_9322);
and U9975 (N_9975,N_9499,N_9283);
nor U9976 (N_9976,N_9049,N_9258);
nor U9977 (N_9977,N_9177,N_9302);
nor U9978 (N_9978,N_9253,N_9375);
nand U9979 (N_9979,N_9213,N_9431);
or U9980 (N_9980,N_9214,N_9467);
nor U9981 (N_9981,N_9096,N_9423);
and U9982 (N_9982,N_9069,N_9132);
nor U9983 (N_9983,N_9377,N_9172);
xor U9984 (N_9984,N_9492,N_9179);
nor U9985 (N_9985,N_9448,N_9013);
nand U9986 (N_9986,N_9271,N_9124);
nor U9987 (N_9987,N_9319,N_9074);
xor U9988 (N_9988,N_9248,N_9316);
xnor U9989 (N_9989,N_9441,N_9127);
nor U9990 (N_9990,N_9376,N_9457);
nor U9991 (N_9991,N_9194,N_9100);
xor U9992 (N_9992,N_9284,N_9157);
and U9993 (N_9993,N_9474,N_9491);
nand U9994 (N_9994,N_9215,N_9412);
nand U9995 (N_9995,N_9106,N_9226);
nand U9996 (N_9996,N_9200,N_9020);
xor U9997 (N_9997,N_9371,N_9446);
and U9998 (N_9998,N_9286,N_9010);
and U9999 (N_9999,N_9140,N_9203);
xnor U10000 (N_10000,N_9952,N_9900);
nand U10001 (N_10001,N_9751,N_9533);
xnor U10002 (N_10002,N_9595,N_9649);
nor U10003 (N_10003,N_9780,N_9733);
xnor U10004 (N_10004,N_9979,N_9862);
xnor U10005 (N_10005,N_9564,N_9870);
nand U10006 (N_10006,N_9568,N_9963);
and U10007 (N_10007,N_9508,N_9708);
or U10008 (N_10008,N_9597,N_9841);
nand U10009 (N_10009,N_9777,N_9662);
nand U10010 (N_10010,N_9660,N_9556);
nor U10011 (N_10011,N_9676,N_9947);
or U10012 (N_10012,N_9656,N_9987);
or U10013 (N_10013,N_9745,N_9640);
and U10014 (N_10014,N_9557,N_9522);
nor U10015 (N_10015,N_9699,N_9525);
nor U10016 (N_10016,N_9757,N_9796);
and U10017 (N_10017,N_9827,N_9726);
nand U10018 (N_10018,N_9860,N_9927);
nor U10019 (N_10019,N_9546,N_9946);
and U10020 (N_10020,N_9545,N_9630);
and U10021 (N_10021,N_9942,N_9552);
nand U10022 (N_10022,N_9550,N_9848);
xor U10023 (N_10023,N_9888,N_9526);
or U10024 (N_10024,N_9746,N_9961);
or U10025 (N_10025,N_9811,N_9655);
and U10026 (N_10026,N_9933,N_9850);
and U10027 (N_10027,N_9750,N_9866);
xor U10028 (N_10028,N_9554,N_9609);
nor U10029 (N_10029,N_9898,N_9964);
nand U10030 (N_10030,N_9578,N_9603);
xnor U10031 (N_10031,N_9692,N_9734);
and U10032 (N_10032,N_9955,N_9853);
or U10033 (N_10033,N_9754,N_9969);
nor U10034 (N_10034,N_9984,N_9803);
and U10035 (N_10035,N_9779,N_9698);
or U10036 (N_10036,N_9788,N_9999);
xnor U10037 (N_10037,N_9527,N_9596);
xnor U10038 (N_10038,N_9911,N_9817);
nand U10039 (N_10039,N_9997,N_9851);
and U10040 (N_10040,N_9667,N_9678);
or U10041 (N_10041,N_9924,N_9759);
nand U10042 (N_10042,N_9572,N_9680);
and U10043 (N_10043,N_9737,N_9614);
and U10044 (N_10044,N_9553,N_9887);
nand U10045 (N_10045,N_9715,N_9886);
and U10046 (N_10046,N_9981,N_9856);
nor U10047 (N_10047,N_9674,N_9602);
nand U10048 (N_10048,N_9790,N_9854);
and U10049 (N_10049,N_9669,N_9926);
nor U10050 (N_10050,N_9507,N_9806);
and U10051 (N_10051,N_9824,N_9760);
nor U10052 (N_10052,N_9565,N_9885);
nor U10053 (N_10053,N_9736,N_9670);
and U10054 (N_10054,N_9989,N_9950);
or U10055 (N_10055,N_9583,N_9558);
xnor U10056 (N_10056,N_9765,N_9835);
nand U10057 (N_10057,N_9551,N_9791);
nor U10058 (N_10058,N_9639,N_9943);
or U10059 (N_10059,N_9991,N_9710);
nand U10060 (N_10060,N_9843,N_9958);
nor U10061 (N_10061,N_9616,N_9787);
and U10062 (N_10062,N_9682,N_9581);
and U10063 (N_10063,N_9706,N_9847);
nor U10064 (N_10064,N_9872,N_9778);
nand U10065 (N_10065,N_9719,N_9618);
xor U10066 (N_10066,N_9543,N_9730);
nor U10067 (N_10067,N_9709,N_9771);
nor U10068 (N_10068,N_9891,N_9819);
nor U10069 (N_10069,N_9769,N_9855);
and U10070 (N_10070,N_9953,N_9901);
nor U10071 (N_10071,N_9668,N_9799);
nand U10072 (N_10072,N_9571,N_9917);
nand U10073 (N_10073,N_9944,N_9727);
and U10074 (N_10074,N_9541,N_9998);
nand U10075 (N_10075,N_9585,N_9586);
or U10076 (N_10076,N_9839,N_9636);
or U10077 (N_10077,N_9812,N_9773);
and U10078 (N_10078,N_9776,N_9500);
or U10079 (N_10079,N_9582,N_9877);
and U10080 (N_10080,N_9818,N_9774);
xnor U10081 (N_10081,N_9875,N_9661);
nand U10082 (N_10082,N_9697,N_9936);
nand U10083 (N_10083,N_9672,N_9923);
nand U10084 (N_10084,N_9717,N_9804);
nor U10085 (N_10085,N_9990,N_9753);
nor U10086 (N_10086,N_9881,N_9664);
nand U10087 (N_10087,N_9988,N_9511);
and U10088 (N_10088,N_9679,N_9895);
nand U10089 (N_10089,N_9645,N_9928);
xnor U10090 (N_10090,N_9693,N_9677);
nand U10091 (N_10091,N_9756,N_9601);
nand U10092 (N_10092,N_9673,N_9642);
nand U10093 (N_10093,N_9702,N_9934);
nor U10094 (N_10094,N_9520,N_9977);
nor U10095 (N_10095,N_9970,N_9535);
or U10096 (N_10096,N_9694,N_9922);
nand U10097 (N_10097,N_9685,N_9834);
nor U10098 (N_10098,N_9782,N_9882);
nand U10099 (N_10099,N_9747,N_9621);
xor U10100 (N_10100,N_9505,N_9577);
xnor U10101 (N_10101,N_9801,N_9718);
xnor U10102 (N_10102,N_9735,N_9657);
xor U10103 (N_10103,N_9975,N_9893);
xor U10104 (N_10104,N_9913,N_9711);
or U10105 (N_10105,N_9532,N_9652);
nand U10106 (N_10106,N_9884,N_9828);
and U10107 (N_10107,N_9721,N_9775);
and U10108 (N_10108,N_9517,N_9896);
nand U10109 (N_10109,N_9620,N_9690);
nand U10110 (N_10110,N_9647,N_9826);
xor U10111 (N_10111,N_9880,N_9570);
xnor U10112 (N_10112,N_9608,N_9837);
or U10113 (N_10113,N_9940,N_9598);
and U10114 (N_10114,N_9524,N_9992);
and U10115 (N_10115,N_9800,N_9744);
nor U10116 (N_10116,N_9523,N_9897);
or U10117 (N_10117,N_9604,N_9611);
nor U10118 (N_10118,N_9874,N_9909);
or U10119 (N_10119,N_9930,N_9764);
nor U10120 (N_10120,N_9643,N_9584);
xnor U10121 (N_10121,N_9861,N_9831);
and U10122 (N_10122,N_9852,N_9894);
nor U10123 (N_10123,N_9613,N_9919);
nand U10124 (N_10124,N_9503,N_9510);
or U10125 (N_10125,N_9589,N_9741);
and U10126 (N_10126,N_9876,N_9986);
nor U10127 (N_10127,N_9842,N_9530);
or U10128 (N_10128,N_9547,N_9729);
and U10129 (N_10129,N_9785,N_9650);
or U10130 (N_10130,N_9575,N_9696);
nor U10131 (N_10131,N_9836,N_9956);
or U10132 (N_10132,N_9939,N_9786);
and U10133 (N_10133,N_9518,N_9907);
or U10134 (N_10134,N_9962,N_9949);
or U10135 (N_10135,N_9606,N_9688);
or U10136 (N_10136,N_9825,N_9629);
xnor U10137 (N_10137,N_9762,N_9529);
or U10138 (N_10138,N_9644,N_9937);
xor U10139 (N_10139,N_9830,N_9797);
or U10140 (N_10140,N_9566,N_9689);
xnor U10141 (N_10141,N_9569,N_9725);
nand U10142 (N_10142,N_9822,N_9903);
or U10143 (N_10143,N_9600,N_9591);
and U10144 (N_10144,N_9789,N_9686);
and U10145 (N_10145,N_9899,N_9592);
nor U10146 (N_10146,N_9627,N_9752);
nor U10147 (N_10147,N_9707,N_9795);
nand U10148 (N_10148,N_9810,N_9599);
xnor U10149 (N_10149,N_9948,N_9637);
and U10150 (N_10150,N_9648,N_9980);
nand U10151 (N_10151,N_9868,N_9829);
and U10152 (N_10152,N_9815,N_9528);
or U10153 (N_10153,N_9610,N_9883);
nor U10154 (N_10154,N_9683,N_9793);
xor U10155 (N_10155,N_9912,N_9982);
xor U10156 (N_10156,N_9513,N_9867);
or U10157 (N_10157,N_9749,N_9954);
or U10158 (N_10158,N_9951,N_9634);
nor U10159 (N_10159,N_9781,N_9857);
xnor U10160 (N_10160,N_9716,N_9701);
and U10161 (N_10161,N_9732,N_9537);
nand U10162 (N_10162,N_9573,N_9763);
nor U10163 (N_10163,N_9869,N_9724);
xor U10164 (N_10164,N_9864,N_9878);
or U10165 (N_10165,N_9814,N_9705);
and U10166 (N_10166,N_9879,N_9914);
nand U10167 (N_10167,N_9720,N_9658);
nor U10168 (N_10168,N_9996,N_9743);
nand U10169 (N_10169,N_9628,N_9574);
and U10170 (N_10170,N_9844,N_9651);
or U10171 (N_10171,N_9972,N_9561);
and U10172 (N_10172,N_9813,N_9904);
nor U10173 (N_10173,N_9873,N_9767);
xnor U10174 (N_10174,N_9742,N_9993);
xnor U10175 (N_10175,N_9784,N_9714);
and U10176 (N_10176,N_9798,N_9536);
or U10177 (N_10177,N_9519,N_9739);
nand U10178 (N_10178,N_9509,N_9671);
and U10179 (N_10179,N_9594,N_9971);
xor U10180 (N_10180,N_9516,N_9612);
or U10181 (N_10181,N_9920,N_9846);
nand U10182 (N_10182,N_9638,N_9712);
nor U10183 (N_10183,N_9973,N_9871);
nor U10184 (N_10184,N_9722,N_9966);
nand U10185 (N_10185,N_9654,N_9653);
nor U10186 (N_10186,N_9770,N_9560);
and U10187 (N_10187,N_9623,N_9695);
nor U10188 (N_10188,N_9563,N_9632);
xor U10189 (N_10189,N_9731,N_9802);
or U10190 (N_10190,N_9580,N_9918);
or U10191 (N_10191,N_9758,N_9579);
or U10192 (N_10192,N_9983,N_9985);
and U10193 (N_10193,N_9816,N_9957);
nand U10194 (N_10194,N_9624,N_9905);
xor U10195 (N_10195,N_9590,N_9995);
xnor U10196 (N_10196,N_9567,N_9663);
xnor U10197 (N_10197,N_9906,N_9723);
nor U10198 (N_10198,N_9755,N_9849);
xor U10199 (N_10199,N_9794,N_9994);
and U10200 (N_10200,N_9504,N_9902);
nor U10201 (N_10201,N_9915,N_9728);
or U10202 (N_10202,N_9666,N_9641);
xnor U10203 (N_10203,N_9840,N_9587);
and U10204 (N_10204,N_9766,N_9687);
xnor U10205 (N_10205,N_9538,N_9821);
xnor U10206 (N_10206,N_9910,N_9617);
nor U10207 (N_10207,N_9514,N_9889);
nor U10208 (N_10208,N_9700,N_9738);
and U10209 (N_10209,N_9968,N_9941);
nor U10210 (N_10210,N_9865,N_9681);
nor U10211 (N_10211,N_9833,N_9626);
nor U10212 (N_10212,N_9978,N_9740);
nand U10213 (N_10213,N_9768,N_9858);
nor U10214 (N_10214,N_9607,N_9615);
or U10215 (N_10215,N_9605,N_9646);
nor U10216 (N_10216,N_9703,N_9967);
or U10217 (N_10217,N_9534,N_9549);
xnor U10218 (N_10218,N_9544,N_9631);
nor U10219 (N_10219,N_9748,N_9761);
nand U10220 (N_10220,N_9823,N_9932);
xor U10221 (N_10221,N_9515,N_9502);
or U10222 (N_10222,N_9562,N_9965);
and U10223 (N_10223,N_9635,N_9931);
or U10224 (N_10224,N_9684,N_9593);
and U10225 (N_10225,N_9704,N_9892);
xor U10226 (N_10226,N_9576,N_9832);
and U10227 (N_10227,N_9805,N_9845);
nor U10228 (N_10228,N_9859,N_9675);
nand U10229 (N_10229,N_9807,N_9935);
and U10230 (N_10230,N_9809,N_9925);
and U10231 (N_10231,N_9908,N_9633);
or U10232 (N_10232,N_9539,N_9921);
nand U10233 (N_10233,N_9890,N_9659);
and U10234 (N_10234,N_9542,N_9506);
xnor U10235 (N_10235,N_9808,N_9783);
xnor U10236 (N_10236,N_9555,N_9976);
nor U10237 (N_10237,N_9691,N_9945);
xnor U10238 (N_10238,N_9512,N_9863);
or U10239 (N_10239,N_9916,N_9838);
nor U10240 (N_10240,N_9521,N_9974);
nor U10241 (N_10241,N_9622,N_9559);
xor U10242 (N_10242,N_9792,N_9548);
and U10243 (N_10243,N_9929,N_9713);
nor U10244 (N_10244,N_9665,N_9501);
or U10245 (N_10245,N_9938,N_9960);
nand U10246 (N_10246,N_9959,N_9531);
xor U10247 (N_10247,N_9540,N_9625);
and U10248 (N_10248,N_9619,N_9588);
and U10249 (N_10249,N_9820,N_9772);
nand U10250 (N_10250,N_9621,N_9946);
and U10251 (N_10251,N_9741,N_9531);
nand U10252 (N_10252,N_9543,N_9723);
and U10253 (N_10253,N_9523,N_9917);
nand U10254 (N_10254,N_9623,N_9864);
or U10255 (N_10255,N_9912,N_9746);
or U10256 (N_10256,N_9632,N_9584);
xnor U10257 (N_10257,N_9504,N_9534);
nand U10258 (N_10258,N_9967,N_9996);
and U10259 (N_10259,N_9783,N_9726);
xnor U10260 (N_10260,N_9762,N_9530);
and U10261 (N_10261,N_9988,N_9713);
xor U10262 (N_10262,N_9807,N_9701);
nor U10263 (N_10263,N_9700,N_9827);
and U10264 (N_10264,N_9909,N_9628);
nor U10265 (N_10265,N_9632,N_9944);
or U10266 (N_10266,N_9662,N_9558);
nand U10267 (N_10267,N_9658,N_9982);
nand U10268 (N_10268,N_9818,N_9931);
xor U10269 (N_10269,N_9916,N_9688);
and U10270 (N_10270,N_9941,N_9828);
nand U10271 (N_10271,N_9980,N_9721);
xor U10272 (N_10272,N_9571,N_9819);
nand U10273 (N_10273,N_9905,N_9874);
nand U10274 (N_10274,N_9692,N_9953);
nand U10275 (N_10275,N_9952,N_9656);
nor U10276 (N_10276,N_9675,N_9960);
xnor U10277 (N_10277,N_9693,N_9938);
xnor U10278 (N_10278,N_9571,N_9716);
nand U10279 (N_10279,N_9618,N_9657);
xor U10280 (N_10280,N_9870,N_9535);
and U10281 (N_10281,N_9567,N_9862);
and U10282 (N_10282,N_9741,N_9679);
or U10283 (N_10283,N_9549,N_9636);
or U10284 (N_10284,N_9589,N_9762);
and U10285 (N_10285,N_9726,N_9904);
nand U10286 (N_10286,N_9653,N_9673);
nand U10287 (N_10287,N_9795,N_9658);
and U10288 (N_10288,N_9614,N_9937);
nand U10289 (N_10289,N_9828,N_9979);
nor U10290 (N_10290,N_9577,N_9918);
nor U10291 (N_10291,N_9802,N_9916);
nand U10292 (N_10292,N_9962,N_9570);
or U10293 (N_10293,N_9594,N_9703);
nor U10294 (N_10294,N_9814,N_9779);
or U10295 (N_10295,N_9776,N_9751);
and U10296 (N_10296,N_9622,N_9834);
or U10297 (N_10297,N_9903,N_9680);
and U10298 (N_10298,N_9930,N_9982);
nor U10299 (N_10299,N_9533,N_9972);
or U10300 (N_10300,N_9786,N_9691);
nand U10301 (N_10301,N_9563,N_9908);
nor U10302 (N_10302,N_9890,N_9671);
nor U10303 (N_10303,N_9758,N_9968);
nand U10304 (N_10304,N_9746,N_9909);
xnor U10305 (N_10305,N_9808,N_9777);
nand U10306 (N_10306,N_9954,N_9871);
nor U10307 (N_10307,N_9642,N_9790);
xor U10308 (N_10308,N_9736,N_9852);
nand U10309 (N_10309,N_9633,N_9610);
and U10310 (N_10310,N_9673,N_9948);
nand U10311 (N_10311,N_9558,N_9507);
nand U10312 (N_10312,N_9843,N_9897);
nand U10313 (N_10313,N_9516,N_9712);
xor U10314 (N_10314,N_9660,N_9986);
and U10315 (N_10315,N_9929,N_9588);
or U10316 (N_10316,N_9608,N_9929);
or U10317 (N_10317,N_9788,N_9852);
xnor U10318 (N_10318,N_9954,N_9735);
xnor U10319 (N_10319,N_9986,N_9812);
xor U10320 (N_10320,N_9820,N_9871);
and U10321 (N_10321,N_9788,N_9699);
nand U10322 (N_10322,N_9998,N_9858);
or U10323 (N_10323,N_9835,N_9592);
nor U10324 (N_10324,N_9798,N_9775);
nor U10325 (N_10325,N_9864,N_9819);
nand U10326 (N_10326,N_9770,N_9950);
and U10327 (N_10327,N_9700,N_9532);
nand U10328 (N_10328,N_9855,N_9529);
xor U10329 (N_10329,N_9667,N_9608);
xor U10330 (N_10330,N_9946,N_9908);
and U10331 (N_10331,N_9582,N_9743);
nor U10332 (N_10332,N_9635,N_9917);
or U10333 (N_10333,N_9868,N_9591);
nand U10334 (N_10334,N_9723,N_9975);
xnor U10335 (N_10335,N_9795,N_9876);
nor U10336 (N_10336,N_9592,N_9629);
or U10337 (N_10337,N_9554,N_9763);
nand U10338 (N_10338,N_9581,N_9968);
and U10339 (N_10339,N_9995,N_9919);
and U10340 (N_10340,N_9823,N_9627);
nor U10341 (N_10341,N_9814,N_9880);
nor U10342 (N_10342,N_9684,N_9630);
nor U10343 (N_10343,N_9836,N_9708);
or U10344 (N_10344,N_9773,N_9850);
or U10345 (N_10345,N_9892,N_9850);
xor U10346 (N_10346,N_9699,N_9884);
nand U10347 (N_10347,N_9743,N_9543);
xor U10348 (N_10348,N_9729,N_9834);
nand U10349 (N_10349,N_9516,N_9617);
or U10350 (N_10350,N_9591,N_9746);
nor U10351 (N_10351,N_9573,N_9839);
and U10352 (N_10352,N_9669,N_9591);
xnor U10353 (N_10353,N_9998,N_9936);
nand U10354 (N_10354,N_9828,N_9573);
or U10355 (N_10355,N_9707,N_9643);
xnor U10356 (N_10356,N_9652,N_9614);
nor U10357 (N_10357,N_9797,N_9779);
or U10358 (N_10358,N_9965,N_9898);
or U10359 (N_10359,N_9855,N_9830);
xor U10360 (N_10360,N_9920,N_9791);
or U10361 (N_10361,N_9868,N_9978);
or U10362 (N_10362,N_9676,N_9877);
or U10363 (N_10363,N_9606,N_9580);
nor U10364 (N_10364,N_9900,N_9568);
xnor U10365 (N_10365,N_9718,N_9748);
or U10366 (N_10366,N_9618,N_9843);
and U10367 (N_10367,N_9515,N_9854);
or U10368 (N_10368,N_9877,N_9816);
and U10369 (N_10369,N_9507,N_9514);
nand U10370 (N_10370,N_9526,N_9592);
nand U10371 (N_10371,N_9801,N_9535);
or U10372 (N_10372,N_9634,N_9826);
nor U10373 (N_10373,N_9895,N_9941);
or U10374 (N_10374,N_9582,N_9869);
nor U10375 (N_10375,N_9874,N_9846);
nor U10376 (N_10376,N_9778,N_9638);
or U10377 (N_10377,N_9575,N_9501);
nand U10378 (N_10378,N_9954,N_9860);
or U10379 (N_10379,N_9971,N_9903);
or U10380 (N_10380,N_9828,N_9660);
and U10381 (N_10381,N_9659,N_9528);
or U10382 (N_10382,N_9755,N_9797);
and U10383 (N_10383,N_9553,N_9763);
or U10384 (N_10384,N_9616,N_9594);
or U10385 (N_10385,N_9594,N_9940);
and U10386 (N_10386,N_9739,N_9703);
nand U10387 (N_10387,N_9553,N_9933);
xnor U10388 (N_10388,N_9749,N_9717);
and U10389 (N_10389,N_9784,N_9605);
or U10390 (N_10390,N_9647,N_9941);
xor U10391 (N_10391,N_9614,N_9747);
nor U10392 (N_10392,N_9667,N_9769);
and U10393 (N_10393,N_9813,N_9643);
nand U10394 (N_10394,N_9935,N_9665);
or U10395 (N_10395,N_9957,N_9857);
and U10396 (N_10396,N_9519,N_9590);
nand U10397 (N_10397,N_9567,N_9925);
and U10398 (N_10398,N_9543,N_9979);
nor U10399 (N_10399,N_9867,N_9799);
and U10400 (N_10400,N_9790,N_9910);
xnor U10401 (N_10401,N_9801,N_9626);
nor U10402 (N_10402,N_9589,N_9914);
xnor U10403 (N_10403,N_9881,N_9865);
nor U10404 (N_10404,N_9672,N_9640);
xnor U10405 (N_10405,N_9679,N_9722);
nor U10406 (N_10406,N_9774,N_9655);
xor U10407 (N_10407,N_9565,N_9580);
nor U10408 (N_10408,N_9645,N_9865);
nor U10409 (N_10409,N_9973,N_9710);
nor U10410 (N_10410,N_9724,N_9893);
or U10411 (N_10411,N_9534,N_9521);
and U10412 (N_10412,N_9938,N_9626);
or U10413 (N_10413,N_9524,N_9851);
xor U10414 (N_10414,N_9808,N_9963);
and U10415 (N_10415,N_9698,N_9507);
or U10416 (N_10416,N_9761,N_9654);
and U10417 (N_10417,N_9990,N_9946);
or U10418 (N_10418,N_9780,N_9648);
nor U10419 (N_10419,N_9899,N_9963);
and U10420 (N_10420,N_9624,N_9760);
nor U10421 (N_10421,N_9981,N_9615);
xnor U10422 (N_10422,N_9811,N_9623);
nand U10423 (N_10423,N_9989,N_9739);
nor U10424 (N_10424,N_9660,N_9708);
or U10425 (N_10425,N_9857,N_9994);
or U10426 (N_10426,N_9697,N_9869);
xor U10427 (N_10427,N_9544,N_9508);
xnor U10428 (N_10428,N_9899,N_9529);
nor U10429 (N_10429,N_9702,N_9896);
nand U10430 (N_10430,N_9500,N_9556);
or U10431 (N_10431,N_9750,N_9762);
xnor U10432 (N_10432,N_9996,N_9649);
xnor U10433 (N_10433,N_9749,N_9626);
xnor U10434 (N_10434,N_9727,N_9800);
nand U10435 (N_10435,N_9590,N_9664);
xor U10436 (N_10436,N_9579,N_9589);
nand U10437 (N_10437,N_9733,N_9642);
and U10438 (N_10438,N_9526,N_9788);
or U10439 (N_10439,N_9823,N_9925);
or U10440 (N_10440,N_9974,N_9599);
and U10441 (N_10441,N_9530,N_9564);
nor U10442 (N_10442,N_9903,N_9884);
or U10443 (N_10443,N_9733,N_9990);
nor U10444 (N_10444,N_9833,N_9877);
nand U10445 (N_10445,N_9673,N_9988);
xor U10446 (N_10446,N_9599,N_9840);
xor U10447 (N_10447,N_9813,N_9744);
nor U10448 (N_10448,N_9759,N_9595);
nand U10449 (N_10449,N_9810,N_9604);
and U10450 (N_10450,N_9938,N_9595);
nor U10451 (N_10451,N_9694,N_9510);
xor U10452 (N_10452,N_9614,N_9959);
nor U10453 (N_10453,N_9535,N_9966);
xnor U10454 (N_10454,N_9533,N_9636);
and U10455 (N_10455,N_9998,N_9775);
or U10456 (N_10456,N_9707,N_9548);
or U10457 (N_10457,N_9896,N_9741);
and U10458 (N_10458,N_9528,N_9934);
nand U10459 (N_10459,N_9764,N_9722);
nor U10460 (N_10460,N_9757,N_9687);
or U10461 (N_10461,N_9708,N_9875);
and U10462 (N_10462,N_9974,N_9847);
nand U10463 (N_10463,N_9987,N_9746);
and U10464 (N_10464,N_9891,N_9534);
nor U10465 (N_10465,N_9951,N_9814);
nor U10466 (N_10466,N_9954,N_9501);
xor U10467 (N_10467,N_9520,N_9923);
xor U10468 (N_10468,N_9854,N_9713);
nor U10469 (N_10469,N_9507,N_9741);
nor U10470 (N_10470,N_9781,N_9865);
and U10471 (N_10471,N_9724,N_9514);
and U10472 (N_10472,N_9553,N_9669);
nand U10473 (N_10473,N_9667,N_9554);
nand U10474 (N_10474,N_9984,N_9930);
xor U10475 (N_10475,N_9859,N_9805);
nand U10476 (N_10476,N_9862,N_9985);
nand U10477 (N_10477,N_9716,N_9549);
xor U10478 (N_10478,N_9790,N_9784);
nand U10479 (N_10479,N_9543,N_9919);
nor U10480 (N_10480,N_9613,N_9608);
xnor U10481 (N_10481,N_9990,N_9672);
or U10482 (N_10482,N_9603,N_9774);
nand U10483 (N_10483,N_9815,N_9665);
nor U10484 (N_10484,N_9741,N_9686);
and U10485 (N_10485,N_9508,N_9721);
or U10486 (N_10486,N_9536,N_9811);
xnor U10487 (N_10487,N_9556,N_9591);
xnor U10488 (N_10488,N_9966,N_9899);
nor U10489 (N_10489,N_9730,N_9731);
or U10490 (N_10490,N_9849,N_9723);
xor U10491 (N_10491,N_9535,N_9905);
xnor U10492 (N_10492,N_9639,N_9959);
or U10493 (N_10493,N_9588,N_9982);
nand U10494 (N_10494,N_9730,N_9973);
xnor U10495 (N_10495,N_9924,N_9653);
xnor U10496 (N_10496,N_9551,N_9748);
xnor U10497 (N_10497,N_9616,N_9967);
nand U10498 (N_10498,N_9577,N_9673);
and U10499 (N_10499,N_9656,N_9568);
or U10500 (N_10500,N_10357,N_10119);
or U10501 (N_10501,N_10011,N_10281);
or U10502 (N_10502,N_10380,N_10309);
or U10503 (N_10503,N_10110,N_10160);
xor U10504 (N_10504,N_10266,N_10081);
nand U10505 (N_10505,N_10220,N_10353);
xnor U10506 (N_10506,N_10225,N_10331);
nor U10507 (N_10507,N_10026,N_10214);
nor U10508 (N_10508,N_10325,N_10207);
xor U10509 (N_10509,N_10072,N_10361);
xor U10510 (N_10510,N_10149,N_10175);
nand U10511 (N_10511,N_10445,N_10365);
nand U10512 (N_10512,N_10157,N_10394);
xor U10513 (N_10513,N_10434,N_10198);
and U10514 (N_10514,N_10320,N_10035);
or U10515 (N_10515,N_10354,N_10262);
or U10516 (N_10516,N_10019,N_10479);
nor U10517 (N_10517,N_10340,N_10187);
and U10518 (N_10518,N_10240,N_10383);
and U10519 (N_10519,N_10116,N_10381);
nor U10520 (N_10520,N_10437,N_10471);
nor U10521 (N_10521,N_10265,N_10291);
xor U10522 (N_10522,N_10447,N_10177);
and U10523 (N_10523,N_10459,N_10310);
or U10524 (N_10524,N_10270,N_10084);
nor U10525 (N_10525,N_10382,N_10347);
nand U10526 (N_10526,N_10128,N_10139);
xnor U10527 (N_10527,N_10478,N_10252);
nand U10528 (N_10528,N_10043,N_10000);
nor U10529 (N_10529,N_10045,N_10206);
nand U10530 (N_10530,N_10080,N_10356);
nor U10531 (N_10531,N_10030,N_10023);
xnor U10532 (N_10532,N_10086,N_10449);
nand U10533 (N_10533,N_10453,N_10372);
nand U10534 (N_10534,N_10341,N_10302);
or U10535 (N_10535,N_10203,N_10275);
and U10536 (N_10536,N_10074,N_10188);
nor U10537 (N_10537,N_10362,N_10371);
xnor U10538 (N_10538,N_10264,N_10488);
xor U10539 (N_10539,N_10260,N_10429);
nor U10540 (N_10540,N_10158,N_10247);
or U10541 (N_10541,N_10232,N_10244);
nand U10542 (N_10542,N_10306,N_10497);
or U10543 (N_10543,N_10173,N_10319);
and U10544 (N_10544,N_10435,N_10192);
and U10545 (N_10545,N_10444,N_10197);
nor U10546 (N_10546,N_10234,N_10415);
and U10547 (N_10547,N_10165,N_10100);
nor U10548 (N_10548,N_10104,N_10055);
nor U10549 (N_10549,N_10031,N_10483);
or U10550 (N_10550,N_10250,N_10370);
xnor U10551 (N_10551,N_10156,N_10374);
xor U10552 (N_10552,N_10287,N_10088);
and U10553 (N_10553,N_10153,N_10059);
or U10554 (N_10554,N_10326,N_10178);
and U10555 (N_10555,N_10248,N_10062);
nand U10556 (N_10556,N_10421,N_10082);
nand U10557 (N_10557,N_10258,N_10036);
nand U10558 (N_10558,N_10295,N_10231);
nor U10559 (N_10559,N_10193,N_10352);
nand U10560 (N_10560,N_10123,N_10179);
xor U10561 (N_10561,N_10235,N_10399);
nand U10562 (N_10562,N_10056,N_10077);
xor U10563 (N_10563,N_10360,N_10268);
nor U10564 (N_10564,N_10273,N_10135);
and U10565 (N_10565,N_10004,N_10422);
nor U10566 (N_10566,N_10425,N_10303);
nor U10567 (N_10567,N_10242,N_10095);
and U10568 (N_10568,N_10057,N_10442);
or U10569 (N_10569,N_10229,N_10141);
nor U10570 (N_10570,N_10473,N_10493);
nand U10571 (N_10571,N_10430,N_10440);
nor U10572 (N_10572,N_10277,N_10106);
nand U10573 (N_10573,N_10046,N_10344);
xnor U10574 (N_10574,N_10317,N_10377);
xor U10575 (N_10575,N_10448,N_10330);
xnor U10576 (N_10576,N_10152,N_10499);
nor U10577 (N_10577,N_10194,N_10114);
or U10578 (N_10578,N_10245,N_10008);
nor U10579 (N_10579,N_10130,N_10020);
and U10580 (N_10580,N_10241,N_10358);
or U10581 (N_10581,N_10454,N_10054);
and U10582 (N_10582,N_10391,N_10064);
nand U10583 (N_10583,N_10301,N_10164);
nand U10584 (N_10584,N_10099,N_10034);
xor U10585 (N_10585,N_10047,N_10070);
or U10586 (N_10586,N_10147,N_10218);
or U10587 (N_10587,N_10006,N_10029);
or U10588 (N_10588,N_10462,N_10044);
and U10589 (N_10589,N_10009,N_10439);
nor U10590 (N_10590,N_10261,N_10233);
nor U10591 (N_10591,N_10313,N_10217);
or U10592 (N_10592,N_10386,N_10398);
or U10593 (N_10593,N_10419,N_10176);
nand U10594 (N_10594,N_10061,N_10170);
xor U10595 (N_10595,N_10468,N_10426);
and U10596 (N_10596,N_10083,N_10005);
or U10597 (N_10597,N_10406,N_10254);
or U10598 (N_10598,N_10085,N_10427);
or U10599 (N_10599,N_10089,N_10167);
or U10600 (N_10600,N_10292,N_10068);
nand U10601 (N_10601,N_10451,N_10414);
xnor U10602 (N_10602,N_10113,N_10073);
and U10603 (N_10603,N_10120,N_10308);
nand U10604 (N_10604,N_10392,N_10485);
and U10605 (N_10605,N_10443,N_10115);
or U10606 (N_10606,N_10002,N_10393);
xor U10607 (N_10607,N_10202,N_10282);
nor U10608 (N_10608,N_10286,N_10490);
nand U10609 (N_10609,N_10132,N_10498);
nor U10610 (N_10610,N_10159,N_10289);
and U10611 (N_10611,N_10373,N_10311);
xnor U10612 (N_10612,N_10142,N_10298);
or U10613 (N_10613,N_10108,N_10090);
or U10614 (N_10614,N_10405,N_10109);
nand U10615 (N_10615,N_10010,N_10375);
or U10616 (N_10616,N_10408,N_10169);
and U10617 (N_10617,N_10323,N_10180);
nand U10618 (N_10618,N_10376,N_10183);
nor U10619 (N_10619,N_10293,N_10125);
xnor U10620 (N_10620,N_10017,N_10369);
and U10621 (N_10621,N_10060,N_10338);
and U10622 (N_10622,N_10257,N_10350);
or U10623 (N_10623,N_10208,N_10144);
or U10624 (N_10624,N_10336,N_10328);
nor U10625 (N_10625,N_10464,N_10129);
or U10626 (N_10626,N_10256,N_10117);
nand U10627 (N_10627,N_10487,N_10413);
nor U10628 (N_10628,N_10297,N_10342);
xor U10629 (N_10629,N_10280,N_10140);
xor U10630 (N_10630,N_10318,N_10307);
and U10631 (N_10631,N_10461,N_10452);
xor U10632 (N_10632,N_10050,N_10096);
and U10633 (N_10633,N_10122,N_10436);
nor U10634 (N_10634,N_10200,N_10463);
nor U10635 (N_10635,N_10033,N_10480);
nand U10636 (N_10636,N_10314,N_10492);
and U10637 (N_10637,N_10205,N_10076);
nand U10638 (N_10638,N_10053,N_10251);
nand U10639 (N_10639,N_10211,N_10032);
and U10640 (N_10640,N_10423,N_10092);
nand U10641 (N_10641,N_10022,N_10335);
or U10642 (N_10642,N_10316,N_10355);
nor U10643 (N_10643,N_10458,N_10486);
nand U10644 (N_10644,N_10037,N_10172);
and U10645 (N_10645,N_10025,N_10038);
and U10646 (N_10646,N_10121,N_10191);
nor U10647 (N_10647,N_10212,N_10027);
nor U10648 (N_10648,N_10329,N_10238);
xor U10649 (N_10649,N_10091,N_10438);
xor U10650 (N_10650,N_10366,N_10168);
xor U10651 (N_10651,N_10278,N_10284);
nor U10652 (N_10652,N_10014,N_10446);
nand U10653 (N_10653,N_10013,N_10040);
or U10654 (N_10654,N_10322,N_10321);
or U10655 (N_10655,N_10327,N_10339);
nand U10656 (N_10656,N_10384,N_10418);
and U10657 (N_10657,N_10223,N_10146);
xnor U10658 (N_10658,N_10174,N_10412);
xnor U10659 (N_10659,N_10288,N_10184);
xnor U10660 (N_10660,N_10199,N_10195);
or U10661 (N_10661,N_10093,N_10118);
or U10662 (N_10662,N_10407,N_10102);
nand U10663 (N_10663,N_10111,N_10171);
or U10664 (N_10664,N_10315,N_10150);
and U10665 (N_10665,N_10397,N_10101);
or U10666 (N_10666,N_10182,N_10334);
nand U10667 (N_10667,N_10465,N_10267);
xor U10668 (N_10668,N_10283,N_10378);
nor U10669 (N_10669,N_10222,N_10400);
xor U10670 (N_10670,N_10276,N_10379);
and U10671 (N_10671,N_10039,N_10484);
or U10672 (N_10672,N_10279,N_10410);
or U10673 (N_10673,N_10098,N_10127);
or U10674 (N_10674,N_10489,N_10126);
xor U10675 (N_10675,N_10403,N_10409);
or U10676 (N_10676,N_10363,N_10432);
xor U10677 (N_10677,N_10243,N_10151);
and U10678 (N_10678,N_10482,N_10263);
and U10679 (N_10679,N_10143,N_10476);
nor U10680 (N_10680,N_10299,N_10097);
and U10681 (N_10681,N_10467,N_10390);
nand U10682 (N_10682,N_10087,N_10071);
xnor U10683 (N_10683,N_10215,N_10349);
and U10684 (N_10684,N_10431,N_10145);
and U10685 (N_10685,N_10201,N_10332);
nand U10686 (N_10686,N_10124,N_10290);
nand U10687 (N_10687,N_10051,N_10166);
xor U10688 (N_10688,N_10253,N_10162);
and U10689 (N_10689,N_10402,N_10204);
xnor U10690 (N_10690,N_10420,N_10337);
and U10691 (N_10691,N_10491,N_10227);
or U10692 (N_10692,N_10213,N_10189);
and U10693 (N_10693,N_10312,N_10075);
and U10694 (N_10694,N_10456,N_10016);
or U10695 (N_10695,N_10343,N_10368);
nand U10696 (N_10696,N_10079,N_10417);
nand U10697 (N_10697,N_10012,N_10163);
and U10698 (N_10698,N_10470,N_10359);
nand U10699 (N_10699,N_10224,N_10494);
nand U10700 (N_10700,N_10185,N_10001);
nand U10701 (N_10701,N_10450,N_10161);
and U10702 (N_10702,N_10351,N_10155);
xnor U10703 (N_10703,N_10069,N_10333);
xnor U10704 (N_10704,N_10255,N_10455);
nand U10705 (N_10705,N_10133,N_10274);
or U10706 (N_10706,N_10018,N_10210);
nor U10707 (N_10707,N_10388,N_10024);
nor U10708 (N_10708,N_10294,N_10041);
nand U10709 (N_10709,N_10495,N_10007);
xor U10710 (N_10710,N_10181,N_10042);
or U10711 (N_10711,N_10209,N_10411);
or U10712 (N_10712,N_10472,N_10496);
xor U10713 (N_10713,N_10131,N_10385);
nor U10714 (N_10714,N_10346,N_10416);
or U10715 (N_10715,N_10249,N_10105);
nor U10716 (N_10716,N_10103,N_10048);
nor U10717 (N_10717,N_10481,N_10052);
or U10718 (N_10718,N_10230,N_10154);
and U10719 (N_10719,N_10457,N_10441);
xnor U10720 (N_10720,N_10049,N_10387);
and U10721 (N_10721,N_10067,N_10389);
nand U10722 (N_10722,N_10186,N_10028);
xor U10723 (N_10723,N_10134,N_10460);
and U10724 (N_10724,N_10364,N_10469);
or U10725 (N_10725,N_10401,N_10239);
nor U10726 (N_10726,N_10246,N_10021);
nand U10727 (N_10727,N_10065,N_10428);
nand U10728 (N_10728,N_10433,N_10474);
xor U10729 (N_10729,N_10424,N_10367);
nor U10730 (N_10730,N_10226,N_10078);
and U10731 (N_10731,N_10272,N_10148);
nor U10732 (N_10732,N_10107,N_10345);
nand U10733 (N_10733,N_10305,N_10466);
nand U10734 (N_10734,N_10015,N_10404);
and U10735 (N_10735,N_10136,N_10196);
nand U10736 (N_10736,N_10237,N_10300);
xor U10737 (N_10737,N_10396,N_10348);
nand U10738 (N_10738,N_10271,N_10236);
and U10739 (N_10739,N_10094,N_10285);
nand U10740 (N_10740,N_10003,N_10324);
and U10741 (N_10741,N_10477,N_10296);
or U10742 (N_10742,N_10138,N_10219);
nor U10743 (N_10743,N_10221,N_10228);
or U10744 (N_10744,N_10137,N_10395);
nor U10745 (N_10745,N_10269,N_10475);
or U10746 (N_10746,N_10216,N_10190);
or U10747 (N_10747,N_10063,N_10058);
and U10748 (N_10748,N_10066,N_10259);
or U10749 (N_10749,N_10304,N_10112);
and U10750 (N_10750,N_10136,N_10042);
nand U10751 (N_10751,N_10143,N_10192);
nor U10752 (N_10752,N_10104,N_10335);
nor U10753 (N_10753,N_10124,N_10111);
and U10754 (N_10754,N_10362,N_10218);
nand U10755 (N_10755,N_10411,N_10287);
and U10756 (N_10756,N_10101,N_10399);
nand U10757 (N_10757,N_10131,N_10064);
nor U10758 (N_10758,N_10336,N_10030);
or U10759 (N_10759,N_10402,N_10164);
nor U10760 (N_10760,N_10316,N_10331);
nor U10761 (N_10761,N_10301,N_10046);
nand U10762 (N_10762,N_10343,N_10413);
xor U10763 (N_10763,N_10288,N_10213);
or U10764 (N_10764,N_10175,N_10449);
nor U10765 (N_10765,N_10379,N_10203);
nor U10766 (N_10766,N_10105,N_10397);
nor U10767 (N_10767,N_10392,N_10491);
xor U10768 (N_10768,N_10134,N_10278);
or U10769 (N_10769,N_10288,N_10209);
or U10770 (N_10770,N_10283,N_10165);
nand U10771 (N_10771,N_10077,N_10033);
nand U10772 (N_10772,N_10470,N_10467);
or U10773 (N_10773,N_10495,N_10289);
and U10774 (N_10774,N_10035,N_10478);
and U10775 (N_10775,N_10144,N_10303);
or U10776 (N_10776,N_10177,N_10186);
nor U10777 (N_10777,N_10339,N_10396);
xor U10778 (N_10778,N_10252,N_10444);
nand U10779 (N_10779,N_10104,N_10475);
xor U10780 (N_10780,N_10193,N_10134);
xor U10781 (N_10781,N_10472,N_10226);
nand U10782 (N_10782,N_10385,N_10313);
or U10783 (N_10783,N_10287,N_10093);
and U10784 (N_10784,N_10159,N_10004);
nand U10785 (N_10785,N_10497,N_10163);
and U10786 (N_10786,N_10316,N_10200);
nor U10787 (N_10787,N_10243,N_10326);
nor U10788 (N_10788,N_10153,N_10184);
nand U10789 (N_10789,N_10377,N_10296);
or U10790 (N_10790,N_10184,N_10362);
nor U10791 (N_10791,N_10228,N_10105);
xor U10792 (N_10792,N_10211,N_10346);
nand U10793 (N_10793,N_10247,N_10356);
nor U10794 (N_10794,N_10464,N_10073);
nand U10795 (N_10795,N_10289,N_10442);
nor U10796 (N_10796,N_10141,N_10496);
nor U10797 (N_10797,N_10433,N_10307);
or U10798 (N_10798,N_10307,N_10406);
nand U10799 (N_10799,N_10397,N_10498);
xor U10800 (N_10800,N_10374,N_10338);
nor U10801 (N_10801,N_10109,N_10043);
xnor U10802 (N_10802,N_10044,N_10006);
nor U10803 (N_10803,N_10303,N_10406);
nand U10804 (N_10804,N_10086,N_10128);
xor U10805 (N_10805,N_10372,N_10051);
and U10806 (N_10806,N_10341,N_10391);
or U10807 (N_10807,N_10167,N_10347);
and U10808 (N_10808,N_10459,N_10400);
nand U10809 (N_10809,N_10139,N_10218);
nand U10810 (N_10810,N_10234,N_10345);
nor U10811 (N_10811,N_10453,N_10480);
nand U10812 (N_10812,N_10325,N_10244);
nand U10813 (N_10813,N_10182,N_10131);
nor U10814 (N_10814,N_10135,N_10262);
nor U10815 (N_10815,N_10198,N_10328);
xor U10816 (N_10816,N_10164,N_10273);
xnor U10817 (N_10817,N_10171,N_10250);
nand U10818 (N_10818,N_10457,N_10069);
nor U10819 (N_10819,N_10440,N_10208);
xnor U10820 (N_10820,N_10358,N_10286);
nor U10821 (N_10821,N_10270,N_10255);
and U10822 (N_10822,N_10263,N_10304);
and U10823 (N_10823,N_10172,N_10148);
nor U10824 (N_10824,N_10061,N_10182);
xor U10825 (N_10825,N_10135,N_10220);
or U10826 (N_10826,N_10062,N_10030);
or U10827 (N_10827,N_10457,N_10237);
or U10828 (N_10828,N_10459,N_10282);
nand U10829 (N_10829,N_10049,N_10170);
nand U10830 (N_10830,N_10372,N_10127);
and U10831 (N_10831,N_10052,N_10145);
or U10832 (N_10832,N_10325,N_10021);
xor U10833 (N_10833,N_10447,N_10498);
and U10834 (N_10834,N_10283,N_10403);
nor U10835 (N_10835,N_10371,N_10135);
xnor U10836 (N_10836,N_10476,N_10372);
nand U10837 (N_10837,N_10200,N_10230);
nor U10838 (N_10838,N_10242,N_10353);
nor U10839 (N_10839,N_10133,N_10301);
or U10840 (N_10840,N_10481,N_10201);
nor U10841 (N_10841,N_10412,N_10165);
nor U10842 (N_10842,N_10406,N_10383);
nand U10843 (N_10843,N_10413,N_10476);
and U10844 (N_10844,N_10054,N_10378);
xnor U10845 (N_10845,N_10046,N_10169);
nand U10846 (N_10846,N_10482,N_10198);
xor U10847 (N_10847,N_10024,N_10312);
nor U10848 (N_10848,N_10483,N_10195);
nor U10849 (N_10849,N_10406,N_10455);
and U10850 (N_10850,N_10113,N_10448);
nand U10851 (N_10851,N_10047,N_10459);
or U10852 (N_10852,N_10305,N_10388);
nor U10853 (N_10853,N_10429,N_10201);
or U10854 (N_10854,N_10399,N_10473);
and U10855 (N_10855,N_10446,N_10317);
and U10856 (N_10856,N_10151,N_10075);
xnor U10857 (N_10857,N_10170,N_10213);
and U10858 (N_10858,N_10027,N_10400);
nor U10859 (N_10859,N_10311,N_10128);
xnor U10860 (N_10860,N_10211,N_10207);
nor U10861 (N_10861,N_10171,N_10097);
xnor U10862 (N_10862,N_10171,N_10068);
and U10863 (N_10863,N_10122,N_10263);
xor U10864 (N_10864,N_10296,N_10247);
nand U10865 (N_10865,N_10467,N_10462);
nand U10866 (N_10866,N_10486,N_10330);
and U10867 (N_10867,N_10170,N_10321);
or U10868 (N_10868,N_10204,N_10113);
and U10869 (N_10869,N_10430,N_10086);
xor U10870 (N_10870,N_10398,N_10151);
nand U10871 (N_10871,N_10045,N_10400);
or U10872 (N_10872,N_10338,N_10475);
or U10873 (N_10873,N_10204,N_10189);
xnor U10874 (N_10874,N_10484,N_10168);
xnor U10875 (N_10875,N_10473,N_10477);
nand U10876 (N_10876,N_10413,N_10341);
nor U10877 (N_10877,N_10436,N_10481);
nor U10878 (N_10878,N_10285,N_10200);
xnor U10879 (N_10879,N_10424,N_10072);
and U10880 (N_10880,N_10060,N_10477);
nor U10881 (N_10881,N_10265,N_10303);
nand U10882 (N_10882,N_10050,N_10301);
and U10883 (N_10883,N_10235,N_10248);
nor U10884 (N_10884,N_10068,N_10128);
nand U10885 (N_10885,N_10387,N_10481);
nor U10886 (N_10886,N_10241,N_10211);
xor U10887 (N_10887,N_10428,N_10223);
and U10888 (N_10888,N_10204,N_10165);
and U10889 (N_10889,N_10389,N_10016);
or U10890 (N_10890,N_10283,N_10244);
and U10891 (N_10891,N_10073,N_10197);
and U10892 (N_10892,N_10157,N_10089);
nor U10893 (N_10893,N_10137,N_10245);
or U10894 (N_10894,N_10375,N_10227);
nand U10895 (N_10895,N_10127,N_10139);
nor U10896 (N_10896,N_10010,N_10198);
nand U10897 (N_10897,N_10214,N_10313);
and U10898 (N_10898,N_10486,N_10085);
or U10899 (N_10899,N_10458,N_10417);
or U10900 (N_10900,N_10238,N_10279);
and U10901 (N_10901,N_10133,N_10180);
nand U10902 (N_10902,N_10216,N_10017);
and U10903 (N_10903,N_10241,N_10104);
xnor U10904 (N_10904,N_10330,N_10009);
and U10905 (N_10905,N_10256,N_10241);
nor U10906 (N_10906,N_10171,N_10286);
nor U10907 (N_10907,N_10117,N_10218);
xor U10908 (N_10908,N_10389,N_10177);
xnor U10909 (N_10909,N_10057,N_10255);
xnor U10910 (N_10910,N_10069,N_10251);
or U10911 (N_10911,N_10345,N_10449);
nor U10912 (N_10912,N_10181,N_10287);
xor U10913 (N_10913,N_10020,N_10479);
nor U10914 (N_10914,N_10164,N_10389);
and U10915 (N_10915,N_10408,N_10498);
or U10916 (N_10916,N_10412,N_10085);
xor U10917 (N_10917,N_10314,N_10457);
xnor U10918 (N_10918,N_10465,N_10096);
and U10919 (N_10919,N_10099,N_10177);
nor U10920 (N_10920,N_10293,N_10057);
or U10921 (N_10921,N_10242,N_10345);
xnor U10922 (N_10922,N_10301,N_10442);
or U10923 (N_10923,N_10256,N_10132);
nand U10924 (N_10924,N_10404,N_10178);
xor U10925 (N_10925,N_10273,N_10375);
nand U10926 (N_10926,N_10032,N_10215);
and U10927 (N_10927,N_10263,N_10302);
and U10928 (N_10928,N_10251,N_10299);
nor U10929 (N_10929,N_10435,N_10138);
or U10930 (N_10930,N_10064,N_10344);
or U10931 (N_10931,N_10405,N_10077);
and U10932 (N_10932,N_10277,N_10468);
and U10933 (N_10933,N_10190,N_10012);
xor U10934 (N_10934,N_10227,N_10170);
xnor U10935 (N_10935,N_10370,N_10220);
or U10936 (N_10936,N_10416,N_10047);
and U10937 (N_10937,N_10239,N_10003);
nand U10938 (N_10938,N_10091,N_10180);
and U10939 (N_10939,N_10260,N_10159);
or U10940 (N_10940,N_10341,N_10138);
nor U10941 (N_10941,N_10254,N_10287);
xnor U10942 (N_10942,N_10017,N_10270);
and U10943 (N_10943,N_10116,N_10119);
nor U10944 (N_10944,N_10438,N_10255);
xor U10945 (N_10945,N_10168,N_10080);
nor U10946 (N_10946,N_10388,N_10355);
or U10947 (N_10947,N_10100,N_10413);
xnor U10948 (N_10948,N_10216,N_10293);
nand U10949 (N_10949,N_10459,N_10059);
xor U10950 (N_10950,N_10435,N_10424);
nand U10951 (N_10951,N_10396,N_10209);
or U10952 (N_10952,N_10037,N_10441);
or U10953 (N_10953,N_10220,N_10245);
or U10954 (N_10954,N_10333,N_10087);
nand U10955 (N_10955,N_10031,N_10090);
and U10956 (N_10956,N_10287,N_10173);
or U10957 (N_10957,N_10372,N_10157);
nand U10958 (N_10958,N_10178,N_10408);
xnor U10959 (N_10959,N_10381,N_10286);
xor U10960 (N_10960,N_10119,N_10217);
nor U10961 (N_10961,N_10382,N_10340);
or U10962 (N_10962,N_10252,N_10446);
nand U10963 (N_10963,N_10435,N_10234);
or U10964 (N_10964,N_10229,N_10048);
nand U10965 (N_10965,N_10425,N_10193);
xnor U10966 (N_10966,N_10218,N_10100);
nand U10967 (N_10967,N_10291,N_10298);
or U10968 (N_10968,N_10003,N_10471);
xnor U10969 (N_10969,N_10247,N_10166);
nor U10970 (N_10970,N_10308,N_10394);
nor U10971 (N_10971,N_10101,N_10109);
nand U10972 (N_10972,N_10457,N_10301);
xnor U10973 (N_10973,N_10204,N_10028);
or U10974 (N_10974,N_10108,N_10328);
and U10975 (N_10975,N_10457,N_10339);
xor U10976 (N_10976,N_10193,N_10078);
xnor U10977 (N_10977,N_10129,N_10310);
nand U10978 (N_10978,N_10401,N_10213);
or U10979 (N_10979,N_10397,N_10318);
nand U10980 (N_10980,N_10061,N_10329);
nor U10981 (N_10981,N_10016,N_10115);
nor U10982 (N_10982,N_10445,N_10235);
nand U10983 (N_10983,N_10387,N_10478);
and U10984 (N_10984,N_10146,N_10113);
and U10985 (N_10985,N_10252,N_10384);
xnor U10986 (N_10986,N_10231,N_10493);
nand U10987 (N_10987,N_10201,N_10340);
or U10988 (N_10988,N_10215,N_10095);
or U10989 (N_10989,N_10274,N_10090);
nor U10990 (N_10990,N_10016,N_10333);
nand U10991 (N_10991,N_10340,N_10033);
xor U10992 (N_10992,N_10245,N_10415);
xor U10993 (N_10993,N_10168,N_10124);
or U10994 (N_10994,N_10284,N_10053);
and U10995 (N_10995,N_10071,N_10176);
xnor U10996 (N_10996,N_10331,N_10394);
nor U10997 (N_10997,N_10400,N_10170);
xnor U10998 (N_10998,N_10213,N_10265);
xnor U10999 (N_10999,N_10429,N_10039);
xnor U11000 (N_11000,N_10683,N_10599);
xor U11001 (N_11001,N_10518,N_10592);
nand U11002 (N_11002,N_10891,N_10932);
and U11003 (N_11003,N_10742,N_10686);
nor U11004 (N_11004,N_10974,N_10637);
xor U11005 (N_11005,N_10602,N_10926);
nor U11006 (N_11006,N_10750,N_10636);
or U11007 (N_11007,N_10813,N_10681);
nand U11008 (N_11008,N_10814,N_10820);
nor U11009 (N_11009,N_10741,N_10783);
and U11010 (N_11010,N_10760,N_10991);
nor U11011 (N_11011,N_10740,N_10650);
nor U11012 (N_11012,N_10990,N_10611);
or U11013 (N_11013,N_10789,N_10770);
xor U11014 (N_11014,N_10981,N_10646);
nor U11015 (N_11015,N_10528,N_10852);
or U11016 (N_11016,N_10615,N_10983);
nand U11017 (N_11017,N_10824,N_10643);
and U11018 (N_11018,N_10875,N_10954);
xnor U11019 (N_11019,N_10840,N_10865);
nand U11020 (N_11020,N_10754,N_10648);
and U11021 (N_11021,N_10745,N_10587);
xor U11022 (N_11022,N_10540,N_10778);
nand U11023 (N_11023,N_10775,N_10589);
nor U11024 (N_11024,N_10657,N_10579);
nor U11025 (N_11025,N_10866,N_10805);
or U11026 (N_11026,N_10804,N_10828);
nor U11027 (N_11027,N_10801,N_10645);
xor U11028 (N_11028,N_10664,N_10919);
xor U11029 (N_11029,N_10997,N_10533);
xor U11030 (N_11030,N_10624,N_10556);
xnor U11031 (N_11031,N_10953,N_10895);
nor U11032 (N_11032,N_10771,N_10934);
nor U11033 (N_11033,N_10774,N_10743);
nor U11034 (N_11034,N_10851,N_10928);
nand U11035 (N_11035,N_10816,N_10790);
nor U11036 (N_11036,N_10605,N_10572);
nand U11037 (N_11037,N_10558,N_10765);
nand U11038 (N_11038,N_10652,N_10780);
nand U11039 (N_11039,N_10662,N_10872);
nand U11040 (N_11040,N_10621,N_10784);
nor U11041 (N_11041,N_10554,N_10702);
or U11042 (N_11042,N_10817,N_10810);
nor U11043 (N_11043,N_10994,N_10673);
and U11044 (N_11044,N_10825,N_10956);
or U11045 (N_11045,N_10786,N_10960);
or U11046 (N_11046,N_10730,N_10695);
nor U11047 (N_11047,N_10710,N_10541);
or U11048 (N_11048,N_10758,N_10534);
and U11049 (N_11049,N_10959,N_10502);
and U11050 (N_11050,N_10992,N_10559);
xnor U11051 (N_11051,N_10985,N_10550);
or U11052 (N_11052,N_10867,N_10627);
nand U11053 (N_11053,N_10588,N_10880);
nor U11054 (N_11054,N_10787,N_10620);
and U11055 (N_11055,N_10958,N_10669);
nand U11056 (N_11056,N_10576,N_10578);
nor U11057 (N_11057,N_10980,N_10670);
xnor U11058 (N_11058,N_10678,N_10649);
nand U11059 (N_11059,N_10516,N_10998);
and U11060 (N_11060,N_10827,N_10939);
nor U11061 (N_11061,N_10967,N_10916);
and U11062 (N_11062,N_10699,N_10922);
nand U11063 (N_11063,N_10715,N_10535);
nor U11064 (N_11064,N_10537,N_10603);
and U11065 (N_11065,N_10655,N_10917);
or U11066 (N_11066,N_10769,N_10856);
and U11067 (N_11067,N_10839,N_10949);
xor U11068 (N_11068,N_10716,N_10545);
xnor U11069 (N_11069,N_10952,N_10906);
xnor U11070 (N_11070,N_10580,N_10526);
xnor U11071 (N_11071,N_10723,N_10694);
or U11072 (N_11072,N_10675,N_10799);
nor U11073 (N_11073,N_10630,N_10788);
and U11074 (N_11074,N_10586,N_10964);
or U11075 (N_11075,N_10547,N_10826);
nand U11076 (N_11076,N_10709,N_10843);
and U11077 (N_11077,N_10849,N_10869);
or U11078 (N_11078,N_10806,N_10667);
or U11079 (N_11079,N_10713,N_10846);
nor U11080 (N_11080,N_10882,N_10961);
nor U11081 (N_11081,N_10698,N_10858);
and U11082 (N_11082,N_10890,N_10910);
nor U11083 (N_11083,N_10968,N_10885);
nor U11084 (N_11084,N_10724,N_10505);
or U11085 (N_11085,N_10688,N_10746);
nand U11086 (N_11086,N_10555,N_10687);
or U11087 (N_11087,N_10888,N_10873);
nor U11088 (N_11088,N_10914,N_10703);
or U11089 (N_11089,N_10501,N_10881);
or U11090 (N_11090,N_10847,N_10947);
or U11091 (N_11091,N_10677,N_10900);
nand U11092 (N_11092,N_10552,N_10779);
or U11093 (N_11093,N_10929,N_10921);
or U11094 (N_11094,N_10762,N_10904);
and U11095 (N_11095,N_10692,N_10530);
xor U11096 (N_11096,N_10564,N_10597);
nor U11097 (N_11097,N_10999,N_10631);
xor U11098 (N_11098,N_10976,N_10642);
xnor U11099 (N_11099,N_10903,N_10864);
nand U11100 (N_11100,N_10835,N_10729);
xnor U11101 (N_11101,N_10823,N_10685);
nand U11102 (N_11102,N_10510,N_10819);
nand U11103 (N_11103,N_10855,N_10924);
nand U11104 (N_11104,N_10728,N_10705);
or U11105 (N_11105,N_10508,N_10608);
xor U11106 (N_11106,N_10720,N_10854);
and U11107 (N_11107,N_10634,N_10595);
nor U11108 (N_11108,N_10701,N_10604);
nor U11109 (N_11109,N_10791,N_10513);
or U11110 (N_11110,N_10766,N_10700);
xnor U11111 (N_11111,N_10719,N_10553);
nand U11112 (N_11112,N_10759,N_10944);
or U11113 (N_11113,N_10767,N_10752);
or U11114 (N_11114,N_10706,N_10818);
and U11115 (N_11115,N_10982,N_10593);
or U11116 (N_11116,N_10811,N_10793);
nand U11117 (N_11117,N_10749,N_10581);
or U11118 (N_11118,N_10876,N_10879);
nand U11119 (N_11119,N_10993,N_10575);
and U11120 (N_11120,N_10978,N_10676);
and U11121 (N_11121,N_10711,N_10629);
and U11122 (N_11122,N_10930,N_10551);
xnor U11123 (N_11123,N_10822,N_10606);
or U11124 (N_11124,N_10697,N_10911);
nand U11125 (N_11125,N_10585,N_10561);
nand U11126 (N_11126,N_10659,N_10731);
nor U11127 (N_11127,N_10563,N_10970);
and U11128 (N_11128,N_10607,N_10514);
or U11129 (N_11129,N_10971,N_10923);
xnor U11130 (N_11130,N_10850,N_10567);
nand U11131 (N_11131,N_10800,N_10529);
and U11132 (N_11132,N_10658,N_10682);
and U11133 (N_11133,N_10965,N_10912);
nor U11134 (N_11134,N_10948,N_10899);
and U11135 (N_11135,N_10509,N_10844);
nor U11136 (N_11136,N_10596,N_10918);
nor U11137 (N_11137,N_10506,N_10772);
or U11138 (N_11138,N_10845,N_10972);
nand U11139 (N_11139,N_10755,N_10957);
nor U11140 (N_11140,N_10834,N_10532);
nand U11141 (N_11141,N_10638,N_10739);
and U11142 (N_11142,N_10647,N_10897);
xor U11143 (N_11143,N_10569,N_10773);
nor U11144 (N_11144,N_10761,N_10747);
and U11145 (N_11145,N_10857,N_10886);
or U11146 (N_11146,N_10654,N_10935);
and U11147 (N_11147,N_10777,N_10598);
nand U11148 (N_11148,N_10656,N_10815);
nor U11149 (N_11149,N_10542,N_10950);
nor U11150 (N_11150,N_10566,N_10557);
and U11151 (N_11151,N_10836,N_10898);
xor U11152 (N_11152,N_10641,N_10617);
nand U11153 (N_11153,N_10623,N_10571);
nor U11154 (N_11154,N_10583,N_10582);
xnor U11155 (N_11155,N_10986,N_10691);
nor U11156 (N_11156,N_10523,N_10616);
and U11157 (N_11157,N_10933,N_10915);
nand U11158 (N_11158,N_10909,N_10901);
nand U11159 (N_11159,N_10539,N_10527);
xor U11160 (N_11160,N_10633,N_10946);
nor U11161 (N_11161,N_10560,N_10871);
nand U11162 (N_11162,N_10768,N_10618);
xor U11163 (N_11163,N_10684,N_10521);
nand U11164 (N_11164,N_10635,N_10896);
nor U11165 (N_11165,N_10883,N_10908);
nand U11166 (N_11166,N_10512,N_10601);
xnor U11167 (N_11167,N_10565,N_10781);
xnor U11168 (N_11168,N_10862,N_10966);
or U11169 (N_11169,N_10500,N_10610);
nor U11170 (N_11170,N_10707,N_10722);
nand U11171 (N_11171,N_10744,N_10853);
nand U11172 (N_11172,N_10809,N_10614);
xnor U11173 (N_11173,N_10507,N_10543);
xnor U11174 (N_11174,N_10712,N_10821);
or U11175 (N_11175,N_10763,N_10661);
xor U11176 (N_11176,N_10831,N_10651);
xor U11177 (N_11177,N_10734,N_10548);
xor U11178 (N_11178,N_10927,N_10977);
or U11179 (N_11179,N_10632,N_10984);
nor U11180 (N_11180,N_10737,N_10546);
nor U11181 (N_11181,N_10708,N_10868);
nand U11182 (N_11182,N_10727,N_10942);
or U11183 (N_11183,N_10996,N_10748);
xnor U11184 (N_11184,N_10726,N_10975);
nand U11185 (N_11185,N_10725,N_10861);
nor U11186 (N_11186,N_10536,N_10884);
nor U11187 (N_11187,N_10902,N_10764);
xnor U11188 (N_11188,N_10570,N_10859);
and U11189 (N_11189,N_10830,N_10798);
or U11190 (N_11190,N_10689,N_10802);
nand U11191 (N_11191,N_10690,N_10938);
xnor U11192 (N_11192,N_10522,N_10628);
or U11193 (N_11193,N_10807,N_10538);
and U11194 (N_11194,N_10622,N_10988);
nor U11195 (N_11195,N_10639,N_10979);
or U11196 (N_11196,N_10794,N_10913);
nand U11197 (N_11197,N_10987,N_10733);
and U11198 (N_11198,N_10892,N_10940);
xnor U11199 (N_11199,N_10613,N_10549);
and U11200 (N_11200,N_10889,N_10738);
and U11201 (N_11201,N_10833,N_10568);
nor U11202 (N_11202,N_10841,N_10753);
or U11203 (N_11203,N_10920,N_10936);
xor U11204 (N_11204,N_10842,N_10562);
and U11205 (N_11205,N_10951,N_10941);
or U11206 (N_11206,N_10925,N_10894);
nor U11207 (N_11207,N_10584,N_10797);
and U11208 (N_11208,N_10625,N_10874);
nand U11209 (N_11209,N_10860,N_10785);
nand U11210 (N_11210,N_10515,N_10665);
and U11211 (N_11211,N_10955,N_10878);
nor U11212 (N_11212,N_10674,N_10525);
nor U11213 (N_11213,N_10504,N_10672);
nand U11214 (N_11214,N_10782,N_10590);
and U11215 (N_11215,N_10544,N_10663);
xnor U11216 (N_11216,N_10600,N_10893);
xor U11217 (N_11217,N_10776,N_10680);
xor U11218 (N_11218,N_10640,N_10995);
or U11219 (N_11219,N_10837,N_10679);
xnor U11220 (N_11220,N_10714,N_10963);
nor U11221 (N_11221,N_10653,N_10644);
xnor U11222 (N_11222,N_10693,N_10573);
nand U11223 (N_11223,N_10511,N_10812);
nand U11224 (N_11224,N_10531,N_10905);
nand U11225 (N_11225,N_10696,N_10907);
and U11226 (N_11226,N_10666,N_10704);
nor U11227 (N_11227,N_10626,N_10668);
and U11228 (N_11228,N_10756,N_10863);
xnor U11229 (N_11229,N_10792,N_10838);
or U11230 (N_11230,N_10732,N_10721);
nor U11231 (N_11231,N_10870,N_10832);
and U11232 (N_11232,N_10612,N_10969);
and U11233 (N_11233,N_10503,N_10660);
xnor U11234 (N_11234,N_10803,N_10594);
and U11235 (N_11235,N_10735,N_10943);
nand U11236 (N_11236,N_10577,N_10751);
and U11237 (N_11237,N_10591,N_10931);
and U11238 (N_11238,N_10796,N_10877);
and U11239 (N_11239,N_10989,N_10520);
nor U11240 (N_11240,N_10808,N_10887);
and U11241 (N_11241,N_10829,N_10619);
xor U11242 (N_11242,N_10973,N_10519);
xnor U11243 (N_11243,N_10524,N_10848);
or U11244 (N_11244,N_10945,N_10574);
and U11245 (N_11245,N_10718,N_10937);
xnor U11246 (N_11246,N_10757,N_10609);
nand U11247 (N_11247,N_10517,N_10671);
nor U11248 (N_11248,N_10962,N_10795);
nand U11249 (N_11249,N_10736,N_10717);
nor U11250 (N_11250,N_10504,N_10535);
xor U11251 (N_11251,N_10552,N_10825);
or U11252 (N_11252,N_10741,N_10945);
and U11253 (N_11253,N_10989,N_10633);
nor U11254 (N_11254,N_10961,N_10890);
xor U11255 (N_11255,N_10984,N_10733);
xnor U11256 (N_11256,N_10551,N_10835);
or U11257 (N_11257,N_10742,N_10834);
nor U11258 (N_11258,N_10812,N_10518);
and U11259 (N_11259,N_10672,N_10750);
or U11260 (N_11260,N_10814,N_10707);
nor U11261 (N_11261,N_10767,N_10504);
and U11262 (N_11262,N_10958,N_10792);
and U11263 (N_11263,N_10781,N_10808);
nand U11264 (N_11264,N_10531,N_10946);
nor U11265 (N_11265,N_10653,N_10714);
nand U11266 (N_11266,N_10548,N_10714);
nand U11267 (N_11267,N_10543,N_10944);
xnor U11268 (N_11268,N_10503,N_10895);
nand U11269 (N_11269,N_10951,N_10927);
or U11270 (N_11270,N_10969,N_10716);
nand U11271 (N_11271,N_10618,N_10770);
nor U11272 (N_11272,N_10547,N_10564);
or U11273 (N_11273,N_10838,N_10795);
nor U11274 (N_11274,N_10585,N_10669);
and U11275 (N_11275,N_10555,N_10755);
nand U11276 (N_11276,N_10718,N_10531);
nor U11277 (N_11277,N_10653,N_10743);
xnor U11278 (N_11278,N_10836,N_10583);
nand U11279 (N_11279,N_10869,N_10934);
nor U11280 (N_11280,N_10742,N_10583);
xnor U11281 (N_11281,N_10553,N_10684);
or U11282 (N_11282,N_10595,N_10672);
nor U11283 (N_11283,N_10621,N_10563);
and U11284 (N_11284,N_10503,N_10843);
nand U11285 (N_11285,N_10927,N_10527);
or U11286 (N_11286,N_10903,N_10611);
xnor U11287 (N_11287,N_10559,N_10930);
nand U11288 (N_11288,N_10621,N_10692);
or U11289 (N_11289,N_10956,N_10580);
nand U11290 (N_11290,N_10656,N_10724);
xnor U11291 (N_11291,N_10781,N_10878);
or U11292 (N_11292,N_10665,N_10871);
and U11293 (N_11293,N_10870,N_10747);
xor U11294 (N_11294,N_10655,N_10715);
nand U11295 (N_11295,N_10813,N_10616);
and U11296 (N_11296,N_10786,N_10599);
xor U11297 (N_11297,N_10702,N_10891);
or U11298 (N_11298,N_10633,N_10548);
nand U11299 (N_11299,N_10713,N_10861);
nor U11300 (N_11300,N_10857,N_10985);
or U11301 (N_11301,N_10786,N_10609);
nand U11302 (N_11302,N_10593,N_10713);
or U11303 (N_11303,N_10894,N_10794);
nand U11304 (N_11304,N_10706,N_10956);
nand U11305 (N_11305,N_10926,N_10502);
xnor U11306 (N_11306,N_10816,N_10826);
xor U11307 (N_11307,N_10546,N_10846);
xor U11308 (N_11308,N_10632,N_10887);
nand U11309 (N_11309,N_10546,N_10560);
or U11310 (N_11310,N_10803,N_10736);
nand U11311 (N_11311,N_10941,N_10641);
or U11312 (N_11312,N_10647,N_10862);
or U11313 (N_11313,N_10639,N_10757);
nor U11314 (N_11314,N_10599,N_10813);
or U11315 (N_11315,N_10903,N_10708);
or U11316 (N_11316,N_10985,N_10558);
xor U11317 (N_11317,N_10710,N_10583);
xnor U11318 (N_11318,N_10575,N_10912);
or U11319 (N_11319,N_10782,N_10764);
or U11320 (N_11320,N_10809,N_10702);
and U11321 (N_11321,N_10897,N_10831);
or U11322 (N_11322,N_10519,N_10801);
nor U11323 (N_11323,N_10790,N_10569);
and U11324 (N_11324,N_10780,N_10871);
nor U11325 (N_11325,N_10972,N_10668);
nand U11326 (N_11326,N_10679,N_10744);
and U11327 (N_11327,N_10608,N_10679);
nor U11328 (N_11328,N_10979,N_10650);
nor U11329 (N_11329,N_10936,N_10896);
nand U11330 (N_11330,N_10912,N_10861);
nand U11331 (N_11331,N_10690,N_10743);
and U11332 (N_11332,N_10605,N_10577);
or U11333 (N_11333,N_10991,N_10698);
or U11334 (N_11334,N_10724,N_10971);
and U11335 (N_11335,N_10786,N_10777);
nor U11336 (N_11336,N_10726,N_10614);
nor U11337 (N_11337,N_10819,N_10895);
xnor U11338 (N_11338,N_10905,N_10571);
and U11339 (N_11339,N_10879,N_10693);
and U11340 (N_11340,N_10953,N_10564);
xnor U11341 (N_11341,N_10583,N_10966);
xnor U11342 (N_11342,N_10712,N_10544);
nor U11343 (N_11343,N_10703,N_10901);
and U11344 (N_11344,N_10520,N_10757);
or U11345 (N_11345,N_10545,N_10728);
or U11346 (N_11346,N_10805,N_10606);
and U11347 (N_11347,N_10925,N_10657);
and U11348 (N_11348,N_10680,N_10758);
nand U11349 (N_11349,N_10665,N_10899);
nand U11350 (N_11350,N_10890,N_10742);
and U11351 (N_11351,N_10990,N_10606);
or U11352 (N_11352,N_10899,N_10652);
nor U11353 (N_11353,N_10675,N_10669);
nand U11354 (N_11354,N_10589,N_10901);
xnor U11355 (N_11355,N_10567,N_10648);
nand U11356 (N_11356,N_10959,N_10993);
nand U11357 (N_11357,N_10646,N_10519);
xnor U11358 (N_11358,N_10604,N_10839);
nor U11359 (N_11359,N_10563,N_10545);
nand U11360 (N_11360,N_10750,N_10891);
xnor U11361 (N_11361,N_10600,N_10629);
or U11362 (N_11362,N_10570,N_10658);
or U11363 (N_11363,N_10507,N_10876);
xnor U11364 (N_11364,N_10886,N_10727);
nor U11365 (N_11365,N_10660,N_10760);
nor U11366 (N_11366,N_10755,N_10700);
nand U11367 (N_11367,N_10544,N_10885);
nand U11368 (N_11368,N_10987,N_10616);
xor U11369 (N_11369,N_10506,N_10709);
nand U11370 (N_11370,N_10853,N_10826);
and U11371 (N_11371,N_10786,N_10858);
nor U11372 (N_11372,N_10629,N_10945);
nand U11373 (N_11373,N_10548,N_10502);
nand U11374 (N_11374,N_10538,N_10759);
nand U11375 (N_11375,N_10766,N_10502);
nor U11376 (N_11376,N_10553,N_10839);
and U11377 (N_11377,N_10602,N_10886);
and U11378 (N_11378,N_10942,N_10794);
and U11379 (N_11379,N_10892,N_10552);
xor U11380 (N_11380,N_10745,N_10608);
or U11381 (N_11381,N_10614,N_10853);
or U11382 (N_11382,N_10874,N_10944);
nand U11383 (N_11383,N_10921,N_10682);
or U11384 (N_11384,N_10704,N_10813);
nand U11385 (N_11385,N_10836,N_10575);
or U11386 (N_11386,N_10582,N_10567);
xor U11387 (N_11387,N_10905,N_10924);
nand U11388 (N_11388,N_10534,N_10589);
nor U11389 (N_11389,N_10525,N_10961);
and U11390 (N_11390,N_10546,N_10777);
or U11391 (N_11391,N_10789,N_10526);
nor U11392 (N_11392,N_10566,N_10714);
nor U11393 (N_11393,N_10805,N_10680);
nor U11394 (N_11394,N_10572,N_10683);
nand U11395 (N_11395,N_10796,N_10836);
nand U11396 (N_11396,N_10906,N_10789);
and U11397 (N_11397,N_10541,N_10557);
or U11398 (N_11398,N_10730,N_10750);
and U11399 (N_11399,N_10772,N_10544);
or U11400 (N_11400,N_10730,N_10816);
nand U11401 (N_11401,N_10674,N_10987);
xor U11402 (N_11402,N_10538,N_10731);
nor U11403 (N_11403,N_10700,N_10582);
nor U11404 (N_11404,N_10530,N_10729);
nor U11405 (N_11405,N_10694,N_10935);
or U11406 (N_11406,N_10954,N_10801);
xnor U11407 (N_11407,N_10613,N_10948);
nand U11408 (N_11408,N_10887,N_10793);
nand U11409 (N_11409,N_10972,N_10746);
and U11410 (N_11410,N_10707,N_10749);
or U11411 (N_11411,N_10903,N_10865);
and U11412 (N_11412,N_10538,N_10675);
nand U11413 (N_11413,N_10552,N_10877);
and U11414 (N_11414,N_10640,N_10550);
xnor U11415 (N_11415,N_10957,N_10878);
and U11416 (N_11416,N_10812,N_10869);
xor U11417 (N_11417,N_10565,N_10668);
and U11418 (N_11418,N_10503,N_10802);
xnor U11419 (N_11419,N_10703,N_10647);
nand U11420 (N_11420,N_10979,N_10575);
nor U11421 (N_11421,N_10873,N_10981);
or U11422 (N_11422,N_10843,N_10757);
nand U11423 (N_11423,N_10717,N_10719);
nor U11424 (N_11424,N_10877,N_10616);
nand U11425 (N_11425,N_10521,N_10622);
nor U11426 (N_11426,N_10516,N_10697);
nand U11427 (N_11427,N_10641,N_10587);
and U11428 (N_11428,N_10790,N_10635);
xor U11429 (N_11429,N_10604,N_10891);
nor U11430 (N_11430,N_10933,N_10797);
xnor U11431 (N_11431,N_10988,N_10924);
nand U11432 (N_11432,N_10898,N_10811);
nor U11433 (N_11433,N_10591,N_10513);
nor U11434 (N_11434,N_10639,N_10688);
and U11435 (N_11435,N_10922,N_10727);
nor U11436 (N_11436,N_10664,N_10819);
or U11437 (N_11437,N_10811,N_10563);
nand U11438 (N_11438,N_10627,N_10586);
nor U11439 (N_11439,N_10893,N_10739);
and U11440 (N_11440,N_10656,N_10553);
xor U11441 (N_11441,N_10749,N_10798);
xor U11442 (N_11442,N_10890,N_10578);
nor U11443 (N_11443,N_10839,N_10821);
nor U11444 (N_11444,N_10881,N_10502);
or U11445 (N_11445,N_10532,N_10906);
nand U11446 (N_11446,N_10705,N_10625);
or U11447 (N_11447,N_10827,N_10655);
and U11448 (N_11448,N_10991,N_10562);
nor U11449 (N_11449,N_10722,N_10644);
or U11450 (N_11450,N_10523,N_10948);
nand U11451 (N_11451,N_10968,N_10725);
nand U11452 (N_11452,N_10519,N_10764);
nand U11453 (N_11453,N_10543,N_10525);
nand U11454 (N_11454,N_10914,N_10525);
and U11455 (N_11455,N_10956,N_10821);
and U11456 (N_11456,N_10947,N_10557);
xnor U11457 (N_11457,N_10582,N_10679);
nor U11458 (N_11458,N_10882,N_10991);
and U11459 (N_11459,N_10975,N_10887);
or U11460 (N_11460,N_10539,N_10531);
or U11461 (N_11461,N_10572,N_10882);
or U11462 (N_11462,N_10789,N_10956);
xor U11463 (N_11463,N_10583,N_10539);
xor U11464 (N_11464,N_10697,N_10887);
or U11465 (N_11465,N_10956,N_10817);
xor U11466 (N_11466,N_10689,N_10675);
nor U11467 (N_11467,N_10922,N_10706);
nand U11468 (N_11468,N_10630,N_10649);
xnor U11469 (N_11469,N_10732,N_10652);
and U11470 (N_11470,N_10517,N_10752);
and U11471 (N_11471,N_10583,N_10774);
nor U11472 (N_11472,N_10810,N_10682);
nand U11473 (N_11473,N_10898,N_10562);
and U11474 (N_11474,N_10662,N_10845);
or U11475 (N_11475,N_10866,N_10961);
nand U11476 (N_11476,N_10712,N_10767);
and U11477 (N_11477,N_10777,N_10983);
xnor U11478 (N_11478,N_10721,N_10766);
and U11479 (N_11479,N_10502,N_10659);
and U11480 (N_11480,N_10812,N_10799);
nor U11481 (N_11481,N_10714,N_10613);
nand U11482 (N_11482,N_10619,N_10592);
nand U11483 (N_11483,N_10764,N_10521);
nand U11484 (N_11484,N_10592,N_10691);
nand U11485 (N_11485,N_10919,N_10594);
nand U11486 (N_11486,N_10768,N_10556);
nor U11487 (N_11487,N_10919,N_10848);
nor U11488 (N_11488,N_10812,N_10597);
nand U11489 (N_11489,N_10681,N_10727);
nor U11490 (N_11490,N_10793,N_10852);
nand U11491 (N_11491,N_10637,N_10692);
nor U11492 (N_11492,N_10679,N_10853);
xnor U11493 (N_11493,N_10908,N_10804);
nand U11494 (N_11494,N_10771,N_10519);
or U11495 (N_11495,N_10666,N_10837);
nor U11496 (N_11496,N_10778,N_10648);
or U11497 (N_11497,N_10986,N_10643);
xor U11498 (N_11498,N_10975,N_10599);
xnor U11499 (N_11499,N_10790,N_10936);
or U11500 (N_11500,N_11105,N_11017);
xnor U11501 (N_11501,N_11455,N_11008);
xor U11502 (N_11502,N_11078,N_11360);
and U11503 (N_11503,N_11386,N_11185);
or U11504 (N_11504,N_11465,N_11183);
nand U11505 (N_11505,N_11088,N_11231);
nor U11506 (N_11506,N_11223,N_11311);
nand U11507 (N_11507,N_11479,N_11257);
nor U11508 (N_11508,N_11038,N_11470);
nand U11509 (N_11509,N_11268,N_11300);
xor U11510 (N_11510,N_11139,N_11137);
or U11511 (N_11511,N_11295,N_11187);
nor U11512 (N_11512,N_11372,N_11224);
nand U11513 (N_11513,N_11288,N_11081);
or U11514 (N_11514,N_11179,N_11128);
or U11515 (N_11515,N_11459,N_11389);
or U11516 (N_11516,N_11043,N_11405);
or U11517 (N_11517,N_11334,N_11358);
nor U11518 (N_11518,N_11423,N_11165);
and U11519 (N_11519,N_11461,N_11339);
and U11520 (N_11520,N_11033,N_11487);
nand U11521 (N_11521,N_11407,N_11271);
xnor U11522 (N_11522,N_11205,N_11316);
xor U11523 (N_11523,N_11041,N_11012);
nand U11524 (N_11524,N_11260,N_11378);
or U11525 (N_11525,N_11091,N_11029);
and U11526 (N_11526,N_11493,N_11480);
nor U11527 (N_11527,N_11049,N_11433);
nor U11528 (N_11528,N_11394,N_11135);
xnor U11529 (N_11529,N_11286,N_11429);
nand U11530 (N_11530,N_11151,N_11208);
nand U11531 (N_11531,N_11471,N_11416);
or U11532 (N_11532,N_11406,N_11190);
and U11533 (N_11533,N_11467,N_11337);
xor U11534 (N_11534,N_11152,N_11004);
nand U11535 (N_11535,N_11198,N_11374);
and U11536 (N_11536,N_11401,N_11212);
nor U11537 (N_11537,N_11228,N_11098);
xor U11538 (N_11538,N_11189,N_11209);
nor U11539 (N_11539,N_11133,N_11166);
nand U11540 (N_11540,N_11227,N_11277);
nand U11541 (N_11541,N_11174,N_11381);
nand U11542 (N_11542,N_11134,N_11248);
and U11543 (N_11543,N_11267,N_11296);
nor U11544 (N_11544,N_11169,N_11379);
nor U11545 (N_11545,N_11236,N_11213);
nand U11546 (N_11546,N_11283,N_11235);
or U11547 (N_11547,N_11168,N_11290);
or U11548 (N_11548,N_11232,N_11246);
and U11549 (N_11549,N_11011,N_11380);
nand U11550 (N_11550,N_11278,N_11454);
or U11551 (N_11551,N_11341,N_11330);
nand U11552 (N_11552,N_11347,N_11097);
nand U11553 (N_11553,N_11320,N_11391);
or U11554 (N_11554,N_11201,N_11426);
xor U11555 (N_11555,N_11154,N_11481);
or U11556 (N_11556,N_11001,N_11450);
nor U11557 (N_11557,N_11425,N_11475);
nor U11558 (N_11558,N_11106,N_11292);
and U11559 (N_11559,N_11448,N_11441);
or U11560 (N_11560,N_11349,N_11181);
and U11561 (N_11561,N_11006,N_11484);
nand U11562 (N_11562,N_11393,N_11101);
nand U11563 (N_11563,N_11039,N_11477);
and U11564 (N_11564,N_11333,N_11009);
nand U11565 (N_11565,N_11331,N_11072);
and U11566 (N_11566,N_11457,N_11304);
and U11567 (N_11567,N_11387,N_11285);
nand U11568 (N_11568,N_11289,N_11023);
nor U11569 (N_11569,N_11392,N_11027);
nand U11570 (N_11570,N_11436,N_11013);
or U11571 (N_11571,N_11469,N_11022);
nor U11572 (N_11572,N_11431,N_11419);
or U11573 (N_11573,N_11269,N_11002);
xor U11574 (N_11574,N_11014,N_11370);
or U11575 (N_11575,N_11282,N_11400);
xnor U11576 (N_11576,N_11335,N_11108);
nor U11577 (N_11577,N_11411,N_11329);
xor U11578 (N_11578,N_11412,N_11144);
or U11579 (N_11579,N_11059,N_11218);
or U11580 (N_11580,N_11308,N_11030);
and U11581 (N_11581,N_11262,N_11453);
nor U11582 (N_11582,N_11353,N_11404);
nand U11583 (N_11583,N_11156,N_11321);
and U11584 (N_11584,N_11395,N_11140);
nor U11585 (N_11585,N_11463,N_11089);
nand U11586 (N_11586,N_11159,N_11415);
or U11587 (N_11587,N_11136,N_11090);
nand U11588 (N_11588,N_11221,N_11015);
nand U11589 (N_11589,N_11397,N_11214);
nand U11590 (N_11590,N_11200,N_11468);
xor U11591 (N_11591,N_11052,N_11068);
nor U11592 (N_11592,N_11344,N_11417);
nor U11593 (N_11593,N_11149,N_11215);
or U11594 (N_11594,N_11279,N_11112);
and U11595 (N_11595,N_11444,N_11003);
or U11596 (N_11596,N_11301,N_11074);
or U11597 (N_11597,N_11146,N_11439);
nor U11598 (N_11598,N_11377,N_11010);
or U11599 (N_11599,N_11026,N_11162);
nand U11600 (N_11600,N_11025,N_11178);
nor U11601 (N_11601,N_11413,N_11371);
nor U11602 (N_11602,N_11414,N_11206);
xnor U11603 (N_11603,N_11297,N_11352);
nor U11604 (N_11604,N_11302,N_11099);
nand U11605 (N_11605,N_11207,N_11061);
or U11606 (N_11606,N_11382,N_11265);
nand U11607 (N_11607,N_11182,N_11366);
or U11608 (N_11608,N_11031,N_11126);
nor U11609 (N_11609,N_11202,N_11298);
xor U11610 (N_11610,N_11238,N_11494);
nor U11611 (N_11611,N_11194,N_11409);
xor U11612 (N_11612,N_11195,N_11109);
nor U11613 (N_11613,N_11186,N_11233);
or U11614 (N_11614,N_11239,N_11045);
and U11615 (N_11615,N_11199,N_11222);
xnor U11616 (N_11616,N_11161,N_11402);
nor U11617 (N_11617,N_11150,N_11067);
or U11618 (N_11618,N_11092,N_11065);
and U11619 (N_11619,N_11388,N_11082);
nand U11620 (N_11620,N_11427,N_11107);
or U11621 (N_11621,N_11491,N_11398);
nand U11622 (N_11622,N_11111,N_11021);
xor U11623 (N_11623,N_11057,N_11087);
nand U11624 (N_11624,N_11259,N_11476);
xor U11625 (N_11625,N_11359,N_11473);
xnor U11626 (N_11626,N_11066,N_11355);
or U11627 (N_11627,N_11390,N_11266);
xnor U11628 (N_11628,N_11251,N_11153);
xor U11629 (N_11629,N_11340,N_11037);
nand U11630 (N_11630,N_11452,N_11119);
or U11631 (N_11631,N_11070,N_11115);
xor U11632 (N_11632,N_11356,N_11080);
nand U11633 (N_11633,N_11142,N_11328);
xnor U11634 (N_11634,N_11141,N_11122);
and U11635 (N_11635,N_11495,N_11310);
or U11636 (N_11636,N_11281,N_11103);
nor U11637 (N_11637,N_11170,N_11244);
and U11638 (N_11638,N_11367,N_11273);
nor U11639 (N_11639,N_11458,N_11184);
nor U11640 (N_11640,N_11164,N_11275);
xor U11641 (N_11641,N_11307,N_11188);
nand U11642 (N_11642,N_11157,N_11451);
nor U11643 (N_11643,N_11250,N_11255);
or U11644 (N_11644,N_11028,N_11102);
or U11645 (N_11645,N_11226,N_11326);
or U11646 (N_11646,N_11132,N_11120);
and U11647 (N_11647,N_11060,N_11193);
and U11648 (N_11648,N_11261,N_11293);
xnor U11649 (N_11649,N_11242,N_11093);
and U11650 (N_11650,N_11483,N_11368);
xnor U11651 (N_11651,N_11264,N_11464);
nand U11652 (N_11652,N_11077,N_11420);
or U11653 (N_11653,N_11210,N_11424);
nor U11654 (N_11654,N_11466,N_11247);
or U11655 (N_11655,N_11270,N_11354);
or U11656 (N_11656,N_11287,N_11249);
nand U11657 (N_11657,N_11440,N_11094);
and U11658 (N_11658,N_11131,N_11138);
or U11659 (N_11659,N_11217,N_11158);
nor U11660 (N_11660,N_11498,N_11113);
nand U11661 (N_11661,N_11376,N_11050);
and U11662 (N_11662,N_11241,N_11034);
and U11663 (N_11663,N_11032,N_11220);
nand U11664 (N_11664,N_11121,N_11410);
nor U11665 (N_11665,N_11348,N_11056);
nand U11666 (N_11666,N_11462,N_11084);
nand U11667 (N_11667,N_11016,N_11042);
xnor U11668 (N_11668,N_11317,N_11234);
nor U11669 (N_11669,N_11143,N_11211);
nand U11670 (N_11670,N_11312,N_11063);
nand U11671 (N_11671,N_11314,N_11237);
or U11672 (N_11672,N_11445,N_11438);
nand U11673 (N_11673,N_11350,N_11305);
or U11674 (N_11674,N_11203,N_11100);
nor U11675 (N_11675,N_11252,N_11005);
or U11676 (N_11676,N_11245,N_11253);
or U11677 (N_11677,N_11129,N_11396);
and U11678 (N_11678,N_11430,N_11125);
and U11679 (N_11679,N_11460,N_11204);
nor U11680 (N_11680,N_11155,N_11299);
xnor U11681 (N_11681,N_11319,N_11075);
or U11682 (N_11682,N_11073,N_11216);
or U11683 (N_11683,N_11171,N_11474);
xor U11684 (N_11684,N_11258,N_11332);
and U11685 (N_11685,N_11361,N_11276);
nor U11686 (N_11686,N_11422,N_11428);
xor U11687 (N_11687,N_11446,N_11083);
xor U11688 (N_11688,N_11116,N_11180);
and U11689 (N_11689,N_11384,N_11338);
nor U11690 (N_11690,N_11054,N_11432);
and U11691 (N_11691,N_11323,N_11434);
nor U11692 (N_11692,N_11291,N_11047);
xor U11693 (N_11693,N_11365,N_11327);
or U11694 (N_11694,N_11325,N_11160);
nor U11695 (N_11695,N_11062,N_11385);
or U11696 (N_11696,N_11117,N_11020);
nor U11697 (N_11697,N_11272,N_11486);
nor U11698 (N_11698,N_11399,N_11167);
nor U11699 (N_11699,N_11053,N_11123);
xnor U11700 (N_11700,N_11256,N_11375);
xnor U11701 (N_11701,N_11024,N_11309);
nand U11702 (N_11702,N_11225,N_11069);
nor U11703 (N_11703,N_11274,N_11254);
nand U11704 (N_11704,N_11369,N_11343);
or U11705 (N_11705,N_11449,N_11342);
xnor U11706 (N_11706,N_11048,N_11364);
xnor U11707 (N_11707,N_11408,N_11000);
nor U11708 (N_11708,N_11315,N_11478);
nand U11709 (N_11709,N_11124,N_11345);
xor U11710 (N_11710,N_11240,N_11497);
or U11711 (N_11711,N_11071,N_11346);
and U11712 (N_11712,N_11148,N_11130);
nand U11713 (N_11713,N_11040,N_11230);
nor U11714 (N_11714,N_11055,N_11303);
or U11715 (N_11715,N_11173,N_11229);
or U11716 (N_11716,N_11177,N_11019);
nand U11717 (N_11717,N_11196,N_11351);
nand U11718 (N_11718,N_11482,N_11362);
nor U11719 (N_11719,N_11064,N_11456);
nand U11720 (N_11720,N_11263,N_11175);
nor U11721 (N_11721,N_11104,N_11163);
nand U11722 (N_11722,N_11145,N_11421);
nand U11723 (N_11723,N_11058,N_11191);
xnor U11724 (N_11724,N_11051,N_11085);
xor U11725 (N_11725,N_11172,N_11007);
xor U11726 (N_11726,N_11018,N_11114);
nand U11727 (N_11727,N_11219,N_11313);
xnor U11728 (N_11728,N_11490,N_11499);
nand U11729 (N_11729,N_11324,N_11363);
xnor U11730 (N_11730,N_11306,N_11418);
and U11731 (N_11731,N_11046,N_11197);
or U11732 (N_11732,N_11294,N_11096);
nor U11733 (N_11733,N_11403,N_11192);
or U11734 (N_11734,N_11447,N_11443);
or U11735 (N_11735,N_11243,N_11147);
and U11736 (N_11736,N_11496,N_11118);
xnor U11737 (N_11737,N_11079,N_11036);
nor U11738 (N_11738,N_11127,N_11280);
nor U11739 (N_11739,N_11086,N_11095);
xor U11740 (N_11740,N_11318,N_11035);
nand U11741 (N_11741,N_11383,N_11489);
nand U11742 (N_11742,N_11284,N_11485);
nand U11743 (N_11743,N_11373,N_11435);
or U11744 (N_11744,N_11357,N_11044);
nand U11745 (N_11745,N_11488,N_11492);
or U11746 (N_11746,N_11336,N_11442);
and U11747 (N_11747,N_11176,N_11437);
or U11748 (N_11748,N_11472,N_11322);
and U11749 (N_11749,N_11110,N_11076);
or U11750 (N_11750,N_11157,N_11426);
xnor U11751 (N_11751,N_11211,N_11080);
and U11752 (N_11752,N_11046,N_11080);
or U11753 (N_11753,N_11360,N_11033);
nand U11754 (N_11754,N_11115,N_11459);
nor U11755 (N_11755,N_11013,N_11156);
nor U11756 (N_11756,N_11006,N_11055);
or U11757 (N_11757,N_11206,N_11070);
nand U11758 (N_11758,N_11013,N_11091);
and U11759 (N_11759,N_11281,N_11074);
or U11760 (N_11760,N_11218,N_11486);
and U11761 (N_11761,N_11441,N_11452);
nand U11762 (N_11762,N_11017,N_11088);
nand U11763 (N_11763,N_11068,N_11072);
xor U11764 (N_11764,N_11229,N_11014);
and U11765 (N_11765,N_11384,N_11077);
or U11766 (N_11766,N_11225,N_11485);
nand U11767 (N_11767,N_11471,N_11472);
xor U11768 (N_11768,N_11392,N_11311);
or U11769 (N_11769,N_11137,N_11234);
and U11770 (N_11770,N_11151,N_11055);
or U11771 (N_11771,N_11332,N_11234);
xnor U11772 (N_11772,N_11111,N_11399);
xnor U11773 (N_11773,N_11064,N_11134);
nor U11774 (N_11774,N_11173,N_11055);
nor U11775 (N_11775,N_11366,N_11381);
nor U11776 (N_11776,N_11414,N_11046);
and U11777 (N_11777,N_11148,N_11247);
xor U11778 (N_11778,N_11269,N_11106);
and U11779 (N_11779,N_11477,N_11282);
xnor U11780 (N_11780,N_11003,N_11131);
xor U11781 (N_11781,N_11132,N_11471);
and U11782 (N_11782,N_11313,N_11156);
nand U11783 (N_11783,N_11328,N_11358);
and U11784 (N_11784,N_11253,N_11447);
nand U11785 (N_11785,N_11157,N_11106);
and U11786 (N_11786,N_11436,N_11219);
and U11787 (N_11787,N_11268,N_11194);
and U11788 (N_11788,N_11281,N_11288);
nand U11789 (N_11789,N_11016,N_11389);
and U11790 (N_11790,N_11098,N_11421);
xnor U11791 (N_11791,N_11285,N_11047);
xor U11792 (N_11792,N_11232,N_11309);
and U11793 (N_11793,N_11370,N_11199);
xnor U11794 (N_11794,N_11168,N_11104);
or U11795 (N_11795,N_11131,N_11081);
xnor U11796 (N_11796,N_11051,N_11019);
or U11797 (N_11797,N_11251,N_11322);
nand U11798 (N_11798,N_11282,N_11316);
nor U11799 (N_11799,N_11401,N_11097);
or U11800 (N_11800,N_11071,N_11334);
nor U11801 (N_11801,N_11064,N_11466);
and U11802 (N_11802,N_11401,N_11061);
xor U11803 (N_11803,N_11000,N_11266);
and U11804 (N_11804,N_11307,N_11310);
nand U11805 (N_11805,N_11268,N_11262);
and U11806 (N_11806,N_11200,N_11160);
xnor U11807 (N_11807,N_11486,N_11348);
xnor U11808 (N_11808,N_11229,N_11414);
nand U11809 (N_11809,N_11112,N_11033);
nor U11810 (N_11810,N_11043,N_11258);
nor U11811 (N_11811,N_11036,N_11498);
nor U11812 (N_11812,N_11221,N_11307);
nor U11813 (N_11813,N_11289,N_11137);
or U11814 (N_11814,N_11046,N_11053);
or U11815 (N_11815,N_11026,N_11117);
nor U11816 (N_11816,N_11409,N_11086);
or U11817 (N_11817,N_11406,N_11132);
xnor U11818 (N_11818,N_11284,N_11031);
nor U11819 (N_11819,N_11257,N_11402);
xor U11820 (N_11820,N_11282,N_11348);
nand U11821 (N_11821,N_11378,N_11499);
and U11822 (N_11822,N_11212,N_11042);
and U11823 (N_11823,N_11231,N_11441);
xor U11824 (N_11824,N_11465,N_11273);
and U11825 (N_11825,N_11327,N_11166);
nand U11826 (N_11826,N_11420,N_11146);
nor U11827 (N_11827,N_11330,N_11421);
and U11828 (N_11828,N_11025,N_11196);
and U11829 (N_11829,N_11285,N_11189);
nor U11830 (N_11830,N_11183,N_11196);
nor U11831 (N_11831,N_11379,N_11021);
nand U11832 (N_11832,N_11343,N_11144);
or U11833 (N_11833,N_11424,N_11026);
or U11834 (N_11834,N_11430,N_11158);
or U11835 (N_11835,N_11244,N_11430);
nand U11836 (N_11836,N_11371,N_11053);
and U11837 (N_11837,N_11064,N_11214);
or U11838 (N_11838,N_11236,N_11303);
xnor U11839 (N_11839,N_11473,N_11228);
and U11840 (N_11840,N_11153,N_11118);
xnor U11841 (N_11841,N_11375,N_11146);
or U11842 (N_11842,N_11331,N_11021);
xor U11843 (N_11843,N_11451,N_11221);
nand U11844 (N_11844,N_11108,N_11162);
nand U11845 (N_11845,N_11005,N_11185);
nand U11846 (N_11846,N_11346,N_11197);
and U11847 (N_11847,N_11097,N_11224);
xor U11848 (N_11848,N_11115,N_11401);
or U11849 (N_11849,N_11142,N_11473);
or U11850 (N_11850,N_11168,N_11349);
nand U11851 (N_11851,N_11145,N_11367);
nand U11852 (N_11852,N_11126,N_11480);
nor U11853 (N_11853,N_11321,N_11096);
nand U11854 (N_11854,N_11039,N_11014);
nand U11855 (N_11855,N_11280,N_11380);
or U11856 (N_11856,N_11325,N_11297);
nor U11857 (N_11857,N_11003,N_11309);
xnor U11858 (N_11858,N_11085,N_11144);
nor U11859 (N_11859,N_11309,N_11180);
xor U11860 (N_11860,N_11139,N_11046);
and U11861 (N_11861,N_11185,N_11204);
nor U11862 (N_11862,N_11176,N_11427);
or U11863 (N_11863,N_11149,N_11328);
nand U11864 (N_11864,N_11217,N_11264);
and U11865 (N_11865,N_11243,N_11119);
xnor U11866 (N_11866,N_11412,N_11374);
nor U11867 (N_11867,N_11180,N_11450);
nand U11868 (N_11868,N_11373,N_11087);
xor U11869 (N_11869,N_11419,N_11200);
or U11870 (N_11870,N_11397,N_11469);
and U11871 (N_11871,N_11433,N_11469);
xor U11872 (N_11872,N_11183,N_11070);
nand U11873 (N_11873,N_11246,N_11099);
xor U11874 (N_11874,N_11307,N_11056);
or U11875 (N_11875,N_11232,N_11207);
or U11876 (N_11876,N_11266,N_11042);
xnor U11877 (N_11877,N_11132,N_11051);
nor U11878 (N_11878,N_11354,N_11353);
nor U11879 (N_11879,N_11475,N_11325);
xnor U11880 (N_11880,N_11288,N_11356);
and U11881 (N_11881,N_11119,N_11212);
and U11882 (N_11882,N_11390,N_11483);
and U11883 (N_11883,N_11367,N_11114);
and U11884 (N_11884,N_11185,N_11225);
or U11885 (N_11885,N_11297,N_11494);
xor U11886 (N_11886,N_11442,N_11271);
nor U11887 (N_11887,N_11104,N_11378);
xor U11888 (N_11888,N_11147,N_11382);
and U11889 (N_11889,N_11089,N_11330);
and U11890 (N_11890,N_11114,N_11271);
and U11891 (N_11891,N_11061,N_11474);
and U11892 (N_11892,N_11287,N_11363);
and U11893 (N_11893,N_11110,N_11405);
xor U11894 (N_11894,N_11139,N_11262);
nor U11895 (N_11895,N_11177,N_11431);
nand U11896 (N_11896,N_11083,N_11208);
xor U11897 (N_11897,N_11115,N_11054);
xor U11898 (N_11898,N_11135,N_11320);
nand U11899 (N_11899,N_11181,N_11392);
nor U11900 (N_11900,N_11220,N_11493);
and U11901 (N_11901,N_11489,N_11398);
xor U11902 (N_11902,N_11048,N_11447);
nor U11903 (N_11903,N_11343,N_11293);
nand U11904 (N_11904,N_11114,N_11090);
nand U11905 (N_11905,N_11336,N_11136);
and U11906 (N_11906,N_11289,N_11339);
nor U11907 (N_11907,N_11318,N_11211);
xor U11908 (N_11908,N_11074,N_11476);
or U11909 (N_11909,N_11282,N_11150);
and U11910 (N_11910,N_11470,N_11479);
xor U11911 (N_11911,N_11356,N_11443);
and U11912 (N_11912,N_11434,N_11070);
nand U11913 (N_11913,N_11300,N_11163);
or U11914 (N_11914,N_11438,N_11011);
nor U11915 (N_11915,N_11292,N_11483);
xnor U11916 (N_11916,N_11072,N_11417);
nor U11917 (N_11917,N_11118,N_11406);
xnor U11918 (N_11918,N_11488,N_11405);
nor U11919 (N_11919,N_11115,N_11037);
or U11920 (N_11920,N_11259,N_11281);
xor U11921 (N_11921,N_11120,N_11110);
or U11922 (N_11922,N_11230,N_11286);
and U11923 (N_11923,N_11286,N_11292);
xor U11924 (N_11924,N_11138,N_11491);
and U11925 (N_11925,N_11106,N_11391);
or U11926 (N_11926,N_11379,N_11229);
and U11927 (N_11927,N_11407,N_11397);
xnor U11928 (N_11928,N_11095,N_11417);
or U11929 (N_11929,N_11040,N_11150);
xnor U11930 (N_11930,N_11380,N_11048);
nor U11931 (N_11931,N_11254,N_11285);
nor U11932 (N_11932,N_11450,N_11391);
nor U11933 (N_11933,N_11076,N_11170);
and U11934 (N_11934,N_11413,N_11417);
or U11935 (N_11935,N_11139,N_11152);
nor U11936 (N_11936,N_11156,N_11290);
nand U11937 (N_11937,N_11006,N_11375);
nor U11938 (N_11938,N_11314,N_11308);
and U11939 (N_11939,N_11287,N_11189);
nand U11940 (N_11940,N_11433,N_11363);
and U11941 (N_11941,N_11303,N_11351);
or U11942 (N_11942,N_11022,N_11430);
nor U11943 (N_11943,N_11140,N_11470);
nand U11944 (N_11944,N_11102,N_11457);
nor U11945 (N_11945,N_11105,N_11022);
or U11946 (N_11946,N_11228,N_11390);
xnor U11947 (N_11947,N_11134,N_11420);
and U11948 (N_11948,N_11174,N_11284);
and U11949 (N_11949,N_11111,N_11458);
and U11950 (N_11950,N_11103,N_11458);
nor U11951 (N_11951,N_11487,N_11143);
or U11952 (N_11952,N_11414,N_11172);
and U11953 (N_11953,N_11110,N_11107);
or U11954 (N_11954,N_11482,N_11290);
and U11955 (N_11955,N_11445,N_11030);
nor U11956 (N_11956,N_11142,N_11115);
or U11957 (N_11957,N_11065,N_11492);
or U11958 (N_11958,N_11119,N_11213);
nor U11959 (N_11959,N_11476,N_11489);
and U11960 (N_11960,N_11208,N_11228);
xor U11961 (N_11961,N_11188,N_11293);
and U11962 (N_11962,N_11373,N_11163);
and U11963 (N_11963,N_11348,N_11077);
or U11964 (N_11964,N_11021,N_11098);
xnor U11965 (N_11965,N_11460,N_11301);
nand U11966 (N_11966,N_11285,N_11415);
or U11967 (N_11967,N_11076,N_11136);
or U11968 (N_11968,N_11393,N_11345);
xor U11969 (N_11969,N_11312,N_11408);
and U11970 (N_11970,N_11171,N_11009);
nand U11971 (N_11971,N_11347,N_11274);
nand U11972 (N_11972,N_11214,N_11283);
and U11973 (N_11973,N_11037,N_11194);
and U11974 (N_11974,N_11492,N_11231);
xnor U11975 (N_11975,N_11059,N_11494);
and U11976 (N_11976,N_11107,N_11309);
and U11977 (N_11977,N_11336,N_11105);
and U11978 (N_11978,N_11420,N_11270);
nor U11979 (N_11979,N_11298,N_11127);
nor U11980 (N_11980,N_11360,N_11018);
xnor U11981 (N_11981,N_11455,N_11399);
or U11982 (N_11982,N_11354,N_11148);
nand U11983 (N_11983,N_11333,N_11279);
nand U11984 (N_11984,N_11029,N_11432);
or U11985 (N_11985,N_11404,N_11100);
or U11986 (N_11986,N_11170,N_11027);
and U11987 (N_11987,N_11450,N_11031);
nor U11988 (N_11988,N_11083,N_11384);
and U11989 (N_11989,N_11129,N_11332);
nor U11990 (N_11990,N_11130,N_11092);
nand U11991 (N_11991,N_11059,N_11438);
nand U11992 (N_11992,N_11491,N_11068);
nand U11993 (N_11993,N_11104,N_11090);
or U11994 (N_11994,N_11078,N_11185);
and U11995 (N_11995,N_11075,N_11130);
nand U11996 (N_11996,N_11291,N_11495);
and U11997 (N_11997,N_11389,N_11044);
and U11998 (N_11998,N_11305,N_11001);
nor U11999 (N_11999,N_11496,N_11225);
nor U12000 (N_12000,N_11648,N_11957);
nand U12001 (N_12001,N_11826,N_11557);
and U12002 (N_12002,N_11909,N_11527);
nand U12003 (N_12003,N_11708,N_11522);
nor U12004 (N_12004,N_11718,N_11612);
and U12005 (N_12005,N_11928,N_11733);
or U12006 (N_12006,N_11625,N_11536);
nor U12007 (N_12007,N_11770,N_11785);
xnor U12008 (N_12008,N_11722,N_11555);
or U12009 (N_12009,N_11745,N_11933);
xor U12010 (N_12010,N_11656,N_11564);
and U12011 (N_12011,N_11758,N_11698);
nor U12012 (N_12012,N_11810,N_11788);
or U12013 (N_12013,N_11927,N_11582);
xor U12014 (N_12014,N_11679,N_11970);
or U12015 (N_12015,N_11647,N_11861);
and U12016 (N_12016,N_11998,N_11920);
nand U12017 (N_12017,N_11993,N_11595);
and U12018 (N_12018,N_11610,N_11585);
and U12019 (N_12019,N_11695,N_11895);
nand U12020 (N_12020,N_11735,N_11680);
and U12021 (N_12021,N_11523,N_11501);
xor U12022 (N_12022,N_11538,N_11635);
nor U12023 (N_12023,N_11976,N_11824);
xnor U12024 (N_12024,N_11596,N_11842);
xor U12025 (N_12025,N_11962,N_11946);
nand U12026 (N_12026,N_11864,N_11812);
and U12027 (N_12027,N_11601,N_11524);
nand U12028 (N_12028,N_11768,N_11556);
nor U12029 (N_12029,N_11593,N_11624);
xor U12030 (N_12030,N_11934,N_11863);
xor U12031 (N_12031,N_11988,N_11664);
and U12032 (N_12032,N_11742,N_11832);
nand U12033 (N_12033,N_11747,N_11953);
nor U12034 (N_12034,N_11713,N_11689);
xnor U12035 (N_12035,N_11836,N_11602);
nand U12036 (N_12036,N_11904,N_11684);
or U12037 (N_12037,N_11534,N_11749);
xnor U12038 (N_12038,N_11731,N_11549);
xor U12039 (N_12039,N_11906,N_11896);
xnor U12040 (N_12040,N_11690,N_11898);
nor U12041 (N_12041,N_11751,N_11592);
xnor U12042 (N_12042,N_11704,N_11821);
and U12043 (N_12043,N_11851,N_11677);
or U12044 (N_12044,N_11782,N_11951);
or U12045 (N_12045,N_11968,N_11702);
xnor U12046 (N_12046,N_11903,N_11880);
xor U12047 (N_12047,N_11545,N_11716);
nor U12048 (N_12048,N_11874,N_11989);
or U12049 (N_12049,N_11719,N_11741);
and U12050 (N_12050,N_11641,N_11644);
or U12051 (N_12051,N_11743,N_11889);
nand U12052 (N_12052,N_11790,N_11567);
nor U12053 (N_12053,N_11655,N_11964);
or U12054 (N_12054,N_11729,N_11653);
nand U12055 (N_12055,N_11971,N_11554);
or U12056 (N_12056,N_11779,N_11769);
nand U12057 (N_12057,N_11759,N_11579);
xnor U12058 (N_12058,N_11691,N_11587);
xor U12059 (N_12059,N_11969,N_11714);
nor U12060 (N_12060,N_11796,N_11738);
and U12061 (N_12061,N_11666,N_11526);
and U12062 (N_12062,N_11780,N_11978);
xnor U12063 (N_12063,N_11760,N_11857);
nor U12064 (N_12064,N_11723,N_11598);
and U12065 (N_12065,N_11607,N_11829);
and U12066 (N_12066,N_11703,N_11887);
nand U12067 (N_12067,N_11915,N_11816);
and U12068 (N_12068,N_11967,N_11542);
nor U12069 (N_12069,N_11809,N_11916);
and U12070 (N_12070,N_11611,N_11762);
xnor U12071 (N_12071,N_11865,N_11817);
or U12072 (N_12072,N_11930,N_11929);
nand U12073 (N_12073,N_11736,N_11616);
nand U12074 (N_12074,N_11649,N_11966);
or U12075 (N_12075,N_11855,N_11528);
xnor U12076 (N_12076,N_11603,N_11900);
or U12077 (N_12077,N_11994,N_11939);
or U12078 (N_12078,N_11921,N_11640);
or U12079 (N_12079,N_11893,N_11717);
nor U12080 (N_12080,N_11618,N_11870);
xor U12081 (N_12081,N_11529,N_11852);
and U12082 (N_12082,N_11654,N_11591);
and U12083 (N_12083,N_11778,N_11533);
xnor U12084 (N_12084,N_11725,N_11688);
nor U12085 (N_12085,N_11667,N_11755);
and U12086 (N_12086,N_11628,N_11818);
and U12087 (N_12087,N_11831,N_11833);
xnor U12088 (N_12088,N_11606,N_11958);
and U12089 (N_12089,N_11840,N_11813);
nand U12090 (N_12090,N_11776,N_11996);
nand U12091 (N_12091,N_11754,N_11795);
and U12092 (N_12092,N_11673,N_11997);
nand U12093 (N_12093,N_11558,N_11662);
and U12094 (N_12094,N_11519,N_11504);
xor U12095 (N_12095,N_11521,N_11925);
xnor U12096 (N_12096,N_11771,N_11604);
nor U12097 (N_12097,N_11746,N_11800);
or U12098 (N_12098,N_11814,N_11726);
nand U12099 (N_12099,N_11897,N_11767);
and U12100 (N_12100,N_11801,N_11634);
or U12101 (N_12101,N_11945,N_11632);
nor U12102 (N_12102,N_11869,N_11918);
or U12103 (N_12103,N_11506,N_11609);
nor U12104 (N_12104,N_11705,N_11561);
xor U12105 (N_12105,N_11982,N_11711);
nor U12106 (N_12106,N_11912,N_11845);
or U12107 (N_12107,N_11763,N_11926);
and U12108 (N_12108,N_11645,N_11671);
xnor U12109 (N_12109,N_11981,N_11669);
nand U12110 (N_12110,N_11959,N_11636);
nor U12111 (N_12111,N_11872,N_11637);
nand U12112 (N_12112,N_11961,N_11910);
nand U12113 (N_12113,N_11737,N_11622);
and U12114 (N_12114,N_11888,N_11942);
nand U12115 (N_12115,N_11772,N_11834);
and U12116 (N_12116,N_11551,N_11871);
nor U12117 (N_12117,N_11943,N_11859);
nand U12118 (N_12118,N_11570,N_11586);
and U12119 (N_12119,N_11999,N_11629);
xnor U12120 (N_12120,N_11894,N_11849);
and U12121 (N_12121,N_11513,N_11947);
or U12122 (N_12122,N_11516,N_11806);
xor U12123 (N_12123,N_11517,N_11547);
xor U12124 (N_12124,N_11908,N_11765);
or U12125 (N_12125,N_11633,N_11507);
nor U12126 (N_12126,N_11948,N_11643);
nor U12127 (N_12127,N_11919,N_11657);
nor U12128 (N_12128,N_11793,N_11709);
xor U12129 (N_12129,N_11573,N_11985);
nand U12130 (N_12130,N_11568,N_11868);
and U12131 (N_12131,N_11590,N_11546);
nand U12132 (N_12132,N_11807,N_11811);
nor U12133 (N_12133,N_11552,N_11954);
xor U12134 (N_12134,N_11562,N_11808);
nand U12135 (N_12135,N_11802,N_11797);
or U12136 (N_12136,N_11617,N_11661);
or U12137 (N_12137,N_11941,N_11581);
or U12138 (N_12138,N_11639,N_11651);
or U12139 (N_12139,N_11697,N_11505);
or U12140 (N_12140,N_11537,N_11752);
and U12141 (N_12141,N_11844,N_11949);
and U12142 (N_12142,N_11935,N_11652);
and U12143 (N_12143,N_11630,N_11975);
xnor U12144 (N_12144,N_11838,N_11509);
nand U12145 (N_12145,N_11599,N_11974);
nor U12146 (N_12146,N_11787,N_11931);
xnor U12147 (N_12147,N_11583,N_11972);
nand U12148 (N_12148,N_11907,N_11901);
and U12149 (N_12149,N_11623,N_11804);
nand U12150 (N_12150,N_11681,N_11823);
and U12151 (N_12151,N_11775,N_11525);
or U12152 (N_12152,N_11761,N_11791);
and U12153 (N_12153,N_11781,N_11531);
xor U12154 (N_12154,N_11753,N_11965);
nand U12155 (N_12155,N_11515,N_11923);
or U12156 (N_12156,N_11685,N_11952);
nand U12157 (N_12157,N_11799,N_11566);
nand U12158 (N_12158,N_11777,N_11905);
nand U12159 (N_12159,N_11783,N_11627);
xor U12160 (N_12160,N_11646,N_11827);
or U12161 (N_12161,N_11944,N_11848);
and U12162 (N_12162,N_11986,N_11532);
and U12163 (N_12163,N_11820,N_11983);
and U12164 (N_12164,N_11543,N_11580);
nand U12165 (N_12165,N_11991,N_11559);
or U12166 (N_12166,N_11854,N_11550);
or U12167 (N_12167,N_11883,N_11511);
xnor U12168 (N_12168,N_11866,N_11879);
xor U12169 (N_12169,N_11675,N_11792);
nor U12170 (N_12170,N_11589,N_11518);
or U12171 (N_12171,N_11502,N_11631);
and U12172 (N_12172,N_11950,N_11597);
nand U12173 (N_12173,N_11715,N_11835);
nand U12174 (N_12174,N_11658,N_11682);
xor U12175 (N_12175,N_11822,N_11839);
and U12176 (N_12176,N_11837,N_11500);
or U12177 (N_12177,N_11774,N_11830);
or U12178 (N_12178,N_11990,N_11608);
xnor U12179 (N_12179,N_11744,N_11825);
nor U12180 (N_12180,N_11913,N_11665);
nor U12181 (N_12181,N_11514,N_11924);
or U12182 (N_12182,N_11756,N_11572);
nand U12183 (N_12183,N_11734,N_11884);
xnor U12184 (N_12184,N_11819,N_11862);
nand U12185 (N_12185,N_11938,N_11720);
and U12186 (N_12186,N_11530,N_11815);
nor U12187 (N_12187,N_11846,N_11860);
nor U12188 (N_12188,N_11701,N_11539);
or U12189 (N_12189,N_11692,N_11541);
and U12190 (N_12190,N_11805,N_11890);
nand U12191 (N_12191,N_11902,N_11620);
xor U12192 (N_12192,N_11694,N_11892);
or U12193 (N_12193,N_11670,N_11973);
nand U12194 (N_12194,N_11732,N_11574);
nand U12195 (N_12195,N_11520,N_11987);
nor U12196 (N_12196,N_11659,N_11668);
nand U12197 (N_12197,N_11748,N_11706);
or U12198 (N_12198,N_11850,N_11563);
xor U12199 (N_12199,N_11914,N_11663);
nor U12200 (N_12200,N_11584,N_11798);
and U12201 (N_12201,N_11979,N_11876);
nor U12202 (N_12202,N_11853,N_11560);
nand U12203 (N_12203,N_11660,N_11512);
and U12204 (N_12204,N_11700,N_11642);
or U12205 (N_12205,N_11786,N_11936);
and U12206 (N_12206,N_11881,N_11984);
nand U12207 (N_12207,N_11605,N_11650);
nor U12208 (N_12208,N_11578,N_11841);
or U12209 (N_12209,N_11977,N_11956);
xor U12210 (N_12210,N_11548,N_11750);
nand U12211 (N_12211,N_11613,N_11867);
or U12212 (N_12212,N_11794,N_11594);
nor U12213 (N_12213,N_11940,N_11693);
nand U12214 (N_12214,N_11882,N_11891);
or U12215 (N_12215,N_11615,N_11687);
nor U12216 (N_12216,N_11773,N_11674);
or U12217 (N_12217,N_11764,N_11676);
nor U12218 (N_12218,N_11686,N_11877);
and U12219 (N_12219,N_11619,N_11728);
nand U12220 (N_12220,N_11721,N_11784);
nor U12221 (N_12221,N_11886,N_11995);
or U12222 (N_12222,N_11856,N_11878);
nand U12223 (N_12223,N_11739,N_11712);
nand U12224 (N_12224,N_11911,N_11540);
xor U12225 (N_12225,N_11535,N_11963);
and U12226 (N_12226,N_11955,N_11727);
nand U12227 (N_12227,N_11508,N_11696);
nor U12228 (N_12228,N_11899,N_11937);
or U12229 (N_12229,N_11510,N_11576);
nor U12230 (N_12230,N_11980,N_11992);
nand U12231 (N_12231,N_11922,N_11626);
xor U12232 (N_12232,N_11544,N_11875);
nand U12233 (N_12233,N_11699,N_11571);
xor U12234 (N_12234,N_11960,N_11724);
and U12235 (N_12235,N_11858,N_11553);
nand U12236 (N_12236,N_11757,N_11789);
nor U12237 (N_12237,N_11873,N_11503);
nand U12238 (N_12238,N_11707,N_11565);
nor U12239 (N_12239,N_11847,N_11917);
or U12240 (N_12240,N_11740,N_11843);
nand U12241 (N_12241,N_11588,N_11683);
nand U12242 (N_12242,N_11621,N_11885);
and U12243 (N_12243,N_11932,N_11577);
xor U12244 (N_12244,N_11730,N_11803);
nor U12245 (N_12245,N_11672,N_11710);
nor U12246 (N_12246,N_11575,N_11600);
nor U12247 (N_12247,N_11638,N_11828);
or U12248 (N_12248,N_11614,N_11766);
or U12249 (N_12249,N_11569,N_11678);
nand U12250 (N_12250,N_11786,N_11999);
and U12251 (N_12251,N_11936,N_11530);
xor U12252 (N_12252,N_11655,N_11760);
nand U12253 (N_12253,N_11793,N_11837);
nor U12254 (N_12254,N_11505,N_11795);
or U12255 (N_12255,N_11809,N_11871);
and U12256 (N_12256,N_11632,N_11536);
nor U12257 (N_12257,N_11906,N_11972);
nor U12258 (N_12258,N_11759,N_11744);
nor U12259 (N_12259,N_11865,N_11929);
and U12260 (N_12260,N_11519,N_11536);
or U12261 (N_12261,N_11505,N_11596);
nor U12262 (N_12262,N_11777,N_11975);
and U12263 (N_12263,N_11837,N_11729);
or U12264 (N_12264,N_11830,N_11910);
nand U12265 (N_12265,N_11796,N_11588);
xnor U12266 (N_12266,N_11735,N_11656);
nor U12267 (N_12267,N_11579,N_11952);
xnor U12268 (N_12268,N_11634,N_11727);
or U12269 (N_12269,N_11734,N_11815);
xnor U12270 (N_12270,N_11791,N_11504);
xor U12271 (N_12271,N_11779,N_11705);
xor U12272 (N_12272,N_11827,N_11585);
and U12273 (N_12273,N_11794,N_11523);
xor U12274 (N_12274,N_11577,N_11785);
and U12275 (N_12275,N_11541,N_11972);
and U12276 (N_12276,N_11791,N_11760);
xor U12277 (N_12277,N_11694,N_11936);
nor U12278 (N_12278,N_11842,N_11640);
xor U12279 (N_12279,N_11820,N_11767);
nor U12280 (N_12280,N_11519,N_11541);
nor U12281 (N_12281,N_11525,N_11740);
nand U12282 (N_12282,N_11520,N_11915);
nand U12283 (N_12283,N_11963,N_11665);
nand U12284 (N_12284,N_11722,N_11782);
nor U12285 (N_12285,N_11756,N_11784);
and U12286 (N_12286,N_11636,N_11761);
xor U12287 (N_12287,N_11782,N_11929);
nor U12288 (N_12288,N_11766,N_11916);
xnor U12289 (N_12289,N_11702,N_11996);
or U12290 (N_12290,N_11570,N_11925);
or U12291 (N_12291,N_11986,N_11502);
or U12292 (N_12292,N_11665,N_11874);
and U12293 (N_12293,N_11684,N_11950);
xnor U12294 (N_12294,N_11667,N_11512);
and U12295 (N_12295,N_11642,N_11761);
and U12296 (N_12296,N_11735,N_11553);
xor U12297 (N_12297,N_11786,N_11738);
nor U12298 (N_12298,N_11783,N_11782);
and U12299 (N_12299,N_11841,N_11549);
nor U12300 (N_12300,N_11582,N_11974);
nand U12301 (N_12301,N_11609,N_11505);
or U12302 (N_12302,N_11604,N_11853);
xnor U12303 (N_12303,N_11800,N_11714);
xor U12304 (N_12304,N_11699,N_11565);
nor U12305 (N_12305,N_11723,N_11612);
and U12306 (N_12306,N_11654,N_11593);
xor U12307 (N_12307,N_11639,N_11702);
nor U12308 (N_12308,N_11912,N_11854);
xor U12309 (N_12309,N_11712,N_11666);
or U12310 (N_12310,N_11508,N_11597);
or U12311 (N_12311,N_11500,N_11975);
or U12312 (N_12312,N_11923,N_11771);
or U12313 (N_12313,N_11695,N_11716);
xor U12314 (N_12314,N_11661,N_11614);
nand U12315 (N_12315,N_11534,N_11923);
or U12316 (N_12316,N_11522,N_11882);
nand U12317 (N_12317,N_11560,N_11722);
nor U12318 (N_12318,N_11583,N_11785);
and U12319 (N_12319,N_11627,N_11730);
or U12320 (N_12320,N_11772,N_11739);
nor U12321 (N_12321,N_11538,N_11752);
nor U12322 (N_12322,N_11608,N_11541);
nor U12323 (N_12323,N_11913,N_11683);
nor U12324 (N_12324,N_11520,N_11717);
and U12325 (N_12325,N_11904,N_11945);
xor U12326 (N_12326,N_11967,N_11528);
and U12327 (N_12327,N_11590,N_11932);
nand U12328 (N_12328,N_11645,N_11988);
or U12329 (N_12329,N_11668,N_11722);
nand U12330 (N_12330,N_11625,N_11679);
and U12331 (N_12331,N_11836,N_11891);
nor U12332 (N_12332,N_11690,N_11910);
xnor U12333 (N_12333,N_11777,N_11538);
nand U12334 (N_12334,N_11638,N_11560);
nor U12335 (N_12335,N_11644,N_11506);
xor U12336 (N_12336,N_11734,N_11567);
and U12337 (N_12337,N_11813,N_11624);
nand U12338 (N_12338,N_11596,N_11899);
or U12339 (N_12339,N_11760,N_11739);
xnor U12340 (N_12340,N_11847,N_11840);
nor U12341 (N_12341,N_11779,N_11838);
nor U12342 (N_12342,N_11900,N_11550);
or U12343 (N_12343,N_11883,N_11725);
nand U12344 (N_12344,N_11859,N_11732);
nand U12345 (N_12345,N_11649,N_11801);
or U12346 (N_12346,N_11622,N_11525);
nand U12347 (N_12347,N_11753,N_11663);
nor U12348 (N_12348,N_11702,N_11507);
and U12349 (N_12349,N_11720,N_11940);
xor U12350 (N_12350,N_11535,N_11671);
or U12351 (N_12351,N_11817,N_11600);
xnor U12352 (N_12352,N_11527,N_11676);
or U12353 (N_12353,N_11525,N_11989);
and U12354 (N_12354,N_11942,N_11553);
xor U12355 (N_12355,N_11896,N_11572);
and U12356 (N_12356,N_11558,N_11523);
xnor U12357 (N_12357,N_11520,N_11605);
nor U12358 (N_12358,N_11978,N_11854);
nor U12359 (N_12359,N_11710,N_11668);
nor U12360 (N_12360,N_11989,N_11983);
and U12361 (N_12361,N_11504,N_11988);
xor U12362 (N_12362,N_11620,N_11968);
or U12363 (N_12363,N_11549,N_11906);
and U12364 (N_12364,N_11663,N_11924);
nand U12365 (N_12365,N_11820,N_11616);
nor U12366 (N_12366,N_11776,N_11569);
or U12367 (N_12367,N_11781,N_11545);
nor U12368 (N_12368,N_11552,N_11589);
and U12369 (N_12369,N_11967,N_11631);
nand U12370 (N_12370,N_11627,N_11905);
nor U12371 (N_12371,N_11809,N_11993);
xor U12372 (N_12372,N_11940,N_11641);
xor U12373 (N_12373,N_11932,N_11848);
xor U12374 (N_12374,N_11853,N_11527);
nor U12375 (N_12375,N_11524,N_11719);
nand U12376 (N_12376,N_11521,N_11765);
or U12377 (N_12377,N_11712,N_11599);
nand U12378 (N_12378,N_11802,N_11671);
nand U12379 (N_12379,N_11602,N_11924);
and U12380 (N_12380,N_11507,N_11824);
or U12381 (N_12381,N_11610,N_11605);
nand U12382 (N_12382,N_11802,N_11639);
nor U12383 (N_12383,N_11927,N_11709);
nor U12384 (N_12384,N_11715,N_11652);
nor U12385 (N_12385,N_11543,N_11794);
nor U12386 (N_12386,N_11855,N_11813);
nand U12387 (N_12387,N_11637,N_11759);
and U12388 (N_12388,N_11795,N_11540);
xnor U12389 (N_12389,N_11661,N_11898);
nor U12390 (N_12390,N_11872,N_11997);
nor U12391 (N_12391,N_11605,N_11845);
nand U12392 (N_12392,N_11551,N_11954);
nor U12393 (N_12393,N_11714,N_11889);
xnor U12394 (N_12394,N_11938,N_11937);
nor U12395 (N_12395,N_11704,N_11544);
nor U12396 (N_12396,N_11991,N_11880);
xor U12397 (N_12397,N_11776,N_11773);
nor U12398 (N_12398,N_11845,N_11851);
xor U12399 (N_12399,N_11585,N_11975);
and U12400 (N_12400,N_11789,N_11919);
nand U12401 (N_12401,N_11996,N_11917);
nand U12402 (N_12402,N_11708,N_11969);
xor U12403 (N_12403,N_11766,N_11830);
or U12404 (N_12404,N_11735,N_11569);
nand U12405 (N_12405,N_11998,N_11518);
and U12406 (N_12406,N_11946,N_11787);
nand U12407 (N_12407,N_11586,N_11709);
or U12408 (N_12408,N_11562,N_11691);
nand U12409 (N_12409,N_11844,N_11891);
or U12410 (N_12410,N_11566,N_11722);
or U12411 (N_12411,N_11864,N_11744);
nor U12412 (N_12412,N_11775,N_11536);
and U12413 (N_12413,N_11721,N_11573);
and U12414 (N_12414,N_11523,N_11552);
nand U12415 (N_12415,N_11640,N_11562);
xnor U12416 (N_12416,N_11973,N_11987);
and U12417 (N_12417,N_11956,N_11852);
nand U12418 (N_12418,N_11900,N_11883);
or U12419 (N_12419,N_11801,N_11947);
nand U12420 (N_12420,N_11955,N_11991);
xor U12421 (N_12421,N_11641,N_11852);
xnor U12422 (N_12422,N_11660,N_11769);
or U12423 (N_12423,N_11970,N_11670);
xnor U12424 (N_12424,N_11713,N_11589);
nor U12425 (N_12425,N_11939,N_11569);
and U12426 (N_12426,N_11632,N_11970);
nor U12427 (N_12427,N_11984,N_11969);
nor U12428 (N_12428,N_11988,N_11861);
and U12429 (N_12429,N_11957,N_11753);
or U12430 (N_12430,N_11885,N_11726);
nand U12431 (N_12431,N_11748,N_11884);
or U12432 (N_12432,N_11744,N_11908);
nor U12433 (N_12433,N_11690,N_11979);
xnor U12434 (N_12434,N_11550,N_11572);
and U12435 (N_12435,N_11916,N_11583);
or U12436 (N_12436,N_11774,N_11631);
and U12437 (N_12437,N_11504,N_11837);
nor U12438 (N_12438,N_11684,N_11752);
xor U12439 (N_12439,N_11664,N_11558);
or U12440 (N_12440,N_11517,N_11965);
nor U12441 (N_12441,N_11804,N_11686);
nand U12442 (N_12442,N_11702,N_11837);
and U12443 (N_12443,N_11922,N_11673);
and U12444 (N_12444,N_11772,N_11558);
nor U12445 (N_12445,N_11607,N_11997);
or U12446 (N_12446,N_11968,N_11952);
xnor U12447 (N_12447,N_11975,N_11505);
nand U12448 (N_12448,N_11502,N_11549);
xnor U12449 (N_12449,N_11866,N_11997);
nand U12450 (N_12450,N_11982,N_11725);
nand U12451 (N_12451,N_11548,N_11607);
nor U12452 (N_12452,N_11757,N_11873);
and U12453 (N_12453,N_11947,N_11826);
and U12454 (N_12454,N_11808,N_11572);
or U12455 (N_12455,N_11794,N_11966);
and U12456 (N_12456,N_11526,N_11767);
and U12457 (N_12457,N_11914,N_11744);
nand U12458 (N_12458,N_11708,N_11812);
xor U12459 (N_12459,N_11823,N_11792);
xnor U12460 (N_12460,N_11520,N_11999);
nand U12461 (N_12461,N_11501,N_11736);
or U12462 (N_12462,N_11820,N_11528);
and U12463 (N_12463,N_11716,N_11553);
and U12464 (N_12464,N_11909,N_11812);
and U12465 (N_12465,N_11905,N_11801);
nor U12466 (N_12466,N_11704,N_11877);
nor U12467 (N_12467,N_11612,N_11757);
or U12468 (N_12468,N_11763,N_11980);
nand U12469 (N_12469,N_11621,N_11725);
or U12470 (N_12470,N_11820,N_11912);
nor U12471 (N_12471,N_11554,N_11791);
nor U12472 (N_12472,N_11764,N_11634);
nor U12473 (N_12473,N_11621,N_11580);
and U12474 (N_12474,N_11707,N_11860);
nand U12475 (N_12475,N_11852,N_11822);
nor U12476 (N_12476,N_11668,N_11919);
or U12477 (N_12477,N_11786,N_11570);
nor U12478 (N_12478,N_11864,N_11641);
nand U12479 (N_12479,N_11667,N_11761);
and U12480 (N_12480,N_11591,N_11949);
xnor U12481 (N_12481,N_11576,N_11678);
or U12482 (N_12482,N_11587,N_11553);
and U12483 (N_12483,N_11734,N_11964);
xor U12484 (N_12484,N_11907,N_11591);
and U12485 (N_12485,N_11850,N_11962);
nand U12486 (N_12486,N_11803,N_11649);
nor U12487 (N_12487,N_11649,N_11845);
xor U12488 (N_12488,N_11555,N_11692);
xor U12489 (N_12489,N_11641,N_11674);
xnor U12490 (N_12490,N_11747,N_11933);
nand U12491 (N_12491,N_11588,N_11913);
nor U12492 (N_12492,N_11579,N_11563);
xor U12493 (N_12493,N_11826,N_11610);
or U12494 (N_12494,N_11987,N_11734);
or U12495 (N_12495,N_11947,N_11528);
nand U12496 (N_12496,N_11506,N_11867);
nor U12497 (N_12497,N_11650,N_11915);
nor U12498 (N_12498,N_11604,N_11538);
and U12499 (N_12499,N_11753,N_11650);
or U12500 (N_12500,N_12434,N_12040);
or U12501 (N_12501,N_12090,N_12102);
xnor U12502 (N_12502,N_12124,N_12180);
nor U12503 (N_12503,N_12373,N_12261);
or U12504 (N_12504,N_12156,N_12143);
and U12505 (N_12505,N_12224,N_12227);
nor U12506 (N_12506,N_12200,N_12312);
nand U12507 (N_12507,N_12053,N_12086);
nand U12508 (N_12508,N_12093,N_12175);
or U12509 (N_12509,N_12337,N_12234);
or U12510 (N_12510,N_12308,N_12207);
and U12511 (N_12511,N_12095,N_12364);
xor U12512 (N_12512,N_12411,N_12088);
and U12513 (N_12513,N_12316,N_12451);
xor U12514 (N_12514,N_12442,N_12035);
and U12515 (N_12515,N_12340,N_12357);
or U12516 (N_12516,N_12375,N_12245);
xnor U12517 (N_12517,N_12336,N_12267);
and U12518 (N_12518,N_12128,N_12454);
and U12519 (N_12519,N_12286,N_12477);
xor U12520 (N_12520,N_12145,N_12325);
or U12521 (N_12521,N_12445,N_12055);
and U12522 (N_12522,N_12253,N_12169);
and U12523 (N_12523,N_12238,N_12423);
or U12524 (N_12524,N_12222,N_12413);
xor U12525 (N_12525,N_12172,N_12057);
nor U12526 (N_12526,N_12187,N_12473);
nand U12527 (N_12527,N_12008,N_12030);
and U12528 (N_12528,N_12044,N_12258);
nor U12529 (N_12529,N_12070,N_12060);
nor U12530 (N_12530,N_12367,N_12067);
and U12531 (N_12531,N_12161,N_12191);
xnor U12532 (N_12532,N_12186,N_12241);
and U12533 (N_12533,N_12299,N_12075);
and U12534 (N_12534,N_12420,N_12449);
xnor U12535 (N_12535,N_12452,N_12397);
or U12536 (N_12536,N_12059,N_12016);
and U12537 (N_12537,N_12365,N_12369);
xor U12538 (N_12538,N_12013,N_12487);
nor U12539 (N_12539,N_12135,N_12460);
or U12540 (N_12540,N_12289,N_12327);
or U12541 (N_12541,N_12326,N_12358);
nand U12542 (N_12542,N_12081,N_12098);
xnor U12543 (N_12543,N_12160,N_12492);
and U12544 (N_12544,N_12415,N_12381);
or U12545 (N_12545,N_12430,N_12361);
nand U12546 (N_12546,N_12484,N_12437);
nand U12547 (N_12547,N_12348,N_12260);
nor U12548 (N_12548,N_12097,N_12400);
and U12549 (N_12549,N_12268,N_12343);
and U12550 (N_12550,N_12410,N_12403);
nand U12551 (N_12551,N_12422,N_12331);
or U12552 (N_12552,N_12388,N_12465);
nor U12553 (N_12553,N_12290,N_12396);
or U12554 (N_12554,N_12401,N_12197);
xor U12555 (N_12555,N_12063,N_12134);
nor U12556 (N_12556,N_12279,N_12037);
or U12557 (N_12557,N_12250,N_12363);
nor U12558 (N_12558,N_12265,N_12303);
nor U12559 (N_12559,N_12116,N_12025);
xor U12560 (N_12560,N_12237,N_12483);
nand U12561 (N_12561,N_12017,N_12216);
xnor U12562 (N_12562,N_12269,N_12402);
nor U12563 (N_12563,N_12218,N_12007);
nor U12564 (N_12564,N_12189,N_12009);
and U12565 (N_12565,N_12125,N_12391);
and U12566 (N_12566,N_12287,N_12211);
nand U12567 (N_12567,N_12352,N_12166);
nand U12568 (N_12568,N_12313,N_12271);
or U12569 (N_12569,N_12274,N_12421);
and U12570 (N_12570,N_12165,N_12104);
or U12571 (N_12571,N_12203,N_12426);
and U12572 (N_12572,N_12469,N_12467);
xnor U12573 (N_12573,N_12333,N_12111);
or U12574 (N_12574,N_12459,N_12176);
nor U12575 (N_12575,N_12285,N_12006);
or U12576 (N_12576,N_12428,N_12170);
nor U12577 (N_12577,N_12223,N_12201);
or U12578 (N_12578,N_12468,N_12034);
and U12579 (N_12579,N_12498,N_12408);
xor U12580 (N_12580,N_12295,N_12202);
xnor U12581 (N_12581,N_12371,N_12491);
or U12582 (N_12582,N_12392,N_12153);
or U12583 (N_12583,N_12259,N_12168);
and U12584 (N_12584,N_12228,N_12334);
and U12585 (N_12585,N_12076,N_12215);
xnor U12586 (N_12586,N_12406,N_12378);
and U12587 (N_12587,N_12366,N_12107);
nor U12588 (N_12588,N_12329,N_12475);
nand U12589 (N_12589,N_12001,N_12317);
and U12590 (N_12590,N_12123,N_12085);
nor U12591 (N_12591,N_12418,N_12065);
nand U12592 (N_12592,N_12069,N_12433);
and U12593 (N_12593,N_12139,N_12281);
or U12594 (N_12594,N_12319,N_12014);
nand U12595 (N_12595,N_12003,N_12417);
nor U12596 (N_12596,N_12026,N_12306);
nor U12597 (N_12597,N_12345,N_12082);
and U12598 (N_12598,N_12377,N_12077);
nand U12599 (N_12599,N_12115,N_12210);
and U12600 (N_12600,N_12004,N_12328);
or U12601 (N_12601,N_12324,N_12194);
or U12602 (N_12602,N_12476,N_12414);
and U12603 (N_12603,N_12471,N_12015);
or U12604 (N_12604,N_12213,N_12072);
xnor U12605 (N_12605,N_12248,N_12438);
and U12606 (N_12606,N_12087,N_12174);
xnor U12607 (N_12607,N_12036,N_12399);
nand U12608 (N_12608,N_12021,N_12141);
nand U12609 (N_12609,N_12243,N_12046);
or U12610 (N_12610,N_12150,N_12131);
nor U12611 (N_12611,N_12395,N_12344);
or U12612 (N_12612,N_12031,N_12148);
nand U12613 (N_12613,N_12188,N_12379);
or U12614 (N_12614,N_12239,N_12220);
xor U12615 (N_12615,N_12011,N_12270);
or U12616 (N_12616,N_12380,N_12184);
nand U12617 (N_12617,N_12350,N_12185);
or U12618 (N_12618,N_12023,N_12493);
xor U12619 (N_12619,N_12162,N_12480);
nand U12620 (N_12620,N_12167,N_12485);
nand U12621 (N_12621,N_12390,N_12440);
or U12622 (N_12622,N_12394,N_12419);
and U12623 (N_12623,N_12147,N_12386);
nor U12624 (N_12624,N_12398,N_12109);
nor U12625 (N_12625,N_12142,N_12425);
nand U12626 (N_12626,N_12120,N_12198);
nand U12627 (N_12627,N_12293,N_12221);
or U12628 (N_12628,N_12355,N_12119);
nand U12629 (N_12629,N_12264,N_12024);
xor U12630 (N_12630,N_12252,N_12247);
nand U12631 (N_12631,N_12195,N_12246);
nor U12632 (N_12632,N_12441,N_12443);
nor U12633 (N_12633,N_12209,N_12226);
xor U12634 (N_12634,N_12049,N_12351);
or U12635 (N_12635,N_12231,N_12407);
xor U12636 (N_12636,N_12229,N_12219);
or U12637 (N_12637,N_12137,N_12262);
and U12638 (N_12638,N_12474,N_12310);
nor U12639 (N_12639,N_12133,N_12020);
nor U12640 (N_12640,N_12117,N_12298);
nand U12641 (N_12641,N_12458,N_12453);
or U12642 (N_12642,N_12305,N_12178);
and U12643 (N_12643,N_12108,N_12318);
nor U12644 (N_12644,N_12029,N_12382);
nor U12645 (N_12645,N_12457,N_12214);
and U12646 (N_12646,N_12126,N_12225);
nand U12647 (N_12647,N_12047,N_12463);
or U12648 (N_12648,N_12376,N_12446);
nand U12649 (N_12649,N_12296,N_12416);
xnor U12650 (N_12650,N_12064,N_12118);
or U12651 (N_12651,N_12335,N_12022);
and U12652 (N_12652,N_12179,N_12230);
nand U12653 (N_12653,N_12456,N_12050);
nand U12654 (N_12654,N_12196,N_12190);
nor U12655 (N_12655,N_12436,N_12347);
and U12656 (N_12656,N_12482,N_12464);
nand U12657 (N_12657,N_12101,N_12346);
or U12658 (N_12658,N_12112,N_12322);
xor U12659 (N_12659,N_12010,N_12171);
nor U12660 (N_12660,N_12283,N_12342);
and U12661 (N_12661,N_12041,N_12429);
or U12662 (N_12662,N_12164,N_12106);
nand U12663 (N_12663,N_12100,N_12462);
nor U12664 (N_12664,N_12489,N_12018);
nor U12665 (N_12665,N_12113,N_12360);
nor U12666 (N_12666,N_12027,N_12159);
nor U12667 (N_12667,N_12424,N_12000);
and U12668 (N_12668,N_12320,N_12256);
xor U12669 (N_12669,N_12080,N_12277);
nor U12670 (N_12670,N_12494,N_12275);
nor U12671 (N_12671,N_12078,N_12193);
or U12672 (N_12672,N_12431,N_12490);
xor U12673 (N_12673,N_12192,N_12300);
nand U12674 (N_12674,N_12427,N_12254);
nor U12675 (N_12675,N_12033,N_12478);
nand U12676 (N_12676,N_12122,N_12071);
nand U12677 (N_12677,N_12461,N_12497);
xor U12678 (N_12678,N_12005,N_12039);
xor U12679 (N_12679,N_12311,N_12199);
or U12680 (N_12680,N_12301,N_12091);
and U12681 (N_12681,N_12205,N_12276);
or U12682 (N_12682,N_12472,N_12404);
xor U12683 (N_12683,N_12292,N_12136);
and U12684 (N_12684,N_12302,N_12177);
nor U12685 (N_12685,N_12251,N_12099);
nand U12686 (N_12686,N_12496,N_12393);
and U12687 (N_12687,N_12240,N_12129);
nor U12688 (N_12688,N_12045,N_12309);
nand U12689 (N_12689,N_12321,N_12233);
nand U12690 (N_12690,N_12151,N_12096);
xnor U12691 (N_12691,N_12236,N_12249);
or U12692 (N_12692,N_12499,N_12323);
and U12693 (N_12693,N_12356,N_12110);
and U12694 (N_12694,N_12084,N_12232);
xor U12695 (N_12695,N_12466,N_12288);
nand U12696 (N_12696,N_12354,N_12470);
nor U12697 (N_12697,N_12448,N_12315);
nor U12698 (N_12698,N_12019,N_12447);
nor U12699 (N_12699,N_12217,N_12073);
xnor U12700 (N_12700,N_12444,N_12338);
xor U12701 (N_12701,N_12304,N_12042);
and U12702 (N_12702,N_12486,N_12173);
or U12703 (N_12703,N_12012,N_12146);
nand U12704 (N_12704,N_12121,N_12183);
nand U12705 (N_12705,N_12370,N_12092);
or U12706 (N_12706,N_12114,N_12389);
xor U12707 (N_12707,N_12479,N_12127);
nor U12708 (N_12708,N_12181,N_12158);
nor U12709 (N_12709,N_12054,N_12103);
nand U12710 (N_12710,N_12038,N_12481);
xnor U12711 (N_12711,N_12330,N_12495);
nand U12712 (N_12712,N_12272,N_12341);
or U12713 (N_12713,N_12435,N_12383);
nand U12714 (N_12714,N_12307,N_12032);
nor U12715 (N_12715,N_12349,N_12079);
or U12716 (N_12716,N_12157,N_12314);
xnor U12717 (N_12717,N_12359,N_12144);
xor U12718 (N_12718,N_12339,N_12094);
nand U12719 (N_12719,N_12273,N_12332);
nand U12720 (N_12720,N_12152,N_12488);
nor U12721 (N_12721,N_12409,N_12294);
nor U12722 (N_12722,N_12242,N_12291);
nor U12723 (N_12723,N_12130,N_12208);
xor U12724 (N_12724,N_12450,N_12455);
xnor U12725 (N_12725,N_12385,N_12282);
nor U12726 (N_12726,N_12235,N_12255);
or U12727 (N_12727,N_12263,N_12083);
nand U12728 (N_12728,N_12138,N_12056);
nor U12729 (N_12729,N_12182,N_12432);
and U12730 (N_12730,N_12002,N_12074);
nand U12731 (N_12731,N_12140,N_12163);
or U12732 (N_12732,N_12058,N_12068);
nor U12733 (N_12733,N_12374,N_12155);
nand U12734 (N_12734,N_12439,N_12052);
and U12735 (N_12735,N_12405,N_12353);
or U12736 (N_12736,N_12154,N_12278);
and U12737 (N_12737,N_12048,N_12297);
and U12738 (N_12738,N_12061,N_12412);
nand U12739 (N_12739,N_12280,N_12028);
and U12740 (N_12740,N_12105,N_12387);
and U12741 (N_12741,N_12368,N_12266);
xnor U12742 (N_12742,N_12204,N_12362);
nand U12743 (N_12743,N_12051,N_12206);
or U12744 (N_12744,N_12257,N_12066);
xor U12745 (N_12745,N_12132,N_12244);
and U12746 (N_12746,N_12089,N_12062);
or U12747 (N_12747,N_12149,N_12212);
xnor U12748 (N_12748,N_12384,N_12372);
nor U12749 (N_12749,N_12043,N_12284);
xnor U12750 (N_12750,N_12006,N_12342);
or U12751 (N_12751,N_12131,N_12077);
nor U12752 (N_12752,N_12309,N_12287);
nor U12753 (N_12753,N_12104,N_12289);
xor U12754 (N_12754,N_12462,N_12429);
nor U12755 (N_12755,N_12111,N_12324);
nand U12756 (N_12756,N_12079,N_12302);
nand U12757 (N_12757,N_12004,N_12210);
nand U12758 (N_12758,N_12410,N_12482);
or U12759 (N_12759,N_12269,N_12321);
or U12760 (N_12760,N_12491,N_12338);
xor U12761 (N_12761,N_12127,N_12261);
and U12762 (N_12762,N_12079,N_12142);
or U12763 (N_12763,N_12143,N_12379);
nor U12764 (N_12764,N_12092,N_12148);
nor U12765 (N_12765,N_12245,N_12247);
xnor U12766 (N_12766,N_12175,N_12329);
nor U12767 (N_12767,N_12211,N_12408);
or U12768 (N_12768,N_12022,N_12113);
nor U12769 (N_12769,N_12265,N_12165);
nand U12770 (N_12770,N_12278,N_12426);
xnor U12771 (N_12771,N_12367,N_12469);
xnor U12772 (N_12772,N_12364,N_12111);
nor U12773 (N_12773,N_12194,N_12343);
nand U12774 (N_12774,N_12413,N_12329);
or U12775 (N_12775,N_12349,N_12017);
nand U12776 (N_12776,N_12456,N_12281);
and U12777 (N_12777,N_12332,N_12159);
and U12778 (N_12778,N_12266,N_12354);
nand U12779 (N_12779,N_12486,N_12076);
nand U12780 (N_12780,N_12252,N_12494);
nor U12781 (N_12781,N_12167,N_12349);
nor U12782 (N_12782,N_12424,N_12279);
nor U12783 (N_12783,N_12407,N_12441);
nand U12784 (N_12784,N_12197,N_12268);
nor U12785 (N_12785,N_12379,N_12344);
nand U12786 (N_12786,N_12160,N_12176);
and U12787 (N_12787,N_12144,N_12198);
xnor U12788 (N_12788,N_12135,N_12330);
xor U12789 (N_12789,N_12075,N_12113);
and U12790 (N_12790,N_12078,N_12320);
and U12791 (N_12791,N_12118,N_12448);
xnor U12792 (N_12792,N_12060,N_12105);
xor U12793 (N_12793,N_12187,N_12270);
and U12794 (N_12794,N_12334,N_12365);
nor U12795 (N_12795,N_12437,N_12315);
nor U12796 (N_12796,N_12085,N_12094);
nand U12797 (N_12797,N_12025,N_12217);
nand U12798 (N_12798,N_12286,N_12292);
nand U12799 (N_12799,N_12194,N_12013);
xnor U12800 (N_12800,N_12036,N_12126);
xnor U12801 (N_12801,N_12338,N_12289);
nand U12802 (N_12802,N_12361,N_12180);
nor U12803 (N_12803,N_12271,N_12155);
or U12804 (N_12804,N_12478,N_12401);
nand U12805 (N_12805,N_12162,N_12377);
and U12806 (N_12806,N_12127,N_12109);
nand U12807 (N_12807,N_12484,N_12478);
xnor U12808 (N_12808,N_12181,N_12381);
and U12809 (N_12809,N_12187,N_12330);
and U12810 (N_12810,N_12189,N_12039);
xnor U12811 (N_12811,N_12275,N_12243);
xor U12812 (N_12812,N_12146,N_12161);
or U12813 (N_12813,N_12176,N_12114);
nor U12814 (N_12814,N_12322,N_12422);
nand U12815 (N_12815,N_12308,N_12350);
nand U12816 (N_12816,N_12346,N_12259);
and U12817 (N_12817,N_12473,N_12013);
or U12818 (N_12818,N_12089,N_12479);
nand U12819 (N_12819,N_12035,N_12070);
nand U12820 (N_12820,N_12285,N_12409);
nand U12821 (N_12821,N_12463,N_12281);
and U12822 (N_12822,N_12152,N_12036);
or U12823 (N_12823,N_12207,N_12172);
nand U12824 (N_12824,N_12203,N_12000);
nand U12825 (N_12825,N_12435,N_12409);
xor U12826 (N_12826,N_12209,N_12046);
and U12827 (N_12827,N_12387,N_12285);
and U12828 (N_12828,N_12304,N_12001);
or U12829 (N_12829,N_12290,N_12047);
nor U12830 (N_12830,N_12429,N_12078);
or U12831 (N_12831,N_12310,N_12171);
nand U12832 (N_12832,N_12202,N_12197);
and U12833 (N_12833,N_12098,N_12200);
xor U12834 (N_12834,N_12232,N_12238);
nor U12835 (N_12835,N_12067,N_12200);
nand U12836 (N_12836,N_12091,N_12049);
nor U12837 (N_12837,N_12003,N_12028);
xnor U12838 (N_12838,N_12229,N_12158);
or U12839 (N_12839,N_12176,N_12434);
nand U12840 (N_12840,N_12379,N_12019);
and U12841 (N_12841,N_12439,N_12016);
or U12842 (N_12842,N_12244,N_12156);
or U12843 (N_12843,N_12130,N_12349);
xor U12844 (N_12844,N_12107,N_12387);
xor U12845 (N_12845,N_12485,N_12453);
xor U12846 (N_12846,N_12197,N_12199);
and U12847 (N_12847,N_12474,N_12422);
and U12848 (N_12848,N_12301,N_12112);
nand U12849 (N_12849,N_12025,N_12449);
xor U12850 (N_12850,N_12064,N_12215);
nand U12851 (N_12851,N_12266,N_12480);
or U12852 (N_12852,N_12231,N_12326);
xor U12853 (N_12853,N_12476,N_12060);
or U12854 (N_12854,N_12135,N_12152);
or U12855 (N_12855,N_12469,N_12176);
nor U12856 (N_12856,N_12444,N_12188);
nand U12857 (N_12857,N_12424,N_12467);
nand U12858 (N_12858,N_12027,N_12290);
and U12859 (N_12859,N_12108,N_12163);
nand U12860 (N_12860,N_12428,N_12265);
or U12861 (N_12861,N_12169,N_12192);
xnor U12862 (N_12862,N_12309,N_12311);
xor U12863 (N_12863,N_12175,N_12145);
and U12864 (N_12864,N_12115,N_12098);
or U12865 (N_12865,N_12295,N_12189);
xor U12866 (N_12866,N_12236,N_12348);
nor U12867 (N_12867,N_12176,N_12375);
or U12868 (N_12868,N_12453,N_12168);
nor U12869 (N_12869,N_12402,N_12452);
nand U12870 (N_12870,N_12349,N_12208);
nor U12871 (N_12871,N_12440,N_12008);
nor U12872 (N_12872,N_12487,N_12498);
and U12873 (N_12873,N_12433,N_12333);
and U12874 (N_12874,N_12141,N_12348);
and U12875 (N_12875,N_12259,N_12108);
nand U12876 (N_12876,N_12234,N_12387);
nor U12877 (N_12877,N_12373,N_12262);
nand U12878 (N_12878,N_12245,N_12099);
xnor U12879 (N_12879,N_12183,N_12487);
and U12880 (N_12880,N_12006,N_12002);
nand U12881 (N_12881,N_12125,N_12034);
nor U12882 (N_12882,N_12429,N_12319);
xnor U12883 (N_12883,N_12447,N_12337);
and U12884 (N_12884,N_12172,N_12378);
and U12885 (N_12885,N_12100,N_12107);
xor U12886 (N_12886,N_12190,N_12311);
xor U12887 (N_12887,N_12226,N_12218);
xnor U12888 (N_12888,N_12470,N_12264);
and U12889 (N_12889,N_12137,N_12354);
and U12890 (N_12890,N_12076,N_12352);
or U12891 (N_12891,N_12012,N_12389);
xnor U12892 (N_12892,N_12054,N_12196);
nor U12893 (N_12893,N_12236,N_12083);
and U12894 (N_12894,N_12063,N_12451);
or U12895 (N_12895,N_12425,N_12375);
xor U12896 (N_12896,N_12214,N_12305);
and U12897 (N_12897,N_12310,N_12279);
or U12898 (N_12898,N_12131,N_12382);
nor U12899 (N_12899,N_12145,N_12334);
or U12900 (N_12900,N_12188,N_12309);
xor U12901 (N_12901,N_12217,N_12277);
xor U12902 (N_12902,N_12378,N_12421);
nand U12903 (N_12903,N_12055,N_12019);
nor U12904 (N_12904,N_12224,N_12035);
and U12905 (N_12905,N_12459,N_12062);
and U12906 (N_12906,N_12391,N_12405);
and U12907 (N_12907,N_12234,N_12351);
nand U12908 (N_12908,N_12120,N_12481);
or U12909 (N_12909,N_12321,N_12122);
nor U12910 (N_12910,N_12224,N_12484);
and U12911 (N_12911,N_12372,N_12277);
xor U12912 (N_12912,N_12387,N_12141);
nand U12913 (N_12913,N_12258,N_12055);
nand U12914 (N_12914,N_12028,N_12187);
and U12915 (N_12915,N_12425,N_12018);
nand U12916 (N_12916,N_12289,N_12056);
nor U12917 (N_12917,N_12302,N_12136);
and U12918 (N_12918,N_12160,N_12088);
nor U12919 (N_12919,N_12244,N_12160);
or U12920 (N_12920,N_12016,N_12122);
nor U12921 (N_12921,N_12219,N_12463);
nor U12922 (N_12922,N_12435,N_12050);
nor U12923 (N_12923,N_12192,N_12084);
xnor U12924 (N_12924,N_12144,N_12042);
xor U12925 (N_12925,N_12254,N_12326);
xnor U12926 (N_12926,N_12033,N_12373);
or U12927 (N_12927,N_12293,N_12342);
nor U12928 (N_12928,N_12251,N_12010);
nor U12929 (N_12929,N_12234,N_12202);
or U12930 (N_12930,N_12184,N_12080);
or U12931 (N_12931,N_12314,N_12404);
and U12932 (N_12932,N_12363,N_12322);
nand U12933 (N_12933,N_12430,N_12224);
and U12934 (N_12934,N_12192,N_12210);
nand U12935 (N_12935,N_12381,N_12444);
and U12936 (N_12936,N_12209,N_12112);
and U12937 (N_12937,N_12118,N_12180);
and U12938 (N_12938,N_12363,N_12494);
or U12939 (N_12939,N_12164,N_12051);
and U12940 (N_12940,N_12149,N_12155);
nand U12941 (N_12941,N_12294,N_12139);
nand U12942 (N_12942,N_12327,N_12374);
nand U12943 (N_12943,N_12359,N_12196);
nor U12944 (N_12944,N_12045,N_12163);
and U12945 (N_12945,N_12149,N_12420);
and U12946 (N_12946,N_12361,N_12202);
or U12947 (N_12947,N_12381,N_12476);
nor U12948 (N_12948,N_12231,N_12441);
nor U12949 (N_12949,N_12341,N_12015);
xnor U12950 (N_12950,N_12300,N_12379);
xnor U12951 (N_12951,N_12267,N_12209);
and U12952 (N_12952,N_12206,N_12417);
and U12953 (N_12953,N_12242,N_12129);
nand U12954 (N_12954,N_12029,N_12191);
nor U12955 (N_12955,N_12497,N_12186);
or U12956 (N_12956,N_12402,N_12482);
or U12957 (N_12957,N_12221,N_12213);
nand U12958 (N_12958,N_12142,N_12454);
or U12959 (N_12959,N_12375,N_12262);
nand U12960 (N_12960,N_12126,N_12390);
or U12961 (N_12961,N_12360,N_12354);
or U12962 (N_12962,N_12350,N_12196);
and U12963 (N_12963,N_12129,N_12259);
and U12964 (N_12964,N_12130,N_12216);
xnor U12965 (N_12965,N_12025,N_12032);
xor U12966 (N_12966,N_12416,N_12468);
or U12967 (N_12967,N_12211,N_12112);
and U12968 (N_12968,N_12204,N_12234);
nor U12969 (N_12969,N_12432,N_12174);
or U12970 (N_12970,N_12468,N_12328);
and U12971 (N_12971,N_12439,N_12028);
xor U12972 (N_12972,N_12276,N_12469);
xor U12973 (N_12973,N_12062,N_12434);
and U12974 (N_12974,N_12484,N_12090);
nor U12975 (N_12975,N_12262,N_12049);
nor U12976 (N_12976,N_12442,N_12211);
nor U12977 (N_12977,N_12385,N_12052);
nand U12978 (N_12978,N_12492,N_12152);
and U12979 (N_12979,N_12016,N_12376);
or U12980 (N_12980,N_12253,N_12220);
or U12981 (N_12981,N_12402,N_12253);
xor U12982 (N_12982,N_12251,N_12309);
and U12983 (N_12983,N_12465,N_12223);
nor U12984 (N_12984,N_12482,N_12458);
xnor U12985 (N_12985,N_12344,N_12405);
and U12986 (N_12986,N_12036,N_12013);
and U12987 (N_12987,N_12047,N_12124);
nor U12988 (N_12988,N_12454,N_12171);
nor U12989 (N_12989,N_12497,N_12457);
or U12990 (N_12990,N_12201,N_12258);
nand U12991 (N_12991,N_12266,N_12248);
and U12992 (N_12992,N_12392,N_12036);
nand U12993 (N_12993,N_12164,N_12028);
or U12994 (N_12994,N_12105,N_12146);
xnor U12995 (N_12995,N_12245,N_12170);
xor U12996 (N_12996,N_12120,N_12204);
nor U12997 (N_12997,N_12328,N_12219);
and U12998 (N_12998,N_12167,N_12392);
xnor U12999 (N_12999,N_12101,N_12212);
or U13000 (N_13000,N_12658,N_12518);
and U13001 (N_13001,N_12997,N_12561);
nand U13002 (N_13002,N_12522,N_12749);
and U13003 (N_13003,N_12849,N_12770);
and U13004 (N_13004,N_12787,N_12694);
nor U13005 (N_13005,N_12819,N_12808);
xor U13006 (N_13006,N_12864,N_12925);
and U13007 (N_13007,N_12521,N_12769);
nor U13008 (N_13008,N_12806,N_12569);
nand U13009 (N_13009,N_12580,N_12516);
and U13010 (N_13010,N_12993,N_12554);
nand U13011 (N_13011,N_12761,N_12861);
nand U13012 (N_13012,N_12591,N_12739);
and U13013 (N_13013,N_12870,N_12623);
nand U13014 (N_13014,N_12840,N_12824);
xor U13015 (N_13015,N_12717,N_12735);
or U13016 (N_13016,N_12611,N_12600);
nor U13017 (N_13017,N_12729,N_12541);
xor U13018 (N_13018,N_12816,N_12697);
or U13019 (N_13019,N_12539,N_12567);
nand U13020 (N_13020,N_12989,N_12716);
or U13021 (N_13021,N_12983,N_12682);
nand U13022 (N_13022,N_12594,N_12820);
or U13023 (N_13023,N_12990,N_12556);
and U13024 (N_13024,N_12551,N_12626);
or U13025 (N_13025,N_12933,N_12951);
and U13026 (N_13026,N_12771,N_12899);
xnor U13027 (N_13027,N_12982,N_12785);
xnor U13028 (N_13028,N_12721,N_12609);
nand U13029 (N_13029,N_12636,N_12776);
xnor U13030 (N_13030,N_12766,N_12881);
or U13031 (N_13031,N_12693,N_12695);
nor U13032 (N_13032,N_12774,N_12577);
and U13033 (N_13033,N_12805,N_12913);
xor U13034 (N_13034,N_12760,N_12773);
xor U13035 (N_13035,N_12886,N_12862);
or U13036 (N_13036,N_12812,N_12972);
xnor U13037 (N_13037,N_12730,N_12944);
or U13038 (N_13038,N_12617,N_12542);
nand U13039 (N_13039,N_12880,N_12549);
nor U13040 (N_13040,N_12723,N_12905);
nand U13041 (N_13041,N_12875,N_12509);
xor U13042 (N_13042,N_12839,N_12614);
and U13043 (N_13043,N_12882,N_12830);
and U13044 (N_13044,N_12575,N_12651);
or U13045 (N_13045,N_12559,N_12775);
and U13046 (N_13046,N_12573,N_12916);
xor U13047 (N_13047,N_12827,N_12911);
nor U13048 (N_13048,N_12991,N_12878);
or U13049 (N_13049,N_12943,N_12505);
nand U13050 (N_13050,N_12858,N_12663);
nor U13051 (N_13051,N_12980,N_12713);
nor U13052 (N_13052,N_12534,N_12842);
nor U13053 (N_13053,N_12999,N_12520);
nand U13054 (N_13054,N_12587,N_12714);
xnor U13055 (N_13055,N_12736,N_12897);
and U13056 (N_13056,N_12867,N_12907);
xnor U13057 (N_13057,N_12523,N_12524);
nor U13058 (N_13058,N_12928,N_12590);
or U13059 (N_13059,N_12866,N_12803);
or U13060 (N_13060,N_12596,N_12661);
or U13061 (N_13061,N_12822,N_12601);
and U13062 (N_13062,N_12583,N_12715);
nand U13063 (N_13063,N_12654,N_12865);
xor U13064 (N_13064,N_12818,N_12835);
xnor U13065 (N_13065,N_12696,N_12826);
nor U13066 (N_13066,N_12637,N_12552);
nand U13067 (N_13067,N_12526,N_12562);
or U13068 (N_13068,N_12978,N_12646);
nor U13069 (N_13069,N_12846,N_12817);
xor U13070 (N_13070,N_12672,N_12802);
nand U13071 (N_13071,N_12550,N_12533);
nor U13072 (N_13072,N_12958,N_12709);
nor U13073 (N_13073,N_12710,N_12772);
and U13074 (N_13074,N_12706,N_12588);
xor U13075 (N_13075,N_12678,N_12922);
xnor U13076 (N_13076,N_12843,N_12608);
or U13077 (N_13077,N_12926,N_12939);
nand U13078 (N_13078,N_12954,N_12506);
and U13079 (N_13079,N_12645,N_12790);
or U13080 (N_13080,N_12971,N_12643);
nor U13081 (N_13081,N_12572,N_12893);
nand U13082 (N_13082,N_12571,N_12987);
and U13083 (N_13083,N_12889,N_12703);
or U13084 (N_13084,N_12935,N_12619);
or U13085 (N_13085,N_12797,N_12850);
and U13086 (N_13086,N_12968,N_12622);
nand U13087 (N_13087,N_12679,N_12910);
xor U13088 (N_13088,N_12758,N_12894);
xor U13089 (N_13089,N_12756,N_12791);
nand U13090 (N_13090,N_12833,N_12501);
or U13091 (N_13091,N_12847,N_12921);
and U13092 (N_13092,N_12510,N_12517);
and U13093 (N_13093,N_12976,N_12741);
and U13094 (N_13094,N_12931,N_12664);
nand U13095 (N_13095,N_12531,N_12720);
or U13096 (N_13096,N_12656,N_12754);
xnor U13097 (N_13097,N_12837,N_12814);
or U13098 (N_13098,N_12854,N_12964);
xnor U13099 (N_13099,N_12634,N_12667);
nand U13100 (N_13100,N_12879,N_12547);
nand U13101 (N_13101,N_12915,N_12638);
xor U13102 (N_13102,N_12901,N_12900);
nor U13103 (N_13103,N_12669,N_12918);
nand U13104 (N_13104,N_12599,N_12810);
nand U13105 (N_13105,N_12869,N_12759);
or U13106 (N_13106,N_12952,N_12597);
xor U13107 (N_13107,N_12752,N_12724);
xor U13108 (N_13108,N_12793,N_12668);
nand U13109 (N_13109,N_12613,N_12953);
or U13110 (N_13110,N_12984,N_12659);
nor U13111 (N_13111,N_12642,N_12692);
xor U13112 (N_13112,N_12537,N_12532);
nand U13113 (N_13113,N_12891,N_12641);
and U13114 (N_13114,N_12650,N_12777);
nand U13115 (N_13115,N_12655,N_12917);
xnor U13116 (N_13116,N_12841,N_12948);
or U13117 (N_13117,N_12582,N_12998);
or U13118 (N_13118,N_12877,N_12941);
xor U13119 (N_13119,N_12592,N_12722);
xor U13120 (N_13120,N_12540,N_12977);
or U13121 (N_13121,N_12783,N_12535);
and U13122 (N_13122,N_12618,N_12662);
xnor U13123 (N_13123,N_12564,N_12852);
nor U13124 (N_13124,N_12868,N_12666);
and U13125 (N_13125,N_12936,N_12887);
nor U13126 (N_13126,N_12825,N_12579);
nor U13127 (N_13127,N_12606,N_12528);
nor U13128 (N_13128,N_12566,N_12848);
xor U13129 (N_13129,N_12512,N_12795);
nand U13130 (N_13130,N_12815,N_12683);
nor U13131 (N_13131,N_12914,N_12538);
nand U13132 (N_13132,N_12653,N_12844);
xnor U13133 (N_13133,N_12734,N_12782);
nand U13134 (N_13134,N_12689,N_12680);
and U13135 (N_13135,N_12831,N_12557);
nor U13136 (N_13136,N_12620,N_12675);
nand U13137 (N_13137,N_12570,N_12504);
or U13138 (N_13138,N_12927,N_12743);
xnor U13139 (N_13139,N_12932,N_12589);
and U13140 (N_13140,N_12823,N_12874);
nor U13141 (N_13141,N_12677,N_12871);
or U13142 (N_13142,N_12553,N_12784);
nand U13143 (N_13143,N_12748,N_12690);
or U13144 (N_13144,N_12727,N_12595);
and U13145 (N_13145,N_12632,N_12718);
nor U13146 (N_13146,N_12781,N_12558);
and U13147 (N_13147,N_12888,N_12644);
nand U13148 (N_13148,N_12786,N_12838);
nor U13149 (N_13149,N_12942,N_12686);
xnor U13150 (N_13150,N_12733,N_12635);
xor U13151 (N_13151,N_12792,N_12704);
nor U13152 (N_13152,N_12799,N_12701);
xor U13153 (N_13153,N_12607,N_12699);
or U13154 (N_13154,N_12707,N_12895);
nor U13155 (N_13155,N_12753,N_12629);
and U13156 (N_13156,N_12975,N_12836);
xnor U13157 (N_13157,N_12708,N_12778);
nor U13158 (N_13158,N_12800,N_12923);
or U13159 (N_13159,N_12625,N_12657);
xor U13160 (N_13160,N_12712,N_12585);
and U13161 (N_13161,N_12647,N_12860);
nor U13162 (N_13162,N_12536,N_12966);
and U13163 (N_13163,N_12890,N_12859);
nand U13164 (N_13164,N_12996,N_12892);
nor U13165 (N_13165,N_12732,N_12832);
xor U13166 (N_13166,N_12593,N_12974);
and U13167 (N_13167,N_12883,N_12568);
xor U13168 (N_13168,N_12970,N_12789);
nand U13169 (N_13169,N_12652,N_12742);
xnor U13170 (N_13170,N_12934,N_12845);
xnor U13171 (N_13171,N_12767,N_12610);
nor U13172 (N_13172,N_12750,N_12962);
or U13173 (N_13173,N_12963,N_12857);
nor U13174 (N_13174,N_12828,N_12515);
or U13175 (N_13175,N_12530,N_12745);
nor U13176 (N_13176,N_12604,N_12670);
nand U13177 (N_13177,N_12648,N_12586);
nand U13178 (N_13178,N_12640,N_12765);
or U13179 (N_13179,N_12853,N_12674);
nor U13180 (N_13180,N_12514,N_12912);
and U13181 (N_13181,N_12967,N_12937);
nand U13182 (N_13182,N_12702,N_12873);
nor U13183 (N_13183,N_12924,N_12973);
nand U13184 (N_13184,N_12957,N_12768);
nor U13185 (N_13185,N_12565,N_12896);
nand U13186 (N_13186,N_12876,N_12906);
xnor U13187 (N_13187,N_12746,N_12950);
or U13188 (N_13188,N_12955,N_12527);
or U13189 (N_13189,N_12929,N_12673);
nand U13190 (N_13190,N_12563,N_12986);
or U13191 (N_13191,N_12605,N_12546);
nor U13192 (N_13192,N_12796,N_12621);
or U13193 (N_13193,N_12738,N_12959);
or U13194 (N_13194,N_12711,N_12574);
xor U13195 (N_13195,N_12633,N_12940);
nand U13196 (N_13196,N_12807,N_12798);
xnor U13197 (N_13197,N_12705,N_12961);
nor U13198 (N_13198,N_12578,N_12856);
and U13199 (N_13199,N_12947,N_12665);
nor U13200 (N_13200,N_12548,N_12904);
xnor U13201 (N_13201,N_12624,N_12603);
nand U13202 (N_13202,N_12903,N_12981);
nand U13203 (N_13203,N_12676,N_12902);
and U13204 (N_13204,N_12930,N_12519);
nor U13205 (N_13205,N_12543,N_12602);
nand U13206 (N_13206,N_12956,N_12872);
nand U13207 (N_13207,N_12855,N_12630);
and U13208 (N_13208,N_12649,N_12884);
and U13209 (N_13209,N_12945,N_12555);
nand U13210 (N_13210,N_12612,N_12513);
nand U13211 (N_13211,N_12687,N_12992);
nand U13212 (N_13212,N_12851,N_12994);
or U13213 (N_13213,N_12794,N_12801);
nor U13214 (N_13214,N_12507,N_12757);
or U13215 (N_13215,N_12755,N_12544);
nor U13216 (N_13216,N_12965,N_12725);
nand U13217 (N_13217,N_12719,N_12885);
and U13218 (N_13218,N_12995,N_12779);
nor U13219 (N_13219,N_12938,N_12685);
xnor U13220 (N_13220,N_12908,N_12737);
and U13221 (N_13221,N_12763,N_12671);
nand U13222 (N_13222,N_12813,N_12698);
xnor U13223 (N_13223,N_12762,N_12691);
nand U13224 (N_13224,N_12511,N_12525);
and U13225 (N_13225,N_12639,N_12960);
xnor U13226 (N_13226,N_12811,N_12660);
and U13227 (N_13227,N_12508,N_12809);
nor U13228 (N_13228,N_12979,N_12764);
and U13229 (N_13229,N_12788,N_12584);
or U13230 (N_13230,N_12804,N_12949);
xor U13231 (N_13231,N_12576,N_12747);
or U13232 (N_13232,N_12829,N_12684);
or U13233 (N_13233,N_12700,N_12728);
nor U13234 (N_13234,N_12780,N_12919);
and U13235 (N_13235,N_12627,N_12969);
xnor U13236 (N_13236,N_12545,N_12726);
nand U13237 (N_13237,N_12744,N_12863);
and U13238 (N_13238,N_12985,N_12834);
nor U13239 (N_13239,N_12560,N_12821);
xnor U13240 (N_13240,N_12500,N_12502);
nand U13241 (N_13241,N_12628,N_12751);
or U13242 (N_13242,N_12631,N_12898);
or U13243 (N_13243,N_12988,N_12616);
or U13244 (N_13244,N_12909,N_12688);
xor U13245 (N_13245,N_12920,N_12529);
nor U13246 (N_13246,N_12681,N_12740);
or U13247 (N_13247,N_12581,N_12503);
nand U13248 (N_13248,N_12598,N_12731);
nor U13249 (N_13249,N_12615,N_12946);
and U13250 (N_13250,N_12715,N_12837);
or U13251 (N_13251,N_12884,N_12690);
and U13252 (N_13252,N_12605,N_12923);
or U13253 (N_13253,N_12569,N_12515);
or U13254 (N_13254,N_12614,N_12709);
xnor U13255 (N_13255,N_12613,N_12680);
and U13256 (N_13256,N_12827,N_12651);
nand U13257 (N_13257,N_12536,N_12763);
nand U13258 (N_13258,N_12762,N_12893);
or U13259 (N_13259,N_12698,N_12773);
nand U13260 (N_13260,N_12636,N_12555);
xnor U13261 (N_13261,N_12811,N_12840);
nor U13262 (N_13262,N_12940,N_12557);
nand U13263 (N_13263,N_12900,N_12651);
nand U13264 (N_13264,N_12884,N_12706);
or U13265 (N_13265,N_12977,N_12848);
and U13266 (N_13266,N_12558,N_12631);
nor U13267 (N_13267,N_12936,N_12825);
nand U13268 (N_13268,N_12932,N_12650);
nor U13269 (N_13269,N_12927,N_12934);
nor U13270 (N_13270,N_12582,N_12514);
or U13271 (N_13271,N_12846,N_12837);
and U13272 (N_13272,N_12912,N_12621);
xor U13273 (N_13273,N_12980,N_12745);
and U13274 (N_13274,N_12879,N_12880);
nor U13275 (N_13275,N_12677,N_12527);
xnor U13276 (N_13276,N_12617,N_12637);
and U13277 (N_13277,N_12635,N_12727);
and U13278 (N_13278,N_12863,N_12552);
and U13279 (N_13279,N_12988,N_12925);
or U13280 (N_13280,N_12887,N_12969);
nor U13281 (N_13281,N_12504,N_12658);
or U13282 (N_13282,N_12753,N_12526);
nand U13283 (N_13283,N_12879,N_12843);
and U13284 (N_13284,N_12730,N_12881);
nand U13285 (N_13285,N_12606,N_12987);
and U13286 (N_13286,N_12588,N_12516);
and U13287 (N_13287,N_12668,N_12972);
xor U13288 (N_13288,N_12671,N_12853);
xnor U13289 (N_13289,N_12559,N_12920);
nand U13290 (N_13290,N_12680,N_12547);
nand U13291 (N_13291,N_12647,N_12579);
nand U13292 (N_13292,N_12546,N_12600);
nand U13293 (N_13293,N_12888,N_12879);
xnor U13294 (N_13294,N_12647,N_12597);
xnor U13295 (N_13295,N_12891,N_12744);
nor U13296 (N_13296,N_12554,N_12570);
nand U13297 (N_13297,N_12805,N_12821);
xor U13298 (N_13298,N_12999,N_12893);
xor U13299 (N_13299,N_12777,N_12739);
xor U13300 (N_13300,N_12515,N_12629);
nand U13301 (N_13301,N_12812,N_12528);
nor U13302 (N_13302,N_12782,N_12644);
nand U13303 (N_13303,N_12787,N_12939);
nor U13304 (N_13304,N_12963,N_12541);
nor U13305 (N_13305,N_12767,N_12711);
and U13306 (N_13306,N_12595,N_12579);
nand U13307 (N_13307,N_12689,N_12772);
and U13308 (N_13308,N_12604,N_12710);
and U13309 (N_13309,N_12954,N_12524);
nor U13310 (N_13310,N_12987,N_12767);
nor U13311 (N_13311,N_12892,N_12547);
and U13312 (N_13312,N_12707,N_12698);
or U13313 (N_13313,N_12818,N_12926);
nor U13314 (N_13314,N_12618,N_12551);
nor U13315 (N_13315,N_12562,N_12530);
xnor U13316 (N_13316,N_12614,N_12633);
xnor U13317 (N_13317,N_12512,N_12537);
or U13318 (N_13318,N_12700,N_12542);
nand U13319 (N_13319,N_12533,N_12924);
xor U13320 (N_13320,N_12610,N_12514);
or U13321 (N_13321,N_12855,N_12750);
or U13322 (N_13322,N_12584,N_12750);
nor U13323 (N_13323,N_12830,N_12518);
nand U13324 (N_13324,N_12745,N_12777);
nor U13325 (N_13325,N_12972,N_12591);
nand U13326 (N_13326,N_12787,N_12623);
nand U13327 (N_13327,N_12586,N_12743);
xor U13328 (N_13328,N_12856,N_12850);
xor U13329 (N_13329,N_12810,N_12806);
and U13330 (N_13330,N_12527,N_12860);
nor U13331 (N_13331,N_12868,N_12796);
and U13332 (N_13332,N_12980,N_12614);
and U13333 (N_13333,N_12551,N_12678);
xor U13334 (N_13334,N_12542,N_12987);
nand U13335 (N_13335,N_12780,N_12728);
nand U13336 (N_13336,N_12502,N_12650);
nand U13337 (N_13337,N_12991,N_12759);
and U13338 (N_13338,N_12852,N_12835);
or U13339 (N_13339,N_12737,N_12838);
nand U13340 (N_13340,N_12882,N_12670);
nor U13341 (N_13341,N_12966,N_12909);
nand U13342 (N_13342,N_12915,N_12725);
nor U13343 (N_13343,N_12986,N_12640);
or U13344 (N_13344,N_12566,N_12660);
nor U13345 (N_13345,N_12549,N_12645);
and U13346 (N_13346,N_12560,N_12852);
or U13347 (N_13347,N_12828,N_12659);
nand U13348 (N_13348,N_12803,N_12562);
and U13349 (N_13349,N_12654,N_12859);
nor U13350 (N_13350,N_12501,N_12999);
and U13351 (N_13351,N_12896,N_12806);
and U13352 (N_13352,N_12536,N_12864);
nand U13353 (N_13353,N_12883,N_12984);
nor U13354 (N_13354,N_12986,N_12577);
nor U13355 (N_13355,N_12554,N_12835);
nor U13356 (N_13356,N_12575,N_12726);
nand U13357 (N_13357,N_12950,N_12750);
xnor U13358 (N_13358,N_12879,N_12818);
nor U13359 (N_13359,N_12519,N_12947);
nand U13360 (N_13360,N_12739,N_12813);
xnor U13361 (N_13361,N_12536,N_12712);
or U13362 (N_13362,N_12881,N_12549);
and U13363 (N_13363,N_12671,N_12683);
and U13364 (N_13364,N_12846,N_12518);
and U13365 (N_13365,N_12852,N_12931);
nand U13366 (N_13366,N_12774,N_12634);
nand U13367 (N_13367,N_12536,N_12761);
nor U13368 (N_13368,N_12682,N_12705);
nand U13369 (N_13369,N_12765,N_12731);
nor U13370 (N_13370,N_12933,N_12652);
or U13371 (N_13371,N_12516,N_12935);
and U13372 (N_13372,N_12996,N_12895);
xor U13373 (N_13373,N_12723,N_12697);
nor U13374 (N_13374,N_12953,N_12515);
xor U13375 (N_13375,N_12566,N_12591);
xnor U13376 (N_13376,N_12617,N_12628);
or U13377 (N_13377,N_12889,N_12949);
or U13378 (N_13378,N_12860,N_12568);
or U13379 (N_13379,N_12636,N_12797);
or U13380 (N_13380,N_12517,N_12807);
and U13381 (N_13381,N_12664,N_12920);
or U13382 (N_13382,N_12768,N_12577);
nor U13383 (N_13383,N_12614,N_12947);
nor U13384 (N_13384,N_12753,N_12898);
and U13385 (N_13385,N_12852,N_12960);
xor U13386 (N_13386,N_12574,N_12800);
nor U13387 (N_13387,N_12954,N_12679);
nor U13388 (N_13388,N_12963,N_12851);
nor U13389 (N_13389,N_12630,N_12816);
and U13390 (N_13390,N_12937,N_12958);
xnor U13391 (N_13391,N_12502,N_12991);
nor U13392 (N_13392,N_12572,N_12881);
and U13393 (N_13393,N_12600,N_12907);
nand U13394 (N_13394,N_12668,N_12824);
or U13395 (N_13395,N_12934,N_12533);
and U13396 (N_13396,N_12772,N_12598);
or U13397 (N_13397,N_12843,N_12623);
or U13398 (N_13398,N_12790,N_12892);
xnor U13399 (N_13399,N_12915,N_12892);
nand U13400 (N_13400,N_12509,N_12827);
nor U13401 (N_13401,N_12894,N_12881);
and U13402 (N_13402,N_12957,N_12745);
or U13403 (N_13403,N_12752,N_12956);
nand U13404 (N_13404,N_12920,N_12902);
xnor U13405 (N_13405,N_12624,N_12715);
nand U13406 (N_13406,N_12942,N_12771);
and U13407 (N_13407,N_12581,N_12593);
nor U13408 (N_13408,N_12602,N_12723);
xnor U13409 (N_13409,N_12885,N_12566);
nor U13410 (N_13410,N_12705,N_12592);
xnor U13411 (N_13411,N_12582,N_12986);
and U13412 (N_13412,N_12914,N_12604);
or U13413 (N_13413,N_12914,N_12646);
and U13414 (N_13414,N_12659,N_12972);
nand U13415 (N_13415,N_12738,N_12589);
or U13416 (N_13416,N_12514,N_12713);
and U13417 (N_13417,N_12858,N_12780);
or U13418 (N_13418,N_12724,N_12582);
nand U13419 (N_13419,N_12834,N_12759);
nand U13420 (N_13420,N_12974,N_12984);
nand U13421 (N_13421,N_12712,N_12923);
and U13422 (N_13422,N_12820,N_12667);
nor U13423 (N_13423,N_12580,N_12810);
xnor U13424 (N_13424,N_12789,N_12765);
nand U13425 (N_13425,N_12690,N_12646);
or U13426 (N_13426,N_12643,N_12725);
and U13427 (N_13427,N_12925,N_12786);
xnor U13428 (N_13428,N_12523,N_12889);
and U13429 (N_13429,N_12930,N_12936);
or U13430 (N_13430,N_12798,N_12873);
or U13431 (N_13431,N_12566,N_12866);
or U13432 (N_13432,N_12958,N_12881);
or U13433 (N_13433,N_12556,N_12558);
nand U13434 (N_13434,N_12858,N_12836);
nand U13435 (N_13435,N_12583,N_12679);
or U13436 (N_13436,N_12770,N_12824);
nor U13437 (N_13437,N_12977,N_12640);
xor U13438 (N_13438,N_12695,N_12767);
nand U13439 (N_13439,N_12509,N_12982);
and U13440 (N_13440,N_12517,N_12625);
and U13441 (N_13441,N_12654,N_12946);
nor U13442 (N_13442,N_12632,N_12760);
xnor U13443 (N_13443,N_12582,N_12939);
or U13444 (N_13444,N_12876,N_12871);
or U13445 (N_13445,N_12997,N_12881);
and U13446 (N_13446,N_12592,N_12825);
or U13447 (N_13447,N_12554,N_12715);
or U13448 (N_13448,N_12748,N_12746);
and U13449 (N_13449,N_12775,N_12772);
and U13450 (N_13450,N_12887,N_12658);
nand U13451 (N_13451,N_12837,N_12623);
nor U13452 (N_13452,N_12961,N_12529);
nor U13453 (N_13453,N_12652,N_12772);
nor U13454 (N_13454,N_12550,N_12920);
xor U13455 (N_13455,N_12516,N_12737);
nand U13456 (N_13456,N_12931,N_12800);
or U13457 (N_13457,N_12921,N_12731);
or U13458 (N_13458,N_12947,N_12907);
nor U13459 (N_13459,N_12971,N_12753);
nand U13460 (N_13460,N_12908,N_12709);
nor U13461 (N_13461,N_12882,N_12657);
xor U13462 (N_13462,N_12655,N_12686);
or U13463 (N_13463,N_12663,N_12929);
nand U13464 (N_13464,N_12743,N_12875);
xor U13465 (N_13465,N_12519,N_12777);
and U13466 (N_13466,N_12624,N_12782);
or U13467 (N_13467,N_12626,N_12681);
or U13468 (N_13468,N_12591,N_12927);
and U13469 (N_13469,N_12891,N_12750);
nand U13470 (N_13470,N_12961,N_12819);
nand U13471 (N_13471,N_12562,N_12554);
xor U13472 (N_13472,N_12935,N_12738);
nand U13473 (N_13473,N_12746,N_12700);
nand U13474 (N_13474,N_12737,N_12596);
nand U13475 (N_13475,N_12911,N_12623);
nand U13476 (N_13476,N_12525,N_12910);
and U13477 (N_13477,N_12976,N_12543);
nand U13478 (N_13478,N_12630,N_12837);
nor U13479 (N_13479,N_12513,N_12729);
xnor U13480 (N_13480,N_12755,N_12523);
nand U13481 (N_13481,N_12928,N_12786);
nand U13482 (N_13482,N_12721,N_12521);
nand U13483 (N_13483,N_12563,N_12568);
nand U13484 (N_13484,N_12584,N_12942);
nand U13485 (N_13485,N_12871,N_12907);
nand U13486 (N_13486,N_12619,N_12866);
and U13487 (N_13487,N_12925,N_12716);
nand U13488 (N_13488,N_12700,N_12801);
nand U13489 (N_13489,N_12976,N_12627);
nand U13490 (N_13490,N_12564,N_12819);
or U13491 (N_13491,N_12852,N_12936);
nand U13492 (N_13492,N_12858,N_12884);
nor U13493 (N_13493,N_12758,N_12685);
and U13494 (N_13494,N_12953,N_12787);
or U13495 (N_13495,N_12510,N_12958);
nor U13496 (N_13496,N_12555,N_12862);
nand U13497 (N_13497,N_12506,N_12994);
nand U13498 (N_13498,N_12826,N_12897);
and U13499 (N_13499,N_12671,N_12749);
nor U13500 (N_13500,N_13221,N_13290);
nor U13501 (N_13501,N_13258,N_13297);
nor U13502 (N_13502,N_13381,N_13322);
nor U13503 (N_13503,N_13261,N_13214);
nand U13504 (N_13504,N_13362,N_13113);
nor U13505 (N_13505,N_13360,N_13382);
nor U13506 (N_13506,N_13013,N_13193);
nor U13507 (N_13507,N_13406,N_13438);
and U13508 (N_13508,N_13153,N_13336);
nand U13509 (N_13509,N_13204,N_13256);
nand U13510 (N_13510,N_13385,N_13146);
xnor U13511 (N_13511,N_13374,N_13288);
or U13512 (N_13512,N_13461,N_13028);
nand U13513 (N_13513,N_13149,N_13138);
nor U13514 (N_13514,N_13430,N_13248);
xnor U13515 (N_13515,N_13283,N_13450);
nand U13516 (N_13516,N_13154,N_13400);
xnor U13517 (N_13517,N_13323,N_13188);
xor U13518 (N_13518,N_13189,N_13464);
or U13519 (N_13519,N_13325,N_13462);
nand U13520 (N_13520,N_13286,N_13407);
xnor U13521 (N_13521,N_13235,N_13492);
nor U13522 (N_13522,N_13303,N_13043);
and U13523 (N_13523,N_13415,N_13165);
or U13524 (N_13524,N_13309,N_13279);
nor U13525 (N_13525,N_13191,N_13140);
xor U13526 (N_13526,N_13349,N_13106);
nor U13527 (N_13527,N_13120,N_13050);
and U13528 (N_13528,N_13240,N_13077);
xor U13529 (N_13529,N_13029,N_13114);
or U13530 (N_13530,N_13367,N_13259);
or U13531 (N_13531,N_13425,N_13321);
xnor U13532 (N_13532,N_13020,N_13163);
xor U13533 (N_13533,N_13408,N_13216);
and U13534 (N_13534,N_13172,N_13122);
nand U13535 (N_13535,N_13411,N_13269);
nor U13536 (N_13536,N_13328,N_13477);
nand U13537 (N_13537,N_13098,N_13257);
and U13538 (N_13538,N_13389,N_13469);
xnor U13539 (N_13539,N_13318,N_13335);
or U13540 (N_13540,N_13068,N_13158);
nand U13541 (N_13541,N_13481,N_13010);
and U13542 (N_13542,N_13368,N_13080);
nor U13543 (N_13543,N_13465,N_13093);
or U13544 (N_13544,N_13420,N_13412);
nand U13545 (N_13545,N_13441,N_13003);
xor U13546 (N_13546,N_13499,N_13075);
nand U13547 (N_13547,N_13126,N_13409);
nor U13548 (N_13548,N_13136,N_13436);
nand U13549 (N_13549,N_13074,N_13363);
nor U13550 (N_13550,N_13118,N_13238);
nand U13551 (N_13551,N_13039,N_13044);
nand U13552 (N_13552,N_13069,N_13317);
and U13553 (N_13553,N_13078,N_13147);
and U13554 (N_13554,N_13372,N_13180);
nand U13555 (N_13555,N_13394,N_13366);
nor U13556 (N_13556,N_13173,N_13311);
nand U13557 (N_13557,N_13466,N_13061);
or U13558 (N_13558,N_13485,N_13038);
nand U13559 (N_13559,N_13179,N_13232);
xor U13560 (N_13560,N_13176,N_13398);
or U13561 (N_13561,N_13159,N_13280);
and U13562 (N_13562,N_13351,N_13255);
or U13563 (N_13563,N_13359,N_13135);
nor U13564 (N_13564,N_13087,N_13222);
nor U13565 (N_13565,N_13373,N_13437);
nor U13566 (N_13566,N_13446,N_13249);
and U13567 (N_13567,N_13234,N_13137);
nand U13568 (N_13568,N_13442,N_13293);
nand U13569 (N_13569,N_13445,N_13081);
nor U13570 (N_13570,N_13205,N_13049);
nand U13571 (N_13571,N_13236,N_13308);
nor U13572 (N_13572,N_13379,N_13211);
and U13573 (N_13573,N_13484,N_13350);
nand U13574 (N_13574,N_13008,N_13353);
nor U13575 (N_13575,N_13427,N_13375);
or U13576 (N_13576,N_13145,N_13117);
xnor U13577 (N_13577,N_13134,N_13181);
nor U13578 (N_13578,N_13162,N_13296);
and U13579 (N_13579,N_13455,N_13105);
nand U13580 (N_13580,N_13094,N_13055);
or U13581 (N_13581,N_13054,N_13210);
and U13582 (N_13582,N_13376,N_13056);
nand U13583 (N_13583,N_13226,N_13027);
xnor U13584 (N_13584,N_13355,N_13183);
or U13585 (N_13585,N_13109,N_13312);
or U13586 (N_13586,N_13058,N_13460);
nand U13587 (N_13587,N_13289,N_13454);
xor U13588 (N_13588,N_13017,N_13313);
xnor U13589 (N_13589,N_13048,N_13202);
nand U13590 (N_13590,N_13433,N_13397);
nand U13591 (N_13591,N_13228,N_13292);
nor U13592 (N_13592,N_13468,N_13219);
nor U13593 (N_13593,N_13199,N_13268);
and U13594 (N_13594,N_13085,N_13042);
or U13595 (N_13595,N_13063,N_13000);
xnor U13596 (N_13596,N_13095,N_13218);
xor U13597 (N_13597,N_13449,N_13340);
and U13598 (N_13598,N_13090,N_13101);
xnor U13599 (N_13599,N_13057,N_13198);
or U13600 (N_13600,N_13267,N_13266);
xor U13601 (N_13601,N_13096,N_13024);
xnor U13602 (N_13602,N_13045,N_13439);
and U13603 (N_13603,N_13476,N_13273);
nor U13604 (N_13604,N_13005,N_13347);
nand U13605 (N_13605,N_13178,N_13060);
nor U13606 (N_13606,N_13016,N_13025);
xnor U13607 (N_13607,N_13348,N_13377);
xnor U13608 (N_13608,N_13144,N_13231);
nand U13609 (N_13609,N_13380,N_13082);
or U13610 (N_13610,N_13151,N_13007);
and U13611 (N_13611,N_13329,N_13316);
xor U13612 (N_13612,N_13285,N_13129);
nor U13613 (N_13613,N_13475,N_13421);
nand U13614 (N_13614,N_13371,N_13130);
nand U13615 (N_13615,N_13343,N_13148);
and U13616 (N_13616,N_13458,N_13486);
or U13617 (N_13617,N_13463,N_13429);
nand U13618 (N_13618,N_13229,N_13459);
nor U13619 (N_13619,N_13456,N_13097);
and U13620 (N_13620,N_13324,N_13496);
xnor U13621 (N_13621,N_13277,N_13295);
or U13622 (N_13622,N_13062,N_13047);
nand U13623 (N_13623,N_13253,N_13209);
nand U13624 (N_13624,N_13300,N_13070);
or U13625 (N_13625,N_13489,N_13124);
nor U13626 (N_13626,N_13370,N_13395);
or U13627 (N_13627,N_13190,N_13051);
nor U13628 (N_13628,N_13391,N_13417);
nand U13629 (N_13629,N_13143,N_13021);
nor U13630 (N_13630,N_13224,N_13107);
or U13631 (N_13631,N_13073,N_13046);
or U13632 (N_13632,N_13012,N_13041);
nor U13633 (N_13633,N_13457,N_13424);
nand U13634 (N_13634,N_13416,N_13006);
nand U13635 (N_13635,N_13497,N_13473);
or U13636 (N_13636,N_13083,N_13015);
or U13637 (N_13637,N_13208,N_13337);
and U13638 (N_13638,N_13037,N_13440);
nor U13639 (N_13639,N_13128,N_13254);
xor U13640 (N_13640,N_13088,N_13092);
and U13641 (N_13641,N_13091,N_13494);
xnor U13642 (N_13642,N_13365,N_13123);
or U13643 (N_13643,N_13213,N_13299);
or U13644 (N_13644,N_13245,N_13184);
xor U13645 (N_13645,N_13166,N_13405);
and U13646 (N_13646,N_13200,N_13393);
nand U13647 (N_13647,N_13423,N_13150);
nand U13648 (N_13648,N_13387,N_13023);
and U13649 (N_13649,N_13401,N_13067);
and U13650 (N_13650,N_13009,N_13197);
nand U13651 (N_13651,N_13033,N_13327);
nor U13652 (N_13652,N_13378,N_13242);
nand U13653 (N_13653,N_13241,N_13342);
xnor U13654 (N_13654,N_13281,N_13170);
and U13655 (N_13655,N_13396,N_13244);
xor U13656 (N_13656,N_13490,N_13444);
or U13657 (N_13657,N_13426,N_13471);
nor U13658 (N_13658,N_13001,N_13326);
xnor U13659 (N_13659,N_13203,N_13142);
nor U13660 (N_13660,N_13125,N_13345);
and U13661 (N_13661,N_13434,N_13186);
and U13662 (N_13662,N_13443,N_13103);
xnor U13663 (N_13663,N_13246,N_13399);
nand U13664 (N_13664,N_13282,N_13152);
xnor U13665 (N_13665,N_13247,N_13495);
or U13666 (N_13666,N_13018,N_13237);
xnor U13667 (N_13667,N_13072,N_13467);
or U13668 (N_13668,N_13390,N_13319);
or U13669 (N_13669,N_13196,N_13115);
xor U13670 (N_13670,N_13291,N_13212);
xnor U13671 (N_13671,N_13104,N_13004);
or U13672 (N_13672,N_13386,N_13334);
or U13673 (N_13673,N_13171,N_13472);
nand U13674 (N_13674,N_13155,N_13089);
or U13675 (N_13675,N_13369,N_13161);
and U13676 (N_13676,N_13356,N_13410);
and U13677 (N_13677,N_13320,N_13315);
and U13678 (N_13678,N_13206,N_13182);
or U13679 (N_13679,N_13435,N_13121);
nor U13680 (N_13680,N_13002,N_13305);
and U13681 (N_13681,N_13265,N_13052);
xnor U13682 (N_13682,N_13064,N_13160);
or U13683 (N_13683,N_13304,N_13341);
or U13684 (N_13684,N_13071,N_13223);
nand U13685 (N_13685,N_13272,N_13331);
and U13686 (N_13686,N_13156,N_13065);
nand U13687 (N_13687,N_13413,N_13086);
nor U13688 (N_13688,N_13307,N_13034);
xnor U13689 (N_13689,N_13243,N_13169);
and U13690 (N_13690,N_13030,N_13491);
xnor U13691 (N_13691,N_13019,N_13402);
or U13692 (N_13692,N_13358,N_13479);
xor U13693 (N_13693,N_13217,N_13357);
nand U13694 (N_13694,N_13195,N_13252);
xnor U13695 (N_13695,N_13333,N_13302);
or U13696 (N_13696,N_13177,N_13164);
xnor U13697 (N_13697,N_13066,N_13230);
nor U13698 (N_13698,N_13059,N_13278);
and U13699 (N_13699,N_13014,N_13157);
xor U13700 (N_13700,N_13201,N_13011);
xnor U13701 (N_13701,N_13493,N_13141);
or U13702 (N_13702,N_13383,N_13036);
nor U13703 (N_13703,N_13276,N_13076);
xnor U13704 (N_13704,N_13225,N_13330);
xnor U13705 (N_13705,N_13275,N_13127);
or U13706 (N_13706,N_13132,N_13298);
nand U13707 (N_13707,N_13262,N_13384);
xnor U13708 (N_13708,N_13470,N_13031);
xor U13709 (N_13709,N_13116,N_13270);
xor U13710 (N_13710,N_13284,N_13451);
nor U13711 (N_13711,N_13239,N_13498);
xnor U13712 (N_13712,N_13185,N_13346);
and U13713 (N_13713,N_13287,N_13428);
nor U13714 (N_13714,N_13022,N_13187);
nor U13715 (N_13715,N_13168,N_13263);
and U13716 (N_13716,N_13175,N_13388);
and U13717 (N_13717,N_13338,N_13301);
nor U13718 (N_13718,N_13306,N_13487);
nand U13719 (N_13719,N_13364,N_13419);
nor U13720 (N_13720,N_13354,N_13079);
xnor U13721 (N_13721,N_13310,N_13431);
xor U13722 (N_13722,N_13131,N_13251);
xnor U13723 (N_13723,N_13332,N_13215);
and U13724 (N_13724,N_13344,N_13482);
nor U13725 (N_13725,N_13119,N_13448);
nor U13726 (N_13726,N_13100,N_13133);
nand U13727 (N_13727,N_13053,N_13110);
nand U13728 (N_13728,N_13207,N_13174);
or U13729 (N_13729,N_13314,N_13271);
xnor U13730 (N_13730,N_13418,N_13260);
nor U13731 (N_13731,N_13361,N_13111);
and U13732 (N_13732,N_13035,N_13483);
or U13733 (N_13733,N_13480,N_13264);
or U13734 (N_13734,N_13026,N_13167);
and U13735 (N_13735,N_13220,N_13404);
nor U13736 (N_13736,N_13099,N_13488);
nor U13737 (N_13737,N_13352,N_13192);
or U13738 (N_13738,N_13422,N_13478);
nor U13739 (N_13739,N_13102,N_13112);
nand U13740 (N_13740,N_13392,N_13339);
xnor U13741 (N_13741,N_13233,N_13139);
and U13742 (N_13742,N_13032,N_13250);
nand U13743 (N_13743,N_13414,N_13474);
or U13744 (N_13744,N_13194,N_13294);
nand U13745 (N_13745,N_13040,N_13274);
or U13746 (N_13746,N_13452,N_13108);
and U13747 (N_13747,N_13084,N_13227);
or U13748 (N_13748,N_13453,N_13432);
nand U13749 (N_13749,N_13447,N_13403);
xor U13750 (N_13750,N_13022,N_13323);
xor U13751 (N_13751,N_13069,N_13044);
nor U13752 (N_13752,N_13123,N_13092);
and U13753 (N_13753,N_13034,N_13349);
xnor U13754 (N_13754,N_13068,N_13266);
or U13755 (N_13755,N_13434,N_13234);
or U13756 (N_13756,N_13406,N_13186);
nor U13757 (N_13757,N_13326,N_13298);
nor U13758 (N_13758,N_13236,N_13291);
xor U13759 (N_13759,N_13464,N_13159);
nor U13760 (N_13760,N_13481,N_13173);
nand U13761 (N_13761,N_13131,N_13031);
and U13762 (N_13762,N_13120,N_13324);
or U13763 (N_13763,N_13311,N_13095);
xnor U13764 (N_13764,N_13415,N_13250);
nand U13765 (N_13765,N_13243,N_13162);
xor U13766 (N_13766,N_13308,N_13357);
or U13767 (N_13767,N_13234,N_13238);
or U13768 (N_13768,N_13210,N_13018);
or U13769 (N_13769,N_13309,N_13354);
nand U13770 (N_13770,N_13319,N_13463);
nor U13771 (N_13771,N_13251,N_13192);
and U13772 (N_13772,N_13141,N_13181);
and U13773 (N_13773,N_13081,N_13077);
xor U13774 (N_13774,N_13279,N_13378);
nor U13775 (N_13775,N_13272,N_13019);
or U13776 (N_13776,N_13098,N_13120);
nor U13777 (N_13777,N_13075,N_13300);
or U13778 (N_13778,N_13048,N_13191);
or U13779 (N_13779,N_13308,N_13449);
xor U13780 (N_13780,N_13169,N_13089);
xnor U13781 (N_13781,N_13466,N_13220);
or U13782 (N_13782,N_13454,N_13338);
nand U13783 (N_13783,N_13419,N_13389);
nor U13784 (N_13784,N_13498,N_13075);
nand U13785 (N_13785,N_13105,N_13308);
nand U13786 (N_13786,N_13452,N_13145);
nor U13787 (N_13787,N_13203,N_13085);
nand U13788 (N_13788,N_13440,N_13279);
and U13789 (N_13789,N_13386,N_13086);
nand U13790 (N_13790,N_13013,N_13197);
xnor U13791 (N_13791,N_13194,N_13334);
or U13792 (N_13792,N_13178,N_13001);
nor U13793 (N_13793,N_13374,N_13164);
xor U13794 (N_13794,N_13444,N_13099);
nand U13795 (N_13795,N_13211,N_13191);
and U13796 (N_13796,N_13190,N_13120);
nor U13797 (N_13797,N_13333,N_13439);
nor U13798 (N_13798,N_13295,N_13153);
nor U13799 (N_13799,N_13054,N_13418);
nor U13800 (N_13800,N_13078,N_13475);
and U13801 (N_13801,N_13062,N_13144);
nor U13802 (N_13802,N_13133,N_13387);
or U13803 (N_13803,N_13464,N_13467);
xor U13804 (N_13804,N_13198,N_13460);
nor U13805 (N_13805,N_13451,N_13480);
xor U13806 (N_13806,N_13002,N_13492);
nand U13807 (N_13807,N_13119,N_13060);
nor U13808 (N_13808,N_13476,N_13005);
or U13809 (N_13809,N_13322,N_13199);
xnor U13810 (N_13810,N_13346,N_13115);
and U13811 (N_13811,N_13079,N_13126);
nand U13812 (N_13812,N_13474,N_13490);
and U13813 (N_13813,N_13288,N_13348);
xnor U13814 (N_13814,N_13203,N_13215);
nor U13815 (N_13815,N_13273,N_13413);
nand U13816 (N_13816,N_13142,N_13187);
xor U13817 (N_13817,N_13321,N_13077);
nor U13818 (N_13818,N_13346,N_13117);
or U13819 (N_13819,N_13419,N_13223);
xnor U13820 (N_13820,N_13222,N_13448);
xor U13821 (N_13821,N_13192,N_13365);
nand U13822 (N_13822,N_13147,N_13474);
nand U13823 (N_13823,N_13059,N_13159);
and U13824 (N_13824,N_13186,N_13358);
or U13825 (N_13825,N_13236,N_13301);
nor U13826 (N_13826,N_13087,N_13486);
and U13827 (N_13827,N_13309,N_13474);
and U13828 (N_13828,N_13014,N_13185);
and U13829 (N_13829,N_13173,N_13422);
nor U13830 (N_13830,N_13017,N_13197);
nor U13831 (N_13831,N_13136,N_13119);
nor U13832 (N_13832,N_13209,N_13146);
nand U13833 (N_13833,N_13075,N_13226);
or U13834 (N_13834,N_13420,N_13241);
nand U13835 (N_13835,N_13195,N_13394);
and U13836 (N_13836,N_13461,N_13010);
and U13837 (N_13837,N_13032,N_13153);
nand U13838 (N_13838,N_13240,N_13158);
nor U13839 (N_13839,N_13033,N_13206);
xor U13840 (N_13840,N_13243,N_13105);
or U13841 (N_13841,N_13468,N_13240);
xor U13842 (N_13842,N_13491,N_13330);
and U13843 (N_13843,N_13416,N_13471);
xor U13844 (N_13844,N_13332,N_13058);
xnor U13845 (N_13845,N_13064,N_13233);
nor U13846 (N_13846,N_13311,N_13071);
xor U13847 (N_13847,N_13365,N_13222);
xnor U13848 (N_13848,N_13488,N_13436);
or U13849 (N_13849,N_13326,N_13472);
and U13850 (N_13850,N_13146,N_13288);
and U13851 (N_13851,N_13164,N_13369);
nor U13852 (N_13852,N_13238,N_13493);
or U13853 (N_13853,N_13325,N_13142);
nor U13854 (N_13854,N_13198,N_13005);
nor U13855 (N_13855,N_13440,N_13340);
xor U13856 (N_13856,N_13145,N_13037);
or U13857 (N_13857,N_13485,N_13001);
xnor U13858 (N_13858,N_13127,N_13172);
nand U13859 (N_13859,N_13469,N_13371);
nor U13860 (N_13860,N_13496,N_13085);
nand U13861 (N_13861,N_13348,N_13389);
or U13862 (N_13862,N_13354,N_13159);
or U13863 (N_13863,N_13342,N_13332);
or U13864 (N_13864,N_13467,N_13329);
nor U13865 (N_13865,N_13294,N_13049);
or U13866 (N_13866,N_13231,N_13186);
xor U13867 (N_13867,N_13020,N_13485);
nand U13868 (N_13868,N_13039,N_13182);
and U13869 (N_13869,N_13082,N_13228);
or U13870 (N_13870,N_13277,N_13466);
xnor U13871 (N_13871,N_13435,N_13289);
xnor U13872 (N_13872,N_13250,N_13467);
or U13873 (N_13873,N_13240,N_13296);
nand U13874 (N_13874,N_13323,N_13085);
nor U13875 (N_13875,N_13489,N_13223);
nand U13876 (N_13876,N_13460,N_13277);
xnor U13877 (N_13877,N_13483,N_13114);
nor U13878 (N_13878,N_13269,N_13424);
xnor U13879 (N_13879,N_13387,N_13468);
and U13880 (N_13880,N_13452,N_13054);
and U13881 (N_13881,N_13109,N_13452);
and U13882 (N_13882,N_13487,N_13461);
nand U13883 (N_13883,N_13262,N_13140);
nand U13884 (N_13884,N_13267,N_13424);
and U13885 (N_13885,N_13289,N_13014);
nand U13886 (N_13886,N_13239,N_13267);
and U13887 (N_13887,N_13106,N_13084);
or U13888 (N_13888,N_13054,N_13145);
and U13889 (N_13889,N_13147,N_13208);
or U13890 (N_13890,N_13209,N_13485);
xor U13891 (N_13891,N_13456,N_13497);
and U13892 (N_13892,N_13433,N_13066);
xor U13893 (N_13893,N_13192,N_13107);
and U13894 (N_13894,N_13154,N_13124);
xnor U13895 (N_13895,N_13344,N_13062);
xnor U13896 (N_13896,N_13062,N_13186);
nand U13897 (N_13897,N_13104,N_13254);
nand U13898 (N_13898,N_13200,N_13292);
nor U13899 (N_13899,N_13271,N_13233);
or U13900 (N_13900,N_13452,N_13014);
nand U13901 (N_13901,N_13237,N_13247);
or U13902 (N_13902,N_13406,N_13247);
xor U13903 (N_13903,N_13364,N_13086);
xor U13904 (N_13904,N_13261,N_13435);
nand U13905 (N_13905,N_13360,N_13177);
and U13906 (N_13906,N_13430,N_13492);
nor U13907 (N_13907,N_13330,N_13487);
nor U13908 (N_13908,N_13083,N_13050);
nor U13909 (N_13909,N_13135,N_13310);
nor U13910 (N_13910,N_13322,N_13413);
and U13911 (N_13911,N_13098,N_13153);
xnor U13912 (N_13912,N_13148,N_13466);
and U13913 (N_13913,N_13441,N_13426);
and U13914 (N_13914,N_13051,N_13283);
xor U13915 (N_13915,N_13459,N_13443);
xor U13916 (N_13916,N_13394,N_13013);
nand U13917 (N_13917,N_13134,N_13410);
xor U13918 (N_13918,N_13391,N_13043);
nand U13919 (N_13919,N_13119,N_13367);
and U13920 (N_13920,N_13477,N_13311);
nor U13921 (N_13921,N_13181,N_13479);
nand U13922 (N_13922,N_13074,N_13210);
or U13923 (N_13923,N_13226,N_13244);
nor U13924 (N_13924,N_13158,N_13472);
xnor U13925 (N_13925,N_13306,N_13441);
xnor U13926 (N_13926,N_13083,N_13196);
or U13927 (N_13927,N_13231,N_13163);
and U13928 (N_13928,N_13446,N_13126);
and U13929 (N_13929,N_13143,N_13150);
xnor U13930 (N_13930,N_13111,N_13476);
nor U13931 (N_13931,N_13430,N_13227);
nor U13932 (N_13932,N_13293,N_13376);
nand U13933 (N_13933,N_13261,N_13048);
and U13934 (N_13934,N_13360,N_13183);
nor U13935 (N_13935,N_13159,N_13008);
or U13936 (N_13936,N_13224,N_13424);
xnor U13937 (N_13937,N_13181,N_13418);
xor U13938 (N_13938,N_13348,N_13363);
and U13939 (N_13939,N_13275,N_13279);
nor U13940 (N_13940,N_13492,N_13374);
or U13941 (N_13941,N_13237,N_13396);
and U13942 (N_13942,N_13259,N_13215);
or U13943 (N_13943,N_13173,N_13210);
or U13944 (N_13944,N_13153,N_13099);
and U13945 (N_13945,N_13178,N_13426);
xor U13946 (N_13946,N_13075,N_13063);
xor U13947 (N_13947,N_13248,N_13401);
xor U13948 (N_13948,N_13440,N_13125);
nor U13949 (N_13949,N_13132,N_13037);
nand U13950 (N_13950,N_13489,N_13371);
xor U13951 (N_13951,N_13214,N_13056);
and U13952 (N_13952,N_13434,N_13225);
nor U13953 (N_13953,N_13019,N_13452);
xnor U13954 (N_13954,N_13155,N_13217);
nor U13955 (N_13955,N_13226,N_13146);
nor U13956 (N_13956,N_13037,N_13370);
xnor U13957 (N_13957,N_13245,N_13006);
or U13958 (N_13958,N_13151,N_13190);
nor U13959 (N_13959,N_13137,N_13402);
xnor U13960 (N_13960,N_13465,N_13499);
and U13961 (N_13961,N_13111,N_13491);
and U13962 (N_13962,N_13094,N_13143);
or U13963 (N_13963,N_13045,N_13142);
or U13964 (N_13964,N_13318,N_13160);
nand U13965 (N_13965,N_13410,N_13404);
or U13966 (N_13966,N_13325,N_13311);
nor U13967 (N_13967,N_13412,N_13443);
xnor U13968 (N_13968,N_13194,N_13394);
and U13969 (N_13969,N_13293,N_13086);
and U13970 (N_13970,N_13047,N_13042);
and U13971 (N_13971,N_13075,N_13264);
nor U13972 (N_13972,N_13455,N_13419);
nand U13973 (N_13973,N_13349,N_13126);
xor U13974 (N_13974,N_13414,N_13110);
nand U13975 (N_13975,N_13179,N_13314);
nor U13976 (N_13976,N_13111,N_13387);
nand U13977 (N_13977,N_13083,N_13388);
nor U13978 (N_13978,N_13487,N_13109);
and U13979 (N_13979,N_13039,N_13468);
or U13980 (N_13980,N_13284,N_13444);
and U13981 (N_13981,N_13389,N_13355);
nor U13982 (N_13982,N_13181,N_13317);
nand U13983 (N_13983,N_13333,N_13073);
and U13984 (N_13984,N_13065,N_13078);
and U13985 (N_13985,N_13364,N_13360);
nand U13986 (N_13986,N_13350,N_13065);
nor U13987 (N_13987,N_13441,N_13450);
nand U13988 (N_13988,N_13332,N_13357);
nand U13989 (N_13989,N_13460,N_13069);
or U13990 (N_13990,N_13438,N_13173);
and U13991 (N_13991,N_13006,N_13440);
and U13992 (N_13992,N_13284,N_13145);
or U13993 (N_13993,N_13438,N_13208);
or U13994 (N_13994,N_13036,N_13006);
or U13995 (N_13995,N_13195,N_13138);
nand U13996 (N_13996,N_13113,N_13267);
nor U13997 (N_13997,N_13358,N_13018);
nand U13998 (N_13998,N_13062,N_13349);
or U13999 (N_13999,N_13114,N_13415);
and U14000 (N_14000,N_13559,N_13814);
or U14001 (N_14001,N_13640,N_13514);
xor U14002 (N_14002,N_13733,N_13724);
or U14003 (N_14003,N_13882,N_13885);
nor U14004 (N_14004,N_13741,N_13549);
xnor U14005 (N_14005,N_13795,N_13786);
nor U14006 (N_14006,N_13967,N_13620);
or U14007 (N_14007,N_13747,N_13803);
xor U14008 (N_14008,N_13515,N_13634);
nor U14009 (N_14009,N_13517,N_13956);
xor U14010 (N_14010,N_13766,N_13941);
xnor U14011 (N_14011,N_13966,N_13943);
xnor U14012 (N_14012,N_13571,N_13719);
nand U14013 (N_14013,N_13772,N_13673);
and U14014 (N_14014,N_13561,N_13734);
or U14015 (N_14015,N_13765,N_13849);
nand U14016 (N_14016,N_13763,N_13847);
nand U14017 (N_14017,N_13852,N_13613);
nand U14018 (N_14018,N_13553,N_13540);
nor U14019 (N_14019,N_13607,N_13609);
nor U14020 (N_14020,N_13915,N_13695);
nand U14021 (N_14021,N_13951,N_13608);
nor U14022 (N_14022,N_13659,N_13868);
or U14023 (N_14023,N_13723,N_13937);
xor U14024 (N_14024,N_13787,N_13703);
nor U14025 (N_14025,N_13872,N_13773);
xor U14026 (N_14026,N_13837,N_13715);
nor U14027 (N_14027,N_13925,N_13725);
xnor U14028 (N_14028,N_13648,N_13845);
or U14029 (N_14029,N_13503,N_13644);
nand U14030 (N_14030,N_13611,N_13585);
nor U14031 (N_14031,N_13797,N_13674);
and U14032 (N_14032,N_13886,N_13546);
nand U14033 (N_14033,N_13898,N_13990);
and U14034 (N_14034,N_13657,N_13841);
nand U14035 (N_14035,N_13756,N_13512);
nor U14036 (N_14036,N_13650,N_13744);
xor U14037 (N_14037,N_13743,N_13897);
or U14038 (N_14038,N_13932,N_13740);
nor U14039 (N_14039,N_13813,N_13569);
and U14040 (N_14040,N_13595,N_13796);
nor U14041 (N_14041,N_13697,N_13875);
or U14042 (N_14042,N_13848,N_13881);
xor U14043 (N_14043,N_13537,N_13985);
or U14044 (N_14044,N_13878,N_13738);
nand U14045 (N_14045,N_13963,N_13919);
xor U14046 (N_14046,N_13682,N_13944);
nor U14047 (N_14047,N_13911,N_13928);
xor U14048 (N_14048,N_13891,N_13679);
nand U14049 (N_14049,N_13681,N_13995);
or U14050 (N_14050,N_13606,N_13564);
xor U14051 (N_14051,N_13808,N_13737);
and U14052 (N_14052,N_13989,N_13572);
xor U14053 (N_14053,N_13950,N_13994);
xnor U14054 (N_14054,N_13807,N_13894);
or U14055 (N_14055,N_13711,N_13533);
nand U14056 (N_14056,N_13843,N_13692);
nand U14057 (N_14057,N_13974,N_13834);
nand U14058 (N_14058,N_13570,N_13769);
nand U14059 (N_14059,N_13999,N_13953);
xnor U14060 (N_14060,N_13699,N_13527);
and U14061 (N_14061,N_13577,N_13982);
xor U14062 (N_14062,N_13506,N_13594);
or U14063 (N_14063,N_13730,N_13904);
xor U14064 (N_14064,N_13854,N_13996);
nor U14065 (N_14065,N_13619,N_13819);
or U14066 (N_14066,N_13713,N_13856);
xor U14067 (N_14067,N_13912,N_13525);
nand U14068 (N_14068,N_13568,N_13850);
nor U14069 (N_14069,N_13718,N_13942);
or U14070 (N_14070,N_13866,N_13810);
nor U14071 (N_14071,N_13516,N_13631);
nor U14072 (N_14072,N_13935,N_13597);
and U14073 (N_14073,N_13930,N_13670);
nor U14074 (N_14074,N_13757,N_13579);
and U14075 (N_14075,N_13704,N_13771);
and U14076 (N_14076,N_13663,N_13785);
xor U14077 (N_14077,N_13983,N_13688);
nand U14078 (N_14078,N_13617,N_13920);
nand U14079 (N_14079,N_13789,N_13735);
and U14080 (N_14080,N_13964,N_13705);
or U14081 (N_14081,N_13584,N_13626);
nor U14082 (N_14082,N_13992,N_13507);
nor U14083 (N_14083,N_13957,N_13702);
nor U14084 (N_14084,N_13598,N_13973);
nor U14085 (N_14085,N_13759,N_13804);
and U14086 (N_14086,N_13976,N_13510);
or U14087 (N_14087,N_13625,N_13916);
nor U14088 (N_14088,N_13914,N_13809);
nand U14089 (N_14089,N_13646,N_13633);
nor U14090 (N_14090,N_13940,N_13690);
nand U14091 (N_14091,N_13788,N_13694);
and U14092 (N_14092,N_13861,N_13874);
and U14093 (N_14093,N_13778,N_13538);
or U14094 (N_14094,N_13521,N_13566);
xor U14095 (N_14095,N_13823,N_13767);
or U14096 (N_14096,N_13884,N_13603);
xnor U14097 (N_14097,N_13906,N_13892);
and U14098 (N_14098,N_13600,N_13717);
nand U14099 (N_14099,N_13913,N_13779);
or U14100 (N_14100,N_13574,N_13981);
nor U14101 (N_14101,N_13632,N_13505);
nor U14102 (N_14102,N_13745,N_13641);
or U14103 (N_14103,N_13899,N_13760);
xor U14104 (N_14104,N_13777,N_13858);
or U14105 (N_14105,N_13918,N_13518);
and U14106 (N_14106,N_13700,N_13986);
xnor U14107 (N_14107,N_13980,N_13877);
nor U14108 (N_14108,N_13667,N_13988);
xor U14109 (N_14109,N_13645,N_13621);
nand U14110 (N_14110,N_13931,N_13802);
or U14111 (N_14111,N_13870,N_13658);
nand U14112 (N_14112,N_13839,N_13676);
and U14113 (N_14113,N_13687,N_13817);
xnor U14114 (N_14114,N_13977,N_13820);
xor U14115 (N_14115,N_13954,N_13677);
or U14116 (N_14116,N_13833,N_13909);
or U14117 (N_14117,N_13706,N_13710);
nor U14118 (N_14118,N_13560,N_13601);
nand U14119 (N_14119,N_13895,N_13825);
or U14120 (N_14120,N_13530,N_13851);
nand U14121 (N_14121,N_13927,N_13661);
or U14122 (N_14122,N_13671,N_13519);
or U14123 (N_14123,N_13534,N_13652);
or U14124 (N_14124,N_13592,N_13979);
nor U14125 (N_14125,N_13924,N_13755);
or U14126 (N_14126,N_13933,N_13922);
or U14127 (N_14127,N_13558,N_13869);
nor U14128 (N_14128,N_13548,N_13776);
xnor U14129 (N_14129,N_13751,N_13859);
or U14130 (N_14130,N_13591,N_13831);
or U14131 (N_14131,N_13800,N_13867);
or U14132 (N_14132,N_13666,N_13712);
xnor U14133 (N_14133,N_13949,N_13665);
or U14134 (N_14134,N_13522,N_13655);
nor U14135 (N_14135,N_13707,N_13835);
nand U14136 (N_14136,N_13984,N_13883);
and U14137 (N_14137,N_13509,N_13781);
nand U14138 (N_14138,N_13660,N_13816);
or U14139 (N_14139,N_13962,N_13552);
or U14140 (N_14140,N_13902,N_13997);
nand U14141 (N_14141,N_13955,N_13536);
or U14142 (N_14142,N_13524,N_13582);
nor U14143 (N_14143,N_13578,N_13589);
nand U14144 (N_14144,N_13840,N_13562);
nand U14145 (N_14145,N_13588,N_13727);
and U14146 (N_14146,N_13969,N_13936);
nand U14147 (N_14147,N_13716,N_13535);
and U14148 (N_14148,N_13662,N_13836);
xnor U14149 (N_14149,N_13624,N_13921);
nor U14150 (N_14150,N_13701,N_13978);
or U14151 (N_14151,N_13842,N_13547);
nor U14152 (N_14152,N_13907,N_13871);
and U14153 (N_14153,N_13961,N_13637);
xnor U14154 (N_14154,N_13770,N_13822);
or U14155 (N_14155,N_13541,N_13513);
and U14156 (N_14156,N_13815,N_13627);
nor U14157 (N_14157,N_13952,N_13501);
or U14158 (N_14158,N_13853,N_13764);
xnor U14159 (N_14159,N_13565,N_13708);
nor U14160 (N_14160,N_13615,N_13805);
xor U14161 (N_14161,N_13829,N_13998);
or U14162 (N_14162,N_13722,N_13946);
xor U14163 (N_14163,N_13623,N_13864);
xor U14164 (N_14164,N_13714,N_13605);
or U14165 (N_14165,N_13865,N_13523);
nor U14166 (N_14166,N_13780,N_13531);
nor U14167 (N_14167,N_13680,N_13968);
xnor U14168 (N_14168,N_13910,N_13826);
and U14169 (N_14169,N_13654,N_13970);
or U14170 (N_14170,N_13664,N_13618);
and U14171 (N_14171,N_13502,N_13721);
or U14172 (N_14172,N_13635,N_13567);
nand U14173 (N_14173,N_13614,N_13539);
xnor U14174 (N_14174,N_13542,N_13873);
nand U14175 (N_14175,N_13855,N_13846);
or U14176 (N_14176,N_13862,N_13917);
and U14177 (N_14177,N_13678,N_13732);
nor U14178 (N_14178,N_13901,N_13728);
xor U14179 (N_14179,N_13975,N_13726);
or U14180 (N_14180,N_13758,N_13739);
or U14181 (N_14181,N_13684,N_13528);
and U14182 (N_14182,N_13863,N_13812);
xnor U14183 (N_14183,N_13628,N_13581);
nor U14184 (N_14184,N_13573,N_13551);
nor U14185 (N_14185,N_13971,N_13508);
nand U14186 (N_14186,N_13934,N_13599);
xnor U14187 (N_14187,N_13500,N_13742);
nand U14188 (N_14188,N_13782,N_13750);
xor U14189 (N_14189,N_13557,N_13686);
or U14190 (N_14190,N_13900,N_13889);
xnor U14191 (N_14191,N_13746,N_13749);
xnor U14192 (N_14192,N_13791,N_13576);
xnor U14193 (N_14193,N_13799,N_13811);
nand U14194 (N_14194,N_13556,N_13893);
or U14195 (N_14195,N_13587,N_13783);
nor U14196 (N_14196,N_13689,N_13938);
xor U14197 (N_14197,N_13948,N_13563);
nand U14198 (N_14198,N_13923,N_13575);
nand U14199 (N_14199,N_13801,N_13880);
or U14200 (N_14200,N_13643,N_13896);
xnor U14201 (N_14201,N_13959,N_13602);
and U14202 (N_14202,N_13775,N_13798);
nand U14203 (N_14203,N_13642,N_13555);
nand U14204 (N_14204,N_13554,N_13720);
nor U14205 (N_14205,N_13832,N_13668);
nor U14206 (N_14206,N_13693,N_13532);
nand U14207 (N_14207,N_13731,N_13806);
nor U14208 (N_14208,N_13818,N_13736);
xnor U14209 (N_14209,N_13972,N_13698);
nor U14210 (N_14210,N_13821,N_13672);
xor U14211 (N_14211,N_13926,N_13748);
and U14212 (N_14212,N_13939,N_13753);
xnor U14213 (N_14213,N_13543,N_13794);
or U14214 (N_14214,N_13828,N_13890);
or U14215 (N_14215,N_13685,N_13593);
and U14216 (N_14216,N_13958,N_13622);
or U14217 (N_14217,N_13929,N_13649);
nor U14218 (N_14218,N_13544,N_13529);
and U14219 (N_14219,N_13857,N_13630);
or U14220 (N_14220,N_13887,N_13792);
or U14221 (N_14221,N_13669,N_13586);
or U14222 (N_14222,N_13691,N_13653);
or U14223 (N_14223,N_13590,N_13656);
or U14224 (N_14224,N_13504,N_13675);
nor U14225 (N_14225,N_13639,N_13762);
nand U14226 (N_14226,N_13784,N_13824);
or U14227 (N_14227,N_13638,N_13888);
xor U14228 (N_14228,N_13830,N_13696);
or U14229 (N_14229,N_13604,N_13987);
nand U14230 (N_14230,N_13729,N_13754);
nand U14231 (N_14231,N_13761,N_13752);
or U14232 (N_14232,N_13879,N_13793);
and U14233 (N_14233,N_13647,N_13860);
xor U14234 (N_14234,N_13960,N_13629);
nor U14235 (N_14235,N_13550,N_13827);
or U14236 (N_14236,N_13636,N_13768);
or U14237 (N_14237,N_13526,N_13965);
nor U14238 (N_14238,N_13616,N_13596);
and U14239 (N_14239,N_13580,N_13947);
or U14240 (N_14240,N_13683,N_13838);
nand U14241 (N_14241,N_13651,N_13520);
nor U14242 (N_14242,N_13583,N_13908);
and U14243 (N_14243,N_13991,N_13945);
and U14244 (N_14244,N_13844,N_13610);
nand U14245 (N_14245,N_13511,N_13709);
xnor U14246 (N_14246,N_13993,N_13612);
xor U14247 (N_14247,N_13545,N_13903);
nand U14248 (N_14248,N_13876,N_13905);
and U14249 (N_14249,N_13790,N_13774);
nor U14250 (N_14250,N_13814,N_13748);
or U14251 (N_14251,N_13987,N_13888);
xnor U14252 (N_14252,N_13612,N_13592);
and U14253 (N_14253,N_13707,N_13922);
nand U14254 (N_14254,N_13876,N_13547);
and U14255 (N_14255,N_13959,N_13965);
nand U14256 (N_14256,N_13738,N_13721);
or U14257 (N_14257,N_13931,N_13638);
or U14258 (N_14258,N_13729,N_13680);
nand U14259 (N_14259,N_13813,N_13711);
xnor U14260 (N_14260,N_13624,N_13662);
nand U14261 (N_14261,N_13852,N_13976);
nand U14262 (N_14262,N_13982,N_13858);
or U14263 (N_14263,N_13865,N_13601);
nand U14264 (N_14264,N_13781,N_13701);
nor U14265 (N_14265,N_13595,N_13930);
nor U14266 (N_14266,N_13867,N_13720);
nand U14267 (N_14267,N_13694,N_13614);
xnor U14268 (N_14268,N_13647,N_13676);
and U14269 (N_14269,N_13887,N_13943);
or U14270 (N_14270,N_13655,N_13928);
or U14271 (N_14271,N_13970,N_13524);
or U14272 (N_14272,N_13899,N_13989);
xnor U14273 (N_14273,N_13689,N_13736);
nor U14274 (N_14274,N_13526,N_13775);
and U14275 (N_14275,N_13549,N_13668);
and U14276 (N_14276,N_13708,N_13501);
nor U14277 (N_14277,N_13663,N_13887);
nand U14278 (N_14278,N_13515,N_13854);
and U14279 (N_14279,N_13646,N_13759);
and U14280 (N_14280,N_13813,N_13641);
or U14281 (N_14281,N_13687,N_13937);
or U14282 (N_14282,N_13501,N_13844);
or U14283 (N_14283,N_13802,N_13673);
nand U14284 (N_14284,N_13593,N_13948);
xnor U14285 (N_14285,N_13565,N_13951);
and U14286 (N_14286,N_13781,N_13619);
or U14287 (N_14287,N_13963,N_13711);
xnor U14288 (N_14288,N_13698,N_13732);
nor U14289 (N_14289,N_13610,N_13986);
and U14290 (N_14290,N_13667,N_13629);
or U14291 (N_14291,N_13724,N_13723);
or U14292 (N_14292,N_13941,N_13818);
or U14293 (N_14293,N_13583,N_13890);
nor U14294 (N_14294,N_13970,N_13504);
xnor U14295 (N_14295,N_13665,N_13688);
nor U14296 (N_14296,N_13942,N_13561);
nor U14297 (N_14297,N_13711,N_13838);
or U14298 (N_14298,N_13514,N_13625);
or U14299 (N_14299,N_13657,N_13713);
nor U14300 (N_14300,N_13884,N_13952);
and U14301 (N_14301,N_13579,N_13541);
and U14302 (N_14302,N_13582,N_13998);
nand U14303 (N_14303,N_13993,N_13947);
xor U14304 (N_14304,N_13683,N_13512);
xor U14305 (N_14305,N_13807,N_13799);
xor U14306 (N_14306,N_13606,N_13521);
xnor U14307 (N_14307,N_13591,N_13566);
xnor U14308 (N_14308,N_13606,N_13737);
nor U14309 (N_14309,N_13570,N_13521);
and U14310 (N_14310,N_13926,N_13634);
or U14311 (N_14311,N_13691,N_13707);
xor U14312 (N_14312,N_13822,N_13941);
nand U14313 (N_14313,N_13818,N_13509);
and U14314 (N_14314,N_13864,N_13752);
xor U14315 (N_14315,N_13863,N_13716);
or U14316 (N_14316,N_13744,N_13700);
or U14317 (N_14317,N_13639,N_13815);
nor U14318 (N_14318,N_13614,N_13941);
xnor U14319 (N_14319,N_13802,N_13730);
nand U14320 (N_14320,N_13787,N_13939);
nand U14321 (N_14321,N_13718,N_13890);
and U14322 (N_14322,N_13846,N_13789);
and U14323 (N_14323,N_13638,N_13881);
or U14324 (N_14324,N_13934,N_13639);
and U14325 (N_14325,N_13557,N_13722);
xnor U14326 (N_14326,N_13971,N_13868);
or U14327 (N_14327,N_13916,N_13537);
and U14328 (N_14328,N_13833,N_13704);
or U14329 (N_14329,N_13563,N_13638);
nor U14330 (N_14330,N_13845,N_13628);
nand U14331 (N_14331,N_13953,N_13679);
xnor U14332 (N_14332,N_13594,N_13658);
and U14333 (N_14333,N_13516,N_13959);
xnor U14334 (N_14334,N_13623,N_13867);
nor U14335 (N_14335,N_13858,N_13928);
or U14336 (N_14336,N_13814,N_13885);
or U14337 (N_14337,N_13626,N_13572);
xor U14338 (N_14338,N_13875,N_13669);
and U14339 (N_14339,N_13606,N_13617);
or U14340 (N_14340,N_13772,N_13691);
or U14341 (N_14341,N_13733,N_13576);
nand U14342 (N_14342,N_13566,N_13836);
and U14343 (N_14343,N_13866,N_13614);
and U14344 (N_14344,N_13884,N_13843);
nand U14345 (N_14345,N_13586,N_13652);
nand U14346 (N_14346,N_13813,N_13603);
or U14347 (N_14347,N_13822,N_13969);
nand U14348 (N_14348,N_13695,N_13855);
xnor U14349 (N_14349,N_13760,N_13765);
nor U14350 (N_14350,N_13896,N_13670);
nor U14351 (N_14351,N_13600,N_13931);
xnor U14352 (N_14352,N_13504,N_13952);
nor U14353 (N_14353,N_13712,N_13652);
nand U14354 (N_14354,N_13672,N_13777);
nand U14355 (N_14355,N_13644,N_13637);
or U14356 (N_14356,N_13595,N_13902);
nor U14357 (N_14357,N_13806,N_13543);
or U14358 (N_14358,N_13987,N_13862);
or U14359 (N_14359,N_13714,N_13675);
nand U14360 (N_14360,N_13969,N_13536);
nor U14361 (N_14361,N_13883,N_13572);
and U14362 (N_14362,N_13725,N_13529);
nor U14363 (N_14363,N_13777,N_13874);
nand U14364 (N_14364,N_13817,N_13905);
nand U14365 (N_14365,N_13742,N_13805);
nand U14366 (N_14366,N_13818,N_13651);
nor U14367 (N_14367,N_13706,N_13751);
xnor U14368 (N_14368,N_13792,N_13611);
xnor U14369 (N_14369,N_13560,N_13914);
and U14370 (N_14370,N_13868,N_13946);
nand U14371 (N_14371,N_13603,N_13664);
nor U14372 (N_14372,N_13508,N_13597);
and U14373 (N_14373,N_13734,N_13950);
xor U14374 (N_14374,N_13576,N_13785);
nand U14375 (N_14375,N_13916,N_13635);
or U14376 (N_14376,N_13609,N_13808);
nand U14377 (N_14377,N_13517,N_13664);
nand U14378 (N_14378,N_13521,N_13534);
nor U14379 (N_14379,N_13834,N_13746);
and U14380 (N_14380,N_13860,N_13792);
nor U14381 (N_14381,N_13828,N_13887);
or U14382 (N_14382,N_13716,N_13531);
or U14383 (N_14383,N_13560,N_13643);
nor U14384 (N_14384,N_13544,N_13872);
and U14385 (N_14385,N_13894,N_13649);
nand U14386 (N_14386,N_13541,N_13999);
xnor U14387 (N_14387,N_13676,N_13905);
nand U14388 (N_14388,N_13986,N_13892);
xnor U14389 (N_14389,N_13802,N_13670);
nand U14390 (N_14390,N_13966,N_13892);
xor U14391 (N_14391,N_13890,N_13615);
and U14392 (N_14392,N_13917,N_13645);
xor U14393 (N_14393,N_13695,N_13994);
nand U14394 (N_14394,N_13506,N_13641);
xor U14395 (N_14395,N_13582,N_13532);
or U14396 (N_14396,N_13716,N_13503);
nand U14397 (N_14397,N_13758,N_13703);
or U14398 (N_14398,N_13557,N_13574);
nand U14399 (N_14399,N_13504,N_13968);
xor U14400 (N_14400,N_13526,N_13688);
or U14401 (N_14401,N_13615,N_13753);
nor U14402 (N_14402,N_13912,N_13904);
nor U14403 (N_14403,N_13828,N_13868);
nand U14404 (N_14404,N_13662,N_13564);
and U14405 (N_14405,N_13505,N_13553);
nand U14406 (N_14406,N_13812,N_13922);
and U14407 (N_14407,N_13955,N_13788);
xor U14408 (N_14408,N_13729,N_13632);
or U14409 (N_14409,N_13660,N_13832);
nor U14410 (N_14410,N_13802,N_13743);
and U14411 (N_14411,N_13849,N_13943);
xnor U14412 (N_14412,N_13501,N_13965);
xor U14413 (N_14413,N_13679,N_13651);
xor U14414 (N_14414,N_13732,N_13757);
nand U14415 (N_14415,N_13602,N_13670);
or U14416 (N_14416,N_13682,N_13598);
nand U14417 (N_14417,N_13749,N_13909);
or U14418 (N_14418,N_13755,N_13852);
xnor U14419 (N_14419,N_13960,N_13530);
and U14420 (N_14420,N_13902,N_13832);
nor U14421 (N_14421,N_13754,N_13762);
or U14422 (N_14422,N_13819,N_13548);
and U14423 (N_14423,N_13730,N_13932);
and U14424 (N_14424,N_13527,N_13829);
nand U14425 (N_14425,N_13919,N_13905);
xor U14426 (N_14426,N_13879,N_13997);
or U14427 (N_14427,N_13753,N_13917);
nor U14428 (N_14428,N_13691,N_13690);
and U14429 (N_14429,N_13806,N_13981);
nand U14430 (N_14430,N_13571,N_13658);
nor U14431 (N_14431,N_13990,N_13722);
xnor U14432 (N_14432,N_13746,N_13677);
xnor U14433 (N_14433,N_13776,N_13847);
nand U14434 (N_14434,N_13835,N_13896);
or U14435 (N_14435,N_13842,N_13527);
xnor U14436 (N_14436,N_13752,N_13591);
nand U14437 (N_14437,N_13732,N_13565);
nor U14438 (N_14438,N_13948,N_13866);
and U14439 (N_14439,N_13708,N_13750);
and U14440 (N_14440,N_13684,N_13679);
nor U14441 (N_14441,N_13826,N_13913);
and U14442 (N_14442,N_13595,N_13897);
or U14443 (N_14443,N_13563,N_13920);
or U14444 (N_14444,N_13782,N_13821);
xor U14445 (N_14445,N_13968,N_13635);
nand U14446 (N_14446,N_13735,N_13947);
and U14447 (N_14447,N_13895,N_13785);
nor U14448 (N_14448,N_13510,N_13612);
nor U14449 (N_14449,N_13947,N_13825);
xor U14450 (N_14450,N_13521,N_13879);
nor U14451 (N_14451,N_13981,N_13614);
nor U14452 (N_14452,N_13824,N_13698);
or U14453 (N_14453,N_13964,N_13788);
and U14454 (N_14454,N_13823,N_13518);
and U14455 (N_14455,N_13798,N_13885);
or U14456 (N_14456,N_13512,N_13948);
xor U14457 (N_14457,N_13754,N_13950);
nand U14458 (N_14458,N_13983,N_13995);
or U14459 (N_14459,N_13868,N_13564);
and U14460 (N_14460,N_13581,N_13903);
xnor U14461 (N_14461,N_13540,N_13935);
nor U14462 (N_14462,N_13913,N_13851);
and U14463 (N_14463,N_13993,N_13941);
or U14464 (N_14464,N_13576,N_13655);
and U14465 (N_14465,N_13537,N_13519);
nor U14466 (N_14466,N_13757,N_13867);
and U14467 (N_14467,N_13541,N_13823);
xnor U14468 (N_14468,N_13592,N_13918);
xor U14469 (N_14469,N_13971,N_13967);
xnor U14470 (N_14470,N_13974,N_13576);
and U14471 (N_14471,N_13765,N_13939);
and U14472 (N_14472,N_13585,N_13828);
xor U14473 (N_14473,N_13869,N_13549);
and U14474 (N_14474,N_13682,N_13524);
nand U14475 (N_14475,N_13828,N_13937);
or U14476 (N_14476,N_13526,N_13808);
and U14477 (N_14477,N_13629,N_13718);
or U14478 (N_14478,N_13943,N_13547);
and U14479 (N_14479,N_13700,N_13616);
or U14480 (N_14480,N_13704,N_13756);
nand U14481 (N_14481,N_13529,N_13696);
xor U14482 (N_14482,N_13918,N_13688);
nor U14483 (N_14483,N_13762,N_13575);
and U14484 (N_14484,N_13570,N_13696);
nand U14485 (N_14485,N_13888,N_13934);
nor U14486 (N_14486,N_13585,N_13980);
and U14487 (N_14487,N_13662,N_13813);
xnor U14488 (N_14488,N_13624,N_13717);
and U14489 (N_14489,N_13684,N_13672);
xnor U14490 (N_14490,N_13937,N_13836);
and U14491 (N_14491,N_13865,N_13510);
xor U14492 (N_14492,N_13534,N_13969);
nand U14493 (N_14493,N_13509,N_13668);
nand U14494 (N_14494,N_13953,N_13793);
nor U14495 (N_14495,N_13893,N_13725);
and U14496 (N_14496,N_13517,N_13791);
or U14497 (N_14497,N_13914,N_13551);
or U14498 (N_14498,N_13675,N_13640);
xnor U14499 (N_14499,N_13959,N_13542);
xor U14500 (N_14500,N_14176,N_14357);
nor U14501 (N_14501,N_14165,N_14474);
xnor U14502 (N_14502,N_14461,N_14154);
nand U14503 (N_14503,N_14393,N_14462);
nand U14504 (N_14504,N_14382,N_14226);
or U14505 (N_14505,N_14005,N_14374);
nand U14506 (N_14506,N_14373,N_14481);
xor U14507 (N_14507,N_14213,N_14451);
xnor U14508 (N_14508,N_14122,N_14046);
nand U14509 (N_14509,N_14204,N_14289);
nand U14510 (N_14510,N_14208,N_14110);
nand U14511 (N_14511,N_14259,N_14116);
nor U14512 (N_14512,N_14106,N_14210);
xor U14513 (N_14513,N_14004,N_14124);
nor U14514 (N_14514,N_14083,N_14491);
nand U14515 (N_14515,N_14472,N_14159);
nand U14516 (N_14516,N_14153,N_14034);
nor U14517 (N_14517,N_14407,N_14042);
and U14518 (N_14518,N_14460,N_14478);
nor U14519 (N_14519,N_14001,N_14468);
or U14520 (N_14520,N_14172,N_14211);
and U14521 (N_14521,N_14156,N_14011);
or U14522 (N_14522,N_14000,N_14418);
or U14523 (N_14523,N_14182,N_14168);
xnor U14524 (N_14524,N_14169,N_14383);
or U14525 (N_14525,N_14400,N_14246);
and U14526 (N_14526,N_14063,N_14184);
nor U14527 (N_14527,N_14024,N_14055);
xnor U14528 (N_14528,N_14157,N_14194);
xor U14529 (N_14529,N_14343,N_14043);
or U14530 (N_14530,N_14327,N_14079);
or U14531 (N_14531,N_14466,N_14145);
nand U14532 (N_14532,N_14359,N_14173);
nor U14533 (N_14533,N_14037,N_14198);
or U14534 (N_14534,N_14085,N_14251);
xnor U14535 (N_14535,N_14202,N_14264);
xor U14536 (N_14536,N_14445,N_14261);
nand U14537 (N_14537,N_14127,N_14052);
xor U14538 (N_14538,N_14488,N_14290);
nor U14539 (N_14539,N_14314,N_14199);
and U14540 (N_14540,N_14029,N_14412);
nor U14541 (N_14541,N_14152,N_14298);
and U14542 (N_14542,N_14395,N_14447);
nor U14543 (N_14543,N_14433,N_14014);
and U14544 (N_14544,N_14380,N_14022);
or U14545 (N_14545,N_14392,N_14366);
nor U14546 (N_14546,N_14054,N_14084);
nor U14547 (N_14547,N_14178,N_14446);
nand U14548 (N_14548,N_14128,N_14015);
nand U14549 (N_14549,N_14492,N_14185);
and U14550 (N_14550,N_14267,N_14317);
nor U14551 (N_14551,N_14191,N_14077);
and U14552 (N_14552,N_14249,N_14436);
nor U14553 (N_14553,N_14097,N_14006);
or U14554 (N_14554,N_14041,N_14448);
and U14555 (N_14555,N_14379,N_14295);
or U14556 (N_14556,N_14170,N_14039);
xor U14557 (N_14557,N_14354,N_14435);
nor U14558 (N_14558,N_14019,N_14141);
and U14559 (N_14559,N_14214,N_14140);
nor U14560 (N_14560,N_14434,N_14403);
or U14561 (N_14561,N_14020,N_14377);
or U14562 (N_14562,N_14269,N_14038);
and U14563 (N_14563,N_14364,N_14371);
xor U14564 (N_14564,N_14304,N_14121);
and U14565 (N_14565,N_14483,N_14337);
and U14566 (N_14566,N_14088,N_14078);
and U14567 (N_14567,N_14353,N_14427);
and U14568 (N_14568,N_14231,N_14081);
xnor U14569 (N_14569,N_14254,N_14033);
and U14570 (N_14570,N_14013,N_14316);
or U14571 (N_14571,N_14312,N_14397);
nor U14572 (N_14572,N_14209,N_14135);
xor U14573 (N_14573,N_14477,N_14007);
or U14574 (N_14574,N_14224,N_14040);
xnor U14575 (N_14575,N_14256,N_14283);
nor U14576 (N_14576,N_14248,N_14469);
or U14577 (N_14577,N_14296,N_14134);
xnor U14578 (N_14578,N_14411,N_14347);
or U14579 (N_14579,N_14105,N_14094);
or U14580 (N_14580,N_14370,N_14276);
or U14581 (N_14581,N_14457,N_14413);
or U14582 (N_14582,N_14167,N_14160);
nand U14583 (N_14583,N_14130,N_14257);
or U14584 (N_14584,N_14439,N_14238);
or U14585 (N_14585,N_14069,N_14301);
nand U14586 (N_14586,N_14220,N_14480);
nor U14587 (N_14587,N_14234,N_14240);
and U14588 (N_14588,N_14065,N_14355);
or U14589 (N_14589,N_14203,N_14268);
nand U14590 (N_14590,N_14287,N_14422);
and U14591 (N_14591,N_14036,N_14440);
nand U14592 (N_14592,N_14023,N_14426);
nand U14593 (N_14593,N_14300,N_14225);
and U14594 (N_14594,N_14281,N_14074);
xnor U14595 (N_14595,N_14275,N_14454);
xnor U14596 (N_14596,N_14060,N_14095);
nor U14597 (N_14597,N_14260,N_14216);
and U14598 (N_14598,N_14093,N_14311);
or U14599 (N_14599,N_14344,N_14218);
xnor U14600 (N_14600,N_14284,N_14192);
or U14601 (N_14601,N_14262,N_14401);
and U14602 (N_14602,N_14297,N_14193);
xnor U14603 (N_14603,N_14201,N_14200);
xor U14604 (N_14604,N_14319,N_14086);
or U14605 (N_14605,N_14385,N_14187);
nor U14606 (N_14606,N_14306,N_14294);
xnor U14607 (N_14607,N_14072,N_14358);
and U14608 (N_14608,N_14195,N_14367);
and U14609 (N_14609,N_14258,N_14067);
xnor U14610 (N_14610,N_14100,N_14498);
nor U14611 (N_14611,N_14031,N_14372);
and U14612 (N_14612,N_14028,N_14292);
and U14613 (N_14613,N_14365,N_14414);
xor U14614 (N_14614,N_14188,N_14302);
or U14615 (N_14615,N_14270,N_14009);
xnor U14616 (N_14616,N_14142,N_14099);
xor U14617 (N_14617,N_14008,N_14323);
or U14618 (N_14618,N_14431,N_14408);
and U14619 (N_14619,N_14398,N_14386);
nor U14620 (N_14620,N_14227,N_14326);
or U14621 (N_14621,N_14125,N_14215);
xnor U14622 (N_14622,N_14376,N_14189);
nor U14623 (N_14623,N_14423,N_14420);
and U14624 (N_14624,N_14114,N_14274);
nor U14625 (N_14625,N_14070,N_14277);
nand U14626 (N_14626,N_14123,N_14010);
or U14627 (N_14627,N_14387,N_14155);
or U14628 (N_14628,N_14432,N_14493);
nor U14629 (N_14629,N_14098,N_14437);
nand U14630 (N_14630,N_14351,N_14416);
xnor U14631 (N_14631,N_14456,N_14196);
or U14632 (N_14632,N_14244,N_14239);
or U14633 (N_14633,N_14402,N_14450);
or U14634 (N_14634,N_14126,N_14050);
nor U14635 (N_14635,N_14349,N_14051);
nand U14636 (N_14636,N_14368,N_14320);
and U14637 (N_14637,N_14489,N_14285);
xnor U14638 (N_14638,N_14229,N_14279);
nor U14639 (N_14639,N_14162,N_14151);
or U14640 (N_14640,N_14419,N_14047);
nand U14641 (N_14641,N_14104,N_14305);
nand U14642 (N_14642,N_14035,N_14076);
nor U14643 (N_14643,N_14389,N_14045);
and U14644 (N_14644,N_14499,N_14137);
and U14645 (N_14645,N_14356,N_14465);
or U14646 (N_14646,N_14363,N_14092);
nor U14647 (N_14647,N_14186,N_14241);
xor U14648 (N_14648,N_14495,N_14091);
and U14649 (N_14649,N_14205,N_14181);
or U14650 (N_14650,N_14061,N_14496);
xnor U14651 (N_14651,N_14293,N_14266);
xor U14652 (N_14652,N_14223,N_14391);
nand U14653 (N_14653,N_14062,N_14321);
and U14654 (N_14654,N_14146,N_14307);
and U14655 (N_14655,N_14102,N_14073);
or U14656 (N_14656,N_14332,N_14149);
or U14657 (N_14657,N_14421,N_14059);
nor U14658 (N_14658,N_14222,N_14103);
xnor U14659 (N_14659,N_14232,N_14441);
nor U14660 (N_14660,N_14030,N_14280);
xor U14661 (N_14661,N_14161,N_14330);
xor U14662 (N_14662,N_14303,N_14068);
or U14663 (N_14663,N_14464,N_14291);
or U14664 (N_14664,N_14331,N_14115);
xor U14665 (N_14665,N_14396,N_14053);
nand U14666 (N_14666,N_14406,N_14082);
or U14667 (N_14667,N_14453,N_14324);
xor U14668 (N_14668,N_14404,N_14148);
nand U14669 (N_14669,N_14475,N_14230);
xnor U14670 (N_14670,N_14417,N_14117);
xnor U14671 (N_14671,N_14428,N_14443);
and U14672 (N_14672,N_14263,N_14335);
xnor U14673 (N_14673,N_14113,N_14096);
nor U14674 (N_14674,N_14197,N_14075);
nand U14675 (N_14675,N_14144,N_14057);
xor U14676 (N_14676,N_14228,N_14452);
or U14677 (N_14677,N_14243,N_14012);
and U14678 (N_14678,N_14252,N_14473);
nand U14679 (N_14679,N_14424,N_14470);
xor U14680 (N_14680,N_14490,N_14265);
xor U14681 (N_14681,N_14484,N_14415);
and U14682 (N_14682,N_14107,N_14467);
or U14683 (N_14683,N_14438,N_14345);
and U14684 (N_14684,N_14147,N_14342);
nor U14685 (N_14685,N_14026,N_14299);
nand U14686 (N_14686,N_14044,N_14494);
or U14687 (N_14687,N_14136,N_14339);
xor U14688 (N_14688,N_14410,N_14390);
nand U14689 (N_14689,N_14212,N_14139);
xnor U14690 (N_14690,N_14058,N_14245);
and U14691 (N_14691,N_14272,N_14325);
or U14692 (N_14692,N_14190,N_14017);
nor U14693 (N_14693,N_14338,N_14233);
and U14694 (N_14694,N_14497,N_14487);
and U14695 (N_14695,N_14361,N_14378);
xor U14696 (N_14696,N_14449,N_14180);
xor U14697 (N_14697,N_14064,N_14164);
nor U14698 (N_14698,N_14341,N_14219);
xor U14699 (N_14699,N_14278,N_14177);
nand U14700 (N_14700,N_14025,N_14352);
or U14701 (N_14701,N_14112,N_14032);
nand U14702 (N_14702,N_14087,N_14131);
and U14703 (N_14703,N_14056,N_14308);
or U14704 (N_14704,N_14409,N_14333);
or U14705 (N_14705,N_14340,N_14016);
and U14706 (N_14706,N_14425,N_14089);
or U14707 (N_14707,N_14271,N_14369);
nand U14708 (N_14708,N_14348,N_14049);
nand U14709 (N_14709,N_14236,N_14071);
and U14710 (N_14710,N_14207,N_14111);
and U14711 (N_14711,N_14101,N_14255);
nand U14712 (N_14712,N_14129,N_14090);
nand U14713 (N_14713,N_14381,N_14150);
nand U14714 (N_14714,N_14179,N_14021);
nor U14715 (N_14715,N_14118,N_14166);
xnor U14716 (N_14716,N_14444,N_14171);
nand U14717 (N_14717,N_14458,N_14429);
nand U14718 (N_14718,N_14328,N_14206);
nand U14719 (N_14719,N_14322,N_14318);
or U14720 (N_14720,N_14399,N_14003);
xor U14721 (N_14721,N_14430,N_14388);
and U14722 (N_14722,N_14242,N_14138);
and U14723 (N_14723,N_14235,N_14108);
xnor U14724 (N_14724,N_14486,N_14217);
or U14725 (N_14725,N_14336,N_14018);
or U14726 (N_14726,N_14384,N_14253);
nor U14727 (N_14727,N_14334,N_14313);
or U14728 (N_14728,N_14066,N_14350);
and U14729 (N_14729,N_14247,N_14309);
nand U14730 (N_14730,N_14476,N_14288);
nor U14731 (N_14731,N_14482,N_14237);
nor U14732 (N_14732,N_14375,N_14479);
nand U14733 (N_14733,N_14471,N_14174);
nor U14734 (N_14734,N_14315,N_14329);
or U14735 (N_14735,N_14459,N_14080);
xor U14736 (N_14736,N_14394,N_14463);
or U14737 (N_14737,N_14163,N_14109);
or U14738 (N_14738,N_14048,N_14143);
or U14739 (N_14739,N_14175,N_14362);
or U14740 (N_14740,N_14286,N_14442);
or U14741 (N_14741,N_14132,N_14405);
xor U14742 (N_14742,N_14183,N_14120);
and U14743 (N_14743,N_14119,N_14455);
xnor U14744 (N_14744,N_14221,N_14282);
or U14745 (N_14745,N_14133,N_14027);
and U14746 (N_14746,N_14273,N_14310);
or U14747 (N_14747,N_14002,N_14158);
nand U14748 (N_14748,N_14485,N_14346);
or U14749 (N_14749,N_14250,N_14360);
nor U14750 (N_14750,N_14423,N_14347);
nand U14751 (N_14751,N_14322,N_14344);
nor U14752 (N_14752,N_14330,N_14461);
nor U14753 (N_14753,N_14284,N_14135);
or U14754 (N_14754,N_14225,N_14373);
nor U14755 (N_14755,N_14448,N_14158);
nand U14756 (N_14756,N_14119,N_14245);
xor U14757 (N_14757,N_14123,N_14100);
nand U14758 (N_14758,N_14353,N_14483);
nand U14759 (N_14759,N_14234,N_14028);
nand U14760 (N_14760,N_14089,N_14409);
and U14761 (N_14761,N_14259,N_14372);
or U14762 (N_14762,N_14130,N_14387);
or U14763 (N_14763,N_14134,N_14408);
or U14764 (N_14764,N_14047,N_14319);
xnor U14765 (N_14765,N_14321,N_14056);
and U14766 (N_14766,N_14416,N_14205);
nand U14767 (N_14767,N_14232,N_14319);
nor U14768 (N_14768,N_14044,N_14066);
nor U14769 (N_14769,N_14315,N_14272);
nor U14770 (N_14770,N_14263,N_14090);
xor U14771 (N_14771,N_14326,N_14324);
nand U14772 (N_14772,N_14102,N_14135);
xnor U14773 (N_14773,N_14099,N_14486);
nand U14774 (N_14774,N_14320,N_14081);
nor U14775 (N_14775,N_14160,N_14036);
xor U14776 (N_14776,N_14491,N_14259);
nor U14777 (N_14777,N_14186,N_14360);
or U14778 (N_14778,N_14495,N_14032);
nand U14779 (N_14779,N_14274,N_14030);
or U14780 (N_14780,N_14132,N_14114);
or U14781 (N_14781,N_14261,N_14040);
xnor U14782 (N_14782,N_14202,N_14493);
xor U14783 (N_14783,N_14180,N_14136);
and U14784 (N_14784,N_14458,N_14273);
or U14785 (N_14785,N_14427,N_14100);
nand U14786 (N_14786,N_14199,N_14379);
nor U14787 (N_14787,N_14395,N_14398);
nor U14788 (N_14788,N_14246,N_14370);
nor U14789 (N_14789,N_14403,N_14144);
and U14790 (N_14790,N_14454,N_14083);
or U14791 (N_14791,N_14320,N_14337);
or U14792 (N_14792,N_14490,N_14206);
nor U14793 (N_14793,N_14075,N_14420);
or U14794 (N_14794,N_14424,N_14126);
or U14795 (N_14795,N_14453,N_14286);
nand U14796 (N_14796,N_14047,N_14375);
nand U14797 (N_14797,N_14056,N_14063);
nand U14798 (N_14798,N_14061,N_14398);
nor U14799 (N_14799,N_14119,N_14109);
nand U14800 (N_14800,N_14273,N_14194);
or U14801 (N_14801,N_14346,N_14081);
or U14802 (N_14802,N_14081,N_14026);
xnor U14803 (N_14803,N_14037,N_14005);
and U14804 (N_14804,N_14491,N_14049);
nor U14805 (N_14805,N_14407,N_14270);
nor U14806 (N_14806,N_14049,N_14343);
nor U14807 (N_14807,N_14205,N_14459);
and U14808 (N_14808,N_14358,N_14429);
nor U14809 (N_14809,N_14253,N_14233);
xor U14810 (N_14810,N_14349,N_14110);
nand U14811 (N_14811,N_14147,N_14473);
nor U14812 (N_14812,N_14156,N_14054);
and U14813 (N_14813,N_14419,N_14207);
xnor U14814 (N_14814,N_14488,N_14351);
nand U14815 (N_14815,N_14071,N_14102);
or U14816 (N_14816,N_14461,N_14365);
or U14817 (N_14817,N_14208,N_14076);
or U14818 (N_14818,N_14106,N_14425);
nand U14819 (N_14819,N_14191,N_14497);
or U14820 (N_14820,N_14402,N_14094);
nor U14821 (N_14821,N_14133,N_14412);
nand U14822 (N_14822,N_14262,N_14041);
nand U14823 (N_14823,N_14253,N_14245);
or U14824 (N_14824,N_14364,N_14490);
and U14825 (N_14825,N_14397,N_14348);
nand U14826 (N_14826,N_14331,N_14204);
or U14827 (N_14827,N_14088,N_14085);
nand U14828 (N_14828,N_14447,N_14164);
nor U14829 (N_14829,N_14084,N_14125);
nand U14830 (N_14830,N_14250,N_14097);
and U14831 (N_14831,N_14055,N_14057);
xor U14832 (N_14832,N_14240,N_14445);
or U14833 (N_14833,N_14262,N_14456);
xor U14834 (N_14834,N_14343,N_14389);
xor U14835 (N_14835,N_14210,N_14396);
and U14836 (N_14836,N_14292,N_14077);
and U14837 (N_14837,N_14164,N_14118);
nand U14838 (N_14838,N_14434,N_14381);
xnor U14839 (N_14839,N_14134,N_14226);
nand U14840 (N_14840,N_14205,N_14021);
nand U14841 (N_14841,N_14342,N_14127);
and U14842 (N_14842,N_14471,N_14414);
xnor U14843 (N_14843,N_14114,N_14437);
nor U14844 (N_14844,N_14250,N_14217);
and U14845 (N_14845,N_14078,N_14126);
and U14846 (N_14846,N_14427,N_14466);
and U14847 (N_14847,N_14481,N_14116);
xor U14848 (N_14848,N_14228,N_14407);
nor U14849 (N_14849,N_14264,N_14406);
nor U14850 (N_14850,N_14391,N_14093);
nand U14851 (N_14851,N_14069,N_14202);
xor U14852 (N_14852,N_14314,N_14174);
nor U14853 (N_14853,N_14362,N_14277);
or U14854 (N_14854,N_14228,N_14196);
or U14855 (N_14855,N_14163,N_14417);
or U14856 (N_14856,N_14366,N_14177);
xor U14857 (N_14857,N_14025,N_14295);
nand U14858 (N_14858,N_14313,N_14205);
nand U14859 (N_14859,N_14265,N_14493);
nand U14860 (N_14860,N_14050,N_14142);
xnor U14861 (N_14861,N_14042,N_14190);
nor U14862 (N_14862,N_14172,N_14160);
nand U14863 (N_14863,N_14181,N_14114);
nor U14864 (N_14864,N_14291,N_14299);
nand U14865 (N_14865,N_14473,N_14370);
and U14866 (N_14866,N_14098,N_14110);
or U14867 (N_14867,N_14356,N_14483);
and U14868 (N_14868,N_14491,N_14462);
nor U14869 (N_14869,N_14489,N_14155);
nor U14870 (N_14870,N_14180,N_14287);
nand U14871 (N_14871,N_14017,N_14169);
or U14872 (N_14872,N_14051,N_14454);
nand U14873 (N_14873,N_14087,N_14399);
and U14874 (N_14874,N_14387,N_14484);
or U14875 (N_14875,N_14427,N_14382);
and U14876 (N_14876,N_14229,N_14380);
nor U14877 (N_14877,N_14391,N_14497);
xnor U14878 (N_14878,N_14417,N_14023);
and U14879 (N_14879,N_14490,N_14199);
and U14880 (N_14880,N_14128,N_14110);
nor U14881 (N_14881,N_14079,N_14461);
and U14882 (N_14882,N_14296,N_14287);
nor U14883 (N_14883,N_14331,N_14448);
nand U14884 (N_14884,N_14473,N_14222);
or U14885 (N_14885,N_14121,N_14182);
or U14886 (N_14886,N_14322,N_14135);
nor U14887 (N_14887,N_14275,N_14293);
and U14888 (N_14888,N_14232,N_14018);
and U14889 (N_14889,N_14369,N_14135);
nand U14890 (N_14890,N_14083,N_14181);
nand U14891 (N_14891,N_14215,N_14269);
xnor U14892 (N_14892,N_14087,N_14079);
xor U14893 (N_14893,N_14125,N_14274);
and U14894 (N_14894,N_14243,N_14077);
xor U14895 (N_14895,N_14179,N_14088);
xnor U14896 (N_14896,N_14214,N_14117);
nor U14897 (N_14897,N_14386,N_14001);
nand U14898 (N_14898,N_14405,N_14165);
or U14899 (N_14899,N_14044,N_14423);
nand U14900 (N_14900,N_14210,N_14163);
and U14901 (N_14901,N_14266,N_14040);
nand U14902 (N_14902,N_14479,N_14005);
and U14903 (N_14903,N_14221,N_14391);
and U14904 (N_14904,N_14104,N_14040);
nand U14905 (N_14905,N_14210,N_14027);
nor U14906 (N_14906,N_14176,N_14244);
or U14907 (N_14907,N_14468,N_14482);
xnor U14908 (N_14908,N_14165,N_14223);
xnor U14909 (N_14909,N_14352,N_14145);
nand U14910 (N_14910,N_14076,N_14234);
or U14911 (N_14911,N_14120,N_14063);
and U14912 (N_14912,N_14122,N_14325);
or U14913 (N_14913,N_14097,N_14067);
nand U14914 (N_14914,N_14329,N_14336);
nor U14915 (N_14915,N_14200,N_14312);
xor U14916 (N_14916,N_14413,N_14215);
nand U14917 (N_14917,N_14403,N_14409);
or U14918 (N_14918,N_14200,N_14007);
nor U14919 (N_14919,N_14183,N_14224);
and U14920 (N_14920,N_14490,N_14397);
nand U14921 (N_14921,N_14311,N_14036);
xor U14922 (N_14922,N_14335,N_14046);
nor U14923 (N_14923,N_14076,N_14401);
nand U14924 (N_14924,N_14205,N_14358);
nand U14925 (N_14925,N_14433,N_14252);
nor U14926 (N_14926,N_14139,N_14458);
nand U14927 (N_14927,N_14053,N_14311);
nor U14928 (N_14928,N_14193,N_14387);
and U14929 (N_14929,N_14014,N_14029);
nand U14930 (N_14930,N_14089,N_14061);
and U14931 (N_14931,N_14305,N_14238);
or U14932 (N_14932,N_14229,N_14177);
nor U14933 (N_14933,N_14018,N_14455);
nand U14934 (N_14934,N_14456,N_14307);
xnor U14935 (N_14935,N_14221,N_14057);
and U14936 (N_14936,N_14275,N_14322);
nand U14937 (N_14937,N_14397,N_14132);
and U14938 (N_14938,N_14226,N_14001);
nor U14939 (N_14939,N_14008,N_14113);
nor U14940 (N_14940,N_14239,N_14432);
nand U14941 (N_14941,N_14084,N_14124);
xor U14942 (N_14942,N_14482,N_14314);
and U14943 (N_14943,N_14279,N_14080);
xor U14944 (N_14944,N_14330,N_14151);
nor U14945 (N_14945,N_14208,N_14198);
nor U14946 (N_14946,N_14292,N_14486);
nand U14947 (N_14947,N_14358,N_14287);
or U14948 (N_14948,N_14068,N_14199);
nand U14949 (N_14949,N_14273,N_14261);
xnor U14950 (N_14950,N_14446,N_14138);
or U14951 (N_14951,N_14337,N_14291);
nand U14952 (N_14952,N_14060,N_14326);
nand U14953 (N_14953,N_14038,N_14195);
xnor U14954 (N_14954,N_14060,N_14164);
xnor U14955 (N_14955,N_14050,N_14481);
and U14956 (N_14956,N_14235,N_14345);
xnor U14957 (N_14957,N_14346,N_14228);
nor U14958 (N_14958,N_14158,N_14245);
nor U14959 (N_14959,N_14057,N_14214);
or U14960 (N_14960,N_14167,N_14103);
nor U14961 (N_14961,N_14377,N_14312);
and U14962 (N_14962,N_14305,N_14177);
and U14963 (N_14963,N_14196,N_14381);
nand U14964 (N_14964,N_14301,N_14206);
and U14965 (N_14965,N_14291,N_14287);
nor U14966 (N_14966,N_14156,N_14281);
nor U14967 (N_14967,N_14451,N_14082);
and U14968 (N_14968,N_14045,N_14176);
nor U14969 (N_14969,N_14297,N_14215);
nor U14970 (N_14970,N_14046,N_14303);
nor U14971 (N_14971,N_14401,N_14230);
or U14972 (N_14972,N_14452,N_14146);
and U14973 (N_14973,N_14296,N_14046);
nand U14974 (N_14974,N_14247,N_14413);
and U14975 (N_14975,N_14179,N_14284);
and U14976 (N_14976,N_14133,N_14311);
xnor U14977 (N_14977,N_14449,N_14297);
nor U14978 (N_14978,N_14267,N_14135);
nand U14979 (N_14979,N_14276,N_14028);
or U14980 (N_14980,N_14006,N_14450);
xor U14981 (N_14981,N_14327,N_14492);
nor U14982 (N_14982,N_14353,N_14008);
nor U14983 (N_14983,N_14301,N_14240);
nor U14984 (N_14984,N_14098,N_14428);
or U14985 (N_14985,N_14417,N_14175);
nand U14986 (N_14986,N_14394,N_14365);
and U14987 (N_14987,N_14366,N_14206);
xor U14988 (N_14988,N_14279,N_14490);
and U14989 (N_14989,N_14001,N_14133);
xnor U14990 (N_14990,N_14071,N_14397);
nand U14991 (N_14991,N_14186,N_14219);
nand U14992 (N_14992,N_14367,N_14269);
nand U14993 (N_14993,N_14479,N_14119);
nor U14994 (N_14994,N_14157,N_14137);
nor U14995 (N_14995,N_14380,N_14324);
and U14996 (N_14996,N_14428,N_14417);
and U14997 (N_14997,N_14172,N_14173);
xor U14998 (N_14998,N_14199,N_14211);
xnor U14999 (N_14999,N_14247,N_14240);
nor U15000 (N_15000,N_14586,N_14732);
nor U15001 (N_15001,N_14944,N_14703);
nor U15002 (N_15002,N_14733,N_14953);
nand U15003 (N_15003,N_14834,N_14699);
xnor U15004 (N_15004,N_14686,N_14937);
nor U15005 (N_15005,N_14745,N_14661);
nor U15006 (N_15006,N_14652,N_14663);
or U15007 (N_15007,N_14889,N_14649);
xor U15008 (N_15008,N_14566,N_14550);
xor U15009 (N_15009,N_14915,N_14867);
nand U15010 (N_15010,N_14601,N_14822);
and U15011 (N_15011,N_14805,N_14910);
nand U15012 (N_15012,N_14752,N_14987);
and U15013 (N_15013,N_14708,N_14885);
or U15014 (N_15014,N_14869,N_14832);
or U15015 (N_15015,N_14780,N_14627);
xnor U15016 (N_15016,N_14786,N_14858);
xnor U15017 (N_15017,N_14777,N_14809);
and U15018 (N_15018,N_14619,N_14818);
nand U15019 (N_15019,N_14782,N_14919);
xnor U15020 (N_15020,N_14602,N_14685);
and U15021 (N_15021,N_14897,N_14784);
or U15022 (N_15022,N_14743,N_14877);
and U15023 (N_15023,N_14861,N_14839);
nor U15024 (N_15024,N_14914,N_14746);
or U15025 (N_15025,N_14640,N_14545);
or U15026 (N_15026,N_14678,N_14501);
and U15027 (N_15027,N_14521,N_14552);
or U15028 (N_15028,N_14544,N_14905);
xnor U15029 (N_15029,N_14995,N_14612);
nand U15030 (N_15030,N_14626,N_14965);
and U15031 (N_15031,N_14622,N_14591);
nand U15032 (N_15032,N_14971,N_14862);
xnor U15033 (N_15033,N_14671,N_14928);
and U15034 (N_15034,N_14924,N_14992);
and U15035 (N_15035,N_14880,N_14578);
nand U15036 (N_15036,N_14581,N_14668);
or U15037 (N_15037,N_14679,N_14765);
nor U15038 (N_15038,N_14962,N_14842);
or U15039 (N_15039,N_14892,N_14674);
nand U15040 (N_15040,N_14943,N_14808);
nor U15041 (N_15041,N_14655,N_14998);
or U15042 (N_15042,N_14868,N_14823);
and U15043 (N_15043,N_14879,N_14875);
nand U15044 (N_15044,N_14583,N_14884);
or U15045 (N_15045,N_14543,N_14511);
xnor U15046 (N_15046,N_14744,N_14701);
nand U15047 (N_15047,N_14532,N_14888);
or U15048 (N_15048,N_14647,N_14956);
or U15049 (N_15049,N_14795,N_14692);
or U15050 (N_15050,N_14579,N_14909);
xor U15051 (N_15051,N_14577,N_14650);
nand U15052 (N_15052,N_14551,N_14694);
or U15053 (N_15053,N_14908,N_14528);
nand U15054 (N_15054,N_14828,N_14604);
and U15055 (N_15055,N_14819,N_14705);
xor U15056 (N_15056,N_14973,N_14712);
nand U15057 (N_15057,N_14955,N_14739);
nand U15058 (N_15058,N_14932,N_14999);
nand U15059 (N_15059,N_14589,N_14680);
and U15060 (N_15060,N_14593,N_14664);
xor U15061 (N_15061,N_14959,N_14632);
nand U15062 (N_15062,N_14850,N_14616);
nand U15063 (N_15063,N_14553,N_14574);
nor U15064 (N_15064,N_14636,N_14523);
xor U15065 (N_15065,N_14548,N_14810);
xor U15066 (N_15066,N_14527,N_14698);
and U15067 (N_15067,N_14524,N_14906);
and U15068 (N_15068,N_14855,N_14886);
and U15069 (N_15069,N_14653,N_14554);
nand U15070 (N_15070,N_14623,N_14558);
and U15071 (N_15071,N_14913,N_14618);
nand U15072 (N_15072,N_14935,N_14917);
xnor U15073 (N_15073,N_14696,N_14563);
or U15074 (N_15074,N_14595,N_14584);
and U15075 (N_15075,N_14568,N_14735);
or U15076 (N_15076,N_14588,N_14714);
nor U15077 (N_15077,N_14723,N_14961);
nand U15078 (N_15078,N_14970,N_14507);
nand U15079 (N_15079,N_14641,N_14547);
and U15080 (N_15080,N_14922,N_14831);
and U15081 (N_15081,N_14951,N_14756);
xor U15082 (N_15082,N_14903,N_14916);
nor U15083 (N_15083,N_14846,N_14534);
nor U15084 (N_15084,N_14871,N_14721);
nor U15085 (N_15085,N_14736,N_14575);
or U15086 (N_15086,N_14630,N_14994);
and U15087 (N_15087,N_14522,N_14603);
or U15088 (N_15088,N_14700,N_14681);
nand U15089 (N_15089,N_14878,N_14695);
nor U15090 (N_15090,N_14946,N_14853);
xnor U15091 (N_15091,N_14991,N_14576);
and U15092 (N_15092,N_14538,N_14654);
nand U15093 (N_15093,N_14900,N_14969);
nor U15094 (N_15094,N_14560,N_14729);
nor U15095 (N_15095,N_14976,N_14975);
or U15096 (N_15096,N_14719,N_14754);
and U15097 (N_15097,N_14631,N_14934);
and U15098 (N_15098,N_14510,N_14741);
and U15099 (N_15099,N_14774,N_14711);
nand U15100 (N_15100,N_14748,N_14557);
nor U15101 (N_15101,N_14675,N_14881);
nand U15102 (N_15102,N_14642,N_14972);
xnor U15103 (N_15103,N_14614,N_14860);
nor U15104 (N_15104,N_14502,N_14787);
and U15105 (N_15105,N_14982,N_14948);
and U15106 (N_15106,N_14830,N_14981);
nor U15107 (N_15107,N_14607,N_14931);
nand U15108 (N_15108,N_14779,N_14738);
or U15109 (N_15109,N_14598,N_14531);
nor U15110 (N_15110,N_14635,N_14911);
nor U15111 (N_15111,N_14565,N_14841);
xnor U15112 (N_15112,N_14725,N_14837);
or U15113 (N_15113,N_14519,N_14728);
xnor U15114 (N_15114,N_14835,N_14540);
and U15115 (N_15115,N_14838,N_14503);
nand U15116 (N_15116,N_14770,N_14791);
xor U15117 (N_15117,N_14793,N_14676);
xor U15118 (N_15118,N_14988,N_14669);
nor U15119 (N_15119,N_14580,N_14573);
or U15120 (N_15120,N_14849,N_14673);
and U15121 (N_15121,N_14517,N_14806);
and U15122 (N_15122,N_14516,N_14968);
or U15123 (N_15123,N_14803,N_14947);
nor U15124 (N_15124,N_14672,N_14542);
or U15125 (N_15125,N_14600,N_14755);
xor U15126 (N_15126,N_14514,N_14559);
and U15127 (N_15127,N_14926,N_14870);
and U15128 (N_15128,N_14824,N_14677);
xor U15129 (N_15129,N_14829,N_14597);
nand U15130 (N_15130,N_14984,N_14771);
nand U15131 (N_15131,N_14762,N_14585);
or U15132 (N_15132,N_14859,N_14785);
xor U15133 (N_15133,N_14772,N_14945);
xor U15134 (N_15134,N_14899,N_14977);
and U15135 (N_15135,N_14512,N_14620);
xnor U15136 (N_15136,N_14920,N_14963);
nor U15137 (N_15137,N_14727,N_14617);
and U15138 (N_15138,N_14891,N_14986);
nor U15139 (N_15139,N_14781,N_14820);
and U15140 (N_15140,N_14907,N_14866);
or U15141 (N_15141,N_14717,N_14561);
nor U15142 (N_15142,N_14940,N_14596);
or U15143 (N_15143,N_14960,N_14556);
and U15144 (N_15144,N_14515,N_14950);
or U15145 (N_15145,N_14776,N_14767);
and U15146 (N_15146,N_14798,N_14590);
or U15147 (N_15147,N_14833,N_14667);
or U15148 (N_15148,N_14904,N_14769);
nand U15149 (N_15149,N_14788,N_14709);
and U15150 (N_15150,N_14792,N_14646);
xor U15151 (N_15151,N_14827,N_14876);
and U15152 (N_15152,N_14742,N_14691);
or U15153 (N_15153,N_14980,N_14638);
and U15154 (N_15154,N_14933,N_14807);
or U15155 (N_15155,N_14857,N_14634);
and U15156 (N_15156,N_14656,N_14958);
nor U15157 (N_15157,N_14500,N_14724);
xor U15158 (N_15158,N_14844,N_14628);
nand U15159 (N_15159,N_14766,N_14582);
and U15160 (N_15160,N_14689,N_14670);
nand U15161 (N_15161,N_14804,N_14865);
and U15162 (N_15162,N_14687,N_14683);
nand U15163 (N_15163,N_14985,N_14525);
nor U15164 (N_15164,N_14845,N_14764);
and U15165 (N_15165,N_14644,N_14570);
or U15166 (N_15166,N_14979,N_14993);
nand U15167 (N_15167,N_14504,N_14821);
nor U15168 (N_15168,N_14882,N_14684);
nand U15169 (N_15169,N_14759,N_14930);
nor U15170 (N_15170,N_14535,N_14873);
nor U15171 (N_15171,N_14657,N_14811);
and U15172 (N_15172,N_14939,N_14802);
and U15173 (N_15173,N_14942,N_14726);
and U15174 (N_15174,N_14760,N_14541);
xnor U15175 (N_15175,N_14513,N_14665);
or U15176 (N_15176,N_14912,N_14624);
nand U15177 (N_15177,N_14957,N_14812);
nor U15178 (N_15178,N_14796,N_14569);
nor U15179 (N_15179,N_14936,N_14989);
xor U15180 (N_15180,N_14996,N_14658);
nor U15181 (N_15181,N_14789,N_14747);
or U15182 (N_15182,N_14800,N_14610);
nor U15183 (N_15183,N_14530,N_14660);
nand U15184 (N_15184,N_14520,N_14768);
or U15185 (N_15185,N_14927,N_14506);
xor U15186 (N_15186,N_14737,N_14509);
or U15187 (N_15187,N_14843,N_14592);
and U15188 (N_15188,N_14901,N_14666);
or U15189 (N_15189,N_14713,N_14949);
xor U15190 (N_15190,N_14826,N_14533);
or U15191 (N_15191,N_14615,N_14983);
nand U15192 (N_15192,N_14763,N_14710);
nand U15193 (N_15193,N_14505,N_14609);
or U15194 (N_15194,N_14757,N_14918);
or U15195 (N_15195,N_14740,N_14790);
nor U15196 (N_15196,N_14990,N_14722);
nor U15197 (N_15197,N_14887,N_14864);
nor U15198 (N_15198,N_14555,N_14606);
nor U15199 (N_15199,N_14707,N_14817);
xnor U15200 (N_15200,N_14613,N_14974);
or U15201 (N_15201,N_14799,N_14704);
or U15202 (N_15202,N_14587,N_14890);
and U15203 (N_15203,N_14536,N_14758);
and U15204 (N_15204,N_14702,N_14750);
or U15205 (N_15205,N_14706,N_14967);
nor U15206 (N_15206,N_14539,N_14651);
nor U15207 (N_15207,N_14761,N_14954);
and U15208 (N_15208,N_14572,N_14852);
nand U15209 (N_15209,N_14693,N_14952);
and U15210 (N_15210,N_14836,N_14938);
nand U15211 (N_15211,N_14716,N_14643);
nand U15212 (N_15212,N_14978,N_14895);
xnor U15213 (N_15213,N_14734,N_14718);
and U15214 (N_15214,N_14863,N_14773);
xor U15215 (N_15215,N_14921,N_14648);
nor U15216 (N_15216,N_14923,N_14848);
xnor U15217 (N_15217,N_14847,N_14872);
nand U15218 (N_15218,N_14751,N_14783);
xor U15219 (N_15219,N_14801,N_14690);
or U15220 (N_15220,N_14625,N_14893);
and U15221 (N_15221,N_14608,N_14688);
or U15222 (N_15222,N_14599,N_14964);
or U15223 (N_15223,N_14546,N_14854);
or U15224 (N_15224,N_14775,N_14797);
or U15225 (N_15225,N_14682,N_14749);
nand U15226 (N_15226,N_14715,N_14902);
and U15227 (N_15227,N_14814,N_14778);
or U15228 (N_15228,N_14605,N_14929);
nor U15229 (N_15229,N_14518,N_14537);
xnor U15230 (N_15230,N_14571,N_14856);
nor U15231 (N_15231,N_14567,N_14549);
or U15232 (N_15232,N_14662,N_14731);
nor U15233 (N_15233,N_14621,N_14697);
nor U15234 (N_15234,N_14894,N_14813);
nor U15235 (N_15235,N_14874,N_14659);
or U15236 (N_15236,N_14896,N_14645);
or U15237 (N_15237,N_14840,N_14629);
nor U15238 (N_15238,N_14637,N_14825);
nand U15239 (N_15239,N_14997,N_14815);
xor U15240 (N_15240,N_14611,N_14529);
and U15241 (N_15241,N_14730,N_14720);
or U15242 (N_15242,N_14633,N_14562);
or U15243 (N_15243,N_14564,N_14883);
xor U15244 (N_15244,N_14753,N_14966);
and U15245 (N_15245,N_14639,N_14851);
or U15246 (N_15246,N_14526,N_14816);
and U15247 (N_15247,N_14594,N_14925);
or U15248 (N_15248,N_14941,N_14794);
nand U15249 (N_15249,N_14898,N_14508);
nand U15250 (N_15250,N_14853,N_14888);
and U15251 (N_15251,N_14730,N_14709);
nand U15252 (N_15252,N_14691,N_14650);
nand U15253 (N_15253,N_14510,N_14700);
xnor U15254 (N_15254,N_14664,N_14564);
and U15255 (N_15255,N_14823,N_14502);
nand U15256 (N_15256,N_14606,N_14638);
or U15257 (N_15257,N_14630,N_14869);
xnor U15258 (N_15258,N_14547,N_14546);
and U15259 (N_15259,N_14812,N_14748);
nor U15260 (N_15260,N_14632,N_14805);
nand U15261 (N_15261,N_14751,N_14800);
nand U15262 (N_15262,N_14709,N_14916);
or U15263 (N_15263,N_14923,N_14595);
nand U15264 (N_15264,N_14785,N_14934);
and U15265 (N_15265,N_14871,N_14958);
xor U15266 (N_15266,N_14704,N_14749);
xor U15267 (N_15267,N_14514,N_14668);
nor U15268 (N_15268,N_14693,N_14502);
and U15269 (N_15269,N_14801,N_14960);
nor U15270 (N_15270,N_14760,N_14622);
nor U15271 (N_15271,N_14914,N_14715);
nor U15272 (N_15272,N_14536,N_14861);
nor U15273 (N_15273,N_14946,N_14769);
xor U15274 (N_15274,N_14725,N_14982);
xor U15275 (N_15275,N_14651,N_14889);
xor U15276 (N_15276,N_14922,N_14849);
nor U15277 (N_15277,N_14701,N_14750);
nand U15278 (N_15278,N_14970,N_14681);
nor U15279 (N_15279,N_14541,N_14780);
nand U15280 (N_15280,N_14617,N_14725);
nand U15281 (N_15281,N_14948,N_14716);
nor U15282 (N_15282,N_14922,N_14997);
nor U15283 (N_15283,N_14954,N_14806);
nand U15284 (N_15284,N_14667,N_14778);
nor U15285 (N_15285,N_14770,N_14853);
nor U15286 (N_15286,N_14536,N_14694);
xnor U15287 (N_15287,N_14615,N_14678);
and U15288 (N_15288,N_14692,N_14662);
nand U15289 (N_15289,N_14931,N_14835);
and U15290 (N_15290,N_14854,N_14931);
nor U15291 (N_15291,N_14625,N_14783);
nor U15292 (N_15292,N_14738,N_14789);
xor U15293 (N_15293,N_14757,N_14954);
nor U15294 (N_15294,N_14819,N_14512);
and U15295 (N_15295,N_14810,N_14611);
or U15296 (N_15296,N_14695,N_14713);
or U15297 (N_15297,N_14620,N_14864);
nand U15298 (N_15298,N_14918,N_14580);
nor U15299 (N_15299,N_14994,N_14520);
or U15300 (N_15300,N_14779,N_14868);
nor U15301 (N_15301,N_14942,N_14888);
and U15302 (N_15302,N_14993,N_14581);
and U15303 (N_15303,N_14908,N_14939);
and U15304 (N_15304,N_14767,N_14861);
and U15305 (N_15305,N_14873,N_14679);
nor U15306 (N_15306,N_14787,N_14757);
nor U15307 (N_15307,N_14861,N_14965);
xor U15308 (N_15308,N_14956,N_14973);
xnor U15309 (N_15309,N_14745,N_14849);
nor U15310 (N_15310,N_14769,N_14948);
nand U15311 (N_15311,N_14695,N_14959);
nor U15312 (N_15312,N_14587,N_14952);
nor U15313 (N_15313,N_14552,N_14528);
nand U15314 (N_15314,N_14921,N_14644);
xnor U15315 (N_15315,N_14823,N_14842);
nand U15316 (N_15316,N_14754,N_14656);
or U15317 (N_15317,N_14853,N_14506);
nand U15318 (N_15318,N_14558,N_14903);
nor U15319 (N_15319,N_14695,N_14810);
nand U15320 (N_15320,N_14765,N_14520);
or U15321 (N_15321,N_14577,N_14977);
or U15322 (N_15322,N_14703,N_14826);
or U15323 (N_15323,N_14960,N_14651);
nor U15324 (N_15324,N_14581,N_14671);
and U15325 (N_15325,N_14553,N_14749);
nor U15326 (N_15326,N_14586,N_14719);
nor U15327 (N_15327,N_14859,N_14753);
nand U15328 (N_15328,N_14522,N_14952);
or U15329 (N_15329,N_14783,N_14609);
nand U15330 (N_15330,N_14881,N_14533);
or U15331 (N_15331,N_14874,N_14644);
or U15332 (N_15332,N_14962,N_14967);
nand U15333 (N_15333,N_14894,N_14769);
nor U15334 (N_15334,N_14505,N_14564);
nand U15335 (N_15335,N_14923,N_14845);
or U15336 (N_15336,N_14668,N_14643);
xnor U15337 (N_15337,N_14582,N_14773);
or U15338 (N_15338,N_14754,N_14652);
or U15339 (N_15339,N_14585,N_14807);
or U15340 (N_15340,N_14662,N_14699);
or U15341 (N_15341,N_14949,N_14842);
xor U15342 (N_15342,N_14768,N_14540);
nor U15343 (N_15343,N_14892,N_14779);
nor U15344 (N_15344,N_14750,N_14544);
nand U15345 (N_15345,N_14812,N_14677);
nand U15346 (N_15346,N_14933,N_14814);
or U15347 (N_15347,N_14528,N_14941);
nor U15348 (N_15348,N_14547,N_14626);
nand U15349 (N_15349,N_14561,N_14563);
nor U15350 (N_15350,N_14902,N_14805);
xnor U15351 (N_15351,N_14983,N_14624);
nor U15352 (N_15352,N_14503,N_14582);
and U15353 (N_15353,N_14936,N_14910);
nand U15354 (N_15354,N_14593,N_14712);
xnor U15355 (N_15355,N_14908,N_14785);
and U15356 (N_15356,N_14765,N_14633);
xor U15357 (N_15357,N_14595,N_14614);
nor U15358 (N_15358,N_14894,N_14953);
or U15359 (N_15359,N_14655,N_14930);
nor U15360 (N_15360,N_14677,N_14776);
nand U15361 (N_15361,N_14755,N_14968);
and U15362 (N_15362,N_14766,N_14847);
or U15363 (N_15363,N_14932,N_14620);
or U15364 (N_15364,N_14954,N_14595);
and U15365 (N_15365,N_14918,N_14592);
nand U15366 (N_15366,N_14611,N_14767);
nand U15367 (N_15367,N_14543,N_14637);
nor U15368 (N_15368,N_14814,N_14929);
and U15369 (N_15369,N_14560,N_14515);
and U15370 (N_15370,N_14959,N_14662);
and U15371 (N_15371,N_14727,N_14845);
or U15372 (N_15372,N_14769,N_14777);
nor U15373 (N_15373,N_14735,N_14565);
and U15374 (N_15374,N_14572,N_14585);
xnor U15375 (N_15375,N_14561,N_14739);
nand U15376 (N_15376,N_14557,N_14869);
nor U15377 (N_15377,N_14987,N_14876);
nand U15378 (N_15378,N_14500,N_14998);
or U15379 (N_15379,N_14831,N_14844);
nor U15380 (N_15380,N_14872,N_14790);
xnor U15381 (N_15381,N_14645,N_14793);
and U15382 (N_15382,N_14921,N_14911);
and U15383 (N_15383,N_14696,N_14747);
or U15384 (N_15384,N_14840,N_14975);
nand U15385 (N_15385,N_14832,N_14909);
nand U15386 (N_15386,N_14667,N_14738);
or U15387 (N_15387,N_14523,N_14640);
nor U15388 (N_15388,N_14662,N_14735);
or U15389 (N_15389,N_14956,N_14951);
nor U15390 (N_15390,N_14977,N_14518);
and U15391 (N_15391,N_14682,N_14872);
xor U15392 (N_15392,N_14994,N_14918);
or U15393 (N_15393,N_14594,N_14908);
nor U15394 (N_15394,N_14827,N_14982);
xor U15395 (N_15395,N_14882,N_14609);
or U15396 (N_15396,N_14934,N_14796);
xnor U15397 (N_15397,N_14661,N_14814);
nand U15398 (N_15398,N_14701,N_14629);
nand U15399 (N_15399,N_14843,N_14503);
nand U15400 (N_15400,N_14823,N_14815);
and U15401 (N_15401,N_14859,N_14628);
and U15402 (N_15402,N_14997,N_14629);
nor U15403 (N_15403,N_14938,N_14614);
xnor U15404 (N_15404,N_14552,N_14631);
and U15405 (N_15405,N_14578,N_14720);
nor U15406 (N_15406,N_14676,N_14625);
nand U15407 (N_15407,N_14609,N_14518);
or U15408 (N_15408,N_14563,N_14886);
and U15409 (N_15409,N_14875,N_14519);
xnor U15410 (N_15410,N_14647,N_14616);
nor U15411 (N_15411,N_14972,N_14760);
xor U15412 (N_15412,N_14538,N_14707);
and U15413 (N_15413,N_14694,N_14581);
or U15414 (N_15414,N_14516,N_14952);
and U15415 (N_15415,N_14594,N_14910);
and U15416 (N_15416,N_14847,N_14868);
xor U15417 (N_15417,N_14553,N_14593);
nand U15418 (N_15418,N_14640,N_14712);
nand U15419 (N_15419,N_14931,N_14605);
nor U15420 (N_15420,N_14965,N_14745);
and U15421 (N_15421,N_14939,N_14747);
xor U15422 (N_15422,N_14559,N_14861);
and U15423 (N_15423,N_14575,N_14612);
nand U15424 (N_15424,N_14950,N_14629);
nand U15425 (N_15425,N_14895,N_14582);
and U15426 (N_15426,N_14741,N_14919);
nor U15427 (N_15427,N_14611,N_14860);
nor U15428 (N_15428,N_14782,N_14836);
nor U15429 (N_15429,N_14959,N_14779);
nand U15430 (N_15430,N_14843,N_14566);
nor U15431 (N_15431,N_14726,N_14869);
nor U15432 (N_15432,N_14865,N_14874);
nor U15433 (N_15433,N_14744,N_14614);
or U15434 (N_15434,N_14869,N_14540);
and U15435 (N_15435,N_14819,N_14661);
or U15436 (N_15436,N_14708,N_14831);
xnor U15437 (N_15437,N_14565,N_14547);
nand U15438 (N_15438,N_14609,N_14747);
and U15439 (N_15439,N_14923,N_14655);
xnor U15440 (N_15440,N_14984,N_14906);
and U15441 (N_15441,N_14550,N_14764);
or U15442 (N_15442,N_14853,N_14769);
or U15443 (N_15443,N_14624,N_14645);
or U15444 (N_15444,N_14959,N_14820);
and U15445 (N_15445,N_14875,N_14666);
or U15446 (N_15446,N_14914,N_14636);
and U15447 (N_15447,N_14594,N_14553);
nor U15448 (N_15448,N_14651,N_14712);
xnor U15449 (N_15449,N_14676,N_14707);
nand U15450 (N_15450,N_14505,N_14567);
and U15451 (N_15451,N_14543,N_14616);
xnor U15452 (N_15452,N_14606,N_14835);
or U15453 (N_15453,N_14592,N_14851);
nor U15454 (N_15454,N_14829,N_14935);
xnor U15455 (N_15455,N_14990,N_14588);
nand U15456 (N_15456,N_14535,N_14588);
nand U15457 (N_15457,N_14935,N_14965);
nand U15458 (N_15458,N_14736,N_14581);
nor U15459 (N_15459,N_14540,N_14973);
nand U15460 (N_15460,N_14997,N_14548);
or U15461 (N_15461,N_14560,N_14979);
nand U15462 (N_15462,N_14819,N_14750);
and U15463 (N_15463,N_14884,N_14922);
nand U15464 (N_15464,N_14570,N_14916);
and U15465 (N_15465,N_14934,N_14640);
or U15466 (N_15466,N_14706,N_14970);
nor U15467 (N_15467,N_14724,N_14692);
nand U15468 (N_15468,N_14775,N_14525);
or U15469 (N_15469,N_14685,N_14507);
or U15470 (N_15470,N_14902,N_14631);
nand U15471 (N_15471,N_14862,N_14776);
nor U15472 (N_15472,N_14833,N_14605);
or U15473 (N_15473,N_14702,N_14891);
or U15474 (N_15474,N_14572,N_14932);
nor U15475 (N_15475,N_14855,N_14576);
and U15476 (N_15476,N_14831,N_14635);
nor U15477 (N_15477,N_14531,N_14920);
and U15478 (N_15478,N_14894,N_14593);
and U15479 (N_15479,N_14711,N_14681);
nor U15480 (N_15480,N_14801,N_14681);
or U15481 (N_15481,N_14591,N_14627);
nor U15482 (N_15482,N_14798,N_14704);
xor U15483 (N_15483,N_14777,N_14890);
or U15484 (N_15484,N_14986,N_14944);
xnor U15485 (N_15485,N_14558,N_14526);
nand U15486 (N_15486,N_14757,N_14721);
nand U15487 (N_15487,N_14777,N_14636);
and U15488 (N_15488,N_14540,N_14790);
or U15489 (N_15489,N_14697,N_14525);
xor U15490 (N_15490,N_14589,N_14778);
and U15491 (N_15491,N_14868,N_14603);
nor U15492 (N_15492,N_14600,N_14724);
or U15493 (N_15493,N_14876,N_14520);
nand U15494 (N_15494,N_14532,N_14868);
xor U15495 (N_15495,N_14881,N_14859);
xnor U15496 (N_15496,N_14853,N_14568);
nand U15497 (N_15497,N_14762,N_14792);
xor U15498 (N_15498,N_14926,N_14950);
and U15499 (N_15499,N_14682,N_14730);
nand U15500 (N_15500,N_15000,N_15333);
nor U15501 (N_15501,N_15475,N_15104);
or U15502 (N_15502,N_15001,N_15062);
nor U15503 (N_15503,N_15384,N_15040);
nor U15504 (N_15504,N_15464,N_15186);
nand U15505 (N_15505,N_15364,N_15382);
or U15506 (N_15506,N_15169,N_15353);
nand U15507 (N_15507,N_15217,N_15248);
nand U15508 (N_15508,N_15401,N_15376);
nor U15509 (N_15509,N_15130,N_15184);
nand U15510 (N_15510,N_15383,N_15146);
or U15511 (N_15511,N_15142,N_15010);
nand U15512 (N_15512,N_15348,N_15386);
or U15513 (N_15513,N_15168,N_15227);
xor U15514 (N_15514,N_15314,N_15312);
nand U15515 (N_15515,N_15499,N_15443);
nand U15516 (N_15516,N_15242,N_15439);
or U15517 (N_15517,N_15153,N_15393);
nor U15518 (N_15518,N_15291,N_15124);
and U15519 (N_15519,N_15273,N_15437);
or U15520 (N_15520,N_15224,N_15021);
nor U15521 (N_15521,N_15230,N_15418);
nand U15522 (N_15522,N_15349,N_15320);
nor U15523 (N_15523,N_15359,N_15252);
or U15524 (N_15524,N_15121,N_15152);
nor U15525 (N_15525,N_15059,N_15448);
or U15526 (N_15526,N_15057,N_15166);
xor U15527 (N_15527,N_15063,N_15022);
nand U15528 (N_15528,N_15163,N_15433);
nand U15529 (N_15529,N_15108,N_15025);
xor U15530 (N_15530,N_15192,N_15127);
nor U15531 (N_15531,N_15061,N_15329);
and U15532 (N_15532,N_15235,N_15373);
and U15533 (N_15533,N_15442,N_15473);
xnor U15534 (N_15534,N_15251,N_15212);
and U15535 (N_15535,N_15189,N_15005);
xnor U15536 (N_15536,N_15197,N_15322);
nand U15537 (N_15537,N_15238,N_15292);
nor U15538 (N_15538,N_15387,N_15255);
nor U15539 (N_15539,N_15222,N_15176);
nor U15540 (N_15540,N_15058,N_15159);
xor U15541 (N_15541,N_15150,N_15385);
nor U15542 (N_15542,N_15027,N_15103);
and U15543 (N_15543,N_15466,N_15096);
or U15544 (N_15544,N_15139,N_15013);
or U15545 (N_15545,N_15321,N_15404);
nor U15546 (N_15546,N_15099,N_15201);
nand U15547 (N_15547,N_15381,N_15380);
xnor U15548 (N_15548,N_15249,N_15165);
and U15549 (N_15549,N_15028,N_15094);
nor U15550 (N_15550,N_15115,N_15421);
nand U15551 (N_15551,N_15431,N_15125);
nor U15552 (N_15552,N_15215,N_15110);
or U15553 (N_15553,N_15424,N_15079);
nor U15554 (N_15554,N_15067,N_15299);
xnor U15555 (N_15555,N_15128,N_15081);
nor U15556 (N_15556,N_15016,N_15438);
nor U15557 (N_15557,N_15225,N_15363);
and U15558 (N_15558,N_15402,N_15428);
xor U15559 (N_15559,N_15318,N_15034);
or U15560 (N_15560,N_15074,N_15145);
and U15561 (N_15561,N_15469,N_15038);
nor U15562 (N_15562,N_15247,N_15253);
nor U15563 (N_15563,N_15307,N_15120);
nand U15564 (N_15564,N_15009,N_15478);
nand U15565 (N_15565,N_15471,N_15472);
nor U15566 (N_15566,N_15164,N_15347);
nand U15567 (N_15567,N_15037,N_15483);
nand U15568 (N_15568,N_15211,N_15411);
nor U15569 (N_15569,N_15129,N_15276);
nor U15570 (N_15570,N_15091,N_15268);
xor U15571 (N_15571,N_15491,N_15123);
nand U15572 (N_15572,N_15277,N_15371);
or U15573 (N_15573,N_15398,N_15098);
or U15574 (N_15574,N_15026,N_15459);
nand U15575 (N_15575,N_15293,N_15427);
nor U15576 (N_15576,N_15178,N_15205);
or U15577 (N_15577,N_15015,N_15107);
nand U15578 (N_15578,N_15114,N_15445);
or U15579 (N_15579,N_15301,N_15374);
or U15580 (N_15580,N_15002,N_15319);
nor U15581 (N_15581,N_15135,N_15368);
or U15582 (N_15582,N_15106,N_15048);
or U15583 (N_15583,N_15213,N_15199);
nand U15584 (N_15584,N_15282,N_15029);
nand U15585 (N_15585,N_15358,N_15423);
xor U15586 (N_15586,N_15350,N_15237);
and U15587 (N_15587,N_15018,N_15298);
or U15588 (N_15588,N_15147,N_15287);
nor U15589 (N_15589,N_15172,N_15181);
or U15590 (N_15590,N_15209,N_15187);
or U15591 (N_15591,N_15461,N_15486);
and U15592 (N_15592,N_15389,N_15269);
or U15593 (N_15593,N_15198,N_15069);
nand U15594 (N_15594,N_15195,N_15066);
nand U15595 (N_15595,N_15162,N_15075);
xor U15596 (N_15596,N_15035,N_15136);
and U15597 (N_15597,N_15304,N_15246);
xor U15598 (N_15598,N_15051,N_15143);
xor U15599 (N_15599,N_15467,N_15148);
xor U15600 (N_15600,N_15258,N_15392);
and U15601 (N_15601,N_15053,N_15216);
xnor U15602 (N_15602,N_15447,N_15378);
nand U15603 (N_15603,N_15126,N_15434);
xnor U15604 (N_15604,N_15167,N_15065);
and U15605 (N_15605,N_15100,N_15315);
xnor U15606 (N_15606,N_15033,N_15432);
xor U15607 (N_15607,N_15451,N_15405);
or U15608 (N_15608,N_15011,N_15444);
and U15609 (N_15609,N_15036,N_15207);
nand U15610 (N_15610,N_15400,N_15295);
or U15611 (N_15611,N_15117,N_15309);
or U15612 (N_15612,N_15245,N_15134);
xnor U15613 (N_15613,N_15446,N_15077);
xnor U15614 (N_15614,N_15236,N_15072);
nand U15615 (N_15615,N_15454,N_15485);
and U15616 (N_15616,N_15297,N_15453);
or U15617 (N_15617,N_15414,N_15468);
xnor U15618 (N_15618,N_15047,N_15019);
or U15619 (N_15619,N_15244,N_15351);
and U15620 (N_15620,N_15416,N_15041);
and U15621 (N_15621,N_15179,N_15030);
and U15622 (N_15622,N_15182,N_15259);
or U15623 (N_15623,N_15306,N_15090);
and U15624 (N_15624,N_15093,N_15221);
or U15625 (N_15625,N_15300,N_15204);
or U15626 (N_15626,N_15313,N_15489);
and U15627 (N_15627,N_15279,N_15233);
nand U15628 (N_15628,N_15390,N_15284);
or U15629 (N_15629,N_15285,N_15281);
xnor U15630 (N_15630,N_15337,N_15458);
xor U15631 (N_15631,N_15003,N_15457);
and U15632 (N_15632,N_15327,N_15267);
nor U15633 (N_15633,N_15484,N_15296);
or U15634 (N_15634,N_15177,N_15497);
nand U15635 (N_15635,N_15156,N_15155);
or U15636 (N_15636,N_15151,N_15495);
nand U15637 (N_15637,N_15365,N_15425);
xor U15638 (N_15638,N_15422,N_15007);
xor U15639 (N_15639,N_15109,N_15006);
or U15640 (N_15640,N_15008,N_15046);
and U15641 (N_15641,N_15289,N_15456);
xor U15642 (N_15642,N_15340,N_15388);
or U15643 (N_15643,N_15157,N_15487);
nor U15644 (N_15644,N_15430,N_15170);
and U15645 (N_15645,N_15426,N_15339);
nand U15646 (N_15646,N_15024,N_15449);
and U15647 (N_15647,N_15052,N_15399);
and U15648 (N_15648,N_15369,N_15362);
nand U15649 (N_15649,N_15133,N_15419);
and U15650 (N_15650,N_15477,N_15316);
or U15651 (N_15651,N_15070,N_15206);
nand U15652 (N_15652,N_15396,N_15455);
nand U15653 (N_15653,N_15012,N_15346);
or U15654 (N_15654,N_15078,N_15326);
xor U15655 (N_15655,N_15218,N_15345);
xnor U15656 (N_15656,N_15479,N_15440);
nand U15657 (N_15657,N_15308,N_15188);
xor U15658 (N_15658,N_15088,N_15290);
and U15659 (N_15659,N_15042,N_15305);
or U15660 (N_15660,N_15240,N_15420);
nor U15661 (N_15661,N_15262,N_15144);
or U15662 (N_15662,N_15004,N_15480);
xnor U15663 (N_15663,N_15089,N_15264);
and U15664 (N_15664,N_15055,N_15482);
or U15665 (N_15665,N_15375,N_15185);
nand U15666 (N_15666,N_15101,N_15085);
or U15667 (N_15667,N_15087,N_15355);
xor U15668 (N_15668,N_15226,N_15325);
nand U15669 (N_15669,N_15095,N_15415);
xnor U15670 (N_15670,N_15496,N_15196);
xnor U15671 (N_15671,N_15223,N_15200);
xnor U15672 (N_15672,N_15372,N_15360);
nor U15673 (N_15673,N_15234,N_15239);
or U15674 (N_15674,N_15083,N_15356);
xnor U15675 (N_15675,N_15272,N_15202);
xor U15676 (N_15676,N_15060,N_15336);
nor U15677 (N_15677,N_15498,N_15241);
and U15678 (N_15678,N_15203,N_15271);
and U15679 (N_15679,N_15450,N_15317);
xnor U15680 (N_15680,N_15334,N_15361);
nor U15681 (N_15681,N_15076,N_15288);
or U15682 (N_15682,N_15250,N_15113);
xnor U15683 (N_15683,N_15014,N_15017);
nand U15684 (N_15684,N_15413,N_15118);
nor U15685 (N_15685,N_15132,N_15131);
and U15686 (N_15686,N_15488,N_15462);
nand U15687 (N_15687,N_15435,N_15045);
and U15688 (N_15688,N_15476,N_15138);
nor U15689 (N_15689,N_15210,N_15180);
nand U15690 (N_15690,N_15474,N_15122);
nor U15691 (N_15691,N_15080,N_15191);
and U15692 (N_15692,N_15441,N_15231);
xnor U15693 (N_15693,N_15119,N_15054);
nand U15694 (N_15694,N_15032,N_15302);
and U15695 (N_15695,N_15116,N_15257);
or U15696 (N_15696,N_15278,N_15232);
and U15697 (N_15697,N_15274,N_15092);
or U15698 (N_15698,N_15228,N_15286);
xnor U15699 (N_15699,N_15260,N_15229);
nor U15700 (N_15700,N_15183,N_15254);
xnor U15701 (N_15701,N_15397,N_15082);
and U15702 (N_15702,N_15370,N_15141);
nor U15703 (N_15703,N_15270,N_15417);
nand U15704 (N_15704,N_15367,N_15214);
and U15705 (N_15705,N_15073,N_15490);
nor U15706 (N_15706,N_15068,N_15294);
nor U15707 (N_15707,N_15311,N_15194);
xor U15708 (N_15708,N_15310,N_15465);
xor U15709 (N_15709,N_15243,N_15330);
and U15710 (N_15710,N_15412,N_15086);
nand U15711 (N_15711,N_15023,N_15190);
nor U15712 (N_15712,N_15429,N_15111);
nand U15713 (N_15713,N_15391,N_15208);
nand U15714 (N_15714,N_15261,N_15344);
nand U15715 (N_15715,N_15377,N_15193);
or U15716 (N_15716,N_15357,N_15071);
nor U15717 (N_15717,N_15050,N_15492);
and U15718 (N_15718,N_15112,N_15043);
nor U15719 (N_15719,N_15049,N_15323);
nor U15720 (N_15720,N_15171,N_15280);
or U15721 (N_15721,N_15064,N_15265);
nand U15722 (N_15722,N_15366,N_15332);
nor U15723 (N_15723,N_15303,N_15493);
and U15724 (N_15724,N_15256,N_15039);
or U15725 (N_15725,N_15328,N_15097);
nand U15726 (N_15726,N_15266,N_15175);
xnor U15727 (N_15727,N_15341,N_15463);
xor U15728 (N_15728,N_15343,N_15470);
nand U15729 (N_15729,N_15452,N_15408);
or U15730 (N_15730,N_15406,N_15494);
or U15731 (N_15731,N_15056,N_15379);
xor U15732 (N_15732,N_15154,N_15084);
or U15733 (N_15733,N_15263,N_15324);
or U15734 (N_15734,N_15220,N_15410);
or U15735 (N_15735,N_15342,N_15044);
or U15736 (N_15736,N_15283,N_15031);
xor U15737 (N_15737,N_15409,N_15219);
nor U15738 (N_15738,N_15102,N_15140);
nand U15739 (N_15739,N_15174,N_15275);
and U15740 (N_15740,N_15158,N_15160);
xnor U15741 (N_15741,N_15394,N_15137);
xor U15742 (N_15742,N_15161,N_15407);
nand U15743 (N_15743,N_15173,N_15395);
nand U15744 (N_15744,N_15149,N_15335);
or U15745 (N_15745,N_15460,N_15403);
xnor U15746 (N_15746,N_15020,N_15354);
or U15747 (N_15747,N_15436,N_15338);
nand U15748 (N_15748,N_15331,N_15352);
xnor U15749 (N_15749,N_15105,N_15481);
nand U15750 (N_15750,N_15187,N_15088);
xnor U15751 (N_15751,N_15026,N_15275);
nor U15752 (N_15752,N_15468,N_15151);
xor U15753 (N_15753,N_15093,N_15496);
or U15754 (N_15754,N_15342,N_15011);
nand U15755 (N_15755,N_15487,N_15313);
and U15756 (N_15756,N_15156,N_15237);
xor U15757 (N_15757,N_15368,N_15484);
and U15758 (N_15758,N_15186,N_15080);
xnor U15759 (N_15759,N_15346,N_15407);
and U15760 (N_15760,N_15454,N_15284);
or U15761 (N_15761,N_15166,N_15294);
and U15762 (N_15762,N_15207,N_15490);
and U15763 (N_15763,N_15379,N_15180);
nand U15764 (N_15764,N_15067,N_15166);
or U15765 (N_15765,N_15117,N_15300);
and U15766 (N_15766,N_15479,N_15238);
or U15767 (N_15767,N_15122,N_15230);
and U15768 (N_15768,N_15430,N_15367);
xor U15769 (N_15769,N_15164,N_15324);
nand U15770 (N_15770,N_15296,N_15440);
nand U15771 (N_15771,N_15174,N_15198);
or U15772 (N_15772,N_15210,N_15438);
and U15773 (N_15773,N_15247,N_15080);
xor U15774 (N_15774,N_15428,N_15383);
nor U15775 (N_15775,N_15018,N_15246);
xor U15776 (N_15776,N_15460,N_15159);
and U15777 (N_15777,N_15434,N_15273);
nand U15778 (N_15778,N_15333,N_15255);
nand U15779 (N_15779,N_15432,N_15467);
nand U15780 (N_15780,N_15249,N_15151);
and U15781 (N_15781,N_15419,N_15458);
nor U15782 (N_15782,N_15021,N_15094);
xor U15783 (N_15783,N_15167,N_15127);
nand U15784 (N_15784,N_15413,N_15262);
or U15785 (N_15785,N_15228,N_15076);
nand U15786 (N_15786,N_15347,N_15334);
and U15787 (N_15787,N_15107,N_15048);
nand U15788 (N_15788,N_15312,N_15018);
xor U15789 (N_15789,N_15067,N_15223);
or U15790 (N_15790,N_15141,N_15225);
xor U15791 (N_15791,N_15316,N_15008);
xor U15792 (N_15792,N_15222,N_15419);
xnor U15793 (N_15793,N_15431,N_15346);
xnor U15794 (N_15794,N_15413,N_15043);
nand U15795 (N_15795,N_15200,N_15127);
xor U15796 (N_15796,N_15389,N_15174);
nor U15797 (N_15797,N_15128,N_15395);
nand U15798 (N_15798,N_15229,N_15021);
nand U15799 (N_15799,N_15059,N_15030);
nor U15800 (N_15800,N_15148,N_15017);
xor U15801 (N_15801,N_15467,N_15227);
or U15802 (N_15802,N_15335,N_15166);
nand U15803 (N_15803,N_15015,N_15121);
nand U15804 (N_15804,N_15171,N_15107);
nand U15805 (N_15805,N_15036,N_15443);
or U15806 (N_15806,N_15342,N_15410);
xor U15807 (N_15807,N_15398,N_15125);
and U15808 (N_15808,N_15308,N_15374);
or U15809 (N_15809,N_15325,N_15034);
and U15810 (N_15810,N_15132,N_15486);
and U15811 (N_15811,N_15481,N_15461);
nand U15812 (N_15812,N_15031,N_15324);
xor U15813 (N_15813,N_15265,N_15462);
nand U15814 (N_15814,N_15290,N_15316);
nor U15815 (N_15815,N_15481,N_15183);
or U15816 (N_15816,N_15036,N_15366);
nand U15817 (N_15817,N_15163,N_15224);
nor U15818 (N_15818,N_15365,N_15287);
nand U15819 (N_15819,N_15360,N_15245);
nor U15820 (N_15820,N_15080,N_15051);
xnor U15821 (N_15821,N_15025,N_15322);
xor U15822 (N_15822,N_15277,N_15259);
and U15823 (N_15823,N_15105,N_15474);
xor U15824 (N_15824,N_15281,N_15434);
or U15825 (N_15825,N_15214,N_15075);
xnor U15826 (N_15826,N_15154,N_15009);
or U15827 (N_15827,N_15317,N_15320);
and U15828 (N_15828,N_15042,N_15301);
xor U15829 (N_15829,N_15124,N_15249);
and U15830 (N_15830,N_15164,N_15255);
xor U15831 (N_15831,N_15390,N_15341);
or U15832 (N_15832,N_15063,N_15019);
xnor U15833 (N_15833,N_15105,N_15322);
and U15834 (N_15834,N_15003,N_15133);
or U15835 (N_15835,N_15168,N_15353);
or U15836 (N_15836,N_15231,N_15079);
xor U15837 (N_15837,N_15109,N_15188);
nand U15838 (N_15838,N_15279,N_15319);
and U15839 (N_15839,N_15351,N_15043);
and U15840 (N_15840,N_15023,N_15273);
or U15841 (N_15841,N_15496,N_15080);
nand U15842 (N_15842,N_15361,N_15197);
nand U15843 (N_15843,N_15283,N_15106);
nor U15844 (N_15844,N_15499,N_15169);
nand U15845 (N_15845,N_15345,N_15145);
nand U15846 (N_15846,N_15063,N_15191);
xor U15847 (N_15847,N_15055,N_15185);
or U15848 (N_15848,N_15445,N_15272);
and U15849 (N_15849,N_15425,N_15087);
nor U15850 (N_15850,N_15030,N_15027);
and U15851 (N_15851,N_15394,N_15489);
xor U15852 (N_15852,N_15085,N_15044);
nor U15853 (N_15853,N_15295,N_15166);
nand U15854 (N_15854,N_15410,N_15005);
xnor U15855 (N_15855,N_15138,N_15410);
xor U15856 (N_15856,N_15087,N_15370);
and U15857 (N_15857,N_15310,N_15311);
nand U15858 (N_15858,N_15225,N_15058);
or U15859 (N_15859,N_15099,N_15396);
and U15860 (N_15860,N_15386,N_15463);
and U15861 (N_15861,N_15081,N_15008);
or U15862 (N_15862,N_15390,N_15081);
and U15863 (N_15863,N_15009,N_15351);
and U15864 (N_15864,N_15264,N_15359);
and U15865 (N_15865,N_15106,N_15017);
nor U15866 (N_15866,N_15024,N_15174);
nor U15867 (N_15867,N_15465,N_15181);
xor U15868 (N_15868,N_15252,N_15312);
or U15869 (N_15869,N_15142,N_15086);
nand U15870 (N_15870,N_15408,N_15194);
and U15871 (N_15871,N_15083,N_15263);
nor U15872 (N_15872,N_15167,N_15351);
nor U15873 (N_15873,N_15044,N_15154);
and U15874 (N_15874,N_15341,N_15174);
nor U15875 (N_15875,N_15114,N_15393);
nand U15876 (N_15876,N_15287,N_15378);
nor U15877 (N_15877,N_15087,N_15071);
or U15878 (N_15878,N_15420,N_15409);
nor U15879 (N_15879,N_15321,N_15251);
nor U15880 (N_15880,N_15045,N_15469);
and U15881 (N_15881,N_15217,N_15032);
and U15882 (N_15882,N_15279,N_15268);
xnor U15883 (N_15883,N_15157,N_15036);
and U15884 (N_15884,N_15197,N_15415);
nor U15885 (N_15885,N_15149,N_15150);
nand U15886 (N_15886,N_15223,N_15406);
and U15887 (N_15887,N_15065,N_15468);
and U15888 (N_15888,N_15385,N_15495);
nand U15889 (N_15889,N_15087,N_15402);
or U15890 (N_15890,N_15438,N_15064);
and U15891 (N_15891,N_15177,N_15224);
or U15892 (N_15892,N_15488,N_15114);
and U15893 (N_15893,N_15152,N_15087);
xor U15894 (N_15894,N_15485,N_15028);
xnor U15895 (N_15895,N_15457,N_15459);
and U15896 (N_15896,N_15296,N_15453);
xor U15897 (N_15897,N_15002,N_15186);
xor U15898 (N_15898,N_15078,N_15270);
and U15899 (N_15899,N_15158,N_15440);
or U15900 (N_15900,N_15163,N_15314);
xnor U15901 (N_15901,N_15075,N_15341);
nor U15902 (N_15902,N_15278,N_15351);
nand U15903 (N_15903,N_15336,N_15337);
nor U15904 (N_15904,N_15075,N_15081);
nand U15905 (N_15905,N_15108,N_15072);
and U15906 (N_15906,N_15150,N_15286);
nor U15907 (N_15907,N_15324,N_15037);
xor U15908 (N_15908,N_15378,N_15262);
xnor U15909 (N_15909,N_15325,N_15261);
xor U15910 (N_15910,N_15160,N_15042);
nand U15911 (N_15911,N_15468,N_15184);
xor U15912 (N_15912,N_15269,N_15451);
nor U15913 (N_15913,N_15480,N_15426);
or U15914 (N_15914,N_15174,N_15181);
or U15915 (N_15915,N_15337,N_15098);
xnor U15916 (N_15916,N_15299,N_15236);
nand U15917 (N_15917,N_15218,N_15337);
xnor U15918 (N_15918,N_15413,N_15195);
nand U15919 (N_15919,N_15148,N_15242);
nor U15920 (N_15920,N_15334,N_15218);
xnor U15921 (N_15921,N_15126,N_15377);
xnor U15922 (N_15922,N_15093,N_15347);
and U15923 (N_15923,N_15457,N_15004);
and U15924 (N_15924,N_15389,N_15278);
and U15925 (N_15925,N_15189,N_15404);
or U15926 (N_15926,N_15043,N_15405);
nor U15927 (N_15927,N_15007,N_15322);
or U15928 (N_15928,N_15448,N_15431);
or U15929 (N_15929,N_15408,N_15278);
or U15930 (N_15930,N_15242,N_15342);
or U15931 (N_15931,N_15263,N_15000);
nand U15932 (N_15932,N_15165,N_15445);
nor U15933 (N_15933,N_15332,N_15286);
xor U15934 (N_15934,N_15466,N_15387);
nand U15935 (N_15935,N_15091,N_15139);
or U15936 (N_15936,N_15173,N_15360);
nand U15937 (N_15937,N_15049,N_15037);
or U15938 (N_15938,N_15489,N_15156);
nand U15939 (N_15939,N_15348,N_15316);
and U15940 (N_15940,N_15029,N_15241);
nand U15941 (N_15941,N_15097,N_15003);
nor U15942 (N_15942,N_15455,N_15346);
and U15943 (N_15943,N_15484,N_15411);
nor U15944 (N_15944,N_15149,N_15038);
and U15945 (N_15945,N_15044,N_15195);
xnor U15946 (N_15946,N_15373,N_15240);
nand U15947 (N_15947,N_15059,N_15435);
and U15948 (N_15948,N_15186,N_15097);
and U15949 (N_15949,N_15362,N_15446);
nor U15950 (N_15950,N_15457,N_15210);
or U15951 (N_15951,N_15160,N_15071);
xor U15952 (N_15952,N_15383,N_15419);
and U15953 (N_15953,N_15012,N_15136);
nor U15954 (N_15954,N_15488,N_15216);
and U15955 (N_15955,N_15160,N_15238);
xor U15956 (N_15956,N_15082,N_15003);
nor U15957 (N_15957,N_15119,N_15183);
and U15958 (N_15958,N_15479,N_15005);
nand U15959 (N_15959,N_15175,N_15344);
xnor U15960 (N_15960,N_15293,N_15383);
or U15961 (N_15961,N_15450,N_15219);
or U15962 (N_15962,N_15342,N_15466);
and U15963 (N_15963,N_15327,N_15143);
nor U15964 (N_15964,N_15335,N_15060);
and U15965 (N_15965,N_15449,N_15068);
nor U15966 (N_15966,N_15084,N_15055);
and U15967 (N_15967,N_15135,N_15319);
or U15968 (N_15968,N_15380,N_15284);
and U15969 (N_15969,N_15242,N_15203);
and U15970 (N_15970,N_15467,N_15315);
nor U15971 (N_15971,N_15049,N_15359);
nor U15972 (N_15972,N_15100,N_15319);
nand U15973 (N_15973,N_15031,N_15113);
nand U15974 (N_15974,N_15398,N_15294);
nand U15975 (N_15975,N_15119,N_15296);
and U15976 (N_15976,N_15242,N_15184);
or U15977 (N_15977,N_15145,N_15305);
and U15978 (N_15978,N_15136,N_15144);
and U15979 (N_15979,N_15019,N_15304);
xor U15980 (N_15980,N_15213,N_15288);
nand U15981 (N_15981,N_15435,N_15077);
xnor U15982 (N_15982,N_15103,N_15038);
xor U15983 (N_15983,N_15042,N_15136);
or U15984 (N_15984,N_15423,N_15227);
or U15985 (N_15985,N_15064,N_15481);
nor U15986 (N_15986,N_15259,N_15369);
nand U15987 (N_15987,N_15238,N_15153);
nand U15988 (N_15988,N_15189,N_15283);
and U15989 (N_15989,N_15232,N_15408);
nor U15990 (N_15990,N_15066,N_15033);
xnor U15991 (N_15991,N_15409,N_15290);
or U15992 (N_15992,N_15100,N_15394);
and U15993 (N_15993,N_15110,N_15330);
nor U15994 (N_15994,N_15430,N_15194);
nor U15995 (N_15995,N_15081,N_15434);
xnor U15996 (N_15996,N_15148,N_15363);
and U15997 (N_15997,N_15019,N_15071);
or U15998 (N_15998,N_15170,N_15301);
or U15999 (N_15999,N_15308,N_15312);
nor U16000 (N_16000,N_15601,N_15831);
or U16001 (N_16001,N_15584,N_15730);
xnor U16002 (N_16002,N_15942,N_15566);
xor U16003 (N_16003,N_15839,N_15746);
nand U16004 (N_16004,N_15852,N_15548);
nand U16005 (N_16005,N_15983,N_15732);
nand U16006 (N_16006,N_15716,N_15575);
nand U16007 (N_16007,N_15937,N_15874);
and U16008 (N_16008,N_15951,N_15868);
and U16009 (N_16009,N_15914,N_15879);
and U16010 (N_16010,N_15545,N_15603);
or U16011 (N_16011,N_15893,N_15501);
or U16012 (N_16012,N_15948,N_15711);
nand U16013 (N_16013,N_15807,N_15974);
xor U16014 (N_16014,N_15749,N_15761);
or U16015 (N_16015,N_15913,N_15826);
xnor U16016 (N_16016,N_15784,N_15591);
or U16017 (N_16017,N_15519,N_15617);
and U16018 (N_16018,N_15631,N_15981);
and U16019 (N_16019,N_15642,N_15835);
and U16020 (N_16020,N_15938,N_15670);
or U16021 (N_16021,N_15659,N_15768);
nand U16022 (N_16022,N_15629,N_15630);
nor U16023 (N_16023,N_15550,N_15558);
or U16024 (N_16024,N_15907,N_15992);
and U16025 (N_16025,N_15627,N_15635);
and U16026 (N_16026,N_15700,N_15865);
or U16027 (N_16027,N_15602,N_15714);
nor U16028 (N_16028,N_15685,N_15718);
or U16029 (N_16029,N_15564,N_15801);
nand U16030 (N_16030,N_15702,N_15921);
nand U16031 (N_16031,N_15653,N_15890);
and U16032 (N_16032,N_15748,N_15939);
xor U16033 (N_16033,N_15594,N_15604);
and U16034 (N_16034,N_15828,N_15689);
nand U16035 (N_16035,N_15579,N_15583);
or U16036 (N_16036,N_15759,N_15504);
xor U16037 (N_16037,N_15643,N_15817);
or U16038 (N_16038,N_15912,N_15894);
nand U16039 (N_16039,N_15561,N_15725);
nor U16040 (N_16040,N_15962,N_15612);
and U16041 (N_16041,N_15622,N_15798);
and U16042 (N_16042,N_15615,N_15936);
xnor U16043 (N_16043,N_15557,N_15553);
and U16044 (N_16044,N_15915,N_15928);
nor U16045 (N_16045,N_15910,N_15903);
nand U16046 (N_16046,N_15559,N_15726);
xor U16047 (N_16047,N_15616,N_15906);
or U16048 (N_16048,N_15802,N_15818);
and U16049 (N_16049,N_15961,N_15986);
nor U16050 (N_16050,N_15592,N_15620);
nor U16051 (N_16051,N_15509,N_15782);
nand U16052 (N_16052,N_15736,N_15883);
or U16053 (N_16053,N_15896,N_15977);
or U16054 (N_16054,N_15658,N_15537);
xor U16055 (N_16055,N_15972,N_15665);
and U16056 (N_16056,N_15688,N_15934);
nor U16057 (N_16057,N_15675,N_15754);
xnor U16058 (N_16058,N_15901,N_15762);
nor U16059 (N_16059,N_15680,N_15851);
nand U16060 (N_16060,N_15699,N_15984);
nand U16061 (N_16061,N_15854,N_15552);
and U16062 (N_16062,N_15963,N_15857);
xor U16063 (N_16063,N_15861,N_15891);
and U16064 (N_16064,N_15796,N_15527);
and U16065 (N_16065,N_15562,N_15646);
and U16066 (N_16066,N_15554,N_15505);
xor U16067 (N_16067,N_15863,N_15930);
nand U16068 (N_16068,N_15809,N_15990);
or U16069 (N_16069,N_15695,N_15590);
or U16070 (N_16070,N_15995,N_15712);
nand U16071 (N_16071,N_15582,N_15740);
nand U16072 (N_16072,N_15727,N_15880);
nor U16073 (N_16073,N_15728,N_15763);
nor U16074 (N_16074,N_15925,N_15926);
nor U16075 (N_16075,N_15833,N_15780);
and U16076 (N_16076,N_15966,N_15701);
or U16077 (N_16077,N_15531,N_15845);
nor U16078 (N_16078,N_15513,N_15904);
nor U16079 (N_16079,N_15713,N_15989);
or U16080 (N_16080,N_15544,N_15955);
xor U16081 (N_16081,N_15674,N_15998);
nand U16082 (N_16082,N_15767,N_15599);
or U16083 (N_16083,N_15673,N_15556);
nand U16084 (N_16084,N_15797,N_15766);
or U16085 (N_16085,N_15535,N_15706);
nand U16086 (N_16086,N_15508,N_15853);
or U16087 (N_16087,N_15729,N_15538);
and U16088 (N_16088,N_15887,N_15844);
nand U16089 (N_16089,N_15618,N_15855);
nand U16090 (N_16090,N_15967,N_15687);
nand U16091 (N_16091,N_15976,N_15521);
xor U16092 (N_16092,N_15637,N_15908);
nor U16093 (N_16093,N_15794,N_15750);
and U16094 (N_16094,N_15657,N_15682);
nor U16095 (N_16095,N_15841,N_15813);
or U16096 (N_16096,N_15741,N_15656);
and U16097 (N_16097,N_15870,N_15823);
xnor U16098 (N_16098,N_15799,N_15842);
nand U16099 (N_16099,N_15805,N_15626);
or U16100 (N_16100,N_15660,N_15946);
nand U16101 (N_16101,N_15507,N_15572);
xor U16102 (N_16102,N_15968,N_15869);
xor U16103 (N_16103,N_15769,N_15994);
xor U16104 (N_16104,N_15882,N_15683);
nand U16105 (N_16105,N_15884,N_15888);
and U16106 (N_16106,N_15667,N_15957);
xnor U16107 (N_16107,N_15811,N_15708);
nand U16108 (N_16108,N_15668,N_15758);
and U16109 (N_16109,N_15650,N_15776);
or U16110 (N_16110,N_15715,N_15515);
xnor U16111 (N_16111,N_15847,N_15563);
nand U16112 (N_16112,N_15771,N_15677);
and U16113 (N_16113,N_15945,N_15614);
xor U16114 (N_16114,N_15722,N_15875);
nor U16115 (N_16115,N_15530,N_15560);
and U16116 (N_16116,N_15541,N_15574);
nand U16117 (N_16117,N_15787,N_15892);
and U16118 (N_16118,N_15819,N_15581);
xnor U16119 (N_16119,N_15929,N_15671);
nand U16120 (N_16120,N_15628,N_15788);
nand U16121 (N_16121,N_15647,N_15872);
nand U16122 (N_16122,N_15518,N_15640);
xor U16123 (N_16123,N_15589,N_15985);
nand U16124 (N_16124,N_15846,N_15940);
nor U16125 (N_16125,N_15570,N_15920);
nor U16126 (N_16126,N_15860,N_15950);
nor U16127 (N_16127,N_15694,N_15909);
nor U16128 (N_16128,N_15676,N_15911);
xnor U16129 (N_16129,N_15954,N_15607);
and U16130 (N_16130,N_15803,N_15684);
or U16131 (N_16131,N_15760,N_15988);
and U16132 (N_16132,N_15698,N_15943);
and U16133 (N_16133,N_15709,N_15704);
nand U16134 (N_16134,N_15619,N_15533);
xor U16135 (N_16135,N_15597,N_15551);
or U16136 (N_16136,N_15720,N_15822);
nand U16137 (N_16137,N_15745,N_15979);
and U16138 (N_16138,N_15546,N_15997);
nand U16139 (N_16139,N_15806,N_15542);
and U16140 (N_16140,N_15931,N_15625);
xnor U16141 (N_16141,N_15744,N_15662);
xor U16142 (N_16142,N_15516,N_15829);
and U16143 (N_16143,N_15696,N_15850);
xnor U16144 (N_16144,N_15502,N_15710);
or U16145 (N_16145,N_15529,N_15881);
nand U16146 (N_16146,N_15593,N_15751);
and U16147 (N_16147,N_15536,N_15532);
nand U16148 (N_16148,N_15568,N_15905);
and U16149 (N_16149,N_15770,N_15789);
and U16150 (N_16150,N_15827,N_15578);
and U16151 (N_16151,N_15927,N_15836);
or U16152 (N_16152,N_15723,N_15949);
xnor U16153 (N_16153,N_15935,N_15547);
xnor U16154 (N_16154,N_15705,N_15980);
or U16155 (N_16155,N_15539,N_15756);
nand U16156 (N_16156,N_15573,N_15524);
xnor U16157 (N_16157,N_15525,N_15686);
xnor U16158 (N_16158,N_15996,N_15843);
nor U16159 (N_16159,N_15969,N_15774);
nor U16160 (N_16160,N_15987,N_15757);
and U16161 (N_16161,N_15735,N_15795);
and U16162 (N_16162,N_15808,N_15849);
nand U16163 (N_16163,N_15555,N_15793);
and U16164 (N_16164,N_15902,N_15743);
nand U16165 (N_16165,N_15821,N_15786);
nand U16166 (N_16166,N_15644,N_15982);
xnor U16167 (N_16167,N_15565,N_15933);
and U16168 (N_16168,N_15810,N_15960);
nand U16169 (N_16169,N_15523,N_15621);
nor U16170 (N_16170,N_15791,N_15649);
xnor U16171 (N_16171,N_15608,N_15959);
and U16172 (N_16172,N_15632,N_15664);
xor U16173 (N_16173,N_15958,N_15666);
xor U16174 (N_16174,N_15975,N_15520);
nand U16175 (N_16175,N_15923,N_15742);
nand U16176 (N_16176,N_15609,N_15777);
or U16177 (N_16177,N_15611,N_15816);
and U16178 (N_16178,N_15733,N_15956);
xor U16179 (N_16179,N_15889,N_15873);
xor U16180 (N_16180,N_15691,N_15895);
nor U16181 (N_16181,N_15511,N_15679);
nand U16182 (N_16182,N_15834,N_15862);
nor U16183 (N_16183,N_15613,N_15991);
nand U16184 (N_16184,N_15815,N_15899);
nor U16185 (N_16185,N_15540,N_15595);
xnor U16186 (N_16186,N_15528,N_15645);
or U16187 (N_16187,N_15824,N_15648);
or U16188 (N_16188,N_15549,N_15944);
xor U16189 (N_16189,N_15503,N_15871);
nor U16190 (N_16190,N_15719,N_15965);
and U16191 (N_16191,N_15918,N_15624);
and U16192 (N_16192,N_15866,N_15898);
nand U16193 (N_16193,N_15970,N_15753);
and U16194 (N_16194,N_15772,N_15993);
or U16195 (N_16195,N_15858,N_15814);
nor U16196 (N_16196,N_15707,N_15623);
nand U16197 (N_16197,N_15678,N_15971);
and U16198 (N_16198,N_15752,N_15681);
and U16199 (N_16199,N_15669,N_15697);
and U16200 (N_16200,N_15577,N_15885);
and U16201 (N_16201,N_15917,N_15932);
nand U16202 (N_16202,N_15543,N_15778);
nand U16203 (N_16203,N_15978,N_15651);
nor U16204 (N_16204,N_15764,N_15999);
and U16205 (N_16205,N_15878,N_15500);
xor U16206 (N_16206,N_15634,N_15567);
nand U16207 (N_16207,N_15877,N_15598);
xor U16208 (N_16208,N_15897,N_15947);
nor U16209 (N_16209,N_15569,N_15526);
xnor U16210 (N_16210,N_15717,N_15864);
nor U16211 (N_16211,N_15941,N_15692);
nand U16212 (N_16212,N_15840,N_15731);
nor U16213 (N_16213,N_15587,N_15639);
and U16214 (N_16214,N_15781,N_15517);
or U16215 (N_16215,N_15641,N_15922);
or U16216 (N_16216,N_15867,N_15652);
nor U16217 (N_16217,N_15952,N_15876);
or U16218 (N_16218,N_15605,N_15973);
and U16219 (N_16219,N_15506,N_15953);
xnor U16220 (N_16220,N_15747,N_15916);
or U16221 (N_16221,N_15690,N_15721);
and U16222 (N_16222,N_15832,N_15633);
and U16223 (N_16223,N_15783,N_15663);
and U16224 (N_16224,N_15512,N_15661);
or U16225 (N_16225,N_15734,N_15800);
and U16226 (N_16226,N_15654,N_15785);
or U16227 (N_16227,N_15724,N_15576);
nand U16228 (N_16228,N_15765,N_15775);
and U16229 (N_16229,N_15886,N_15606);
and U16230 (N_16230,N_15790,N_15859);
xnor U16231 (N_16231,N_15773,N_15825);
xor U16232 (N_16232,N_15514,N_15534);
nor U16233 (N_16233,N_15596,N_15755);
xnor U16234 (N_16234,N_15655,N_15820);
nor U16235 (N_16235,N_15600,N_15703);
nand U16236 (N_16236,N_15856,N_15571);
and U16237 (N_16237,N_15919,N_15522);
nand U16238 (N_16238,N_15792,N_15738);
or U16239 (N_16239,N_15693,N_15672);
and U16240 (N_16240,N_15739,N_15830);
nor U16241 (N_16241,N_15585,N_15924);
xor U16242 (N_16242,N_15610,N_15737);
or U16243 (N_16243,N_15838,N_15812);
or U16244 (N_16244,N_15804,N_15638);
or U16245 (N_16245,N_15779,N_15837);
or U16246 (N_16246,N_15510,N_15848);
xor U16247 (N_16247,N_15588,N_15900);
or U16248 (N_16248,N_15580,N_15636);
xnor U16249 (N_16249,N_15964,N_15586);
nand U16250 (N_16250,N_15630,N_15685);
or U16251 (N_16251,N_15697,N_15521);
xnor U16252 (N_16252,N_15808,N_15794);
nand U16253 (N_16253,N_15642,N_15750);
or U16254 (N_16254,N_15639,N_15730);
nor U16255 (N_16255,N_15601,N_15568);
and U16256 (N_16256,N_15746,N_15718);
or U16257 (N_16257,N_15992,N_15958);
nor U16258 (N_16258,N_15801,N_15893);
or U16259 (N_16259,N_15726,N_15758);
and U16260 (N_16260,N_15768,N_15706);
nor U16261 (N_16261,N_15811,N_15501);
or U16262 (N_16262,N_15514,N_15932);
xnor U16263 (N_16263,N_15588,N_15562);
xor U16264 (N_16264,N_15802,N_15585);
nor U16265 (N_16265,N_15894,N_15727);
nor U16266 (N_16266,N_15864,N_15566);
or U16267 (N_16267,N_15653,N_15782);
nor U16268 (N_16268,N_15575,N_15948);
and U16269 (N_16269,N_15656,N_15633);
and U16270 (N_16270,N_15740,N_15542);
nand U16271 (N_16271,N_15597,N_15592);
or U16272 (N_16272,N_15979,N_15771);
and U16273 (N_16273,N_15843,N_15826);
nand U16274 (N_16274,N_15685,N_15514);
nand U16275 (N_16275,N_15867,N_15900);
nor U16276 (N_16276,N_15865,N_15590);
and U16277 (N_16277,N_15503,N_15727);
nand U16278 (N_16278,N_15673,N_15711);
and U16279 (N_16279,N_15719,N_15733);
and U16280 (N_16280,N_15643,N_15710);
nor U16281 (N_16281,N_15509,N_15838);
xnor U16282 (N_16282,N_15736,N_15608);
and U16283 (N_16283,N_15504,N_15525);
nand U16284 (N_16284,N_15565,N_15641);
and U16285 (N_16285,N_15665,N_15987);
or U16286 (N_16286,N_15819,N_15835);
and U16287 (N_16287,N_15909,N_15637);
and U16288 (N_16288,N_15566,N_15687);
nor U16289 (N_16289,N_15899,N_15744);
nor U16290 (N_16290,N_15632,N_15703);
nor U16291 (N_16291,N_15582,N_15842);
xnor U16292 (N_16292,N_15544,N_15704);
nand U16293 (N_16293,N_15546,N_15799);
xnor U16294 (N_16294,N_15917,N_15957);
nor U16295 (N_16295,N_15572,N_15711);
or U16296 (N_16296,N_15966,N_15749);
and U16297 (N_16297,N_15679,N_15965);
nand U16298 (N_16298,N_15981,N_15945);
xnor U16299 (N_16299,N_15716,N_15786);
and U16300 (N_16300,N_15922,N_15804);
and U16301 (N_16301,N_15595,N_15808);
or U16302 (N_16302,N_15902,N_15857);
or U16303 (N_16303,N_15695,N_15507);
or U16304 (N_16304,N_15813,N_15866);
xnor U16305 (N_16305,N_15747,N_15796);
or U16306 (N_16306,N_15870,N_15951);
or U16307 (N_16307,N_15553,N_15661);
xnor U16308 (N_16308,N_15578,N_15969);
and U16309 (N_16309,N_15837,N_15519);
nor U16310 (N_16310,N_15755,N_15820);
nand U16311 (N_16311,N_15636,N_15682);
nor U16312 (N_16312,N_15784,N_15557);
and U16313 (N_16313,N_15705,N_15541);
or U16314 (N_16314,N_15616,N_15773);
xor U16315 (N_16315,N_15685,N_15785);
nand U16316 (N_16316,N_15655,N_15572);
or U16317 (N_16317,N_15888,N_15675);
or U16318 (N_16318,N_15519,N_15649);
nand U16319 (N_16319,N_15588,N_15949);
nor U16320 (N_16320,N_15568,N_15735);
or U16321 (N_16321,N_15798,N_15831);
and U16322 (N_16322,N_15846,N_15671);
nand U16323 (N_16323,N_15964,N_15527);
or U16324 (N_16324,N_15692,N_15891);
nor U16325 (N_16325,N_15688,N_15732);
or U16326 (N_16326,N_15694,N_15780);
and U16327 (N_16327,N_15519,N_15906);
and U16328 (N_16328,N_15894,N_15679);
nor U16329 (N_16329,N_15990,N_15774);
and U16330 (N_16330,N_15726,N_15707);
or U16331 (N_16331,N_15532,N_15535);
or U16332 (N_16332,N_15889,N_15823);
xor U16333 (N_16333,N_15716,N_15515);
xor U16334 (N_16334,N_15645,N_15569);
and U16335 (N_16335,N_15526,N_15584);
nor U16336 (N_16336,N_15579,N_15601);
or U16337 (N_16337,N_15725,N_15931);
or U16338 (N_16338,N_15759,N_15644);
nor U16339 (N_16339,N_15715,N_15735);
or U16340 (N_16340,N_15568,N_15878);
or U16341 (N_16341,N_15919,N_15805);
xor U16342 (N_16342,N_15656,N_15623);
or U16343 (N_16343,N_15962,N_15879);
or U16344 (N_16344,N_15838,N_15949);
xor U16345 (N_16345,N_15714,N_15924);
and U16346 (N_16346,N_15560,N_15744);
nor U16347 (N_16347,N_15732,N_15876);
nand U16348 (N_16348,N_15934,N_15738);
and U16349 (N_16349,N_15947,N_15704);
nand U16350 (N_16350,N_15588,N_15635);
xnor U16351 (N_16351,N_15960,N_15883);
nor U16352 (N_16352,N_15570,N_15798);
nor U16353 (N_16353,N_15594,N_15630);
nor U16354 (N_16354,N_15982,N_15774);
or U16355 (N_16355,N_15885,N_15792);
nor U16356 (N_16356,N_15533,N_15514);
nor U16357 (N_16357,N_15736,N_15807);
nand U16358 (N_16358,N_15623,N_15586);
nor U16359 (N_16359,N_15971,N_15754);
or U16360 (N_16360,N_15993,N_15886);
nor U16361 (N_16361,N_15612,N_15933);
or U16362 (N_16362,N_15989,N_15531);
and U16363 (N_16363,N_15949,N_15505);
or U16364 (N_16364,N_15852,N_15970);
and U16365 (N_16365,N_15572,N_15802);
nand U16366 (N_16366,N_15656,N_15812);
nor U16367 (N_16367,N_15857,N_15638);
or U16368 (N_16368,N_15866,N_15618);
nand U16369 (N_16369,N_15939,N_15694);
and U16370 (N_16370,N_15813,N_15653);
and U16371 (N_16371,N_15578,N_15789);
or U16372 (N_16372,N_15782,N_15903);
nor U16373 (N_16373,N_15563,N_15719);
nand U16374 (N_16374,N_15757,N_15634);
and U16375 (N_16375,N_15722,N_15950);
and U16376 (N_16376,N_15727,N_15711);
and U16377 (N_16377,N_15677,N_15856);
and U16378 (N_16378,N_15800,N_15572);
xor U16379 (N_16379,N_15697,N_15961);
nand U16380 (N_16380,N_15579,N_15705);
nand U16381 (N_16381,N_15903,N_15743);
or U16382 (N_16382,N_15944,N_15959);
or U16383 (N_16383,N_15978,N_15773);
xor U16384 (N_16384,N_15514,N_15634);
and U16385 (N_16385,N_15889,N_15895);
xnor U16386 (N_16386,N_15979,N_15973);
xnor U16387 (N_16387,N_15782,N_15858);
and U16388 (N_16388,N_15664,N_15571);
and U16389 (N_16389,N_15822,N_15890);
and U16390 (N_16390,N_15632,N_15914);
nand U16391 (N_16391,N_15563,N_15567);
or U16392 (N_16392,N_15812,N_15865);
and U16393 (N_16393,N_15725,N_15685);
nor U16394 (N_16394,N_15743,N_15706);
xor U16395 (N_16395,N_15921,N_15518);
and U16396 (N_16396,N_15625,N_15783);
or U16397 (N_16397,N_15898,N_15834);
nor U16398 (N_16398,N_15511,N_15876);
xnor U16399 (N_16399,N_15708,N_15772);
and U16400 (N_16400,N_15576,N_15569);
or U16401 (N_16401,N_15707,N_15593);
nor U16402 (N_16402,N_15703,N_15572);
xor U16403 (N_16403,N_15731,N_15883);
xor U16404 (N_16404,N_15683,N_15875);
and U16405 (N_16405,N_15648,N_15680);
xor U16406 (N_16406,N_15701,N_15990);
xor U16407 (N_16407,N_15753,N_15587);
nor U16408 (N_16408,N_15745,N_15940);
nand U16409 (N_16409,N_15830,N_15623);
and U16410 (N_16410,N_15603,N_15692);
or U16411 (N_16411,N_15840,N_15650);
or U16412 (N_16412,N_15965,N_15553);
xor U16413 (N_16413,N_15952,N_15548);
nand U16414 (N_16414,N_15520,N_15551);
and U16415 (N_16415,N_15846,N_15668);
xor U16416 (N_16416,N_15583,N_15849);
nand U16417 (N_16417,N_15659,N_15512);
or U16418 (N_16418,N_15771,N_15724);
nand U16419 (N_16419,N_15633,N_15693);
nand U16420 (N_16420,N_15594,N_15685);
and U16421 (N_16421,N_15847,N_15696);
xor U16422 (N_16422,N_15610,N_15992);
nor U16423 (N_16423,N_15750,N_15804);
and U16424 (N_16424,N_15745,N_15855);
nor U16425 (N_16425,N_15572,N_15674);
or U16426 (N_16426,N_15756,N_15726);
nand U16427 (N_16427,N_15694,N_15781);
nor U16428 (N_16428,N_15796,N_15750);
nor U16429 (N_16429,N_15988,N_15678);
xnor U16430 (N_16430,N_15932,N_15896);
nor U16431 (N_16431,N_15606,N_15779);
nor U16432 (N_16432,N_15982,N_15504);
and U16433 (N_16433,N_15842,N_15551);
nor U16434 (N_16434,N_15523,N_15851);
or U16435 (N_16435,N_15687,N_15780);
or U16436 (N_16436,N_15863,N_15655);
nor U16437 (N_16437,N_15623,N_15908);
nor U16438 (N_16438,N_15787,N_15537);
xor U16439 (N_16439,N_15984,N_15727);
and U16440 (N_16440,N_15680,N_15968);
and U16441 (N_16441,N_15986,N_15876);
nand U16442 (N_16442,N_15655,N_15940);
nand U16443 (N_16443,N_15966,N_15930);
nand U16444 (N_16444,N_15882,N_15690);
nor U16445 (N_16445,N_15948,N_15799);
and U16446 (N_16446,N_15506,N_15589);
or U16447 (N_16447,N_15535,N_15696);
xor U16448 (N_16448,N_15572,N_15549);
nor U16449 (N_16449,N_15774,N_15930);
and U16450 (N_16450,N_15698,N_15530);
and U16451 (N_16451,N_15782,N_15799);
and U16452 (N_16452,N_15629,N_15770);
or U16453 (N_16453,N_15878,N_15717);
and U16454 (N_16454,N_15952,N_15532);
xnor U16455 (N_16455,N_15716,N_15610);
or U16456 (N_16456,N_15590,N_15734);
and U16457 (N_16457,N_15821,N_15647);
and U16458 (N_16458,N_15901,N_15888);
nand U16459 (N_16459,N_15906,N_15967);
nand U16460 (N_16460,N_15560,N_15631);
xnor U16461 (N_16461,N_15761,N_15805);
xor U16462 (N_16462,N_15679,N_15861);
nand U16463 (N_16463,N_15894,N_15516);
and U16464 (N_16464,N_15713,N_15650);
xnor U16465 (N_16465,N_15583,N_15944);
or U16466 (N_16466,N_15665,N_15670);
nand U16467 (N_16467,N_15900,N_15544);
and U16468 (N_16468,N_15696,N_15725);
nand U16469 (N_16469,N_15667,N_15688);
or U16470 (N_16470,N_15991,N_15901);
and U16471 (N_16471,N_15797,N_15854);
or U16472 (N_16472,N_15957,N_15993);
and U16473 (N_16473,N_15950,N_15951);
xnor U16474 (N_16474,N_15977,N_15716);
nor U16475 (N_16475,N_15777,N_15907);
and U16476 (N_16476,N_15850,N_15526);
nand U16477 (N_16477,N_15812,N_15891);
and U16478 (N_16478,N_15880,N_15675);
xor U16479 (N_16479,N_15719,N_15649);
xnor U16480 (N_16480,N_15697,N_15843);
nor U16481 (N_16481,N_15963,N_15600);
or U16482 (N_16482,N_15916,N_15850);
nand U16483 (N_16483,N_15767,N_15937);
nand U16484 (N_16484,N_15571,N_15735);
xnor U16485 (N_16485,N_15673,N_15625);
or U16486 (N_16486,N_15789,N_15597);
and U16487 (N_16487,N_15891,N_15642);
and U16488 (N_16488,N_15915,N_15878);
nand U16489 (N_16489,N_15878,N_15929);
nand U16490 (N_16490,N_15714,N_15973);
nand U16491 (N_16491,N_15679,N_15751);
xnor U16492 (N_16492,N_15810,N_15906);
nor U16493 (N_16493,N_15818,N_15829);
nand U16494 (N_16494,N_15962,N_15972);
nand U16495 (N_16495,N_15914,N_15679);
and U16496 (N_16496,N_15713,N_15778);
xnor U16497 (N_16497,N_15930,N_15847);
and U16498 (N_16498,N_15961,N_15644);
nand U16499 (N_16499,N_15849,N_15983);
nand U16500 (N_16500,N_16452,N_16447);
xnor U16501 (N_16501,N_16275,N_16337);
nand U16502 (N_16502,N_16062,N_16176);
or U16503 (N_16503,N_16123,N_16496);
and U16504 (N_16504,N_16222,N_16201);
and U16505 (N_16505,N_16375,N_16475);
nor U16506 (N_16506,N_16157,N_16048);
or U16507 (N_16507,N_16122,N_16465);
nor U16508 (N_16508,N_16232,N_16033);
and U16509 (N_16509,N_16369,N_16494);
xnor U16510 (N_16510,N_16329,N_16274);
nor U16511 (N_16511,N_16249,N_16117);
and U16512 (N_16512,N_16282,N_16046);
and U16513 (N_16513,N_16394,N_16011);
nor U16514 (N_16514,N_16351,N_16059);
xnor U16515 (N_16515,N_16445,N_16039);
nor U16516 (N_16516,N_16359,N_16199);
xor U16517 (N_16517,N_16373,N_16102);
and U16518 (N_16518,N_16243,N_16271);
nor U16519 (N_16519,N_16185,N_16081);
or U16520 (N_16520,N_16101,N_16418);
and U16521 (N_16521,N_16365,N_16319);
or U16522 (N_16522,N_16367,N_16245);
xor U16523 (N_16523,N_16323,N_16404);
nand U16524 (N_16524,N_16118,N_16137);
nand U16525 (N_16525,N_16415,N_16435);
or U16526 (N_16526,N_16024,N_16175);
xnor U16527 (N_16527,N_16299,N_16053);
and U16528 (N_16528,N_16170,N_16076);
and U16529 (N_16529,N_16142,N_16135);
nand U16530 (N_16530,N_16023,N_16128);
and U16531 (N_16531,N_16223,N_16090);
nand U16532 (N_16532,N_16491,N_16110);
nor U16533 (N_16533,N_16001,N_16289);
nand U16534 (N_16534,N_16200,N_16013);
nand U16535 (N_16535,N_16119,N_16397);
xnor U16536 (N_16536,N_16487,N_16019);
nand U16537 (N_16537,N_16092,N_16287);
nor U16538 (N_16538,N_16253,N_16309);
nand U16539 (N_16539,N_16348,N_16094);
nand U16540 (N_16540,N_16156,N_16058);
or U16541 (N_16541,N_16111,N_16332);
nand U16542 (N_16542,N_16364,N_16313);
nor U16543 (N_16543,N_16462,N_16043);
and U16544 (N_16544,N_16100,N_16163);
nor U16545 (N_16545,N_16458,N_16261);
and U16546 (N_16546,N_16315,N_16455);
nor U16547 (N_16547,N_16012,N_16064);
nand U16548 (N_16548,N_16207,N_16103);
nand U16549 (N_16549,N_16036,N_16326);
nor U16550 (N_16550,N_16027,N_16010);
nand U16551 (N_16551,N_16087,N_16008);
nor U16552 (N_16552,N_16352,N_16162);
nand U16553 (N_16553,N_16390,N_16318);
nand U16554 (N_16554,N_16000,N_16141);
xnor U16555 (N_16555,N_16400,N_16338);
nor U16556 (N_16556,N_16166,N_16035);
and U16557 (N_16557,N_16218,N_16264);
or U16558 (N_16558,N_16234,N_16386);
nand U16559 (N_16559,N_16003,N_16448);
and U16560 (N_16560,N_16235,N_16181);
nor U16561 (N_16561,N_16335,N_16422);
xor U16562 (N_16562,N_16481,N_16247);
and U16563 (N_16563,N_16417,N_16290);
and U16564 (N_16564,N_16263,N_16120);
and U16565 (N_16565,N_16099,N_16252);
nand U16566 (N_16566,N_16322,N_16408);
nor U16567 (N_16567,N_16317,N_16380);
xor U16568 (N_16568,N_16073,N_16196);
and U16569 (N_16569,N_16072,N_16440);
or U16570 (N_16570,N_16211,N_16026);
nor U16571 (N_16571,N_16069,N_16421);
or U16572 (N_16572,N_16324,N_16344);
and U16573 (N_16573,N_16083,N_16231);
xnor U16574 (N_16574,N_16066,N_16198);
and U16575 (N_16575,N_16442,N_16437);
or U16576 (N_16576,N_16341,N_16186);
or U16577 (N_16577,N_16124,N_16457);
xor U16578 (N_16578,N_16071,N_16424);
nand U16579 (N_16579,N_16106,N_16431);
nor U16580 (N_16580,N_16333,N_16041);
nor U16581 (N_16581,N_16342,N_16314);
or U16582 (N_16582,N_16070,N_16398);
nor U16583 (N_16583,N_16444,N_16038);
xor U16584 (N_16584,N_16302,N_16089);
nor U16585 (N_16585,N_16349,N_16460);
and U16586 (N_16586,N_16391,N_16149);
nor U16587 (N_16587,N_16086,N_16433);
xor U16588 (N_16588,N_16405,N_16480);
nor U16589 (N_16589,N_16063,N_16187);
nor U16590 (N_16590,N_16206,N_16273);
nand U16591 (N_16591,N_16214,N_16055);
nor U16592 (N_16592,N_16096,N_16009);
nand U16593 (N_16593,N_16340,N_16169);
nand U16594 (N_16594,N_16416,N_16014);
and U16595 (N_16595,N_16459,N_16125);
or U16596 (N_16596,N_16174,N_16469);
and U16597 (N_16597,N_16130,N_16229);
nor U16598 (N_16598,N_16188,N_16366);
xor U16599 (N_16599,N_16280,N_16242);
nor U16600 (N_16600,N_16297,N_16401);
or U16601 (N_16601,N_16184,N_16042);
nor U16602 (N_16602,N_16197,N_16138);
or U16603 (N_16603,N_16237,N_16032);
nor U16604 (N_16604,N_16483,N_16443);
nand U16605 (N_16605,N_16116,N_16387);
nor U16606 (N_16606,N_16126,N_16230);
xor U16607 (N_16607,N_16370,N_16361);
nor U16608 (N_16608,N_16093,N_16121);
or U16609 (N_16609,N_16461,N_16078);
xor U16610 (N_16610,N_16220,N_16224);
nor U16611 (N_16611,N_16429,N_16129);
nor U16612 (N_16612,N_16478,N_16152);
xor U16613 (N_16613,N_16489,N_16392);
and U16614 (N_16614,N_16383,N_16419);
xor U16615 (N_16615,N_16148,N_16316);
or U16616 (N_16616,N_16473,N_16388);
nor U16617 (N_16617,N_16015,N_16239);
nand U16618 (N_16618,N_16384,N_16004);
xor U16619 (N_16619,N_16449,N_16258);
nand U16620 (N_16620,N_16044,N_16250);
and U16621 (N_16621,N_16212,N_16493);
and U16622 (N_16622,N_16131,N_16031);
and U16623 (N_16623,N_16262,N_16045);
and U16624 (N_16624,N_16077,N_16283);
nand U16625 (N_16625,N_16407,N_16439);
or U16626 (N_16626,N_16084,N_16293);
and U16627 (N_16627,N_16021,N_16269);
and U16628 (N_16628,N_16098,N_16385);
or U16629 (N_16629,N_16238,N_16029);
nor U16630 (N_16630,N_16007,N_16311);
nand U16631 (N_16631,N_16018,N_16298);
xnor U16632 (N_16632,N_16074,N_16466);
nand U16633 (N_16633,N_16410,N_16147);
xnor U16634 (N_16634,N_16037,N_16436);
xnor U16635 (N_16635,N_16272,N_16374);
and U16636 (N_16636,N_16260,N_16372);
nor U16637 (N_16637,N_16056,N_16371);
or U16638 (N_16638,N_16308,N_16345);
xnor U16639 (N_16639,N_16158,N_16307);
xor U16640 (N_16640,N_16217,N_16306);
xor U16641 (N_16641,N_16267,N_16379);
and U16642 (N_16642,N_16355,N_16434);
xor U16643 (N_16643,N_16266,N_16358);
nand U16644 (N_16644,N_16143,N_16017);
nand U16645 (N_16645,N_16310,N_16301);
nor U16646 (N_16646,N_16403,N_16294);
nand U16647 (N_16647,N_16040,N_16277);
and U16648 (N_16648,N_16104,N_16382);
nand U16649 (N_16649,N_16192,N_16080);
nand U16650 (N_16650,N_16381,N_16168);
xnor U16651 (N_16651,N_16068,N_16492);
nor U16652 (N_16652,N_16303,N_16354);
and U16653 (N_16653,N_16225,N_16346);
xnor U16654 (N_16654,N_16414,N_16095);
nand U16655 (N_16655,N_16105,N_16179);
xnor U16656 (N_16656,N_16164,N_16278);
and U16657 (N_16657,N_16088,N_16482);
or U16658 (N_16658,N_16476,N_16360);
and U16659 (N_16659,N_16296,N_16195);
and U16660 (N_16660,N_16304,N_16079);
nor U16661 (N_16661,N_16336,N_16114);
xor U16662 (N_16662,N_16171,N_16050);
nand U16663 (N_16663,N_16497,N_16210);
or U16664 (N_16664,N_16155,N_16178);
xor U16665 (N_16665,N_16312,N_16109);
xor U16666 (N_16666,N_16057,N_16172);
xor U16667 (N_16667,N_16488,N_16464);
xnor U16668 (N_16668,N_16474,N_16331);
or U16669 (N_16669,N_16065,N_16446);
xnor U16670 (N_16670,N_16305,N_16426);
nand U16671 (N_16671,N_16291,N_16165);
xor U16672 (N_16672,N_16256,N_16226);
nor U16673 (N_16673,N_16159,N_16353);
xor U16674 (N_16674,N_16328,N_16281);
nor U16675 (N_16675,N_16265,N_16276);
xnor U16676 (N_16676,N_16485,N_16194);
and U16677 (N_16677,N_16246,N_16052);
nor U16678 (N_16678,N_16115,N_16241);
or U16679 (N_16679,N_16216,N_16425);
or U16680 (N_16680,N_16049,N_16451);
and U16681 (N_16681,N_16413,N_16132);
nor U16682 (N_16682,N_16054,N_16396);
xor U16683 (N_16683,N_16005,N_16362);
xor U16684 (N_16684,N_16034,N_16288);
nand U16685 (N_16685,N_16209,N_16330);
xor U16686 (N_16686,N_16020,N_16472);
xnor U16687 (N_16687,N_16395,N_16183);
nor U16688 (N_16688,N_16204,N_16484);
nor U16689 (N_16689,N_16409,N_16161);
xor U16690 (N_16690,N_16240,N_16471);
and U16691 (N_16691,N_16180,N_16146);
and U16692 (N_16692,N_16325,N_16219);
and U16693 (N_16693,N_16423,N_16002);
nand U16694 (N_16694,N_16479,N_16393);
nand U16695 (N_16695,N_16368,N_16025);
nand U16696 (N_16696,N_16430,N_16327);
and U16697 (N_16697,N_16486,N_16270);
xor U16698 (N_16698,N_16160,N_16082);
nand U16699 (N_16699,N_16127,N_16300);
nand U16700 (N_16700,N_16259,N_16402);
xnor U16701 (N_16701,N_16467,N_16406);
or U16702 (N_16702,N_16133,N_16279);
xor U16703 (N_16703,N_16295,N_16182);
xor U16704 (N_16704,N_16257,N_16244);
and U16705 (N_16705,N_16075,N_16499);
and U16706 (N_16706,N_16051,N_16347);
xnor U16707 (N_16707,N_16399,N_16215);
xor U16708 (N_16708,N_16498,N_16228);
nand U16709 (N_16709,N_16006,N_16251);
nor U16710 (N_16710,N_16134,N_16173);
and U16711 (N_16711,N_16468,N_16284);
nand U16712 (N_16712,N_16420,N_16236);
or U16713 (N_16713,N_16470,N_16193);
and U16714 (N_16714,N_16136,N_16190);
and U16715 (N_16715,N_16463,N_16213);
and U16716 (N_16716,N_16067,N_16097);
xnor U16717 (N_16717,N_16016,N_16203);
xor U16718 (N_16718,N_16233,N_16357);
or U16719 (N_16719,N_16438,N_16060);
or U16720 (N_16720,N_16144,N_16145);
and U16721 (N_16721,N_16085,N_16150);
nand U16722 (N_16722,N_16450,N_16022);
xor U16723 (N_16723,N_16107,N_16208);
xor U16724 (N_16724,N_16113,N_16140);
and U16725 (N_16725,N_16292,N_16167);
xnor U16726 (N_16726,N_16454,N_16320);
or U16727 (N_16727,N_16376,N_16453);
nor U16728 (N_16728,N_16412,N_16378);
nor U16729 (N_16729,N_16177,N_16248);
nor U16730 (N_16730,N_16411,N_16030);
or U16731 (N_16731,N_16321,N_16028);
and U16732 (N_16732,N_16334,N_16427);
xnor U16733 (N_16733,N_16490,N_16151);
nor U16734 (N_16734,N_16227,N_16154);
nand U16735 (N_16735,N_16091,N_16356);
and U16736 (N_16736,N_16495,N_16432);
or U16737 (N_16737,N_16268,N_16254);
xnor U16738 (N_16738,N_16112,N_16047);
or U16739 (N_16739,N_16061,N_16389);
nor U16740 (N_16740,N_16286,N_16221);
xnor U16741 (N_16741,N_16205,N_16153);
nand U16742 (N_16742,N_16477,N_16191);
or U16743 (N_16743,N_16456,N_16202);
xor U16744 (N_16744,N_16139,N_16350);
nor U16745 (N_16745,N_16363,N_16255);
nand U16746 (N_16746,N_16343,N_16428);
xor U16747 (N_16747,N_16377,N_16339);
nand U16748 (N_16748,N_16441,N_16189);
nand U16749 (N_16749,N_16285,N_16108);
nand U16750 (N_16750,N_16087,N_16294);
and U16751 (N_16751,N_16203,N_16488);
nor U16752 (N_16752,N_16288,N_16385);
xor U16753 (N_16753,N_16370,N_16020);
nor U16754 (N_16754,N_16435,N_16287);
and U16755 (N_16755,N_16133,N_16125);
nor U16756 (N_16756,N_16498,N_16404);
or U16757 (N_16757,N_16341,N_16316);
nand U16758 (N_16758,N_16430,N_16467);
xor U16759 (N_16759,N_16452,N_16297);
and U16760 (N_16760,N_16048,N_16457);
nor U16761 (N_16761,N_16027,N_16375);
or U16762 (N_16762,N_16295,N_16395);
or U16763 (N_16763,N_16155,N_16397);
nor U16764 (N_16764,N_16098,N_16398);
nand U16765 (N_16765,N_16319,N_16368);
and U16766 (N_16766,N_16459,N_16463);
nand U16767 (N_16767,N_16107,N_16165);
nand U16768 (N_16768,N_16188,N_16126);
nand U16769 (N_16769,N_16402,N_16049);
nor U16770 (N_16770,N_16045,N_16114);
nand U16771 (N_16771,N_16391,N_16406);
and U16772 (N_16772,N_16477,N_16158);
or U16773 (N_16773,N_16376,N_16484);
nand U16774 (N_16774,N_16400,N_16462);
and U16775 (N_16775,N_16116,N_16173);
xor U16776 (N_16776,N_16344,N_16210);
and U16777 (N_16777,N_16466,N_16027);
xor U16778 (N_16778,N_16461,N_16103);
and U16779 (N_16779,N_16475,N_16040);
and U16780 (N_16780,N_16466,N_16161);
nand U16781 (N_16781,N_16067,N_16292);
xnor U16782 (N_16782,N_16042,N_16256);
nand U16783 (N_16783,N_16285,N_16005);
nor U16784 (N_16784,N_16177,N_16314);
xor U16785 (N_16785,N_16398,N_16353);
nor U16786 (N_16786,N_16367,N_16274);
or U16787 (N_16787,N_16248,N_16011);
xor U16788 (N_16788,N_16406,N_16054);
or U16789 (N_16789,N_16243,N_16445);
xnor U16790 (N_16790,N_16442,N_16156);
nand U16791 (N_16791,N_16209,N_16476);
nand U16792 (N_16792,N_16364,N_16081);
nor U16793 (N_16793,N_16444,N_16014);
nor U16794 (N_16794,N_16491,N_16208);
xor U16795 (N_16795,N_16358,N_16036);
xnor U16796 (N_16796,N_16284,N_16479);
xor U16797 (N_16797,N_16342,N_16265);
nand U16798 (N_16798,N_16251,N_16118);
or U16799 (N_16799,N_16271,N_16075);
xor U16800 (N_16800,N_16312,N_16260);
and U16801 (N_16801,N_16173,N_16386);
and U16802 (N_16802,N_16432,N_16425);
nor U16803 (N_16803,N_16108,N_16380);
xor U16804 (N_16804,N_16085,N_16342);
and U16805 (N_16805,N_16245,N_16321);
xor U16806 (N_16806,N_16157,N_16487);
nand U16807 (N_16807,N_16230,N_16006);
and U16808 (N_16808,N_16260,N_16382);
xnor U16809 (N_16809,N_16168,N_16191);
nor U16810 (N_16810,N_16298,N_16471);
and U16811 (N_16811,N_16237,N_16047);
or U16812 (N_16812,N_16048,N_16086);
nand U16813 (N_16813,N_16045,N_16142);
or U16814 (N_16814,N_16050,N_16163);
nand U16815 (N_16815,N_16130,N_16330);
nor U16816 (N_16816,N_16130,N_16422);
xnor U16817 (N_16817,N_16384,N_16100);
nand U16818 (N_16818,N_16214,N_16116);
xnor U16819 (N_16819,N_16443,N_16099);
or U16820 (N_16820,N_16238,N_16447);
nor U16821 (N_16821,N_16230,N_16185);
or U16822 (N_16822,N_16035,N_16364);
nor U16823 (N_16823,N_16289,N_16266);
and U16824 (N_16824,N_16190,N_16161);
nand U16825 (N_16825,N_16020,N_16368);
xor U16826 (N_16826,N_16335,N_16128);
nor U16827 (N_16827,N_16466,N_16146);
or U16828 (N_16828,N_16306,N_16493);
nor U16829 (N_16829,N_16312,N_16342);
xnor U16830 (N_16830,N_16356,N_16005);
xnor U16831 (N_16831,N_16421,N_16255);
xor U16832 (N_16832,N_16185,N_16359);
and U16833 (N_16833,N_16496,N_16192);
nor U16834 (N_16834,N_16475,N_16394);
xnor U16835 (N_16835,N_16492,N_16398);
xor U16836 (N_16836,N_16342,N_16480);
or U16837 (N_16837,N_16150,N_16456);
and U16838 (N_16838,N_16308,N_16083);
or U16839 (N_16839,N_16430,N_16421);
nand U16840 (N_16840,N_16418,N_16397);
or U16841 (N_16841,N_16173,N_16442);
xor U16842 (N_16842,N_16314,N_16052);
xnor U16843 (N_16843,N_16385,N_16071);
nor U16844 (N_16844,N_16406,N_16296);
and U16845 (N_16845,N_16328,N_16441);
xor U16846 (N_16846,N_16248,N_16423);
and U16847 (N_16847,N_16283,N_16387);
nor U16848 (N_16848,N_16021,N_16158);
nand U16849 (N_16849,N_16096,N_16034);
nor U16850 (N_16850,N_16207,N_16184);
nor U16851 (N_16851,N_16017,N_16326);
nand U16852 (N_16852,N_16270,N_16113);
xor U16853 (N_16853,N_16468,N_16283);
or U16854 (N_16854,N_16457,N_16142);
xor U16855 (N_16855,N_16168,N_16436);
nor U16856 (N_16856,N_16155,N_16460);
nor U16857 (N_16857,N_16466,N_16311);
nand U16858 (N_16858,N_16243,N_16393);
or U16859 (N_16859,N_16218,N_16062);
nor U16860 (N_16860,N_16272,N_16136);
xor U16861 (N_16861,N_16406,N_16067);
xor U16862 (N_16862,N_16225,N_16438);
and U16863 (N_16863,N_16365,N_16119);
nand U16864 (N_16864,N_16086,N_16405);
or U16865 (N_16865,N_16118,N_16102);
nor U16866 (N_16866,N_16062,N_16339);
nor U16867 (N_16867,N_16291,N_16198);
xor U16868 (N_16868,N_16274,N_16319);
xor U16869 (N_16869,N_16186,N_16096);
nand U16870 (N_16870,N_16030,N_16033);
nor U16871 (N_16871,N_16219,N_16192);
or U16872 (N_16872,N_16066,N_16430);
and U16873 (N_16873,N_16164,N_16318);
or U16874 (N_16874,N_16264,N_16407);
xnor U16875 (N_16875,N_16012,N_16219);
or U16876 (N_16876,N_16486,N_16037);
xor U16877 (N_16877,N_16355,N_16335);
and U16878 (N_16878,N_16061,N_16164);
nand U16879 (N_16879,N_16320,N_16280);
xnor U16880 (N_16880,N_16127,N_16042);
nand U16881 (N_16881,N_16337,N_16340);
nor U16882 (N_16882,N_16374,N_16132);
nor U16883 (N_16883,N_16444,N_16334);
or U16884 (N_16884,N_16031,N_16401);
nand U16885 (N_16885,N_16124,N_16185);
or U16886 (N_16886,N_16384,N_16185);
nand U16887 (N_16887,N_16397,N_16031);
or U16888 (N_16888,N_16288,N_16323);
xor U16889 (N_16889,N_16467,N_16083);
or U16890 (N_16890,N_16035,N_16175);
xnor U16891 (N_16891,N_16324,N_16367);
and U16892 (N_16892,N_16261,N_16487);
nand U16893 (N_16893,N_16205,N_16294);
nor U16894 (N_16894,N_16130,N_16480);
and U16895 (N_16895,N_16408,N_16193);
or U16896 (N_16896,N_16192,N_16282);
and U16897 (N_16897,N_16124,N_16491);
nand U16898 (N_16898,N_16129,N_16371);
nor U16899 (N_16899,N_16204,N_16086);
and U16900 (N_16900,N_16371,N_16269);
nand U16901 (N_16901,N_16410,N_16105);
or U16902 (N_16902,N_16226,N_16286);
xor U16903 (N_16903,N_16359,N_16156);
and U16904 (N_16904,N_16129,N_16409);
xnor U16905 (N_16905,N_16187,N_16267);
or U16906 (N_16906,N_16277,N_16499);
nor U16907 (N_16907,N_16458,N_16237);
and U16908 (N_16908,N_16414,N_16145);
xnor U16909 (N_16909,N_16423,N_16393);
xor U16910 (N_16910,N_16250,N_16148);
or U16911 (N_16911,N_16308,N_16406);
nand U16912 (N_16912,N_16126,N_16119);
or U16913 (N_16913,N_16160,N_16025);
and U16914 (N_16914,N_16181,N_16161);
nand U16915 (N_16915,N_16305,N_16226);
nand U16916 (N_16916,N_16326,N_16199);
xor U16917 (N_16917,N_16228,N_16032);
or U16918 (N_16918,N_16098,N_16384);
or U16919 (N_16919,N_16366,N_16310);
xor U16920 (N_16920,N_16098,N_16379);
nand U16921 (N_16921,N_16343,N_16437);
and U16922 (N_16922,N_16131,N_16061);
nor U16923 (N_16923,N_16176,N_16084);
or U16924 (N_16924,N_16106,N_16469);
xor U16925 (N_16925,N_16494,N_16140);
or U16926 (N_16926,N_16120,N_16278);
nand U16927 (N_16927,N_16000,N_16151);
and U16928 (N_16928,N_16314,N_16315);
nor U16929 (N_16929,N_16399,N_16184);
xor U16930 (N_16930,N_16122,N_16396);
nor U16931 (N_16931,N_16390,N_16069);
nor U16932 (N_16932,N_16126,N_16051);
nor U16933 (N_16933,N_16074,N_16048);
and U16934 (N_16934,N_16232,N_16426);
nor U16935 (N_16935,N_16017,N_16223);
xnor U16936 (N_16936,N_16097,N_16046);
and U16937 (N_16937,N_16303,N_16424);
and U16938 (N_16938,N_16247,N_16314);
xnor U16939 (N_16939,N_16473,N_16415);
or U16940 (N_16940,N_16134,N_16458);
nand U16941 (N_16941,N_16399,N_16435);
and U16942 (N_16942,N_16237,N_16126);
nor U16943 (N_16943,N_16316,N_16195);
nand U16944 (N_16944,N_16124,N_16430);
xor U16945 (N_16945,N_16453,N_16175);
and U16946 (N_16946,N_16065,N_16284);
nor U16947 (N_16947,N_16041,N_16357);
nand U16948 (N_16948,N_16426,N_16209);
nor U16949 (N_16949,N_16396,N_16139);
nand U16950 (N_16950,N_16443,N_16416);
xor U16951 (N_16951,N_16188,N_16167);
or U16952 (N_16952,N_16398,N_16025);
xor U16953 (N_16953,N_16227,N_16170);
xnor U16954 (N_16954,N_16373,N_16108);
and U16955 (N_16955,N_16213,N_16299);
or U16956 (N_16956,N_16093,N_16477);
and U16957 (N_16957,N_16227,N_16267);
and U16958 (N_16958,N_16095,N_16186);
nand U16959 (N_16959,N_16379,N_16200);
nand U16960 (N_16960,N_16158,N_16372);
nor U16961 (N_16961,N_16061,N_16476);
xnor U16962 (N_16962,N_16010,N_16281);
nor U16963 (N_16963,N_16460,N_16429);
nor U16964 (N_16964,N_16488,N_16170);
nor U16965 (N_16965,N_16118,N_16252);
nor U16966 (N_16966,N_16035,N_16146);
nand U16967 (N_16967,N_16452,N_16078);
or U16968 (N_16968,N_16022,N_16025);
xnor U16969 (N_16969,N_16032,N_16176);
nor U16970 (N_16970,N_16474,N_16112);
xor U16971 (N_16971,N_16361,N_16043);
nor U16972 (N_16972,N_16258,N_16438);
xnor U16973 (N_16973,N_16150,N_16311);
xor U16974 (N_16974,N_16270,N_16326);
or U16975 (N_16975,N_16175,N_16288);
and U16976 (N_16976,N_16197,N_16401);
and U16977 (N_16977,N_16039,N_16052);
and U16978 (N_16978,N_16484,N_16437);
nand U16979 (N_16979,N_16301,N_16023);
nor U16980 (N_16980,N_16409,N_16205);
nor U16981 (N_16981,N_16448,N_16038);
xnor U16982 (N_16982,N_16309,N_16318);
nor U16983 (N_16983,N_16491,N_16302);
nor U16984 (N_16984,N_16274,N_16125);
xnor U16985 (N_16985,N_16136,N_16295);
nand U16986 (N_16986,N_16258,N_16356);
nand U16987 (N_16987,N_16116,N_16163);
or U16988 (N_16988,N_16411,N_16492);
nand U16989 (N_16989,N_16160,N_16074);
and U16990 (N_16990,N_16323,N_16172);
xor U16991 (N_16991,N_16388,N_16344);
nand U16992 (N_16992,N_16370,N_16146);
nand U16993 (N_16993,N_16369,N_16174);
and U16994 (N_16994,N_16308,N_16132);
and U16995 (N_16995,N_16245,N_16100);
nand U16996 (N_16996,N_16238,N_16207);
nor U16997 (N_16997,N_16260,N_16098);
and U16998 (N_16998,N_16491,N_16449);
or U16999 (N_16999,N_16132,N_16155);
or U17000 (N_17000,N_16698,N_16781);
xor U17001 (N_17001,N_16909,N_16949);
nor U17002 (N_17002,N_16750,N_16992);
and U17003 (N_17003,N_16879,N_16617);
nor U17004 (N_17004,N_16504,N_16688);
nand U17005 (N_17005,N_16711,N_16842);
nor U17006 (N_17006,N_16985,N_16720);
nand U17007 (N_17007,N_16527,N_16924);
or U17008 (N_17008,N_16989,N_16564);
xor U17009 (N_17009,N_16818,N_16956);
or U17010 (N_17010,N_16948,N_16636);
xor U17011 (N_17011,N_16647,N_16746);
xor U17012 (N_17012,N_16601,N_16667);
xor U17013 (N_17013,N_16893,N_16975);
or U17014 (N_17014,N_16969,N_16925);
nand U17015 (N_17015,N_16904,N_16990);
and U17016 (N_17016,N_16680,N_16537);
and U17017 (N_17017,N_16870,N_16913);
nor U17018 (N_17018,N_16703,N_16999);
or U17019 (N_17019,N_16863,N_16886);
nor U17020 (N_17020,N_16816,N_16559);
nand U17021 (N_17021,N_16613,N_16916);
and U17022 (N_17022,N_16691,N_16858);
xor U17023 (N_17023,N_16779,N_16815);
nor U17024 (N_17024,N_16534,N_16809);
and U17025 (N_17025,N_16629,N_16812);
nor U17026 (N_17026,N_16915,N_16853);
nand U17027 (N_17027,N_16709,N_16821);
xor U17028 (N_17028,N_16957,N_16681);
xnor U17029 (N_17029,N_16503,N_16529);
xnor U17030 (N_17030,N_16888,N_16766);
nor U17031 (N_17031,N_16825,N_16973);
nand U17032 (N_17032,N_16618,N_16943);
and U17033 (N_17033,N_16862,N_16906);
nor U17034 (N_17034,N_16683,N_16631);
xnor U17035 (N_17035,N_16979,N_16525);
nor U17036 (N_17036,N_16612,N_16951);
and U17037 (N_17037,N_16621,N_16744);
and U17038 (N_17038,N_16823,N_16546);
nand U17039 (N_17039,N_16582,N_16715);
and U17040 (N_17040,N_16988,N_16843);
nand U17041 (N_17041,N_16895,N_16742);
nor U17042 (N_17042,N_16847,N_16995);
and U17043 (N_17043,N_16811,N_16541);
nor U17044 (N_17044,N_16731,N_16649);
or U17045 (N_17045,N_16581,N_16996);
xnor U17046 (N_17046,N_16512,N_16623);
nand U17047 (N_17047,N_16814,N_16937);
and U17048 (N_17048,N_16826,N_16550);
or U17049 (N_17049,N_16539,N_16577);
nor U17050 (N_17050,N_16699,N_16603);
or U17051 (N_17051,N_16628,N_16807);
xnor U17052 (N_17052,N_16508,N_16579);
nor U17053 (N_17053,N_16762,N_16782);
nand U17054 (N_17054,N_16902,N_16876);
or U17055 (N_17055,N_16773,N_16976);
nor U17056 (N_17056,N_16686,N_16810);
and U17057 (N_17057,N_16509,N_16675);
xor U17058 (N_17058,N_16903,N_16569);
or U17059 (N_17059,N_16729,N_16808);
xnor U17060 (N_17060,N_16935,N_16993);
and U17061 (N_17061,N_16650,N_16638);
nand U17062 (N_17062,N_16608,N_16566);
nor U17063 (N_17063,N_16834,N_16748);
nand U17064 (N_17064,N_16502,N_16947);
or U17065 (N_17065,N_16590,N_16955);
nor U17066 (N_17066,N_16760,N_16963);
or U17067 (N_17067,N_16830,N_16604);
nor U17068 (N_17068,N_16706,N_16668);
and U17069 (N_17069,N_16751,N_16580);
nand U17070 (N_17070,N_16648,N_16684);
or U17071 (N_17071,N_16934,N_16936);
or U17072 (N_17072,N_16733,N_16802);
xnor U17073 (N_17073,N_16739,N_16994);
nand U17074 (N_17074,N_16987,N_16515);
nor U17075 (N_17075,N_16970,N_16548);
nand U17076 (N_17076,N_16828,N_16849);
nor U17077 (N_17077,N_16789,N_16929);
and U17078 (N_17078,N_16506,N_16726);
and U17079 (N_17079,N_16772,N_16953);
xnor U17080 (N_17080,N_16869,N_16797);
nand U17081 (N_17081,N_16908,N_16767);
or U17082 (N_17082,N_16846,N_16761);
and U17083 (N_17083,N_16792,N_16778);
and U17084 (N_17084,N_16714,N_16555);
nor U17085 (N_17085,N_16661,N_16697);
xnor U17086 (N_17086,N_16759,N_16605);
nand U17087 (N_17087,N_16927,N_16907);
nand U17088 (N_17088,N_16662,N_16875);
xor U17089 (N_17089,N_16672,N_16620);
nor U17090 (N_17090,N_16511,N_16551);
nor U17091 (N_17091,N_16896,N_16984);
xnor U17092 (N_17092,N_16864,N_16597);
nand U17093 (N_17093,N_16928,N_16513);
and U17094 (N_17094,N_16837,N_16839);
xnor U17095 (N_17095,N_16754,N_16911);
or U17096 (N_17096,N_16942,N_16645);
or U17097 (N_17097,N_16570,N_16793);
or U17098 (N_17098,N_16941,N_16632);
xor U17099 (N_17099,N_16777,N_16595);
nor U17100 (N_17100,N_16769,N_16840);
xor U17101 (N_17101,N_16594,N_16881);
xnor U17102 (N_17102,N_16930,N_16644);
or U17103 (N_17103,N_16642,N_16861);
xor U17104 (N_17104,N_16655,N_16866);
nand U17105 (N_17105,N_16798,N_16982);
nor U17106 (N_17106,N_16931,N_16889);
nor U17107 (N_17107,N_16678,N_16961);
and U17108 (N_17108,N_16855,N_16557);
or U17109 (N_17109,N_16874,N_16673);
xnor U17110 (N_17110,N_16517,N_16532);
and U17111 (N_17111,N_16630,N_16890);
or U17112 (N_17112,N_16817,N_16521);
or U17113 (N_17113,N_16721,N_16967);
xor U17114 (N_17114,N_16757,N_16901);
nand U17115 (N_17115,N_16801,N_16880);
nor U17116 (N_17116,N_16624,N_16724);
and U17117 (N_17117,N_16905,N_16845);
and U17118 (N_17118,N_16554,N_16659);
or U17119 (N_17119,N_16526,N_16685);
xor U17120 (N_17120,N_16938,N_16510);
and U17121 (N_17121,N_16894,N_16519);
xnor U17122 (N_17122,N_16696,N_16585);
nor U17123 (N_17123,N_16983,N_16552);
xor U17124 (N_17124,N_16633,N_16922);
or U17125 (N_17125,N_16799,N_16516);
xor U17126 (N_17126,N_16713,N_16653);
nand U17127 (N_17127,N_16707,N_16600);
and U17128 (N_17128,N_16669,N_16584);
nand U17129 (N_17129,N_16820,N_16932);
nand U17130 (N_17130,N_16587,N_16663);
xnor U17131 (N_17131,N_16591,N_16528);
or U17132 (N_17132,N_16567,N_16921);
xnor U17133 (N_17133,N_16806,N_16614);
xnor U17134 (N_17134,N_16553,N_16791);
or U17135 (N_17135,N_16944,N_16701);
and U17136 (N_17136,N_16568,N_16523);
xnor U17137 (N_17137,N_16609,N_16736);
nor U17138 (N_17138,N_16920,N_16883);
xnor U17139 (N_17139,N_16966,N_16573);
nor U17140 (N_17140,N_16664,N_16787);
nand U17141 (N_17141,N_16737,N_16844);
nand U17142 (N_17142,N_16968,N_16933);
xnor U17143 (N_17143,N_16674,N_16705);
and U17144 (N_17144,N_16602,N_16514);
nand U17145 (N_17145,N_16563,N_16615);
or U17146 (N_17146,N_16940,N_16851);
nor U17147 (N_17147,N_16606,N_16877);
nand U17148 (N_17148,N_16848,N_16852);
nor U17149 (N_17149,N_16946,N_16693);
xor U17150 (N_17150,N_16538,N_16639);
nand U17151 (N_17151,N_16919,N_16575);
nor U17152 (N_17152,N_16670,N_16803);
or U17153 (N_17153,N_16657,N_16872);
nand U17154 (N_17154,N_16898,N_16959);
nand U17155 (N_17155,N_16592,N_16939);
xnor U17156 (N_17156,N_16780,N_16687);
nor U17157 (N_17157,N_16900,N_16794);
nand U17158 (N_17158,N_16796,N_16868);
and U17159 (N_17159,N_16640,N_16813);
nand U17160 (N_17160,N_16710,N_16980);
nor U17161 (N_17161,N_16704,N_16531);
and U17162 (N_17162,N_16634,N_16700);
nand U17163 (N_17163,N_16676,N_16571);
and U17164 (N_17164,N_16954,N_16841);
or U17165 (N_17165,N_16835,N_16611);
nor U17166 (N_17166,N_16785,N_16836);
nand U17167 (N_17167,N_16923,N_16882);
nor U17168 (N_17168,N_16771,N_16583);
xnor U17169 (N_17169,N_16740,N_16960);
xnor U17170 (N_17170,N_16912,N_16505);
or U17171 (N_17171,N_16690,N_16758);
and U17172 (N_17172,N_16914,N_16660);
nand U17173 (N_17173,N_16658,N_16520);
nand U17174 (N_17174,N_16540,N_16501);
and U17175 (N_17175,N_16530,N_16945);
or U17176 (N_17176,N_16745,N_16694);
nor U17177 (N_17177,N_16965,N_16977);
xnor U17178 (N_17178,N_16734,N_16986);
xor U17179 (N_17179,N_16997,N_16518);
nand U17180 (N_17180,N_16776,N_16565);
or U17181 (N_17181,N_16593,N_16790);
and U17182 (N_17182,N_16784,N_16626);
nor U17183 (N_17183,N_16832,N_16749);
or U17184 (N_17184,N_16543,N_16770);
or U17185 (N_17185,N_16646,N_16556);
or U17186 (N_17186,N_16610,N_16562);
xor U17187 (N_17187,N_16524,N_16910);
xor U17188 (N_17188,N_16533,N_16926);
or U17189 (N_17189,N_16522,N_16560);
nor U17190 (N_17190,N_16755,N_16651);
xor U17191 (N_17191,N_16666,N_16718);
xor U17192 (N_17192,N_16692,N_16884);
or U17193 (N_17193,N_16574,N_16682);
nor U17194 (N_17194,N_16730,N_16800);
xnor U17195 (N_17195,N_16544,N_16865);
nand U17196 (N_17196,N_16578,N_16616);
or U17197 (N_17197,N_16738,N_16671);
nand U17198 (N_17198,N_16827,N_16747);
nand U17199 (N_17199,N_16854,N_16804);
nor U17200 (N_17200,N_16743,N_16978);
nand U17201 (N_17201,N_16607,N_16829);
or U17202 (N_17202,N_16656,N_16561);
nor U17203 (N_17203,N_16765,N_16637);
xnor U17204 (N_17204,N_16735,N_16856);
xnor U17205 (N_17205,N_16981,N_16897);
nand U17206 (N_17206,N_16619,N_16665);
nor U17207 (N_17207,N_16598,N_16622);
nor U17208 (N_17208,N_16971,N_16857);
nand U17209 (N_17209,N_16599,N_16652);
xnor U17210 (N_17210,N_16958,N_16962);
nor U17211 (N_17211,N_16887,N_16867);
and U17212 (N_17212,N_16991,N_16822);
nor U17213 (N_17213,N_16586,N_16643);
and U17214 (N_17214,N_16795,N_16819);
and U17215 (N_17215,N_16917,N_16741);
xnor U17216 (N_17216,N_16732,N_16918);
nand U17217 (N_17217,N_16859,N_16891);
nand U17218 (N_17218,N_16878,N_16727);
and U17219 (N_17219,N_16952,N_16572);
nor U17220 (N_17220,N_16871,N_16625);
xnor U17221 (N_17221,N_16850,N_16974);
xor U17222 (N_17222,N_16764,N_16775);
xor U17223 (N_17223,N_16717,N_16833);
or U17224 (N_17224,N_16860,N_16627);
xor U17225 (N_17225,N_16535,N_16725);
nand U17226 (N_17226,N_16824,N_16596);
nor U17227 (N_17227,N_16753,N_16752);
or U17228 (N_17228,N_16549,N_16722);
xor U17229 (N_17229,N_16679,N_16702);
or U17230 (N_17230,N_16899,N_16589);
nor U17231 (N_17231,N_16774,N_16788);
xnor U17232 (N_17232,N_16805,N_16695);
and U17233 (N_17233,N_16723,N_16545);
nor U17234 (N_17234,N_16500,N_16558);
xnor U17235 (N_17235,N_16950,N_16712);
and U17236 (N_17236,N_16972,N_16654);
nor U17237 (N_17237,N_16542,N_16838);
xnor U17238 (N_17238,N_16635,N_16576);
xor U17239 (N_17239,N_16885,N_16786);
nand U17240 (N_17240,N_16728,N_16719);
xor U17241 (N_17241,N_16641,N_16873);
and U17242 (N_17242,N_16677,N_16507);
nor U17243 (N_17243,N_16768,N_16689);
or U17244 (N_17244,N_16783,N_16892);
xor U17245 (N_17245,N_16536,N_16547);
or U17246 (N_17246,N_16708,N_16998);
and U17247 (N_17247,N_16831,N_16588);
xor U17248 (N_17248,N_16964,N_16716);
xnor U17249 (N_17249,N_16763,N_16756);
and U17250 (N_17250,N_16875,N_16519);
and U17251 (N_17251,N_16586,N_16746);
and U17252 (N_17252,N_16920,N_16859);
or U17253 (N_17253,N_16744,N_16955);
and U17254 (N_17254,N_16586,N_16773);
or U17255 (N_17255,N_16913,N_16951);
or U17256 (N_17256,N_16729,N_16989);
nor U17257 (N_17257,N_16849,N_16715);
xnor U17258 (N_17258,N_16919,N_16847);
nand U17259 (N_17259,N_16811,N_16787);
and U17260 (N_17260,N_16851,N_16935);
nor U17261 (N_17261,N_16544,N_16711);
nand U17262 (N_17262,N_16721,N_16815);
or U17263 (N_17263,N_16820,N_16949);
nand U17264 (N_17264,N_16662,N_16755);
xor U17265 (N_17265,N_16535,N_16919);
or U17266 (N_17266,N_16873,N_16972);
or U17267 (N_17267,N_16597,N_16801);
or U17268 (N_17268,N_16675,N_16577);
nand U17269 (N_17269,N_16617,N_16895);
and U17270 (N_17270,N_16908,N_16762);
nand U17271 (N_17271,N_16806,N_16668);
and U17272 (N_17272,N_16918,N_16815);
xnor U17273 (N_17273,N_16691,N_16599);
nor U17274 (N_17274,N_16601,N_16761);
xor U17275 (N_17275,N_16610,N_16992);
nand U17276 (N_17276,N_16866,N_16972);
nor U17277 (N_17277,N_16710,N_16896);
or U17278 (N_17278,N_16849,N_16854);
and U17279 (N_17279,N_16637,N_16676);
nand U17280 (N_17280,N_16912,N_16822);
or U17281 (N_17281,N_16578,N_16951);
nor U17282 (N_17282,N_16661,N_16863);
and U17283 (N_17283,N_16848,N_16807);
or U17284 (N_17284,N_16748,N_16969);
nor U17285 (N_17285,N_16562,N_16833);
or U17286 (N_17286,N_16912,N_16762);
and U17287 (N_17287,N_16907,N_16669);
or U17288 (N_17288,N_16720,N_16996);
nand U17289 (N_17289,N_16586,N_16567);
nand U17290 (N_17290,N_16711,N_16875);
or U17291 (N_17291,N_16923,N_16799);
xnor U17292 (N_17292,N_16975,N_16656);
and U17293 (N_17293,N_16976,N_16616);
and U17294 (N_17294,N_16849,N_16935);
nor U17295 (N_17295,N_16641,N_16856);
nor U17296 (N_17296,N_16634,N_16571);
or U17297 (N_17297,N_16549,N_16627);
nor U17298 (N_17298,N_16702,N_16532);
nand U17299 (N_17299,N_16627,N_16562);
xor U17300 (N_17300,N_16563,N_16829);
xor U17301 (N_17301,N_16995,N_16693);
nand U17302 (N_17302,N_16996,N_16675);
nor U17303 (N_17303,N_16860,N_16787);
and U17304 (N_17304,N_16570,N_16982);
or U17305 (N_17305,N_16851,N_16915);
or U17306 (N_17306,N_16988,N_16856);
or U17307 (N_17307,N_16994,N_16842);
xor U17308 (N_17308,N_16964,N_16505);
and U17309 (N_17309,N_16991,N_16764);
or U17310 (N_17310,N_16548,N_16973);
or U17311 (N_17311,N_16682,N_16634);
and U17312 (N_17312,N_16802,N_16794);
nand U17313 (N_17313,N_16562,N_16944);
nand U17314 (N_17314,N_16768,N_16541);
nor U17315 (N_17315,N_16501,N_16762);
or U17316 (N_17316,N_16508,N_16689);
nor U17317 (N_17317,N_16594,N_16554);
nor U17318 (N_17318,N_16858,N_16681);
xnor U17319 (N_17319,N_16985,N_16652);
or U17320 (N_17320,N_16827,N_16562);
and U17321 (N_17321,N_16866,N_16555);
nand U17322 (N_17322,N_16849,N_16868);
nand U17323 (N_17323,N_16957,N_16952);
xnor U17324 (N_17324,N_16686,N_16681);
and U17325 (N_17325,N_16701,N_16823);
xnor U17326 (N_17326,N_16740,N_16803);
nand U17327 (N_17327,N_16694,N_16827);
nand U17328 (N_17328,N_16503,N_16554);
xor U17329 (N_17329,N_16502,N_16825);
nand U17330 (N_17330,N_16739,N_16552);
and U17331 (N_17331,N_16599,N_16573);
and U17332 (N_17332,N_16608,N_16734);
nor U17333 (N_17333,N_16586,N_16908);
xor U17334 (N_17334,N_16590,N_16632);
or U17335 (N_17335,N_16894,N_16935);
and U17336 (N_17336,N_16847,N_16599);
xnor U17337 (N_17337,N_16993,N_16924);
xor U17338 (N_17338,N_16919,N_16537);
nand U17339 (N_17339,N_16668,N_16968);
and U17340 (N_17340,N_16692,N_16829);
or U17341 (N_17341,N_16539,N_16819);
and U17342 (N_17342,N_16997,N_16510);
and U17343 (N_17343,N_16567,N_16555);
nor U17344 (N_17344,N_16763,N_16818);
and U17345 (N_17345,N_16560,N_16825);
xnor U17346 (N_17346,N_16852,N_16821);
nand U17347 (N_17347,N_16915,N_16685);
or U17348 (N_17348,N_16807,N_16818);
xor U17349 (N_17349,N_16511,N_16743);
nand U17350 (N_17350,N_16995,N_16938);
xor U17351 (N_17351,N_16553,N_16720);
or U17352 (N_17352,N_16912,N_16986);
nand U17353 (N_17353,N_16696,N_16982);
xor U17354 (N_17354,N_16862,N_16987);
or U17355 (N_17355,N_16785,N_16879);
xor U17356 (N_17356,N_16639,N_16896);
nor U17357 (N_17357,N_16684,N_16959);
nor U17358 (N_17358,N_16600,N_16922);
xor U17359 (N_17359,N_16732,N_16879);
and U17360 (N_17360,N_16540,N_16774);
nor U17361 (N_17361,N_16683,N_16606);
nand U17362 (N_17362,N_16624,N_16778);
nor U17363 (N_17363,N_16593,N_16777);
or U17364 (N_17364,N_16919,N_16678);
nand U17365 (N_17365,N_16716,N_16689);
nand U17366 (N_17366,N_16862,N_16746);
or U17367 (N_17367,N_16646,N_16633);
nor U17368 (N_17368,N_16501,N_16802);
xor U17369 (N_17369,N_16610,N_16809);
or U17370 (N_17370,N_16710,N_16526);
nand U17371 (N_17371,N_16760,N_16872);
and U17372 (N_17372,N_16946,N_16917);
and U17373 (N_17373,N_16800,N_16892);
xnor U17374 (N_17374,N_16553,N_16892);
nand U17375 (N_17375,N_16818,N_16551);
xor U17376 (N_17376,N_16880,N_16940);
xor U17377 (N_17377,N_16998,N_16746);
nor U17378 (N_17378,N_16897,N_16895);
and U17379 (N_17379,N_16551,N_16592);
nand U17380 (N_17380,N_16793,N_16856);
or U17381 (N_17381,N_16742,N_16520);
nand U17382 (N_17382,N_16955,N_16664);
and U17383 (N_17383,N_16580,N_16786);
nor U17384 (N_17384,N_16792,N_16815);
and U17385 (N_17385,N_16947,N_16537);
xor U17386 (N_17386,N_16646,N_16532);
nand U17387 (N_17387,N_16866,N_16837);
xnor U17388 (N_17388,N_16715,N_16781);
and U17389 (N_17389,N_16857,N_16555);
nor U17390 (N_17390,N_16525,N_16640);
or U17391 (N_17391,N_16958,N_16945);
nor U17392 (N_17392,N_16610,N_16503);
or U17393 (N_17393,N_16512,N_16956);
and U17394 (N_17394,N_16962,N_16879);
nand U17395 (N_17395,N_16758,N_16748);
or U17396 (N_17396,N_16660,N_16833);
nor U17397 (N_17397,N_16982,N_16604);
nand U17398 (N_17398,N_16852,N_16912);
nor U17399 (N_17399,N_16998,N_16658);
nand U17400 (N_17400,N_16787,N_16573);
nor U17401 (N_17401,N_16579,N_16683);
and U17402 (N_17402,N_16916,N_16725);
or U17403 (N_17403,N_16644,N_16822);
xor U17404 (N_17404,N_16515,N_16927);
xor U17405 (N_17405,N_16934,N_16967);
or U17406 (N_17406,N_16671,N_16934);
nor U17407 (N_17407,N_16815,N_16505);
xor U17408 (N_17408,N_16881,N_16529);
xnor U17409 (N_17409,N_16781,N_16878);
nand U17410 (N_17410,N_16639,N_16913);
or U17411 (N_17411,N_16818,N_16557);
xor U17412 (N_17412,N_16557,N_16985);
or U17413 (N_17413,N_16776,N_16846);
nand U17414 (N_17414,N_16954,N_16867);
and U17415 (N_17415,N_16569,N_16587);
xnor U17416 (N_17416,N_16926,N_16874);
nand U17417 (N_17417,N_16519,N_16957);
nand U17418 (N_17418,N_16700,N_16583);
xnor U17419 (N_17419,N_16866,N_16971);
nand U17420 (N_17420,N_16754,N_16728);
or U17421 (N_17421,N_16994,N_16619);
nand U17422 (N_17422,N_16501,N_16615);
and U17423 (N_17423,N_16513,N_16749);
nand U17424 (N_17424,N_16834,N_16799);
nor U17425 (N_17425,N_16607,N_16866);
xor U17426 (N_17426,N_16724,N_16973);
or U17427 (N_17427,N_16987,N_16840);
nand U17428 (N_17428,N_16927,N_16577);
or U17429 (N_17429,N_16862,N_16930);
and U17430 (N_17430,N_16817,N_16853);
nand U17431 (N_17431,N_16732,N_16768);
or U17432 (N_17432,N_16613,N_16766);
or U17433 (N_17433,N_16781,N_16947);
or U17434 (N_17434,N_16996,N_16990);
and U17435 (N_17435,N_16862,N_16712);
nor U17436 (N_17436,N_16796,N_16506);
or U17437 (N_17437,N_16554,N_16994);
and U17438 (N_17438,N_16572,N_16806);
xnor U17439 (N_17439,N_16556,N_16747);
nand U17440 (N_17440,N_16728,N_16911);
nor U17441 (N_17441,N_16934,N_16756);
nor U17442 (N_17442,N_16573,N_16985);
nor U17443 (N_17443,N_16888,N_16791);
xnor U17444 (N_17444,N_16551,N_16949);
nor U17445 (N_17445,N_16648,N_16755);
xor U17446 (N_17446,N_16635,N_16730);
nand U17447 (N_17447,N_16818,N_16553);
xnor U17448 (N_17448,N_16686,N_16583);
xor U17449 (N_17449,N_16603,N_16722);
or U17450 (N_17450,N_16562,N_16619);
nand U17451 (N_17451,N_16765,N_16904);
nand U17452 (N_17452,N_16974,N_16838);
and U17453 (N_17453,N_16702,N_16947);
or U17454 (N_17454,N_16917,N_16759);
or U17455 (N_17455,N_16853,N_16923);
xnor U17456 (N_17456,N_16972,N_16963);
or U17457 (N_17457,N_16903,N_16966);
nor U17458 (N_17458,N_16928,N_16622);
and U17459 (N_17459,N_16559,N_16656);
xor U17460 (N_17460,N_16690,N_16634);
nor U17461 (N_17461,N_16699,N_16630);
nor U17462 (N_17462,N_16528,N_16665);
or U17463 (N_17463,N_16553,N_16718);
xor U17464 (N_17464,N_16982,N_16565);
xnor U17465 (N_17465,N_16645,N_16844);
and U17466 (N_17466,N_16603,N_16901);
xnor U17467 (N_17467,N_16735,N_16850);
xor U17468 (N_17468,N_16674,N_16514);
xnor U17469 (N_17469,N_16809,N_16664);
and U17470 (N_17470,N_16519,N_16776);
xor U17471 (N_17471,N_16949,N_16936);
and U17472 (N_17472,N_16737,N_16722);
nor U17473 (N_17473,N_16563,N_16964);
or U17474 (N_17474,N_16731,N_16536);
nor U17475 (N_17475,N_16663,N_16712);
nand U17476 (N_17476,N_16673,N_16804);
nand U17477 (N_17477,N_16788,N_16670);
and U17478 (N_17478,N_16538,N_16998);
xor U17479 (N_17479,N_16646,N_16685);
xnor U17480 (N_17480,N_16555,N_16950);
or U17481 (N_17481,N_16795,N_16791);
nor U17482 (N_17482,N_16860,N_16917);
and U17483 (N_17483,N_16578,N_16932);
or U17484 (N_17484,N_16884,N_16900);
and U17485 (N_17485,N_16633,N_16736);
xnor U17486 (N_17486,N_16667,N_16869);
and U17487 (N_17487,N_16638,N_16525);
xnor U17488 (N_17488,N_16528,N_16547);
and U17489 (N_17489,N_16521,N_16678);
and U17490 (N_17490,N_16983,N_16686);
and U17491 (N_17491,N_16763,N_16929);
and U17492 (N_17492,N_16885,N_16702);
or U17493 (N_17493,N_16720,N_16637);
xnor U17494 (N_17494,N_16793,N_16749);
and U17495 (N_17495,N_16969,N_16573);
or U17496 (N_17496,N_16994,N_16526);
and U17497 (N_17497,N_16706,N_16874);
xnor U17498 (N_17498,N_16810,N_16644);
nand U17499 (N_17499,N_16896,N_16954);
and U17500 (N_17500,N_17218,N_17240);
and U17501 (N_17501,N_17290,N_17353);
nor U17502 (N_17502,N_17485,N_17411);
xor U17503 (N_17503,N_17378,N_17320);
and U17504 (N_17504,N_17158,N_17117);
nor U17505 (N_17505,N_17054,N_17136);
xnor U17506 (N_17506,N_17396,N_17326);
nand U17507 (N_17507,N_17060,N_17357);
and U17508 (N_17508,N_17424,N_17224);
or U17509 (N_17509,N_17147,N_17022);
nor U17510 (N_17510,N_17385,N_17341);
xor U17511 (N_17511,N_17072,N_17305);
xnor U17512 (N_17512,N_17495,N_17186);
nand U17513 (N_17513,N_17171,N_17464);
nand U17514 (N_17514,N_17467,N_17456);
nor U17515 (N_17515,N_17225,N_17263);
nor U17516 (N_17516,N_17313,N_17484);
nand U17517 (N_17517,N_17355,N_17428);
xnor U17518 (N_17518,N_17232,N_17333);
or U17519 (N_17519,N_17414,N_17001);
or U17520 (N_17520,N_17322,N_17262);
nor U17521 (N_17521,N_17102,N_17479);
nand U17522 (N_17522,N_17024,N_17159);
nand U17523 (N_17523,N_17079,N_17468);
or U17524 (N_17524,N_17365,N_17113);
nand U17525 (N_17525,N_17036,N_17403);
xor U17526 (N_17526,N_17366,N_17329);
nor U17527 (N_17527,N_17033,N_17324);
or U17528 (N_17528,N_17198,N_17166);
and U17529 (N_17529,N_17392,N_17384);
nand U17530 (N_17530,N_17111,N_17459);
nand U17531 (N_17531,N_17139,N_17144);
and U17532 (N_17532,N_17243,N_17478);
or U17533 (N_17533,N_17220,N_17150);
nand U17534 (N_17534,N_17071,N_17463);
nand U17535 (N_17535,N_17181,N_17372);
and U17536 (N_17536,N_17439,N_17156);
or U17537 (N_17537,N_17020,N_17006);
nor U17538 (N_17538,N_17344,N_17406);
xor U17539 (N_17539,N_17109,N_17330);
or U17540 (N_17540,N_17004,N_17000);
nand U17541 (N_17541,N_17394,N_17399);
or U17542 (N_17542,N_17048,N_17032);
nor U17543 (N_17543,N_17073,N_17053);
nand U17544 (N_17544,N_17300,N_17162);
xnor U17545 (N_17545,N_17078,N_17420);
or U17546 (N_17546,N_17319,N_17462);
nand U17547 (N_17547,N_17261,N_17301);
nor U17548 (N_17548,N_17165,N_17309);
nor U17549 (N_17549,N_17371,N_17405);
xnor U17550 (N_17550,N_17238,N_17276);
nand U17551 (N_17551,N_17303,N_17021);
nor U17552 (N_17552,N_17321,N_17223);
xnor U17553 (N_17553,N_17148,N_17254);
nor U17554 (N_17554,N_17059,N_17057);
nand U17555 (N_17555,N_17266,N_17027);
or U17556 (N_17556,N_17483,N_17297);
and U17557 (N_17557,N_17140,N_17310);
xor U17558 (N_17558,N_17245,N_17077);
xor U17559 (N_17559,N_17193,N_17412);
nand U17560 (N_17560,N_17489,N_17207);
or U17561 (N_17561,N_17012,N_17304);
and U17562 (N_17562,N_17028,N_17242);
nand U17563 (N_17563,N_17432,N_17358);
xor U17564 (N_17564,N_17143,N_17334);
or U17565 (N_17565,N_17093,N_17317);
and U17566 (N_17566,N_17041,N_17393);
or U17567 (N_17567,N_17130,N_17096);
or U17568 (N_17568,N_17375,N_17058);
xnor U17569 (N_17569,N_17445,N_17256);
or U17570 (N_17570,N_17349,N_17362);
or U17571 (N_17571,N_17444,N_17241);
xor U17572 (N_17572,N_17381,N_17338);
xor U17573 (N_17573,N_17308,N_17327);
nor U17574 (N_17574,N_17189,N_17034);
nor U17575 (N_17575,N_17473,N_17451);
xor U17576 (N_17576,N_17315,N_17236);
and U17577 (N_17577,N_17101,N_17257);
nor U17578 (N_17578,N_17114,N_17452);
nand U17579 (N_17579,N_17044,N_17348);
xnor U17580 (N_17580,N_17448,N_17170);
xor U17581 (N_17581,N_17360,N_17110);
nand U17582 (N_17582,N_17202,N_17342);
and U17583 (N_17583,N_17450,N_17088);
xnor U17584 (N_17584,N_17318,N_17107);
nand U17585 (N_17585,N_17328,N_17002);
xor U17586 (N_17586,N_17226,N_17345);
nor U17587 (N_17587,N_17269,N_17499);
xor U17588 (N_17588,N_17260,N_17486);
and U17589 (N_17589,N_17208,N_17354);
xnor U17590 (N_17590,N_17472,N_17426);
or U17591 (N_17591,N_17373,N_17227);
nand U17592 (N_17592,N_17183,N_17106);
or U17593 (N_17593,N_17296,N_17292);
xor U17594 (N_17594,N_17124,N_17359);
nand U17595 (N_17595,N_17434,N_17142);
or U17596 (N_17596,N_17010,N_17281);
or U17597 (N_17597,N_17474,N_17298);
xor U17598 (N_17598,N_17215,N_17285);
and U17599 (N_17599,N_17052,N_17350);
nand U17600 (N_17600,N_17383,N_17168);
nor U17601 (N_17601,N_17339,N_17201);
and U17602 (N_17602,N_17336,N_17274);
nor U17603 (N_17603,N_17476,N_17194);
nand U17604 (N_17604,N_17013,N_17419);
and U17605 (N_17605,N_17176,N_17233);
and U17606 (N_17606,N_17442,N_17237);
nand U17607 (N_17607,N_17294,N_17118);
xnor U17608 (N_17608,N_17047,N_17154);
nor U17609 (N_17609,N_17205,N_17031);
or U17610 (N_17610,N_17160,N_17417);
nor U17611 (N_17611,N_17137,N_17427);
xnor U17612 (N_17612,N_17061,N_17014);
or U17613 (N_17613,N_17248,N_17407);
or U17614 (N_17614,N_17086,N_17457);
nand U17615 (N_17615,N_17045,N_17216);
and U17616 (N_17616,N_17128,N_17374);
xnor U17617 (N_17617,N_17095,N_17075);
or U17618 (N_17618,N_17461,N_17090);
or U17619 (N_17619,N_17413,N_17410);
or U17620 (N_17620,N_17164,N_17370);
and U17621 (N_17621,N_17286,N_17066);
nand U17622 (N_17622,N_17219,N_17307);
and U17623 (N_17623,N_17367,N_17446);
nand U17624 (N_17624,N_17376,N_17173);
nor U17625 (N_17625,N_17222,N_17312);
nor U17626 (N_17626,N_17469,N_17449);
and U17627 (N_17627,N_17108,N_17440);
or U17628 (N_17628,N_17015,N_17038);
nand U17629 (N_17629,N_17480,N_17465);
nand U17630 (N_17630,N_17389,N_17284);
xnor U17631 (N_17631,N_17155,N_17259);
xnor U17632 (N_17632,N_17163,N_17258);
and U17633 (N_17633,N_17040,N_17100);
nor U17634 (N_17634,N_17351,N_17184);
nand U17635 (N_17635,N_17453,N_17404);
nand U17636 (N_17636,N_17084,N_17488);
nor U17637 (N_17637,N_17049,N_17221);
xnor U17638 (N_17638,N_17119,N_17007);
nor U17639 (N_17639,N_17239,N_17429);
or U17640 (N_17640,N_17092,N_17234);
nand U17641 (N_17641,N_17085,N_17134);
nand U17642 (N_17642,N_17120,N_17203);
or U17643 (N_17643,N_17364,N_17011);
and U17644 (N_17644,N_17125,N_17390);
nand U17645 (N_17645,N_17029,N_17246);
xnor U17646 (N_17646,N_17074,N_17408);
and U17647 (N_17647,N_17431,N_17065);
xor U17648 (N_17648,N_17493,N_17206);
or U17649 (N_17649,N_17423,N_17196);
nor U17650 (N_17650,N_17018,N_17430);
or U17651 (N_17651,N_17487,N_17089);
xor U17652 (N_17652,N_17352,N_17231);
and U17653 (N_17653,N_17454,N_17212);
nand U17654 (N_17654,N_17082,N_17282);
xnor U17655 (N_17655,N_17332,N_17083);
or U17656 (N_17656,N_17149,N_17008);
and U17657 (N_17657,N_17217,N_17293);
and U17658 (N_17658,N_17331,N_17172);
and U17659 (N_17659,N_17081,N_17200);
and U17660 (N_17660,N_17076,N_17035);
nand U17661 (N_17661,N_17116,N_17123);
or U17662 (N_17662,N_17187,N_17409);
nand U17663 (N_17663,N_17094,N_17311);
xnor U17664 (N_17664,N_17347,N_17497);
or U17665 (N_17665,N_17279,N_17380);
xnor U17666 (N_17666,N_17275,N_17152);
or U17667 (N_17667,N_17030,N_17127);
or U17668 (N_17668,N_17135,N_17017);
nand U17669 (N_17669,N_17270,N_17122);
nor U17670 (N_17670,N_17368,N_17306);
or U17671 (N_17671,N_17255,N_17167);
and U17672 (N_17672,N_17210,N_17115);
nor U17673 (N_17673,N_17447,N_17126);
or U17674 (N_17674,N_17314,N_17498);
nand U17675 (N_17675,N_17199,N_17067);
xor U17676 (N_17676,N_17046,N_17400);
and U17677 (N_17677,N_17415,N_17069);
or U17678 (N_17678,N_17195,N_17153);
nand U17679 (N_17679,N_17460,N_17490);
nor U17680 (N_17680,N_17250,N_17491);
nor U17681 (N_17681,N_17401,N_17063);
or U17682 (N_17682,N_17477,N_17174);
nand U17683 (N_17683,N_17441,N_17228);
nor U17684 (N_17684,N_17112,N_17235);
xor U17685 (N_17685,N_17051,N_17151);
or U17686 (N_17686,N_17131,N_17455);
and U17687 (N_17687,N_17191,N_17190);
or U17688 (N_17688,N_17443,N_17481);
xnor U17689 (N_17689,N_17070,N_17099);
and U17690 (N_17690,N_17356,N_17204);
nor U17691 (N_17691,N_17026,N_17388);
nor U17692 (N_17692,N_17299,N_17175);
nand U17693 (N_17693,N_17087,N_17050);
or U17694 (N_17694,N_17494,N_17105);
xnor U17695 (N_17695,N_17492,N_17252);
xor U17696 (N_17696,N_17161,N_17418);
nand U17697 (N_17697,N_17346,N_17230);
and U17698 (N_17698,N_17340,N_17277);
nor U17699 (N_17699,N_17379,N_17387);
or U17700 (N_17700,N_17271,N_17391);
or U17701 (N_17701,N_17253,N_17129);
nand U17702 (N_17702,N_17211,N_17138);
nand U17703 (N_17703,N_17482,N_17132);
or U17704 (N_17704,N_17104,N_17343);
xor U17705 (N_17705,N_17188,N_17386);
nand U17706 (N_17706,N_17361,N_17146);
nand U17707 (N_17707,N_17425,N_17283);
xnor U17708 (N_17708,N_17422,N_17062);
or U17709 (N_17709,N_17295,N_17398);
nand U17710 (N_17710,N_17005,N_17023);
and U17711 (N_17711,N_17169,N_17278);
xor U17712 (N_17712,N_17178,N_17251);
or U17713 (N_17713,N_17325,N_17302);
nor U17714 (N_17714,N_17080,N_17185);
nand U17715 (N_17715,N_17435,N_17265);
nor U17716 (N_17716,N_17141,N_17337);
or U17717 (N_17717,N_17369,N_17475);
nor U17718 (N_17718,N_17496,N_17402);
nand U17719 (N_17719,N_17397,N_17470);
nand U17720 (N_17720,N_17180,N_17064);
xor U17721 (N_17721,N_17229,N_17471);
and U17722 (N_17722,N_17009,N_17280);
and U17723 (N_17723,N_17316,N_17323);
or U17724 (N_17724,N_17433,N_17272);
nor U17725 (N_17725,N_17039,N_17043);
and U17726 (N_17726,N_17068,N_17133);
nor U17727 (N_17727,N_17416,N_17377);
xnor U17728 (N_17728,N_17264,N_17395);
xnor U17729 (N_17729,N_17363,N_17025);
xor U17730 (N_17730,N_17091,N_17056);
or U17731 (N_17731,N_17247,N_17288);
and U17732 (N_17732,N_17016,N_17438);
nand U17733 (N_17733,N_17157,N_17273);
or U17734 (N_17734,N_17003,N_17209);
xnor U17735 (N_17735,N_17098,N_17436);
xor U17736 (N_17736,N_17466,N_17268);
or U17737 (N_17737,N_17249,N_17213);
xor U17738 (N_17738,N_17289,N_17197);
nand U17739 (N_17739,N_17244,N_17019);
or U17740 (N_17740,N_17382,N_17182);
or U17741 (N_17741,N_17335,N_17421);
and U17742 (N_17742,N_17121,N_17179);
xor U17743 (N_17743,N_17287,N_17145);
nand U17744 (N_17744,N_17037,N_17103);
xor U17745 (N_17745,N_17192,N_17042);
and U17746 (N_17746,N_17177,N_17437);
xnor U17747 (N_17747,N_17291,N_17458);
nand U17748 (N_17748,N_17055,N_17097);
nand U17749 (N_17749,N_17267,N_17214);
xor U17750 (N_17750,N_17148,N_17231);
and U17751 (N_17751,N_17336,N_17272);
nor U17752 (N_17752,N_17470,N_17308);
nor U17753 (N_17753,N_17286,N_17259);
nor U17754 (N_17754,N_17170,N_17079);
nor U17755 (N_17755,N_17490,N_17313);
nor U17756 (N_17756,N_17347,N_17047);
xnor U17757 (N_17757,N_17138,N_17265);
and U17758 (N_17758,N_17498,N_17435);
nor U17759 (N_17759,N_17356,N_17445);
nor U17760 (N_17760,N_17056,N_17344);
and U17761 (N_17761,N_17424,N_17050);
nand U17762 (N_17762,N_17361,N_17330);
xor U17763 (N_17763,N_17131,N_17406);
and U17764 (N_17764,N_17160,N_17294);
and U17765 (N_17765,N_17383,N_17109);
and U17766 (N_17766,N_17020,N_17247);
nor U17767 (N_17767,N_17232,N_17473);
nor U17768 (N_17768,N_17359,N_17362);
and U17769 (N_17769,N_17302,N_17238);
or U17770 (N_17770,N_17083,N_17177);
or U17771 (N_17771,N_17061,N_17467);
nor U17772 (N_17772,N_17278,N_17394);
nand U17773 (N_17773,N_17387,N_17485);
xor U17774 (N_17774,N_17097,N_17224);
nor U17775 (N_17775,N_17406,N_17013);
nor U17776 (N_17776,N_17177,N_17297);
and U17777 (N_17777,N_17389,N_17084);
xor U17778 (N_17778,N_17413,N_17403);
nor U17779 (N_17779,N_17477,N_17084);
xnor U17780 (N_17780,N_17201,N_17378);
or U17781 (N_17781,N_17102,N_17265);
nand U17782 (N_17782,N_17202,N_17494);
nor U17783 (N_17783,N_17213,N_17425);
and U17784 (N_17784,N_17264,N_17281);
and U17785 (N_17785,N_17423,N_17286);
nor U17786 (N_17786,N_17165,N_17252);
nand U17787 (N_17787,N_17034,N_17241);
or U17788 (N_17788,N_17372,N_17295);
and U17789 (N_17789,N_17251,N_17041);
nand U17790 (N_17790,N_17432,N_17074);
and U17791 (N_17791,N_17411,N_17160);
or U17792 (N_17792,N_17025,N_17250);
and U17793 (N_17793,N_17182,N_17110);
or U17794 (N_17794,N_17466,N_17263);
nand U17795 (N_17795,N_17437,N_17296);
xnor U17796 (N_17796,N_17483,N_17466);
and U17797 (N_17797,N_17017,N_17083);
nor U17798 (N_17798,N_17315,N_17043);
xnor U17799 (N_17799,N_17250,N_17001);
or U17800 (N_17800,N_17257,N_17217);
nand U17801 (N_17801,N_17141,N_17460);
nor U17802 (N_17802,N_17279,N_17361);
or U17803 (N_17803,N_17373,N_17231);
xnor U17804 (N_17804,N_17314,N_17280);
nor U17805 (N_17805,N_17191,N_17285);
xnor U17806 (N_17806,N_17054,N_17375);
xnor U17807 (N_17807,N_17312,N_17223);
nor U17808 (N_17808,N_17109,N_17359);
nor U17809 (N_17809,N_17027,N_17157);
xnor U17810 (N_17810,N_17218,N_17471);
xnor U17811 (N_17811,N_17076,N_17353);
nor U17812 (N_17812,N_17173,N_17453);
and U17813 (N_17813,N_17320,N_17181);
and U17814 (N_17814,N_17434,N_17499);
xor U17815 (N_17815,N_17227,N_17322);
and U17816 (N_17816,N_17442,N_17151);
or U17817 (N_17817,N_17122,N_17496);
nor U17818 (N_17818,N_17172,N_17136);
nor U17819 (N_17819,N_17307,N_17109);
nor U17820 (N_17820,N_17239,N_17389);
or U17821 (N_17821,N_17063,N_17405);
nand U17822 (N_17822,N_17309,N_17315);
xor U17823 (N_17823,N_17147,N_17438);
xnor U17824 (N_17824,N_17471,N_17345);
and U17825 (N_17825,N_17092,N_17260);
and U17826 (N_17826,N_17334,N_17298);
or U17827 (N_17827,N_17445,N_17465);
nand U17828 (N_17828,N_17471,N_17284);
nor U17829 (N_17829,N_17212,N_17290);
or U17830 (N_17830,N_17307,N_17401);
and U17831 (N_17831,N_17387,N_17099);
nand U17832 (N_17832,N_17228,N_17031);
nor U17833 (N_17833,N_17386,N_17152);
or U17834 (N_17834,N_17029,N_17303);
or U17835 (N_17835,N_17166,N_17313);
xnor U17836 (N_17836,N_17419,N_17094);
nand U17837 (N_17837,N_17179,N_17174);
or U17838 (N_17838,N_17125,N_17494);
xor U17839 (N_17839,N_17468,N_17113);
xor U17840 (N_17840,N_17228,N_17224);
and U17841 (N_17841,N_17252,N_17412);
nor U17842 (N_17842,N_17364,N_17473);
nor U17843 (N_17843,N_17256,N_17491);
or U17844 (N_17844,N_17312,N_17246);
nand U17845 (N_17845,N_17045,N_17444);
and U17846 (N_17846,N_17397,N_17066);
nand U17847 (N_17847,N_17404,N_17354);
xor U17848 (N_17848,N_17012,N_17007);
nor U17849 (N_17849,N_17392,N_17284);
or U17850 (N_17850,N_17300,N_17188);
xor U17851 (N_17851,N_17468,N_17149);
and U17852 (N_17852,N_17192,N_17152);
xor U17853 (N_17853,N_17351,N_17421);
and U17854 (N_17854,N_17384,N_17387);
nand U17855 (N_17855,N_17158,N_17494);
and U17856 (N_17856,N_17006,N_17151);
xnor U17857 (N_17857,N_17000,N_17221);
and U17858 (N_17858,N_17447,N_17256);
nand U17859 (N_17859,N_17179,N_17028);
nor U17860 (N_17860,N_17191,N_17067);
and U17861 (N_17861,N_17054,N_17359);
xor U17862 (N_17862,N_17217,N_17008);
nor U17863 (N_17863,N_17441,N_17178);
nor U17864 (N_17864,N_17416,N_17030);
or U17865 (N_17865,N_17075,N_17446);
nand U17866 (N_17866,N_17037,N_17250);
xnor U17867 (N_17867,N_17148,N_17356);
nand U17868 (N_17868,N_17195,N_17122);
or U17869 (N_17869,N_17212,N_17425);
nor U17870 (N_17870,N_17363,N_17212);
xor U17871 (N_17871,N_17491,N_17316);
xnor U17872 (N_17872,N_17255,N_17097);
and U17873 (N_17873,N_17349,N_17360);
and U17874 (N_17874,N_17355,N_17292);
nor U17875 (N_17875,N_17158,N_17441);
or U17876 (N_17876,N_17216,N_17258);
and U17877 (N_17877,N_17492,N_17464);
nor U17878 (N_17878,N_17224,N_17295);
and U17879 (N_17879,N_17207,N_17382);
and U17880 (N_17880,N_17106,N_17020);
or U17881 (N_17881,N_17285,N_17009);
nor U17882 (N_17882,N_17064,N_17020);
nor U17883 (N_17883,N_17406,N_17448);
nor U17884 (N_17884,N_17368,N_17124);
nand U17885 (N_17885,N_17298,N_17477);
nand U17886 (N_17886,N_17128,N_17290);
and U17887 (N_17887,N_17185,N_17286);
nor U17888 (N_17888,N_17313,N_17156);
nor U17889 (N_17889,N_17263,N_17297);
xor U17890 (N_17890,N_17018,N_17324);
nand U17891 (N_17891,N_17487,N_17351);
nor U17892 (N_17892,N_17293,N_17413);
nor U17893 (N_17893,N_17480,N_17153);
nand U17894 (N_17894,N_17465,N_17069);
or U17895 (N_17895,N_17281,N_17323);
or U17896 (N_17896,N_17348,N_17163);
nand U17897 (N_17897,N_17390,N_17475);
and U17898 (N_17898,N_17070,N_17175);
or U17899 (N_17899,N_17228,N_17062);
or U17900 (N_17900,N_17395,N_17367);
or U17901 (N_17901,N_17193,N_17085);
nand U17902 (N_17902,N_17234,N_17305);
nor U17903 (N_17903,N_17305,N_17309);
nor U17904 (N_17904,N_17472,N_17487);
nor U17905 (N_17905,N_17397,N_17358);
or U17906 (N_17906,N_17118,N_17192);
nand U17907 (N_17907,N_17214,N_17149);
xnor U17908 (N_17908,N_17216,N_17081);
nor U17909 (N_17909,N_17292,N_17105);
or U17910 (N_17910,N_17101,N_17468);
nor U17911 (N_17911,N_17308,N_17324);
xnor U17912 (N_17912,N_17308,N_17409);
xor U17913 (N_17913,N_17293,N_17382);
nor U17914 (N_17914,N_17232,N_17086);
nand U17915 (N_17915,N_17492,N_17232);
and U17916 (N_17916,N_17209,N_17328);
or U17917 (N_17917,N_17236,N_17469);
nand U17918 (N_17918,N_17086,N_17238);
nor U17919 (N_17919,N_17464,N_17105);
or U17920 (N_17920,N_17427,N_17340);
or U17921 (N_17921,N_17357,N_17432);
nor U17922 (N_17922,N_17164,N_17294);
nand U17923 (N_17923,N_17297,N_17203);
nor U17924 (N_17924,N_17311,N_17283);
xor U17925 (N_17925,N_17296,N_17250);
and U17926 (N_17926,N_17066,N_17117);
and U17927 (N_17927,N_17201,N_17462);
or U17928 (N_17928,N_17258,N_17299);
xnor U17929 (N_17929,N_17252,N_17227);
and U17930 (N_17930,N_17491,N_17311);
xor U17931 (N_17931,N_17107,N_17090);
nor U17932 (N_17932,N_17207,N_17231);
or U17933 (N_17933,N_17049,N_17393);
and U17934 (N_17934,N_17027,N_17095);
xnor U17935 (N_17935,N_17328,N_17395);
and U17936 (N_17936,N_17149,N_17020);
or U17937 (N_17937,N_17342,N_17482);
and U17938 (N_17938,N_17203,N_17492);
xnor U17939 (N_17939,N_17399,N_17402);
nor U17940 (N_17940,N_17426,N_17321);
or U17941 (N_17941,N_17463,N_17360);
xor U17942 (N_17942,N_17468,N_17381);
nor U17943 (N_17943,N_17477,N_17250);
xnor U17944 (N_17944,N_17006,N_17204);
nor U17945 (N_17945,N_17029,N_17261);
nand U17946 (N_17946,N_17244,N_17107);
or U17947 (N_17947,N_17383,N_17321);
xor U17948 (N_17948,N_17462,N_17408);
nand U17949 (N_17949,N_17041,N_17440);
xnor U17950 (N_17950,N_17458,N_17483);
and U17951 (N_17951,N_17269,N_17238);
or U17952 (N_17952,N_17251,N_17304);
and U17953 (N_17953,N_17342,N_17087);
nor U17954 (N_17954,N_17308,N_17217);
nor U17955 (N_17955,N_17442,N_17203);
nor U17956 (N_17956,N_17490,N_17497);
and U17957 (N_17957,N_17363,N_17056);
and U17958 (N_17958,N_17194,N_17128);
or U17959 (N_17959,N_17128,N_17093);
or U17960 (N_17960,N_17461,N_17172);
xnor U17961 (N_17961,N_17031,N_17275);
xor U17962 (N_17962,N_17472,N_17458);
nor U17963 (N_17963,N_17080,N_17124);
or U17964 (N_17964,N_17496,N_17464);
and U17965 (N_17965,N_17408,N_17125);
nor U17966 (N_17966,N_17486,N_17266);
nand U17967 (N_17967,N_17188,N_17289);
xor U17968 (N_17968,N_17300,N_17336);
xor U17969 (N_17969,N_17237,N_17058);
or U17970 (N_17970,N_17367,N_17037);
xor U17971 (N_17971,N_17068,N_17192);
nand U17972 (N_17972,N_17386,N_17216);
and U17973 (N_17973,N_17275,N_17262);
nand U17974 (N_17974,N_17335,N_17430);
and U17975 (N_17975,N_17305,N_17079);
and U17976 (N_17976,N_17338,N_17375);
xor U17977 (N_17977,N_17173,N_17308);
xor U17978 (N_17978,N_17227,N_17456);
xor U17979 (N_17979,N_17251,N_17025);
xor U17980 (N_17980,N_17440,N_17497);
xnor U17981 (N_17981,N_17334,N_17181);
xor U17982 (N_17982,N_17006,N_17471);
nor U17983 (N_17983,N_17421,N_17118);
nor U17984 (N_17984,N_17040,N_17281);
xor U17985 (N_17985,N_17088,N_17014);
nand U17986 (N_17986,N_17282,N_17287);
xnor U17987 (N_17987,N_17033,N_17382);
nand U17988 (N_17988,N_17127,N_17485);
and U17989 (N_17989,N_17121,N_17186);
nand U17990 (N_17990,N_17387,N_17123);
and U17991 (N_17991,N_17334,N_17152);
and U17992 (N_17992,N_17280,N_17321);
nand U17993 (N_17993,N_17261,N_17344);
xnor U17994 (N_17994,N_17095,N_17133);
and U17995 (N_17995,N_17043,N_17328);
and U17996 (N_17996,N_17345,N_17365);
or U17997 (N_17997,N_17342,N_17344);
xnor U17998 (N_17998,N_17105,N_17288);
xnor U17999 (N_17999,N_17331,N_17243);
or U18000 (N_18000,N_17866,N_17708);
xnor U18001 (N_18001,N_17578,N_17731);
and U18002 (N_18002,N_17887,N_17624);
xor U18003 (N_18003,N_17553,N_17995);
nand U18004 (N_18004,N_17765,N_17853);
and U18005 (N_18005,N_17780,N_17689);
nor U18006 (N_18006,N_17598,N_17620);
and U18007 (N_18007,N_17536,N_17631);
and U18008 (N_18008,N_17908,N_17874);
or U18009 (N_18009,N_17792,N_17519);
nand U18010 (N_18010,N_17936,N_17638);
and U18011 (N_18011,N_17834,N_17895);
or U18012 (N_18012,N_17750,N_17757);
xor U18013 (N_18013,N_17974,N_17685);
nand U18014 (N_18014,N_17891,N_17919);
nor U18015 (N_18015,N_17705,N_17715);
and U18016 (N_18016,N_17819,N_17978);
and U18017 (N_18017,N_17735,N_17863);
or U18018 (N_18018,N_17982,N_17660);
and U18019 (N_18019,N_17861,N_17881);
nand U18020 (N_18020,N_17827,N_17549);
or U18021 (N_18021,N_17928,N_17611);
nand U18022 (N_18022,N_17589,N_17503);
nand U18023 (N_18023,N_17957,N_17865);
or U18024 (N_18024,N_17640,N_17544);
nor U18025 (N_18025,N_17949,N_17602);
nand U18026 (N_18026,N_17634,N_17858);
or U18027 (N_18027,N_17730,N_17667);
or U18028 (N_18028,N_17644,N_17524);
nand U18029 (N_18029,N_17561,N_17828);
nand U18030 (N_18030,N_17622,N_17783);
xnor U18031 (N_18031,N_17605,N_17944);
and U18032 (N_18032,N_17740,N_17693);
nand U18033 (N_18033,N_17522,N_17885);
or U18034 (N_18034,N_17969,N_17502);
or U18035 (N_18035,N_17684,N_17851);
nor U18036 (N_18036,N_17569,N_17784);
nand U18037 (N_18037,N_17512,N_17545);
or U18038 (N_18038,N_17674,N_17746);
nand U18039 (N_18039,N_17896,N_17666);
or U18040 (N_18040,N_17527,N_17902);
nor U18041 (N_18041,N_17954,N_17894);
xor U18042 (N_18042,N_17556,N_17655);
nand U18043 (N_18043,N_17868,N_17617);
nand U18044 (N_18044,N_17927,N_17651);
or U18045 (N_18045,N_17682,N_17976);
or U18046 (N_18046,N_17805,N_17809);
and U18047 (N_18047,N_17504,N_17639);
nand U18048 (N_18048,N_17714,N_17738);
nand U18049 (N_18049,N_17900,N_17755);
nor U18050 (N_18050,N_17506,N_17794);
or U18051 (N_18051,N_17511,N_17897);
or U18052 (N_18052,N_17745,N_17647);
nand U18053 (N_18053,N_17787,N_17539);
or U18054 (N_18054,N_17628,N_17642);
or U18055 (N_18055,N_17546,N_17837);
xnor U18056 (N_18056,N_17802,N_17641);
xnor U18057 (N_18057,N_17867,N_17615);
and U18058 (N_18058,N_17547,N_17904);
and U18059 (N_18059,N_17878,N_17905);
nand U18060 (N_18060,N_17998,N_17618);
and U18061 (N_18061,N_17652,N_17669);
xnor U18062 (N_18062,N_17654,N_17948);
or U18063 (N_18063,N_17576,N_17820);
nor U18064 (N_18064,N_17763,N_17818);
and U18065 (N_18065,N_17807,N_17525);
nand U18066 (N_18066,N_17847,N_17993);
xnor U18067 (N_18067,N_17515,N_17764);
or U18068 (N_18068,N_17562,N_17612);
nor U18069 (N_18069,N_17626,N_17958);
and U18070 (N_18070,N_17729,N_17687);
nor U18071 (N_18071,N_17899,N_17676);
or U18072 (N_18072,N_17945,N_17889);
nand U18073 (N_18073,N_17718,N_17580);
nand U18074 (N_18074,N_17924,N_17788);
nor U18075 (N_18075,N_17529,N_17778);
nor U18076 (N_18076,N_17551,N_17532);
and U18077 (N_18077,N_17907,N_17681);
nand U18078 (N_18078,N_17931,N_17850);
or U18079 (N_18079,N_17725,N_17796);
or U18080 (N_18080,N_17762,N_17513);
nor U18081 (N_18081,N_17776,N_17721);
and U18082 (N_18082,N_17943,N_17645);
nor U18083 (N_18083,N_17988,N_17839);
xor U18084 (N_18084,N_17803,N_17559);
or U18085 (N_18085,N_17842,N_17747);
and U18086 (N_18086,N_17930,N_17629);
xor U18087 (N_18087,N_17781,N_17859);
and U18088 (N_18088,N_17552,N_17816);
nor U18089 (N_18089,N_17711,N_17694);
nor U18090 (N_18090,N_17686,N_17806);
nor U18091 (N_18091,N_17588,N_17980);
and U18092 (N_18092,N_17779,N_17507);
xnor U18093 (N_18093,N_17953,N_17968);
or U18094 (N_18094,N_17538,N_17723);
xor U18095 (N_18095,N_17929,N_17883);
nand U18096 (N_18096,N_17751,N_17987);
nor U18097 (N_18097,N_17548,N_17966);
nand U18098 (N_18098,N_17756,N_17841);
or U18099 (N_18099,N_17554,N_17650);
nor U18100 (N_18100,N_17661,N_17568);
nand U18101 (N_18101,N_17659,N_17633);
nor U18102 (N_18102,N_17772,N_17630);
nor U18103 (N_18103,N_17508,N_17619);
or U18104 (N_18104,N_17767,N_17679);
and U18105 (N_18105,N_17872,N_17844);
xor U18106 (N_18106,N_17962,N_17994);
or U18107 (N_18107,N_17935,N_17862);
or U18108 (N_18108,N_17753,N_17520);
nor U18109 (N_18109,N_17845,N_17594);
nor U18110 (N_18110,N_17759,N_17910);
nor U18111 (N_18111,N_17574,N_17918);
xnor U18112 (N_18112,N_17952,N_17593);
or U18113 (N_18113,N_17955,N_17632);
xnor U18114 (N_18114,N_17939,N_17848);
nand U18115 (N_18115,N_17600,N_17610);
or U18116 (N_18116,N_17608,N_17852);
and U18117 (N_18117,N_17604,N_17663);
or U18118 (N_18118,N_17912,N_17956);
xor U18119 (N_18119,N_17986,N_17701);
nor U18120 (N_18120,N_17728,N_17571);
nand U18121 (N_18121,N_17843,N_17592);
or U18122 (N_18122,N_17830,N_17880);
nand U18123 (N_18123,N_17585,N_17603);
xnor U18124 (N_18124,N_17977,N_17543);
and U18125 (N_18125,N_17849,N_17744);
and U18126 (N_18126,N_17786,N_17664);
or U18127 (N_18127,N_17586,N_17517);
xor U18128 (N_18128,N_17704,N_17742);
xor U18129 (N_18129,N_17879,N_17906);
and U18130 (N_18130,N_17683,N_17675);
or U18131 (N_18131,N_17656,N_17983);
xor U18132 (N_18132,N_17771,N_17926);
nor U18133 (N_18133,N_17814,N_17570);
xor U18134 (N_18134,N_17692,N_17719);
nor U18135 (N_18135,N_17903,N_17609);
and U18136 (N_18136,N_17505,N_17500);
nand U18137 (N_18137,N_17710,N_17599);
or U18138 (N_18138,N_17768,N_17775);
or U18139 (N_18139,N_17793,N_17812);
nor U18140 (N_18140,N_17657,N_17668);
nand U18141 (N_18141,N_17825,N_17791);
nor U18142 (N_18142,N_17960,N_17871);
or U18143 (N_18143,N_17886,N_17530);
or U18144 (N_18144,N_17785,N_17990);
xnor U18145 (N_18145,N_17898,N_17916);
xor U18146 (N_18146,N_17736,N_17560);
nand U18147 (N_18147,N_17971,N_17923);
and U18148 (N_18148,N_17521,N_17933);
xnor U18149 (N_18149,N_17643,N_17777);
nand U18150 (N_18150,N_17575,N_17558);
or U18151 (N_18151,N_17909,N_17648);
nand U18152 (N_18152,N_17846,N_17790);
xnor U18153 (N_18153,N_17797,N_17514);
nor U18154 (N_18154,N_17869,N_17563);
xor U18155 (N_18155,N_17717,N_17917);
and U18156 (N_18156,N_17550,N_17537);
xnor U18157 (N_18157,N_17699,N_17613);
and U18158 (N_18158,N_17915,N_17702);
nand U18159 (N_18159,N_17534,N_17516);
nand U18160 (N_18160,N_17733,N_17541);
nor U18161 (N_18161,N_17965,N_17607);
or U18162 (N_18162,N_17596,N_17673);
and U18163 (N_18163,N_17739,N_17698);
xor U18164 (N_18164,N_17709,N_17566);
nor U18165 (N_18165,N_17985,N_17542);
and U18166 (N_18166,N_17587,N_17726);
nor U18167 (N_18167,N_17614,N_17581);
xor U18168 (N_18168,N_17691,N_17590);
and U18169 (N_18169,N_17811,N_17813);
nand U18170 (N_18170,N_17975,N_17950);
nor U18171 (N_18171,N_17821,N_17857);
or U18172 (N_18172,N_17690,N_17509);
and U18173 (N_18173,N_17680,N_17942);
nor U18174 (N_18174,N_17579,N_17959);
nor U18175 (N_18175,N_17817,N_17760);
nor U18176 (N_18176,N_17913,N_17829);
nor U18177 (N_18177,N_17637,N_17672);
nand U18178 (N_18178,N_17724,N_17662);
and U18179 (N_18179,N_17947,N_17967);
or U18180 (N_18180,N_17695,N_17557);
nor U18181 (N_18181,N_17732,N_17727);
nor U18182 (N_18182,N_17951,N_17884);
nand U18183 (N_18183,N_17540,N_17523);
nor U18184 (N_18184,N_17623,N_17749);
nand U18185 (N_18185,N_17716,N_17892);
nand U18186 (N_18186,N_17703,N_17555);
or U18187 (N_18187,N_17914,N_17621);
xor U18188 (N_18188,N_17981,N_17782);
xor U18189 (N_18189,N_17510,N_17646);
xor U18190 (N_18190,N_17526,N_17946);
xnor U18191 (N_18191,N_17815,N_17810);
and U18192 (N_18192,N_17528,N_17597);
and U18193 (N_18193,N_17582,N_17577);
and U18194 (N_18194,N_17635,N_17770);
or U18195 (N_18195,N_17921,N_17743);
nor U18196 (N_18196,N_17970,N_17808);
xnor U18197 (N_18197,N_17932,N_17713);
and U18198 (N_18198,N_17583,N_17737);
nand U18199 (N_18199,N_17761,N_17769);
nand U18200 (N_18200,N_17888,N_17573);
xor U18201 (N_18201,N_17636,N_17697);
or U18202 (N_18202,N_17855,N_17748);
or U18203 (N_18203,N_17961,N_17973);
xnor U18204 (N_18204,N_17856,N_17832);
nor U18205 (N_18205,N_17937,N_17670);
and U18206 (N_18206,N_17653,N_17696);
or U18207 (N_18207,N_17840,N_17773);
xnor U18208 (N_18208,N_17567,N_17911);
xor U18209 (N_18209,N_17616,N_17700);
nor U18210 (N_18210,N_17671,N_17501);
and U18211 (N_18211,N_17925,N_17999);
nand U18212 (N_18212,N_17875,N_17860);
xnor U18213 (N_18213,N_17940,N_17838);
nand U18214 (N_18214,N_17922,N_17722);
xnor U18215 (N_18215,N_17535,N_17707);
nor U18216 (N_18216,N_17824,N_17758);
or U18217 (N_18217,N_17997,N_17893);
nor U18218 (N_18218,N_17572,N_17833);
xor U18219 (N_18219,N_17564,N_17677);
nor U18220 (N_18220,N_17800,N_17890);
xnor U18221 (N_18221,N_17789,N_17984);
xnor U18222 (N_18222,N_17996,N_17658);
nor U18223 (N_18223,N_17795,N_17804);
or U18224 (N_18224,N_17864,N_17678);
nor U18225 (N_18225,N_17606,N_17991);
xor U18226 (N_18226,N_17531,N_17752);
and U18227 (N_18227,N_17882,N_17754);
nor U18228 (N_18228,N_17774,N_17901);
nor U18229 (N_18229,N_17720,N_17741);
and U18230 (N_18230,N_17877,N_17873);
xnor U18231 (N_18231,N_17533,N_17766);
xnor U18232 (N_18232,N_17665,N_17835);
xor U18233 (N_18233,N_17822,N_17627);
nor U18234 (N_18234,N_17979,N_17823);
nand U18235 (N_18235,N_17938,N_17876);
nand U18236 (N_18236,N_17601,N_17712);
or U18237 (N_18237,N_17565,N_17920);
xnor U18238 (N_18238,N_17992,N_17836);
nor U18239 (N_18239,N_17798,N_17518);
nor U18240 (N_18240,N_17831,N_17854);
nor U18241 (N_18241,N_17595,N_17584);
or U18242 (N_18242,N_17649,N_17934);
or U18243 (N_18243,N_17870,N_17972);
nand U18244 (N_18244,N_17591,N_17964);
or U18245 (N_18245,N_17688,N_17801);
nand U18246 (N_18246,N_17734,N_17706);
nor U18247 (N_18247,N_17941,N_17963);
and U18248 (N_18248,N_17826,N_17989);
nand U18249 (N_18249,N_17799,N_17625);
nor U18250 (N_18250,N_17626,N_17838);
or U18251 (N_18251,N_17868,N_17907);
nor U18252 (N_18252,N_17687,N_17793);
nor U18253 (N_18253,N_17964,N_17501);
nor U18254 (N_18254,N_17706,N_17767);
nand U18255 (N_18255,N_17577,N_17567);
and U18256 (N_18256,N_17816,N_17932);
nand U18257 (N_18257,N_17871,N_17908);
xor U18258 (N_18258,N_17986,N_17537);
nor U18259 (N_18259,N_17724,N_17940);
nand U18260 (N_18260,N_17767,N_17683);
and U18261 (N_18261,N_17558,N_17726);
nor U18262 (N_18262,N_17522,N_17698);
xnor U18263 (N_18263,N_17742,N_17605);
or U18264 (N_18264,N_17536,N_17928);
xor U18265 (N_18265,N_17564,N_17750);
or U18266 (N_18266,N_17853,N_17516);
and U18267 (N_18267,N_17651,N_17579);
xnor U18268 (N_18268,N_17984,N_17674);
nor U18269 (N_18269,N_17564,N_17799);
and U18270 (N_18270,N_17549,N_17868);
and U18271 (N_18271,N_17512,N_17754);
nand U18272 (N_18272,N_17955,N_17902);
nor U18273 (N_18273,N_17959,N_17930);
xnor U18274 (N_18274,N_17580,N_17663);
or U18275 (N_18275,N_17678,N_17892);
and U18276 (N_18276,N_17930,N_17717);
and U18277 (N_18277,N_17938,N_17581);
nor U18278 (N_18278,N_17656,N_17518);
or U18279 (N_18279,N_17844,N_17506);
nor U18280 (N_18280,N_17707,N_17567);
nor U18281 (N_18281,N_17822,N_17743);
xor U18282 (N_18282,N_17942,N_17745);
and U18283 (N_18283,N_17955,N_17969);
nor U18284 (N_18284,N_17710,N_17910);
nor U18285 (N_18285,N_17606,N_17536);
xor U18286 (N_18286,N_17988,N_17750);
and U18287 (N_18287,N_17709,N_17846);
and U18288 (N_18288,N_17646,N_17523);
or U18289 (N_18289,N_17782,N_17806);
and U18290 (N_18290,N_17896,N_17888);
and U18291 (N_18291,N_17623,N_17958);
and U18292 (N_18292,N_17752,N_17677);
and U18293 (N_18293,N_17783,N_17557);
nor U18294 (N_18294,N_17854,N_17516);
or U18295 (N_18295,N_17708,N_17725);
and U18296 (N_18296,N_17957,N_17758);
and U18297 (N_18297,N_17644,N_17897);
xor U18298 (N_18298,N_17896,N_17867);
or U18299 (N_18299,N_17581,N_17989);
nor U18300 (N_18300,N_17775,N_17558);
and U18301 (N_18301,N_17657,N_17958);
nand U18302 (N_18302,N_17631,N_17705);
nand U18303 (N_18303,N_17547,N_17672);
xor U18304 (N_18304,N_17712,N_17635);
nand U18305 (N_18305,N_17570,N_17580);
nor U18306 (N_18306,N_17705,N_17572);
nor U18307 (N_18307,N_17844,N_17607);
and U18308 (N_18308,N_17546,N_17654);
or U18309 (N_18309,N_17726,N_17731);
nor U18310 (N_18310,N_17772,N_17800);
nand U18311 (N_18311,N_17948,N_17617);
nor U18312 (N_18312,N_17617,N_17508);
nand U18313 (N_18313,N_17527,N_17768);
or U18314 (N_18314,N_17563,N_17561);
or U18315 (N_18315,N_17911,N_17789);
and U18316 (N_18316,N_17790,N_17928);
nand U18317 (N_18317,N_17603,N_17956);
xor U18318 (N_18318,N_17672,N_17817);
nand U18319 (N_18319,N_17646,N_17897);
nand U18320 (N_18320,N_17778,N_17686);
nand U18321 (N_18321,N_17591,N_17755);
or U18322 (N_18322,N_17715,N_17829);
nand U18323 (N_18323,N_17661,N_17760);
nand U18324 (N_18324,N_17768,N_17935);
nor U18325 (N_18325,N_17946,N_17583);
nand U18326 (N_18326,N_17975,N_17890);
and U18327 (N_18327,N_17792,N_17590);
nor U18328 (N_18328,N_17782,N_17976);
and U18329 (N_18329,N_17541,N_17603);
or U18330 (N_18330,N_17557,N_17506);
nor U18331 (N_18331,N_17504,N_17569);
nand U18332 (N_18332,N_17830,N_17611);
nor U18333 (N_18333,N_17934,N_17561);
and U18334 (N_18334,N_17607,N_17929);
xor U18335 (N_18335,N_17541,N_17814);
xnor U18336 (N_18336,N_17882,N_17835);
and U18337 (N_18337,N_17551,N_17799);
nor U18338 (N_18338,N_17823,N_17867);
nand U18339 (N_18339,N_17585,N_17928);
nor U18340 (N_18340,N_17793,N_17760);
nor U18341 (N_18341,N_17521,N_17880);
nor U18342 (N_18342,N_17514,N_17936);
nor U18343 (N_18343,N_17907,N_17876);
nor U18344 (N_18344,N_17693,N_17831);
nand U18345 (N_18345,N_17640,N_17564);
nand U18346 (N_18346,N_17681,N_17608);
xor U18347 (N_18347,N_17691,N_17566);
and U18348 (N_18348,N_17659,N_17655);
xor U18349 (N_18349,N_17842,N_17731);
xnor U18350 (N_18350,N_17782,N_17871);
xor U18351 (N_18351,N_17847,N_17611);
xnor U18352 (N_18352,N_17867,N_17922);
xor U18353 (N_18353,N_17987,N_17761);
nand U18354 (N_18354,N_17619,N_17512);
nor U18355 (N_18355,N_17917,N_17770);
or U18356 (N_18356,N_17927,N_17638);
nor U18357 (N_18357,N_17887,N_17660);
nor U18358 (N_18358,N_17770,N_17610);
nor U18359 (N_18359,N_17796,N_17735);
nand U18360 (N_18360,N_17654,N_17824);
and U18361 (N_18361,N_17701,N_17774);
nand U18362 (N_18362,N_17561,N_17986);
nand U18363 (N_18363,N_17669,N_17594);
and U18364 (N_18364,N_17694,N_17905);
nand U18365 (N_18365,N_17736,N_17784);
and U18366 (N_18366,N_17746,N_17526);
nor U18367 (N_18367,N_17868,N_17611);
nand U18368 (N_18368,N_17803,N_17935);
nor U18369 (N_18369,N_17517,N_17833);
and U18370 (N_18370,N_17699,N_17536);
nand U18371 (N_18371,N_17582,N_17726);
xor U18372 (N_18372,N_17676,N_17580);
nor U18373 (N_18373,N_17933,N_17852);
or U18374 (N_18374,N_17725,N_17676);
nand U18375 (N_18375,N_17545,N_17862);
nand U18376 (N_18376,N_17597,N_17729);
xnor U18377 (N_18377,N_17840,N_17575);
xnor U18378 (N_18378,N_17751,N_17786);
or U18379 (N_18379,N_17892,N_17970);
nand U18380 (N_18380,N_17527,N_17611);
nand U18381 (N_18381,N_17715,N_17904);
nand U18382 (N_18382,N_17989,N_17623);
nand U18383 (N_18383,N_17852,N_17648);
nor U18384 (N_18384,N_17507,N_17575);
nand U18385 (N_18385,N_17574,N_17996);
nand U18386 (N_18386,N_17783,N_17872);
and U18387 (N_18387,N_17789,N_17615);
or U18388 (N_18388,N_17936,N_17901);
xnor U18389 (N_18389,N_17910,N_17750);
or U18390 (N_18390,N_17986,N_17906);
nand U18391 (N_18391,N_17653,N_17917);
xor U18392 (N_18392,N_17509,N_17795);
nor U18393 (N_18393,N_17663,N_17979);
nand U18394 (N_18394,N_17566,N_17840);
and U18395 (N_18395,N_17716,N_17897);
xnor U18396 (N_18396,N_17628,N_17611);
xor U18397 (N_18397,N_17884,N_17746);
nor U18398 (N_18398,N_17556,N_17708);
nor U18399 (N_18399,N_17710,N_17582);
xor U18400 (N_18400,N_17916,N_17549);
xor U18401 (N_18401,N_17769,N_17891);
nand U18402 (N_18402,N_17876,N_17638);
nand U18403 (N_18403,N_17890,N_17879);
or U18404 (N_18404,N_17547,N_17829);
nand U18405 (N_18405,N_17983,N_17984);
nor U18406 (N_18406,N_17726,N_17910);
nand U18407 (N_18407,N_17884,N_17638);
nor U18408 (N_18408,N_17609,N_17516);
and U18409 (N_18409,N_17897,N_17978);
and U18410 (N_18410,N_17560,N_17887);
and U18411 (N_18411,N_17730,N_17826);
xor U18412 (N_18412,N_17848,N_17558);
xnor U18413 (N_18413,N_17502,N_17631);
and U18414 (N_18414,N_17783,N_17555);
or U18415 (N_18415,N_17948,N_17873);
nand U18416 (N_18416,N_17791,N_17540);
and U18417 (N_18417,N_17633,N_17942);
nor U18418 (N_18418,N_17616,N_17505);
or U18419 (N_18419,N_17567,N_17533);
or U18420 (N_18420,N_17949,N_17777);
nor U18421 (N_18421,N_17688,N_17893);
xnor U18422 (N_18422,N_17683,N_17765);
and U18423 (N_18423,N_17827,N_17503);
nand U18424 (N_18424,N_17787,N_17502);
or U18425 (N_18425,N_17808,N_17812);
xnor U18426 (N_18426,N_17637,N_17696);
xor U18427 (N_18427,N_17561,N_17820);
nor U18428 (N_18428,N_17717,N_17540);
nor U18429 (N_18429,N_17505,N_17881);
nand U18430 (N_18430,N_17991,N_17570);
xnor U18431 (N_18431,N_17725,N_17512);
and U18432 (N_18432,N_17679,N_17812);
xor U18433 (N_18433,N_17718,N_17861);
or U18434 (N_18434,N_17919,N_17859);
xor U18435 (N_18435,N_17771,N_17575);
xor U18436 (N_18436,N_17609,N_17933);
and U18437 (N_18437,N_17896,N_17752);
nor U18438 (N_18438,N_17957,N_17742);
and U18439 (N_18439,N_17516,N_17600);
nand U18440 (N_18440,N_17946,N_17675);
nand U18441 (N_18441,N_17825,N_17926);
nor U18442 (N_18442,N_17841,N_17942);
xor U18443 (N_18443,N_17757,N_17903);
or U18444 (N_18444,N_17750,N_17841);
nor U18445 (N_18445,N_17869,N_17986);
xor U18446 (N_18446,N_17762,N_17612);
nand U18447 (N_18447,N_17964,N_17924);
xor U18448 (N_18448,N_17776,N_17697);
nor U18449 (N_18449,N_17815,N_17634);
nor U18450 (N_18450,N_17564,N_17567);
nor U18451 (N_18451,N_17682,N_17574);
nor U18452 (N_18452,N_17975,N_17578);
and U18453 (N_18453,N_17544,N_17769);
or U18454 (N_18454,N_17564,N_17511);
nor U18455 (N_18455,N_17647,N_17940);
or U18456 (N_18456,N_17614,N_17938);
and U18457 (N_18457,N_17608,N_17974);
xnor U18458 (N_18458,N_17517,N_17952);
nand U18459 (N_18459,N_17508,N_17592);
xnor U18460 (N_18460,N_17930,N_17537);
xor U18461 (N_18461,N_17842,N_17827);
xor U18462 (N_18462,N_17649,N_17662);
or U18463 (N_18463,N_17645,N_17552);
and U18464 (N_18464,N_17814,N_17938);
nor U18465 (N_18465,N_17817,N_17908);
nor U18466 (N_18466,N_17904,N_17742);
or U18467 (N_18467,N_17519,N_17913);
xnor U18468 (N_18468,N_17813,N_17670);
or U18469 (N_18469,N_17988,N_17940);
and U18470 (N_18470,N_17698,N_17503);
or U18471 (N_18471,N_17874,N_17682);
xnor U18472 (N_18472,N_17594,N_17774);
xor U18473 (N_18473,N_17909,N_17964);
nor U18474 (N_18474,N_17744,N_17721);
xor U18475 (N_18475,N_17504,N_17604);
and U18476 (N_18476,N_17535,N_17714);
nand U18477 (N_18477,N_17923,N_17972);
or U18478 (N_18478,N_17728,N_17634);
and U18479 (N_18479,N_17969,N_17582);
xnor U18480 (N_18480,N_17976,N_17515);
nand U18481 (N_18481,N_17773,N_17581);
nor U18482 (N_18482,N_17551,N_17780);
or U18483 (N_18483,N_17694,N_17663);
nor U18484 (N_18484,N_17687,N_17933);
nand U18485 (N_18485,N_17710,N_17851);
or U18486 (N_18486,N_17547,N_17614);
nor U18487 (N_18487,N_17598,N_17922);
and U18488 (N_18488,N_17744,N_17628);
nor U18489 (N_18489,N_17943,N_17852);
xor U18490 (N_18490,N_17962,N_17991);
nor U18491 (N_18491,N_17691,N_17611);
and U18492 (N_18492,N_17661,N_17917);
or U18493 (N_18493,N_17791,N_17581);
xor U18494 (N_18494,N_17529,N_17889);
xnor U18495 (N_18495,N_17556,N_17764);
nor U18496 (N_18496,N_17686,N_17785);
or U18497 (N_18497,N_17973,N_17645);
xor U18498 (N_18498,N_17998,N_17602);
nor U18499 (N_18499,N_17735,N_17746);
xnor U18500 (N_18500,N_18310,N_18402);
nor U18501 (N_18501,N_18321,N_18173);
nand U18502 (N_18502,N_18341,N_18216);
or U18503 (N_18503,N_18292,N_18200);
or U18504 (N_18504,N_18209,N_18232);
and U18505 (N_18505,N_18248,N_18165);
nor U18506 (N_18506,N_18083,N_18231);
or U18507 (N_18507,N_18376,N_18096);
xor U18508 (N_18508,N_18259,N_18426);
and U18509 (N_18509,N_18311,N_18499);
xor U18510 (N_18510,N_18485,N_18410);
and U18511 (N_18511,N_18496,N_18421);
and U18512 (N_18512,N_18015,N_18475);
xnor U18513 (N_18513,N_18117,N_18278);
nor U18514 (N_18514,N_18211,N_18283);
or U18515 (N_18515,N_18188,N_18328);
or U18516 (N_18516,N_18220,N_18023);
and U18517 (N_18517,N_18425,N_18000);
or U18518 (N_18518,N_18408,N_18057);
nand U18519 (N_18519,N_18084,N_18423);
nand U18520 (N_18520,N_18448,N_18466);
nand U18521 (N_18521,N_18281,N_18071);
nand U18522 (N_18522,N_18093,N_18396);
xor U18523 (N_18523,N_18178,N_18493);
and U18524 (N_18524,N_18401,N_18214);
and U18525 (N_18525,N_18136,N_18424);
nand U18526 (N_18526,N_18450,N_18403);
nand U18527 (N_18527,N_18462,N_18004);
and U18528 (N_18528,N_18454,N_18273);
and U18529 (N_18529,N_18108,N_18438);
xnor U18530 (N_18530,N_18102,N_18050);
nor U18531 (N_18531,N_18497,N_18308);
and U18532 (N_18532,N_18204,N_18110);
xor U18533 (N_18533,N_18033,N_18250);
xnor U18534 (N_18534,N_18467,N_18063);
nor U18535 (N_18535,N_18460,N_18003);
nor U18536 (N_18536,N_18360,N_18413);
nand U18537 (N_18537,N_18293,N_18115);
and U18538 (N_18538,N_18473,N_18304);
or U18539 (N_18539,N_18106,N_18353);
nor U18540 (N_18540,N_18458,N_18352);
or U18541 (N_18541,N_18103,N_18290);
xnor U18542 (N_18542,N_18205,N_18262);
nand U18543 (N_18543,N_18088,N_18447);
nand U18544 (N_18544,N_18149,N_18195);
nand U18545 (N_18545,N_18040,N_18335);
nor U18546 (N_18546,N_18021,N_18182);
nand U18547 (N_18547,N_18480,N_18097);
nor U18548 (N_18548,N_18197,N_18068);
and U18549 (N_18549,N_18457,N_18201);
nor U18550 (N_18550,N_18064,N_18449);
nand U18551 (N_18551,N_18477,N_18268);
xnor U18552 (N_18552,N_18430,N_18065);
nand U18553 (N_18553,N_18280,N_18150);
xor U18554 (N_18554,N_18285,N_18339);
xnor U18555 (N_18555,N_18130,N_18440);
or U18556 (N_18556,N_18052,N_18370);
nand U18557 (N_18557,N_18443,N_18092);
nand U18558 (N_18558,N_18406,N_18212);
nand U18559 (N_18559,N_18446,N_18427);
nand U18560 (N_18560,N_18364,N_18038);
and U18561 (N_18561,N_18238,N_18398);
xnor U18562 (N_18562,N_18081,N_18010);
xnor U18563 (N_18563,N_18476,N_18251);
nand U18564 (N_18564,N_18288,N_18354);
nand U18565 (N_18565,N_18078,N_18126);
xor U18566 (N_18566,N_18367,N_18279);
nor U18567 (N_18567,N_18349,N_18305);
nor U18568 (N_18568,N_18193,N_18207);
nand U18569 (N_18569,N_18163,N_18313);
nor U18570 (N_18570,N_18124,N_18433);
xnor U18571 (N_18571,N_18488,N_18069);
xor U18572 (N_18572,N_18487,N_18148);
nand U18573 (N_18573,N_18159,N_18019);
xor U18574 (N_18574,N_18435,N_18388);
or U18575 (N_18575,N_18346,N_18415);
nor U18576 (N_18576,N_18428,N_18012);
xnor U18577 (N_18577,N_18158,N_18384);
xnor U18578 (N_18578,N_18157,N_18419);
nor U18579 (N_18579,N_18241,N_18374);
or U18580 (N_18580,N_18380,N_18274);
nand U18581 (N_18581,N_18317,N_18191);
nor U18582 (N_18582,N_18302,N_18468);
nand U18583 (N_18583,N_18162,N_18061);
xnor U18584 (N_18584,N_18330,N_18121);
nor U18585 (N_18585,N_18392,N_18147);
and U18586 (N_18586,N_18323,N_18048);
and U18587 (N_18587,N_18486,N_18383);
nor U18588 (N_18588,N_18414,N_18287);
or U18589 (N_18589,N_18264,N_18405);
nand U18590 (N_18590,N_18490,N_18138);
xnor U18591 (N_18591,N_18306,N_18483);
and U18592 (N_18592,N_18153,N_18243);
and U18593 (N_18593,N_18261,N_18263);
or U18594 (N_18594,N_18361,N_18347);
nor U18595 (N_18595,N_18340,N_18309);
xnor U18596 (N_18596,N_18312,N_18336);
nand U18597 (N_18597,N_18289,N_18058);
nor U18598 (N_18598,N_18412,N_18337);
nor U18599 (N_18599,N_18385,N_18176);
xor U18600 (N_18600,N_18420,N_18472);
or U18601 (N_18601,N_18331,N_18080);
and U18602 (N_18602,N_18436,N_18253);
xnor U18603 (N_18603,N_18318,N_18011);
nor U18604 (N_18604,N_18495,N_18391);
nand U18605 (N_18605,N_18217,N_18066);
nand U18606 (N_18606,N_18186,N_18465);
and U18607 (N_18607,N_18301,N_18053);
nor U18608 (N_18608,N_18027,N_18123);
nor U18609 (N_18609,N_18369,N_18422);
and U18610 (N_18610,N_18375,N_18351);
nor U18611 (N_18611,N_18016,N_18152);
xor U18612 (N_18612,N_18177,N_18169);
and U18613 (N_18613,N_18332,N_18164);
or U18614 (N_18614,N_18120,N_18345);
nor U18615 (N_18615,N_18362,N_18082);
nand U18616 (N_18616,N_18297,N_18041);
xor U18617 (N_18617,N_18258,N_18439);
xnor U18618 (N_18618,N_18269,N_18389);
nand U18619 (N_18619,N_18154,N_18111);
or U18620 (N_18620,N_18464,N_18194);
xnor U18621 (N_18621,N_18007,N_18031);
or U18622 (N_18622,N_18039,N_18355);
nand U18623 (N_18623,N_18125,N_18245);
xor U18624 (N_18624,N_18416,N_18067);
xor U18625 (N_18625,N_18218,N_18042);
xnor U18626 (N_18626,N_18073,N_18128);
nor U18627 (N_18627,N_18118,N_18079);
nand U18628 (N_18628,N_18129,N_18075);
or U18629 (N_18629,N_18418,N_18333);
nand U18630 (N_18630,N_18455,N_18046);
and U18631 (N_18631,N_18479,N_18030);
or U18632 (N_18632,N_18070,N_18113);
nand U18633 (N_18633,N_18225,N_18094);
nand U18634 (N_18634,N_18470,N_18303);
or U18635 (N_18635,N_18431,N_18127);
xnor U18636 (N_18636,N_18114,N_18358);
nand U18637 (N_18637,N_18397,N_18399);
nand U18638 (N_18638,N_18377,N_18095);
or U18639 (N_18639,N_18144,N_18394);
nor U18640 (N_18640,N_18298,N_18235);
and U18641 (N_18641,N_18295,N_18180);
xnor U18642 (N_18642,N_18456,N_18257);
or U18643 (N_18643,N_18233,N_18112);
and U18644 (N_18644,N_18270,N_18090);
nor U18645 (N_18645,N_18219,N_18286);
and U18646 (N_18646,N_18469,N_18453);
nor U18647 (N_18647,N_18168,N_18184);
nor U18648 (N_18648,N_18206,N_18008);
nand U18649 (N_18649,N_18109,N_18085);
nand U18650 (N_18650,N_18028,N_18196);
nand U18651 (N_18651,N_18441,N_18051);
nand U18652 (N_18652,N_18087,N_18276);
xor U18653 (N_18653,N_18224,N_18277);
xnor U18654 (N_18654,N_18284,N_18091);
xor U18655 (N_18655,N_18244,N_18463);
and U18656 (N_18656,N_18227,N_18020);
nand U18657 (N_18657,N_18307,N_18272);
and U18658 (N_18658,N_18265,N_18478);
nor U18659 (N_18659,N_18252,N_18100);
or U18660 (N_18660,N_18009,N_18494);
or U18661 (N_18661,N_18407,N_18296);
nor U18662 (N_18662,N_18359,N_18132);
or U18663 (N_18663,N_18045,N_18179);
xnor U18664 (N_18664,N_18036,N_18215);
and U18665 (N_18665,N_18099,N_18035);
xnor U18666 (N_18666,N_18137,N_18043);
or U18667 (N_18667,N_18239,N_18135);
nor U18668 (N_18668,N_18199,N_18342);
nor U18669 (N_18669,N_18255,N_18322);
nand U18670 (N_18670,N_18379,N_18260);
xnor U18671 (N_18671,N_18185,N_18017);
or U18672 (N_18672,N_18229,N_18022);
and U18673 (N_18673,N_18237,N_18300);
and U18674 (N_18674,N_18208,N_18481);
nand U18675 (N_18675,N_18242,N_18146);
or U18676 (N_18676,N_18086,N_18381);
nand U18677 (N_18677,N_18437,N_18240);
xor U18678 (N_18678,N_18056,N_18356);
xnor U18679 (N_18679,N_18172,N_18025);
nand U18680 (N_18680,N_18089,N_18059);
nand U18681 (N_18681,N_18267,N_18002);
nor U18682 (N_18682,N_18282,N_18107);
nand U18683 (N_18683,N_18160,N_18266);
nor U18684 (N_18684,N_18174,N_18451);
nand U18685 (N_18685,N_18387,N_18062);
or U18686 (N_18686,N_18432,N_18249);
or U18687 (N_18687,N_18325,N_18452);
xor U18688 (N_18688,N_18116,N_18343);
or U18689 (N_18689,N_18213,N_18210);
xor U18690 (N_18690,N_18101,N_18029);
xnor U18691 (N_18691,N_18393,N_18324);
nor U18692 (N_18692,N_18183,N_18371);
and U18693 (N_18693,N_18498,N_18156);
nand U18694 (N_18694,N_18034,N_18026);
nor U18695 (N_18695,N_18357,N_18489);
nor U18696 (N_18696,N_18143,N_18192);
or U18697 (N_18697,N_18429,N_18032);
nor U18698 (N_18698,N_18366,N_18044);
nor U18699 (N_18699,N_18400,N_18134);
xor U18700 (N_18700,N_18291,N_18098);
or U18701 (N_18701,N_18417,N_18350);
or U18702 (N_18702,N_18491,N_18319);
nor U18703 (N_18703,N_18049,N_18254);
and U18704 (N_18704,N_18326,N_18378);
nor U18705 (N_18705,N_18072,N_18459);
and U18706 (N_18706,N_18014,N_18329);
or U18707 (N_18707,N_18492,N_18334);
and U18708 (N_18708,N_18203,N_18236);
xor U18709 (N_18709,N_18442,N_18409);
xnor U18710 (N_18710,N_18372,N_18434);
nand U18711 (N_18711,N_18054,N_18404);
xor U18712 (N_18712,N_18175,N_18181);
nand U18713 (N_18713,N_18390,N_18077);
or U18714 (N_18714,N_18256,N_18226);
nor U18715 (N_18715,N_18348,N_18133);
or U18716 (N_18716,N_18018,N_18167);
and U18717 (N_18717,N_18024,N_18474);
and U18718 (N_18718,N_18141,N_18131);
or U18719 (N_18719,N_18395,N_18228);
nand U18720 (N_18720,N_18320,N_18373);
and U18721 (N_18721,N_18060,N_18365);
xor U18722 (N_18722,N_18013,N_18461);
and U18723 (N_18723,N_18338,N_18161);
nand U18724 (N_18724,N_18104,N_18247);
or U18725 (N_18725,N_18151,N_18445);
and U18726 (N_18726,N_18202,N_18316);
nand U18727 (N_18727,N_18187,N_18119);
and U18728 (N_18728,N_18166,N_18246);
and U18729 (N_18729,N_18222,N_18140);
nand U18730 (N_18730,N_18344,N_18444);
nand U18731 (N_18731,N_18299,N_18368);
xnor U18732 (N_18732,N_18411,N_18190);
or U18733 (N_18733,N_18005,N_18327);
or U18734 (N_18734,N_18382,N_18006);
nand U18735 (N_18735,N_18198,N_18074);
or U18736 (N_18736,N_18294,N_18363);
nor U18737 (N_18737,N_18275,N_18484);
and U18738 (N_18738,N_18386,N_18122);
nor U18739 (N_18739,N_18189,N_18170);
or U18740 (N_18740,N_18314,N_18223);
nor U18741 (N_18741,N_18047,N_18105);
xnor U18742 (N_18742,N_18155,N_18145);
xor U18743 (N_18743,N_18271,N_18055);
xnor U18744 (N_18744,N_18230,N_18234);
and U18745 (N_18745,N_18142,N_18001);
nand U18746 (N_18746,N_18471,N_18171);
nand U18747 (N_18747,N_18037,N_18076);
xnor U18748 (N_18748,N_18221,N_18315);
or U18749 (N_18749,N_18139,N_18482);
nor U18750 (N_18750,N_18278,N_18007);
or U18751 (N_18751,N_18402,N_18367);
nand U18752 (N_18752,N_18122,N_18014);
nor U18753 (N_18753,N_18340,N_18079);
xor U18754 (N_18754,N_18488,N_18403);
xnor U18755 (N_18755,N_18010,N_18150);
and U18756 (N_18756,N_18390,N_18394);
or U18757 (N_18757,N_18337,N_18421);
nand U18758 (N_18758,N_18462,N_18019);
and U18759 (N_18759,N_18432,N_18072);
and U18760 (N_18760,N_18028,N_18494);
nand U18761 (N_18761,N_18115,N_18384);
xor U18762 (N_18762,N_18172,N_18058);
nand U18763 (N_18763,N_18427,N_18347);
and U18764 (N_18764,N_18246,N_18277);
nor U18765 (N_18765,N_18086,N_18211);
xor U18766 (N_18766,N_18329,N_18320);
nand U18767 (N_18767,N_18231,N_18401);
and U18768 (N_18768,N_18306,N_18037);
nand U18769 (N_18769,N_18328,N_18350);
nor U18770 (N_18770,N_18089,N_18136);
or U18771 (N_18771,N_18128,N_18032);
and U18772 (N_18772,N_18036,N_18149);
nor U18773 (N_18773,N_18126,N_18041);
and U18774 (N_18774,N_18119,N_18177);
or U18775 (N_18775,N_18385,N_18255);
nand U18776 (N_18776,N_18060,N_18466);
and U18777 (N_18777,N_18076,N_18172);
nor U18778 (N_18778,N_18362,N_18312);
xnor U18779 (N_18779,N_18406,N_18118);
nor U18780 (N_18780,N_18299,N_18209);
and U18781 (N_18781,N_18056,N_18429);
nor U18782 (N_18782,N_18036,N_18289);
or U18783 (N_18783,N_18375,N_18010);
or U18784 (N_18784,N_18326,N_18198);
nand U18785 (N_18785,N_18416,N_18326);
xor U18786 (N_18786,N_18346,N_18318);
and U18787 (N_18787,N_18187,N_18480);
or U18788 (N_18788,N_18215,N_18378);
xor U18789 (N_18789,N_18096,N_18450);
nor U18790 (N_18790,N_18066,N_18468);
or U18791 (N_18791,N_18049,N_18125);
nand U18792 (N_18792,N_18352,N_18197);
xor U18793 (N_18793,N_18052,N_18463);
and U18794 (N_18794,N_18478,N_18168);
or U18795 (N_18795,N_18051,N_18100);
xnor U18796 (N_18796,N_18036,N_18123);
xor U18797 (N_18797,N_18109,N_18289);
nand U18798 (N_18798,N_18300,N_18421);
and U18799 (N_18799,N_18048,N_18256);
nor U18800 (N_18800,N_18465,N_18016);
xnor U18801 (N_18801,N_18181,N_18230);
nand U18802 (N_18802,N_18314,N_18034);
nor U18803 (N_18803,N_18175,N_18362);
and U18804 (N_18804,N_18481,N_18404);
nor U18805 (N_18805,N_18405,N_18006);
or U18806 (N_18806,N_18157,N_18319);
xnor U18807 (N_18807,N_18474,N_18327);
nand U18808 (N_18808,N_18304,N_18387);
and U18809 (N_18809,N_18013,N_18444);
or U18810 (N_18810,N_18445,N_18484);
xor U18811 (N_18811,N_18475,N_18400);
xnor U18812 (N_18812,N_18411,N_18178);
xor U18813 (N_18813,N_18064,N_18007);
and U18814 (N_18814,N_18165,N_18091);
nor U18815 (N_18815,N_18349,N_18381);
or U18816 (N_18816,N_18164,N_18160);
or U18817 (N_18817,N_18160,N_18473);
nand U18818 (N_18818,N_18211,N_18225);
and U18819 (N_18819,N_18381,N_18315);
and U18820 (N_18820,N_18373,N_18494);
and U18821 (N_18821,N_18491,N_18342);
and U18822 (N_18822,N_18467,N_18098);
xor U18823 (N_18823,N_18414,N_18347);
nor U18824 (N_18824,N_18104,N_18344);
and U18825 (N_18825,N_18262,N_18097);
or U18826 (N_18826,N_18365,N_18414);
or U18827 (N_18827,N_18356,N_18156);
and U18828 (N_18828,N_18473,N_18376);
nand U18829 (N_18829,N_18176,N_18381);
nand U18830 (N_18830,N_18180,N_18179);
and U18831 (N_18831,N_18359,N_18226);
or U18832 (N_18832,N_18498,N_18174);
xor U18833 (N_18833,N_18202,N_18201);
or U18834 (N_18834,N_18367,N_18071);
nand U18835 (N_18835,N_18456,N_18345);
and U18836 (N_18836,N_18447,N_18047);
nand U18837 (N_18837,N_18471,N_18219);
xor U18838 (N_18838,N_18277,N_18359);
or U18839 (N_18839,N_18335,N_18253);
nor U18840 (N_18840,N_18282,N_18156);
or U18841 (N_18841,N_18027,N_18158);
and U18842 (N_18842,N_18001,N_18452);
nor U18843 (N_18843,N_18396,N_18218);
or U18844 (N_18844,N_18203,N_18475);
and U18845 (N_18845,N_18337,N_18257);
or U18846 (N_18846,N_18177,N_18348);
or U18847 (N_18847,N_18270,N_18296);
nor U18848 (N_18848,N_18015,N_18024);
nor U18849 (N_18849,N_18435,N_18185);
nand U18850 (N_18850,N_18274,N_18181);
xor U18851 (N_18851,N_18193,N_18425);
or U18852 (N_18852,N_18319,N_18293);
nor U18853 (N_18853,N_18243,N_18378);
and U18854 (N_18854,N_18039,N_18010);
or U18855 (N_18855,N_18159,N_18077);
and U18856 (N_18856,N_18338,N_18283);
or U18857 (N_18857,N_18141,N_18333);
xor U18858 (N_18858,N_18018,N_18215);
nor U18859 (N_18859,N_18395,N_18191);
xor U18860 (N_18860,N_18415,N_18446);
and U18861 (N_18861,N_18055,N_18207);
and U18862 (N_18862,N_18459,N_18295);
and U18863 (N_18863,N_18152,N_18442);
xor U18864 (N_18864,N_18446,N_18067);
nor U18865 (N_18865,N_18064,N_18191);
or U18866 (N_18866,N_18374,N_18122);
and U18867 (N_18867,N_18492,N_18004);
nand U18868 (N_18868,N_18422,N_18428);
xnor U18869 (N_18869,N_18381,N_18211);
nor U18870 (N_18870,N_18079,N_18341);
xor U18871 (N_18871,N_18351,N_18162);
nand U18872 (N_18872,N_18021,N_18221);
xnor U18873 (N_18873,N_18338,N_18444);
xor U18874 (N_18874,N_18441,N_18042);
nand U18875 (N_18875,N_18452,N_18073);
nand U18876 (N_18876,N_18199,N_18047);
nand U18877 (N_18877,N_18007,N_18213);
and U18878 (N_18878,N_18317,N_18296);
xor U18879 (N_18879,N_18042,N_18140);
or U18880 (N_18880,N_18339,N_18265);
nor U18881 (N_18881,N_18026,N_18041);
and U18882 (N_18882,N_18108,N_18104);
nor U18883 (N_18883,N_18200,N_18220);
nor U18884 (N_18884,N_18141,N_18102);
nor U18885 (N_18885,N_18297,N_18499);
or U18886 (N_18886,N_18403,N_18418);
or U18887 (N_18887,N_18279,N_18106);
xnor U18888 (N_18888,N_18418,N_18440);
nand U18889 (N_18889,N_18364,N_18155);
xnor U18890 (N_18890,N_18477,N_18397);
and U18891 (N_18891,N_18410,N_18246);
nor U18892 (N_18892,N_18212,N_18131);
or U18893 (N_18893,N_18413,N_18072);
xor U18894 (N_18894,N_18175,N_18131);
or U18895 (N_18895,N_18419,N_18287);
or U18896 (N_18896,N_18322,N_18084);
nand U18897 (N_18897,N_18073,N_18052);
xnor U18898 (N_18898,N_18047,N_18107);
xor U18899 (N_18899,N_18186,N_18099);
and U18900 (N_18900,N_18493,N_18355);
nor U18901 (N_18901,N_18121,N_18270);
nand U18902 (N_18902,N_18226,N_18076);
nor U18903 (N_18903,N_18081,N_18210);
nor U18904 (N_18904,N_18404,N_18420);
and U18905 (N_18905,N_18292,N_18304);
and U18906 (N_18906,N_18468,N_18410);
or U18907 (N_18907,N_18253,N_18456);
nor U18908 (N_18908,N_18052,N_18321);
or U18909 (N_18909,N_18263,N_18428);
nand U18910 (N_18910,N_18340,N_18251);
or U18911 (N_18911,N_18253,N_18357);
nand U18912 (N_18912,N_18482,N_18328);
and U18913 (N_18913,N_18061,N_18276);
nand U18914 (N_18914,N_18372,N_18222);
nand U18915 (N_18915,N_18022,N_18416);
and U18916 (N_18916,N_18362,N_18473);
nor U18917 (N_18917,N_18168,N_18384);
nand U18918 (N_18918,N_18395,N_18370);
and U18919 (N_18919,N_18171,N_18249);
or U18920 (N_18920,N_18190,N_18452);
or U18921 (N_18921,N_18243,N_18472);
nand U18922 (N_18922,N_18019,N_18480);
or U18923 (N_18923,N_18428,N_18287);
nor U18924 (N_18924,N_18180,N_18338);
nand U18925 (N_18925,N_18478,N_18211);
and U18926 (N_18926,N_18140,N_18070);
nand U18927 (N_18927,N_18499,N_18369);
nand U18928 (N_18928,N_18444,N_18397);
or U18929 (N_18929,N_18281,N_18058);
or U18930 (N_18930,N_18034,N_18343);
and U18931 (N_18931,N_18457,N_18015);
nand U18932 (N_18932,N_18480,N_18431);
or U18933 (N_18933,N_18481,N_18416);
and U18934 (N_18934,N_18498,N_18366);
xor U18935 (N_18935,N_18007,N_18448);
or U18936 (N_18936,N_18095,N_18471);
nor U18937 (N_18937,N_18311,N_18140);
or U18938 (N_18938,N_18402,N_18412);
xor U18939 (N_18939,N_18216,N_18398);
xnor U18940 (N_18940,N_18402,N_18020);
xnor U18941 (N_18941,N_18421,N_18135);
or U18942 (N_18942,N_18165,N_18159);
and U18943 (N_18943,N_18482,N_18121);
nor U18944 (N_18944,N_18162,N_18033);
or U18945 (N_18945,N_18241,N_18378);
or U18946 (N_18946,N_18470,N_18455);
xnor U18947 (N_18947,N_18208,N_18088);
and U18948 (N_18948,N_18426,N_18013);
or U18949 (N_18949,N_18360,N_18463);
nand U18950 (N_18950,N_18083,N_18408);
xnor U18951 (N_18951,N_18224,N_18009);
nor U18952 (N_18952,N_18495,N_18437);
or U18953 (N_18953,N_18005,N_18097);
or U18954 (N_18954,N_18161,N_18258);
xor U18955 (N_18955,N_18161,N_18042);
xnor U18956 (N_18956,N_18415,N_18453);
xnor U18957 (N_18957,N_18321,N_18042);
xnor U18958 (N_18958,N_18273,N_18272);
and U18959 (N_18959,N_18380,N_18233);
xor U18960 (N_18960,N_18019,N_18104);
and U18961 (N_18961,N_18006,N_18012);
or U18962 (N_18962,N_18067,N_18268);
or U18963 (N_18963,N_18309,N_18115);
xnor U18964 (N_18964,N_18018,N_18005);
xor U18965 (N_18965,N_18425,N_18098);
and U18966 (N_18966,N_18237,N_18375);
xor U18967 (N_18967,N_18161,N_18495);
or U18968 (N_18968,N_18130,N_18268);
xnor U18969 (N_18969,N_18344,N_18096);
and U18970 (N_18970,N_18171,N_18368);
or U18971 (N_18971,N_18431,N_18089);
or U18972 (N_18972,N_18212,N_18408);
and U18973 (N_18973,N_18127,N_18252);
xor U18974 (N_18974,N_18424,N_18480);
or U18975 (N_18975,N_18163,N_18426);
and U18976 (N_18976,N_18235,N_18439);
nand U18977 (N_18977,N_18077,N_18105);
or U18978 (N_18978,N_18140,N_18016);
nand U18979 (N_18979,N_18175,N_18154);
or U18980 (N_18980,N_18473,N_18173);
and U18981 (N_18981,N_18226,N_18163);
and U18982 (N_18982,N_18002,N_18465);
or U18983 (N_18983,N_18276,N_18114);
nand U18984 (N_18984,N_18250,N_18170);
xor U18985 (N_18985,N_18294,N_18139);
and U18986 (N_18986,N_18189,N_18113);
or U18987 (N_18987,N_18335,N_18318);
xor U18988 (N_18988,N_18367,N_18467);
nor U18989 (N_18989,N_18217,N_18133);
or U18990 (N_18990,N_18490,N_18155);
and U18991 (N_18991,N_18242,N_18257);
or U18992 (N_18992,N_18062,N_18296);
nand U18993 (N_18993,N_18464,N_18400);
or U18994 (N_18994,N_18476,N_18356);
xor U18995 (N_18995,N_18073,N_18168);
xnor U18996 (N_18996,N_18246,N_18087);
or U18997 (N_18997,N_18360,N_18069);
nor U18998 (N_18998,N_18230,N_18205);
xor U18999 (N_18999,N_18040,N_18495);
nand U19000 (N_19000,N_18643,N_18866);
nand U19001 (N_19001,N_18845,N_18848);
nand U19002 (N_19002,N_18506,N_18989);
and U19003 (N_19003,N_18668,N_18929);
nor U19004 (N_19004,N_18798,N_18540);
and U19005 (N_19005,N_18712,N_18867);
nor U19006 (N_19006,N_18700,N_18896);
and U19007 (N_19007,N_18727,N_18874);
xnor U19008 (N_19008,N_18942,N_18534);
or U19009 (N_19009,N_18614,N_18851);
nand U19010 (N_19010,N_18588,N_18817);
and U19011 (N_19011,N_18559,N_18505);
nor U19012 (N_19012,N_18608,N_18923);
nor U19013 (N_19013,N_18598,N_18714);
and U19014 (N_19014,N_18770,N_18587);
and U19015 (N_19015,N_18699,N_18926);
xor U19016 (N_19016,N_18751,N_18584);
or U19017 (N_19017,N_18887,N_18661);
xnor U19018 (N_19018,N_18791,N_18600);
and U19019 (N_19019,N_18597,N_18790);
nand U19020 (N_19020,N_18758,N_18579);
or U19021 (N_19021,N_18935,N_18806);
xor U19022 (N_19022,N_18696,N_18580);
xor U19023 (N_19023,N_18826,N_18581);
xnor U19024 (N_19024,N_18898,N_18748);
or U19025 (N_19025,N_18960,N_18735);
nor U19026 (N_19026,N_18911,N_18841);
nand U19027 (N_19027,N_18992,N_18880);
and U19028 (N_19028,N_18738,N_18897);
or U19029 (N_19029,N_18623,N_18919);
nor U19030 (N_19030,N_18634,N_18788);
xnor U19031 (N_19031,N_18517,N_18903);
xor U19032 (N_19032,N_18629,N_18596);
or U19033 (N_19033,N_18924,N_18739);
and U19034 (N_19034,N_18914,N_18552);
and U19035 (N_19035,N_18594,N_18778);
nor U19036 (N_19036,N_18829,N_18538);
and U19037 (N_19037,N_18892,N_18564);
nor U19038 (N_19038,N_18721,N_18977);
and U19039 (N_19039,N_18516,N_18681);
nor U19040 (N_19040,N_18503,N_18905);
xnor U19041 (N_19041,N_18901,N_18818);
nor U19042 (N_19042,N_18764,N_18884);
nor U19043 (N_19043,N_18906,N_18653);
nand U19044 (N_19044,N_18842,N_18938);
or U19045 (N_19045,N_18998,N_18780);
or U19046 (N_19046,N_18967,N_18613);
nor U19047 (N_19047,N_18976,N_18895);
nand U19048 (N_19048,N_18774,N_18563);
nor U19049 (N_19049,N_18946,N_18719);
and U19050 (N_19050,N_18843,N_18646);
and U19051 (N_19051,N_18692,N_18978);
nand U19052 (N_19052,N_18768,N_18888);
xor U19053 (N_19053,N_18827,N_18678);
nand U19054 (N_19054,N_18518,N_18834);
or U19055 (N_19055,N_18511,N_18627);
xor U19056 (N_19056,N_18514,N_18785);
and U19057 (N_19057,N_18548,N_18837);
nor U19058 (N_19058,N_18805,N_18708);
or U19059 (N_19059,N_18592,N_18607);
and U19060 (N_19060,N_18686,N_18889);
or U19061 (N_19061,N_18756,N_18711);
xnor U19062 (N_19062,N_18986,N_18951);
xor U19063 (N_19063,N_18822,N_18713);
xnor U19064 (N_19064,N_18955,N_18695);
xor U19065 (N_19065,N_18971,N_18804);
xor U19066 (N_19066,N_18979,N_18773);
xnor U19067 (N_19067,N_18754,N_18513);
xnor U19068 (N_19068,N_18647,N_18502);
and U19069 (N_19069,N_18939,N_18900);
and U19070 (N_19070,N_18945,N_18922);
xnor U19071 (N_19071,N_18752,N_18562);
nand U19072 (N_19072,N_18832,N_18932);
nor U19073 (N_19073,N_18617,N_18725);
nor U19074 (N_19074,N_18726,N_18852);
nor U19075 (N_19075,N_18801,N_18730);
nand U19076 (N_19076,N_18861,N_18720);
xor U19077 (N_19077,N_18966,N_18674);
nand U19078 (N_19078,N_18876,N_18544);
nand U19079 (N_19079,N_18676,N_18606);
and U19080 (N_19080,N_18797,N_18512);
and U19081 (N_19081,N_18793,N_18537);
nand U19082 (N_19082,N_18515,N_18999);
or U19083 (N_19083,N_18991,N_18621);
nor U19084 (N_19084,N_18704,N_18715);
or U19085 (N_19085,N_18941,N_18523);
and U19086 (N_19086,N_18716,N_18850);
nand U19087 (N_19087,N_18765,N_18839);
xnor U19088 (N_19088,N_18710,N_18777);
nor U19089 (N_19089,N_18599,N_18844);
xor U19090 (N_19090,N_18500,N_18728);
and U19091 (N_19091,N_18632,N_18509);
or U19092 (N_19092,N_18891,N_18859);
xnor U19093 (N_19093,N_18753,N_18741);
or U19094 (N_19094,N_18959,N_18747);
nor U19095 (N_19095,N_18742,N_18988);
or U19096 (N_19096,N_18664,N_18640);
nor U19097 (N_19097,N_18908,N_18916);
and U19098 (N_19098,N_18644,N_18807);
nand U19099 (N_19099,N_18749,N_18729);
nor U19100 (N_19100,N_18902,N_18616);
or U19101 (N_19101,N_18904,N_18795);
nand U19102 (N_19102,N_18821,N_18882);
and U19103 (N_19103,N_18995,N_18682);
nor U19104 (N_19104,N_18542,N_18763);
and U19105 (N_19105,N_18803,N_18501);
xnor U19106 (N_19106,N_18810,N_18928);
xnor U19107 (N_19107,N_18820,N_18636);
nor U19108 (N_19108,N_18786,N_18886);
xnor U19109 (N_19109,N_18553,N_18865);
xor U19110 (N_19110,N_18931,N_18853);
nor U19111 (N_19111,N_18863,N_18650);
or U19112 (N_19112,N_18583,N_18521);
nand U19113 (N_19113,N_18799,N_18648);
nand U19114 (N_19114,N_18990,N_18968);
xnor U19115 (N_19115,N_18560,N_18994);
and U19116 (N_19116,N_18556,N_18925);
nand U19117 (N_19117,N_18860,N_18655);
xor U19118 (N_19118,N_18857,N_18781);
and U19119 (N_19119,N_18718,N_18809);
nand U19120 (N_19120,N_18618,N_18740);
and U19121 (N_19121,N_18524,N_18937);
and U19122 (N_19122,N_18947,N_18528);
or U19123 (N_19123,N_18709,N_18525);
nor U19124 (N_19124,N_18964,N_18586);
and U19125 (N_19125,N_18645,N_18881);
nor U19126 (N_19126,N_18766,N_18706);
nand U19127 (N_19127,N_18944,N_18543);
nor U19128 (N_19128,N_18894,N_18870);
and U19129 (N_19129,N_18918,N_18535);
or U19130 (N_19130,N_18557,N_18577);
xnor U19131 (N_19131,N_18943,N_18574);
or U19132 (N_19132,N_18522,N_18776);
and U19133 (N_19133,N_18771,N_18917);
nor U19134 (N_19134,N_18800,N_18687);
nor U19135 (N_19135,N_18659,N_18641);
nand U19136 (N_19136,N_18642,N_18769);
xnor U19137 (N_19137,N_18657,N_18536);
or U19138 (N_19138,N_18762,N_18934);
nand U19139 (N_19139,N_18656,N_18984);
and U19140 (N_19140,N_18529,N_18745);
xnor U19141 (N_19141,N_18520,N_18701);
and U19142 (N_19142,N_18877,N_18566);
and U19143 (N_19143,N_18912,N_18933);
or U19144 (N_19144,N_18733,N_18705);
nand U19145 (N_19145,N_18662,N_18619);
and U19146 (N_19146,N_18746,N_18831);
nor U19147 (N_19147,N_18972,N_18554);
xor U19148 (N_19148,N_18633,N_18508);
nor U19149 (N_19149,N_18958,N_18603);
and U19150 (N_19150,N_18823,N_18993);
and U19151 (N_19151,N_18759,N_18734);
nand U19152 (N_19152,N_18651,N_18983);
nor U19153 (N_19153,N_18787,N_18590);
nor U19154 (N_19154,N_18825,N_18789);
xnor U19155 (N_19155,N_18875,N_18915);
xor U19156 (N_19156,N_18585,N_18847);
nand U19157 (N_19157,N_18907,N_18812);
nor U19158 (N_19158,N_18626,N_18920);
or U19159 (N_19159,N_18610,N_18737);
and U19160 (N_19160,N_18814,N_18833);
nand U19161 (N_19161,N_18675,N_18702);
or U19162 (N_19162,N_18975,N_18872);
or U19163 (N_19163,N_18808,N_18707);
and U19164 (N_19164,N_18802,N_18673);
or U19165 (N_19165,N_18660,N_18813);
nor U19166 (N_19166,N_18568,N_18504);
or U19167 (N_19167,N_18816,N_18601);
xor U19168 (N_19168,N_18796,N_18824);
nor U19169 (N_19169,N_18899,N_18927);
nand U19170 (N_19170,N_18551,N_18684);
xnor U19171 (N_19171,N_18638,N_18576);
xor U19172 (N_19172,N_18772,N_18957);
nor U19173 (N_19173,N_18873,N_18565);
and U19174 (N_19174,N_18663,N_18609);
or U19175 (N_19175,N_18724,N_18703);
nand U19176 (N_19176,N_18555,N_18539);
and U19177 (N_19177,N_18996,N_18910);
xor U19178 (N_19178,N_18667,N_18624);
and U19179 (N_19179,N_18654,N_18890);
and U19180 (N_19180,N_18864,N_18533);
nand U19181 (N_19181,N_18602,N_18982);
xor U19182 (N_19182,N_18893,N_18604);
or U19183 (N_19183,N_18963,N_18591);
nor U19184 (N_19184,N_18828,N_18507);
nand U19185 (N_19185,N_18985,N_18854);
nor U19186 (N_19186,N_18558,N_18575);
or U19187 (N_19187,N_18878,N_18541);
nand U19188 (N_19188,N_18589,N_18611);
and U19189 (N_19189,N_18697,N_18547);
nand U19190 (N_19190,N_18973,N_18775);
or U19191 (N_19191,N_18858,N_18694);
and U19192 (N_19192,N_18997,N_18970);
or U19193 (N_19193,N_18936,N_18569);
nand U19194 (N_19194,N_18570,N_18838);
nand U19195 (N_19195,N_18862,N_18783);
nor U19196 (N_19196,N_18593,N_18671);
nand U19197 (N_19197,N_18595,N_18732);
nor U19198 (N_19198,N_18649,N_18652);
nand U19199 (N_19199,N_18869,N_18909);
and U19200 (N_19200,N_18981,N_18689);
or U19201 (N_19201,N_18669,N_18974);
xnor U19202 (N_19202,N_18578,N_18830);
xnor U19203 (N_19203,N_18677,N_18605);
nor U19204 (N_19204,N_18693,N_18717);
nand U19205 (N_19205,N_18620,N_18879);
nand U19206 (N_19206,N_18690,N_18962);
nor U19207 (N_19207,N_18840,N_18952);
nor U19208 (N_19208,N_18639,N_18582);
xnor U19209 (N_19209,N_18761,N_18849);
or U19210 (N_19210,N_18622,N_18868);
nor U19211 (N_19211,N_18856,N_18546);
xnor U19212 (N_19212,N_18519,N_18965);
and U19213 (N_19213,N_18680,N_18950);
or U19214 (N_19214,N_18625,N_18631);
or U19215 (N_19215,N_18571,N_18630);
or U19216 (N_19216,N_18956,N_18628);
nor U19217 (N_19217,N_18736,N_18961);
nor U19218 (N_19218,N_18871,N_18510);
nor U19219 (N_19219,N_18921,N_18637);
and U19220 (N_19220,N_18954,N_18672);
nor U19221 (N_19221,N_18635,N_18811);
nand U19222 (N_19222,N_18930,N_18683);
nor U19223 (N_19223,N_18527,N_18750);
nand U19224 (N_19224,N_18691,N_18685);
and U19225 (N_19225,N_18567,N_18782);
and U19226 (N_19226,N_18670,N_18744);
nor U19227 (N_19227,N_18836,N_18679);
or U19228 (N_19228,N_18794,N_18784);
xor U19229 (N_19229,N_18698,N_18835);
nor U19230 (N_19230,N_18612,N_18530);
nand U19231 (N_19231,N_18767,N_18815);
nand U19232 (N_19232,N_18757,N_18987);
and U19233 (N_19233,N_18723,N_18940);
and U19234 (N_19234,N_18666,N_18855);
or U19235 (N_19235,N_18953,N_18913);
and U19236 (N_19236,N_18819,N_18779);
xor U19237 (N_19237,N_18549,N_18526);
and U19238 (N_19238,N_18722,N_18550);
xor U19239 (N_19239,N_18846,N_18948);
or U19240 (N_19240,N_18883,N_18665);
or U19241 (N_19241,N_18949,N_18792);
and U19242 (N_19242,N_18969,N_18755);
nand U19243 (N_19243,N_18561,N_18731);
and U19244 (N_19244,N_18688,N_18573);
and U19245 (N_19245,N_18658,N_18743);
nor U19246 (N_19246,N_18572,N_18615);
and U19247 (N_19247,N_18760,N_18531);
or U19248 (N_19248,N_18885,N_18532);
or U19249 (N_19249,N_18980,N_18545);
nor U19250 (N_19250,N_18897,N_18502);
nand U19251 (N_19251,N_18909,N_18918);
xor U19252 (N_19252,N_18640,N_18579);
nand U19253 (N_19253,N_18675,N_18722);
xor U19254 (N_19254,N_18868,N_18715);
or U19255 (N_19255,N_18959,N_18673);
nand U19256 (N_19256,N_18573,N_18773);
nand U19257 (N_19257,N_18781,N_18748);
nor U19258 (N_19258,N_18551,N_18997);
or U19259 (N_19259,N_18796,N_18523);
xnor U19260 (N_19260,N_18819,N_18718);
xnor U19261 (N_19261,N_18748,N_18951);
xnor U19262 (N_19262,N_18605,N_18544);
or U19263 (N_19263,N_18640,N_18747);
nand U19264 (N_19264,N_18796,N_18772);
nand U19265 (N_19265,N_18755,N_18711);
nor U19266 (N_19266,N_18959,N_18671);
nand U19267 (N_19267,N_18506,N_18599);
or U19268 (N_19268,N_18886,N_18586);
nor U19269 (N_19269,N_18880,N_18897);
or U19270 (N_19270,N_18869,N_18789);
or U19271 (N_19271,N_18863,N_18869);
or U19272 (N_19272,N_18778,N_18940);
xnor U19273 (N_19273,N_18925,N_18948);
nand U19274 (N_19274,N_18608,N_18893);
nand U19275 (N_19275,N_18695,N_18712);
or U19276 (N_19276,N_18570,N_18670);
and U19277 (N_19277,N_18976,N_18840);
nand U19278 (N_19278,N_18679,N_18605);
or U19279 (N_19279,N_18996,N_18694);
xor U19280 (N_19280,N_18734,N_18629);
nor U19281 (N_19281,N_18940,N_18757);
and U19282 (N_19282,N_18984,N_18683);
and U19283 (N_19283,N_18517,N_18779);
or U19284 (N_19284,N_18877,N_18794);
and U19285 (N_19285,N_18665,N_18865);
nand U19286 (N_19286,N_18583,N_18998);
or U19287 (N_19287,N_18586,N_18603);
or U19288 (N_19288,N_18936,N_18521);
xor U19289 (N_19289,N_18837,N_18804);
and U19290 (N_19290,N_18524,N_18783);
xnor U19291 (N_19291,N_18539,N_18797);
nand U19292 (N_19292,N_18967,N_18850);
or U19293 (N_19293,N_18545,N_18641);
nand U19294 (N_19294,N_18730,N_18568);
nor U19295 (N_19295,N_18634,N_18802);
nor U19296 (N_19296,N_18922,N_18970);
xor U19297 (N_19297,N_18504,N_18836);
xnor U19298 (N_19298,N_18693,N_18724);
xnor U19299 (N_19299,N_18548,N_18633);
nor U19300 (N_19300,N_18737,N_18738);
and U19301 (N_19301,N_18994,N_18878);
nor U19302 (N_19302,N_18680,N_18854);
or U19303 (N_19303,N_18802,N_18886);
or U19304 (N_19304,N_18693,N_18572);
nor U19305 (N_19305,N_18756,N_18840);
xor U19306 (N_19306,N_18959,N_18773);
xor U19307 (N_19307,N_18638,N_18872);
nor U19308 (N_19308,N_18694,N_18734);
xnor U19309 (N_19309,N_18500,N_18682);
nand U19310 (N_19310,N_18849,N_18920);
nor U19311 (N_19311,N_18830,N_18681);
nor U19312 (N_19312,N_18944,N_18817);
nand U19313 (N_19313,N_18633,N_18945);
xor U19314 (N_19314,N_18624,N_18817);
and U19315 (N_19315,N_18811,N_18576);
xnor U19316 (N_19316,N_18869,N_18589);
or U19317 (N_19317,N_18998,N_18537);
nor U19318 (N_19318,N_18675,N_18872);
and U19319 (N_19319,N_18851,N_18860);
xnor U19320 (N_19320,N_18966,N_18752);
nand U19321 (N_19321,N_18757,N_18713);
nand U19322 (N_19322,N_18941,N_18648);
and U19323 (N_19323,N_18700,N_18824);
and U19324 (N_19324,N_18842,N_18730);
nand U19325 (N_19325,N_18733,N_18724);
nor U19326 (N_19326,N_18955,N_18614);
nand U19327 (N_19327,N_18688,N_18592);
xnor U19328 (N_19328,N_18745,N_18786);
nor U19329 (N_19329,N_18675,N_18951);
nand U19330 (N_19330,N_18892,N_18760);
nor U19331 (N_19331,N_18858,N_18629);
and U19332 (N_19332,N_18786,N_18989);
nand U19333 (N_19333,N_18715,N_18731);
nand U19334 (N_19334,N_18523,N_18982);
or U19335 (N_19335,N_18964,N_18750);
or U19336 (N_19336,N_18881,N_18616);
xnor U19337 (N_19337,N_18541,N_18883);
nand U19338 (N_19338,N_18527,N_18676);
nor U19339 (N_19339,N_18936,N_18937);
or U19340 (N_19340,N_18849,N_18913);
or U19341 (N_19341,N_18763,N_18859);
or U19342 (N_19342,N_18546,N_18847);
xor U19343 (N_19343,N_18661,N_18533);
and U19344 (N_19344,N_18861,N_18793);
and U19345 (N_19345,N_18799,N_18610);
and U19346 (N_19346,N_18852,N_18554);
and U19347 (N_19347,N_18759,N_18569);
and U19348 (N_19348,N_18751,N_18719);
nand U19349 (N_19349,N_18719,N_18866);
xor U19350 (N_19350,N_18889,N_18694);
nor U19351 (N_19351,N_18739,N_18630);
nand U19352 (N_19352,N_18693,N_18685);
nor U19353 (N_19353,N_18897,N_18806);
and U19354 (N_19354,N_18559,N_18551);
xnor U19355 (N_19355,N_18696,N_18677);
nand U19356 (N_19356,N_18528,N_18803);
and U19357 (N_19357,N_18567,N_18571);
nor U19358 (N_19358,N_18746,N_18888);
xor U19359 (N_19359,N_18939,N_18617);
xnor U19360 (N_19360,N_18555,N_18666);
and U19361 (N_19361,N_18719,N_18593);
xnor U19362 (N_19362,N_18574,N_18631);
or U19363 (N_19363,N_18856,N_18921);
nor U19364 (N_19364,N_18833,N_18768);
and U19365 (N_19365,N_18622,N_18785);
nor U19366 (N_19366,N_18844,N_18576);
nor U19367 (N_19367,N_18680,N_18920);
nor U19368 (N_19368,N_18569,N_18943);
nand U19369 (N_19369,N_18962,N_18698);
or U19370 (N_19370,N_18665,N_18944);
xnor U19371 (N_19371,N_18807,N_18717);
nor U19372 (N_19372,N_18684,N_18538);
nor U19373 (N_19373,N_18993,N_18920);
nand U19374 (N_19374,N_18811,N_18998);
nor U19375 (N_19375,N_18692,N_18660);
xor U19376 (N_19376,N_18781,N_18562);
and U19377 (N_19377,N_18752,N_18787);
nor U19378 (N_19378,N_18646,N_18518);
nor U19379 (N_19379,N_18743,N_18604);
nor U19380 (N_19380,N_18611,N_18945);
and U19381 (N_19381,N_18960,N_18928);
or U19382 (N_19382,N_18826,N_18721);
nand U19383 (N_19383,N_18842,N_18547);
or U19384 (N_19384,N_18521,N_18743);
nor U19385 (N_19385,N_18784,N_18756);
or U19386 (N_19386,N_18829,N_18965);
or U19387 (N_19387,N_18658,N_18551);
nor U19388 (N_19388,N_18903,N_18915);
xor U19389 (N_19389,N_18785,N_18910);
nor U19390 (N_19390,N_18735,N_18527);
and U19391 (N_19391,N_18563,N_18901);
xnor U19392 (N_19392,N_18653,N_18680);
nor U19393 (N_19393,N_18849,N_18576);
or U19394 (N_19394,N_18863,N_18872);
xor U19395 (N_19395,N_18514,N_18649);
and U19396 (N_19396,N_18979,N_18594);
or U19397 (N_19397,N_18922,N_18604);
nor U19398 (N_19398,N_18521,N_18866);
nand U19399 (N_19399,N_18994,N_18959);
or U19400 (N_19400,N_18541,N_18793);
xnor U19401 (N_19401,N_18553,N_18942);
nor U19402 (N_19402,N_18668,N_18667);
or U19403 (N_19403,N_18560,N_18537);
nor U19404 (N_19404,N_18937,N_18905);
or U19405 (N_19405,N_18606,N_18966);
or U19406 (N_19406,N_18761,N_18756);
nand U19407 (N_19407,N_18837,N_18511);
nor U19408 (N_19408,N_18611,N_18771);
nor U19409 (N_19409,N_18800,N_18866);
and U19410 (N_19410,N_18562,N_18815);
nor U19411 (N_19411,N_18566,N_18901);
nand U19412 (N_19412,N_18894,N_18865);
or U19413 (N_19413,N_18877,N_18684);
and U19414 (N_19414,N_18849,N_18781);
and U19415 (N_19415,N_18835,N_18989);
and U19416 (N_19416,N_18642,N_18988);
or U19417 (N_19417,N_18840,N_18748);
xor U19418 (N_19418,N_18900,N_18931);
and U19419 (N_19419,N_18956,N_18902);
xnor U19420 (N_19420,N_18857,N_18636);
or U19421 (N_19421,N_18948,N_18899);
nor U19422 (N_19422,N_18683,N_18895);
nor U19423 (N_19423,N_18791,N_18593);
or U19424 (N_19424,N_18653,N_18889);
nand U19425 (N_19425,N_18564,N_18528);
xnor U19426 (N_19426,N_18825,N_18764);
nor U19427 (N_19427,N_18709,N_18853);
nor U19428 (N_19428,N_18708,N_18948);
and U19429 (N_19429,N_18798,N_18634);
nor U19430 (N_19430,N_18770,N_18911);
nand U19431 (N_19431,N_18590,N_18729);
nand U19432 (N_19432,N_18760,N_18911);
and U19433 (N_19433,N_18994,N_18601);
nor U19434 (N_19434,N_18808,N_18820);
xnor U19435 (N_19435,N_18854,N_18537);
xor U19436 (N_19436,N_18951,N_18709);
xnor U19437 (N_19437,N_18916,N_18969);
and U19438 (N_19438,N_18975,N_18736);
or U19439 (N_19439,N_18696,N_18658);
xor U19440 (N_19440,N_18526,N_18590);
or U19441 (N_19441,N_18660,N_18606);
nor U19442 (N_19442,N_18947,N_18877);
nor U19443 (N_19443,N_18890,N_18692);
xor U19444 (N_19444,N_18614,N_18861);
nor U19445 (N_19445,N_18874,N_18628);
or U19446 (N_19446,N_18942,N_18529);
and U19447 (N_19447,N_18836,N_18877);
nand U19448 (N_19448,N_18520,N_18738);
xor U19449 (N_19449,N_18900,N_18798);
and U19450 (N_19450,N_18818,N_18632);
xor U19451 (N_19451,N_18895,N_18866);
or U19452 (N_19452,N_18501,N_18636);
nor U19453 (N_19453,N_18751,N_18703);
and U19454 (N_19454,N_18795,N_18941);
xnor U19455 (N_19455,N_18596,N_18956);
nor U19456 (N_19456,N_18668,N_18671);
nor U19457 (N_19457,N_18745,N_18804);
and U19458 (N_19458,N_18824,N_18502);
nor U19459 (N_19459,N_18563,N_18722);
nand U19460 (N_19460,N_18860,N_18576);
and U19461 (N_19461,N_18707,N_18539);
nor U19462 (N_19462,N_18666,N_18706);
and U19463 (N_19463,N_18803,N_18586);
nor U19464 (N_19464,N_18698,N_18975);
xor U19465 (N_19465,N_18757,N_18712);
xnor U19466 (N_19466,N_18759,N_18541);
nor U19467 (N_19467,N_18791,N_18869);
nor U19468 (N_19468,N_18984,N_18814);
nand U19469 (N_19469,N_18689,N_18672);
or U19470 (N_19470,N_18891,N_18605);
or U19471 (N_19471,N_18850,N_18824);
nand U19472 (N_19472,N_18964,N_18869);
or U19473 (N_19473,N_18947,N_18583);
or U19474 (N_19474,N_18890,N_18900);
xor U19475 (N_19475,N_18715,N_18618);
nor U19476 (N_19476,N_18940,N_18794);
nor U19477 (N_19477,N_18811,N_18694);
or U19478 (N_19478,N_18993,N_18515);
xnor U19479 (N_19479,N_18661,N_18864);
and U19480 (N_19480,N_18686,N_18881);
and U19481 (N_19481,N_18982,N_18731);
nor U19482 (N_19482,N_18602,N_18705);
and U19483 (N_19483,N_18926,N_18603);
nor U19484 (N_19484,N_18888,N_18764);
and U19485 (N_19485,N_18689,N_18678);
and U19486 (N_19486,N_18931,N_18997);
or U19487 (N_19487,N_18969,N_18936);
nor U19488 (N_19488,N_18950,N_18908);
nand U19489 (N_19489,N_18633,N_18950);
xnor U19490 (N_19490,N_18999,N_18584);
and U19491 (N_19491,N_18996,N_18715);
or U19492 (N_19492,N_18517,N_18641);
nor U19493 (N_19493,N_18743,N_18613);
nor U19494 (N_19494,N_18812,N_18891);
or U19495 (N_19495,N_18569,N_18967);
or U19496 (N_19496,N_18698,N_18804);
xnor U19497 (N_19497,N_18685,N_18922);
or U19498 (N_19498,N_18768,N_18764);
or U19499 (N_19499,N_18572,N_18877);
nor U19500 (N_19500,N_19152,N_19183);
and U19501 (N_19501,N_19460,N_19025);
nand U19502 (N_19502,N_19039,N_19060);
nand U19503 (N_19503,N_19229,N_19361);
or U19504 (N_19504,N_19096,N_19150);
and U19505 (N_19505,N_19018,N_19443);
xnor U19506 (N_19506,N_19478,N_19357);
and U19507 (N_19507,N_19250,N_19132);
nor U19508 (N_19508,N_19270,N_19212);
or U19509 (N_19509,N_19027,N_19348);
and U19510 (N_19510,N_19123,N_19404);
or U19511 (N_19511,N_19490,N_19251);
and U19512 (N_19512,N_19344,N_19078);
nor U19513 (N_19513,N_19484,N_19493);
and U19514 (N_19514,N_19035,N_19492);
nor U19515 (N_19515,N_19408,N_19365);
xor U19516 (N_19516,N_19059,N_19378);
and U19517 (N_19517,N_19353,N_19068);
xnor U19518 (N_19518,N_19214,N_19444);
nand U19519 (N_19519,N_19433,N_19128);
and U19520 (N_19520,N_19127,N_19049);
or U19521 (N_19521,N_19189,N_19446);
or U19522 (N_19522,N_19358,N_19331);
xor U19523 (N_19523,N_19261,N_19439);
nor U19524 (N_19524,N_19436,N_19188);
or U19525 (N_19525,N_19120,N_19376);
xor U19526 (N_19526,N_19418,N_19090);
xnor U19527 (N_19527,N_19073,N_19240);
xnor U19528 (N_19528,N_19031,N_19021);
or U19529 (N_19529,N_19368,N_19165);
and U19530 (N_19530,N_19017,N_19317);
or U19531 (N_19531,N_19464,N_19466);
nor U19532 (N_19532,N_19015,N_19161);
nand U19533 (N_19533,N_19101,N_19156);
or U19534 (N_19534,N_19461,N_19327);
and U19535 (N_19535,N_19177,N_19019);
xnor U19536 (N_19536,N_19205,N_19431);
nor U19537 (N_19537,N_19372,N_19472);
xor U19538 (N_19538,N_19405,N_19497);
or U19539 (N_19539,N_19275,N_19070);
or U19540 (N_19540,N_19076,N_19098);
xnor U19541 (N_19541,N_19005,N_19476);
or U19542 (N_19542,N_19412,N_19028);
or U19543 (N_19543,N_19263,N_19211);
or U19544 (N_19544,N_19370,N_19075);
nor U19545 (N_19545,N_19350,N_19245);
xnor U19546 (N_19546,N_19080,N_19091);
nor U19547 (N_19547,N_19465,N_19232);
nand U19548 (N_19548,N_19224,N_19193);
or U19549 (N_19549,N_19118,N_19360);
xor U19550 (N_19550,N_19470,N_19299);
nor U19551 (N_19551,N_19174,N_19238);
and U19552 (N_19552,N_19410,N_19341);
and U19553 (N_19553,N_19155,N_19323);
and U19554 (N_19554,N_19169,N_19064);
nor U19555 (N_19555,N_19151,N_19011);
nand U19556 (N_19556,N_19382,N_19312);
nor U19557 (N_19557,N_19416,N_19434);
xnor U19558 (N_19558,N_19399,N_19255);
or U19559 (N_19559,N_19103,N_19475);
nor U19560 (N_19560,N_19029,N_19373);
and U19561 (N_19561,N_19053,N_19225);
nand U19562 (N_19562,N_19398,N_19283);
nor U19563 (N_19563,N_19311,N_19402);
nand U19564 (N_19564,N_19253,N_19095);
or U19565 (N_19565,N_19202,N_19149);
nand U19566 (N_19566,N_19289,N_19236);
nand U19567 (N_19567,N_19292,N_19326);
nor U19568 (N_19568,N_19087,N_19142);
and U19569 (N_19569,N_19257,N_19206);
and U19570 (N_19570,N_19097,N_19030);
and U19571 (N_19571,N_19131,N_19159);
nand U19572 (N_19572,N_19221,N_19305);
xor U19573 (N_19573,N_19249,N_19425);
nand U19574 (N_19574,N_19279,N_19204);
or U19575 (N_19575,N_19298,N_19172);
xor U19576 (N_19576,N_19109,N_19459);
or U19577 (N_19577,N_19483,N_19141);
xor U19578 (N_19578,N_19429,N_19247);
nand U19579 (N_19579,N_19072,N_19296);
and U19580 (N_19580,N_19194,N_19414);
and U19581 (N_19581,N_19044,N_19387);
or U19582 (N_19582,N_19208,N_19220);
and U19583 (N_19583,N_19364,N_19215);
nor U19584 (N_19584,N_19456,N_19138);
xor U19585 (N_19585,N_19084,N_19010);
nand U19586 (N_19586,N_19145,N_19187);
xor U19587 (N_19587,N_19040,N_19033);
or U19588 (N_19588,N_19244,N_19020);
nor U19589 (N_19589,N_19394,N_19494);
xor U19590 (N_19590,N_19036,N_19351);
or U19591 (N_19591,N_19200,N_19432);
nor U19592 (N_19592,N_19014,N_19280);
and U19593 (N_19593,N_19302,N_19467);
nor U19594 (N_19594,N_19393,N_19337);
xnor U19595 (N_19595,N_19316,N_19003);
and U19596 (N_19596,N_19451,N_19210);
and U19597 (N_19597,N_19117,N_19181);
nor U19598 (N_19598,N_19157,N_19207);
nand U19599 (N_19599,N_19310,N_19479);
nand U19600 (N_19600,N_19108,N_19486);
and U19601 (N_19601,N_19314,N_19306);
nand U19602 (N_19602,N_19498,N_19260);
nand U19603 (N_19603,N_19496,N_19377);
or U19604 (N_19604,N_19241,N_19171);
nor U19605 (N_19605,N_19111,N_19162);
and U19606 (N_19606,N_19092,N_19457);
nand U19607 (N_19607,N_19288,N_19175);
and U19608 (N_19608,N_19153,N_19160);
nor U19609 (N_19609,N_19233,N_19166);
nand U19610 (N_19610,N_19234,N_19058);
or U19611 (N_19611,N_19178,N_19334);
nand U19612 (N_19612,N_19158,N_19321);
nor U19613 (N_19613,N_19421,N_19170);
xnor U19614 (N_19614,N_19458,N_19196);
nor U19615 (N_19615,N_19422,N_19216);
or U19616 (N_19616,N_19054,N_19026);
nor U19617 (N_19617,N_19329,N_19235);
xnor U19618 (N_19618,N_19455,N_19413);
nand U19619 (N_19619,N_19340,N_19300);
and U19620 (N_19620,N_19093,N_19391);
or U19621 (N_19621,N_19066,N_19012);
nor U19622 (N_19622,N_19488,N_19309);
and U19623 (N_19623,N_19185,N_19006);
and U19624 (N_19624,N_19315,N_19385);
and U19625 (N_19625,N_19230,N_19007);
nor U19626 (N_19626,N_19223,N_19441);
xnor U19627 (N_19627,N_19154,N_19146);
and U19628 (N_19628,N_19386,N_19148);
or U19629 (N_19629,N_19190,N_19231);
and U19630 (N_19630,N_19081,N_19065);
nor U19631 (N_19631,N_19445,N_19367);
or U19632 (N_19632,N_19400,N_19083);
and U19633 (N_19633,N_19002,N_19411);
or U19634 (N_19634,N_19415,N_19375);
or U19635 (N_19635,N_19342,N_19034);
or U19636 (N_19636,N_19469,N_19038);
or U19637 (N_19637,N_19480,N_19287);
nor U19638 (N_19638,N_19045,N_19004);
or U19639 (N_19639,N_19048,N_19116);
or U19640 (N_19640,N_19099,N_19126);
or U19641 (N_19641,N_19499,N_19063);
or U19642 (N_19642,N_19228,N_19359);
or U19643 (N_19643,N_19392,N_19055);
xor U19644 (N_19644,N_19403,N_19167);
nand U19645 (N_19645,N_19285,N_19114);
and U19646 (N_19646,N_19435,N_19173);
nand U19647 (N_19647,N_19071,N_19105);
or U19648 (N_19648,N_19143,N_19136);
and U19649 (N_19649,N_19395,N_19354);
nand U19650 (N_19650,N_19213,N_19086);
nor U19651 (N_19651,N_19452,N_19121);
and U19652 (N_19652,N_19369,N_19265);
nand U19653 (N_19653,N_19267,N_19226);
nor U19654 (N_19654,N_19390,N_19450);
xor U19655 (N_19655,N_19407,N_19428);
or U19656 (N_19656,N_19176,N_19102);
nor U19657 (N_19657,N_19266,N_19009);
xor U19658 (N_19658,N_19104,N_19366);
or U19659 (N_19659,N_19140,N_19198);
and U19660 (N_19660,N_19352,N_19164);
and U19661 (N_19661,N_19243,N_19124);
or U19662 (N_19662,N_19339,N_19277);
and U19663 (N_19663,N_19088,N_19082);
or U19664 (N_19664,N_19381,N_19282);
xnor U19665 (N_19665,N_19333,N_19318);
nand U19666 (N_19666,N_19453,N_19325);
nor U19667 (N_19667,N_19023,N_19454);
and U19668 (N_19668,N_19384,N_19113);
or U19669 (N_19669,N_19135,N_19191);
xor U19670 (N_19670,N_19423,N_19089);
nor U19671 (N_19671,N_19262,N_19284);
and U19672 (N_19672,N_19345,N_19290);
or U19673 (N_19673,N_19301,N_19122);
xnor U19674 (N_19674,N_19374,N_19192);
and U19675 (N_19675,N_19074,N_19319);
and U19676 (N_19676,N_19248,N_19179);
and U19677 (N_19677,N_19383,N_19056);
nand U19678 (N_19678,N_19069,N_19438);
xor U19679 (N_19679,N_19022,N_19379);
or U19680 (N_19680,N_19491,N_19471);
or U19681 (N_19681,N_19129,N_19426);
xor U19682 (N_19682,N_19349,N_19217);
nor U19683 (N_19683,N_19037,N_19106);
or U19684 (N_19684,N_19406,N_19050);
or U19685 (N_19685,N_19272,N_19042);
or U19686 (N_19686,N_19297,N_19303);
and U19687 (N_19687,N_19420,N_19330);
nand U19688 (N_19688,N_19100,N_19184);
nor U19689 (N_19689,N_19447,N_19313);
or U19690 (N_19690,N_19481,N_19147);
nor U19691 (N_19691,N_19258,N_19335);
nand U19692 (N_19692,N_19079,N_19473);
or U19693 (N_19693,N_19139,N_19409);
xnor U19694 (N_19694,N_19041,N_19362);
xnor U19695 (N_19695,N_19067,N_19448);
nand U19696 (N_19696,N_19252,N_19237);
and U19697 (N_19697,N_19427,N_19324);
and U19698 (N_19698,N_19242,N_19201);
and U19699 (N_19699,N_19485,N_19489);
nand U19700 (N_19700,N_19032,N_19264);
and U19701 (N_19701,N_19195,N_19094);
nand U19702 (N_19702,N_19008,N_19013);
xor U19703 (N_19703,N_19462,N_19371);
nand U19704 (N_19704,N_19168,N_19278);
or U19705 (N_19705,N_19062,N_19273);
nand U19706 (N_19706,N_19218,N_19293);
and U19707 (N_19707,N_19380,N_19199);
and U19708 (N_19708,N_19107,N_19442);
or U19709 (N_19709,N_19449,N_19125);
xor U19710 (N_19710,N_19222,N_19307);
xnor U19711 (N_19711,N_19430,N_19197);
or U19712 (N_19712,N_19047,N_19137);
nor U19713 (N_19713,N_19363,N_19269);
and U19714 (N_19714,N_19052,N_19209);
or U19715 (N_19715,N_19468,N_19332);
xor U19716 (N_19716,N_19322,N_19396);
and U19717 (N_19717,N_19051,N_19268);
nor U19718 (N_19718,N_19061,N_19239);
or U19719 (N_19719,N_19227,N_19336);
xor U19720 (N_19720,N_19437,N_19046);
nor U19721 (N_19721,N_19308,N_19203);
nor U19722 (N_19722,N_19115,N_19182);
or U19723 (N_19723,N_19417,N_19487);
or U19724 (N_19724,N_19256,N_19440);
nand U19725 (N_19725,N_19424,N_19133);
xnor U19726 (N_19726,N_19043,N_19495);
nor U19727 (N_19727,N_19016,N_19355);
and U19728 (N_19728,N_19291,N_19295);
and U19729 (N_19729,N_19271,N_19338);
or U19730 (N_19730,N_19130,N_19419);
nor U19731 (N_19731,N_19000,N_19294);
nand U19732 (N_19732,N_19119,N_19246);
or U19733 (N_19733,N_19144,N_19389);
xnor U19734 (N_19734,N_19085,N_19259);
and U19735 (N_19735,N_19463,N_19281);
or U19736 (N_19736,N_19057,N_19343);
xnor U19737 (N_19737,N_19219,N_19474);
nand U19738 (N_19738,N_19001,N_19328);
nand U19739 (N_19739,N_19347,N_19077);
nand U19740 (N_19740,N_19254,N_19110);
and U19741 (N_19741,N_19346,N_19482);
nand U19742 (N_19742,N_19477,N_19286);
and U19743 (N_19743,N_19276,N_19320);
and U19744 (N_19744,N_19024,N_19180);
nor U19745 (N_19745,N_19134,N_19397);
or U19746 (N_19746,N_19388,N_19304);
nand U19747 (N_19747,N_19356,N_19274);
xnor U19748 (N_19748,N_19401,N_19112);
xor U19749 (N_19749,N_19186,N_19163);
nor U19750 (N_19750,N_19394,N_19122);
and U19751 (N_19751,N_19280,N_19247);
nand U19752 (N_19752,N_19034,N_19305);
nor U19753 (N_19753,N_19381,N_19129);
nand U19754 (N_19754,N_19287,N_19156);
or U19755 (N_19755,N_19240,N_19353);
xor U19756 (N_19756,N_19341,N_19412);
and U19757 (N_19757,N_19495,N_19187);
nor U19758 (N_19758,N_19344,N_19045);
and U19759 (N_19759,N_19313,N_19158);
nand U19760 (N_19760,N_19072,N_19000);
nor U19761 (N_19761,N_19074,N_19084);
or U19762 (N_19762,N_19159,N_19023);
or U19763 (N_19763,N_19196,N_19275);
nor U19764 (N_19764,N_19070,N_19420);
xnor U19765 (N_19765,N_19394,N_19170);
nand U19766 (N_19766,N_19488,N_19377);
or U19767 (N_19767,N_19447,N_19364);
or U19768 (N_19768,N_19165,N_19452);
nor U19769 (N_19769,N_19265,N_19011);
xor U19770 (N_19770,N_19322,N_19119);
or U19771 (N_19771,N_19239,N_19260);
and U19772 (N_19772,N_19059,N_19323);
xor U19773 (N_19773,N_19071,N_19290);
xor U19774 (N_19774,N_19144,N_19042);
nor U19775 (N_19775,N_19234,N_19265);
nor U19776 (N_19776,N_19242,N_19303);
or U19777 (N_19777,N_19474,N_19110);
xnor U19778 (N_19778,N_19128,N_19367);
nand U19779 (N_19779,N_19397,N_19315);
nor U19780 (N_19780,N_19417,N_19267);
and U19781 (N_19781,N_19310,N_19459);
or U19782 (N_19782,N_19411,N_19452);
nor U19783 (N_19783,N_19158,N_19161);
or U19784 (N_19784,N_19221,N_19202);
nor U19785 (N_19785,N_19095,N_19365);
xor U19786 (N_19786,N_19129,N_19118);
or U19787 (N_19787,N_19284,N_19429);
xor U19788 (N_19788,N_19046,N_19175);
nor U19789 (N_19789,N_19340,N_19212);
nand U19790 (N_19790,N_19399,N_19233);
nor U19791 (N_19791,N_19268,N_19343);
or U19792 (N_19792,N_19046,N_19236);
and U19793 (N_19793,N_19175,N_19196);
nand U19794 (N_19794,N_19444,N_19263);
xnor U19795 (N_19795,N_19340,N_19057);
or U19796 (N_19796,N_19267,N_19358);
or U19797 (N_19797,N_19443,N_19276);
nor U19798 (N_19798,N_19469,N_19464);
or U19799 (N_19799,N_19223,N_19016);
nand U19800 (N_19800,N_19220,N_19126);
xnor U19801 (N_19801,N_19195,N_19064);
and U19802 (N_19802,N_19352,N_19341);
nand U19803 (N_19803,N_19360,N_19160);
nand U19804 (N_19804,N_19401,N_19072);
and U19805 (N_19805,N_19304,N_19274);
and U19806 (N_19806,N_19322,N_19404);
xnor U19807 (N_19807,N_19466,N_19015);
nor U19808 (N_19808,N_19197,N_19402);
xor U19809 (N_19809,N_19337,N_19175);
nand U19810 (N_19810,N_19486,N_19416);
or U19811 (N_19811,N_19354,N_19318);
nor U19812 (N_19812,N_19072,N_19271);
and U19813 (N_19813,N_19128,N_19382);
xnor U19814 (N_19814,N_19017,N_19102);
and U19815 (N_19815,N_19074,N_19242);
nand U19816 (N_19816,N_19272,N_19327);
and U19817 (N_19817,N_19407,N_19481);
or U19818 (N_19818,N_19312,N_19178);
nor U19819 (N_19819,N_19369,N_19370);
nand U19820 (N_19820,N_19090,N_19429);
and U19821 (N_19821,N_19384,N_19419);
or U19822 (N_19822,N_19367,N_19156);
nor U19823 (N_19823,N_19239,N_19217);
nand U19824 (N_19824,N_19244,N_19035);
xnor U19825 (N_19825,N_19268,N_19353);
xor U19826 (N_19826,N_19260,N_19315);
nor U19827 (N_19827,N_19469,N_19050);
or U19828 (N_19828,N_19339,N_19344);
xor U19829 (N_19829,N_19065,N_19198);
or U19830 (N_19830,N_19025,N_19219);
xnor U19831 (N_19831,N_19421,N_19376);
and U19832 (N_19832,N_19088,N_19293);
nand U19833 (N_19833,N_19374,N_19013);
nand U19834 (N_19834,N_19308,N_19343);
and U19835 (N_19835,N_19232,N_19356);
nand U19836 (N_19836,N_19128,N_19472);
nor U19837 (N_19837,N_19045,N_19030);
or U19838 (N_19838,N_19103,N_19307);
and U19839 (N_19839,N_19223,N_19297);
or U19840 (N_19840,N_19125,N_19355);
nor U19841 (N_19841,N_19249,N_19283);
and U19842 (N_19842,N_19392,N_19487);
nand U19843 (N_19843,N_19172,N_19335);
nor U19844 (N_19844,N_19035,N_19375);
or U19845 (N_19845,N_19183,N_19062);
and U19846 (N_19846,N_19302,N_19091);
or U19847 (N_19847,N_19147,N_19130);
or U19848 (N_19848,N_19414,N_19321);
xor U19849 (N_19849,N_19386,N_19459);
nand U19850 (N_19850,N_19040,N_19380);
or U19851 (N_19851,N_19375,N_19169);
nor U19852 (N_19852,N_19301,N_19360);
and U19853 (N_19853,N_19448,N_19290);
nand U19854 (N_19854,N_19389,N_19437);
xnor U19855 (N_19855,N_19190,N_19002);
xnor U19856 (N_19856,N_19495,N_19236);
and U19857 (N_19857,N_19230,N_19325);
and U19858 (N_19858,N_19062,N_19088);
nand U19859 (N_19859,N_19205,N_19252);
or U19860 (N_19860,N_19043,N_19307);
nand U19861 (N_19861,N_19473,N_19325);
or U19862 (N_19862,N_19165,N_19336);
xnor U19863 (N_19863,N_19250,N_19170);
nand U19864 (N_19864,N_19366,N_19349);
or U19865 (N_19865,N_19054,N_19085);
nor U19866 (N_19866,N_19365,N_19177);
or U19867 (N_19867,N_19008,N_19166);
nor U19868 (N_19868,N_19233,N_19117);
and U19869 (N_19869,N_19099,N_19326);
or U19870 (N_19870,N_19298,N_19312);
nand U19871 (N_19871,N_19387,N_19112);
nand U19872 (N_19872,N_19266,N_19400);
or U19873 (N_19873,N_19489,N_19376);
nor U19874 (N_19874,N_19138,N_19100);
or U19875 (N_19875,N_19433,N_19343);
and U19876 (N_19876,N_19144,N_19090);
nor U19877 (N_19877,N_19053,N_19437);
and U19878 (N_19878,N_19403,N_19069);
nand U19879 (N_19879,N_19080,N_19359);
nand U19880 (N_19880,N_19105,N_19259);
nor U19881 (N_19881,N_19199,N_19330);
or U19882 (N_19882,N_19073,N_19222);
or U19883 (N_19883,N_19163,N_19410);
nor U19884 (N_19884,N_19113,N_19228);
nand U19885 (N_19885,N_19421,N_19129);
and U19886 (N_19886,N_19143,N_19490);
xnor U19887 (N_19887,N_19383,N_19195);
nand U19888 (N_19888,N_19300,N_19250);
xor U19889 (N_19889,N_19179,N_19339);
nand U19890 (N_19890,N_19095,N_19192);
nor U19891 (N_19891,N_19296,N_19284);
or U19892 (N_19892,N_19009,N_19132);
nor U19893 (N_19893,N_19151,N_19122);
or U19894 (N_19894,N_19499,N_19251);
nand U19895 (N_19895,N_19262,N_19050);
nor U19896 (N_19896,N_19474,N_19126);
and U19897 (N_19897,N_19230,N_19429);
nand U19898 (N_19898,N_19408,N_19024);
nor U19899 (N_19899,N_19149,N_19361);
nand U19900 (N_19900,N_19032,N_19194);
nand U19901 (N_19901,N_19450,N_19058);
nor U19902 (N_19902,N_19361,N_19170);
xnor U19903 (N_19903,N_19331,N_19206);
and U19904 (N_19904,N_19109,N_19322);
xor U19905 (N_19905,N_19300,N_19063);
and U19906 (N_19906,N_19279,N_19261);
or U19907 (N_19907,N_19470,N_19447);
or U19908 (N_19908,N_19096,N_19358);
and U19909 (N_19909,N_19136,N_19173);
nand U19910 (N_19910,N_19284,N_19353);
nand U19911 (N_19911,N_19033,N_19002);
nand U19912 (N_19912,N_19111,N_19453);
and U19913 (N_19913,N_19179,N_19019);
and U19914 (N_19914,N_19292,N_19344);
and U19915 (N_19915,N_19199,N_19490);
or U19916 (N_19916,N_19287,N_19033);
nand U19917 (N_19917,N_19157,N_19117);
and U19918 (N_19918,N_19332,N_19189);
and U19919 (N_19919,N_19069,N_19355);
nand U19920 (N_19920,N_19217,N_19096);
nor U19921 (N_19921,N_19388,N_19203);
or U19922 (N_19922,N_19109,N_19449);
nand U19923 (N_19923,N_19477,N_19032);
and U19924 (N_19924,N_19039,N_19267);
nand U19925 (N_19925,N_19192,N_19001);
nand U19926 (N_19926,N_19123,N_19100);
nand U19927 (N_19927,N_19261,N_19108);
nor U19928 (N_19928,N_19322,N_19198);
and U19929 (N_19929,N_19445,N_19021);
or U19930 (N_19930,N_19369,N_19077);
or U19931 (N_19931,N_19046,N_19294);
nand U19932 (N_19932,N_19343,N_19312);
nor U19933 (N_19933,N_19364,N_19465);
nand U19934 (N_19934,N_19461,N_19204);
xnor U19935 (N_19935,N_19001,N_19079);
nand U19936 (N_19936,N_19246,N_19143);
nor U19937 (N_19937,N_19171,N_19179);
nand U19938 (N_19938,N_19091,N_19112);
xnor U19939 (N_19939,N_19192,N_19279);
nand U19940 (N_19940,N_19345,N_19061);
nor U19941 (N_19941,N_19004,N_19017);
xnor U19942 (N_19942,N_19033,N_19425);
and U19943 (N_19943,N_19098,N_19309);
nor U19944 (N_19944,N_19345,N_19388);
xor U19945 (N_19945,N_19469,N_19489);
nand U19946 (N_19946,N_19167,N_19366);
nor U19947 (N_19947,N_19185,N_19052);
nor U19948 (N_19948,N_19068,N_19021);
nand U19949 (N_19949,N_19017,N_19177);
xor U19950 (N_19950,N_19088,N_19105);
nor U19951 (N_19951,N_19001,N_19026);
xnor U19952 (N_19952,N_19149,N_19066);
nand U19953 (N_19953,N_19290,N_19020);
or U19954 (N_19954,N_19333,N_19205);
xnor U19955 (N_19955,N_19166,N_19186);
nand U19956 (N_19956,N_19486,N_19018);
and U19957 (N_19957,N_19032,N_19471);
nand U19958 (N_19958,N_19311,N_19262);
nand U19959 (N_19959,N_19404,N_19325);
nand U19960 (N_19960,N_19181,N_19213);
xor U19961 (N_19961,N_19275,N_19058);
or U19962 (N_19962,N_19419,N_19037);
nor U19963 (N_19963,N_19274,N_19473);
xor U19964 (N_19964,N_19004,N_19342);
and U19965 (N_19965,N_19129,N_19366);
nor U19966 (N_19966,N_19185,N_19337);
and U19967 (N_19967,N_19303,N_19407);
nand U19968 (N_19968,N_19335,N_19327);
nand U19969 (N_19969,N_19459,N_19456);
or U19970 (N_19970,N_19093,N_19026);
or U19971 (N_19971,N_19076,N_19075);
or U19972 (N_19972,N_19095,N_19190);
or U19973 (N_19973,N_19237,N_19196);
and U19974 (N_19974,N_19351,N_19055);
xor U19975 (N_19975,N_19170,N_19150);
and U19976 (N_19976,N_19437,N_19166);
nand U19977 (N_19977,N_19026,N_19410);
and U19978 (N_19978,N_19422,N_19220);
xnor U19979 (N_19979,N_19295,N_19328);
xor U19980 (N_19980,N_19059,N_19495);
nor U19981 (N_19981,N_19406,N_19316);
nor U19982 (N_19982,N_19266,N_19236);
and U19983 (N_19983,N_19171,N_19362);
nand U19984 (N_19984,N_19089,N_19207);
and U19985 (N_19985,N_19056,N_19451);
nor U19986 (N_19986,N_19425,N_19196);
nor U19987 (N_19987,N_19082,N_19063);
or U19988 (N_19988,N_19166,N_19176);
nor U19989 (N_19989,N_19058,N_19029);
or U19990 (N_19990,N_19322,N_19383);
or U19991 (N_19991,N_19499,N_19352);
and U19992 (N_19992,N_19108,N_19259);
or U19993 (N_19993,N_19117,N_19047);
nand U19994 (N_19994,N_19491,N_19194);
and U19995 (N_19995,N_19218,N_19093);
or U19996 (N_19996,N_19374,N_19426);
nor U19997 (N_19997,N_19107,N_19217);
xnor U19998 (N_19998,N_19231,N_19233);
nand U19999 (N_19999,N_19454,N_19396);
nor U20000 (N_20000,N_19736,N_19520);
and U20001 (N_20001,N_19578,N_19928);
xnor U20002 (N_20002,N_19511,N_19505);
nand U20003 (N_20003,N_19605,N_19715);
or U20004 (N_20004,N_19844,N_19757);
or U20005 (N_20005,N_19965,N_19506);
nand U20006 (N_20006,N_19557,N_19532);
or U20007 (N_20007,N_19921,N_19555);
xnor U20008 (N_20008,N_19608,N_19606);
nor U20009 (N_20009,N_19722,N_19577);
xor U20010 (N_20010,N_19961,N_19684);
and U20011 (N_20011,N_19912,N_19543);
or U20012 (N_20012,N_19616,N_19818);
and U20013 (N_20013,N_19907,N_19859);
or U20014 (N_20014,N_19647,N_19840);
and U20015 (N_20015,N_19937,N_19791);
xnor U20016 (N_20016,N_19966,N_19622);
nand U20017 (N_20017,N_19696,N_19995);
nor U20018 (N_20018,N_19914,N_19645);
xnor U20019 (N_20019,N_19801,N_19979);
and U20020 (N_20020,N_19533,N_19933);
or U20021 (N_20021,N_19565,N_19724);
nor U20022 (N_20022,N_19944,N_19864);
xor U20023 (N_20023,N_19703,N_19594);
xor U20024 (N_20024,N_19688,N_19666);
nor U20025 (N_20025,N_19895,N_19670);
and U20026 (N_20026,N_19737,N_19892);
or U20027 (N_20027,N_19519,N_19780);
xor U20028 (N_20028,N_19887,N_19627);
xnor U20029 (N_20029,N_19659,N_19985);
or U20030 (N_20030,N_19669,N_19925);
nor U20031 (N_20031,N_19819,N_19676);
or U20032 (N_20032,N_19509,N_19689);
or U20033 (N_20033,N_19711,N_19618);
xor U20034 (N_20034,N_19894,N_19850);
or U20035 (N_20035,N_19570,N_19752);
nor U20036 (N_20036,N_19805,N_19623);
nand U20037 (N_20037,N_19504,N_19759);
and U20038 (N_20038,N_19994,N_19528);
xor U20039 (N_20039,N_19651,N_19571);
and U20040 (N_20040,N_19734,N_19704);
xnor U20041 (N_20041,N_19663,N_19766);
nand U20042 (N_20042,N_19628,N_19513);
and U20043 (N_20043,N_19716,N_19603);
or U20044 (N_20044,N_19554,N_19807);
nand U20045 (N_20045,N_19640,N_19595);
nand U20046 (N_20046,N_19566,N_19839);
or U20047 (N_20047,N_19920,N_19542);
or U20048 (N_20048,N_19833,N_19707);
nor U20049 (N_20049,N_19799,N_19861);
and U20050 (N_20050,N_19870,N_19899);
and U20051 (N_20051,N_19888,N_19891);
nand U20052 (N_20052,N_19730,N_19910);
nand U20053 (N_20053,N_19815,N_19694);
xnor U20054 (N_20054,N_19817,N_19526);
nor U20055 (N_20055,N_19885,N_19916);
nand U20056 (N_20056,N_19770,N_19569);
and U20057 (N_20057,N_19990,N_19792);
or U20058 (N_20058,N_19869,N_19573);
xnor U20059 (N_20059,N_19556,N_19946);
and U20060 (N_20060,N_19638,N_19604);
nor U20061 (N_20061,N_19889,N_19681);
or U20062 (N_20062,N_19559,N_19539);
xor U20063 (N_20063,N_19738,N_19545);
or U20064 (N_20064,N_19584,N_19970);
nor U20065 (N_20065,N_19726,N_19596);
or U20066 (N_20066,N_19827,N_19739);
nand U20067 (N_20067,N_19846,N_19862);
and U20068 (N_20068,N_19612,N_19560);
nor U20069 (N_20069,N_19562,N_19636);
and U20070 (N_20070,N_19593,N_19834);
nor U20071 (N_20071,N_19968,N_19656);
xnor U20072 (N_20072,N_19664,N_19754);
nor U20073 (N_20073,N_19607,N_19789);
nand U20074 (N_20074,N_19989,N_19837);
nor U20075 (N_20075,N_19794,N_19587);
and U20076 (N_20076,N_19843,N_19976);
or U20077 (N_20077,N_19808,N_19691);
and U20078 (N_20078,N_19963,N_19880);
nor U20079 (N_20079,N_19810,N_19598);
nand U20080 (N_20080,N_19779,N_19948);
or U20081 (N_20081,N_19633,N_19708);
or U20082 (N_20082,N_19515,N_19508);
and U20083 (N_20083,N_19918,N_19875);
nand U20084 (N_20084,N_19929,N_19953);
or U20085 (N_20085,N_19854,N_19599);
or U20086 (N_20086,N_19547,N_19909);
nor U20087 (N_20087,N_19583,N_19753);
xor U20088 (N_20088,N_19853,N_19702);
or U20089 (N_20089,N_19855,N_19790);
or U20090 (N_20090,N_19732,N_19776);
and U20091 (N_20091,N_19580,N_19822);
nor U20092 (N_20092,N_19997,N_19709);
xor U20093 (N_20093,N_19958,N_19905);
nor U20094 (N_20094,N_19524,N_19969);
nor U20095 (N_20095,N_19553,N_19535);
or U20096 (N_20096,N_19728,N_19660);
and U20097 (N_20097,N_19574,N_19549);
or U20098 (N_20098,N_19922,N_19673);
and U20099 (N_20099,N_19537,N_19624);
xnor U20100 (N_20100,N_19959,N_19873);
and U20101 (N_20101,N_19802,N_19936);
or U20102 (N_20102,N_19939,N_19761);
or U20103 (N_20103,N_19522,N_19591);
xnor U20104 (N_20104,N_19783,N_19652);
nor U20105 (N_20105,N_19649,N_19646);
or U20106 (N_20106,N_19725,N_19956);
nor U20107 (N_20107,N_19534,N_19592);
nand U20108 (N_20108,N_19540,N_19886);
and U20109 (N_20109,N_19721,N_19809);
and U20110 (N_20110,N_19881,N_19816);
nand U20111 (N_20111,N_19654,N_19823);
and U20112 (N_20112,N_19723,N_19697);
or U20113 (N_20113,N_19575,N_19988);
or U20114 (N_20114,N_19778,N_19590);
nand U20115 (N_20115,N_19878,N_19617);
nand U20116 (N_20116,N_19782,N_19984);
and U20117 (N_20117,N_19576,N_19635);
nor U20118 (N_20118,N_19973,N_19619);
or U20119 (N_20119,N_19765,N_19686);
xnor U20120 (N_20120,N_19643,N_19856);
xor U20121 (N_20121,N_19804,N_19986);
and U20122 (N_20122,N_19865,N_19767);
or U20123 (N_20123,N_19814,N_19763);
nor U20124 (N_20124,N_19983,N_19964);
nand U20125 (N_20125,N_19831,N_19842);
and U20126 (N_20126,N_19629,N_19678);
and U20127 (N_20127,N_19991,N_19655);
nand U20128 (N_20128,N_19706,N_19877);
nand U20129 (N_20129,N_19650,N_19858);
and U20130 (N_20130,N_19719,N_19762);
nor U20131 (N_20131,N_19589,N_19981);
and U20132 (N_20132,N_19527,N_19987);
or U20133 (N_20133,N_19631,N_19733);
and U20134 (N_20134,N_19924,N_19741);
xnor U20135 (N_20135,N_19586,N_19897);
or U20136 (N_20136,N_19851,N_19915);
xnor U20137 (N_20137,N_19876,N_19942);
nand U20138 (N_20138,N_19551,N_19943);
nor U20139 (N_20139,N_19516,N_19582);
xnor U20140 (N_20140,N_19938,N_19755);
nand U20141 (N_20141,N_19552,N_19829);
xor U20142 (N_20142,N_19683,N_19777);
xor U20143 (N_20143,N_19567,N_19751);
nor U20144 (N_20144,N_19698,N_19685);
nor U20145 (N_20145,N_19680,N_19867);
nand U20146 (N_20146,N_19919,N_19525);
and U20147 (N_20147,N_19720,N_19917);
and U20148 (N_20148,N_19879,N_19625);
xor U20149 (N_20149,N_19501,N_19860);
nand U20150 (N_20150,N_19671,N_19731);
xnor U20151 (N_20151,N_19531,N_19771);
nor U20152 (N_20152,N_19695,N_19620);
and U20153 (N_20153,N_19967,N_19700);
xor U20154 (N_20154,N_19658,N_19800);
xnor U20155 (N_20155,N_19847,N_19538);
or U20156 (N_20156,N_19502,N_19911);
nor U20157 (N_20157,N_19940,N_19713);
and U20158 (N_20158,N_19871,N_19932);
nand U20159 (N_20159,N_19675,N_19714);
nand U20160 (N_20160,N_19821,N_19746);
nor U20161 (N_20161,N_19848,N_19903);
xor U20162 (N_20162,N_19896,N_19644);
or U20163 (N_20163,N_19507,N_19634);
nand U20164 (N_20164,N_19836,N_19518);
xor U20165 (N_20165,N_19826,N_19597);
nor U20166 (N_20166,N_19906,N_19908);
nor U20167 (N_20167,N_19977,N_19874);
or U20168 (N_20168,N_19744,N_19774);
nor U20169 (N_20169,N_19931,N_19529);
and U20170 (N_20170,N_19661,N_19665);
xor U20171 (N_20171,N_19996,N_19900);
and U20172 (N_20172,N_19639,N_19787);
xor U20173 (N_20173,N_19824,N_19945);
or U20174 (N_20174,N_19610,N_19747);
nand U20175 (N_20175,N_19949,N_19803);
and U20176 (N_20176,N_19841,N_19630);
nor U20177 (N_20177,N_19999,N_19668);
and U20178 (N_20178,N_19677,N_19784);
nor U20179 (N_20179,N_19868,N_19561);
xor U20180 (N_20180,N_19793,N_19530);
or U20181 (N_20181,N_19692,N_19934);
or U20182 (N_20182,N_19500,N_19712);
or U20183 (N_20183,N_19572,N_19884);
nor U20184 (N_20184,N_19813,N_19718);
nor U20185 (N_20185,N_19971,N_19993);
nand U20186 (N_20186,N_19514,N_19653);
nand U20187 (N_20187,N_19788,N_19611);
and U20188 (N_20188,N_19890,N_19563);
nand U20189 (N_20189,N_19954,N_19835);
nor U20190 (N_20190,N_19764,N_19972);
or U20191 (N_20191,N_19512,N_19564);
and U20192 (N_20192,N_19705,N_19693);
and U20193 (N_20193,N_19626,N_19773);
or U20194 (N_20194,N_19588,N_19998);
nand U20195 (N_20195,N_19935,N_19786);
nand U20196 (N_20196,N_19975,N_19541);
or U20197 (N_20197,N_19883,N_19690);
nand U20198 (N_20198,N_19710,N_19558);
nor U20199 (N_20199,N_19775,N_19717);
nor U20200 (N_20200,N_19830,N_19893);
or U20201 (N_20201,N_19863,N_19548);
nor U20202 (N_20202,N_19510,N_19760);
or U20203 (N_20203,N_19898,N_19820);
nor U20204 (N_20204,N_19632,N_19621);
nor U20205 (N_20205,N_19828,N_19769);
xor U20206 (N_20206,N_19796,N_19901);
nor U20207 (N_20207,N_19641,N_19952);
nor U20208 (N_20208,N_19679,N_19785);
xnor U20209 (N_20209,N_19648,N_19585);
xor U20210 (N_20210,N_19568,N_19682);
nand U20211 (N_20211,N_19749,N_19756);
nor U20212 (N_20212,N_19546,N_19735);
nor U20213 (N_20213,N_19904,N_19923);
and U20214 (N_20214,N_19951,N_19536);
and U20215 (N_20215,N_19615,N_19947);
xor U20216 (N_20216,N_19740,N_19849);
and U20217 (N_20217,N_19614,N_19978);
nor U20218 (N_20218,N_19642,N_19503);
and U20219 (N_20219,N_19613,N_19980);
and U20220 (N_20220,N_19550,N_19962);
xnor U20221 (N_20221,N_19930,N_19517);
or U20222 (N_20222,N_19806,N_19667);
nor U20223 (N_20223,N_19982,N_19795);
or U20224 (N_20224,N_19872,N_19637);
nand U20225 (N_20225,N_19974,N_19672);
or U20226 (N_20226,N_19882,N_19609);
and U20227 (N_20227,N_19742,N_19772);
and U20228 (N_20228,N_19866,N_19602);
nand U20229 (N_20229,N_19992,N_19927);
xnor U20230 (N_20230,N_19523,N_19674);
or U20231 (N_20231,N_19687,N_19600);
xnor U20232 (N_20232,N_19955,N_19902);
xor U20233 (N_20233,N_19950,N_19926);
and U20234 (N_20234,N_19812,N_19743);
xor U20235 (N_20235,N_19781,N_19913);
xor U20236 (N_20236,N_19662,N_19832);
nor U20237 (N_20237,N_19521,N_19579);
xor U20238 (N_20238,N_19941,N_19798);
xnor U20239 (N_20239,N_19758,N_19544);
xor U20240 (N_20240,N_19729,N_19581);
nor U20241 (N_20241,N_19960,N_19838);
xor U20242 (N_20242,N_19957,N_19852);
or U20243 (N_20243,N_19657,N_19701);
xor U20244 (N_20244,N_19825,N_19748);
nor U20245 (N_20245,N_19857,N_19745);
or U20246 (N_20246,N_19797,N_19811);
nor U20247 (N_20247,N_19601,N_19699);
nor U20248 (N_20248,N_19845,N_19750);
nand U20249 (N_20249,N_19727,N_19768);
xnor U20250 (N_20250,N_19877,N_19689);
and U20251 (N_20251,N_19819,N_19729);
nor U20252 (N_20252,N_19643,N_19605);
nor U20253 (N_20253,N_19906,N_19857);
xnor U20254 (N_20254,N_19528,N_19531);
or U20255 (N_20255,N_19644,N_19926);
nand U20256 (N_20256,N_19666,N_19533);
or U20257 (N_20257,N_19511,N_19733);
nor U20258 (N_20258,N_19667,N_19905);
and U20259 (N_20259,N_19741,N_19813);
nand U20260 (N_20260,N_19778,N_19962);
nor U20261 (N_20261,N_19529,N_19934);
xnor U20262 (N_20262,N_19950,N_19627);
nand U20263 (N_20263,N_19962,N_19708);
or U20264 (N_20264,N_19848,N_19532);
and U20265 (N_20265,N_19652,N_19560);
and U20266 (N_20266,N_19757,N_19808);
xnor U20267 (N_20267,N_19989,N_19541);
nor U20268 (N_20268,N_19803,N_19580);
nand U20269 (N_20269,N_19950,N_19555);
or U20270 (N_20270,N_19569,N_19960);
xor U20271 (N_20271,N_19605,N_19631);
nor U20272 (N_20272,N_19579,N_19897);
nor U20273 (N_20273,N_19820,N_19702);
nor U20274 (N_20274,N_19998,N_19808);
nor U20275 (N_20275,N_19945,N_19667);
and U20276 (N_20276,N_19889,N_19689);
nor U20277 (N_20277,N_19945,N_19628);
nand U20278 (N_20278,N_19730,N_19807);
and U20279 (N_20279,N_19615,N_19787);
and U20280 (N_20280,N_19884,N_19886);
nor U20281 (N_20281,N_19526,N_19771);
xnor U20282 (N_20282,N_19914,N_19898);
nor U20283 (N_20283,N_19794,N_19675);
and U20284 (N_20284,N_19508,N_19533);
and U20285 (N_20285,N_19583,N_19584);
nand U20286 (N_20286,N_19756,N_19507);
nor U20287 (N_20287,N_19961,N_19861);
xor U20288 (N_20288,N_19647,N_19763);
or U20289 (N_20289,N_19805,N_19853);
or U20290 (N_20290,N_19846,N_19705);
nor U20291 (N_20291,N_19662,N_19727);
nand U20292 (N_20292,N_19988,N_19500);
nand U20293 (N_20293,N_19662,N_19695);
xor U20294 (N_20294,N_19866,N_19517);
nor U20295 (N_20295,N_19804,N_19658);
or U20296 (N_20296,N_19543,N_19633);
or U20297 (N_20297,N_19528,N_19975);
nand U20298 (N_20298,N_19950,N_19530);
nor U20299 (N_20299,N_19806,N_19793);
nand U20300 (N_20300,N_19818,N_19995);
xor U20301 (N_20301,N_19808,N_19988);
nand U20302 (N_20302,N_19529,N_19835);
or U20303 (N_20303,N_19815,N_19877);
nor U20304 (N_20304,N_19736,N_19654);
and U20305 (N_20305,N_19592,N_19618);
and U20306 (N_20306,N_19620,N_19704);
xnor U20307 (N_20307,N_19530,N_19853);
xor U20308 (N_20308,N_19837,N_19727);
nand U20309 (N_20309,N_19597,N_19623);
xor U20310 (N_20310,N_19942,N_19967);
and U20311 (N_20311,N_19612,N_19533);
xnor U20312 (N_20312,N_19950,N_19664);
nand U20313 (N_20313,N_19874,N_19713);
nor U20314 (N_20314,N_19544,N_19915);
xor U20315 (N_20315,N_19527,N_19707);
nand U20316 (N_20316,N_19608,N_19780);
or U20317 (N_20317,N_19881,N_19776);
xnor U20318 (N_20318,N_19584,N_19742);
or U20319 (N_20319,N_19557,N_19764);
or U20320 (N_20320,N_19695,N_19505);
nor U20321 (N_20321,N_19666,N_19836);
or U20322 (N_20322,N_19508,N_19710);
nor U20323 (N_20323,N_19509,N_19893);
nor U20324 (N_20324,N_19686,N_19729);
or U20325 (N_20325,N_19938,N_19697);
xnor U20326 (N_20326,N_19842,N_19912);
and U20327 (N_20327,N_19768,N_19712);
nand U20328 (N_20328,N_19685,N_19967);
nor U20329 (N_20329,N_19911,N_19940);
nor U20330 (N_20330,N_19844,N_19920);
nor U20331 (N_20331,N_19838,N_19902);
or U20332 (N_20332,N_19739,N_19738);
nand U20333 (N_20333,N_19639,N_19885);
nor U20334 (N_20334,N_19817,N_19688);
xnor U20335 (N_20335,N_19959,N_19685);
nand U20336 (N_20336,N_19950,N_19684);
or U20337 (N_20337,N_19947,N_19742);
or U20338 (N_20338,N_19736,N_19507);
and U20339 (N_20339,N_19702,N_19600);
and U20340 (N_20340,N_19817,N_19785);
or U20341 (N_20341,N_19924,N_19691);
xnor U20342 (N_20342,N_19844,N_19805);
nand U20343 (N_20343,N_19813,N_19772);
and U20344 (N_20344,N_19990,N_19503);
nand U20345 (N_20345,N_19582,N_19703);
nor U20346 (N_20346,N_19970,N_19857);
nor U20347 (N_20347,N_19561,N_19726);
and U20348 (N_20348,N_19758,N_19941);
nor U20349 (N_20349,N_19987,N_19938);
nor U20350 (N_20350,N_19712,N_19986);
and U20351 (N_20351,N_19949,N_19636);
xnor U20352 (N_20352,N_19893,N_19673);
xor U20353 (N_20353,N_19616,N_19751);
xnor U20354 (N_20354,N_19748,N_19969);
or U20355 (N_20355,N_19665,N_19569);
nor U20356 (N_20356,N_19558,N_19863);
or U20357 (N_20357,N_19762,N_19863);
nand U20358 (N_20358,N_19703,N_19810);
nand U20359 (N_20359,N_19970,N_19601);
xor U20360 (N_20360,N_19790,N_19834);
and U20361 (N_20361,N_19645,N_19776);
nor U20362 (N_20362,N_19507,N_19920);
nor U20363 (N_20363,N_19866,N_19772);
or U20364 (N_20364,N_19613,N_19877);
nor U20365 (N_20365,N_19674,N_19591);
nor U20366 (N_20366,N_19859,N_19547);
and U20367 (N_20367,N_19554,N_19844);
xor U20368 (N_20368,N_19527,N_19563);
nor U20369 (N_20369,N_19501,N_19882);
xnor U20370 (N_20370,N_19721,N_19521);
and U20371 (N_20371,N_19954,N_19731);
or U20372 (N_20372,N_19804,N_19796);
and U20373 (N_20373,N_19685,N_19735);
nand U20374 (N_20374,N_19586,N_19528);
xor U20375 (N_20375,N_19533,N_19837);
nand U20376 (N_20376,N_19578,N_19748);
and U20377 (N_20377,N_19821,N_19573);
xnor U20378 (N_20378,N_19721,N_19766);
xor U20379 (N_20379,N_19972,N_19703);
or U20380 (N_20380,N_19897,N_19964);
or U20381 (N_20381,N_19510,N_19654);
xor U20382 (N_20382,N_19811,N_19834);
xnor U20383 (N_20383,N_19921,N_19653);
nand U20384 (N_20384,N_19704,N_19641);
and U20385 (N_20385,N_19711,N_19830);
xnor U20386 (N_20386,N_19987,N_19866);
nand U20387 (N_20387,N_19709,N_19771);
and U20388 (N_20388,N_19676,N_19773);
nand U20389 (N_20389,N_19642,N_19812);
and U20390 (N_20390,N_19520,N_19681);
nor U20391 (N_20391,N_19872,N_19629);
nor U20392 (N_20392,N_19876,N_19905);
xnor U20393 (N_20393,N_19682,N_19964);
or U20394 (N_20394,N_19698,N_19565);
and U20395 (N_20395,N_19717,N_19540);
xor U20396 (N_20396,N_19690,N_19586);
nor U20397 (N_20397,N_19763,N_19751);
nand U20398 (N_20398,N_19777,N_19989);
xnor U20399 (N_20399,N_19536,N_19910);
nor U20400 (N_20400,N_19916,N_19893);
nand U20401 (N_20401,N_19979,N_19737);
or U20402 (N_20402,N_19506,N_19580);
nand U20403 (N_20403,N_19817,N_19660);
and U20404 (N_20404,N_19821,N_19919);
nand U20405 (N_20405,N_19677,N_19653);
xor U20406 (N_20406,N_19584,N_19603);
xor U20407 (N_20407,N_19547,N_19602);
nor U20408 (N_20408,N_19784,N_19944);
xnor U20409 (N_20409,N_19823,N_19843);
xor U20410 (N_20410,N_19590,N_19544);
nor U20411 (N_20411,N_19984,N_19571);
and U20412 (N_20412,N_19892,N_19569);
nor U20413 (N_20413,N_19996,N_19530);
nand U20414 (N_20414,N_19955,N_19617);
and U20415 (N_20415,N_19939,N_19621);
nor U20416 (N_20416,N_19622,N_19808);
nor U20417 (N_20417,N_19816,N_19796);
xor U20418 (N_20418,N_19600,N_19947);
nor U20419 (N_20419,N_19958,N_19854);
or U20420 (N_20420,N_19776,N_19970);
nor U20421 (N_20421,N_19628,N_19621);
nor U20422 (N_20422,N_19680,N_19742);
xor U20423 (N_20423,N_19522,N_19579);
xor U20424 (N_20424,N_19704,N_19672);
or U20425 (N_20425,N_19832,N_19842);
and U20426 (N_20426,N_19907,N_19629);
or U20427 (N_20427,N_19942,N_19859);
xor U20428 (N_20428,N_19565,N_19546);
and U20429 (N_20429,N_19568,N_19641);
or U20430 (N_20430,N_19657,N_19524);
nor U20431 (N_20431,N_19619,N_19935);
and U20432 (N_20432,N_19623,N_19541);
and U20433 (N_20433,N_19893,N_19798);
or U20434 (N_20434,N_19797,N_19887);
nor U20435 (N_20435,N_19516,N_19653);
or U20436 (N_20436,N_19634,N_19774);
or U20437 (N_20437,N_19715,N_19836);
and U20438 (N_20438,N_19572,N_19909);
and U20439 (N_20439,N_19765,N_19700);
xor U20440 (N_20440,N_19576,N_19665);
xor U20441 (N_20441,N_19855,N_19803);
nand U20442 (N_20442,N_19523,N_19635);
nor U20443 (N_20443,N_19828,N_19837);
nand U20444 (N_20444,N_19769,N_19968);
nand U20445 (N_20445,N_19955,N_19590);
nor U20446 (N_20446,N_19559,N_19766);
nor U20447 (N_20447,N_19879,N_19906);
nor U20448 (N_20448,N_19710,N_19936);
and U20449 (N_20449,N_19983,N_19534);
xnor U20450 (N_20450,N_19789,N_19626);
nor U20451 (N_20451,N_19732,N_19728);
or U20452 (N_20452,N_19640,N_19581);
xnor U20453 (N_20453,N_19690,N_19603);
and U20454 (N_20454,N_19686,N_19531);
nand U20455 (N_20455,N_19850,N_19783);
and U20456 (N_20456,N_19774,N_19830);
and U20457 (N_20457,N_19893,N_19915);
nand U20458 (N_20458,N_19917,N_19708);
nor U20459 (N_20459,N_19857,N_19747);
or U20460 (N_20460,N_19955,N_19925);
and U20461 (N_20461,N_19691,N_19778);
or U20462 (N_20462,N_19989,N_19538);
and U20463 (N_20463,N_19620,N_19724);
nand U20464 (N_20464,N_19802,N_19699);
nor U20465 (N_20465,N_19693,N_19613);
xor U20466 (N_20466,N_19727,N_19950);
and U20467 (N_20467,N_19636,N_19885);
nor U20468 (N_20468,N_19678,N_19828);
nand U20469 (N_20469,N_19982,N_19552);
nor U20470 (N_20470,N_19901,N_19882);
and U20471 (N_20471,N_19760,N_19968);
nand U20472 (N_20472,N_19675,N_19896);
and U20473 (N_20473,N_19852,N_19759);
nor U20474 (N_20474,N_19526,N_19539);
nor U20475 (N_20475,N_19801,N_19864);
and U20476 (N_20476,N_19558,N_19719);
or U20477 (N_20477,N_19532,N_19906);
nor U20478 (N_20478,N_19664,N_19896);
and U20479 (N_20479,N_19884,N_19869);
nand U20480 (N_20480,N_19530,N_19887);
or U20481 (N_20481,N_19966,N_19687);
nand U20482 (N_20482,N_19883,N_19742);
nor U20483 (N_20483,N_19720,N_19669);
nor U20484 (N_20484,N_19617,N_19723);
nand U20485 (N_20485,N_19891,N_19827);
xnor U20486 (N_20486,N_19623,N_19844);
or U20487 (N_20487,N_19586,N_19543);
nand U20488 (N_20488,N_19559,N_19715);
or U20489 (N_20489,N_19965,N_19939);
xnor U20490 (N_20490,N_19837,N_19831);
xor U20491 (N_20491,N_19648,N_19759);
and U20492 (N_20492,N_19998,N_19981);
or U20493 (N_20493,N_19595,N_19864);
nor U20494 (N_20494,N_19804,N_19645);
or U20495 (N_20495,N_19674,N_19866);
nand U20496 (N_20496,N_19716,N_19900);
nand U20497 (N_20497,N_19624,N_19960);
xor U20498 (N_20498,N_19742,N_19892);
nor U20499 (N_20499,N_19750,N_19714);
nor U20500 (N_20500,N_20113,N_20188);
nor U20501 (N_20501,N_20258,N_20271);
or U20502 (N_20502,N_20210,N_20087);
nor U20503 (N_20503,N_20160,N_20240);
xor U20504 (N_20504,N_20373,N_20082);
nor U20505 (N_20505,N_20030,N_20083);
xor U20506 (N_20506,N_20004,N_20498);
nand U20507 (N_20507,N_20039,N_20261);
nand U20508 (N_20508,N_20419,N_20380);
nand U20509 (N_20509,N_20161,N_20178);
nand U20510 (N_20510,N_20095,N_20396);
and U20511 (N_20511,N_20464,N_20156);
nor U20512 (N_20512,N_20018,N_20260);
or U20513 (N_20513,N_20143,N_20385);
or U20514 (N_20514,N_20387,N_20356);
and U20515 (N_20515,N_20345,N_20237);
or U20516 (N_20516,N_20218,N_20448);
and U20517 (N_20517,N_20068,N_20036);
nand U20518 (N_20518,N_20140,N_20180);
xnor U20519 (N_20519,N_20475,N_20220);
nand U20520 (N_20520,N_20050,N_20031);
nor U20521 (N_20521,N_20395,N_20438);
nand U20522 (N_20522,N_20459,N_20032);
nand U20523 (N_20523,N_20442,N_20250);
or U20524 (N_20524,N_20219,N_20342);
xor U20525 (N_20525,N_20192,N_20348);
or U20526 (N_20526,N_20425,N_20055);
or U20527 (N_20527,N_20064,N_20299);
and U20528 (N_20528,N_20303,N_20381);
and U20529 (N_20529,N_20386,N_20462);
xnor U20530 (N_20530,N_20417,N_20231);
and U20531 (N_20531,N_20499,N_20114);
or U20532 (N_20532,N_20158,N_20024);
xnor U20533 (N_20533,N_20202,N_20277);
or U20534 (N_20534,N_20078,N_20027);
or U20535 (N_20535,N_20293,N_20135);
nand U20536 (N_20536,N_20089,N_20205);
and U20537 (N_20537,N_20097,N_20040);
nand U20538 (N_20538,N_20347,N_20067);
xor U20539 (N_20539,N_20301,N_20228);
nand U20540 (N_20540,N_20246,N_20094);
or U20541 (N_20541,N_20150,N_20165);
and U20542 (N_20542,N_20069,N_20129);
nand U20543 (N_20543,N_20447,N_20330);
and U20544 (N_20544,N_20080,N_20096);
xnor U20545 (N_20545,N_20035,N_20195);
or U20546 (N_20546,N_20247,N_20496);
xor U20547 (N_20547,N_20304,N_20355);
nor U20548 (N_20548,N_20422,N_20481);
nor U20549 (N_20549,N_20057,N_20189);
xnor U20550 (N_20550,N_20429,N_20492);
and U20551 (N_20551,N_20168,N_20051);
xor U20552 (N_20552,N_20077,N_20130);
xor U20553 (N_20553,N_20398,N_20430);
or U20554 (N_20554,N_20349,N_20333);
or U20555 (N_20555,N_20019,N_20213);
nand U20556 (N_20556,N_20029,N_20230);
nor U20557 (N_20557,N_20343,N_20361);
xnor U20558 (N_20558,N_20340,N_20073);
or U20559 (N_20559,N_20365,N_20369);
nor U20560 (N_20560,N_20206,N_20358);
or U20561 (N_20561,N_20233,N_20289);
xor U20562 (N_20562,N_20444,N_20245);
nor U20563 (N_20563,N_20125,N_20332);
nor U20564 (N_20564,N_20242,N_20460);
xnor U20565 (N_20565,N_20187,N_20106);
xnor U20566 (N_20566,N_20485,N_20063);
nand U20567 (N_20567,N_20001,N_20028);
and U20568 (N_20568,N_20312,N_20098);
xor U20569 (N_20569,N_20434,N_20015);
or U20570 (N_20570,N_20437,N_20414);
nand U20571 (N_20571,N_20043,N_20139);
xnor U20572 (N_20572,N_20486,N_20421);
xnor U20573 (N_20573,N_20463,N_20487);
nand U20574 (N_20574,N_20415,N_20477);
and U20575 (N_20575,N_20428,N_20453);
and U20576 (N_20576,N_20426,N_20391);
and U20577 (N_20577,N_20166,N_20173);
and U20578 (N_20578,N_20167,N_20127);
or U20579 (N_20579,N_20427,N_20059);
xor U20580 (N_20580,N_20257,N_20320);
xnor U20581 (N_20581,N_20280,N_20182);
xnor U20582 (N_20582,N_20283,N_20424);
xnor U20583 (N_20583,N_20270,N_20466);
nand U20584 (N_20584,N_20093,N_20132);
xor U20585 (N_20585,N_20164,N_20241);
nand U20586 (N_20586,N_20159,N_20013);
or U20587 (N_20587,N_20389,N_20351);
xor U20588 (N_20588,N_20134,N_20359);
and U20589 (N_20589,N_20222,N_20201);
or U20590 (N_20590,N_20234,N_20314);
nand U20591 (N_20591,N_20184,N_20402);
and U20592 (N_20592,N_20441,N_20163);
nand U20593 (N_20593,N_20061,N_20108);
nand U20594 (N_20594,N_20374,N_20384);
nand U20595 (N_20595,N_20149,N_20153);
or U20596 (N_20596,N_20144,N_20062);
nor U20597 (N_20597,N_20081,N_20232);
nand U20598 (N_20598,N_20099,N_20409);
nor U20599 (N_20599,N_20316,N_20190);
and U20600 (N_20600,N_20038,N_20196);
or U20601 (N_20601,N_20199,N_20243);
xnor U20602 (N_20602,N_20116,N_20104);
xnor U20603 (N_20603,N_20341,N_20394);
or U20604 (N_20604,N_20103,N_20070);
xor U20605 (N_20605,N_20305,N_20123);
xor U20606 (N_20606,N_20121,N_20450);
or U20607 (N_20607,N_20408,N_20091);
nand U20608 (N_20608,N_20334,N_20457);
or U20609 (N_20609,N_20468,N_20276);
nor U20610 (N_20610,N_20364,N_20439);
and U20611 (N_20611,N_20290,N_20480);
nand U20612 (N_20612,N_20319,N_20177);
nor U20613 (N_20613,N_20212,N_20399);
nor U20614 (N_20614,N_20251,N_20045);
nor U20615 (N_20615,N_20269,N_20294);
and U20616 (N_20616,N_20151,N_20327);
and U20617 (N_20617,N_20155,N_20357);
nor U20618 (N_20618,N_20313,N_20476);
nand U20619 (N_20619,N_20054,N_20344);
and U20620 (N_20620,N_20474,N_20109);
or U20621 (N_20621,N_20445,N_20090);
or U20622 (N_20622,N_20397,N_20076);
xnor U20623 (N_20623,N_20286,N_20420);
xor U20624 (N_20624,N_20092,N_20490);
or U20625 (N_20625,N_20413,N_20401);
xor U20626 (N_20626,N_20371,N_20204);
nor U20627 (N_20627,N_20047,N_20236);
xnor U20628 (N_20628,N_20449,N_20472);
xnor U20629 (N_20629,N_20221,N_20382);
or U20630 (N_20630,N_20010,N_20203);
nand U20631 (N_20631,N_20086,N_20009);
nor U20632 (N_20632,N_20186,N_20298);
xor U20633 (N_20633,N_20041,N_20454);
xor U20634 (N_20634,N_20238,N_20056);
nand U20635 (N_20635,N_20366,N_20388);
xnor U20636 (N_20636,N_20265,N_20405);
or U20637 (N_20637,N_20458,N_20052);
nor U20638 (N_20638,N_20363,N_20249);
and U20639 (N_20639,N_20263,N_20321);
nand U20640 (N_20640,N_20179,N_20211);
nor U20641 (N_20641,N_20208,N_20215);
and U20642 (N_20642,N_20488,N_20037);
and U20643 (N_20643,N_20049,N_20229);
xnor U20644 (N_20644,N_20217,N_20279);
nor U20645 (N_20645,N_20058,N_20295);
xor U20646 (N_20646,N_20372,N_20171);
and U20647 (N_20647,N_20074,N_20119);
or U20648 (N_20648,N_20354,N_20491);
nor U20649 (N_20649,N_20467,N_20138);
or U20650 (N_20650,N_20157,N_20141);
nand U20651 (N_20651,N_20446,N_20022);
or U20652 (N_20652,N_20350,N_20297);
or U20653 (N_20653,N_20335,N_20065);
and U20654 (N_20654,N_20193,N_20259);
nor U20655 (N_20655,N_20407,N_20310);
xor U20656 (N_20656,N_20469,N_20110);
and U20657 (N_20657,N_20336,N_20255);
xor U20658 (N_20658,N_20275,N_20390);
nand U20659 (N_20659,N_20185,N_20197);
xor U20660 (N_20660,N_20066,N_20432);
xor U20661 (N_20661,N_20044,N_20148);
nand U20662 (N_20662,N_20128,N_20003);
nor U20663 (N_20663,N_20346,N_20254);
or U20664 (N_20664,N_20273,N_20403);
and U20665 (N_20665,N_20465,N_20026);
or U20666 (N_20666,N_20470,N_20360);
xnor U20667 (N_20667,N_20456,N_20262);
and U20668 (N_20668,N_20007,N_20324);
and U20669 (N_20669,N_20183,N_20495);
nand U20670 (N_20670,N_20410,N_20025);
and U20671 (N_20671,N_20433,N_20112);
nor U20672 (N_20672,N_20226,N_20331);
and U20673 (N_20673,N_20473,N_20014);
or U20674 (N_20674,N_20147,N_20216);
and U20675 (N_20675,N_20315,N_20281);
nor U20676 (N_20676,N_20338,N_20339);
nor U20677 (N_20677,N_20431,N_20284);
or U20678 (N_20678,N_20017,N_20411);
nand U20679 (N_20679,N_20124,N_20483);
xor U20680 (N_20680,N_20300,N_20337);
and U20681 (N_20681,N_20383,N_20256);
nand U20682 (N_20682,N_20272,N_20367);
and U20683 (N_20683,N_20309,N_20227);
xnor U20684 (N_20684,N_20006,N_20489);
xnor U20685 (N_20685,N_20060,N_20072);
xor U20686 (N_20686,N_20033,N_20000);
nand U20687 (N_20687,N_20377,N_20461);
xor U20688 (N_20688,N_20322,N_20136);
and U20689 (N_20689,N_20170,N_20253);
nor U20690 (N_20690,N_20326,N_20034);
and U20691 (N_20691,N_20406,N_20176);
and U20692 (N_20692,N_20484,N_20362);
or U20693 (N_20693,N_20085,N_20478);
xor U20694 (N_20694,N_20002,N_20131);
nor U20695 (N_20695,N_20107,N_20115);
or U20696 (N_20696,N_20443,N_20207);
nor U20697 (N_20697,N_20235,N_20376);
xnor U20698 (N_20698,N_20042,N_20370);
xor U20699 (N_20699,N_20323,N_20102);
and U20700 (N_20700,N_20225,N_20393);
nor U20701 (N_20701,N_20021,N_20296);
xnor U20702 (N_20702,N_20325,N_20418);
and U20703 (N_20703,N_20046,N_20311);
nand U20704 (N_20704,N_20005,N_20088);
nor U20705 (N_20705,N_20306,N_20146);
or U20706 (N_20706,N_20126,N_20172);
xnor U20707 (N_20707,N_20169,N_20048);
and U20708 (N_20708,N_20142,N_20368);
or U20709 (N_20709,N_20302,N_20264);
nor U20710 (N_20710,N_20117,N_20266);
nor U20711 (N_20711,N_20137,N_20423);
and U20712 (N_20712,N_20194,N_20224);
nand U20713 (N_20713,N_20353,N_20400);
nand U20714 (N_20714,N_20223,N_20118);
and U20715 (N_20715,N_20120,N_20023);
xnor U20716 (N_20716,N_20452,N_20133);
nand U20717 (N_20717,N_20451,N_20282);
or U20718 (N_20718,N_20455,N_20267);
xor U20719 (N_20719,N_20174,N_20152);
nor U20720 (N_20720,N_20497,N_20436);
and U20721 (N_20721,N_20122,N_20175);
nor U20722 (N_20722,N_20317,N_20493);
and U20723 (N_20723,N_20214,N_20071);
nor U20724 (N_20724,N_20191,N_20111);
nand U20725 (N_20725,N_20318,N_20200);
or U20726 (N_20726,N_20209,N_20244);
nand U20727 (N_20727,N_20145,N_20412);
xnor U20728 (N_20728,N_20162,N_20239);
or U20729 (N_20729,N_20416,N_20011);
xor U20730 (N_20730,N_20375,N_20329);
and U20731 (N_20731,N_20328,N_20105);
nor U20732 (N_20732,N_20482,N_20079);
nor U20733 (N_20733,N_20435,N_20274);
and U20734 (N_20734,N_20252,N_20378);
nand U20735 (N_20735,N_20154,N_20292);
xor U20736 (N_20736,N_20101,N_20404);
nor U20737 (N_20737,N_20198,N_20288);
nand U20738 (N_20738,N_20287,N_20352);
nor U20739 (N_20739,N_20100,N_20392);
or U20740 (N_20740,N_20084,N_20053);
and U20741 (N_20741,N_20278,N_20075);
and U20742 (N_20742,N_20285,N_20268);
xor U20743 (N_20743,N_20479,N_20008);
or U20744 (N_20744,N_20020,N_20379);
nor U20745 (N_20745,N_20471,N_20181);
nand U20746 (N_20746,N_20291,N_20440);
or U20747 (N_20747,N_20248,N_20494);
or U20748 (N_20748,N_20307,N_20308);
nor U20749 (N_20749,N_20016,N_20012);
and U20750 (N_20750,N_20327,N_20298);
and U20751 (N_20751,N_20028,N_20380);
or U20752 (N_20752,N_20062,N_20032);
nand U20753 (N_20753,N_20263,N_20204);
or U20754 (N_20754,N_20029,N_20074);
or U20755 (N_20755,N_20235,N_20284);
nor U20756 (N_20756,N_20066,N_20103);
or U20757 (N_20757,N_20419,N_20040);
or U20758 (N_20758,N_20411,N_20275);
xor U20759 (N_20759,N_20035,N_20138);
nor U20760 (N_20760,N_20463,N_20430);
and U20761 (N_20761,N_20249,N_20220);
or U20762 (N_20762,N_20405,N_20166);
xor U20763 (N_20763,N_20162,N_20003);
and U20764 (N_20764,N_20100,N_20418);
or U20765 (N_20765,N_20100,N_20197);
and U20766 (N_20766,N_20492,N_20091);
and U20767 (N_20767,N_20297,N_20443);
xnor U20768 (N_20768,N_20378,N_20279);
nor U20769 (N_20769,N_20033,N_20293);
and U20770 (N_20770,N_20100,N_20428);
xnor U20771 (N_20771,N_20317,N_20222);
nand U20772 (N_20772,N_20296,N_20090);
xor U20773 (N_20773,N_20327,N_20107);
and U20774 (N_20774,N_20242,N_20255);
xnor U20775 (N_20775,N_20195,N_20280);
xnor U20776 (N_20776,N_20429,N_20312);
xor U20777 (N_20777,N_20153,N_20399);
nand U20778 (N_20778,N_20318,N_20454);
and U20779 (N_20779,N_20284,N_20361);
xnor U20780 (N_20780,N_20228,N_20132);
xor U20781 (N_20781,N_20396,N_20137);
and U20782 (N_20782,N_20000,N_20340);
or U20783 (N_20783,N_20179,N_20162);
nor U20784 (N_20784,N_20381,N_20435);
nand U20785 (N_20785,N_20120,N_20264);
nand U20786 (N_20786,N_20445,N_20043);
nand U20787 (N_20787,N_20483,N_20294);
xnor U20788 (N_20788,N_20452,N_20454);
or U20789 (N_20789,N_20415,N_20183);
nor U20790 (N_20790,N_20148,N_20314);
and U20791 (N_20791,N_20295,N_20065);
or U20792 (N_20792,N_20304,N_20290);
xor U20793 (N_20793,N_20314,N_20343);
and U20794 (N_20794,N_20050,N_20039);
xor U20795 (N_20795,N_20262,N_20290);
or U20796 (N_20796,N_20258,N_20354);
xor U20797 (N_20797,N_20471,N_20022);
and U20798 (N_20798,N_20129,N_20392);
or U20799 (N_20799,N_20087,N_20176);
nand U20800 (N_20800,N_20153,N_20368);
and U20801 (N_20801,N_20355,N_20092);
nor U20802 (N_20802,N_20388,N_20429);
nand U20803 (N_20803,N_20096,N_20365);
or U20804 (N_20804,N_20131,N_20273);
nor U20805 (N_20805,N_20312,N_20277);
nand U20806 (N_20806,N_20320,N_20217);
xor U20807 (N_20807,N_20117,N_20222);
and U20808 (N_20808,N_20468,N_20040);
nor U20809 (N_20809,N_20414,N_20245);
nand U20810 (N_20810,N_20273,N_20113);
nor U20811 (N_20811,N_20454,N_20334);
nor U20812 (N_20812,N_20230,N_20158);
xnor U20813 (N_20813,N_20266,N_20278);
nand U20814 (N_20814,N_20164,N_20016);
and U20815 (N_20815,N_20332,N_20282);
or U20816 (N_20816,N_20390,N_20139);
nor U20817 (N_20817,N_20000,N_20167);
and U20818 (N_20818,N_20354,N_20140);
nor U20819 (N_20819,N_20180,N_20069);
or U20820 (N_20820,N_20061,N_20361);
and U20821 (N_20821,N_20244,N_20173);
xor U20822 (N_20822,N_20159,N_20045);
or U20823 (N_20823,N_20050,N_20030);
or U20824 (N_20824,N_20092,N_20427);
nor U20825 (N_20825,N_20203,N_20069);
nor U20826 (N_20826,N_20343,N_20396);
or U20827 (N_20827,N_20039,N_20211);
nand U20828 (N_20828,N_20291,N_20254);
and U20829 (N_20829,N_20157,N_20497);
or U20830 (N_20830,N_20498,N_20347);
nor U20831 (N_20831,N_20073,N_20039);
and U20832 (N_20832,N_20101,N_20238);
nor U20833 (N_20833,N_20399,N_20309);
or U20834 (N_20834,N_20305,N_20154);
nor U20835 (N_20835,N_20092,N_20005);
nor U20836 (N_20836,N_20477,N_20468);
nor U20837 (N_20837,N_20120,N_20421);
nand U20838 (N_20838,N_20408,N_20038);
and U20839 (N_20839,N_20171,N_20217);
or U20840 (N_20840,N_20177,N_20463);
nand U20841 (N_20841,N_20390,N_20300);
nor U20842 (N_20842,N_20173,N_20414);
xnor U20843 (N_20843,N_20493,N_20159);
nor U20844 (N_20844,N_20004,N_20294);
nor U20845 (N_20845,N_20031,N_20049);
nor U20846 (N_20846,N_20386,N_20392);
nor U20847 (N_20847,N_20493,N_20110);
or U20848 (N_20848,N_20417,N_20333);
nor U20849 (N_20849,N_20271,N_20224);
xnor U20850 (N_20850,N_20319,N_20215);
nor U20851 (N_20851,N_20421,N_20143);
nand U20852 (N_20852,N_20247,N_20022);
and U20853 (N_20853,N_20178,N_20231);
nor U20854 (N_20854,N_20149,N_20035);
and U20855 (N_20855,N_20170,N_20230);
nand U20856 (N_20856,N_20313,N_20368);
and U20857 (N_20857,N_20102,N_20125);
xor U20858 (N_20858,N_20030,N_20146);
and U20859 (N_20859,N_20499,N_20034);
nand U20860 (N_20860,N_20075,N_20294);
xor U20861 (N_20861,N_20499,N_20270);
or U20862 (N_20862,N_20235,N_20181);
and U20863 (N_20863,N_20495,N_20213);
xor U20864 (N_20864,N_20037,N_20118);
or U20865 (N_20865,N_20094,N_20035);
and U20866 (N_20866,N_20132,N_20074);
or U20867 (N_20867,N_20035,N_20307);
nor U20868 (N_20868,N_20431,N_20263);
nor U20869 (N_20869,N_20404,N_20288);
or U20870 (N_20870,N_20403,N_20155);
or U20871 (N_20871,N_20134,N_20146);
and U20872 (N_20872,N_20194,N_20416);
xnor U20873 (N_20873,N_20407,N_20441);
and U20874 (N_20874,N_20370,N_20399);
nand U20875 (N_20875,N_20272,N_20043);
and U20876 (N_20876,N_20423,N_20357);
and U20877 (N_20877,N_20078,N_20095);
or U20878 (N_20878,N_20329,N_20155);
nor U20879 (N_20879,N_20410,N_20462);
nand U20880 (N_20880,N_20177,N_20196);
or U20881 (N_20881,N_20147,N_20231);
or U20882 (N_20882,N_20046,N_20200);
nand U20883 (N_20883,N_20005,N_20449);
xor U20884 (N_20884,N_20198,N_20390);
or U20885 (N_20885,N_20161,N_20374);
nor U20886 (N_20886,N_20468,N_20222);
nor U20887 (N_20887,N_20131,N_20078);
or U20888 (N_20888,N_20496,N_20245);
and U20889 (N_20889,N_20390,N_20057);
xor U20890 (N_20890,N_20147,N_20022);
nor U20891 (N_20891,N_20277,N_20093);
xor U20892 (N_20892,N_20407,N_20228);
or U20893 (N_20893,N_20380,N_20094);
and U20894 (N_20894,N_20467,N_20341);
xnor U20895 (N_20895,N_20057,N_20295);
nand U20896 (N_20896,N_20210,N_20113);
xor U20897 (N_20897,N_20182,N_20164);
nand U20898 (N_20898,N_20198,N_20182);
or U20899 (N_20899,N_20416,N_20130);
and U20900 (N_20900,N_20007,N_20328);
xnor U20901 (N_20901,N_20178,N_20453);
nand U20902 (N_20902,N_20022,N_20391);
or U20903 (N_20903,N_20067,N_20394);
nor U20904 (N_20904,N_20210,N_20364);
xor U20905 (N_20905,N_20476,N_20082);
xnor U20906 (N_20906,N_20096,N_20122);
nor U20907 (N_20907,N_20245,N_20111);
and U20908 (N_20908,N_20277,N_20192);
and U20909 (N_20909,N_20468,N_20249);
or U20910 (N_20910,N_20232,N_20472);
or U20911 (N_20911,N_20178,N_20333);
and U20912 (N_20912,N_20382,N_20400);
and U20913 (N_20913,N_20369,N_20080);
and U20914 (N_20914,N_20034,N_20001);
nand U20915 (N_20915,N_20300,N_20401);
and U20916 (N_20916,N_20147,N_20127);
and U20917 (N_20917,N_20185,N_20436);
xnor U20918 (N_20918,N_20255,N_20246);
nor U20919 (N_20919,N_20013,N_20279);
nor U20920 (N_20920,N_20174,N_20148);
xnor U20921 (N_20921,N_20005,N_20464);
xor U20922 (N_20922,N_20003,N_20287);
nand U20923 (N_20923,N_20453,N_20104);
nand U20924 (N_20924,N_20120,N_20407);
nand U20925 (N_20925,N_20229,N_20286);
xor U20926 (N_20926,N_20344,N_20215);
xnor U20927 (N_20927,N_20374,N_20286);
nand U20928 (N_20928,N_20481,N_20204);
xnor U20929 (N_20929,N_20421,N_20407);
or U20930 (N_20930,N_20152,N_20234);
and U20931 (N_20931,N_20222,N_20028);
nor U20932 (N_20932,N_20476,N_20163);
nor U20933 (N_20933,N_20247,N_20374);
or U20934 (N_20934,N_20279,N_20169);
and U20935 (N_20935,N_20472,N_20421);
and U20936 (N_20936,N_20305,N_20244);
or U20937 (N_20937,N_20242,N_20381);
nor U20938 (N_20938,N_20410,N_20238);
and U20939 (N_20939,N_20467,N_20111);
xnor U20940 (N_20940,N_20235,N_20436);
nand U20941 (N_20941,N_20205,N_20023);
or U20942 (N_20942,N_20023,N_20377);
or U20943 (N_20943,N_20078,N_20349);
nor U20944 (N_20944,N_20476,N_20087);
or U20945 (N_20945,N_20353,N_20025);
xor U20946 (N_20946,N_20403,N_20186);
and U20947 (N_20947,N_20169,N_20168);
xor U20948 (N_20948,N_20243,N_20201);
and U20949 (N_20949,N_20026,N_20350);
nor U20950 (N_20950,N_20289,N_20439);
nand U20951 (N_20951,N_20426,N_20192);
xnor U20952 (N_20952,N_20252,N_20057);
nand U20953 (N_20953,N_20166,N_20048);
nor U20954 (N_20954,N_20424,N_20022);
nand U20955 (N_20955,N_20026,N_20191);
nor U20956 (N_20956,N_20078,N_20480);
nor U20957 (N_20957,N_20168,N_20133);
nand U20958 (N_20958,N_20188,N_20152);
xnor U20959 (N_20959,N_20213,N_20438);
xor U20960 (N_20960,N_20392,N_20384);
xor U20961 (N_20961,N_20379,N_20384);
and U20962 (N_20962,N_20177,N_20261);
and U20963 (N_20963,N_20154,N_20229);
and U20964 (N_20964,N_20378,N_20147);
or U20965 (N_20965,N_20495,N_20098);
nor U20966 (N_20966,N_20479,N_20123);
nor U20967 (N_20967,N_20384,N_20033);
or U20968 (N_20968,N_20410,N_20358);
or U20969 (N_20969,N_20445,N_20153);
and U20970 (N_20970,N_20238,N_20165);
or U20971 (N_20971,N_20194,N_20388);
or U20972 (N_20972,N_20345,N_20413);
or U20973 (N_20973,N_20249,N_20050);
or U20974 (N_20974,N_20149,N_20257);
or U20975 (N_20975,N_20256,N_20138);
and U20976 (N_20976,N_20222,N_20121);
nor U20977 (N_20977,N_20476,N_20055);
and U20978 (N_20978,N_20174,N_20036);
nor U20979 (N_20979,N_20263,N_20158);
nor U20980 (N_20980,N_20025,N_20307);
nand U20981 (N_20981,N_20341,N_20015);
or U20982 (N_20982,N_20111,N_20434);
xor U20983 (N_20983,N_20133,N_20296);
or U20984 (N_20984,N_20479,N_20167);
xor U20985 (N_20985,N_20205,N_20210);
nand U20986 (N_20986,N_20002,N_20012);
or U20987 (N_20987,N_20009,N_20328);
xor U20988 (N_20988,N_20166,N_20392);
nor U20989 (N_20989,N_20142,N_20249);
nand U20990 (N_20990,N_20277,N_20261);
nor U20991 (N_20991,N_20069,N_20350);
xnor U20992 (N_20992,N_20228,N_20253);
and U20993 (N_20993,N_20447,N_20155);
nand U20994 (N_20994,N_20001,N_20355);
nand U20995 (N_20995,N_20043,N_20251);
nor U20996 (N_20996,N_20220,N_20311);
nor U20997 (N_20997,N_20169,N_20260);
and U20998 (N_20998,N_20075,N_20025);
nand U20999 (N_20999,N_20407,N_20232);
nand U21000 (N_21000,N_20956,N_20914);
or U21001 (N_21001,N_20942,N_20553);
or U21002 (N_21002,N_20945,N_20814);
xnor U21003 (N_21003,N_20534,N_20824);
and U21004 (N_21004,N_20744,N_20665);
nand U21005 (N_21005,N_20782,N_20677);
and U21006 (N_21006,N_20607,N_20793);
nand U21007 (N_21007,N_20909,N_20660);
and U21008 (N_21008,N_20523,N_20880);
and U21009 (N_21009,N_20687,N_20969);
nor U21010 (N_21010,N_20784,N_20825);
xnor U21011 (N_21011,N_20542,N_20941);
and U21012 (N_21012,N_20767,N_20890);
and U21013 (N_21013,N_20990,N_20549);
nand U21014 (N_21014,N_20540,N_20512);
and U21015 (N_21015,N_20902,N_20551);
and U21016 (N_21016,N_20577,N_20883);
nand U21017 (N_21017,N_20723,N_20895);
xor U21018 (N_21018,N_20800,N_20799);
xor U21019 (N_21019,N_20650,N_20694);
xor U21020 (N_21020,N_20507,N_20750);
and U21021 (N_21021,N_20718,N_20834);
nand U21022 (N_21022,N_20501,N_20541);
nand U21023 (N_21023,N_20866,N_20773);
or U21024 (N_21024,N_20778,N_20755);
xnor U21025 (N_21025,N_20746,N_20869);
and U21026 (N_21026,N_20823,N_20878);
nand U21027 (N_21027,N_20719,N_20545);
or U21028 (N_21028,N_20818,N_20528);
nand U21029 (N_21029,N_20735,N_20884);
and U21030 (N_21030,N_20522,N_20612);
xnor U21031 (N_21031,N_20882,N_20666);
and U21032 (N_21032,N_20768,N_20554);
and U21033 (N_21033,N_20770,N_20872);
nor U21034 (N_21034,N_20525,N_20937);
and U21035 (N_21035,N_20916,N_20819);
and U21036 (N_21036,N_20751,N_20888);
and U21037 (N_21037,N_20864,N_20550);
nor U21038 (N_21038,N_20568,N_20785);
nand U21039 (N_21039,N_20691,N_20900);
nor U21040 (N_21040,N_20739,N_20935);
nand U21041 (N_21041,N_20924,N_20874);
nand U21042 (N_21042,N_20727,N_20989);
or U21043 (N_21043,N_20926,N_20981);
nor U21044 (N_21044,N_20961,N_20983);
and U21045 (N_21045,N_20844,N_20645);
xnor U21046 (N_21046,N_20986,N_20901);
xor U21047 (N_21047,N_20630,N_20529);
nand U21048 (N_21048,N_20663,N_20736);
and U21049 (N_21049,N_20609,N_20920);
xnor U21050 (N_21050,N_20829,N_20594);
xnor U21051 (N_21051,N_20646,N_20603);
and U21052 (N_21052,N_20991,N_20688);
nor U21053 (N_21053,N_20859,N_20978);
xor U21054 (N_21054,N_20759,N_20711);
and U21055 (N_21055,N_20740,N_20985);
xnor U21056 (N_21056,N_20537,N_20947);
xnor U21057 (N_21057,N_20634,N_20641);
nor U21058 (N_21058,N_20939,N_20669);
and U21059 (N_21059,N_20912,N_20514);
and U21060 (N_21060,N_20838,N_20976);
nor U21061 (N_21061,N_20801,N_20911);
nand U21062 (N_21062,N_20854,N_20853);
and U21063 (N_21063,N_20629,N_20552);
xnor U21064 (N_21064,N_20720,N_20959);
nand U21065 (N_21065,N_20997,N_20724);
and U21066 (N_21066,N_20597,N_20813);
nand U21067 (N_21067,N_20865,N_20973);
or U21068 (N_21068,N_20531,N_20567);
and U21069 (N_21069,N_20970,N_20995);
or U21070 (N_21070,N_20810,N_20886);
and U21071 (N_21071,N_20993,N_20876);
or U21072 (N_21072,N_20671,N_20557);
and U21073 (N_21073,N_20692,N_20667);
or U21074 (N_21074,N_20615,N_20606);
or U21075 (N_21075,N_20526,N_20563);
xor U21076 (N_21076,N_20836,N_20530);
or U21077 (N_21077,N_20828,N_20925);
or U21078 (N_21078,N_20946,N_20633);
or U21079 (N_21079,N_20599,N_20808);
nand U21080 (N_21080,N_20710,N_20915);
nor U21081 (N_21081,N_20849,N_20613);
and U21082 (N_21082,N_20678,N_20602);
nand U21083 (N_21083,N_20572,N_20658);
nor U21084 (N_21084,N_20732,N_20717);
xor U21085 (N_21085,N_20611,N_20538);
and U21086 (N_21086,N_20581,N_20835);
and U21087 (N_21087,N_20972,N_20675);
and U21088 (N_21088,N_20753,N_20802);
or U21089 (N_21089,N_20579,N_20730);
xor U21090 (N_21090,N_20757,N_20521);
nand U21091 (N_21091,N_20620,N_20680);
nand U21092 (N_21092,N_20604,N_20682);
nor U21093 (N_21093,N_20776,N_20566);
nor U21094 (N_21094,N_20845,N_20578);
xnor U21095 (N_21095,N_20725,N_20932);
nand U21096 (N_21096,N_20737,N_20811);
or U21097 (N_21097,N_20816,N_20875);
nor U21098 (N_21098,N_20940,N_20592);
xor U21099 (N_21099,N_20714,N_20949);
nor U21100 (N_21100,N_20651,N_20787);
and U21101 (N_21101,N_20994,N_20846);
xnor U21102 (N_21102,N_20928,N_20574);
nor U21103 (N_21103,N_20575,N_20943);
or U21104 (N_21104,N_20795,N_20786);
and U21105 (N_21105,N_20765,N_20860);
xnor U21106 (N_21106,N_20975,N_20952);
xnor U21107 (N_21107,N_20798,N_20504);
xnor U21108 (N_21108,N_20857,N_20547);
nor U21109 (N_21109,N_20841,N_20631);
xor U21110 (N_21110,N_20520,N_20833);
nand U21111 (N_21111,N_20571,N_20506);
or U21112 (N_21112,N_20964,N_20585);
xnor U21113 (N_21113,N_20674,N_20618);
nand U21114 (N_21114,N_20546,N_20950);
nand U21115 (N_21115,N_20992,N_20861);
nor U21116 (N_21116,N_20622,N_20556);
or U21117 (N_21117,N_20754,N_20636);
xnor U21118 (N_21118,N_20870,N_20511);
nor U21119 (N_21119,N_20683,N_20930);
or U21120 (N_21120,N_20858,N_20502);
xor U21121 (N_21121,N_20938,N_20974);
and U21122 (N_21122,N_20790,N_20748);
and U21123 (N_21123,N_20806,N_20764);
xnor U21124 (N_21124,N_20623,N_20960);
nand U21125 (N_21125,N_20643,N_20593);
or U21126 (N_21126,N_20536,N_20804);
nor U21127 (N_21127,N_20758,N_20713);
and U21128 (N_21128,N_20769,N_20519);
and U21129 (N_21129,N_20805,N_20684);
xnor U21130 (N_21130,N_20703,N_20771);
xor U21131 (N_21131,N_20923,N_20967);
nor U21132 (N_21132,N_20905,N_20681);
nand U21133 (N_21133,N_20775,N_20624);
or U21134 (N_21134,N_20569,N_20716);
or U21135 (N_21135,N_20591,N_20918);
xor U21136 (N_21136,N_20570,N_20999);
xor U21137 (N_21137,N_20722,N_20826);
nor U21138 (N_21138,N_20936,N_20689);
or U21139 (N_21139,N_20982,N_20850);
or U21140 (N_21140,N_20792,N_20686);
nand U21141 (N_21141,N_20893,N_20543);
nor U21142 (N_21142,N_20517,N_20933);
and U21143 (N_21143,N_20873,N_20596);
nand U21144 (N_21144,N_20852,N_20913);
or U21145 (N_21145,N_20734,N_20505);
xnor U21146 (N_21146,N_20867,N_20702);
nor U21147 (N_21147,N_20774,N_20639);
nand U21148 (N_21148,N_20934,N_20837);
nand U21149 (N_21149,N_20695,N_20555);
and U21150 (N_21150,N_20662,N_20701);
nor U21151 (N_21151,N_20715,N_20621);
and U21152 (N_21152,N_20743,N_20668);
nor U21153 (N_21153,N_20707,N_20598);
and U21154 (N_21154,N_20820,N_20610);
xor U21155 (N_21155,N_20708,N_20733);
nor U21156 (N_21156,N_20963,N_20752);
and U21157 (N_21157,N_20693,N_20697);
or U21158 (N_21158,N_20560,N_20712);
nor U21159 (N_21159,N_20919,N_20608);
xor U21160 (N_21160,N_20863,N_20562);
nor U21161 (N_21161,N_20679,N_20855);
and U21162 (N_21162,N_20781,N_20500);
xor U21163 (N_21163,N_20847,N_20565);
or U21164 (N_21164,N_20627,N_20524);
and U21165 (N_21165,N_20640,N_20953);
xnor U21166 (N_21166,N_20894,N_20605);
nand U21167 (N_21167,N_20513,N_20929);
nor U21168 (N_21168,N_20908,N_20616);
nand U21169 (N_21169,N_20601,N_20851);
or U21170 (N_21170,N_20791,N_20588);
xor U21171 (N_21171,N_20772,N_20644);
or U21172 (N_21172,N_20661,N_20968);
or U21173 (N_21173,N_20656,N_20654);
nand U21174 (N_21174,N_20921,N_20797);
nor U21175 (N_21175,N_20544,N_20922);
or U21176 (N_21176,N_20831,N_20822);
nand U21177 (N_21177,N_20780,N_20626);
nor U21178 (N_21178,N_20580,N_20700);
xnor U21179 (N_21179,N_20906,N_20971);
or U21180 (N_21180,N_20955,N_20887);
nor U21181 (N_21181,N_20762,N_20659);
and U21182 (N_21182,N_20706,N_20788);
or U21183 (N_21183,N_20817,N_20516);
xor U21184 (N_21184,N_20564,N_20761);
xor U21185 (N_21185,N_20948,N_20696);
and U21186 (N_21186,N_20510,N_20527);
xnor U21187 (N_21187,N_20614,N_20548);
and U21188 (N_21188,N_20907,N_20903);
nor U21189 (N_21189,N_20904,N_20879);
nand U21190 (N_21190,N_20533,N_20862);
or U21191 (N_21191,N_20595,N_20877);
nor U21192 (N_21192,N_20657,N_20789);
xor U21193 (N_21193,N_20515,N_20897);
xnor U21194 (N_21194,N_20632,N_20655);
or U21195 (N_21195,N_20705,N_20741);
xor U21196 (N_21196,N_20619,N_20582);
nand U21197 (N_21197,N_20889,N_20891);
or U21198 (N_21198,N_20649,N_20518);
or U21199 (N_21199,N_20996,N_20868);
or U21200 (N_21200,N_20709,N_20951);
xor U21201 (N_21201,N_20910,N_20638);
nor U21202 (N_21202,N_20881,N_20600);
xor U21203 (N_21203,N_20721,N_20962);
nand U21204 (N_21204,N_20728,N_20742);
or U21205 (N_21205,N_20535,N_20731);
nor U21206 (N_21206,N_20830,N_20508);
or U21207 (N_21207,N_20803,N_20763);
or U21208 (N_21208,N_20954,N_20815);
and U21209 (N_21209,N_20573,N_20977);
or U21210 (N_21210,N_20998,N_20625);
or U21211 (N_21211,N_20589,N_20503);
and U21212 (N_21212,N_20783,N_20617);
nor U21213 (N_21213,N_20777,N_20747);
and U21214 (N_21214,N_20749,N_20637);
or U21215 (N_21215,N_20979,N_20840);
and U21216 (N_21216,N_20704,N_20885);
or U21217 (N_21217,N_20647,N_20583);
nand U21218 (N_21218,N_20726,N_20584);
xnor U21219 (N_21219,N_20539,N_20871);
or U21220 (N_21220,N_20685,N_20586);
nand U21221 (N_21221,N_20832,N_20738);
or U21222 (N_21222,N_20756,N_20842);
and U21223 (N_21223,N_20690,N_20558);
xor U21224 (N_21224,N_20965,N_20984);
xnor U21225 (N_21225,N_20559,N_20896);
nor U21226 (N_21226,N_20848,N_20821);
xnor U21227 (N_21227,N_20899,N_20729);
nor U21228 (N_21228,N_20779,N_20794);
or U21229 (N_21229,N_20587,N_20898);
and U21230 (N_21230,N_20927,N_20839);
and U21231 (N_21231,N_20628,N_20698);
xor U21232 (N_21232,N_20699,N_20673);
xor U21233 (N_21233,N_20532,N_20635);
nand U21234 (N_21234,N_20760,N_20648);
or U21235 (N_21235,N_20796,N_20980);
nor U21236 (N_21236,N_20988,N_20944);
or U21237 (N_21237,N_20652,N_20590);
and U21238 (N_21238,N_20827,N_20561);
xor U21239 (N_21239,N_20766,N_20812);
and U21240 (N_21240,N_20672,N_20807);
or U21241 (N_21241,N_20670,N_20676);
xor U21242 (N_21242,N_20664,N_20653);
xor U21243 (N_21243,N_20576,N_20957);
xnor U21244 (N_21244,N_20931,N_20987);
nand U21245 (N_21245,N_20892,N_20958);
xnor U21246 (N_21246,N_20809,N_20509);
or U21247 (N_21247,N_20642,N_20917);
or U21248 (N_21248,N_20745,N_20843);
or U21249 (N_21249,N_20856,N_20966);
or U21250 (N_21250,N_20969,N_20610);
or U21251 (N_21251,N_20794,N_20853);
xnor U21252 (N_21252,N_20851,N_20748);
or U21253 (N_21253,N_20973,N_20792);
and U21254 (N_21254,N_20970,N_20597);
xor U21255 (N_21255,N_20597,N_20609);
nand U21256 (N_21256,N_20852,N_20597);
xor U21257 (N_21257,N_20761,N_20914);
nand U21258 (N_21258,N_20660,N_20646);
xnor U21259 (N_21259,N_20535,N_20645);
or U21260 (N_21260,N_20724,N_20825);
xor U21261 (N_21261,N_20756,N_20522);
or U21262 (N_21262,N_20813,N_20677);
and U21263 (N_21263,N_20768,N_20953);
or U21264 (N_21264,N_20514,N_20783);
xor U21265 (N_21265,N_20755,N_20641);
or U21266 (N_21266,N_20683,N_20622);
or U21267 (N_21267,N_20769,N_20610);
xor U21268 (N_21268,N_20954,N_20532);
xor U21269 (N_21269,N_20620,N_20794);
nor U21270 (N_21270,N_20907,N_20866);
nand U21271 (N_21271,N_20788,N_20987);
and U21272 (N_21272,N_20813,N_20957);
nand U21273 (N_21273,N_20562,N_20592);
xnor U21274 (N_21274,N_20828,N_20998);
xnor U21275 (N_21275,N_20571,N_20808);
xnor U21276 (N_21276,N_20539,N_20624);
and U21277 (N_21277,N_20702,N_20743);
xor U21278 (N_21278,N_20978,N_20998);
or U21279 (N_21279,N_20586,N_20800);
and U21280 (N_21280,N_20949,N_20718);
xnor U21281 (N_21281,N_20794,N_20542);
nand U21282 (N_21282,N_20918,N_20869);
nor U21283 (N_21283,N_20940,N_20521);
nor U21284 (N_21284,N_20924,N_20970);
xor U21285 (N_21285,N_20744,N_20750);
and U21286 (N_21286,N_20760,N_20999);
and U21287 (N_21287,N_20814,N_20993);
and U21288 (N_21288,N_20561,N_20828);
nand U21289 (N_21289,N_20921,N_20869);
nor U21290 (N_21290,N_20956,N_20612);
xnor U21291 (N_21291,N_20732,N_20606);
or U21292 (N_21292,N_20979,N_20678);
nor U21293 (N_21293,N_20663,N_20588);
nand U21294 (N_21294,N_20509,N_20862);
nor U21295 (N_21295,N_20596,N_20503);
and U21296 (N_21296,N_20953,N_20923);
nand U21297 (N_21297,N_20675,N_20745);
or U21298 (N_21298,N_20907,N_20794);
xor U21299 (N_21299,N_20886,N_20763);
nor U21300 (N_21300,N_20628,N_20965);
nor U21301 (N_21301,N_20843,N_20580);
or U21302 (N_21302,N_20787,N_20918);
xor U21303 (N_21303,N_20551,N_20959);
or U21304 (N_21304,N_20982,N_20845);
nor U21305 (N_21305,N_20597,N_20591);
xor U21306 (N_21306,N_20750,N_20753);
xor U21307 (N_21307,N_20815,N_20531);
or U21308 (N_21308,N_20906,N_20782);
nand U21309 (N_21309,N_20661,N_20659);
nand U21310 (N_21310,N_20825,N_20792);
xnor U21311 (N_21311,N_20666,N_20699);
nor U21312 (N_21312,N_20965,N_20662);
nor U21313 (N_21313,N_20873,N_20597);
xnor U21314 (N_21314,N_20898,N_20828);
and U21315 (N_21315,N_20876,N_20619);
xnor U21316 (N_21316,N_20538,N_20737);
nor U21317 (N_21317,N_20546,N_20866);
xnor U21318 (N_21318,N_20937,N_20691);
or U21319 (N_21319,N_20708,N_20953);
and U21320 (N_21320,N_20937,N_20882);
nor U21321 (N_21321,N_20534,N_20996);
xor U21322 (N_21322,N_20909,N_20630);
and U21323 (N_21323,N_20910,N_20593);
nand U21324 (N_21324,N_20960,N_20711);
nor U21325 (N_21325,N_20665,N_20628);
nand U21326 (N_21326,N_20959,N_20934);
xnor U21327 (N_21327,N_20931,N_20643);
nand U21328 (N_21328,N_20909,N_20904);
nor U21329 (N_21329,N_20626,N_20852);
nand U21330 (N_21330,N_20834,N_20880);
or U21331 (N_21331,N_20552,N_20711);
and U21332 (N_21332,N_20524,N_20535);
nand U21333 (N_21333,N_20621,N_20702);
nor U21334 (N_21334,N_20904,N_20882);
or U21335 (N_21335,N_20862,N_20947);
and U21336 (N_21336,N_20583,N_20562);
xor U21337 (N_21337,N_20925,N_20617);
xor U21338 (N_21338,N_20555,N_20822);
or U21339 (N_21339,N_20604,N_20571);
xnor U21340 (N_21340,N_20594,N_20947);
or U21341 (N_21341,N_20836,N_20534);
nor U21342 (N_21342,N_20941,N_20994);
or U21343 (N_21343,N_20903,N_20613);
and U21344 (N_21344,N_20582,N_20947);
or U21345 (N_21345,N_20660,N_20612);
or U21346 (N_21346,N_20986,N_20807);
and U21347 (N_21347,N_20666,N_20607);
nor U21348 (N_21348,N_20871,N_20508);
nor U21349 (N_21349,N_20549,N_20951);
xor U21350 (N_21350,N_20582,N_20745);
nor U21351 (N_21351,N_20801,N_20864);
nor U21352 (N_21352,N_20940,N_20522);
and U21353 (N_21353,N_20699,N_20710);
nand U21354 (N_21354,N_20899,N_20717);
or U21355 (N_21355,N_20706,N_20669);
nand U21356 (N_21356,N_20560,N_20825);
xor U21357 (N_21357,N_20561,N_20720);
or U21358 (N_21358,N_20514,N_20680);
xnor U21359 (N_21359,N_20782,N_20644);
xor U21360 (N_21360,N_20872,N_20737);
or U21361 (N_21361,N_20724,N_20779);
xnor U21362 (N_21362,N_20654,N_20734);
nand U21363 (N_21363,N_20928,N_20701);
xor U21364 (N_21364,N_20840,N_20880);
nand U21365 (N_21365,N_20654,N_20964);
nor U21366 (N_21366,N_20897,N_20872);
nand U21367 (N_21367,N_20825,N_20631);
and U21368 (N_21368,N_20749,N_20512);
nand U21369 (N_21369,N_20794,N_20511);
xor U21370 (N_21370,N_20697,N_20645);
nor U21371 (N_21371,N_20600,N_20929);
xor U21372 (N_21372,N_20611,N_20671);
and U21373 (N_21373,N_20891,N_20573);
nand U21374 (N_21374,N_20978,N_20882);
nand U21375 (N_21375,N_20506,N_20589);
or U21376 (N_21376,N_20563,N_20776);
or U21377 (N_21377,N_20888,N_20574);
xor U21378 (N_21378,N_20659,N_20741);
xor U21379 (N_21379,N_20578,N_20635);
and U21380 (N_21380,N_20832,N_20577);
nand U21381 (N_21381,N_20566,N_20786);
nand U21382 (N_21382,N_20907,N_20708);
nand U21383 (N_21383,N_20933,N_20869);
xnor U21384 (N_21384,N_20645,N_20815);
or U21385 (N_21385,N_20540,N_20666);
nand U21386 (N_21386,N_20922,N_20652);
nand U21387 (N_21387,N_20734,N_20708);
nand U21388 (N_21388,N_20562,N_20801);
or U21389 (N_21389,N_20874,N_20960);
nand U21390 (N_21390,N_20612,N_20741);
or U21391 (N_21391,N_20736,N_20807);
nand U21392 (N_21392,N_20607,N_20631);
nor U21393 (N_21393,N_20950,N_20562);
nand U21394 (N_21394,N_20528,N_20681);
nor U21395 (N_21395,N_20706,N_20757);
and U21396 (N_21396,N_20919,N_20968);
or U21397 (N_21397,N_20956,N_20508);
xnor U21398 (N_21398,N_20843,N_20800);
and U21399 (N_21399,N_20903,N_20906);
or U21400 (N_21400,N_20982,N_20943);
and U21401 (N_21401,N_20603,N_20892);
and U21402 (N_21402,N_20863,N_20518);
nand U21403 (N_21403,N_20704,N_20807);
nand U21404 (N_21404,N_20928,N_20923);
and U21405 (N_21405,N_20681,N_20546);
nor U21406 (N_21406,N_20824,N_20749);
nand U21407 (N_21407,N_20695,N_20751);
xor U21408 (N_21408,N_20799,N_20673);
and U21409 (N_21409,N_20603,N_20705);
xnor U21410 (N_21410,N_20676,N_20722);
and U21411 (N_21411,N_20690,N_20588);
xnor U21412 (N_21412,N_20893,N_20870);
or U21413 (N_21413,N_20508,N_20971);
nand U21414 (N_21414,N_20566,N_20783);
nor U21415 (N_21415,N_20720,N_20635);
xnor U21416 (N_21416,N_20586,N_20596);
or U21417 (N_21417,N_20718,N_20532);
or U21418 (N_21418,N_20849,N_20877);
nor U21419 (N_21419,N_20725,N_20513);
or U21420 (N_21420,N_20877,N_20605);
xnor U21421 (N_21421,N_20779,N_20950);
or U21422 (N_21422,N_20762,N_20917);
nor U21423 (N_21423,N_20969,N_20758);
or U21424 (N_21424,N_20675,N_20637);
nor U21425 (N_21425,N_20814,N_20870);
xnor U21426 (N_21426,N_20841,N_20880);
nand U21427 (N_21427,N_20754,N_20881);
and U21428 (N_21428,N_20584,N_20994);
nor U21429 (N_21429,N_20574,N_20973);
or U21430 (N_21430,N_20838,N_20500);
nor U21431 (N_21431,N_20929,N_20940);
nand U21432 (N_21432,N_20765,N_20682);
nand U21433 (N_21433,N_20952,N_20728);
or U21434 (N_21434,N_20719,N_20875);
or U21435 (N_21435,N_20995,N_20738);
xnor U21436 (N_21436,N_20726,N_20602);
nor U21437 (N_21437,N_20815,N_20561);
nand U21438 (N_21438,N_20932,N_20615);
nand U21439 (N_21439,N_20666,N_20614);
and U21440 (N_21440,N_20647,N_20635);
nor U21441 (N_21441,N_20565,N_20603);
xor U21442 (N_21442,N_20948,N_20655);
xor U21443 (N_21443,N_20902,N_20897);
or U21444 (N_21444,N_20718,N_20798);
nand U21445 (N_21445,N_20926,N_20849);
or U21446 (N_21446,N_20955,N_20681);
nor U21447 (N_21447,N_20652,N_20924);
nor U21448 (N_21448,N_20777,N_20768);
xnor U21449 (N_21449,N_20840,N_20667);
or U21450 (N_21450,N_20866,N_20650);
nor U21451 (N_21451,N_20651,N_20752);
and U21452 (N_21452,N_20648,N_20946);
or U21453 (N_21453,N_20592,N_20661);
nor U21454 (N_21454,N_20616,N_20943);
and U21455 (N_21455,N_20742,N_20700);
and U21456 (N_21456,N_20969,N_20993);
xor U21457 (N_21457,N_20583,N_20792);
nand U21458 (N_21458,N_20623,N_20535);
and U21459 (N_21459,N_20783,N_20572);
or U21460 (N_21460,N_20976,N_20734);
nand U21461 (N_21461,N_20896,N_20748);
or U21462 (N_21462,N_20629,N_20648);
or U21463 (N_21463,N_20514,N_20867);
nand U21464 (N_21464,N_20805,N_20733);
nand U21465 (N_21465,N_20944,N_20641);
nor U21466 (N_21466,N_20776,N_20890);
nand U21467 (N_21467,N_20771,N_20637);
xnor U21468 (N_21468,N_20789,N_20711);
or U21469 (N_21469,N_20855,N_20649);
nand U21470 (N_21470,N_20715,N_20661);
xor U21471 (N_21471,N_20817,N_20921);
nor U21472 (N_21472,N_20528,N_20548);
or U21473 (N_21473,N_20831,N_20998);
nand U21474 (N_21474,N_20967,N_20570);
or U21475 (N_21475,N_20520,N_20921);
xnor U21476 (N_21476,N_20865,N_20998);
or U21477 (N_21477,N_20985,N_20504);
and U21478 (N_21478,N_20584,N_20791);
and U21479 (N_21479,N_20658,N_20873);
and U21480 (N_21480,N_20758,N_20737);
nor U21481 (N_21481,N_20601,N_20679);
nand U21482 (N_21482,N_20976,N_20779);
and U21483 (N_21483,N_20736,N_20835);
xnor U21484 (N_21484,N_20848,N_20646);
xor U21485 (N_21485,N_20568,N_20942);
and U21486 (N_21486,N_20999,N_20715);
nor U21487 (N_21487,N_20816,N_20839);
and U21488 (N_21488,N_20615,N_20899);
nand U21489 (N_21489,N_20963,N_20797);
and U21490 (N_21490,N_20760,N_20969);
nand U21491 (N_21491,N_20640,N_20831);
and U21492 (N_21492,N_20551,N_20937);
and U21493 (N_21493,N_20946,N_20699);
nand U21494 (N_21494,N_20891,N_20947);
and U21495 (N_21495,N_20982,N_20966);
and U21496 (N_21496,N_20735,N_20893);
xnor U21497 (N_21497,N_20762,N_20529);
xor U21498 (N_21498,N_20598,N_20653);
and U21499 (N_21499,N_20681,N_20527);
xor U21500 (N_21500,N_21267,N_21378);
xor U21501 (N_21501,N_21051,N_21295);
xor U21502 (N_21502,N_21494,N_21213);
and U21503 (N_21503,N_21036,N_21177);
nand U21504 (N_21504,N_21286,N_21194);
and U21505 (N_21505,N_21081,N_21485);
and U21506 (N_21506,N_21143,N_21134);
xor U21507 (N_21507,N_21262,N_21329);
and U21508 (N_21508,N_21006,N_21482);
and U21509 (N_21509,N_21359,N_21137);
or U21510 (N_21510,N_21303,N_21129);
nor U21511 (N_21511,N_21476,N_21342);
or U21512 (N_21512,N_21061,N_21164);
nor U21513 (N_21513,N_21448,N_21268);
xor U21514 (N_21514,N_21108,N_21018);
and U21515 (N_21515,N_21096,N_21106);
and U21516 (N_21516,N_21073,N_21151);
and U21517 (N_21517,N_21016,N_21305);
or U21518 (N_21518,N_21150,N_21351);
or U21519 (N_21519,N_21462,N_21477);
nor U21520 (N_21520,N_21426,N_21316);
and U21521 (N_21521,N_21092,N_21178);
xor U21522 (N_21522,N_21419,N_21408);
nand U21523 (N_21523,N_21389,N_21029);
or U21524 (N_21524,N_21290,N_21079);
or U21525 (N_21525,N_21373,N_21019);
nor U21526 (N_21526,N_21376,N_21261);
nor U21527 (N_21527,N_21112,N_21043);
xor U21528 (N_21528,N_21272,N_21049);
or U21529 (N_21529,N_21350,N_21001);
nor U21530 (N_21530,N_21105,N_21269);
xnor U21531 (N_21531,N_21136,N_21153);
nor U21532 (N_21532,N_21443,N_21495);
nor U21533 (N_21533,N_21384,N_21201);
xor U21534 (N_21534,N_21028,N_21420);
and U21535 (N_21535,N_21364,N_21457);
xnor U21536 (N_21536,N_21042,N_21460);
or U21537 (N_21537,N_21375,N_21124);
nand U21538 (N_21538,N_21149,N_21089);
nor U21539 (N_21539,N_21047,N_21370);
nor U21540 (N_21540,N_21025,N_21191);
nand U21541 (N_21541,N_21343,N_21474);
and U21542 (N_21542,N_21117,N_21155);
or U21543 (N_21543,N_21087,N_21287);
and U21544 (N_21544,N_21398,N_21406);
nor U21545 (N_21545,N_21205,N_21352);
nor U21546 (N_21546,N_21496,N_21162);
or U21547 (N_21547,N_21392,N_21035);
or U21548 (N_21548,N_21447,N_21312);
xnor U21549 (N_21549,N_21218,N_21413);
nand U21550 (N_21550,N_21078,N_21257);
or U21551 (N_21551,N_21169,N_21004);
nand U21552 (N_21552,N_21363,N_21015);
nand U21553 (N_21553,N_21390,N_21196);
xor U21554 (N_21554,N_21265,N_21439);
nor U21555 (N_21555,N_21119,N_21291);
and U21556 (N_21556,N_21057,N_21469);
or U21557 (N_21557,N_21454,N_21031);
nand U21558 (N_21558,N_21338,N_21039);
nor U21559 (N_21559,N_21012,N_21479);
nand U21560 (N_21560,N_21297,N_21311);
and U21561 (N_21561,N_21000,N_21484);
xor U21562 (N_21562,N_21386,N_21279);
or U21563 (N_21563,N_21103,N_21217);
nor U21564 (N_21564,N_21030,N_21052);
nor U21565 (N_21565,N_21102,N_21385);
or U21566 (N_21566,N_21266,N_21409);
or U21567 (N_21567,N_21307,N_21491);
nand U21568 (N_21568,N_21422,N_21412);
xnor U21569 (N_21569,N_21308,N_21202);
nand U21570 (N_21570,N_21161,N_21046);
nor U21571 (N_21571,N_21063,N_21333);
nor U21572 (N_21572,N_21327,N_21365);
xor U21573 (N_21573,N_21313,N_21034);
nand U21574 (N_21574,N_21349,N_21487);
or U21575 (N_21575,N_21104,N_21499);
nand U21576 (N_21576,N_21374,N_21240);
or U21577 (N_21577,N_21357,N_21256);
and U21578 (N_21578,N_21423,N_21187);
or U21579 (N_21579,N_21247,N_21284);
and U21580 (N_21580,N_21315,N_21038);
nand U21581 (N_21581,N_21174,N_21172);
nor U21582 (N_21582,N_21442,N_21417);
or U21583 (N_21583,N_21190,N_21159);
or U21584 (N_21584,N_21416,N_21395);
nor U21585 (N_21585,N_21055,N_21361);
and U21586 (N_21586,N_21465,N_21271);
nor U21587 (N_21587,N_21399,N_21347);
and U21588 (N_21588,N_21253,N_21192);
nand U21589 (N_21589,N_21339,N_21074);
xnor U21590 (N_21590,N_21017,N_21450);
nor U21591 (N_21591,N_21014,N_21090);
and U21592 (N_21592,N_21110,N_21148);
nand U21593 (N_21593,N_21387,N_21180);
nor U21594 (N_21594,N_21170,N_21072);
xor U21595 (N_21595,N_21360,N_21250);
nor U21596 (N_21596,N_21324,N_21430);
and U21597 (N_21597,N_21421,N_21139);
nand U21598 (N_21598,N_21372,N_21446);
xor U21599 (N_21599,N_21002,N_21126);
xnor U21600 (N_21600,N_21223,N_21152);
xnor U21601 (N_21601,N_21381,N_21344);
or U21602 (N_21602,N_21280,N_21277);
nor U21603 (N_21603,N_21182,N_21093);
or U21604 (N_21604,N_21492,N_21179);
or U21605 (N_21605,N_21122,N_21157);
or U21606 (N_21606,N_21032,N_21466);
or U21607 (N_21607,N_21451,N_21237);
and U21608 (N_21608,N_21227,N_21383);
and U21609 (N_21609,N_21310,N_21296);
or U21610 (N_21610,N_21220,N_21239);
and U21611 (N_21611,N_21070,N_21082);
nand U21612 (N_21612,N_21397,N_21435);
or U21613 (N_21613,N_21197,N_21255);
nor U21614 (N_21614,N_21044,N_21130);
nand U21615 (N_21615,N_21283,N_21299);
nor U21616 (N_21616,N_21405,N_21473);
nand U21617 (N_21617,N_21175,N_21438);
or U21618 (N_21618,N_21084,N_21478);
and U21619 (N_21619,N_21185,N_21125);
nor U21620 (N_21620,N_21432,N_21234);
nor U21621 (N_21621,N_21254,N_21418);
or U21622 (N_21622,N_21354,N_21285);
xor U21623 (N_21623,N_21011,N_21453);
or U21624 (N_21624,N_21123,N_21188);
xnor U21625 (N_21625,N_21212,N_21075);
nor U21626 (N_21626,N_21210,N_21068);
xor U21627 (N_21627,N_21238,N_21449);
xnor U21628 (N_21628,N_21216,N_21245);
nor U21629 (N_21629,N_21366,N_21230);
or U21630 (N_21630,N_21132,N_21281);
nor U21631 (N_21631,N_21241,N_21160);
or U21632 (N_21632,N_21027,N_21244);
nor U21633 (N_21633,N_21204,N_21067);
nor U21634 (N_21634,N_21024,N_21135);
or U21635 (N_21635,N_21226,N_21353);
nand U21636 (N_21636,N_21401,N_21101);
and U21637 (N_21637,N_21293,N_21382);
nand U21638 (N_21638,N_21400,N_21058);
and U21639 (N_21639,N_21071,N_21128);
nor U21640 (N_21640,N_21222,N_21133);
nand U21641 (N_21641,N_21207,N_21320);
and U21642 (N_21642,N_21113,N_21048);
nor U21643 (N_21643,N_21371,N_21193);
nor U21644 (N_21644,N_21424,N_21183);
and U21645 (N_21645,N_21322,N_21379);
nor U21646 (N_21646,N_21270,N_21471);
nand U21647 (N_21647,N_21472,N_21037);
xnor U21648 (N_21648,N_21041,N_21340);
nor U21649 (N_21649,N_21116,N_21414);
nand U21650 (N_21650,N_21236,N_21452);
or U21651 (N_21651,N_21489,N_21437);
or U21652 (N_21652,N_21273,N_21211);
xnor U21653 (N_21653,N_21053,N_21358);
or U21654 (N_21654,N_21334,N_21208);
or U21655 (N_21655,N_21294,N_21186);
nand U21656 (N_21656,N_21224,N_21062);
xor U21657 (N_21657,N_21242,N_21335);
nor U21658 (N_21658,N_21306,N_21114);
or U21659 (N_21659,N_21225,N_21168);
or U21660 (N_21660,N_21121,N_21428);
or U21661 (N_21661,N_21147,N_21402);
or U21662 (N_21662,N_21411,N_21325);
and U21663 (N_21663,N_21083,N_21377);
nor U21664 (N_21664,N_21431,N_21127);
nor U21665 (N_21665,N_21263,N_21059);
nand U21666 (N_21666,N_21429,N_21198);
xnor U21667 (N_21667,N_21498,N_21336);
nand U21668 (N_21668,N_21301,N_21171);
nand U21669 (N_21669,N_21369,N_21380);
nor U21670 (N_21670,N_21203,N_21445);
nor U21671 (N_21671,N_21156,N_21138);
and U21672 (N_21672,N_21362,N_21278);
and U21673 (N_21673,N_21050,N_21154);
xor U21674 (N_21674,N_21463,N_21199);
nor U21675 (N_21675,N_21109,N_21013);
and U21676 (N_21676,N_21060,N_21323);
nand U21677 (N_21677,N_21056,N_21480);
nand U21678 (N_21678,N_21464,N_21142);
xnor U21679 (N_21679,N_21228,N_21022);
or U21680 (N_21680,N_21348,N_21302);
xnor U21681 (N_21681,N_21209,N_21167);
or U21682 (N_21682,N_21097,N_21440);
and U21683 (N_21683,N_21094,N_21003);
nor U21684 (N_21684,N_21131,N_21243);
xor U21685 (N_21685,N_21140,N_21163);
nand U21686 (N_21686,N_21231,N_21020);
nor U21687 (N_21687,N_21355,N_21189);
nand U21688 (N_21688,N_21066,N_21248);
nor U21689 (N_21689,N_21252,N_21118);
nand U21690 (N_21690,N_21337,N_21076);
xor U21691 (N_21691,N_21318,N_21077);
and U21692 (N_21692,N_21393,N_21332);
xor U21693 (N_21693,N_21314,N_21069);
xor U21694 (N_21694,N_21095,N_21394);
xor U21695 (N_21695,N_21493,N_21425);
xnor U21696 (N_21696,N_21274,N_21005);
xnor U21697 (N_21697,N_21176,N_21195);
nor U21698 (N_21698,N_21214,N_21391);
xor U21699 (N_21699,N_21215,N_21388);
nand U21700 (N_21700,N_21475,N_21396);
nor U21701 (N_21701,N_21497,N_21404);
nand U21702 (N_21702,N_21483,N_21321);
nor U21703 (N_21703,N_21008,N_21080);
xor U21704 (N_21704,N_21184,N_21433);
or U21705 (N_21705,N_21260,N_21100);
xor U21706 (N_21706,N_21065,N_21300);
xnor U21707 (N_21707,N_21099,N_21407);
nor U21708 (N_21708,N_21166,N_21319);
nor U21709 (N_21709,N_21367,N_21023);
or U21710 (N_21710,N_21326,N_21459);
xor U21711 (N_21711,N_21276,N_21467);
nand U21712 (N_21712,N_21249,N_21330);
and U21713 (N_21713,N_21298,N_21470);
xnor U21714 (N_21714,N_21200,N_21331);
xnor U21715 (N_21715,N_21085,N_21289);
nor U21716 (N_21716,N_21455,N_21251);
and U21717 (N_21717,N_21064,N_21054);
and U21718 (N_21718,N_21088,N_21441);
or U21719 (N_21719,N_21468,N_21232);
nor U21720 (N_21720,N_21009,N_21107);
nor U21721 (N_21721,N_21146,N_21007);
nand U21722 (N_21722,N_21282,N_21111);
nor U21723 (N_21723,N_21403,N_21246);
nor U21724 (N_21724,N_21144,N_21021);
nor U21725 (N_21725,N_21456,N_21341);
nor U21726 (N_21726,N_21288,N_21026);
or U21727 (N_21727,N_21206,N_21173);
xnor U21728 (N_21728,N_21219,N_21309);
nand U21729 (N_21729,N_21010,N_21275);
nor U21730 (N_21730,N_21436,N_21045);
and U21731 (N_21731,N_21141,N_21415);
or U21732 (N_21732,N_21481,N_21345);
nor U21733 (N_21733,N_21040,N_21346);
nor U21734 (N_21734,N_21221,N_21098);
or U21735 (N_21735,N_21165,N_21258);
nand U21736 (N_21736,N_21410,N_21488);
nor U21737 (N_21737,N_21229,N_21145);
xor U21738 (N_21738,N_21235,N_21086);
nand U21739 (N_21739,N_21158,N_21356);
or U21740 (N_21740,N_21115,N_21490);
nand U21741 (N_21741,N_21427,N_21368);
and U21742 (N_21742,N_21444,N_21264);
nand U21743 (N_21743,N_21328,N_21461);
and U21744 (N_21744,N_21091,N_21486);
nand U21745 (N_21745,N_21259,N_21434);
xor U21746 (N_21746,N_21292,N_21458);
xnor U21747 (N_21747,N_21033,N_21233);
nor U21748 (N_21748,N_21120,N_21181);
and U21749 (N_21749,N_21317,N_21304);
or U21750 (N_21750,N_21218,N_21164);
or U21751 (N_21751,N_21075,N_21367);
nand U21752 (N_21752,N_21273,N_21228);
nor U21753 (N_21753,N_21425,N_21158);
or U21754 (N_21754,N_21103,N_21131);
and U21755 (N_21755,N_21453,N_21208);
nor U21756 (N_21756,N_21189,N_21404);
nor U21757 (N_21757,N_21461,N_21032);
or U21758 (N_21758,N_21452,N_21258);
nor U21759 (N_21759,N_21189,N_21420);
nor U21760 (N_21760,N_21336,N_21086);
nand U21761 (N_21761,N_21396,N_21083);
xor U21762 (N_21762,N_21218,N_21457);
and U21763 (N_21763,N_21082,N_21137);
nor U21764 (N_21764,N_21055,N_21028);
and U21765 (N_21765,N_21211,N_21227);
and U21766 (N_21766,N_21473,N_21002);
nand U21767 (N_21767,N_21141,N_21007);
or U21768 (N_21768,N_21450,N_21385);
xor U21769 (N_21769,N_21482,N_21103);
xor U21770 (N_21770,N_21184,N_21050);
nand U21771 (N_21771,N_21044,N_21205);
or U21772 (N_21772,N_21363,N_21041);
and U21773 (N_21773,N_21125,N_21040);
and U21774 (N_21774,N_21477,N_21273);
xor U21775 (N_21775,N_21234,N_21126);
and U21776 (N_21776,N_21272,N_21002);
and U21777 (N_21777,N_21400,N_21208);
nand U21778 (N_21778,N_21330,N_21456);
and U21779 (N_21779,N_21310,N_21092);
or U21780 (N_21780,N_21386,N_21329);
xor U21781 (N_21781,N_21315,N_21447);
xor U21782 (N_21782,N_21466,N_21474);
nand U21783 (N_21783,N_21222,N_21367);
nand U21784 (N_21784,N_21433,N_21423);
and U21785 (N_21785,N_21096,N_21293);
xor U21786 (N_21786,N_21210,N_21166);
nor U21787 (N_21787,N_21197,N_21136);
or U21788 (N_21788,N_21346,N_21205);
nand U21789 (N_21789,N_21288,N_21330);
xnor U21790 (N_21790,N_21051,N_21400);
or U21791 (N_21791,N_21496,N_21254);
and U21792 (N_21792,N_21497,N_21280);
or U21793 (N_21793,N_21247,N_21403);
nor U21794 (N_21794,N_21282,N_21040);
nor U21795 (N_21795,N_21161,N_21024);
and U21796 (N_21796,N_21061,N_21025);
xnor U21797 (N_21797,N_21068,N_21026);
and U21798 (N_21798,N_21332,N_21322);
or U21799 (N_21799,N_21096,N_21167);
nor U21800 (N_21800,N_21437,N_21446);
xnor U21801 (N_21801,N_21450,N_21214);
nand U21802 (N_21802,N_21380,N_21471);
nand U21803 (N_21803,N_21012,N_21120);
xor U21804 (N_21804,N_21100,N_21068);
and U21805 (N_21805,N_21130,N_21141);
nand U21806 (N_21806,N_21248,N_21215);
xnor U21807 (N_21807,N_21215,N_21039);
xor U21808 (N_21808,N_21487,N_21022);
nand U21809 (N_21809,N_21291,N_21391);
xnor U21810 (N_21810,N_21056,N_21150);
or U21811 (N_21811,N_21028,N_21107);
or U21812 (N_21812,N_21489,N_21296);
or U21813 (N_21813,N_21047,N_21441);
and U21814 (N_21814,N_21424,N_21061);
nor U21815 (N_21815,N_21116,N_21010);
nor U21816 (N_21816,N_21175,N_21367);
nor U21817 (N_21817,N_21077,N_21275);
and U21818 (N_21818,N_21389,N_21254);
nor U21819 (N_21819,N_21322,N_21098);
xor U21820 (N_21820,N_21458,N_21073);
nand U21821 (N_21821,N_21228,N_21114);
xnor U21822 (N_21822,N_21163,N_21294);
nor U21823 (N_21823,N_21498,N_21232);
nand U21824 (N_21824,N_21192,N_21259);
and U21825 (N_21825,N_21315,N_21230);
or U21826 (N_21826,N_21483,N_21369);
or U21827 (N_21827,N_21126,N_21473);
or U21828 (N_21828,N_21092,N_21295);
xnor U21829 (N_21829,N_21239,N_21330);
xnor U21830 (N_21830,N_21297,N_21338);
nand U21831 (N_21831,N_21154,N_21351);
and U21832 (N_21832,N_21070,N_21286);
nor U21833 (N_21833,N_21181,N_21077);
or U21834 (N_21834,N_21350,N_21456);
nor U21835 (N_21835,N_21287,N_21410);
xnor U21836 (N_21836,N_21050,N_21010);
xnor U21837 (N_21837,N_21090,N_21300);
xnor U21838 (N_21838,N_21286,N_21395);
and U21839 (N_21839,N_21080,N_21158);
nor U21840 (N_21840,N_21403,N_21356);
and U21841 (N_21841,N_21172,N_21408);
xor U21842 (N_21842,N_21001,N_21070);
xnor U21843 (N_21843,N_21008,N_21052);
nor U21844 (N_21844,N_21058,N_21374);
nor U21845 (N_21845,N_21243,N_21323);
nand U21846 (N_21846,N_21162,N_21100);
nor U21847 (N_21847,N_21283,N_21158);
xnor U21848 (N_21848,N_21430,N_21006);
xnor U21849 (N_21849,N_21289,N_21187);
or U21850 (N_21850,N_21396,N_21106);
and U21851 (N_21851,N_21212,N_21473);
xor U21852 (N_21852,N_21256,N_21156);
or U21853 (N_21853,N_21469,N_21321);
nand U21854 (N_21854,N_21285,N_21318);
xor U21855 (N_21855,N_21382,N_21022);
or U21856 (N_21856,N_21347,N_21040);
xor U21857 (N_21857,N_21489,N_21201);
nand U21858 (N_21858,N_21106,N_21207);
nor U21859 (N_21859,N_21132,N_21475);
or U21860 (N_21860,N_21000,N_21245);
nor U21861 (N_21861,N_21387,N_21008);
nand U21862 (N_21862,N_21291,N_21121);
nand U21863 (N_21863,N_21485,N_21058);
nor U21864 (N_21864,N_21129,N_21183);
nand U21865 (N_21865,N_21235,N_21385);
nand U21866 (N_21866,N_21489,N_21165);
nand U21867 (N_21867,N_21478,N_21228);
nand U21868 (N_21868,N_21225,N_21236);
nand U21869 (N_21869,N_21039,N_21185);
nand U21870 (N_21870,N_21241,N_21046);
nor U21871 (N_21871,N_21030,N_21373);
or U21872 (N_21872,N_21139,N_21461);
nor U21873 (N_21873,N_21338,N_21433);
nand U21874 (N_21874,N_21177,N_21477);
or U21875 (N_21875,N_21315,N_21092);
or U21876 (N_21876,N_21484,N_21457);
or U21877 (N_21877,N_21356,N_21068);
or U21878 (N_21878,N_21167,N_21276);
and U21879 (N_21879,N_21176,N_21491);
xnor U21880 (N_21880,N_21088,N_21203);
nor U21881 (N_21881,N_21141,N_21323);
xnor U21882 (N_21882,N_21425,N_21076);
and U21883 (N_21883,N_21352,N_21025);
nor U21884 (N_21884,N_21491,N_21053);
nand U21885 (N_21885,N_21327,N_21269);
nor U21886 (N_21886,N_21368,N_21052);
nand U21887 (N_21887,N_21148,N_21033);
and U21888 (N_21888,N_21069,N_21468);
and U21889 (N_21889,N_21070,N_21152);
nand U21890 (N_21890,N_21440,N_21123);
xnor U21891 (N_21891,N_21048,N_21416);
xor U21892 (N_21892,N_21256,N_21375);
or U21893 (N_21893,N_21029,N_21175);
xnor U21894 (N_21894,N_21405,N_21259);
nand U21895 (N_21895,N_21263,N_21233);
nand U21896 (N_21896,N_21120,N_21036);
xor U21897 (N_21897,N_21223,N_21433);
nand U21898 (N_21898,N_21200,N_21494);
and U21899 (N_21899,N_21090,N_21231);
nand U21900 (N_21900,N_21210,N_21224);
or U21901 (N_21901,N_21381,N_21452);
or U21902 (N_21902,N_21038,N_21359);
nand U21903 (N_21903,N_21135,N_21233);
and U21904 (N_21904,N_21034,N_21017);
xor U21905 (N_21905,N_21288,N_21304);
and U21906 (N_21906,N_21104,N_21408);
xor U21907 (N_21907,N_21422,N_21326);
nor U21908 (N_21908,N_21204,N_21119);
xnor U21909 (N_21909,N_21205,N_21131);
or U21910 (N_21910,N_21086,N_21455);
nand U21911 (N_21911,N_21197,N_21352);
xnor U21912 (N_21912,N_21365,N_21480);
nor U21913 (N_21913,N_21209,N_21299);
xnor U21914 (N_21914,N_21442,N_21339);
nand U21915 (N_21915,N_21067,N_21317);
and U21916 (N_21916,N_21490,N_21374);
xnor U21917 (N_21917,N_21090,N_21362);
and U21918 (N_21918,N_21378,N_21093);
and U21919 (N_21919,N_21171,N_21152);
or U21920 (N_21920,N_21228,N_21376);
nand U21921 (N_21921,N_21180,N_21153);
nand U21922 (N_21922,N_21172,N_21387);
xnor U21923 (N_21923,N_21274,N_21192);
xor U21924 (N_21924,N_21085,N_21444);
xor U21925 (N_21925,N_21240,N_21298);
nor U21926 (N_21926,N_21419,N_21005);
or U21927 (N_21927,N_21306,N_21076);
nor U21928 (N_21928,N_21254,N_21440);
nor U21929 (N_21929,N_21198,N_21079);
or U21930 (N_21930,N_21083,N_21458);
nor U21931 (N_21931,N_21476,N_21281);
and U21932 (N_21932,N_21063,N_21131);
and U21933 (N_21933,N_21017,N_21033);
nor U21934 (N_21934,N_21492,N_21457);
nor U21935 (N_21935,N_21443,N_21060);
or U21936 (N_21936,N_21362,N_21111);
nor U21937 (N_21937,N_21309,N_21397);
and U21938 (N_21938,N_21059,N_21224);
nand U21939 (N_21939,N_21206,N_21350);
or U21940 (N_21940,N_21236,N_21255);
xnor U21941 (N_21941,N_21321,N_21155);
and U21942 (N_21942,N_21424,N_21089);
or U21943 (N_21943,N_21423,N_21427);
or U21944 (N_21944,N_21295,N_21085);
and U21945 (N_21945,N_21132,N_21362);
nand U21946 (N_21946,N_21385,N_21334);
nand U21947 (N_21947,N_21035,N_21416);
nor U21948 (N_21948,N_21242,N_21067);
or U21949 (N_21949,N_21329,N_21484);
nand U21950 (N_21950,N_21463,N_21145);
nand U21951 (N_21951,N_21218,N_21376);
or U21952 (N_21952,N_21484,N_21289);
nand U21953 (N_21953,N_21052,N_21073);
xor U21954 (N_21954,N_21025,N_21007);
nand U21955 (N_21955,N_21224,N_21271);
or U21956 (N_21956,N_21322,N_21309);
nand U21957 (N_21957,N_21206,N_21480);
xor U21958 (N_21958,N_21265,N_21048);
or U21959 (N_21959,N_21274,N_21100);
and U21960 (N_21960,N_21225,N_21421);
xnor U21961 (N_21961,N_21041,N_21251);
or U21962 (N_21962,N_21473,N_21377);
and U21963 (N_21963,N_21039,N_21443);
or U21964 (N_21964,N_21438,N_21267);
xor U21965 (N_21965,N_21012,N_21184);
and U21966 (N_21966,N_21013,N_21191);
nand U21967 (N_21967,N_21427,N_21032);
nand U21968 (N_21968,N_21015,N_21284);
and U21969 (N_21969,N_21324,N_21472);
nand U21970 (N_21970,N_21071,N_21237);
and U21971 (N_21971,N_21139,N_21343);
and U21972 (N_21972,N_21440,N_21488);
nand U21973 (N_21973,N_21419,N_21062);
xor U21974 (N_21974,N_21499,N_21408);
xnor U21975 (N_21975,N_21478,N_21280);
nor U21976 (N_21976,N_21278,N_21454);
nor U21977 (N_21977,N_21437,N_21310);
and U21978 (N_21978,N_21427,N_21272);
and U21979 (N_21979,N_21237,N_21050);
nor U21980 (N_21980,N_21343,N_21393);
nand U21981 (N_21981,N_21196,N_21385);
nor U21982 (N_21982,N_21162,N_21369);
xor U21983 (N_21983,N_21347,N_21124);
or U21984 (N_21984,N_21267,N_21135);
or U21985 (N_21985,N_21019,N_21423);
and U21986 (N_21986,N_21441,N_21383);
and U21987 (N_21987,N_21235,N_21443);
and U21988 (N_21988,N_21359,N_21058);
nor U21989 (N_21989,N_21342,N_21429);
and U21990 (N_21990,N_21057,N_21010);
nor U21991 (N_21991,N_21442,N_21009);
nor U21992 (N_21992,N_21407,N_21015);
nor U21993 (N_21993,N_21430,N_21033);
nor U21994 (N_21994,N_21032,N_21158);
nand U21995 (N_21995,N_21133,N_21240);
or U21996 (N_21996,N_21159,N_21186);
nand U21997 (N_21997,N_21405,N_21367);
xor U21998 (N_21998,N_21259,N_21111);
or U21999 (N_21999,N_21270,N_21226);
nor U22000 (N_22000,N_21534,N_21977);
nand U22001 (N_22001,N_21595,N_21758);
xnor U22002 (N_22002,N_21726,N_21675);
nor U22003 (N_22003,N_21916,N_21562);
and U22004 (N_22004,N_21502,N_21770);
nor U22005 (N_22005,N_21721,N_21827);
or U22006 (N_22006,N_21983,N_21926);
nor U22007 (N_22007,N_21563,N_21570);
nor U22008 (N_22008,N_21897,N_21915);
xor U22009 (N_22009,N_21564,N_21814);
nor U22010 (N_22010,N_21628,N_21727);
or U22011 (N_22011,N_21875,N_21906);
xnor U22012 (N_22012,N_21512,N_21792);
nor U22013 (N_22013,N_21995,N_21852);
nand U22014 (N_22014,N_21962,N_21691);
and U22015 (N_22015,N_21781,N_21637);
or U22016 (N_22016,N_21524,N_21924);
and U22017 (N_22017,N_21687,N_21971);
nand U22018 (N_22018,N_21544,N_21677);
nor U22019 (N_22019,N_21937,N_21704);
and U22020 (N_22020,N_21881,N_21829);
nand U22021 (N_22021,N_21813,N_21606);
or U22022 (N_22022,N_21766,N_21907);
or U22023 (N_22023,N_21561,N_21550);
nand U22024 (N_22024,N_21988,N_21627);
nand U22025 (N_22025,N_21948,N_21608);
or U22026 (N_22026,N_21670,N_21543);
xor U22027 (N_22027,N_21690,N_21892);
nand U22028 (N_22028,N_21588,N_21902);
xor U22029 (N_22029,N_21879,N_21755);
and U22030 (N_22030,N_21894,N_21530);
xnor U22031 (N_22031,N_21982,N_21750);
nand U22032 (N_22032,N_21749,N_21836);
nand U22033 (N_22033,N_21617,N_21643);
and U22034 (N_22034,N_21692,N_21993);
nand U22035 (N_22035,N_21854,N_21735);
nor U22036 (N_22036,N_21508,N_21669);
nand U22037 (N_22037,N_21647,N_21644);
nor U22038 (N_22038,N_21934,N_21659);
xnor U22039 (N_22039,N_21753,N_21972);
nand U22040 (N_22040,N_21509,N_21600);
xnor U22041 (N_22041,N_21652,N_21837);
nand U22042 (N_22042,N_21985,N_21678);
xnor U22043 (N_22043,N_21999,N_21701);
or U22044 (N_22044,N_21807,N_21519);
nand U22045 (N_22045,N_21604,N_21980);
nor U22046 (N_22046,N_21861,N_21855);
nor U22047 (N_22047,N_21525,N_21905);
xnor U22048 (N_22048,N_21674,N_21707);
nor U22049 (N_22049,N_21865,N_21660);
nor U22050 (N_22050,N_21506,N_21858);
nand U22051 (N_22051,N_21762,N_21812);
or U22052 (N_22052,N_21532,N_21953);
and U22053 (N_22053,N_21739,N_21918);
nand U22054 (N_22054,N_21803,N_21733);
xnor U22055 (N_22055,N_21997,N_21996);
or U22056 (N_22056,N_21682,N_21956);
nand U22057 (N_22057,N_21901,N_21624);
nand U22058 (N_22058,N_21540,N_21752);
nor U22059 (N_22059,N_21898,N_21783);
nor U22060 (N_22060,N_21516,N_21870);
xnor U22061 (N_22061,N_21789,N_21715);
xnor U22062 (N_22062,N_21947,N_21941);
nand U22063 (N_22063,N_21683,N_21969);
and U22064 (N_22064,N_21922,N_21945);
nor U22065 (N_22065,N_21642,N_21976);
xnor U22066 (N_22066,N_21695,N_21528);
or U22067 (N_22067,N_21859,N_21848);
xor U22068 (N_22068,N_21869,N_21793);
nor U22069 (N_22069,N_21613,N_21957);
xnor U22070 (N_22070,N_21640,N_21621);
nor U22071 (N_22071,N_21574,N_21790);
or U22072 (N_22072,N_21705,N_21620);
nor U22073 (N_22073,N_21984,N_21594);
or U22074 (N_22074,N_21679,N_21919);
nor U22075 (N_22075,N_21602,N_21830);
and U22076 (N_22076,N_21787,N_21741);
and U22077 (N_22077,N_21951,N_21936);
nand U22078 (N_22078,N_21834,N_21863);
nor U22079 (N_22079,N_21746,N_21522);
and U22080 (N_22080,N_21759,N_21754);
nor U22081 (N_22081,N_21603,N_21719);
and U22082 (N_22082,N_21992,N_21587);
nor U22083 (N_22083,N_21514,N_21895);
xnor U22084 (N_22084,N_21850,N_21538);
xor U22085 (N_22085,N_21943,N_21541);
xnor U22086 (N_22086,N_21504,N_21559);
xnor U22087 (N_22087,N_21709,N_21968);
xor U22088 (N_22088,N_21625,N_21772);
xor U22089 (N_22089,N_21843,N_21839);
xnor U22090 (N_22090,N_21648,N_21761);
xor U22091 (N_22091,N_21927,N_21586);
xor U22092 (N_22092,N_21964,N_21661);
nor U22093 (N_22093,N_21886,N_21501);
nor U22094 (N_22094,N_21728,N_21884);
nand U22095 (N_22095,N_21638,N_21649);
xnor U22096 (N_22096,N_21819,N_21515);
or U22097 (N_22097,N_21979,N_21663);
or U22098 (N_22098,N_21605,N_21856);
or U22099 (N_22099,N_21929,N_21584);
xnor U22100 (N_22100,N_21511,N_21725);
nor U22101 (N_22101,N_21517,N_21801);
and U22102 (N_22102,N_21928,N_21656);
or U22103 (N_22103,N_21802,N_21536);
or U22104 (N_22104,N_21986,N_21558);
nand U22105 (N_22105,N_21713,N_21958);
or U22106 (N_22106,N_21533,N_21944);
nand U22107 (N_22107,N_21629,N_21805);
or U22108 (N_22108,N_21763,N_21526);
or U22109 (N_22109,N_21824,N_21622);
and U22110 (N_22110,N_21871,N_21903);
xnor U22111 (N_22111,N_21932,N_21589);
nand U22112 (N_22112,N_21828,N_21880);
nor U22113 (N_22113,N_21745,N_21645);
nor U22114 (N_22114,N_21811,N_21998);
or U22115 (N_22115,N_21833,N_21655);
nor U22116 (N_22116,N_21592,N_21662);
and U22117 (N_22117,N_21917,N_21966);
nor U22118 (N_22118,N_21568,N_21842);
nand U22119 (N_22119,N_21942,N_21867);
and U22120 (N_22120,N_21612,N_21940);
nor U22121 (N_22121,N_21959,N_21954);
and U22122 (N_22122,N_21712,N_21731);
nor U22123 (N_22123,N_21900,N_21885);
or U22124 (N_22124,N_21791,N_21553);
nor U22125 (N_22125,N_21684,N_21706);
and U22126 (N_22126,N_21653,N_21641);
or U22127 (N_22127,N_21702,N_21777);
nor U22128 (N_22128,N_21809,N_21673);
nor U22129 (N_22129,N_21989,N_21665);
or U22130 (N_22130,N_21711,N_21694);
xnor U22131 (N_22131,N_21569,N_21551);
nand U22132 (N_22132,N_21639,N_21930);
nor U22133 (N_22133,N_21714,N_21887);
and U22134 (N_22134,N_21717,N_21831);
or U22135 (N_22135,N_21557,N_21838);
or U22136 (N_22136,N_21596,N_21667);
nand U22137 (N_22137,N_21862,N_21573);
xor U22138 (N_22138,N_21780,N_21878);
and U22139 (N_22139,N_21832,N_21732);
and U22140 (N_22140,N_21693,N_21967);
nor U22141 (N_22141,N_21666,N_21632);
xor U22142 (N_22142,N_21730,N_21910);
and U22143 (N_22143,N_21555,N_21591);
xnor U22144 (N_22144,N_21935,N_21974);
xor U22145 (N_22145,N_21877,N_21529);
xor U22146 (N_22146,N_21668,N_21868);
nor U22147 (N_22147,N_21537,N_21912);
nor U22148 (N_22148,N_21883,N_21841);
nor U22149 (N_22149,N_21891,N_21981);
xnor U22150 (N_22150,N_21821,N_21527);
xnor U22151 (N_22151,N_21688,N_21565);
nor U22152 (N_22152,N_21576,N_21575);
or U22153 (N_22153,N_21866,N_21521);
xnor U22154 (N_22154,N_21896,N_21775);
nand U22155 (N_22155,N_21931,N_21990);
and U22156 (N_22156,N_21938,N_21657);
xnor U22157 (N_22157,N_21840,N_21611);
nor U22158 (N_22158,N_21994,N_21946);
nor U22159 (N_22159,N_21788,N_21925);
xnor U22160 (N_22160,N_21742,N_21808);
or U22161 (N_22161,N_21864,N_21939);
nand U22162 (N_22162,N_21955,N_21546);
xor U22163 (N_22163,N_21718,N_21510);
nor U22164 (N_22164,N_21991,N_21699);
nand U22165 (N_22165,N_21796,N_21823);
nand U22166 (N_22166,N_21609,N_21744);
nand U22167 (N_22167,N_21820,N_21631);
nor U22168 (N_22168,N_21961,N_21876);
or U22169 (N_22169,N_21797,N_21610);
xnor U22170 (N_22170,N_21676,N_21582);
and U22171 (N_22171,N_21874,N_21810);
nor U22172 (N_22172,N_21978,N_21952);
or U22173 (N_22173,N_21720,N_21554);
and U22174 (N_22174,N_21724,N_21580);
xnor U22175 (N_22175,N_21571,N_21549);
nand U22176 (N_22176,N_21716,N_21654);
and U22177 (N_22177,N_21882,N_21520);
or U22178 (N_22178,N_21548,N_21723);
and U22179 (N_22179,N_21736,N_21740);
nand U22180 (N_22180,N_21963,N_21646);
or U22181 (N_22181,N_21578,N_21703);
or U22182 (N_22182,N_21768,N_21773);
nor U22183 (N_22183,N_21556,N_21748);
or U22184 (N_22184,N_21960,N_21626);
and U22185 (N_22185,N_21698,N_21597);
or U22186 (N_22186,N_21970,N_21598);
and U22187 (N_22187,N_21531,N_21923);
and U22188 (N_22188,N_21686,N_21616);
xor U22189 (N_22189,N_21806,N_21633);
xnor U22190 (N_22190,N_21623,N_21784);
nor U22191 (N_22191,N_21835,N_21904);
or U22192 (N_22192,N_21671,N_21817);
nor U22193 (N_22193,N_21794,N_21685);
or U22194 (N_22194,N_21585,N_21844);
and U22195 (N_22195,N_21581,N_21975);
and U22196 (N_22196,N_21756,N_21888);
or U22197 (N_22197,N_21503,N_21743);
nand U22198 (N_22198,N_21920,N_21889);
or U22199 (N_22199,N_21590,N_21764);
nand U22200 (N_22200,N_21710,N_21542);
nand U22201 (N_22201,N_21615,N_21729);
nand U22202 (N_22202,N_21618,N_21872);
nand U22203 (N_22203,N_21816,N_21851);
nand U22204 (N_22204,N_21607,N_21579);
xnor U22205 (N_22205,N_21547,N_21765);
xnor U22206 (N_22206,N_21760,N_21696);
xnor U22207 (N_22207,N_21630,N_21507);
or U22208 (N_22208,N_21846,N_21689);
and U22209 (N_22209,N_21577,N_21893);
nand U22210 (N_22210,N_21751,N_21545);
nand U22211 (N_22211,N_21847,N_21518);
nor U22212 (N_22212,N_21965,N_21853);
nand U22213 (N_22213,N_21908,N_21672);
nor U22214 (N_22214,N_21815,N_21769);
and U22215 (N_22215,N_21505,N_21914);
nor U22216 (N_22216,N_21798,N_21973);
nor U22217 (N_22217,N_21890,N_21800);
or U22218 (N_22218,N_21566,N_21795);
and U22219 (N_22219,N_21500,N_21635);
and U22220 (N_22220,N_21658,N_21785);
nand U22221 (N_22221,N_21681,N_21949);
and U22222 (N_22222,N_21734,N_21767);
xnor U22223 (N_22223,N_21737,N_21513);
nor U22224 (N_22224,N_21697,N_21747);
and U22225 (N_22225,N_21804,N_21523);
nand U22226 (N_22226,N_21539,N_21987);
or U22227 (N_22227,N_21757,N_21651);
or U22228 (N_22228,N_21722,N_21799);
xnor U22229 (N_22229,N_21664,N_21650);
xnor U22230 (N_22230,N_21552,N_21825);
nand U22231 (N_22231,N_21680,N_21860);
nor U22232 (N_22232,N_21636,N_21700);
nor U22233 (N_22233,N_21567,N_21822);
and U22234 (N_22234,N_21849,N_21913);
or U22235 (N_22235,N_21771,N_21778);
xor U22236 (N_22236,N_21933,N_21779);
or U22237 (N_22237,N_21776,N_21857);
nor U22238 (N_22238,N_21535,N_21911);
xnor U22239 (N_22239,N_21738,N_21818);
xor U22240 (N_22240,N_21786,N_21873);
and U22241 (N_22241,N_21950,N_21599);
nor U22242 (N_22242,N_21619,N_21774);
and U22243 (N_22243,N_21909,N_21634);
xnor U22244 (N_22244,N_21782,N_21899);
or U22245 (N_22245,N_21845,N_21826);
or U22246 (N_22246,N_21593,N_21614);
and U22247 (N_22247,N_21921,N_21560);
xor U22248 (N_22248,N_21572,N_21583);
and U22249 (N_22249,N_21601,N_21708);
or U22250 (N_22250,N_21932,N_21857);
nand U22251 (N_22251,N_21909,N_21532);
nand U22252 (N_22252,N_21998,N_21552);
nor U22253 (N_22253,N_21924,N_21723);
and U22254 (N_22254,N_21797,N_21979);
and U22255 (N_22255,N_21509,N_21577);
nor U22256 (N_22256,N_21782,N_21833);
or U22257 (N_22257,N_21856,N_21740);
and U22258 (N_22258,N_21784,N_21514);
and U22259 (N_22259,N_21590,N_21660);
or U22260 (N_22260,N_21746,N_21756);
nor U22261 (N_22261,N_21677,N_21703);
nor U22262 (N_22262,N_21959,N_21977);
and U22263 (N_22263,N_21583,N_21797);
nand U22264 (N_22264,N_21566,N_21578);
and U22265 (N_22265,N_21931,N_21711);
nor U22266 (N_22266,N_21561,N_21838);
nand U22267 (N_22267,N_21764,N_21680);
and U22268 (N_22268,N_21507,N_21906);
and U22269 (N_22269,N_21801,N_21510);
and U22270 (N_22270,N_21852,N_21591);
nor U22271 (N_22271,N_21713,N_21994);
xor U22272 (N_22272,N_21582,N_21780);
and U22273 (N_22273,N_21832,N_21538);
or U22274 (N_22274,N_21576,N_21810);
nand U22275 (N_22275,N_21519,N_21852);
or U22276 (N_22276,N_21800,N_21670);
nand U22277 (N_22277,N_21932,N_21934);
or U22278 (N_22278,N_21863,N_21892);
nand U22279 (N_22279,N_21951,N_21968);
and U22280 (N_22280,N_21554,N_21534);
nor U22281 (N_22281,N_21721,N_21953);
and U22282 (N_22282,N_21614,N_21797);
nor U22283 (N_22283,N_21603,N_21980);
and U22284 (N_22284,N_21824,N_21556);
xor U22285 (N_22285,N_21695,N_21922);
and U22286 (N_22286,N_21987,N_21504);
or U22287 (N_22287,N_21845,N_21858);
nor U22288 (N_22288,N_21674,N_21758);
or U22289 (N_22289,N_21510,N_21903);
nor U22290 (N_22290,N_21977,N_21775);
and U22291 (N_22291,N_21869,N_21798);
nor U22292 (N_22292,N_21682,N_21529);
or U22293 (N_22293,N_21545,N_21930);
nor U22294 (N_22294,N_21669,N_21618);
xnor U22295 (N_22295,N_21681,N_21542);
nor U22296 (N_22296,N_21651,N_21991);
nor U22297 (N_22297,N_21727,N_21954);
or U22298 (N_22298,N_21834,N_21939);
and U22299 (N_22299,N_21525,N_21743);
or U22300 (N_22300,N_21876,N_21820);
xor U22301 (N_22301,N_21555,N_21973);
xnor U22302 (N_22302,N_21922,N_21520);
or U22303 (N_22303,N_21929,N_21864);
or U22304 (N_22304,N_21776,N_21772);
nand U22305 (N_22305,N_21872,N_21622);
nand U22306 (N_22306,N_21524,N_21502);
or U22307 (N_22307,N_21673,N_21845);
nor U22308 (N_22308,N_21863,N_21733);
or U22309 (N_22309,N_21637,N_21764);
xnor U22310 (N_22310,N_21805,N_21902);
or U22311 (N_22311,N_21705,N_21671);
or U22312 (N_22312,N_21936,N_21882);
nor U22313 (N_22313,N_21900,N_21967);
or U22314 (N_22314,N_21982,N_21521);
nor U22315 (N_22315,N_21752,N_21677);
and U22316 (N_22316,N_21529,N_21789);
or U22317 (N_22317,N_21942,N_21819);
nor U22318 (N_22318,N_21588,N_21538);
and U22319 (N_22319,N_21600,N_21687);
or U22320 (N_22320,N_21708,N_21597);
and U22321 (N_22321,N_21545,N_21521);
and U22322 (N_22322,N_21774,N_21688);
nor U22323 (N_22323,N_21876,N_21534);
xor U22324 (N_22324,N_21744,N_21592);
nor U22325 (N_22325,N_21538,N_21649);
nor U22326 (N_22326,N_21699,N_21696);
and U22327 (N_22327,N_21623,N_21796);
xor U22328 (N_22328,N_21864,N_21633);
nand U22329 (N_22329,N_21671,N_21894);
or U22330 (N_22330,N_21787,N_21988);
or U22331 (N_22331,N_21604,N_21871);
xnor U22332 (N_22332,N_21817,N_21909);
and U22333 (N_22333,N_21824,N_21600);
nand U22334 (N_22334,N_21692,N_21593);
and U22335 (N_22335,N_21755,N_21926);
nor U22336 (N_22336,N_21533,N_21520);
nor U22337 (N_22337,N_21582,N_21508);
nor U22338 (N_22338,N_21623,N_21656);
xnor U22339 (N_22339,N_21915,N_21680);
nor U22340 (N_22340,N_21714,N_21744);
and U22341 (N_22341,N_21655,N_21870);
and U22342 (N_22342,N_21596,N_21932);
or U22343 (N_22343,N_21937,N_21567);
and U22344 (N_22344,N_21505,N_21830);
xor U22345 (N_22345,N_21859,N_21629);
xnor U22346 (N_22346,N_21941,N_21788);
xnor U22347 (N_22347,N_21943,N_21749);
nand U22348 (N_22348,N_21743,N_21618);
or U22349 (N_22349,N_21990,N_21833);
xor U22350 (N_22350,N_21834,N_21594);
xor U22351 (N_22351,N_21554,N_21598);
and U22352 (N_22352,N_21740,N_21538);
xor U22353 (N_22353,N_21704,N_21570);
or U22354 (N_22354,N_21963,N_21815);
nor U22355 (N_22355,N_21689,N_21966);
nor U22356 (N_22356,N_21998,N_21710);
nand U22357 (N_22357,N_21652,N_21808);
xnor U22358 (N_22358,N_21889,N_21565);
xor U22359 (N_22359,N_21683,N_21870);
nor U22360 (N_22360,N_21939,N_21661);
or U22361 (N_22361,N_21892,N_21765);
or U22362 (N_22362,N_21572,N_21640);
nand U22363 (N_22363,N_21887,N_21825);
nor U22364 (N_22364,N_21795,N_21831);
or U22365 (N_22365,N_21638,N_21827);
nand U22366 (N_22366,N_21555,N_21552);
or U22367 (N_22367,N_21885,N_21611);
and U22368 (N_22368,N_21823,N_21568);
and U22369 (N_22369,N_21819,N_21529);
xor U22370 (N_22370,N_21845,N_21752);
and U22371 (N_22371,N_21972,N_21749);
and U22372 (N_22372,N_21651,N_21532);
nor U22373 (N_22373,N_21910,N_21759);
nor U22374 (N_22374,N_21534,N_21968);
or U22375 (N_22375,N_21549,N_21650);
nand U22376 (N_22376,N_21816,N_21507);
and U22377 (N_22377,N_21888,N_21604);
xnor U22378 (N_22378,N_21929,N_21845);
nor U22379 (N_22379,N_21966,N_21714);
nor U22380 (N_22380,N_21578,N_21512);
nor U22381 (N_22381,N_21770,N_21861);
nor U22382 (N_22382,N_21720,N_21779);
nor U22383 (N_22383,N_21783,N_21980);
and U22384 (N_22384,N_21894,N_21679);
or U22385 (N_22385,N_21757,N_21533);
nor U22386 (N_22386,N_21960,N_21980);
or U22387 (N_22387,N_21911,N_21966);
nand U22388 (N_22388,N_21608,N_21831);
and U22389 (N_22389,N_21507,N_21876);
or U22390 (N_22390,N_21628,N_21815);
or U22391 (N_22391,N_21825,N_21900);
or U22392 (N_22392,N_21558,N_21834);
nor U22393 (N_22393,N_21892,N_21783);
xnor U22394 (N_22394,N_21892,N_21617);
or U22395 (N_22395,N_21840,N_21905);
nor U22396 (N_22396,N_21911,N_21525);
and U22397 (N_22397,N_21580,N_21504);
or U22398 (N_22398,N_21996,N_21836);
xor U22399 (N_22399,N_21759,N_21933);
and U22400 (N_22400,N_21938,N_21590);
or U22401 (N_22401,N_21531,N_21928);
nand U22402 (N_22402,N_21942,N_21568);
or U22403 (N_22403,N_21910,N_21924);
and U22404 (N_22404,N_21982,N_21933);
or U22405 (N_22405,N_21787,N_21837);
nor U22406 (N_22406,N_21846,N_21806);
nor U22407 (N_22407,N_21912,N_21666);
xnor U22408 (N_22408,N_21615,N_21781);
and U22409 (N_22409,N_21952,N_21530);
nand U22410 (N_22410,N_21816,N_21548);
or U22411 (N_22411,N_21526,N_21698);
xnor U22412 (N_22412,N_21661,N_21892);
nand U22413 (N_22413,N_21872,N_21800);
xor U22414 (N_22414,N_21672,N_21763);
or U22415 (N_22415,N_21960,N_21795);
and U22416 (N_22416,N_21814,N_21703);
xnor U22417 (N_22417,N_21603,N_21833);
and U22418 (N_22418,N_21508,N_21600);
xor U22419 (N_22419,N_21959,N_21692);
nor U22420 (N_22420,N_21865,N_21548);
nand U22421 (N_22421,N_21742,N_21533);
nand U22422 (N_22422,N_21906,N_21866);
nor U22423 (N_22423,N_21530,N_21773);
and U22424 (N_22424,N_21760,N_21579);
nand U22425 (N_22425,N_21690,N_21593);
and U22426 (N_22426,N_21790,N_21692);
nand U22427 (N_22427,N_21609,N_21594);
or U22428 (N_22428,N_21792,N_21598);
nor U22429 (N_22429,N_21768,N_21703);
xor U22430 (N_22430,N_21529,N_21842);
or U22431 (N_22431,N_21897,N_21994);
nand U22432 (N_22432,N_21536,N_21752);
or U22433 (N_22433,N_21718,N_21689);
or U22434 (N_22434,N_21662,N_21502);
xor U22435 (N_22435,N_21887,N_21623);
or U22436 (N_22436,N_21721,N_21770);
or U22437 (N_22437,N_21711,N_21845);
xnor U22438 (N_22438,N_21818,N_21563);
and U22439 (N_22439,N_21934,N_21707);
and U22440 (N_22440,N_21862,N_21846);
and U22441 (N_22441,N_21829,N_21705);
xor U22442 (N_22442,N_21626,N_21502);
nand U22443 (N_22443,N_21605,N_21727);
and U22444 (N_22444,N_21504,N_21890);
and U22445 (N_22445,N_21936,N_21859);
or U22446 (N_22446,N_21533,N_21995);
or U22447 (N_22447,N_21977,N_21966);
nor U22448 (N_22448,N_21993,N_21734);
or U22449 (N_22449,N_21917,N_21984);
xnor U22450 (N_22450,N_21832,N_21808);
nor U22451 (N_22451,N_21915,N_21773);
xnor U22452 (N_22452,N_21753,N_21789);
and U22453 (N_22453,N_21771,N_21565);
nor U22454 (N_22454,N_21974,N_21516);
or U22455 (N_22455,N_21817,N_21989);
or U22456 (N_22456,N_21783,N_21849);
xor U22457 (N_22457,N_21709,N_21872);
and U22458 (N_22458,N_21531,N_21749);
nand U22459 (N_22459,N_21546,N_21659);
xnor U22460 (N_22460,N_21582,N_21860);
nor U22461 (N_22461,N_21929,N_21602);
and U22462 (N_22462,N_21672,N_21572);
nor U22463 (N_22463,N_21927,N_21903);
xor U22464 (N_22464,N_21951,N_21783);
nand U22465 (N_22465,N_21554,N_21501);
or U22466 (N_22466,N_21933,N_21979);
or U22467 (N_22467,N_21563,N_21691);
or U22468 (N_22468,N_21703,N_21517);
xnor U22469 (N_22469,N_21622,N_21507);
and U22470 (N_22470,N_21539,N_21525);
nor U22471 (N_22471,N_21695,N_21628);
and U22472 (N_22472,N_21598,N_21631);
nand U22473 (N_22473,N_21551,N_21749);
nand U22474 (N_22474,N_21547,N_21893);
xnor U22475 (N_22475,N_21722,N_21800);
nor U22476 (N_22476,N_21673,N_21716);
nand U22477 (N_22477,N_21901,N_21921);
or U22478 (N_22478,N_21768,N_21531);
nor U22479 (N_22479,N_21976,N_21726);
or U22480 (N_22480,N_21912,N_21740);
xor U22481 (N_22481,N_21792,N_21970);
or U22482 (N_22482,N_21578,N_21875);
xor U22483 (N_22483,N_21502,N_21928);
and U22484 (N_22484,N_21565,N_21779);
xor U22485 (N_22485,N_21983,N_21944);
and U22486 (N_22486,N_21676,N_21672);
or U22487 (N_22487,N_21668,N_21859);
nor U22488 (N_22488,N_21827,N_21543);
or U22489 (N_22489,N_21769,N_21500);
and U22490 (N_22490,N_21893,N_21846);
or U22491 (N_22491,N_21658,N_21556);
and U22492 (N_22492,N_21982,N_21601);
nor U22493 (N_22493,N_21829,N_21797);
or U22494 (N_22494,N_21610,N_21802);
or U22495 (N_22495,N_21718,N_21834);
nor U22496 (N_22496,N_21796,N_21957);
xnor U22497 (N_22497,N_21758,N_21930);
xnor U22498 (N_22498,N_21952,N_21779);
xor U22499 (N_22499,N_21905,N_21649);
nand U22500 (N_22500,N_22378,N_22481);
xnor U22501 (N_22501,N_22075,N_22036);
nor U22502 (N_22502,N_22346,N_22277);
nor U22503 (N_22503,N_22003,N_22086);
and U22504 (N_22504,N_22441,N_22002);
nand U22505 (N_22505,N_22436,N_22280);
nand U22506 (N_22506,N_22097,N_22491);
nor U22507 (N_22507,N_22094,N_22389);
and U22508 (N_22508,N_22178,N_22234);
and U22509 (N_22509,N_22259,N_22463);
nand U22510 (N_22510,N_22046,N_22454);
and U22511 (N_22511,N_22394,N_22477);
xor U22512 (N_22512,N_22239,N_22130);
or U22513 (N_22513,N_22254,N_22348);
or U22514 (N_22514,N_22054,N_22453);
or U22515 (N_22515,N_22123,N_22141);
nor U22516 (N_22516,N_22290,N_22332);
xor U22517 (N_22517,N_22139,N_22342);
or U22518 (N_22518,N_22373,N_22474);
nor U22519 (N_22519,N_22063,N_22048);
nor U22520 (N_22520,N_22150,N_22319);
and U22521 (N_22521,N_22037,N_22228);
and U22522 (N_22522,N_22371,N_22146);
nor U22523 (N_22523,N_22038,N_22349);
nand U22524 (N_22524,N_22308,N_22118);
xnor U22525 (N_22525,N_22102,N_22187);
nor U22526 (N_22526,N_22096,N_22467);
nand U22527 (N_22527,N_22471,N_22266);
or U22528 (N_22528,N_22238,N_22461);
or U22529 (N_22529,N_22232,N_22242);
nand U22530 (N_22530,N_22320,N_22338);
or U22531 (N_22531,N_22257,N_22128);
nor U22532 (N_22532,N_22240,N_22489);
xor U22533 (N_22533,N_22093,N_22482);
or U22534 (N_22534,N_22050,N_22060);
and U22535 (N_22535,N_22412,N_22044);
or U22536 (N_22536,N_22137,N_22111);
xnor U22537 (N_22537,N_22397,N_22370);
nand U22538 (N_22538,N_22161,N_22487);
xor U22539 (N_22539,N_22227,N_22143);
and U22540 (N_22540,N_22388,N_22419);
nor U22541 (N_22541,N_22034,N_22466);
or U22542 (N_22542,N_22088,N_22233);
nand U22543 (N_22543,N_22306,N_22104);
or U22544 (N_22544,N_22458,N_22212);
or U22545 (N_22545,N_22116,N_22399);
xnor U22546 (N_22546,N_22084,N_22082);
and U22547 (N_22547,N_22149,N_22327);
and U22548 (N_22548,N_22425,N_22005);
nand U22549 (N_22549,N_22087,N_22427);
xnor U22550 (N_22550,N_22330,N_22208);
nand U22551 (N_22551,N_22494,N_22127);
xor U22552 (N_22552,N_22179,N_22032);
xnor U22553 (N_22553,N_22249,N_22193);
and U22554 (N_22554,N_22076,N_22424);
xor U22555 (N_22555,N_22016,N_22169);
and U22556 (N_22556,N_22080,N_22194);
or U22557 (N_22557,N_22231,N_22056);
or U22558 (N_22558,N_22386,N_22019);
or U22559 (N_22559,N_22070,N_22451);
or U22560 (N_22560,N_22288,N_22243);
nand U22561 (N_22561,N_22433,N_22011);
or U22562 (N_22562,N_22113,N_22405);
or U22563 (N_22563,N_22354,N_22432);
nor U22564 (N_22564,N_22160,N_22421);
or U22565 (N_22565,N_22068,N_22183);
or U22566 (N_22566,N_22331,N_22335);
xnor U22567 (N_22567,N_22138,N_22140);
and U22568 (N_22568,N_22055,N_22449);
nor U22569 (N_22569,N_22291,N_22058);
and U22570 (N_22570,N_22101,N_22017);
nor U22571 (N_22571,N_22091,N_22448);
or U22572 (N_22572,N_22316,N_22000);
or U22573 (N_22573,N_22013,N_22099);
nor U22574 (N_22574,N_22196,N_22192);
nor U22575 (N_22575,N_22269,N_22365);
or U22576 (N_22576,N_22457,N_22109);
or U22577 (N_22577,N_22301,N_22476);
nor U22578 (N_22578,N_22153,N_22337);
nor U22579 (N_22579,N_22081,N_22434);
and U22580 (N_22580,N_22163,N_22031);
or U22581 (N_22581,N_22490,N_22384);
and U22582 (N_22582,N_22041,N_22224);
xnor U22583 (N_22583,N_22030,N_22355);
nor U22584 (N_22584,N_22237,N_22112);
nand U22585 (N_22585,N_22184,N_22006);
nor U22586 (N_22586,N_22195,N_22106);
nor U22587 (N_22587,N_22162,N_22014);
nor U22588 (N_22588,N_22148,N_22326);
xnor U22589 (N_22589,N_22340,N_22136);
and U22590 (N_22590,N_22374,N_22008);
or U22591 (N_22591,N_22012,N_22176);
xnor U22592 (N_22592,N_22430,N_22159);
and U22593 (N_22593,N_22318,N_22324);
xnor U22594 (N_22594,N_22411,N_22429);
nand U22595 (N_22595,N_22125,N_22428);
nor U22596 (N_22596,N_22189,N_22217);
nand U22597 (N_22597,N_22049,N_22083);
nand U22598 (N_22598,N_22135,N_22317);
xor U22599 (N_22599,N_22040,N_22360);
nor U22600 (N_22600,N_22133,N_22214);
and U22601 (N_22601,N_22473,N_22278);
nor U22602 (N_22602,N_22283,N_22376);
xor U22603 (N_22603,N_22268,N_22416);
nor U22604 (N_22604,N_22039,N_22276);
or U22605 (N_22605,N_22312,N_22334);
or U22606 (N_22606,N_22270,N_22156);
nand U22607 (N_22607,N_22236,N_22444);
nor U22608 (N_22608,N_22368,N_22252);
nor U22609 (N_22609,N_22062,N_22078);
or U22610 (N_22610,N_22251,N_22390);
and U22611 (N_22611,N_22447,N_22413);
or U22612 (N_22612,N_22459,N_22171);
or U22613 (N_22613,N_22119,N_22170);
or U22614 (N_22614,N_22307,N_22166);
xnor U22615 (N_22615,N_22035,N_22213);
or U22616 (N_22616,N_22007,N_22498);
nor U22617 (N_22617,N_22381,N_22328);
nor U22618 (N_22618,N_22158,N_22061);
xnor U22619 (N_22619,N_22379,N_22377);
or U22620 (N_22620,N_22085,N_22464);
nor U22621 (N_22621,N_22406,N_22391);
or U22622 (N_22622,N_22216,N_22296);
xor U22623 (N_22623,N_22356,N_22369);
xor U22624 (N_22624,N_22485,N_22226);
or U22625 (N_22625,N_22345,N_22418);
nor U22626 (N_22626,N_22336,N_22387);
nand U22627 (N_22627,N_22190,N_22366);
nand U22628 (N_22628,N_22359,N_22339);
or U22629 (N_22629,N_22281,N_22333);
or U22630 (N_22630,N_22262,N_22175);
nand U22631 (N_22631,N_22244,N_22470);
and U22632 (N_22632,N_22465,N_22051);
and U22633 (N_22633,N_22486,N_22205);
or U22634 (N_22634,N_22004,N_22066);
nor U22635 (N_22635,N_22261,N_22154);
and U22636 (N_22636,N_22472,N_22015);
xor U22637 (N_22637,N_22478,N_22009);
and U22638 (N_22638,N_22230,N_22462);
and U22639 (N_22639,N_22253,N_22396);
nor U22640 (N_22640,N_22435,N_22298);
nand U22641 (N_22641,N_22185,N_22495);
nand U22642 (N_22642,N_22404,N_22198);
nand U22643 (N_22643,N_22279,N_22392);
nor U22644 (N_22644,N_22071,N_22199);
or U22645 (N_22645,N_22053,N_22284);
nand U22646 (N_22646,N_22382,N_22393);
xor U22647 (N_22647,N_22285,N_22028);
nor U22648 (N_22648,N_22426,N_22303);
xnor U22649 (N_22649,N_22311,N_22151);
or U22650 (N_22650,N_22247,N_22442);
or U22651 (N_22651,N_22264,N_22010);
xnor U22652 (N_22652,N_22440,N_22452);
or U22653 (N_22653,N_22206,N_22181);
nand U22654 (N_22654,N_22351,N_22245);
xor U22655 (N_22655,N_22410,N_22289);
nor U22656 (N_22656,N_22493,N_22124);
and U22657 (N_22657,N_22201,N_22045);
nor U22658 (N_22658,N_22165,N_22114);
and U22659 (N_22659,N_22282,N_22321);
nor U22660 (N_22660,N_22177,N_22409);
nand U22661 (N_22661,N_22267,N_22431);
nor U22662 (N_22662,N_22021,N_22222);
or U22663 (N_22663,N_22408,N_22001);
or U22664 (N_22664,N_22023,N_22287);
nand U22665 (N_22665,N_22152,N_22069);
nor U22666 (N_22666,N_22100,N_22380);
nor U22667 (N_22667,N_22414,N_22455);
nand U22668 (N_22668,N_22203,N_22357);
or U22669 (N_22669,N_22142,N_22157);
nand U22670 (N_22670,N_22188,N_22353);
nor U22671 (N_22671,N_22367,N_22042);
xor U22672 (N_22672,N_22126,N_22469);
and U22673 (N_22673,N_22246,N_22313);
nand U22674 (N_22674,N_22173,N_22225);
nand U22675 (N_22675,N_22347,N_22372);
nor U22676 (N_22676,N_22167,N_22438);
xnor U22677 (N_22677,N_22155,N_22026);
or U22678 (N_22678,N_22072,N_22274);
nor U22679 (N_22679,N_22025,N_22344);
and U22680 (N_22680,N_22375,N_22098);
nand U22681 (N_22681,N_22286,N_22092);
or U22682 (N_22682,N_22383,N_22300);
or U22683 (N_22683,N_22122,N_22197);
xnor U22684 (N_22684,N_22121,N_22297);
xor U22685 (N_22685,N_22027,N_22202);
and U22686 (N_22686,N_22499,N_22299);
nand U22687 (N_22687,N_22350,N_22089);
nor U22688 (N_22688,N_22263,N_22302);
xor U22689 (N_22689,N_22131,N_22029);
xnor U22690 (N_22690,N_22132,N_22358);
or U22691 (N_22691,N_22107,N_22241);
nor U22692 (N_22692,N_22310,N_22445);
nand U22693 (N_22693,N_22095,N_22295);
and U22694 (N_22694,N_22484,N_22215);
nand U22695 (N_22695,N_22292,N_22210);
nor U22696 (N_22696,N_22147,N_22400);
nor U22697 (N_22697,N_22497,N_22077);
and U22698 (N_22698,N_22129,N_22401);
xor U22699 (N_22699,N_22018,N_22479);
nor U22700 (N_22700,N_22304,N_22090);
and U22701 (N_22701,N_22052,N_22398);
nand U22702 (N_22702,N_22073,N_22271);
nor U22703 (N_22703,N_22108,N_22204);
xor U22704 (N_22704,N_22255,N_22260);
and U22705 (N_22705,N_22322,N_22024);
nor U22706 (N_22706,N_22103,N_22174);
nor U22707 (N_22707,N_22117,N_22407);
xnor U22708 (N_22708,N_22415,N_22420);
nand U22709 (N_22709,N_22219,N_22067);
nor U22710 (N_22710,N_22043,N_22172);
or U22711 (N_22711,N_22422,N_22220);
nor U22712 (N_22712,N_22315,N_22065);
nor U22713 (N_22713,N_22492,N_22164);
nand U22714 (N_22714,N_22120,N_22456);
nor U22715 (N_22715,N_22074,N_22218);
xnor U22716 (N_22716,N_22229,N_22402);
nor U22717 (N_22717,N_22475,N_22273);
or U22718 (N_22718,N_22079,N_22305);
nand U22719 (N_22719,N_22446,N_22110);
xnor U22720 (N_22720,N_22460,N_22343);
xnor U22721 (N_22721,N_22115,N_22145);
and U22722 (N_22722,N_22134,N_22309);
and U22723 (N_22723,N_22423,N_22314);
nand U22724 (N_22724,N_22483,N_22480);
nor U22725 (N_22725,N_22057,N_22258);
nor U22726 (N_22726,N_22186,N_22275);
nor U22727 (N_22727,N_22144,N_22033);
or U22728 (N_22728,N_22437,N_22105);
nand U22729 (N_22729,N_22325,N_22221);
nor U22730 (N_22730,N_22250,N_22064);
xor U22731 (N_22731,N_22182,N_22293);
and U22732 (N_22732,N_22209,N_22180);
nand U22733 (N_22733,N_22200,N_22265);
xnor U22734 (N_22734,N_22047,N_22272);
and U22735 (N_22735,N_22352,N_22361);
xor U22736 (N_22736,N_22450,N_22211);
xor U22737 (N_22737,N_22020,N_22022);
nor U22738 (N_22738,N_22439,N_22362);
or U22739 (N_22739,N_22363,N_22403);
nand U22740 (N_22740,N_22329,N_22191);
xnor U22741 (N_22741,N_22168,N_22385);
nand U22742 (N_22742,N_22417,N_22468);
nand U22743 (N_22743,N_22207,N_22256);
nand U22744 (N_22744,N_22248,N_22395);
nand U22745 (N_22745,N_22443,N_22323);
xor U22746 (N_22746,N_22235,N_22223);
and U22747 (N_22747,N_22364,N_22496);
nand U22748 (N_22748,N_22488,N_22059);
and U22749 (N_22749,N_22294,N_22341);
nand U22750 (N_22750,N_22480,N_22150);
and U22751 (N_22751,N_22164,N_22220);
or U22752 (N_22752,N_22023,N_22178);
or U22753 (N_22753,N_22081,N_22115);
nand U22754 (N_22754,N_22257,N_22237);
nand U22755 (N_22755,N_22217,N_22427);
and U22756 (N_22756,N_22192,N_22037);
nand U22757 (N_22757,N_22209,N_22426);
xor U22758 (N_22758,N_22308,N_22111);
nand U22759 (N_22759,N_22034,N_22245);
nor U22760 (N_22760,N_22085,N_22262);
nand U22761 (N_22761,N_22460,N_22486);
nand U22762 (N_22762,N_22216,N_22051);
or U22763 (N_22763,N_22346,N_22393);
and U22764 (N_22764,N_22222,N_22098);
or U22765 (N_22765,N_22118,N_22396);
or U22766 (N_22766,N_22165,N_22464);
nand U22767 (N_22767,N_22476,N_22100);
and U22768 (N_22768,N_22206,N_22021);
xnor U22769 (N_22769,N_22288,N_22485);
nand U22770 (N_22770,N_22284,N_22406);
and U22771 (N_22771,N_22401,N_22221);
and U22772 (N_22772,N_22319,N_22069);
nor U22773 (N_22773,N_22128,N_22285);
nor U22774 (N_22774,N_22093,N_22023);
nand U22775 (N_22775,N_22438,N_22036);
nand U22776 (N_22776,N_22000,N_22464);
xor U22777 (N_22777,N_22247,N_22352);
nand U22778 (N_22778,N_22264,N_22109);
nand U22779 (N_22779,N_22303,N_22089);
xor U22780 (N_22780,N_22356,N_22437);
nor U22781 (N_22781,N_22227,N_22040);
nor U22782 (N_22782,N_22346,N_22193);
and U22783 (N_22783,N_22010,N_22042);
nor U22784 (N_22784,N_22343,N_22064);
or U22785 (N_22785,N_22368,N_22423);
xor U22786 (N_22786,N_22236,N_22154);
nand U22787 (N_22787,N_22041,N_22373);
and U22788 (N_22788,N_22102,N_22174);
nand U22789 (N_22789,N_22324,N_22053);
nor U22790 (N_22790,N_22414,N_22259);
xnor U22791 (N_22791,N_22405,N_22129);
nor U22792 (N_22792,N_22423,N_22202);
nand U22793 (N_22793,N_22281,N_22073);
nor U22794 (N_22794,N_22184,N_22168);
nand U22795 (N_22795,N_22066,N_22489);
xor U22796 (N_22796,N_22418,N_22482);
nand U22797 (N_22797,N_22453,N_22460);
nor U22798 (N_22798,N_22258,N_22382);
or U22799 (N_22799,N_22029,N_22484);
or U22800 (N_22800,N_22301,N_22364);
nor U22801 (N_22801,N_22368,N_22474);
and U22802 (N_22802,N_22418,N_22190);
nand U22803 (N_22803,N_22440,N_22123);
nand U22804 (N_22804,N_22487,N_22268);
xor U22805 (N_22805,N_22248,N_22442);
nor U22806 (N_22806,N_22123,N_22226);
xnor U22807 (N_22807,N_22288,N_22483);
or U22808 (N_22808,N_22099,N_22472);
xnor U22809 (N_22809,N_22073,N_22294);
xnor U22810 (N_22810,N_22412,N_22483);
and U22811 (N_22811,N_22439,N_22126);
xnor U22812 (N_22812,N_22113,N_22438);
xor U22813 (N_22813,N_22148,N_22015);
and U22814 (N_22814,N_22242,N_22113);
nor U22815 (N_22815,N_22218,N_22287);
and U22816 (N_22816,N_22348,N_22137);
and U22817 (N_22817,N_22449,N_22199);
or U22818 (N_22818,N_22448,N_22379);
and U22819 (N_22819,N_22057,N_22354);
nand U22820 (N_22820,N_22243,N_22479);
xor U22821 (N_22821,N_22238,N_22270);
and U22822 (N_22822,N_22397,N_22209);
xnor U22823 (N_22823,N_22048,N_22159);
and U22824 (N_22824,N_22455,N_22328);
nand U22825 (N_22825,N_22087,N_22438);
or U22826 (N_22826,N_22064,N_22358);
or U22827 (N_22827,N_22094,N_22475);
xor U22828 (N_22828,N_22293,N_22317);
and U22829 (N_22829,N_22147,N_22027);
nand U22830 (N_22830,N_22334,N_22281);
nand U22831 (N_22831,N_22323,N_22134);
and U22832 (N_22832,N_22372,N_22322);
nor U22833 (N_22833,N_22257,N_22320);
nor U22834 (N_22834,N_22251,N_22100);
and U22835 (N_22835,N_22485,N_22050);
nor U22836 (N_22836,N_22099,N_22142);
nor U22837 (N_22837,N_22035,N_22495);
or U22838 (N_22838,N_22039,N_22242);
nor U22839 (N_22839,N_22486,N_22376);
nand U22840 (N_22840,N_22401,N_22229);
xor U22841 (N_22841,N_22118,N_22131);
nand U22842 (N_22842,N_22128,N_22057);
and U22843 (N_22843,N_22305,N_22240);
nor U22844 (N_22844,N_22008,N_22042);
xor U22845 (N_22845,N_22345,N_22389);
xnor U22846 (N_22846,N_22476,N_22394);
or U22847 (N_22847,N_22310,N_22316);
xnor U22848 (N_22848,N_22401,N_22374);
nand U22849 (N_22849,N_22358,N_22429);
nor U22850 (N_22850,N_22271,N_22163);
nand U22851 (N_22851,N_22341,N_22329);
nand U22852 (N_22852,N_22342,N_22203);
and U22853 (N_22853,N_22361,N_22310);
xnor U22854 (N_22854,N_22247,N_22478);
nor U22855 (N_22855,N_22096,N_22066);
xnor U22856 (N_22856,N_22320,N_22180);
and U22857 (N_22857,N_22441,N_22052);
and U22858 (N_22858,N_22023,N_22051);
or U22859 (N_22859,N_22124,N_22411);
nand U22860 (N_22860,N_22438,N_22094);
and U22861 (N_22861,N_22345,N_22079);
nand U22862 (N_22862,N_22335,N_22002);
and U22863 (N_22863,N_22398,N_22219);
and U22864 (N_22864,N_22188,N_22036);
xnor U22865 (N_22865,N_22356,N_22222);
or U22866 (N_22866,N_22357,N_22487);
xnor U22867 (N_22867,N_22125,N_22466);
or U22868 (N_22868,N_22194,N_22020);
or U22869 (N_22869,N_22498,N_22003);
nor U22870 (N_22870,N_22127,N_22270);
nor U22871 (N_22871,N_22378,N_22407);
nand U22872 (N_22872,N_22402,N_22116);
or U22873 (N_22873,N_22175,N_22052);
and U22874 (N_22874,N_22263,N_22348);
nand U22875 (N_22875,N_22169,N_22329);
xnor U22876 (N_22876,N_22231,N_22441);
nand U22877 (N_22877,N_22163,N_22089);
xor U22878 (N_22878,N_22042,N_22120);
nor U22879 (N_22879,N_22097,N_22380);
or U22880 (N_22880,N_22066,N_22128);
nor U22881 (N_22881,N_22491,N_22171);
nor U22882 (N_22882,N_22020,N_22001);
or U22883 (N_22883,N_22278,N_22326);
nor U22884 (N_22884,N_22475,N_22137);
nor U22885 (N_22885,N_22479,N_22180);
and U22886 (N_22886,N_22153,N_22219);
nand U22887 (N_22887,N_22316,N_22470);
or U22888 (N_22888,N_22469,N_22083);
nor U22889 (N_22889,N_22460,N_22235);
xor U22890 (N_22890,N_22000,N_22498);
and U22891 (N_22891,N_22361,N_22258);
nor U22892 (N_22892,N_22176,N_22308);
xnor U22893 (N_22893,N_22401,N_22277);
and U22894 (N_22894,N_22334,N_22291);
xor U22895 (N_22895,N_22224,N_22248);
nor U22896 (N_22896,N_22493,N_22398);
and U22897 (N_22897,N_22490,N_22416);
nand U22898 (N_22898,N_22177,N_22482);
nand U22899 (N_22899,N_22394,N_22237);
or U22900 (N_22900,N_22482,N_22408);
nor U22901 (N_22901,N_22009,N_22123);
xnor U22902 (N_22902,N_22373,N_22389);
and U22903 (N_22903,N_22368,N_22301);
nand U22904 (N_22904,N_22031,N_22137);
xnor U22905 (N_22905,N_22195,N_22357);
xnor U22906 (N_22906,N_22407,N_22160);
nand U22907 (N_22907,N_22379,N_22484);
nand U22908 (N_22908,N_22401,N_22413);
nor U22909 (N_22909,N_22484,N_22214);
nor U22910 (N_22910,N_22129,N_22375);
nor U22911 (N_22911,N_22144,N_22081);
nand U22912 (N_22912,N_22341,N_22029);
nor U22913 (N_22913,N_22242,N_22160);
or U22914 (N_22914,N_22428,N_22414);
and U22915 (N_22915,N_22421,N_22022);
nor U22916 (N_22916,N_22483,N_22382);
nor U22917 (N_22917,N_22358,N_22180);
and U22918 (N_22918,N_22060,N_22169);
xor U22919 (N_22919,N_22133,N_22052);
or U22920 (N_22920,N_22002,N_22063);
or U22921 (N_22921,N_22396,N_22476);
or U22922 (N_22922,N_22372,N_22189);
nand U22923 (N_22923,N_22227,N_22342);
or U22924 (N_22924,N_22008,N_22445);
and U22925 (N_22925,N_22038,N_22070);
xor U22926 (N_22926,N_22191,N_22474);
nor U22927 (N_22927,N_22442,N_22062);
xnor U22928 (N_22928,N_22325,N_22435);
xnor U22929 (N_22929,N_22242,N_22444);
xnor U22930 (N_22930,N_22119,N_22101);
nor U22931 (N_22931,N_22119,N_22059);
and U22932 (N_22932,N_22011,N_22384);
nand U22933 (N_22933,N_22094,N_22465);
or U22934 (N_22934,N_22299,N_22388);
or U22935 (N_22935,N_22027,N_22353);
or U22936 (N_22936,N_22257,N_22206);
nand U22937 (N_22937,N_22281,N_22061);
nor U22938 (N_22938,N_22168,N_22196);
xnor U22939 (N_22939,N_22224,N_22424);
xnor U22940 (N_22940,N_22002,N_22352);
xor U22941 (N_22941,N_22091,N_22169);
nor U22942 (N_22942,N_22400,N_22044);
nor U22943 (N_22943,N_22138,N_22250);
or U22944 (N_22944,N_22085,N_22008);
and U22945 (N_22945,N_22046,N_22117);
nand U22946 (N_22946,N_22374,N_22341);
or U22947 (N_22947,N_22231,N_22413);
xor U22948 (N_22948,N_22208,N_22011);
nand U22949 (N_22949,N_22104,N_22333);
nand U22950 (N_22950,N_22110,N_22163);
xor U22951 (N_22951,N_22414,N_22232);
xor U22952 (N_22952,N_22439,N_22360);
and U22953 (N_22953,N_22190,N_22319);
or U22954 (N_22954,N_22321,N_22280);
xnor U22955 (N_22955,N_22226,N_22272);
or U22956 (N_22956,N_22271,N_22260);
nor U22957 (N_22957,N_22128,N_22326);
nand U22958 (N_22958,N_22180,N_22032);
or U22959 (N_22959,N_22196,N_22405);
xor U22960 (N_22960,N_22068,N_22248);
or U22961 (N_22961,N_22332,N_22331);
nor U22962 (N_22962,N_22262,N_22239);
or U22963 (N_22963,N_22476,N_22387);
or U22964 (N_22964,N_22141,N_22092);
nor U22965 (N_22965,N_22302,N_22477);
nand U22966 (N_22966,N_22492,N_22452);
xor U22967 (N_22967,N_22216,N_22122);
and U22968 (N_22968,N_22298,N_22073);
and U22969 (N_22969,N_22101,N_22066);
or U22970 (N_22970,N_22340,N_22427);
nand U22971 (N_22971,N_22198,N_22226);
xnor U22972 (N_22972,N_22394,N_22463);
nor U22973 (N_22973,N_22298,N_22283);
nand U22974 (N_22974,N_22488,N_22258);
nor U22975 (N_22975,N_22211,N_22468);
and U22976 (N_22976,N_22098,N_22115);
and U22977 (N_22977,N_22192,N_22141);
nand U22978 (N_22978,N_22252,N_22256);
nor U22979 (N_22979,N_22411,N_22033);
and U22980 (N_22980,N_22386,N_22320);
xnor U22981 (N_22981,N_22413,N_22206);
nor U22982 (N_22982,N_22275,N_22375);
nand U22983 (N_22983,N_22315,N_22264);
and U22984 (N_22984,N_22456,N_22208);
or U22985 (N_22985,N_22089,N_22227);
or U22986 (N_22986,N_22475,N_22353);
nand U22987 (N_22987,N_22082,N_22283);
nor U22988 (N_22988,N_22398,N_22266);
nand U22989 (N_22989,N_22035,N_22353);
xnor U22990 (N_22990,N_22062,N_22176);
nor U22991 (N_22991,N_22207,N_22402);
or U22992 (N_22992,N_22203,N_22241);
xnor U22993 (N_22993,N_22288,N_22077);
nand U22994 (N_22994,N_22289,N_22290);
and U22995 (N_22995,N_22430,N_22250);
nand U22996 (N_22996,N_22263,N_22369);
or U22997 (N_22997,N_22067,N_22374);
and U22998 (N_22998,N_22031,N_22047);
nor U22999 (N_22999,N_22495,N_22082);
or U23000 (N_23000,N_22694,N_22716);
and U23001 (N_23001,N_22921,N_22788);
xor U23002 (N_23002,N_22608,N_22665);
nor U23003 (N_23003,N_22505,N_22658);
nand U23004 (N_23004,N_22832,N_22689);
xor U23005 (N_23005,N_22939,N_22666);
nor U23006 (N_23006,N_22806,N_22985);
xnor U23007 (N_23007,N_22710,N_22873);
and U23008 (N_23008,N_22834,N_22726);
nand U23009 (N_23009,N_22643,N_22762);
nor U23010 (N_23010,N_22894,N_22769);
xnor U23011 (N_23011,N_22979,N_22811);
xor U23012 (N_23012,N_22838,N_22548);
nand U23013 (N_23013,N_22787,N_22882);
nand U23014 (N_23014,N_22656,N_22872);
nor U23015 (N_23015,N_22594,N_22853);
nor U23016 (N_23016,N_22518,N_22639);
xnor U23017 (N_23017,N_22720,N_22786);
and U23018 (N_23018,N_22622,N_22630);
xnor U23019 (N_23019,N_22502,N_22708);
nor U23020 (N_23020,N_22699,N_22794);
or U23021 (N_23021,N_22755,N_22839);
nor U23022 (N_23022,N_22638,N_22581);
or U23023 (N_23023,N_22856,N_22766);
and U23024 (N_23024,N_22750,N_22655);
and U23025 (N_23025,N_22947,N_22893);
or U23026 (N_23026,N_22702,N_22761);
xnor U23027 (N_23027,N_22628,N_22956);
xnor U23028 (N_23028,N_22654,N_22558);
nand U23029 (N_23029,N_22513,N_22852);
and U23030 (N_23030,N_22529,N_22718);
nor U23031 (N_23031,N_22841,N_22751);
or U23032 (N_23032,N_22791,N_22728);
nand U23033 (N_23033,N_22647,N_22908);
xnor U23034 (N_23034,N_22779,N_22793);
nand U23035 (N_23035,N_22919,N_22538);
xor U23036 (N_23036,N_22936,N_22542);
and U23037 (N_23037,N_22596,N_22574);
nor U23038 (N_23038,N_22583,N_22764);
or U23039 (N_23039,N_22900,N_22732);
or U23040 (N_23040,N_22822,N_22920);
or U23041 (N_23041,N_22661,N_22990);
xnor U23042 (N_23042,N_22859,N_22589);
xnor U23043 (N_23043,N_22773,N_22931);
nand U23044 (N_23044,N_22996,N_22911);
nand U23045 (N_23045,N_22831,N_22539);
nand U23046 (N_23046,N_22560,N_22901);
or U23047 (N_23047,N_22714,N_22753);
xor U23048 (N_23048,N_22519,N_22818);
or U23049 (N_23049,N_22933,N_22632);
xnor U23050 (N_23050,N_22826,N_22633);
or U23051 (N_23051,N_22734,N_22587);
or U23052 (N_23052,N_22974,N_22951);
or U23053 (N_23053,N_22557,N_22846);
nor U23054 (N_23054,N_22625,N_22544);
nor U23055 (N_23055,N_22902,N_22892);
xnor U23056 (N_23056,N_22799,N_22644);
nor U23057 (N_23057,N_22566,N_22515);
and U23058 (N_23058,N_22964,N_22783);
and U23059 (N_23059,N_22845,N_22877);
nand U23060 (N_23060,N_22657,N_22789);
nor U23061 (N_23061,N_22819,N_22646);
nor U23062 (N_23062,N_22676,N_22512);
and U23063 (N_23063,N_22631,N_22813);
xor U23064 (N_23064,N_22526,N_22912);
xnor U23065 (N_23065,N_22627,N_22567);
xnor U23066 (N_23066,N_22994,N_22896);
xor U23067 (N_23067,N_22705,N_22562);
and U23068 (N_23068,N_22966,N_22770);
and U23069 (N_23069,N_22747,N_22508);
nor U23070 (N_23070,N_22506,N_22550);
xor U23071 (N_23071,N_22805,N_22615);
nand U23072 (N_23072,N_22855,N_22815);
nor U23073 (N_23073,N_22523,N_22532);
nand U23074 (N_23074,N_22723,N_22642);
and U23075 (N_23075,N_22667,N_22800);
xnor U23076 (N_23076,N_22686,N_22565);
nor U23077 (N_23077,N_22944,N_22778);
nor U23078 (N_23078,N_22934,N_22978);
and U23079 (N_23079,N_22520,N_22537);
xnor U23080 (N_23080,N_22678,N_22957);
nand U23081 (N_23081,N_22953,N_22555);
nor U23082 (N_23082,N_22807,N_22975);
nor U23083 (N_23083,N_22521,N_22850);
nor U23084 (N_23084,N_22591,N_22878);
nor U23085 (N_23085,N_22942,N_22925);
nand U23086 (N_23086,N_22932,N_22808);
nand U23087 (N_23087,N_22854,N_22918);
xnor U23088 (N_23088,N_22849,N_22823);
xor U23089 (N_23089,N_22559,N_22943);
xor U23090 (N_23090,N_22669,N_22692);
nor U23091 (N_23091,N_22814,N_22593);
or U23092 (N_23092,N_22636,N_22829);
nor U23093 (N_23093,N_22758,N_22679);
xnor U23094 (N_23094,N_22745,N_22511);
nand U23095 (N_23095,N_22879,N_22713);
nor U23096 (N_23096,N_22570,N_22672);
nor U23097 (N_23097,N_22835,N_22775);
and U23098 (N_23098,N_22662,N_22746);
or U23099 (N_23099,N_22968,N_22917);
nand U23100 (N_23100,N_22916,N_22701);
and U23101 (N_23101,N_22564,N_22561);
and U23102 (N_23102,N_22599,N_22965);
xnor U23103 (N_23103,N_22578,N_22743);
nand U23104 (N_23104,N_22610,N_22652);
xor U23105 (N_23105,N_22637,N_22906);
and U23106 (N_23106,N_22533,N_22851);
nand U23107 (N_23107,N_22759,N_22929);
xor U23108 (N_23108,N_22740,N_22576);
nand U23109 (N_23109,N_22884,N_22527);
xor U23110 (N_23110,N_22602,N_22735);
nor U23111 (N_23111,N_22954,N_22618);
xor U23112 (N_23112,N_22897,N_22992);
xnor U23113 (N_23113,N_22691,N_22827);
xnor U23114 (N_23114,N_22650,N_22863);
nor U23115 (N_23115,N_22660,N_22771);
or U23116 (N_23116,N_22757,N_22999);
or U23117 (N_23117,N_22712,N_22952);
nor U23118 (N_23118,N_22802,N_22648);
nor U23119 (N_23119,N_22619,N_22704);
xnor U23120 (N_23120,N_22817,N_22821);
or U23121 (N_23121,N_22828,N_22510);
nor U23122 (N_23122,N_22895,N_22541);
nand U23123 (N_23123,N_22795,N_22616);
and U23124 (N_23124,N_22858,N_22626);
or U23125 (N_23125,N_22780,N_22812);
and U23126 (N_23126,N_22962,N_22698);
nor U23127 (N_23127,N_22963,N_22703);
and U23128 (N_23128,N_22837,N_22913);
nor U23129 (N_23129,N_22717,N_22781);
nor U23130 (N_23130,N_22514,N_22722);
nand U23131 (N_23131,N_22867,N_22641);
xor U23132 (N_23132,N_22848,N_22977);
and U23133 (N_23133,N_22898,N_22733);
nand U23134 (N_23134,N_22986,N_22836);
xor U23135 (N_23135,N_22634,N_22959);
nand U23136 (N_23136,N_22792,N_22765);
and U23137 (N_23137,N_22534,N_22971);
xnor U23138 (N_23138,N_22991,N_22603);
nand U23139 (N_23139,N_22531,N_22605);
xnor U23140 (N_23140,N_22730,N_22801);
nand U23141 (N_23141,N_22960,N_22798);
or U23142 (N_23142,N_22707,N_22530);
xnor U23143 (N_23143,N_22680,N_22993);
nand U23144 (N_23144,N_22535,N_22609);
nor U23145 (N_23145,N_22958,N_22653);
nand U23146 (N_23146,N_22763,N_22946);
and U23147 (N_23147,N_22972,N_22738);
or U23148 (N_23148,N_22937,N_22681);
nand U23149 (N_23149,N_22905,N_22597);
xor U23150 (N_23150,N_22592,N_22997);
or U23151 (N_23151,N_22973,N_22736);
nor U23152 (N_23152,N_22899,N_22804);
or U23153 (N_23153,N_22737,N_22961);
or U23154 (N_23154,N_22928,N_22674);
nor U23155 (N_23155,N_22843,N_22553);
or U23156 (N_23156,N_22888,N_22989);
or U23157 (N_23157,N_22768,N_22987);
or U23158 (N_23158,N_22721,N_22741);
or U23159 (N_23159,N_22682,N_22824);
and U23160 (N_23160,N_22725,N_22865);
nand U23161 (N_23161,N_22784,N_22607);
nor U23162 (N_23162,N_22885,N_22549);
xor U23163 (N_23163,N_22938,N_22777);
and U23164 (N_23164,N_22909,N_22910);
nand U23165 (N_23165,N_22744,N_22543);
xnor U23166 (N_23166,N_22904,N_22577);
xor U23167 (N_23167,N_22677,N_22890);
nand U23168 (N_23168,N_22673,N_22575);
nand U23169 (N_23169,N_22860,N_22955);
or U23170 (N_23170,N_22983,N_22687);
xnor U23171 (N_23171,N_22606,N_22926);
nand U23172 (N_23172,N_22748,N_22797);
xor U23173 (N_23173,N_22785,N_22727);
or U23174 (N_23174,N_22940,N_22825);
nand U23175 (N_23175,N_22923,N_22924);
xnor U23176 (N_23176,N_22949,N_22772);
and U23177 (N_23177,N_22668,N_22640);
xnor U23178 (N_23178,N_22585,N_22528);
or U23179 (N_23179,N_22945,N_22871);
xor U23180 (N_23180,N_22590,N_22715);
xor U23181 (N_23181,N_22941,N_22995);
or U23182 (N_23182,N_22980,N_22988);
or U23183 (N_23183,N_22907,N_22790);
xor U23184 (N_23184,N_22545,N_22803);
or U23185 (N_23185,N_22588,N_22711);
nor U23186 (N_23186,N_22922,N_22840);
xor U23187 (N_23187,N_22820,N_22731);
xnor U23188 (N_23188,N_22614,N_22579);
nor U23189 (N_23189,N_22684,N_22875);
and U23190 (N_23190,N_22876,N_22927);
xor U23191 (N_23191,N_22967,N_22861);
nor U23192 (N_23192,N_22675,N_22649);
and U23193 (N_23193,N_22970,N_22883);
xnor U23194 (N_23194,N_22580,N_22729);
and U23195 (N_23195,N_22874,N_22930);
xnor U23196 (N_23196,N_22584,N_22754);
nor U23197 (N_23197,N_22645,N_22500);
and U23198 (N_23198,N_22948,N_22551);
nand U23199 (N_23199,N_22774,N_22889);
nor U23200 (N_23200,N_22671,N_22796);
and U23201 (N_23201,N_22696,N_22864);
nand U23202 (N_23202,N_22891,N_22914);
nand U23203 (N_23203,N_22546,N_22572);
xnor U23204 (N_23204,N_22695,N_22776);
or U23205 (N_23205,N_22868,N_22880);
nor U23206 (N_23206,N_22620,N_22767);
nor U23207 (N_23207,N_22659,N_22844);
nand U23208 (N_23208,N_22709,N_22552);
nor U23209 (N_23209,N_22866,N_22582);
nand U23210 (N_23210,N_22816,N_22915);
nor U23211 (N_23211,N_22756,N_22516);
nor U23212 (N_23212,N_22700,N_22664);
nand U23213 (N_23213,N_22611,N_22569);
nor U23214 (N_23214,N_22501,N_22683);
xor U23215 (N_23215,N_22556,N_22685);
nor U23216 (N_23216,N_22624,N_22706);
nand U23217 (N_23217,N_22598,N_22719);
nand U23218 (N_23218,N_22604,N_22749);
or U23219 (N_23219,N_22830,N_22935);
xnor U23220 (N_23220,N_22629,N_22623);
nor U23221 (N_23221,N_22870,N_22547);
xnor U23222 (N_23222,N_22503,N_22507);
nor U23223 (N_23223,N_22670,N_22524);
nand U23224 (N_23224,N_22842,N_22571);
or U23225 (N_23225,N_22862,N_22847);
xnor U23226 (N_23226,N_22554,N_22976);
and U23227 (N_23227,N_22886,N_22950);
xnor U23228 (N_23228,N_22568,N_22663);
or U23229 (N_23229,N_22810,N_22525);
nor U23230 (N_23230,N_22509,N_22981);
nand U23231 (N_23231,N_22688,N_22739);
and U23232 (N_23232,N_22612,N_22617);
nand U23233 (N_23233,N_22613,N_22690);
xnor U23234 (N_23234,N_22522,N_22724);
and U23235 (N_23235,N_22651,N_22998);
xor U23236 (N_23236,N_22969,N_22517);
or U23237 (N_23237,N_22693,N_22601);
nor U23238 (N_23238,N_22573,N_22504);
and U23239 (N_23239,N_22984,N_22540);
nor U23240 (N_23240,N_22982,N_22857);
xnor U23241 (N_23241,N_22595,N_22621);
nor U23242 (N_23242,N_22869,N_22809);
xor U23243 (N_23243,N_22600,N_22887);
or U23244 (N_23244,N_22742,N_22635);
or U23245 (N_23245,N_22752,N_22782);
nor U23246 (N_23246,N_22536,N_22697);
xor U23247 (N_23247,N_22833,N_22760);
nand U23248 (N_23248,N_22881,N_22563);
nand U23249 (N_23249,N_22586,N_22903);
nand U23250 (N_23250,N_22971,N_22519);
and U23251 (N_23251,N_22613,N_22799);
and U23252 (N_23252,N_22680,N_22900);
and U23253 (N_23253,N_22992,N_22670);
nor U23254 (N_23254,N_22513,N_22544);
and U23255 (N_23255,N_22976,N_22857);
xnor U23256 (N_23256,N_22593,N_22886);
xnor U23257 (N_23257,N_22814,N_22606);
nor U23258 (N_23258,N_22742,N_22773);
or U23259 (N_23259,N_22815,N_22936);
and U23260 (N_23260,N_22838,N_22839);
and U23261 (N_23261,N_22904,N_22989);
xnor U23262 (N_23262,N_22998,N_22531);
nor U23263 (N_23263,N_22859,N_22844);
or U23264 (N_23264,N_22576,N_22536);
or U23265 (N_23265,N_22808,N_22575);
nand U23266 (N_23266,N_22818,N_22641);
or U23267 (N_23267,N_22727,N_22590);
nor U23268 (N_23268,N_22581,N_22577);
nor U23269 (N_23269,N_22963,N_22718);
or U23270 (N_23270,N_22582,N_22542);
nand U23271 (N_23271,N_22947,N_22716);
or U23272 (N_23272,N_22521,N_22846);
or U23273 (N_23273,N_22902,N_22815);
nand U23274 (N_23274,N_22946,N_22708);
or U23275 (N_23275,N_22835,N_22731);
or U23276 (N_23276,N_22676,N_22819);
nor U23277 (N_23277,N_22502,N_22751);
nor U23278 (N_23278,N_22962,N_22563);
nand U23279 (N_23279,N_22819,N_22756);
nor U23280 (N_23280,N_22580,N_22627);
nand U23281 (N_23281,N_22989,N_22998);
or U23282 (N_23282,N_22825,N_22767);
and U23283 (N_23283,N_22618,N_22662);
or U23284 (N_23284,N_22984,N_22516);
nor U23285 (N_23285,N_22718,N_22510);
nor U23286 (N_23286,N_22941,N_22631);
xnor U23287 (N_23287,N_22790,N_22973);
and U23288 (N_23288,N_22774,N_22831);
or U23289 (N_23289,N_22942,N_22747);
nand U23290 (N_23290,N_22738,N_22980);
and U23291 (N_23291,N_22752,N_22651);
nand U23292 (N_23292,N_22687,N_22623);
nor U23293 (N_23293,N_22647,N_22976);
xnor U23294 (N_23294,N_22991,N_22614);
nor U23295 (N_23295,N_22837,N_22849);
xnor U23296 (N_23296,N_22898,N_22878);
xnor U23297 (N_23297,N_22928,N_22586);
or U23298 (N_23298,N_22991,N_22907);
xor U23299 (N_23299,N_22617,N_22902);
nand U23300 (N_23300,N_22748,N_22877);
and U23301 (N_23301,N_22626,N_22739);
nor U23302 (N_23302,N_22937,N_22799);
or U23303 (N_23303,N_22653,N_22752);
nand U23304 (N_23304,N_22857,N_22556);
or U23305 (N_23305,N_22919,N_22630);
xnor U23306 (N_23306,N_22780,N_22536);
xnor U23307 (N_23307,N_22741,N_22892);
and U23308 (N_23308,N_22802,N_22587);
nand U23309 (N_23309,N_22822,N_22890);
xor U23310 (N_23310,N_22749,N_22847);
xnor U23311 (N_23311,N_22676,N_22960);
nor U23312 (N_23312,N_22821,N_22543);
nand U23313 (N_23313,N_22508,N_22985);
and U23314 (N_23314,N_22665,N_22727);
xor U23315 (N_23315,N_22680,N_22891);
xnor U23316 (N_23316,N_22886,N_22584);
or U23317 (N_23317,N_22774,N_22612);
xnor U23318 (N_23318,N_22878,N_22851);
nand U23319 (N_23319,N_22869,N_22659);
nand U23320 (N_23320,N_22659,N_22705);
and U23321 (N_23321,N_22582,N_22726);
or U23322 (N_23322,N_22965,N_22912);
or U23323 (N_23323,N_22945,N_22803);
nor U23324 (N_23324,N_22866,N_22642);
nand U23325 (N_23325,N_22543,N_22951);
and U23326 (N_23326,N_22508,N_22858);
nor U23327 (N_23327,N_22698,N_22586);
and U23328 (N_23328,N_22904,N_22670);
and U23329 (N_23329,N_22639,N_22700);
or U23330 (N_23330,N_22798,N_22708);
and U23331 (N_23331,N_22562,N_22524);
or U23332 (N_23332,N_22792,N_22997);
xor U23333 (N_23333,N_22659,N_22874);
and U23334 (N_23334,N_22962,N_22794);
and U23335 (N_23335,N_22855,N_22771);
nand U23336 (N_23336,N_22851,N_22933);
and U23337 (N_23337,N_22835,N_22858);
nand U23338 (N_23338,N_22740,N_22590);
nand U23339 (N_23339,N_22674,N_22807);
nor U23340 (N_23340,N_22558,N_22832);
xnor U23341 (N_23341,N_22897,N_22840);
nand U23342 (N_23342,N_22965,N_22791);
or U23343 (N_23343,N_22847,N_22835);
or U23344 (N_23344,N_22562,N_22568);
or U23345 (N_23345,N_22887,N_22664);
or U23346 (N_23346,N_22634,N_22898);
nand U23347 (N_23347,N_22579,N_22702);
or U23348 (N_23348,N_22813,N_22686);
or U23349 (N_23349,N_22679,N_22518);
xor U23350 (N_23350,N_22747,N_22518);
xor U23351 (N_23351,N_22585,N_22504);
or U23352 (N_23352,N_22807,N_22737);
and U23353 (N_23353,N_22820,N_22978);
xnor U23354 (N_23354,N_22597,N_22841);
nor U23355 (N_23355,N_22680,N_22911);
or U23356 (N_23356,N_22789,N_22533);
or U23357 (N_23357,N_22546,N_22636);
or U23358 (N_23358,N_22933,N_22713);
or U23359 (N_23359,N_22942,N_22721);
nand U23360 (N_23360,N_22540,N_22585);
nor U23361 (N_23361,N_22840,N_22873);
xor U23362 (N_23362,N_22652,N_22695);
xor U23363 (N_23363,N_22738,N_22958);
xnor U23364 (N_23364,N_22768,N_22594);
or U23365 (N_23365,N_22977,N_22980);
or U23366 (N_23366,N_22984,N_22773);
and U23367 (N_23367,N_22718,N_22989);
nand U23368 (N_23368,N_22990,N_22978);
nor U23369 (N_23369,N_22993,N_22685);
nor U23370 (N_23370,N_22797,N_22928);
or U23371 (N_23371,N_22775,N_22719);
nand U23372 (N_23372,N_22506,N_22562);
and U23373 (N_23373,N_22721,N_22924);
or U23374 (N_23374,N_22598,N_22996);
and U23375 (N_23375,N_22538,N_22858);
and U23376 (N_23376,N_22793,N_22692);
xnor U23377 (N_23377,N_22796,N_22988);
and U23378 (N_23378,N_22952,N_22646);
or U23379 (N_23379,N_22897,N_22874);
xnor U23380 (N_23380,N_22543,N_22628);
and U23381 (N_23381,N_22757,N_22602);
nand U23382 (N_23382,N_22647,N_22808);
and U23383 (N_23383,N_22650,N_22893);
or U23384 (N_23384,N_22727,N_22972);
and U23385 (N_23385,N_22750,N_22795);
xnor U23386 (N_23386,N_22608,N_22793);
nand U23387 (N_23387,N_22615,N_22528);
xnor U23388 (N_23388,N_22774,N_22993);
or U23389 (N_23389,N_22576,N_22544);
xnor U23390 (N_23390,N_22587,N_22867);
xor U23391 (N_23391,N_22700,N_22747);
and U23392 (N_23392,N_22844,N_22917);
nand U23393 (N_23393,N_22829,N_22720);
nand U23394 (N_23394,N_22789,N_22574);
or U23395 (N_23395,N_22536,N_22761);
or U23396 (N_23396,N_22967,N_22669);
nor U23397 (N_23397,N_22630,N_22606);
nor U23398 (N_23398,N_22806,N_22812);
and U23399 (N_23399,N_22648,N_22565);
xor U23400 (N_23400,N_22924,N_22994);
and U23401 (N_23401,N_22805,N_22646);
nand U23402 (N_23402,N_22868,N_22693);
nor U23403 (N_23403,N_22866,N_22691);
nand U23404 (N_23404,N_22962,N_22711);
or U23405 (N_23405,N_22692,N_22586);
xor U23406 (N_23406,N_22547,N_22948);
nor U23407 (N_23407,N_22541,N_22791);
xor U23408 (N_23408,N_22644,N_22526);
or U23409 (N_23409,N_22939,N_22601);
xor U23410 (N_23410,N_22941,N_22750);
nor U23411 (N_23411,N_22675,N_22836);
xnor U23412 (N_23412,N_22783,N_22882);
nor U23413 (N_23413,N_22702,N_22539);
and U23414 (N_23414,N_22675,N_22917);
nor U23415 (N_23415,N_22933,N_22805);
nand U23416 (N_23416,N_22987,N_22704);
or U23417 (N_23417,N_22925,N_22614);
and U23418 (N_23418,N_22972,N_22769);
and U23419 (N_23419,N_22746,N_22963);
nand U23420 (N_23420,N_22812,N_22537);
xnor U23421 (N_23421,N_22975,N_22969);
or U23422 (N_23422,N_22729,N_22694);
nand U23423 (N_23423,N_22669,N_22895);
xor U23424 (N_23424,N_22851,N_22576);
and U23425 (N_23425,N_22653,N_22740);
nor U23426 (N_23426,N_22575,N_22508);
or U23427 (N_23427,N_22639,N_22978);
nand U23428 (N_23428,N_22945,N_22928);
or U23429 (N_23429,N_22655,N_22900);
xnor U23430 (N_23430,N_22541,N_22581);
nor U23431 (N_23431,N_22749,N_22846);
and U23432 (N_23432,N_22885,N_22681);
nand U23433 (N_23433,N_22519,N_22697);
and U23434 (N_23434,N_22737,N_22931);
and U23435 (N_23435,N_22589,N_22749);
and U23436 (N_23436,N_22863,N_22864);
and U23437 (N_23437,N_22542,N_22559);
xor U23438 (N_23438,N_22916,N_22741);
and U23439 (N_23439,N_22688,N_22895);
nand U23440 (N_23440,N_22820,N_22652);
and U23441 (N_23441,N_22731,N_22887);
xor U23442 (N_23442,N_22516,N_22812);
xor U23443 (N_23443,N_22829,N_22526);
nand U23444 (N_23444,N_22883,N_22757);
and U23445 (N_23445,N_22940,N_22871);
or U23446 (N_23446,N_22993,N_22661);
nor U23447 (N_23447,N_22965,N_22880);
nand U23448 (N_23448,N_22787,N_22687);
and U23449 (N_23449,N_22646,N_22714);
or U23450 (N_23450,N_22920,N_22615);
nor U23451 (N_23451,N_22919,N_22549);
and U23452 (N_23452,N_22663,N_22833);
or U23453 (N_23453,N_22886,N_22782);
xnor U23454 (N_23454,N_22747,N_22991);
and U23455 (N_23455,N_22609,N_22540);
nand U23456 (N_23456,N_22827,N_22958);
xnor U23457 (N_23457,N_22777,N_22960);
xor U23458 (N_23458,N_22915,N_22814);
or U23459 (N_23459,N_22643,N_22995);
nor U23460 (N_23460,N_22947,N_22571);
nand U23461 (N_23461,N_22830,N_22557);
xnor U23462 (N_23462,N_22598,N_22768);
or U23463 (N_23463,N_22907,N_22776);
nor U23464 (N_23464,N_22864,N_22832);
xnor U23465 (N_23465,N_22666,N_22560);
nor U23466 (N_23466,N_22577,N_22538);
or U23467 (N_23467,N_22632,N_22819);
nor U23468 (N_23468,N_22695,N_22750);
and U23469 (N_23469,N_22724,N_22979);
nand U23470 (N_23470,N_22835,N_22809);
nand U23471 (N_23471,N_22842,N_22607);
xor U23472 (N_23472,N_22870,N_22519);
xor U23473 (N_23473,N_22945,N_22807);
nor U23474 (N_23474,N_22887,N_22685);
and U23475 (N_23475,N_22916,N_22526);
or U23476 (N_23476,N_22552,N_22635);
or U23477 (N_23477,N_22951,N_22647);
xnor U23478 (N_23478,N_22792,N_22543);
xor U23479 (N_23479,N_22817,N_22807);
and U23480 (N_23480,N_22874,N_22994);
and U23481 (N_23481,N_22863,N_22848);
nor U23482 (N_23482,N_22974,N_22697);
or U23483 (N_23483,N_22670,N_22629);
xnor U23484 (N_23484,N_22960,N_22921);
xor U23485 (N_23485,N_22994,N_22848);
xnor U23486 (N_23486,N_22736,N_22757);
nor U23487 (N_23487,N_22555,N_22604);
or U23488 (N_23488,N_22511,N_22743);
nand U23489 (N_23489,N_22742,N_22636);
and U23490 (N_23490,N_22788,N_22706);
nor U23491 (N_23491,N_22997,N_22849);
or U23492 (N_23492,N_22892,N_22672);
nor U23493 (N_23493,N_22910,N_22899);
xnor U23494 (N_23494,N_22848,N_22661);
and U23495 (N_23495,N_22591,N_22694);
and U23496 (N_23496,N_22803,N_22861);
or U23497 (N_23497,N_22641,N_22845);
and U23498 (N_23498,N_22715,N_22699);
nand U23499 (N_23499,N_22769,N_22926);
xor U23500 (N_23500,N_23043,N_23492);
nand U23501 (N_23501,N_23366,N_23219);
and U23502 (N_23502,N_23063,N_23186);
nand U23503 (N_23503,N_23049,N_23406);
or U23504 (N_23504,N_23298,N_23344);
xnor U23505 (N_23505,N_23073,N_23323);
nor U23506 (N_23506,N_23267,N_23170);
xor U23507 (N_23507,N_23211,N_23295);
xor U23508 (N_23508,N_23081,N_23355);
and U23509 (N_23509,N_23411,N_23475);
and U23510 (N_23510,N_23490,N_23131);
or U23511 (N_23511,N_23104,N_23258);
xor U23512 (N_23512,N_23433,N_23383);
nand U23513 (N_23513,N_23239,N_23398);
nand U23514 (N_23514,N_23487,N_23044);
nor U23515 (N_23515,N_23498,N_23294);
xnor U23516 (N_23516,N_23201,N_23385);
xor U23517 (N_23517,N_23160,N_23233);
nand U23518 (N_23518,N_23285,N_23351);
xor U23519 (N_23519,N_23362,N_23273);
xnor U23520 (N_23520,N_23336,N_23332);
nor U23521 (N_23521,N_23140,N_23126);
and U23522 (N_23522,N_23051,N_23471);
nand U23523 (N_23523,N_23256,N_23269);
nor U23524 (N_23524,N_23265,N_23427);
or U23525 (N_23525,N_23138,N_23486);
nor U23526 (N_23526,N_23047,N_23390);
nor U23527 (N_23527,N_23112,N_23062);
nand U23528 (N_23528,N_23464,N_23177);
or U23529 (N_23529,N_23036,N_23455);
and U23530 (N_23530,N_23147,N_23228);
and U23531 (N_23531,N_23139,N_23234);
or U23532 (N_23532,N_23397,N_23013);
xnor U23533 (N_23533,N_23283,N_23071);
xnor U23534 (N_23534,N_23320,N_23064);
xnor U23535 (N_23535,N_23156,N_23286);
nor U23536 (N_23536,N_23200,N_23114);
and U23537 (N_23537,N_23472,N_23018);
and U23538 (N_23538,N_23252,N_23457);
or U23539 (N_23539,N_23148,N_23082);
nand U23540 (N_23540,N_23491,N_23105);
or U23541 (N_23541,N_23137,N_23149);
or U23542 (N_23542,N_23038,N_23000);
and U23543 (N_23543,N_23128,N_23442);
and U23544 (N_23544,N_23226,N_23374);
nand U23545 (N_23545,N_23015,N_23447);
or U23546 (N_23546,N_23399,N_23422);
nand U23547 (N_23547,N_23244,N_23032);
nor U23548 (N_23548,N_23317,N_23180);
nand U23549 (N_23549,N_23263,N_23040);
or U23550 (N_23550,N_23431,N_23257);
xnor U23551 (N_23551,N_23477,N_23430);
nand U23552 (N_23552,N_23438,N_23277);
nand U23553 (N_23553,N_23495,N_23246);
nand U23554 (N_23554,N_23094,N_23021);
nand U23555 (N_23555,N_23004,N_23150);
nor U23556 (N_23556,N_23005,N_23087);
or U23557 (N_23557,N_23307,N_23299);
xnor U23558 (N_23558,N_23347,N_23067);
or U23559 (N_23559,N_23291,N_23225);
nand U23560 (N_23560,N_23353,N_23189);
xnor U23561 (N_23561,N_23202,N_23454);
nand U23562 (N_23562,N_23023,N_23297);
nor U23563 (N_23563,N_23407,N_23006);
nor U23564 (N_23564,N_23065,N_23035);
nand U23565 (N_23565,N_23496,N_23394);
and U23566 (N_23566,N_23145,N_23412);
and U23567 (N_23567,N_23152,N_23016);
and U23568 (N_23568,N_23345,N_23250);
and U23569 (N_23569,N_23441,N_23480);
nor U23570 (N_23570,N_23079,N_23003);
or U23571 (N_23571,N_23260,N_23264);
or U23572 (N_23572,N_23382,N_23088);
and U23573 (N_23573,N_23135,N_23426);
nor U23574 (N_23574,N_23077,N_23236);
or U23575 (N_23575,N_23174,N_23384);
xnor U23576 (N_23576,N_23127,N_23381);
nor U23577 (N_23577,N_23130,N_23227);
and U23578 (N_23578,N_23279,N_23237);
nor U23579 (N_23579,N_23074,N_23388);
xor U23580 (N_23580,N_23474,N_23059);
nand U23581 (N_23581,N_23042,N_23334);
and U23582 (N_23582,N_23162,N_23371);
nand U23583 (N_23583,N_23330,N_23499);
nand U23584 (N_23584,N_23254,N_23253);
or U23585 (N_23585,N_23377,N_23415);
nor U23586 (N_23586,N_23497,N_23343);
nand U23587 (N_23587,N_23274,N_23363);
or U23588 (N_23588,N_23421,N_23197);
or U23589 (N_23589,N_23403,N_23448);
nand U23590 (N_23590,N_23117,N_23419);
nor U23591 (N_23591,N_23066,N_23194);
nor U23592 (N_23592,N_23292,N_23316);
nor U23593 (N_23593,N_23359,N_23303);
nor U23594 (N_23594,N_23091,N_23181);
nand U23595 (N_23595,N_23466,N_23488);
or U23596 (N_23596,N_23187,N_23108);
nor U23597 (N_23597,N_23360,N_23123);
or U23598 (N_23598,N_23103,N_23208);
or U23599 (N_23599,N_23439,N_23107);
and U23600 (N_23600,N_23163,N_23270);
or U23601 (N_23601,N_23259,N_23461);
and U23602 (N_23602,N_23012,N_23031);
nor U23603 (N_23603,N_23075,N_23481);
nor U23604 (N_23604,N_23207,N_23408);
xnor U23605 (N_23605,N_23161,N_23098);
or U23606 (N_23606,N_23241,N_23240);
nor U23607 (N_23607,N_23052,N_23235);
or U23608 (N_23608,N_23251,N_23095);
xnor U23609 (N_23609,N_23232,N_23453);
or U23610 (N_23610,N_23078,N_23056);
or U23611 (N_23611,N_23282,N_23296);
and U23612 (N_23612,N_23440,N_23166);
xnor U23613 (N_23613,N_23178,N_23167);
xor U23614 (N_23614,N_23218,N_23121);
xor U23615 (N_23615,N_23272,N_23190);
xnor U23616 (N_23616,N_23357,N_23155);
xnor U23617 (N_23617,N_23185,N_23468);
or U23618 (N_23618,N_23300,N_23312);
nand U23619 (N_23619,N_23308,N_23302);
nor U23620 (N_23620,N_23379,N_23093);
nor U23621 (N_23621,N_23048,N_23395);
and U23622 (N_23622,N_23168,N_23165);
nand U23623 (N_23623,N_23324,N_23281);
or U23624 (N_23624,N_23055,N_23276);
nand U23625 (N_23625,N_23169,N_23340);
xnor U23626 (N_23626,N_23428,N_23255);
or U23627 (N_23627,N_23389,N_23084);
nor U23628 (N_23628,N_23060,N_23376);
nand U23629 (N_23629,N_23310,N_23204);
nand U23630 (N_23630,N_23171,N_23230);
or U23631 (N_23631,N_23070,N_23460);
nand U23632 (N_23632,N_23293,N_23311);
or U23633 (N_23633,N_23322,N_23444);
xor U23634 (N_23634,N_23482,N_23159);
nand U23635 (N_23635,N_23205,N_23304);
or U23636 (N_23636,N_23008,N_23248);
and U23637 (N_23637,N_23026,N_23425);
xnor U23638 (N_23638,N_23215,N_23364);
xnor U23639 (N_23639,N_23418,N_23305);
xnor U23640 (N_23640,N_23212,N_23321);
and U23641 (N_23641,N_23420,N_23154);
xnor U23642 (N_23642,N_23125,N_23493);
and U23643 (N_23643,N_23375,N_23280);
and U23644 (N_23644,N_23306,N_23456);
or U23645 (N_23645,N_23446,N_23086);
xnor U23646 (N_23646,N_23367,N_23229);
nand U23647 (N_23647,N_23266,N_23132);
nor U23648 (N_23648,N_23452,N_23409);
nor U23649 (N_23649,N_23096,N_23120);
nand U23650 (N_23650,N_23097,N_23039);
and U23651 (N_23651,N_23157,N_23053);
nand U23652 (N_23652,N_23405,N_23476);
or U23653 (N_23653,N_23172,N_23247);
nand U23654 (N_23654,N_23262,N_23494);
or U23655 (N_23655,N_23069,N_23058);
xnor U23656 (N_23656,N_23467,N_23313);
and U23657 (N_23657,N_23118,N_23243);
or U23658 (N_23658,N_23356,N_23002);
or U23659 (N_23659,N_23393,N_23102);
nand U23660 (N_23660,N_23319,N_23144);
nand U23661 (N_23661,N_23315,N_23220);
xnor U23662 (N_23662,N_23068,N_23136);
or U23663 (N_23663,N_23231,N_23119);
or U23664 (N_23664,N_23027,N_23268);
or U23665 (N_23665,N_23416,N_23338);
xnor U23666 (N_23666,N_23432,N_23436);
and U23667 (N_23667,N_23326,N_23478);
nor U23668 (N_23668,N_23184,N_23349);
and U23669 (N_23669,N_23115,N_23361);
nor U23670 (N_23670,N_23214,N_23443);
nor U23671 (N_23671,N_23209,N_23141);
nor U23672 (N_23672,N_23116,N_23124);
nand U23673 (N_23673,N_23033,N_23470);
nor U23674 (N_23674,N_23007,N_23458);
and U23675 (N_23675,N_23301,N_23224);
and U23676 (N_23676,N_23057,N_23372);
nor U23677 (N_23677,N_23271,N_23216);
xnor U23678 (N_23678,N_23245,N_23451);
and U23679 (N_23679,N_23459,N_23391);
or U23680 (N_23680,N_23024,N_23348);
nand U23681 (N_23681,N_23401,N_23182);
nor U23682 (N_23682,N_23223,N_23191);
or U23683 (N_23683,N_23196,N_23373);
and U23684 (N_23684,N_23198,N_23176);
nor U23685 (N_23685,N_23080,N_23142);
nand U23686 (N_23686,N_23188,N_23369);
nand U23687 (N_23687,N_23146,N_23333);
nand U23688 (N_23688,N_23350,N_23378);
or U23689 (N_23689,N_23370,N_23358);
and U23690 (N_23690,N_23179,N_23473);
xnor U23691 (N_23691,N_23484,N_23337);
nor U23692 (N_23692,N_23396,N_23109);
nor U23693 (N_23693,N_23164,N_23354);
xor U23694 (N_23694,N_23489,N_23175);
and U23695 (N_23695,N_23089,N_23392);
xor U23696 (N_23696,N_23203,N_23099);
nand U23697 (N_23697,N_23404,N_23045);
or U23698 (N_23698,N_23028,N_23054);
nor U23699 (N_23699,N_23380,N_23110);
nand U23700 (N_23700,N_23287,N_23485);
nand U23701 (N_23701,N_23022,N_23106);
nand U23702 (N_23702,N_23242,N_23206);
xor U23703 (N_23703,N_23331,N_23037);
nand U23704 (N_23704,N_23402,N_23129);
and U23705 (N_23705,N_23314,N_23193);
xor U23706 (N_23706,N_23173,N_23429);
nor U23707 (N_23707,N_23365,N_23221);
nor U23708 (N_23708,N_23386,N_23025);
xnor U23709 (N_23709,N_23009,N_23434);
nand U23710 (N_23710,N_23424,N_23083);
nand U23711 (N_23711,N_23011,N_23183);
and U23712 (N_23712,N_23111,N_23050);
nand U23713 (N_23713,N_23041,N_23100);
or U23714 (N_23714,N_23090,N_23462);
nor U23715 (N_23715,N_23469,N_23450);
xor U23716 (N_23716,N_23261,N_23213);
nor U23717 (N_23717,N_23010,N_23133);
xor U23718 (N_23718,N_23387,N_23342);
nor U23719 (N_23719,N_23122,N_23143);
and U23720 (N_23720,N_23329,N_23072);
xnor U23721 (N_23721,N_23076,N_23238);
and U23722 (N_23722,N_23275,N_23046);
nor U23723 (N_23723,N_23019,N_23437);
nor U23724 (N_23724,N_23034,N_23217);
nand U23725 (N_23725,N_23309,N_23288);
nor U23726 (N_23726,N_23085,N_23423);
and U23727 (N_23727,N_23327,N_23290);
nor U23728 (N_23728,N_23029,N_23134);
xor U23729 (N_23729,N_23092,N_23335);
nand U23730 (N_23730,N_23030,N_23284);
and U23731 (N_23731,N_23410,N_23328);
nor U23732 (N_23732,N_23479,N_23014);
nand U23733 (N_23733,N_23222,N_23289);
and U23734 (N_23734,N_23325,N_23195);
nor U23735 (N_23735,N_23061,N_23368);
or U23736 (N_23736,N_23417,N_23192);
nor U23737 (N_23737,N_23017,N_23101);
or U23738 (N_23738,N_23400,N_23001);
or U23739 (N_23739,N_23278,N_23483);
and U23740 (N_23740,N_23414,N_23249);
and U23741 (N_23741,N_23020,N_23449);
nor U23742 (N_23742,N_23465,N_23199);
nor U23743 (N_23743,N_23341,N_23352);
nor U23744 (N_23744,N_23463,N_23210);
or U23745 (N_23745,N_23158,N_23435);
or U23746 (N_23746,N_23445,N_23113);
nand U23747 (N_23747,N_23151,N_23153);
nor U23748 (N_23748,N_23413,N_23339);
xnor U23749 (N_23749,N_23346,N_23318);
nor U23750 (N_23750,N_23476,N_23417);
nor U23751 (N_23751,N_23294,N_23260);
nand U23752 (N_23752,N_23225,N_23303);
or U23753 (N_23753,N_23059,N_23463);
or U23754 (N_23754,N_23385,N_23124);
xnor U23755 (N_23755,N_23183,N_23385);
nor U23756 (N_23756,N_23195,N_23037);
nand U23757 (N_23757,N_23339,N_23427);
xor U23758 (N_23758,N_23170,N_23009);
xor U23759 (N_23759,N_23467,N_23108);
xnor U23760 (N_23760,N_23454,N_23288);
or U23761 (N_23761,N_23050,N_23327);
xor U23762 (N_23762,N_23345,N_23362);
or U23763 (N_23763,N_23093,N_23459);
nand U23764 (N_23764,N_23034,N_23055);
nand U23765 (N_23765,N_23491,N_23442);
nor U23766 (N_23766,N_23001,N_23179);
or U23767 (N_23767,N_23408,N_23449);
or U23768 (N_23768,N_23474,N_23005);
nor U23769 (N_23769,N_23474,N_23068);
xor U23770 (N_23770,N_23365,N_23170);
nor U23771 (N_23771,N_23135,N_23347);
nand U23772 (N_23772,N_23052,N_23225);
xnor U23773 (N_23773,N_23363,N_23452);
nand U23774 (N_23774,N_23008,N_23061);
xnor U23775 (N_23775,N_23210,N_23433);
or U23776 (N_23776,N_23217,N_23276);
nand U23777 (N_23777,N_23365,N_23166);
or U23778 (N_23778,N_23364,N_23128);
nor U23779 (N_23779,N_23301,N_23252);
xor U23780 (N_23780,N_23396,N_23235);
nand U23781 (N_23781,N_23376,N_23175);
and U23782 (N_23782,N_23286,N_23249);
or U23783 (N_23783,N_23451,N_23181);
xnor U23784 (N_23784,N_23218,N_23360);
nand U23785 (N_23785,N_23405,N_23244);
nand U23786 (N_23786,N_23182,N_23076);
or U23787 (N_23787,N_23262,N_23114);
xnor U23788 (N_23788,N_23478,N_23366);
and U23789 (N_23789,N_23349,N_23015);
and U23790 (N_23790,N_23195,N_23407);
and U23791 (N_23791,N_23062,N_23372);
nor U23792 (N_23792,N_23259,N_23239);
or U23793 (N_23793,N_23247,N_23362);
nand U23794 (N_23794,N_23201,N_23329);
or U23795 (N_23795,N_23432,N_23183);
xnor U23796 (N_23796,N_23393,N_23035);
nand U23797 (N_23797,N_23142,N_23343);
nor U23798 (N_23798,N_23387,N_23066);
nand U23799 (N_23799,N_23293,N_23053);
nor U23800 (N_23800,N_23489,N_23415);
nand U23801 (N_23801,N_23007,N_23132);
xnor U23802 (N_23802,N_23394,N_23014);
nor U23803 (N_23803,N_23117,N_23368);
nor U23804 (N_23804,N_23229,N_23407);
xor U23805 (N_23805,N_23403,N_23336);
xnor U23806 (N_23806,N_23099,N_23430);
and U23807 (N_23807,N_23187,N_23498);
and U23808 (N_23808,N_23168,N_23188);
xnor U23809 (N_23809,N_23086,N_23272);
nand U23810 (N_23810,N_23437,N_23070);
nand U23811 (N_23811,N_23324,N_23466);
or U23812 (N_23812,N_23433,N_23419);
xnor U23813 (N_23813,N_23367,N_23240);
xnor U23814 (N_23814,N_23281,N_23204);
nand U23815 (N_23815,N_23238,N_23320);
nand U23816 (N_23816,N_23375,N_23008);
xor U23817 (N_23817,N_23498,N_23254);
nand U23818 (N_23818,N_23341,N_23105);
xnor U23819 (N_23819,N_23251,N_23340);
nor U23820 (N_23820,N_23384,N_23064);
nand U23821 (N_23821,N_23452,N_23013);
nor U23822 (N_23822,N_23042,N_23486);
nand U23823 (N_23823,N_23021,N_23174);
and U23824 (N_23824,N_23195,N_23200);
and U23825 (N_23825,N_23228,N_23046);
nor U23826 (N_23826,N_23056,N_23007);
nand U23827 (N_23827,N_23098,N_23483);
xnor U23828 (N_23828,N_23071,N_23228);
and U23829 (N_23829,N_23183,N_23076);
xnor U23830 (N_23830,N_23052,N_23430);
nor U23831 (N_23831,N_23018,N_23181);
xor U23832 (N_23832,N_23223,N_23389);
or U23833 (N_23833,N_23440,N_23487);
nor U23834 (N_23834,N_23066,N_23248);
nand U23835 (N_23835,N_23305,N_23034);
or U23836 (N_23836,N_23077,N_23303);
or U23837 (N_23837,N_23190,N_23105);
or U23838 (N_23838,N_23154,N_23290);
nand U23839 (N_23839,N_23322,N_23181);
xor U23840 (N_23840,N_23366,N_23197);
xor U23841 (N_23841,N_23459,N_23299);
nand U23842 (N_23842,N_23304,N_23029);
or U23843 (N_23843,N_23372,N_23491);
and U23844 (N_23844,N_23152,N_23025);
xnor U23845 (N_23845,N_23208,N_23271);
or U23846 (N_23846,N_23419,N_23174);
and U23847 (N_23847,N_23022,N_23025);
or U23848 (N_23848,N_23389,N_23025);
and U23849 (N_23849,N_23135,N_23351);
and U23850 (N_23850,N_23488,N_23383);
and U23851 (N_23851,N_23209,N_23391);
nand U23852 (N_23852,N_23306,N_23491);
or U23853 (N_23853,N_23266,N_23392);
nor U23854 (N_23854,N_23495,N_23140);
or U23855 (N_23855,N_23140,N_23153);
nand U23856 (N_23856,N_23248,N_23106);
or U23857 (N_23857,N_23053,N_23338);
or U23858 (N_23858,N_23079,N_23416);
nor U23859 (N_23859,N_23125,N_23126);
and U23860 (N_23860,N_23305,N_23434);
nor U23861 (N_23861,N_23412,N_23257);
nand U23862 (N_23862,N_23124,N_23355);
nand U23863 (N_23863,N_23427,N_23037);
and U23864 (N_23864,N_23154,N_23359);
xor U23865 (N_23865,N_23080,N_23207);
nand U23866 (N_23866,N_23046,N_23086);
xor U23867 (N_23867,N_23285,N_23074);
nand U23868 (N_23868,N_23210,N_23301);
nand U23869 (N_23869,N_23243,N_23215);
nand U23870 (N_23870,N_23452,N_23360);
or U23871 (N_23871,N_23028,N_23250);
or U23872 (N_23872,N_23186,N_23034);
nor U23873 (N_23873,N_23266,N_23181);
or U23874 (N_23874,N_23099,N_23003);
nand U23875 (N_23875,N_23276,N_23250);
xnor U23876 (N_23876,N_23150,N_23212);
nand U23877 (N_23877,N_23149,N_23479);
nand U23878 (N_23878,N_23173,N_23425);
and U23879 (N_23879,N_23379,N_23411);
nor U23880 (N_23880,N_23115,N_23289);
nor U23881 (N_23881,N_23483,N_23294);
xor U23882 (N_23882,N_23062,N_23383);
and U23883 (N_23883,N_23447,N_23401);
or U23884 (N_23884,N_23426,N_23377);
and U23885 (N_23885,N_23357,N_23041);
nand U23886 (N_23886,N_23004,N_23466);
xor U23887 (N_23887,N_23279,N_23040);
xnor U23888 (N_23888,N_23312,N_23047);
nand U23889 (N_23889,N_23339,N_23139);
or U23890 (N_23890,N_23060,N_23210);
xnor U23891 (N_23891,N_23386,N_23093);
or U23892 (N_23892,N_23270,N_23203);
or U23893 (N_23893,N_23401,N_23050);
or U23894 (N_23894,N_23251,N_23252);
or U23895 (N_23895,N_23096,N_23422);
nor U23896 (N_23896,N_23412,N_23317);
nor U23897 (N_23897,N_23147,N_23178);
nor U23898 (N_23898,N_23420,N_23045);
or U23899 (N_23899,N_23226,N_23196);
or U23900 (N_23900,N_23496,N_23157);
or U23901 (N_23901,N_23426,N_23218);
xor U23902 (N_23902,N_23105,N_23122);
or U23903 (N_23903,N_23059,N_23170);
and U23904 (N_23904,N_23169,N_23491);
xor U23905 (N_23905,N_23112,N_23299);
nand U23906 (N_23906,N_23343,N_23177);
nand U23907 (N_23907,N_23341,N_23316);
or U23908 (N_23908,N_23277,N_23261);
nand U23909 (N_23909,N_23412,N_23378);
nand U23910 (N_23910,N_23364,N_23376);
nand U23911 (N_23911,N_23233,N_23188);
nand U23912 (N_23912,N_23010,N_23344);
or U23913 (N_23913,N_23052,N_23349);
and U23914 (N_23914,N_23211,N_23439);
nand U23915 (N_23915,N_23063,N_23108);
nor U23916 (N_23916,N_23206,N_23488);
nand U23917 (N_23917,N_23397,N_23284);
or U23918 (N_23918,N_23178,N_23492);
nor U23919 (N_23919,N_23337,N_23091);
nor U23920 (N_23920,N_23254,N_23125);
nand U23921 (N_23921,N_23309,N_23270);
xnor U23922 (N_23922,N_23495,N_23384);
nand U23923 (N_23923,N_23293,N_23192);
xnor U23924 (N_23924,N_23073,N_23197);
and U23925 (N_23925,N_23337,N_23442);
or U23926 (N_23926,N_23084,N_23234);
xnor U23927 (N_23927,N_23045,N_23490);
xnor U23928 (N_23928,N_23494,N_23396);
nand U23929 (N_23929,N_23095,N_23345);
nand U23930 (N_23930,N_23444,N_23477);
and U23931 (N_23931,N_23374,N_23428);
nand U23932 (N_23932,N_23362,N_23354);
nor U23933 (N_23933,N_23250,N_23003);
nor U23934 (N_23934,N_23417,N_23277);
nand U23935 (N_23935,N_23417,N_23470);
nor U23936 (N_23936,N_23188,N_23485);
and U23937 (N_23937,N_23198,N_23002);
nor U23938 (N_23938,N_23374,N_23335);
xor U23939 (N_23939,N_23323,N_23197);
and U23940 (N_23940,N_23449,N_23133);
and U23941 (N_23941,N_23283,N_23370);
or U23942 (N_23942,N_23221,N_23320);
or U23943 (N_23943,N_23098,N_23240);
nand U23944 (N_23944,N_23183,N_23134);
xor U23945 (N_23945,N_23389,N_23411);
and U23946 (N_23946,N_23372,N_23100);
or U23947 (N_23947,N_23482,N_23037);
nor U23948 (N_23948,N_23308,N_23105);
nand U23949 (N_23949,N_23348,N_23387);
xor U23950 (N_23950,N_23200,N_23113);
or U23951 (N_23951,N_23329,N_23256);
nor U23952 (N_23952,N_23013,N_23197);
xor U23953 (N_23953,N_23119,N_23162);
and U23954 (N_23954,N_23066,N_23329);
xnor U23955 (N_23955,N_23160,N_23147);
nor U23956 (N_23956,N_23477,N_23034);
or U23957 (N_23957,N_23216,N_23230);
or U23958 (N_23958,N_23353,N_23192);
xor U23959 (N_23959,N_23069,N_23479);
xor U23960 (N_23960,N_23309,N_23023);
xor U23961 (N_23961,N_23059,N_23149);
nand U23962 (N_23962,N_23281,N_23025);
xnor U23963 (N_23963,N_23106,N_23290);
nand U23964 (N_23964,N_23144,N_23389);
or U23965 (N_23965,N_23052,N_23283);
nor U23966 (N_23966,N_23061,N_23206);
and U23967 (N_23967,N_23307,N_23127);
and U23968 (N_23968,N_23071,N_23067);
and U23969 (N_23969,N_23056,N_23102);
nand U23970 (N_23970,N_23146,N_23271);
or U23971 (N_23971,N_23071,N_23176);
nand U23972 (N_23972,N_23032,N_23461);
nand U23973 (N_23973,N_23106,N_23094);
nand U23974 (N_23974,N_23303,N_23498);
and U23975 (N_23975,N_23328,N_23284);
xnor U23976 (N_23976,N_23186,N_23199);
and U23977 (N_23977,N_23223,N_23467);
and U23978 (N_23978,N_23052,N_23030);
xor U23979 (N_23979,N_23448,N_23268);
xnor U23980 (N_23980,N_23478,N_23199);
xnor U23981 (N_23981,N_23050,N_23187);
or U23982 (N_23982,N_23182,N_23146);
or U23983 (N_23983,N_23494,N_23110);
xnor U23984 (N_23984,N_23226,N_23360);
xnor U23985 (N_23985,N_23432,N_23351);
or U23986 (N_23986,N_23272,N_23327);
xnor U23987 (N_23987,N_23447,N_23058);
or U23988 (N_23988,N_23323,N_23211);
nor U23989 (N_23989,N_23098,N_23388);
nand U23990 (N_23990,N_23441,N_23016);
and U23991 (N_23991,N_23223,N_23224);
nand U23992 (N_23992,N_23233,N_23016);
xor U23993 (N_23993,N_23427,N_23060);
xnor U23994 (N_23994,N_23426,N_23187);
or U23995 (N_23995,N_23019,N_23414);
xor U23996 (N_23996,N_23044,N_23232);
or U23997 (N_23997,N_23092,N_23184);
or U23998 (N_23998,N_23167,N_23084);
nor U23999 (N_23999,N_23207,N_23099);
nand U24000 (N_24000,N_23575,N_23852);
and U24001 (N_24001,N_23760,N_23579);
nand U24002 (N_24002,N_23952,N_23652);
nor U24003 (N_24003,N_23746,N_23784);
and U24004 (N_24004,N_23881,N_23797);
nor U24005 (N_24005,N_23820,N_23933);
nand U24006 (N_24006,N_23866,N_23566);
nor U24007 (N_24007,N_23741,N_23774);
and U24008 (N_24008,N_23752,N_23620);
xor U24009 (N_24009,N_23546,N_23674);
or U24010 (N_24010,N_23902,N_23993);
and U24011 (N_24011,N_23920,N_23813);
xor U24012 (N_24012,N_23505,N_23925);
xnor U24013 (N_24013,N_23529,N_23709);
nand U24014 (N_24014,N_23814,N_23560);
nand U24015 (N_24015,N_23851,N_23842);
and U24016 (N_24016,N_23795,N_23959);
or U24017 (N_24017,N_23834,N_23829);
xnor U24018 (N_24018,N_23670,N_23544);
xor U24019 (N_24019,N_23901,N_23998);
or U24020 (N_24020,N_23808,N_23922);
and U24021 (N_24021,N_23754,N_23504);
or U24022 (N_24022,N_23703,N_23898);
nor U24023 (N_24023,N_23833,N_23605);
nor U24024 (N_24024,N_23695,N_23590);
nor U24025 (N_24025,N_23728,N_23608);
and U24026 (N_24026,N_23916,N_23651);
nor U24027 (N_24027,N_23937,N_23525);
xor U24028 (N_24028,N_23982,N_23981);
or U24029 (N_24029,N_23569,N_23715);
xor U24030 (N_24030,N_23841,N_23618);
nand U24031 (N_24031,N_23750,N_23923);
xor U24032 (N_24032,N_23989,N_23592);
and U24033 (N_24033,N_23509,N_23938);
and U24034 (N_24034,N_23997,N_23751);
nand U24035 (N_24035,N_23532,N_23664);
xnor U24036 (N_24036,N_23966,N_23817);
nand U24037 (N_24037,N_23671,N_23656);
and U24038 (N_24038,N_23800,N_23921);
xnor U24039 (N_24039,N_23619,N_23684);
xor U24040 (N_24040,N_23976,N_23734);
xnor U24041 (N_24041,N_23697,N_23819);
nor U24042 (N_24042,N_23617,N_23791);
or U24043 (N_24043,N_23642,N_23588);
nand U24044 (N_24044,N_23578,N_23700);
nor U24045 (N_24045,N_23957,N_23869);
nand U24046 (N_24046,N_23726,N_23847);
nand U24047 (N_24047,N_23984,N_23731);
xnor U24048 (N_24048,N_23634,N_23767);
nor U24049 (N_24049,N_23538,N_23553);
nand U24050 (N_24050,N_23971,N_23837);
xnor U24051 (N_24051,N_23850,N_23517);
and U24052 (N_24052,N_23650,N_23948);
nor U24053 (N_24053,N_23706,N_23843);
or U24054 (N_24054,N_23615,N_23811);
nor U24055 (N_24055,N_23968,N_23704);
or U24056 (N_24056,N_23707,N_23864);
or U24057 (N_24057,N_23939,N_23806);
xnor U24058 (N_24058,N_23687,N_23961);
xnor U24059 (N_24059,N_23717,N_23798);
and U24060 (N_24060,N_23994,N_23978);
nand U24061 (N_24061,N_23649,N_23551);
xor U24062 (N_24062,N_23780,N_23533);
or U24063 (N_24063,N_23882,N_23637);
xnor U24064 (N_24064,N_23844,N_23522);
xnor U24065 (N_24065,N_23802,N_23679);
nand U24066 (N_24066,N_23963,N_23911);
or U24067 (N_24067,N_23807,N_23770);
or U24068 (N_24068,N_23555,N_23536);
xnor U24069 (N_24069,N_23613,N_23904);
and U24070 (N_24070,N_23614,N_23556);
or U24071 (N_24071,N_23849,N_23738);
nand U24072 (N_24072,N_23768,N_23875);
nand U24073 (N_24073,N_23860,N_23794);
and U24074 (N_24074,N_23520,N_23861);
or U24075 (N_24075,N_23924,N_23756);
or U24076 (N_24076,N_23992,N_23762);
nand U24077 (N_24077,N_23960,N_23534);
xor U24078 (N_24078,N_23668,N_23627);
nor U24079 (N_24079,N_23776,N_23962);
or U24080 (N_24080,N_23694,N_23683);
xor U24081 (N_24081,N_23822,N_23660);
nor U24082 (N_24082,N_23600,N_23836);
nor U24083 (N_24083,N_23724,N_23507);
or U24084 (N_24084,N_23908,N_23720);
xnor U24085 (N_24085,N_23931,N_23698);
xor U24086 (N_24086,N_23732,N_23586);
or U24087 (N_24087,N_23779,N_23910);
nor U24088 (N_24088,N_23990,N_23688);
nor U24089 (N_24089,N_23714,N_23644);
or U24090 (N_24090,N_23603,N_23543);
and U24091 (N_24091,N_23677,N_23718);
nand U24092 (N_24092,N_23624,N_23975);
nor U24093 (N_24093,N_23789,N_23635);
nand U24094 (N_24094,N_23643,N_23540);
or U24095 (N_24095,N_23895,N_23596);
nor U24096 (N_24096,N_23545,N_23893);
nand U24097 (N_24097,N_23782,N_23748);
nor U24098 (N_24098,N_23628,N_23725);
or U24099 (N_24099,N_23854,N_23705);
and U24100 (N_24100,N_23744,N_23577);
xnor U24101 (N_24101,N_23599,N_23828);
xnor U24102 (N_24102,N_23803,N_23737);
nand U24103 (N_24103,N_23763,N_23810);
nor U24104 (N_24104,N_23740,N_23874);
xnor U24105 (N_24105,N_23610,N_23884);
nor U24106 (N_24106,N_23712,N_23796);
xor U24107 (N_24107,N_23988,N_23940);
xnor U24108 (N_24108,N_23974,N_23799);
and U24109 (N_24109,N_23502,N_23879);
nor U24110 (N_24110,N_23769,N_23735);
and U24111 (N_24111,N_23859,N_23891);
or U24112 (N_24112,N_23580,N_23573);
nand U24113 (N_24113,N_23870,N_23805);
and U24114 (N_24114,N_23629,N_23572);
nor U24115 (N_24115,N_23640,N_23742);
or U24116 (N_24116,N_23838,N_23500);
xnor U24117 (N_24117,N_23766,N_23680);
xnor U24118 (N_24118,N_23793,N_23858);
xor U24119 (N_24119,N_23669,N_23815);
nand U24120 (N_24120,N_23863,N_23835);
nand U24121 (N_24121,N_23778,N_23995);
or U24122 (N_24122,N_23818,N_23542);
or U24123 (N_24123,N_23749,N_23787);
nand U24124 (N_24124,N_23845,N_23999);
nor U24125 (N_24125,N_23661,N_23773);
nand U24126 (N_24126,N_23826,N_23755);
and U24127 (N_24127,N_23730,N_23515);
nand U24128 (N_24128,N_23945,N_23658);
nand U24129 (N_24129,N_23979,N_23591);
xor U24130 (N_24130,N_23987,N_23672);
nor U24131 (N_24131,N_23693,N_23840);
nor U24132 (N_24132,N_23927,N_23567);
or U24133 (N_24133,N_23785,N_23561);
xor U24134 (N_24134,N_23777,N_23513);
and U24135 (N_24135,N_23903,N_23936);
or U24136 (N_24136,N_23899,N_23606);
nor U24137 (N_24137,N_23878,N_23953);
and U24138 (N_24138,N_23956,N_23871);
or U24139 (N_24139,N_23523,N_23722);
and U24140 (N_24140,N_23954,N_23886);
xnor U24141 (N_24141,N_23535,N_23900);
xor U24142 (N_24142,N_23934,N_23885);
xor U24143 (N_24143,N_23865,N_23689);
or U24144 (N_24144,N_23930,N_23675);
or U24145 (N_24145,N_23648,N_23665);
and U24146 (N_24146,N_23510,N_23530);
nand U24147 (N_24147,N_23832,N_23639);
xor U24148 (N_24148,N_23616,N_23761);
nor U24149 (N_24149,N_23623,N_23926);
or U24150 (N_24150,N_23846,N_23554);
nand U24151 (N_24151,N_23857,N_23589);
nand U24152 (N_24152,N_23559,N_23662);
xor U24153 (N_24153,N_23611,N_23654);
and U24154 (N_24154,N_23950,N_23631);
and U24155 (N_24155,N_23757,N_23663);
or U24156 (N_24156,N_23699,N_23565);
xor U24157 (N_24157,N_23682,N_23892);
xnor U24158 (N_24158,N_23594,N_23514);
or U24159 (N_24159,N_23621,N_23919);
and U24160 (N_24160,N_23636,N_23583);
xnor U24161 (N_24161,N_23969,N_23653);
nand U24162 (N_24162,N_23716,N_23702);
nor U24163 (N_24163,N_23681,N_23537);
nand U24164 (N_24164,N_23853,N_23991);
nor U24165 (N_24165,N_23856,N_23501);
nor U24166 (N_24166,N_23827,N_23512);
or U24167 (N_24167,N_23967,N_23873);
nor U24168 (N_24168,N_23753,N_23701);
and U24169 (N_24169,N_23980,N_23977);
or U24170 (N_24170,N_23915,N_23585);
xor U24171 (N_24171,N_23888,N_23563);
and U24172 (N_24172,N_23907,N_23625);
nand U24173 (N_24173,N_23964,N_23788);
nor U24174 (N_24174,N_23801,N_23867);
nand U24175 (N_24175,N_23876,N_23595);
nor U24176 (N_24176,N_23632,N_23887);
and U24177 (N_24177,N_23521,N_23771);
or U24178 (N_24178,N_23508,N_23912);
xnor U24179 (N_24179,N_23986,N_23719);
and U24180 (N_24180,N_23790,N_23526);
nand U24181 (N_24181,N_23511,N_23727);
or U24182 (N_24182,N_23983,N_23909);
or U24183 (N_24183,N_23552,N_23574);
and U24184 (N_24184,N_23913,N_23929);
nor U24185 (N_24185,N_23759,N_23758);
and U24186 (N_24186,N_23710,N_23676);
nand U24187 (N_24187,N_23576,N_23612);
nor U24188 (N_24188,N_23816,N_23985);
xnor U24189 (N_24189,N_23872,N_23582);
nor U24190 (N_24190,N_23692,N_23868);
nand U24191 (N_24191,N_23647,N_23633);
xor U24192 (N_24192,N_23764,N_23713);
xnor U24193 (N_24193,N_23862,N_23729);
nor U24194 (N_24194,N_23733,N_23678);
nor U24195 (N_24195,N_23972,N_23955);
and U24196 (N_24196,N_23944,N_23570);
or U24197 (N_24197,N_23889,N_23519);
nand U24198 (N_24198,N_23932,N_23549);
or U24199 (N_24199,N_23593,N_23890);
or U24200 (N_24200,N_23584,N_23550);
nor U24201 (N_24201,N_23942,N_23638);
or U24202 (N_24202,N_23691,N_23839);
nor U24203 (N_24203,N_23503,N_23918);
nand U24204 (N_24204,N_23792,N_23809);
or U24205 (N_24205,N_23848,N_23831);
and U24206 (N_24206,N_23928,N_23685);
nor U24207 (N_24207,N_23965,N_23877);
or U24208 (N_24208,N_23597,N_23765);
nand U24209 (N_24209,N_23548,N_23721);
nor U24210 (N_24210,N_23547,N_23996);
xnor U24211 (N_24211,N_23609,N_23823);
and U24212 (N_24212,N_23527,N_23666);
or U24213 (N_24213,N_23739,N_23747);
nor U24214 (N_24214,N_23558,N_23896);
nand U24215 (N_24215,N_23906,N_23736);
or U24216 (N_24216,N_23905,N_23673);
and U24217 (N_24217,N_23506,N_23943);
and U24218 (N_24218,N_23528,N_23970);
xnor U24219 (N_24219,N_23564,N_23821);
nand U24220 (N_24220,N_23825,N_23686);
or U24221 (N_24221,N_23781,N_23783);
and U24222 (N_24222,N_23897,N_23541);
xnor U24223 (N_24223,N_23708,N_23696);
nand U24224 (N_24224,N_23946,N_23743);
or U24225 (N_24225,N_23601,N_23659);
xnor U24226 (N_24226,N_23883,N_23745);
and U24227 (N_24227,N_23646,N_23973);
nand U24228 (N_24228,N_23723,N_23951);
nor U24229 (N_24229,N_23604,N_23562);
and U24230 (N_24230,N_23775,N_23935);
nor U24231 (N_24231,N_23812,N_23657);
and U24232 (N_24232,N_23772,N_23645);
or U24233 (N_24233,N_23581,N_23622);
or U24234 (N_24234,N_23518,N_23524);
nor U24235 (N_24235,N_23531,N_23949);
xnor U24236 (N_24236,N_23786,N_23958);
nor U24237 (N_24237,N_23602,N_23568);
nor U24238 (N_24238,N_23587,N_23941);
and U24239 (N_24239,N_23626,N_23630);
nand U24240 (N_24240,N_23557,N_23855);
and U24241 (N_24241,N_23804,N_23571);
nor U24242 (N_24242,N_23516,N_23947);
and U24243 (N_24243,N_23894,N_23917);
or U24244 (N_24244,N_23598,N_23824);
and U24245 (N_24245,N_23914,N_23655);
xor U24246 (N_24246,N_23539,N_23690);
nor U24247 (N_24247,N_23667,N_23607);
or U24248 (N_24248,N_23830,N_23641);
or U24249 (N_24249,N_23880,N_23711);
xor U24250 (N_24250,N_23904,N_23730);
nor U24251 (N_24251,N_23883,N_23785);
or U24252 (N_24252,N_23521,N_23931);
xnor U24253 (N_24253,N_23897,N_23772);
and U24254 (N_24254,N_23626,N_23684);
nand U24255 (N_24255,N_23999,N_23531);
nor U24256 (N_24256,N_23942,N_23814);
nor U24257 (N_24257,N_23655,N_23701);
and U24258 (N_24258,N_23649,N_23729);
nor U24259 (N_24259,N_23794,N_23687);
xor U24260 (N_24260,N_23573,N_23727);
nor U24261 (N_24261,N_23870,N_23639);
nor U24262 (N_24262,N_23992,N_23765);
nand U24263 (N_24263,N_23977,N_23842);
nand U24264 (N_24264,N_23727,N_23837);
nand U24265 (N_24265,N_23519,N_23966);
nand U24266 (N_24266,N_23927,N_23912);
xnor U24267 (N_24267,N_23656,N_23634);
and U24268 (N_24268,N_23609,N_23906);
nor U24269 (N_24269,N_23761,N_23827);
nand U24270 (N_24270,N_23820,N_23602);
nor U24271 (N_24271,N_23554,N_23743);
xnor U24272 (N_24272,N_23973,N_23590);
or U24273 (N_24273,N_23570,N_23653);
nand U24274 (N_24274,N_23973,N_23570);
or U24275 (N_24275,N_23908,N_23819);
and U24276 (N_24276,N_23943,N_23707);
or U24277 (N_24277,N_23973,N_23955);
xnor U24278 (N_24278,N_23632,N_23908);
and U24279 (N_24279,N_23890,N_23626);
xor U24280 (N_24280,N_23760,N_23914);
and U24281 (N_24281,N_23833,N_23511);
nand U24282 (N_24282,N_23990,N_23658);
xor U24283 (N_24283,N_23927,N_23984);
nor U24284 (N_24284,N_23933,N_23523);
nor U24285 (N_24285,N_23716,N_23549);
xnor U24286 (N_24286,N_23833,N_23972);
or U24287 (N_24287,N_23752,N_23956);
xnor U24288 (N_24288,N_23851,N_23996);
nand U24289 (N_24289,N_23639,N_23607);
and U24290 (N_24290,N_23575,N_23556);
or U24291 (N_24291,N_23826,N_23725);
and U24292 (N_24292,N_23545,N_23514);
or U24293 (N_24293,N_23707,N_23831);
nor U24294 (N_24294,N_23835,N_23634);
nand U24295 (N_24295,N_23644,N_23687);
xnor U24296 (N_24296,N_23938,N_23842);
nand U24297 (N_24297,N_23701,N_23529);
or U24298 (N_24298,N_23599,N_23607);
nor U24299 (N_24299,N_23716,N_23588);
xor U24300 (N_24300,N_23925,N_23691);
nand U24301 (N_24301,N_23587,N_23588);
and U24302 (N_24302,N_23928,N_23977);
or U24303 (N_24303,N_23650,N_23723);
nand U24304 (N_24304,N_23968,N_23569);
nand U24305 (N_24305,N_23634,N_23806);
xor U24306 (N_24306,N_23688,N_23652);
and U24307 (N_24307,N_23511,N_23524);
or U24308 (N_24308,N_23786,N_23874);
or U24309 (N_24309,N_23754,N_23582);
xnor U24310 (N_24310,N_23955,N_23680);
and U24311 (N_24311,N_23920,N_23704);
or U24312 (N_24312,N_23668,N_23637);
xor U24313 (N_24313,N_23951,N_23560);
and U24314 (N_24314,N_23568,N_23854);
and U24315 (N_24315,N_23565,N_23883);
or U24316 (N_24316,N_23992,N_23526);
and U24317 (N_24317,N_23727,N_23916);
nor U24318 (N_24318,N_23674,N_23689);
xor U24319 (N_24319,N_23756,N_23996);
nand U24320 (N_24320,N_23711,N_23766);
or U24321 (N_24321,N_23702,N_23667);
or U24322 (N_24322,N_23955,N_23745);
or U24323 (N_24323,N_23682,N_23582);
nand U24324 (N_24324,N_23848,N_23898);
and U24325 (N_24325,N_23727,N_23990);
nor U24326 (N_24326,N_23800,N_23736);
nand U24327 (N_24327,N_23950,N_23985);
nand U24328 (N_24328,N_23781,N_23518);
or U24329 (N_24329,N_23950,N_23880);
nand U24330 (N_24330,N_23506,N_23982);
or U24331 (N_24331,N_23821,N_23994);
and U24332 (N_24332,N_23998,N_23919);
and U24333 (N_24333,N_23791,N_23741);
and U24334 (N_24334,N_23938,N_23945);
xnor U24335 (N_24335,N_23712,N_23871);
or U24336 (N_24336,N_23990,N_23756);
nand U24337 (N_24337,N_23675,N_23688);
nand U24338 (N_24338,N_23707,N_23630);
and U24339 (N_24339,N_23927,N_23875);
or U24340 (N_24340,N_23941,N_23630);
or U24341 (N_24341,N_23878,N_23836);
or U24342 (N_24342,N_23751,N_23898);
and U24343 (N_24343,N_23782,N_23639);
or U24344 (N_24344,N_23714,N_23972);
xnor U24345 (N_24345,N_23564,N_23863);
or U24346 (N_24346,N_23511,N_23703);
or U24347 (N_24347,N_23568,N_23643);
nand U24348 (N_24348,N_23626,N_23606);
or U24349 (N_24349,N_23937,N_23909);
nand U24350 (N_24350,N_23691,N_23556);
xor U24351 (N_24351,N_23773,N_23949);
or U24352 (N_24352,N_23807,N_23615);
nand U24353 (N_24353,N_23758,N_23687);
or U24354 (N_24354,N_23976,N_23553);
or U24355 (N_24355,N_23537,N_23773);
or U24356 (N_24356,N_23516,N_23555);
or U24357 (N_24357,N_23519,N_23553);
nor U24358 (N_24358,N_23963,N_23828);
nand U24359 (N_24359,N_23650,N_23586);
nand U24360 (N_24360,N_23621,N_23699);
and U24361 (N_24361,N_23933,N_23831);
xnor U24362 (N_24362,N_23665,N_23569);
nor U24363 (N_24363,N_23867,N_23820);
xor U24364 (N_24364,N_23900,N_23655);
xor U24365 (N_24365,N_23836,N_23734);
and U24366 (N_24366,N_23688,N_23908);
nor U24367 (N_24367,N_23652,N_23580);
nor U24368 (N_24368,N_23981,N_23825);
nand U24369 (N_24369,N_23630,N_23817);
nor U24370 (N_24370,N_23682,N_23520);
xor U24371 (N_24371,N_23532,N_23540);
nor U24372 (N_24372,N_23517,N_23503);
and U24373 (N_24373,N_23612,N_23566);
nor U24374 (N_24374,N_23584,N_23645);
or U24375 (N_24375,N_23858,N_23866);
xnor U24376 (N_24376,N_23727,N_23623);
nand U24377 (N_24377,N_23677,N_23562);
nand U24378 (N_24378,N_23594,N_23551);
or U24379 (N_24379,N_23652,N_23662);
nand U24380 (N_24380,N_23761,N_23883);
nand U24381 (N_24381,N_23649,N_23614);
nand U24382 (N_24382,N_23605,N_23722);
or U24383 (N_24383,N_23645,N_23501);
nand U24384 (N_24384,N_23754,N_23891);
or U24385 (N_24385,N_23558,N_23623);
nand U24386 (N_24386,N_23766,N_23616);
nor U24387 (N_24387,N_23541,N_23743);
xnor U24388 (N_24388,N_23810,N_23824);
xnor U24389 (N_24389,N_23816,N_23621);
nand U24390 (N_24390,N_23705,N_23756);
and U24391 (N_24391,N_23742,N_23806);
nor U24392 (N_24392,N_23963,N_23600);
nor U24393 (N_24393,N_23657,N_23935);
nor U24394 (N_24394,N_23805,N_23603);
nor U24395 (N_24395,N_23942,N_23990);
nand U24396 (N_24396,N_23659,N_23762);
or U24397 (N_24397,N_23611,N_23652);
nand U24398 (N_24398,N_23530,N_23548);
and U24399 (N_24399,N_23710,N_23969);
and U24400 (N_24400,N_23709,N_23954);
or U24401 (N_24401,N_23761,N_23735);
nand U24402 (N_24402,N_23622,N_23990);
nor U24403 (N_24403,N_23585,N_23972);
nand U24404 (N_24404,N_23791,N_23699);
xnor U24405 (N_24405,N_23908,N_23544);
and U24406 (N_24406,N_23638,N_23814);
nor U24407 (N_24407,N_23793,N_23534);
and U24408 (N_24408,N_23717,N_23628);
nand U24409 (N_24409,N_23947,N_23641);
xor U24410 (N_24410,N_23777,N_23633);
or U24411 (N_24411,N_23732,N_23857);
xnor U24412 (N_24412,N_23888,N_23836);
nor U24413 (N_24413,N_23605,N_23534);
or U24414 (N_24414,N_23683,N_23836);
nand U24415 (N_24415,N_23553,N_23506);
nand U24416 (N_24416,N_23877,N_23564);
xor U24417 (N_24417,N_23951,N_23749);
and U24418 (N_24418,N_23572,N_23566);
xor U24419 (N_24419,N_23513,N_23955);
and U24420 (N_24420,N_23909,N_23987);
or U24421 (N_24421,N_23727,N_23564);
and U24422 (N_24422,N_23876,N_23653);
and U24423 (N_24423,N_23736,N_23920);
and U24424 (N_24424,N_23538,N_23902);
or U24425 (N_24425,N_23924,N_23836);
and U24426 (N_24426,N_23725,N_23578);
xor U24427 (N_24427,N_23567,N_23601);
and U24428 (N_24428,N_23650,N_23868);
or U24429 (N_24429,N_23726,N_23777);
xnor U24430 (N_24430,N_23672,N_23703);
or U24431 (N_24431,N_23532,N_23698);
and U24432 (N_24432,N_23694,N_23533);
and U24433 (N_24433,N_23743,N_23650);
xor U24434 (N_24434,N_23512,N_23789);
and U24435 (N_24435,N_23511,N_23567);
or U24436 (N_24436,N_23767,N_23997);
nor U24437 (N_24437,N_23761,N_23601);
xor U24438 (N_24438,N_23967,N_23587);
nand U24439 (N_24439,N_23724,N_23552);
nand U24440 (N_24440,N_23578,N_23879);
and U24441 (N_24441,N_23568,N_23982);
or U24442 (N_24442,N_23791,N_23640);
nand U24443 (N_24443,N_23585,N_23537);
or U24444 (N_24444,N_23929,N_23811);
nor U24445 (N_24445,N_23772,N_23563);
or U24446 (N_24446,N_23553,N_23803);
xnor U24447 (N_24447,N_23804,N_23831);
nand U24448 (N_24448,N_23996,N_23562);
nor U24449 (N_24449,N_23884,N_23730);
xor U24450 (N_24450,N_23965,N_23533);
and U24451 (N_24451,N_23572,N_23527);
xor U24452 (N_24452,N_23723,N_23821);
nor U24453 (N_24453,N_23780,N_23802);
or U24454 (N_24454,N_23927,N_23660);
and U24455 (N_24455,N_23762,N_23920);
or U24456 (N_24456,N_23588,N_23697);
nand U24457 (N_24457,N_23507,N_23537);
xor U24458 (N_24458,N_23685,N_23752);
xor U24459 (N_24459,N_23521,N_23523);
nor U24460 (N_24460,N_23535,N_23564);
xnor U24461 (N_24461,N_23544,N_23920);
xor U24462 (N_24462,N_23530,N_23699);
xor U24463 (N_24463,N_23601,N_23558);
or U24464 (N_24464,N_23764,N_23999);
nand U24465 (N_24465,N_23575,N_23589);
or U24466 (N_24466,N_23856,N_23549);
nand U24467 (N_24467,N_23898,N_23728);
or U24468 (N_24468,N_23936,N_23848);
nor U24469 (N_24469,N_23970,N_23782);
or U24470 (N_24470,N_23970,N_23705);
and U24471 (N_24471,N_23995,N_23821);
nor U24472 (N_24472,N_23959,N_23751);
xnor U24473 (N_24473,N_23802,N_23676);
or U24474 (N_24474,N_23571,N_23699);
xnor U24475 (N_24475,N_23707,N_23788);
xor U24476 (N_24476,N_23994,N_23697);
xnor U24477 (N_24477,N_23789,N_23994);
and U24478 (N_24478,N_23948,N_23509);
xnor U24479 (N_24479,N_23965,N_23637);
nand U24480 (N_24480,N_23624,N_23831);
nand U24481 (N_24481,N_23540,N_23691);
nand U24482 (N_24482,N_23800,N_23780);
xor U24483 (N_24483,N_23621,N_23793);
or U24484 (N_24484,N_23817,N_23536);
nor U24485 (N_24485,N_23588,N_23725);
nor U24486 (N_24486,N_23646,N_23746);
nand U24487 (N_24487,N_23561,N_23884);
or U24488 (N_24488,N_23608,N_23621);
xor U24489 (N_24489,N_23943,N_23933);
xor U24490 (N_24490,N_23809,N_23728);
nor U24491 (N_24491,N_23775,N_23563);
xor U24492 (N_24492,N_23795,N_23975);
xnor U24493 (N_24493,N_23574,N_23875);
xor U24494 (N_24494,N_23661,N_23936);
or U24495 (N_24495,N_23948,N_23512);
xnor U24496 (N_24496,N_23628,N_23542);
and U24497 (N_24497,N_23687,N_23779);
and U24498 (N_24498,N_23909,N_23784);
or U24499 (N_24499,N_23816,N_23687);
or U24500 (N_24500,N_24087,N_24218);
or U24501 (N_24501,N_24134,N_24421);
xor U24502 (N_24502,N_24227,N_24092);
or U24503 (N_24503,N_24058,N_24033);
or U24504 (N_24504,N_24283,N_24246);
nor U24505 (N_24505,N_24075,N_24106);
nand U24506 (N_24506,N_24153,N_24312);
or U24507 (N_24507,N_24128,N_24279);
xnor U24508 (N_24508,N_24047,N_24369);
nor U24509 (N_24509,N_24298,N_24146);
or U24510 (N_24510,N_24456,N_24014);
xor U24511 (N_24511,N_24296,N_24322);
and U24512 (N_24512,N_24142,N_24301);
xor U24513 (N_24513,N_24090,N_24072);
nor U24514 (N_24514,N_24374,N_24193);
and U24515 (N_24515,N_24306,N_24163);
and U24516 (N_24516,N_24052,N_24171);
and U24517 (N_24517,N_24310,N_24044);
nand U24518 (N_24518,N_24045,N_24414);
or U24519 (N_24519,N_24156,N_24139);
nand U24520 (N_24520,N_24049,N_24416);
nand U24521 (N_24521,N_24140,N_24463);
xor U24522 (N_24522,N_24173,N_24332);
xnor U24523 (N_24523,N_24431,N_24239);
nor U24524 (N_24524,N_24459,N_24125);
and U24525 (N_24525,N_24133,N_24401);
nand U24526 (N_24526,N_24483,N_24126);
and U24527 (N_24527,N_24390,N_24223);
or U24528 (N_24528,N_24215,N_24340);
and U24529 (N_24529,N_24445,N_24064);
nand U24530 (N_24530,N_24222,N_24138);
or U24531 (N_24531,N_24288,N_24285);
and U24532 (N_24532,N_24229,N_24041);
and U24533 (N_24533,N_24260,N_24023);
or U24534 (N_24534,N_24268,N_24162);
nor U24535 (N_24535,N_24497,N_24417);
nor U24536 (N_24536,N_24355,N_24358);
nand U24537 (N_24537,N_24124,N_24247);
and U24538 (N_24538,N_24315,N_24429);
nor U24539 (N_24539,N_24293,N_24253);
xnor U24540 (N_24540,N_24423,N_24099);
or U24541 (N_24541,N_24011,N_24016);
nand U24542 (N_24542,N_24377,N_24078);
xnor U24543 (N_24543,N_24337,N_24498);
xor U24544 (N_24544,N_24378,N_24418);
nand U24545 (N_24545,N_24206,N_24149);
nor U24546 (N_24546,N_24034,N_24096);
xor U24547 (N_24547,N_24453,N_24376);
xnor U24548 (N_24548,N_24076,N_24110);
nand U24549 (N_24549,N_24307,N_24244);
nor U24550 (N_24550,N_24342,N_24385);
and U24551 (N_24551,N_24339,N_24480);
or U24552 (N_24552,N_24176,N_24172);
nor U24553 (N_24553,N_24074,N_24018);
or U24554 (N_24554,N_24238,N_24248);
nor U24555 (N_24555,N_24136,N_24028);
nor U24556 (N_24556,N_24413,N_24084);
or U24557 (N_24557,N_24115,N_24422);
or U24558 (N_24558,N_24079,N_24294);
nand U24559 (N_24559,N_24119,N_24321);
and U24560 (N_24560,N_24118,N_24179);
xnor U24561 (N_24561,N_24302,N_24123);
nor U24562 (N_24562,N_24211,N_24365);
nand U24563 (N_24563,N_24435,N_24353);
nor U24564 (N_24564,N_24132,N_24205);
xor U24565 (N_24565,N_24252,N_24000);
and U24566 (N_24566,N_24392,N_24344);
xor U24567 (N_24567,N_24187,N_24207);
nor U24568 (N_24568,N_24001,N_24221);
and U24569 (N_24569,N_24089,N_24212);
or U24570 (N_24570,N_24116,N_24462);
nor U24571 (N_24571,N_24346,N_24236);
nand U24572 (N_24572,N_24281,N_24166);
and U24573 (N_24573,N_24448,N_24408);
xnor U24574 (N_24574,N_24083,N_24261);
and U24575 (N_24575,N_24224,N_24046);
nor U24576 (N_24576,N_24277,N_24237);
nand U24577 (N_24577,N_24481,N_24190);
xor U24578 (N_24578,N_24476,N_24402);
nor U24579 (N_24579,N_24254,N_24325);
or U24580 (N_24580,N_24270,N_24061);
nor U24581 (N_24581,N_24466,N_24347);
and U24582 (N_24582,N_24318,N_24164);
and U24583 (N_24583,N_24407,N_24330);
nand U24584 (N_24584,N_24487,N_24005);
nor U24585 (N_24585,N_24472,N_24366);
xor U24586 (N_24586,N_24305,N_24495);
and U24587 (N_24587,N_24471,N_24251);
and U24588 (N_24588,N_24372,N_24428);
and U24589 (N_24589,N_24051,N_24059);
or U24590 (N_24590,N_24112,N_24147);
xor U24591 (N_24591,N_24313,N_24181);
or U24592 (N_24592,N_24220,N_24002);
and U24593 (N_24593,N_24452,N_24454);
nand U24594 (N_24594,N_24160,N_24067);
xnor U24595 (N_24595,N_24255,N_24286);
and U24596 (N_24596,N_24314,N_24333);
xor U24597 (N_24597,N_24444,N_24077);
xnor U24598 (N_24598,N_24434,N_24424);
nor U24599 (N_24599,N_24289,N_24108);
xor U24600 (N_24600,N_24437,N_24157);
or U24601 (N_24601,N_24432,N_24183);
or U24602 (N_24602,N_24299,N_24042);
nand U24603 (N_24603,N_24451,N_24264);
nor U24604 (N_24604,N_24290,N_24039);
or U24605 (N_24605,N_24219,N_24331);
nand U24606 (N_24606,N_24109,N_24175);
nor U24607 (N_24607,N_24027,N_24391);
xnor U24608 (N_24608,N_24113,N_24216);
and U24609 (N_24609,N_24273,N_24240);
or U24610 (N_24610,N_24383,N_24213);
nand U24611 (N_24611,N_24209,N_24017);
nand U24612 (N_24612,N_24103,N_24271);
or U24613 (N_24613,N_24419,N_24159);
xor U24614 (N_24614,N_24121,N_24282);
and U24615 (N_24615,N_24478,N_24371);
nor U24616 (N_24616,N_24105,N_24415);
and U24617 (N_24617,N_24150,N_24488);
or U24618 (N_24618,N_24029,N_24447);
nor U24619 (N_24619,N_24093,N_24359);
or U24620 (N_24620,N_24026,N_24102);
and U24621 (N_24621,N_24405,N_24329);
and U24622 (N_24622,N_24111,N_24309);
nor U24623 (N_24623,N_24430,N_24354);
xnor U24624 (N_24624,N_24461,N_24040);
xor U24625 (N_24625,N_24272,N_24137);
xor U24626 (N_24626,N_24019,N_24024);
and U24627 (N_24627,N_24086,N_24069);
nor U24628 (N_24628,N_24228,N_24465);
nor U24629 (N_24629,N_24335,N_24085);
xor U24630 (N_24630,N_24122,N_24144);
nor U24631 (N_24631,N_24154,N_24152);
or U24632 (N_24632,N_24436,N_24441);
nor U24633 (N_24633,N_24263,N_24449);
and U24634 (N_24634,N_24311,N_24217);
xnor U24635 (N_24635,N_24012,N_24101);
and U24636 (N_24636,N_24182,N_24097);
and U24637 (N_24637,N_24233,N_24158);
xnor U24638 (N_24638,N_24174,N_24384);
nand U24639 (N_24639,N_24258,N_24323);
nor U24640 (N_24640,N_24155,N_24245);
xnor U24641 (N_24641,N_24393,N_24007);
nor U24642 (N_24642,N_24492,N_24013);
nand U24643 (N_24643,N_24100,N_24485);
and U24644 (N_24644,N_24010,N_24491);
nor U24645 (N_24645,N_24180,N_24457);
and U24646 (N_24646,N_24243,N_24479);
and U24647 (N_24647,N_24095,N_24030);
nand U24648 (N_24648,N_24278,N_24203);
nand U24649 (N_24649,N_24235,N_24396);
nor U24650 (N_24650,N_24326,N_24357);
and U24651 (N_24651,N_24370,N_24427);
or U24652 (N_24652,N_24364,N_24367);
and U24653 (N_24653,N_24231,N_24470);
and U24654 (N_24654,N_24360,N_24053);
xnor U24655 (N_24655,N_24328,N_24442);
nand U24656 (N_24656,N_24494,N_24208);
nand U24657 (N_24657,N_24015,N_24184);
or U24658 (N_24658,N_24386,N_24161);
xor U24659 (N_24659,N_24398,N_24382);
and U24660 (N_24660,N_24343,N_24114);
nand U24661 (N_24661,N_24274,N_24199);
nor U24662 (N_24662,N_24308,N_24300);
nand U24663 (N_24663,N_24141,N_24275);
nor U24664 (N_24664,N_24256,N_24022);
xnor U24665 (N_24665,N_24189,N_24048);
nor U24666 (N_24666,N_24130,N_24458);
and U24667 (N_24667,N_24127,N_24440);
nor U24668 (N_24668,N_24167,N_24433);
and U24669 (N_24669,N_24259,N_24151);
or U24670 (N_24670,N_24484,N_24284);
and U24671 (N_24671,N_24129,N_24350);
nand U24672 (N_24672,N_24412,N_24295);
nand U24673 (N_24673,N_24406,N_24426);
or U24674 (N_24674,N_24020,N_24241);
or U24675 (N_24675,N_24320,N_24063);
xnor U24676 (N_24676,N_24473,N_24071);
xnor U24677 (N_24677,N_24474,N_24352);
and U24678 (N_24678,N_24368,N_24410);
nor U24679 (N_24679,N_24185,N_24351);
xor U24680 (N_24680,N_24009,N_24450);
xnor U24681 (N_24681,N_24204,N_24165);
xnor U24682 (N_24682,N_24081,N_24266);
and U24683 (N_24683,N_24008,N_24006);
or U24684 (N_24684,N_24265,N_24066);
nand U24685 (N_24685,N_24361,N_24334);
xnor U24686 (N_24686,N_24276,N_24191);
nand U24687 (N_24687,N_24094,N_24131);
or U24688 (N_24688,N_24356,N_24198);
xor U24689 (N_24689,N_24316,N_24338);
and U24690 (N_24690,N_24091,N_24196);
nor U24691 (N_24691,N_24345,N_24003);
nand U24692 (N_24692,N_24168,N_24327);
and U24693 (N_24693,N_24395,N_24055);
nand U24694 (N_24694,N_24201,N_24186);
nand U24695 (N_24695,N_24057,N_24060);
nand U24696 (N_24696,N_24135,N_24192);
and U24697 (N_24697,N_24467,N_24249);
nor U24698 (N_24698,N_24036,N_24230);
nor U24699 (N_24699,N_24032,N_24194);
nor U24700 (N_24700,N_24280,N_24303);
xor U24701 (N_24701,N_24065,N_24287);
or U24702 (N_24702,N_24037,N_24399);
or U24703 (N_24703,N_24070,N_24490);
or U24704 (N_24704,N_24225,N_24088);
xor U24705 (N_24705,N_24496,N_24242);
xnor U24706 (N_24706,N_24202,N_24319);
and U24707 (N_24707,N_24304,N_24297);
nand U24708 (N_24708,N_24317,N_24439);
xnor U24709 (N_24709,N_24397,N_24043);
xnor U24710 (N_24710,N_24292,N_24438);
nor U24711 (N_24711,N_24460,N_24050);
nand U24712 (N_24712,N_24362,N_24403);
nand U24713 (N_24713,N_24269,N_24262);
nand U24714 (N_24714,N_24250,N_24486);
or U24715 (N_24715,N_24468,N_24054);
xnor U24716 (N_24716,N_24336,N_24232);
nor U24717 (N_24717,N_24062,N_24031);
nand U24718 (N_24718,N_24420,N_24143);
and U24719 (N_24719,N_24200,N_24080);
and U24720 (N_24720,N_24082,N_24475);
and U24721 (N_24721,N_24145,N_24499);
and U24722 (N_24722,N_24464,N_24170);
nand U24723 (N_24723,N_24341,N_24379);
and U24724 (N_24724,N_24446,N_24493);
nor U24725 (N_24725,N_24195,N_24349);
nor U24726 (N_24726,N_24469,N_24120);
xor U24727 (N_24727,N_24098,N_24400);
xnor U24728 (N_24728,N_24169,N_24394);
or U24729 (N_24729,N_24226,N_24363);
nor U24730 (N_24730,N_24409,N_24068);
and U24731 (N_24731,N_24257,N_24178);
nand U24732 (N_24732,N_24489,N_24188);
or U24733 (N_24733,N_24056,N_24388);
nor U24734 (N_24734,N_24482,N_24348);
or U24735 (N_24735,N_24177,N_24117);
xor U24736 (N_24736,N_24107,N_24375);
xnor U24737 (N_24737,N_24373,N_24234);
xnor U24738 (N_24738,N_24291,N_24148);
xor U24739 (N_24739,N_24404,N_24380);
xnor U24740 (N_24740,N_24387,N_24267);
nor U24741 (N_24741,N_24025,N_24411);
nand U24742 (N_24742,N_24210,N_24425);
and U24743 (N_24743,N_24021,N_24477);
or U24744 (N_24744,N_24214,N_24324);
xor U24745 (N_24745,N_24035,N_24381);
nand U24746 (N_24746,N_24197,N_24455);
nand U24747 (N_24747,N_24104,N_24073);
and U24748 (N_24748,N_24389,N_24038);
nand U24749 (N_24749,N_24443,N_24004);
or U24750 (N_24750,N_24370,N_24476);
nand U24751 (N_24751,N_24203,N_24243);
or U24752 (N_24752,N_24193,N_24002);
nor U24753 (N_24753,N_24149,N_24163);
or U24754 (N_24754,N_24384,N_24187);
and U24755 (N_24755,N_24386,N_24447);
xor U24756 (N_24756,N_24324,N_24054);
nand U24757 (N_24757,N_24305,N_24399);
nand U24758 (N_24758,N_24006,N_24495);
or U24759 (N_24759,N_24198,N_24377);
xnor U24760 (N_24760,N_24004,N_24213);
and U24761 (N_24761,N_24267,N_24309);
and U24762 (N_24762,N_24421,N_24419);
and U24763 (N_24763,N_24361,N_24146);
nand U24764 (N_24764,N_24376,N_24448);
or U24765 (N_24765,N_24282,N_24483);
nand U24766 (N_24766,N_24208,N_24240);
xor U24767 (N_24767,N_24320,N_24382);
or U24768 (N_24768,N_24413,N_24137);
nor U24769 (N_24769,N_24385,N_24269);
xor U24770 (N_24770,N_24317,N_24206);
nor U24771 (N_24771,N_24331,N_24210);
nor U24772 (N_24772,N_24374,N_24021);
or U24773 (N_24773,N_24168,N_24084);
nor U24774 (N_24774,N_24378,N_24230);
and U24775 (N_24775,N_24163,N_24464);
xnor U24776 (N_24776,N_24361,N_24319);
and U24777 (N_24777,N_24082,N_24314);
nor U24778 (N_24778,N_24017,N_24161);
or U24779 (N_24779,N_24256,N_24237);
nor U24780 (N_24780,N_24379,N_24161);
xnor U24781 (N_24781,N_24100,N_24352);
nand U24782 (N_24782,N_24203,N_24008);
and U24783 (N_24783,N_24115,N_24128);
nand U24784 (N_24784,N_24057,N_24332);
xor U24785 (N_24785,N_24461,N_24289);
nor U24786 (N_24786,N_24004,N_24034);
nor U24787 (N_24787,N_24204,N_24231);
xnor U24788 (N_24788,N_24476,N_24368);
xor U24789 (N_24789,N_24116,N_24299);
and U24790 (N_24790,N_24446,N_24371);
nand U24791 (N_24791,N_24442,N_24287);
xor U24792 (N_24792,N_24181,N_24392);
and U24793 (N_24793,N_24191,N_24360);
and U24794 (N_24794,N_24082,N_24175);
nor U24795 (N_24795,N_24030,N_24484);
or U24796 (N_24796,N_24273,N_24109);
or U24797 (N_24797,N_24428,N_24357);
or U24798 (N_24798,N_24359,N_24444);
xnor U24799 (N_24799,N_24320,N_24094);
nor U24800 (N_24800,N_24366,N_24099);
nor U24801 (N_24801,N_24112,N_24437);
nor U24802 (N_24802,N_24449,N_24170);
nand U24803 (N_24803,N_24186,N_24013);
or U24804 (N_24804,N_24314,N_24419);
nand U24805 (N_24805,N_24075,N_24300);
xnor U24806 (N_24806,N_24005,N_24379);
and U24807 (N_24807,N_24055,N_24248);
nor U24808 (N_24808,N_24061,N_24224);
nor U24809 (N_24809,N_24495,N_24161);
nor U24810 (N_24810,N_24319,N_24359);
and U24811 (N_24811,N_24470,N_24361);
xnor U24812 (N_24812,N_24255,N_24414);
xnor U24813 (N_24813,N_24104,N_24152);
and U24814 (N_24814,N_24111,N_24303);
xnor U24815 (N_24815,N_24014,N_24108);
or U24816 (N_24816,N_24333,N_24082);
nand U24817 (N_24817,N_24450,N_24173);
nor U24818 (N_24818,N_24453,N_24067);
nor U24819 (N_24819,N_24481,N_24311);
nor U24820 (N_24820,N_24383,N_24360);
xor U24821 (N_24821,N_24468,N_24318);
xor U24822 (N_24822,N_24362,N_24295);
xor U24823 (N_24823,N_24381,N_24362);
xnor U24824 (N_24824,N_24339,N_24030);
xor U24825 (N_24825,N_24453,N_24035);
or U24826 (N_24826,N_24320,N_24013);
or U24827 (N_24827,N_24082,N_24376);
nand U24828 (N_24828,N_24313,N_24318);
nand U24829 (N_24829,N_24140,N_24219);
and U24830 (N_24830,N_24084,N_24469);
and U24831 (N_24831,N_24003,N_24067);
nand U24832 (N_24832,N_24052,N_24207);
xor U24833 (N_24833,N_24182,N_24491);
nor U24834 (N_24834,N_24476,N_24401);
and U24835 (N_24835,N_24126,N_24273);
and U24836 (N_24836,N_24485,N_24239);
or U24837 (N_24837,N_24100,N_24126);
xnor U24838 (N_24838,N_24290,N_24425);
nor U24839 (N_24839,N_24153,N_24304);
xnor U24840 (N_24840,N_24231,N_24004);
or U24841 (N_24841,N_24460,N_24486);
or U24842 (N_24842,N_24402,N_24438);
nor U24843 (N_24843,N_24233,N_24240);
nand U24844 (N_24844,N_24221,N_24078);
xor U24845 (N_24845,N_24011,N_24167);
or U24846 (N_24846,N_24409,N_24259);
nand U24847 (N_24847,N_24456,N_24096);
nand U24848 (N_24848,N_24079,N_24210);
xor U24849 (N_24849,N_24020,N_24193);
nand U24850 (N_24850,N_24465,N_24341);
or U24851 (N_24851,N_24221,N_24486);
and U24852 (N_24852,N_24011,N_24213);
nand U24853 (N_24853,N_24014,N_24337);
or U24854 (N_24854,N_24177,N_24118);
nor U24855 (N_24855,N_24021,N_24479);
or U24856 (N_24856,N_24467,N_24176);
xor U24857 (N_24857,N_24475,N_24424);
xor U24858 (N_24858,N_24070,N_24341);
xor U24859 (N_24859,N_24490,N_24027);
nand U24860 (N_24860,N_24481,N_24074);
and U24861 (N_24861,N_24223,N_24437);
and U24862 (N_24862,N_24209,N_24021);
and U24863 (N_24863,N_24368,N_24214);
xnor U24864 (N_24864,N_24483,N_24481);
and U24865 (N_24865,N_24092,N_24013);
nor U24866 (N_24866,N_24017,N_24405);
and U24867 (N_24867,N_24022,N_24484);
xnor U24868 (N_24868,N_24263,N_24340);
xnor U24869 (N_24869,N_24114,N_24390);
and U24870 (N_24870,N_24175,N_24140);
nor U24871 (N_24871,N_24393,N_24351);
xnor U24872 (N_24872,N_24005,N_24475);
nand U24873 (N_24873,N_24015,N_24401);
nor U24874 (N_24874,N_24377,N_24444);
or U24875 (N_24875,N_24423,N_24095);
and U24876 (N_24876,N_24268,N_24294);
and U24877 (N_24877,N_24461,N_24184);
nand U24878 (N_24878,N_24444,N_24447);
nand U24879 (N_24879,N_24076,N_24099);
or U24880 (N_24880,N_24435,N_24285);
and U24881 (N_24881,N_24146,N_24255);
and U24882 (N_24882,N_24258,N_24157);
nor U24883 (N_24883,N_24078,N_24486);
nor U24884 (N_24884,N_24401,N_24408);
or U24885 (N_24885,N_24050,N_24254);
or U24886 (N_24886,N_24303,N_24334);
nor U24887 (N_24887,N_24236,N_24415);
and U24888 (N_24888,N_24409,N_24191);
and U24889 (N_24889,N_24070,N_24363);
nor U24890 (N_24890,N_24252,N_24351);
nor U24891 (N_24891,N_24361,N_24291);
and U24892 (N_24892,N_24348,N_24406);
and U24893 (N_24893,N_24259,N_24161);
nor U24894 (N_24894,N_24149,N_24302);
and U24895 (N_24895,N_24460,N_24492);
and U24896 (N_24896,N_24374,N_24161);
nor U24897 (N_24897,N_24196,N_24170);
xor U24898 (N_24898,N_24152,N_24264);
or U24899 (N_24899,N_24489,N_24494);
nand U24900 (N_24900,N_24050,N_24445);
xor U24901 (N_24901,N_24404,N_24206);
xnor U24902 (N_24902,N_24300,N_24367);
or U24903 (N_24903,N_24052,N_24154);
or U24904 (N_24904,N_24441,N_24342);
or U24905 (N_24905,N_24155,N_24199);
xor U24906 (N_24906,N_24349,N_24219);
nor U24907 (N_24907,N_24216,N_24120);
or U24908 (N_24908,N_24028,N_24498);
nor U24909 (N_24909,N_24024,N_24485);
xor U24910 (N_24910,N_24193,N_24413);
nand U24911 (N_24911,N_24250,N_24186);
nor U24912 (N_24912,N_24435,N_24278);
nor U24913 (N_24913,N_24391,N_24338);
nor U24914 (N_24914,N_24239,N_24451);
nor U24915 (N_24915,N_24144,N_24117);
nor U24916 (N_24916,N_24298,N_24208);
and U24917 (N_24917,N_24249,N_24362);
xnor U24918 (N_24918,N_24098,N_24489);
nor U24919 (N_24919,N_24255,N_24206);
nand U24920 (N_24920,N_24477,N_24240);
or U24921 (N_24921,N_24159,N_24399);
nor U24922 (N_24922,N_24066,N_24401);
and U24923 (N_24923,N_24418,N_24465);
nor U24924 (N_24924,N_24472,N_24425);
xor U24925 (N_24925,N_24269,N_24328);
nor U24926 (N_24926,N_24167,N_24307);
nand U24927 (N_24927,N_24246,N_24160);
and U24928 (N_24928,N_24090,N_24261);
or U24929 (N_24929,N_24046,N_24331);
or U24930 (N_24930,N_24019,N_24162);
and U24931 (N_24931,N_24403,N_24491);
nand U24932 (N_24932,N_24130,N_24378);
nand U24933 (N_24933,N_24084,N_24144);
nor U24934 (N_24934,N_24420,N_24459);
nor U24935 (N_24935,N_24410,N_24022);
nand U24936 (N_24936,N_24244,N_24452);
nand U24937 (N_24937,N_24155,N_24394);
nand U24938 (N_24938,N_24422,N_24198);
nand U24939 (N_24939,N_24402,N_24001);
xnor U24940 (N_24940,N_24381,N_24036);
xor U24941 (N_24941,N_24224,N_24238);
nor U24942 (N_24942,N_24063,N_24161);
and U24943 (N_24943,N_24068,N_24273);
nor U24944 (N_24944,N_24210,N_24048);
nor U24945 (N_24945,N_24213,N_24349);
or U24946 (N_24946,N_24199,N_24012);
nand U24947 (N_24947,N_24121,N_24180);
and U24948 (N_24948,N_24377,N_24312);
nor U24949 (N_24949,N_24009,N_24369);
nand U24950 (N_24950,N_24477,N_24058);
nand U24951 (N_24951,N_24117,N_24160);
xor U24952 (N_24952,N_24412,N_24307);
nor U24953 (N_24953,N_24318,N_24087);
or U24954 (N_24954,N_24287,N_24000);
nor U24955 (N_24955,N_24147,N_24011);
nor U24956 (N_24956,N_24021,N_24460);
xor U24957 (N_24957,N_24363,N_24196);
and U24958 (N_24958,N_24030,N_24272);
nor U24959 (N_24959,N_24209,N_24346);
nand U24960 (N_24960,N_24437,N_24472);
and U24961 (N_24961,N_24223,N_24452);
nor U24962 (N_24962,N_24172,N_24464);
or U24963 (N_24963,N_24095,N_24437);
nor U24964 (N_24964,N_24158,N_24062);
or U24965 (N_24965,N_24033,N_24055);
nand U24966 (N_24966,N_24016,N_24012);
or U24967 (N_24967,N_24470,N_24389);
xnor U24968 (N_24968,N_24463,N_24279);
or U24969 (N_24969,N_24132,N_24098);
nand U24970 (N_24970,N_24395,N_24033);
nand U24971 (N_24971,N_24200,N_24228);
nand U24972 (N_24972,N_24081,N_24296);
xnor U24973 (N_24973,N_24444,N_24333);
and U24974 (N_24974,N_24134,N_24433);
or U24975 (N_24975,N_24037,N_24283);
and U24976 (N_24976,N_24138,N_24315);
or U24977 (N_24977,N_24066,N_24025);
or U24978 (N_24978,N_24242,N_24471);
xnor U24979 (N_24979,N_24193,N_24060);
and U24980 (N_24980,N_24127,N_24409);
and U24981 (N_24981,N_24299,N_24219);
or U24982 (N_24982,N_24460,N_24266);
nand U24983 (N_24983,N_24049,N_24076);
or U24984 (N_24984,N_24444,N_24279);
and U24985 (N_24985,N_24153,N_24093);
or U24986 (N_24986,N_24312,N_24006);
or U24987 (N_24987,N_24329,N_24347);
and U24988 (N_24988,N_24216,N_24191);
nand U24989 (N_24989,N_24249,N_24185);
or U24990 (N_24990,N_24460,N_24271);
and U24991 (N_24991,N_24260,N_24086);
xnor U24992 (N_24992,N_24178,N_24276);
nand U24993 (N_24993,N_24141,N_24185);
xor U24994 (N_24994,N_24344,N_24487);
xnor U24995 (N_24995,N_24076,N_24281);
xor U24996 (N_24996,N_24167,N_24424);
xnor U24997 (N_24997,N_24371,N_24176);
and U24998 (N_24998,N_24224,N_24055);
nor U24999 (N_24999,N_24034,N_24308);
and U25000 (N_25000,N_24757,N_24641);
or U25001 (N_25001,N_24889,N_24514);
and U25002 (N_25002,N_24811,N_24752);
nand U25003 (N_25003,N_24666,N_24942);
or U25004 (N_25004,N_24740,N_24878);
nor U25005 (N_25005,N_24973,N_24772);
and U25006 (N_25006,N_24638,N_24927);
xor U25007 (N_25007,N_24997,N_24901);
or U25008 (N_25008,N_24921,N_24763);
and U25009 (N_25009,N_24711,N_24827);
nand U25010 (N_25010,N_24646,N_24817);
nand U25011 (N_25011,N_24516,N_24855);
and U25012 (N_25012,N_24785,N_24593);
nor U25013 (N_25013,N_24599,N_24939);
and U25014 (N_25014,N_24710,N_24963);
xnor U25015 (N_25015,N_24664,N_24581);
nor U25016 (N_25016,N_24836,N_24911);
or U25017 (N_25017,N_24844,N_24510);
nor U25018 (N_25018,N_24649,N_24934);
or U25019 (N_25019,N_24610,N_24737);
or U25020 (N_25020,N_24764,N_24841);
nand U25021 (N_25021,N_24854,N_24789);
and U25022 (N_25022,N_24684,N_24578);
xor U25023 (N_25023,N_24801,N_24794);
nor U25024 (N_25024,N_24781,N_24637);
or U25025 (N_25025,N_24598,N_24659);
or U25026 (N_25026,N_24832,N_24777);
nor U25027 (N_25027,N_24948,N_24550);
xor U25028 (N_25028,N_24813,N_24962);
nor U25029 (N_25029,N_24651,N_24564);
nand U25030 (N_25030,N_24833,N_24863);
xor U25031 (N_25031,N_24748,N_24688);
nand U25032 (N_25032,N_24562,N_24515);
or U25033 (N_25033,N_24650,N_24584);
or U25034 (N_25034,N_24814,N_24970);
nor U25035 (N_25035,N_24912,N_24891);
and U25036 (N_25036,N_24546,N_24782);
or U25037 (N_25037,N_24968,N_24604);
and U25038 (N_25038,N_24791,N_24850);
nor U25039 (N_25039,N_24852,N_24956);
xnor U25040 (N_25040,N_24609,N_24582);
or U25041 (N_25041,N_24930,N_24790);
nor U25042 (N_25042,N_24605,N_24544);
nor U25043 (N_25043,N_24858,N_24591);
nand U25044 (N_25044,N_24741,N_24634);
nor U25045 (N_25045,N_24835,N_24671);
and U25046 (N_25046,N_24861,N_24769);
xor U25047 (N_25047,N_24916,N_24503);
nand U25048 (N_25048,N_24834,N_24992);
or U25049 (N_25049,N_24828,N_24837);
and U25050 (N_25050,N_24635,N_24502);
or U25051 (N_25051,N_24954,N_24877);
xnor U25052 (N_25052,N_24991,N_24935);
or U25053 (N_25053,N_24686,N_24856);
nand U25054 (N_25054,N_24938,N_24917);
or U25055 (N_25055,N_24627,N_24829);
nor U25056 (N_25056,N_24642,N_24888);
nor U25057 (N_25057,N_24571,N_24862);
xnor U25058 (N_25058,N_24818,N_24613);
xnor U25059 (N_25059,N_24631,N_24668);
nor U25060 (N_25060,N_24848,N_24788);
and U25061 (N_25061,N_24590,N_24778);
and U25062 (N_25062,N_24719,N_24966);
nor U25063 (N_25063,N_24923,N_24774);
xor U25064 (N_25064,N_24972,N_24745);
nor U25065 (N_25065,N_24595,N_24577);
nor U25066 (N_25066,N_24853,N_24821);
and U25067 (N_25067,N_24816,N_24674);
xnor U25068 (N_25068,N_24527,N_24949);
xor U25069 (N_25069,N_24670,N_24880);
or U25070 (N_25070,N_24569,N_24644);
nor U25071 (N_25071,N_24952,N_24867);
xnor U25072 (N_25072,N_24602,N_24770);
nand U25073 (N_25073,N_24755,N_24507);
nor U25074 (N_25074,N_24708,N_24932);
or U25075 (N_25075,N_24753,N_24509);
nor U25076 (N_25076,N_24695,N_24565);
xor U25077 (N_25077,N_24504,N_24890);
and U25078 (N_25078,N_24730,N_24693);
nor U25079 (N_25079,N_24760,N_24596);
nand U25080 (N_25080,N_24716,N_24606);
nor U25081 (N_25081,N_24698,N_24756);
or U25082 (N_25082,N_24720,N_24802);
nand U25083 (N_25083,N_24902,N_24908);
nor U25084 (N_25084,N_24614,N_24554);
nand U25085 (N_25085,N_24603,N_24920);
or U25086 (N_25086,N_24971,N_24979);
xnor U25087 (N_25087,N_24725,N_24667);
nand U25088 (N_25088,N_24758,N_24946);
nand U25089 (N_25089,N_24586,N_24661);
nor U25090 (N_25090,N_24714,N_24784);
nand U25091 (N_25091,N_24903,N_24857);
xor U25092 (N_25092,N_24898,N_24665);
nand U25093 (N_25093,N_24709,N_24640);
nor U25094 (N_25094,N_24995,N_24553);
or U25095 (N_25095,N_24563,N_24983);
nor U25096 (N_25096,N_24924,N_24780);
nand U25097 (N_25097,N_24628,N_24933);
or U25098 (N_25098,N_24851,N_24925);
xor U25099 (N_25099,N_24636,N_24712);
xor U25100 (N_25100,N_24506,N_24558);
nor U25101 (N_25101,N_24623,N_24587);
and U25102 (N_25102,N_24608,N_24705);
xor U25103 (N_25103,N_24690,N_24704);
xnor U25104 (N_25104,N_24570,N_24803);
or U25105 (N_25105,N_24842,N_24579);
nor U25106 (N_25106,N_24568,N_24574);
xor U25107 (N_25107,N_24677,N_24822);
xnor U25108 (N_25108,N_24588,N_24798);
nand U25109 (N_25109,N_24715,N_24887);
nand U25110 (N_25110,N_24860,N_24965);
xnor U25111 (N_25111,N_24820,N_24696);
or U25112 (N_25112,N_24697,N_24618);
and U25113 (N_25113,N_24776,N_24922);
xor U25114 (N_25114,N_24687,N_24999);
nand U25115 (N_25115,N_24551,N_24950);
or U25116 (N_25116,N_24626,N_24975);
nand U25117 (N_25117,N_24530,N_24919);
nor U25118 (N_25118,N_24654,N_24976);
nand U25119 (N_25119,N_24539,N_24957);
nor U25120 (N_25120,N_24542,N_24994);
or U25121 (N_25121,N_24703,N_24918);
nand U25122 (N_25122,N_24731,N_24726);
and U25123 (N_25123,N_24663,N_24682);
nand U25124 (N_25124,N_24771,N_24520);
or U25125 (N_25125,N_24944,N_24985);
nand U25126 (N_25126,N_24727,N_24875);
or U25127 (N_25127,N_24617,N_24859);
or U25128 (N_25128,N_24967,N_24589);
nor U25129 (N_25129,N_24762,N_24940);
xor U25130 (N_25130,N_24532,N_24679);
xor U25131 (N_25131,N_24910,N_24980);
nand U25132 (N_25132,N_24787,N_24724);
nand U25133 (N_25133,N_24534,N_24914);
xnor U25134 (N_25134,N_24525,N_24786);
nor U25135 (N_25135,N_24978,N_24797);
and U25136 (N_25136,N_24945,N_24846);
nor U25137 (N_25137,N_24879,N_24669);
nor U25138 (N_25138,N_24865,N_24713);
and U25139 (N_25139,N_24528,N_24807);
nand U25140 (N_25140,N_24961,N_24678);
xor U25141 (N_25141,N_24573,N_24557);
or U25142 (N_25142,N_24556,N_24612);
xnor U25143 (N_25143,N_24773,N_24585);
and U25144 (N_25144,N_24658,N_24899);
nand U25145 (N_25145,N_24630,N_24611);
xor U25146 (N_25146,N_24621,N_24744);
or U25147 (N_25147,N_24815,N_24597);
nand U25148 (N_25148,N_24524,N_24907);
nand U25149 (N_25149,N_24750,N_24518);
xnor U25150 (N_25150,N_24826,N_24793);
nand U25151 (N_25151,N_24894,N_24873);
or U25152 (N_25152,N_24735,N_24733);
xnor U25153 (N_25153,N_24960,N_24531);
nor U25154 (N_25154,N_24984,N_24548);
nor U25155 (N_25155,N_24600,N_24694);
nand U25156 (N_25156,N_24819,N_24915);
nand U25157 (N_25157,N_24529,N_24652);
and U25158 (N_25158,N_24900,N_24882);
xor U25159 (N_25159,N_24812,N_24931);
or U25160 (N_25160,N_24988,N_24691);
nand U25161 (N_25161,N_24974,N_24870);
or U25162 (N_25162,N_24700,N_24517);
nand U25163 (N_25163,N_24619,N_24702);
nand U25164 (N_25164,N_24683,N_24536);
xor U25165 (N_25165,N_24883,N_24876);
xor U25166 (N_25166,N_24512,N_24721);
xnor U25167 (N_25167,N_24996,N_24871);
nand U25168 (N_25168,N_24729,N_24936);
nor U25169 (N_25169,N_24808,N_24576);
and U25170 (N_25170,N_24625,N_24673);
xnor U25171 (N_25171,N_24959,N_24655);
nand U25172 (N_25172,N_24643,N_24566);
nand U25173 (N_25173,N_24739,N_24718);
or U25174 (N_25174,N_24869,N_24657);
or U25175 (N_25175,N_24624,N_24537);
nor U25176 (N_25176,N_24926,N_24982);
nand U25177 (N_25177,N_24904,N_24541);
or U25178 (N_25178,N_24656,N_24977);
xor U25179 (N_25179,N_24723,N_24897);
nor U25180 (N_25180,N_24706,N_24672);
nand U25181 (N_25181,N_24552,N_24511);
nand U25182 (N_25182,N_24805,N_24840);
or U25183 (N_25183,N_24500,N_24759);
xnor U25184 (N_25184,N_24754,N_24761);
and U25185 (N_25185,N_24601,N_24549);
and U25186 (N_25186,N_24779,N_24806);
or U25187 (N_25187,N_24543,N_24620);
xor U25188 (N_25188,N_24799,N_24955);
and U25189 (N_25189,N_24538,N_24743);
nor U25190 (N_25190,N_24707,N_24660);
or U25191 (N_25191,N_24580,N_24847);
xnor U25192 (N_25192,N_24885,N_24804);
and U25193 (N_25193,N_24993,N_24749);
xnor U25194 (N_25194,N_24639,N_24969);
nand U25195 (N_25195,N_24717,N_24738);
xnor U25196 (N_25196,N_24800,N_24909);
nand U25197 (N_25197,N_24747,N_24824);
nand U25198 (N_25198,N_24689,N_24522);
and U25199 (N_25199,N_24559,N_24521);
nand U25200 (N_25200,N_24555,N_24701);
xor U25201 (N_25201,N_24839,N_24872);
and U25202 (N_25202,N_24575,N_24526);
xor U25203 (N_25203,N_24746,N_24728);
or U25204 (N_25204,N_24645,N_24662);
nor U25205 (N_25205,N_24647,N_24675);
or U25206 (N_25206,N_24767,N_24864);
xor U25207 (N_25207,N_24893,N_24886);
and U25208 (N_25208,N_24986,N_24892);
nand U25209 (N_25209,N_24622,N_24722);
and U25210 (N_25210,N_24906,N_24567);
nor U25211 (N_25211,N_24895,N_24583);
or U25212 (N_25212,N_24866,N_24685);
or U25213 (N_25213,N_24981,N_24884);
or U25214 (N_25214,N_24998,N_24929);
and U25215 (N_25215,N_24615,N_24681);
nor U25216 (N_25216,N_24947,N_24937);
and U25217 (N_25217,N_24941,N_24849);
xnor U25218 (N_25218,N_24913,N_24616);
or U25219 (N_25219,N_24523,N_24783);
xnor U25220 (N_25220,N_24958,N_24648);
nor U25221 (N_25221,N_24845,N_24629);
and U25222 (N_25222,N_24928,N_24868);
or U25223 (N_25223,N_24953,N_24632);
xor U25224 (N_25224,N_24987,N_24823);
nor U25225 (N_25225,N_24676,N_24736);
nand U25226 (N_25226,N_24734,N_24572);
or U25227 (N_25227,N_24809,N_24796);
and U25228 (N_25228,N_24692,N_24519);
nor U25229 (N_25229,N_24843,N_24508);
nand U25230 (N_25230,N_24680,N_24545);
nor U25231 (N_25231,N_24768,N_24775);
nand U25232 (N_25232,N_24513,N_24990);
and U25233 (N_25233,N_24766,N_24594);
xor U25234 (N_25234,N_24964,N_24831);
xnor U25235 (N_25235,N_24633,N_24830);
nor U25236 (N_25236,N_24607,N_24825);
and U25237 (N_25237,N_24533,N_24592);
nor U25238 (N_25238,N_24547,N_24881);
nand U25239 (N_25239,N_24810,N_24732);
nor U25240 (N_25240,N_24699,N_24838);
nand U25241 (N_25241,N_24989,N_24742);
nand U25242 (N_25242,N_24505,N_24501);
and U25243 (N_25243,N_24951,N_24561);
xor U25244 (N_25244,N_24874,N_24751);
nand U25245 (N_25245,N_24905,N_24765);
and U25246 (N_25246,N_24540,N_24795);
nand U25247 (N_25247,N_24896,N_24653);
nor U25248 (N_25248,N_24560,N_24535);
nor U25249 (N_25249,N_24792,N_24943);
xnor U25250 (N_25250,N_24712,N_24771);
nand U25251 (N_25251,N_24512,N_24929);
or U25252 (N_25252,N_24587,N_24771);
nand U25253 (N_25253,N_24598,N_24547);
nor U25254 (N_25254,N_24979,N_24985);
or U25255 (N_25255,N_24749,N_24916);
nand U25256 (N_25256,N_24896,N_24684);
and U25257 (N_25257,N_24600,N_24949);
or U25258 (N_25258,N_24724,N_24923);
nor U25259 (N_25259,N_24518,N_24659);
xnor U25260 (N_25260,N_24969,N_24771);
and U25261 (N_25261,N_24855,N_24759);
or U25262 (N_25262,N_24956,N_24994);
xor U25263 (N_25263,N_24858,N_24860);
xnor U25264 (N_25264,N_24740,N_24945);
or U25265 (N_25265,N_24569,N_24793);
and U25266 (N_25266,N_24679,N_24787);
and U25267 (N_25267,N_24780,N_24839);
nor U25268 (N_25268,N_24697,N_24507);
or U25269 (N_25269,N_24784,N_24908);
xnor U25270 (N_25270,N_24861,N_24566);
nand U25271 (N_25271,N_24803,N_24643);
nand U25272 (N_25272,N_24672,N_24560);
nor U25273 (N_25273,N_24543,N_24790);
xnor U25274 (N_25274,N_24961,N_24687);
xor U25275 (N_25275,N_24554,N_24563);
and U25276 (N_25276,N_24951,N_24732);
xnor U25277 (N_25277,N_24716,N_24709);
nand U25278 (N_25278,N_24739,N_24618);
nor U25279 (N_25279,N_24691,N_24985);
nor U25280 (N_25280,N_24943,N_24732);
nand U25281 (N_25281,N_24608,N_24855);
xor U25282 (N_25282,N_24988,N_24741);
xnor U25283 (N_25283,N_24629,N_24614);
and U25284 (N_25284,N_24944,N_24513);
nand U25285 (N_25285,N_24671,N_24961);
or U25286 (N_25286,N_24694,N_24603);
nand U25287 (N_25287,N_24988,N_24737);
xnor U25288 (N_25288,N_24938,N_24845);
nand U25289 (N_25289,N_24724,N_24846);
xnor U25290 (N_25290,N_24726,N_24808);
nor U25291 (N_25291,N_24661,N_24916);
and U25292 (N_25292,N_24728,N_24639);
nand U25293 (N_25293,N_24973,N_24757);
and U25294 (N_25294,N_24637,N_24993);
nand U25295 (N_25295,N_24684,N_24792);
or U25296 (N_25296,N_24888,N_24977);
xnor U25297 (N_25297,N_24683,N_24965);
nor U25298 (N_25298,N_24552,N_24624);
or U25299 (N_25299,N_24821,N_24565);
or U25300 (N_25300,N_24696,N_24985);
or U25301 (N_25301,N_24568,N_24632);
or U25302 (N_25302,N_24780,N_24980);
nand U25303 (N_25303,N_24790,N_24617);
xnor U25304 (N_25304,N_24894,N_24906);
nor U25305 (N_25305,N_24589,N_24937);
nor U25306 (N_25306,N_24685,N_24840);
xor U25307 (N_25307,N_24639,N_24925);
and U25308 (N_25308,N_24759,N_24832);
or U25309 (N_25309,N_24973,N_24921);
nand U25310 (N_25310,N_24808,N_24577);
xnor U25311 (N_25311,N_24715,N_24773);
nand U25312 (N_25312,N_24938,N_24591);
nand U25313 (N_25313,N_24531,N_24602);
or U25314 (N_25314,N_24567,N_24633);
xor U25315 (N_25315,N_24600,N_24718);
nor U25316 (N_25316,N_24863,N_24877);
or U25317 (N_25317,N_24699,N_24757);
or U25318 (N_25318,N_24719,N_24931);
or U25319 (N_25319,N_24829,N_24556);
xnor U25320 (N_25320,N_24584,N_24992);
and U25321 (N_25321,N_24501,N_24622);
and U25322 (N_25322,N_24703,N_24951);
and U25323 (N_25323,N_24684,N_24543);
nor U25324 (N_25324,N_24978,N_24633);
or U25325 (N_25325,N_24675,N_24592);
and U25326 (N_25326,N_24757,N_24749);
and U25327 (N_25327,N_24707,N_24528);
nor U25328 (N_25328,N_24571,N_24930);
or U25329 (N_25329,N_24835,N_24657);
and U25330 (N_25330,N_24912,N_24585);
xor U25331 (N_25331,N_24898,N_24812);
and U25332 (N_25332,N_24912,N_24999);
nor U25333 (N_25333,N_24693,N_24574);
nor U25334 (N_25334,N_24566,N_24876);
or U25335 (N_25335,N_24766,N_24829);
nand U25336 (N_25336,N_24974,N_24964);
nand U25337 (N_25337,N_24631,N_24812);
or U25338 (N_25338,N_24594,N_24724);
and U25339 (N_25339,N_24875,N_24558);
nor U25340 (N_25340,N_24776,N_24818);
and U25341 (N_25341,N_24915,N_24646);
or U25342 (N_25342,N_24984,N_24814);
nand U25343 (N_25343,N_24827,N_24627);
nor U25344 (N_25344,N_24823,N_24902);
xor U25345 (N_25345,N_24735,N_24852);
nand U25346 (N_25346,N_24863,N_24577);
and U25347 (N_25347,N_24636,N_24566);
and U25348 (N_25348,N_24635,N_24990);
nor U25349 (N_25349,N_24939,N_24644);
or U25350 (N_25350,N_24673,N_24516);
and U25351 (N_25351,N_24704,N_24803);
or U25352 (N_25352,N_24947,N_24653);
nor U25353 (N_25353,N_24790,N_24674);
and U25354 (N_25354,N_24628,N_24859);
or U25355 (N_25355,N_24914,N_24697);
or U25356 (N_25356,N_24931,N_24583);
or U25357 (N_25357,N_24901,N_24786);
and U25358 (N_25358,N_24853,N_24900);
xor U25359 (N_25359,N_24656,N_24690);
nor U25360 (N_25360,N_24545,N_24776);
nand U25361 (N_25361,N_24928,N_24647);
or U25362 (N_25362,N_24957,N_24762);
xor U25363 (N_25363,N_24951,N_24664);
and U25364 (N_25364,N_24812,N_24838);
xor U25365 (N_25365,N_24996,N_24536);
nand U25366 (N_25366,N_24697,N_24741);
or U25367 (N_25367,N_24782,N_24935);
nor U25368 (N_25368,N_24830,N_24723);
and U25369 (N_25369,N_24602,N_24836);
nand U25370 (N_25370,N_24604,N_24513);
or U25371 (N_25371,N_24521,N_24869);
xnor U25372 (N_25372,N_24816,N_24632);
and U25373 (N_25373,N_24850,N_24690);
or U25374 (N_25374,N_24614,N_24838);
and U25375 (N_25375,N_24549,N_24825);
or U25376 (N_25376,N_24948,N_24515);
and U25377 (N_25377,N_24920,N_24904);
nand U25378 (N_25378,N_24602,N_24659);
nor U25379 (N_25379,N_24957,N_24532);
or U25380 (N_25380,N_24565,N_24936);
xnor U25381 (N_25381,N_24845,N_24777);
and U25382 (N_25382,N_24563,N_24743);
or U25383 (N_25383,N_24940,N_24721);
xor U25384 (N_25384,N_24714,N_24800);
nor U25385 (N_25385,N_24827,N_24990);
nor U25386 (N_25386,N_24503,N_24692);
and U25387 (N_25387,N_24627,N_24571);
nor U25388 (N_25388,N_24518,N_24810);
or U25389 (N_25389,N_24853,N_24588);
and U25390 (N_25390,N_24617,N_24566);
or U25391 (N_25391,N_24658,N_24674);
nor U25392 (N_25392,N_24651,N_24603);
nor U25393 (N_25393,N_24724,N_24582);
nand U25394 (N_25394,N_24632,N_24866);
nor U25395 (N_25395,N_24630,N_24679);
nand U25396 (N_25396,N_24577,N_24909);
nand U25397 (N_25397,N_24957,N_24603);
and U25398 (N_25398,N_24615,N_24894);
or U25399 (N_25399,N_24666,N_24816);
or U25400 (N_25400,N_24622,N_24779);
and U25401 (N_25401,N_24552,N_24892);
nor U25402 (N_25402,N_24904,N_24663);
and U25403 (N_25403,N_24772,N_24750);
nand U25404 (N_25404,N_24895,N_24555);
nor U25405 (N_25405,N_24709,N_24767);
or U25406 (N_25406,N_24667,N_24669);
nor U25407 (N_25407,N_24655,N_24537);
nand U25408 (N_25408,N_24769,N_24567);
and U25409 (N_25409,N_24906,N_24708);
and U25410 (N_25410,N_24744,N_24507);
nand U25411 (N_25411,N_24520,N_24841);
nor U25412 (N_25412,N_24775,N_24647);
xor U25413 (N_25413,N_24738,N_24808);
and U25414 (N_25414,N_24806,N_24594);
or U25415 (N_25415,N_24528,N_24505);
nor U25416 (N_25416,N_24706,N_24941);
or U25417 (N_25417,N_24656,N_24935);
nor U25418 (N_25418,N_24967,N_24772);
or U25419 (N_25419,N_24829,N_24896);
nor U25420 (N_25420,N_24953,N_24684);
nand U25421 (N_25421,N_24980,N_24640);
and U25422 (N_25422,N_24838,N_24502);
nand U25423 (N_25423,N_24789,N_24646);
nor U25424 (N_25424,N_24542,N_24633);
nor U25425 (N_25425,N_24716,N_24519);
or U25426 (N_25426,N_24552,N_24633);
and U25427 (N_25427,N_24961,N_24852);
and U25428 (N_25428,N_24992,N_24526);
xnor U25429 (N_25429,N_24551,N_24673);
nor U25430 (N_25430,N_24951,N_24937);
xor U25431 (N_25431,N_24806,N_24653);
nor U25432 (N_25432,N_24901,N_24817);
and U25433 (N_25433,N_24937,N_24527);
xor U25434 (N_25434,N_24534,N_24564);
xor U25435 (N_25435,N_24835,N_24676);
nand U25436 (N_25436,N_24768,N_24725);
nand U25437 (N_25437,N_24910,N_24671);
nand U25438 (N_25438,N_24982,N_24541);
xnor U25439 (N_25439,N_24894,N_24971);
and U25440 (N_25440,N_24737,N_24584);
xor U25441 (N_25441,N_24964,N_24798);
and U25442 (N_25442,N_24978,N_24752);
or U25443 (N_25443,N_24668,N_24752);
and U25444 (N_25444,N_24814,N_24993);
nor U25445 (N_25445,N_24939,N_24514);
nor U25446 (N_25446,N_24968,N_24937);
and U25447 (N_25447,N_24962,N_24849);
or U25448 (N_25448,N_24753,N_24580);
xnor U25449 (N_25449,N_24831,N_24921);
nor U25450 (N_25450,N_24732,N_24851);
xor U25451 (N_25451,N_24936,N_24533);
and U25452 (N_25452,N_24624,N_24770);
and U25453 (N_25453,N_24633,N_24787);
and U25454 (N_25454,N_24593,N_24530);
xor U25455 (N_25455,N_24601,N_24578);
xnor U25456 (N_25456,N_24888,N_24884);
nand U25457 (N_25457,N_24791,N_24619);
and U25458 (N_25458,N_24865,N_24981);
nand U25459 (N_25459,N_24692,N_24853);
and U25460 (N_25460,N_24910,N_24543);
xor U25461 (N_25461,N_24758,N_24799);
or U25462 (N_25462,N_24851,N_24961);
or U25463 (N_25463,N_24786,N_24642);
nand U25464 (N_25464,N_24585,N_24979);
or U25465 (N_25465,N_24880,N_24590);
or U25466 (N_25466,N_24981,N_24926);
nor U25467 (N_25467,N_24932,N_24623);
nor U25468 (N_25468,N_24937,N_24995);
nor U25469 (N_25469,N_24955,N_24780);
nand U25470 (N_25470,N_24585,N_24879);
nor U25471 (N_25471,N_24832,N_24704);
or U25472 (N_25472,N_24722,N_24846);
xnor U25473 (N_25473,N_24694,N_24662);
or U25474 (N_25474,N_24885,N_24788);
nor U25475 (N_25475,N_24805,N_24533);
xor U25476 (N_25476,N_24925,N_24759);
or U25477 (N_25477,N_24945,N_24589);
nand U25478 (N_25478,N_24714,N_24876);
xnor U25479 (N_25479,N_24764,N_24598);
nand U25480 (N_25480,N_24723,N_24764);
nor U25481 (N_25481,N_24642,N_24747);
nand U25482 (N_25482,N_24844,N_24914);
and U25483 (N_25483,N_24687,N_24977);
xor U25484 (N_25484,N_24779,N_24740);
nand U25485 (N_25485,N_24898,N_24575);
nor U25486 (N_25486,N_24724,N_24716);
nor U25487 (N_25487,N_24923,N_24546);
and U25488 (N_25488,N_24785,N_24661);
nand U25489 (N_25489,N_24687,N_24805);
nor U25490 (N_25490,N_24703,N_24595);
or U25491 (N_25491,N_24935,N_24831);
nor U25492 (N_25492,N_24863,N_24641);
nor U25493 (N_25493,N_24735,N_24611);
xor U25494 (N_25494,N_24696,N_24617);
nor U25495 (N_25495,N_24504,N_24894);
xor U25496 (N_25496,N_24795,N_24766);
nor U25497 (N_25497,N_24562,N_24696);
or U25498 (N_25498,N_24806,N_24532);
nand U25499 (N_25499,N_24625,N_24588);
xnor U25500 (N_25500,N_25030,N_25122);
xor U25501 (N_25501,N_25357,N_25338);
nor U25502 (N_25502,N_25285,N_25067);
nand U25503 (N_25503,N_25039,N_25135);
nand U25504 (N_25504,N_25430,N_25372);
nor U25505 (N_25505,N_25295,N_25180);
xor U25506 (N_25506,N_25016,N_25167);
and U25507 (N_25507,N_25490,N_25223);
and U25508 (N_25508,N_25044,N_25025);
nor U25509 (N_25509,N_25464,N_25255);
nor U25510 (N_25510,N_25446,N_25365);
nor U25511 (N_25511,N_25475,N_25179);
xor U25512 (N_25512,N_25029,N_25071);
xnor U25513 (N_25513,N_25184,N_25352);
nor U25514 (N_25514,N_25283,N_25075);
nor U25515 (N_25515,N_25217,N_25459);
and U25516 (N_25516,N_25380,N_25163);
or U25517 (N_25517,N_25387,N_25381);
xor U25518 (N_25518,N_25341,N_25236);
nand U25519 (N_25519,N_25378,N_25031);
xor U25520 (N_25520,N_25328,N_25248);
or U25521 (N_25521,N_25336,N_25262);
nand U25522 (N_25522,N_25403,N_25073);
xnor U25523 (N_25523,N_25054,N_25226);
xnor U25524 (N_25524,N_25414,N_25144);
nor U25525 (N_25525,N_25488,N_25245);
nor U25526 (N_25526,N_25186,N_25363);
and U25527 (N_25527,N_25438,N_25118);
or U25528 (N_25528,N_25251,N_25420);
and U25529 (N_25529,N_25242,N_25492);
nand U25530 (N_25530,N_25162,N_25158);
and U25531 (N_25531,N_25389,N_25423);
nor U25532 (N_25532,N_25287,N_25280);
or U25533 (N_25533,N_25219,N_25308);
nand U25534 (N_25534,N_25270,N_25155);
xnor U25535 (N_25535,N_25457,N_25436);
nor U25536 (N_25536,N_25193,N_25001);
nand U25537 (N_25537,N_25188,N_25078);
and U25538 (N_25538,N_25337,N_25126);
and U25539 (N_25539,N_25116,N_25413);
or U25540 (N_25540,N_25474,N_25173);
or U25541 (N_25541,N_25063,N_25159);
xnor U25542 (N_25542,N_25222,N_25291);
nand U25543 (N_25543,N_25407,N_25410);
nand U25544 (N_25544,N_25312,N_25318);
and U25545 (N_25545,N_25320,N_25297);
nor U25546 (N_25546,N_25383,N_25115);
or U25547 (N_25547,N_25244,N_25136);
or U25548 (N_25548,N_25290,N_25334);
or U25549 (N_25549,N_25323,N_25092);
nor U25550 (N_25550,N_25349,N_25482);
nand U25551 (N_25551,N_25429,N_25125);
and U25552 (N_25552,N_25398,N_25002);
or U25553 (N_25553,N_25360,N_25012);
xor U25554 (N_25554,N_25061,N_25281);
or U25555 (N_25555,N_25463,N_25424);
or U25556 (N_25556,N_25443,N_25294);
nor U25557 (N_25557,N_25160,N_25182);
or U25558 (N_25558,N_25271,N_25028);
and U25559 (N_25559,N_25119,N_25469);
nand U25560 (N_25560,N_25239,N_25348);
and U25561 (N_25561,N_25487,N_25289);
nand U25562 (N_25562,N_25204,N_25279);
or U25563 (N_25563,N_25485,N_25276);
xnor U25564 (N_25564,N_25342,N_25174);
and U25565 (N_25565,N_25235,N_25010);
nand U25566 (N_25566,N_25267,N_25168);
xor U25567 (N_25567,N_25339,N_25109);
nand U25568 (N_25568,N_25120,N_25497);
and U25569 (N_25569,N_25057,N_25089);
xor U25570 (N_25570,N_25307,N_25178);
or U25571 (N_25571,N_25298,N_25422);
nand U25572 (N_25572,N_25189,N_25134);
and U25573 (N_25573,N_25011,N_25264);
and U25574 (N_25574,N_25077,N_25364);
nor U25575 (N_25575,N_25213,N_25055);
or U25576 (N_25576,N_25456,N_25220);
nor U25577 (N_25577,N_25099,N_25278);
nor U25578 (N_25578,N_25129,N_25008);
nand U25579 (N_25579,N_25228,N_25444);
nor U25580 (N_25580,N_25201,N_25088);
xor U25581 (N_25581,N_25056,N_25140);
or U25582 (N_25582,N_25361,N_25254);
nand U25583 (N_25583,N_25166,N_25038);
nand U25584 (N_25584,N_25081,N_25000);
xor U25585 (N_25585,N_25395,N_25154);
and U25586 (N_25586,N_25074,N_25151);
or U25587 (N_25587,N_25326,N_25448);
and U25588 (N_25588,N_25198,N_25232);
nor U25589 (N_25589,N_25227,N_25241);
nor U25590 (N_25590,N_25246,N_25354);
and U25591 (N_25591,N_25453,N_25440);
or U25592 (N_25592,N_25368,N_25455);
nor U25593 (N_25593,N_25494,N_25371);
nor U25594 (N_25594,N_25468,N_25411);
nor U25595 (N_25595,N_25147,N_25133);
nor U25596 (N_25596,N_25311,N_25209);
or U25597 (N_25597,N_25268,N_25142);
xor U25598 (N_25598,N_25121,N_25392);
xor U25599 (N_25599,N_25181,N_25141);
xor U25600 (N_25600,N_25176,N_25417);
and U25601 (N_25601,N_25305,N_25489);
or U25602 (N_25602,N_25356,N_25317);
or U25603 (N_25603,N_25149,N_25024);
or U25604 (N_25604,N_25385,N_25304);
nor U25605 (N_25605,N_25231,N_25384);
or U25606 (N_25606,N_25401,N_25259);
and U25607 (N_25607,N_25237,N_25185);
and U25608 (N_25608,N_25022,N_25406);
nor U25609 (N_25609,N_25230,N_25053);
or U25610 (N_25610,N_25316,N_25172);
or U25611 (N_25611,N_25019,N_25052);
xor U25612 (N_25612,N_25351,N_25415);
xor U25613 (N_25613,N_25156,N_25132);
xnor U25614 (N_25614,N_25036,N_25388);
nor U25615 (N_25615,N_25393,N_25284);
xor U25616 (N_25616,N_25037,N_25458);
nand U25617 (N_25617,N_25353,N_25493);
nor U25618 (N_25618,N_25131,N_25322);
and U25619 (N_25619,N_25369,N_25009);
nor U25620 (N_25620,N_25343,N_25203);
xor U25621 (N_25621,N_25145,N_25476);
nor U25622 (N_25622,N_25293,N_25451);
nor U25623 (N_25623,N_25441,N_25080);
xor U25624 (N_25624,N_25138,N_25359);
xor U25625 (N_25625,N_25299,N_25419);
nor U25626 (N_25626,N_25064,N_25153);
nor U25627 (N_25627,N_25402,N_25470);
nor U25628 (N_25628,N_25397,N_25199);
nand U25629 (N_25629,N_25362,N_25005);
nor U25630 (N_25630,N_25471,N_25187);
or U25631 (N_25631,N_25041,N_25164);
or U25632 (N_25632,N_25137,N_25086);
or U25633 (N_25633,N_25247,N_25333);
xor U25634 (N_25634,N_25252,N_25048);
nor U25635 (N_25635,N_25068,N_25421);
or U25636 (N_25636,N_25026,N_25047);
or U25637 (N_25637,N_25192,N_25197);
nand U25638 (N_25638,N_25321,N_25331);
and U25639 (N_25639,N_25060,N_25175);
xor U25640 (N_25640,N_25288,N_25096);
xnor U25641 (N_25641,N_25069,N_25218);
or U25642 (N_25642,N_25114,N_25366);
nor U25643 (N_25643,N_25396,N_25152);
or U25644 (N_25644,N_25108,N_25094);
and U25645 (N_25645,N_25085,N_25146);
nand U25646 (N_25646,N_25447,N_25426);
or U25647 (N_25647,N_25206,N_25325);
and U25648 (N_25648,N_25486,N_25275);
or U25649 (N_25649,N_25087,N_25100);
nand U25650 (N_25650,N_25496,N_25258);
or U25651 (N_25651,N_25079,N_25309);
and U25652 (N_25652,N_25499,N_25327);
nor U25653 (N_25653,N_25059,N_25212);
and U25654 (N_25654,N_25382,N_25434);
nand U25655 (N_25655,N_25106,N_25452);
nand U25656 (N_25656,N_25329,N_25310);
nand U25657 (N_25657,N_25404,N_25435);
and U25658 (N_25658,N_25082,N_25263);
nand U25659 (N_25659,N_25340,N_25277);
or U25660 (N_25660,N_25240,N_25183);
nor U25661 (N_25661,N_25195,N_25211);
and U25662 (N_25662,N_25437,N_25257);
or U25663 (N_25663,N_25070,N_25405);
xor U25664 (N_25664,N_25233,N_25105);
nor U25665 (N_25665,N_25479,N_25472);
and U25666 (N_25666,N_25045,N_25139);
or U25667 (N_25667,N_25004,N_25427);
and U25668 (N_25668,N_25196,N_25098);
and U25669 (N_25669,N_25449,N_25358);
nor U25670 (N_25670,N_25101,N_25225);
xor U25671 (N_25671,N_25300,N_25097);
nor U25672 (N_25672,N_25083,N_25350);
nand U25673 (N_25673,N_25386,N_25051);
or U25674 (N_25674,N_25202,N_25095);
nand U25675 (N_25675,N_25110,N_25208);
xor U25676 (N_25676,N_25399,N_25177);
nor U25677 (N_25677,N_25130,N_25046);
nand U25678 (N_25678,N_25161,N_25104);
nor U25679 (N_25679,N_25260,N_25150);
and U25680 (N_25680,N_25439,N_25273);
nand U25681 (N_25681,N_25454,N_25091);
and U25682 (N_25682,N_25123,N_25390);
nand U25683 (N_25683,N_25391,N_25170);
or U25684 (N_25684,N_25296,N_25332);
and U25685 (N_25685,N_25207,N_25450);
nand U25686 (N_25686,N_25473,N_25127);
and U25687 (N_25687,N_25076,N_25214);
and U25688 (N_25688,N_25072,N_25165);
and U25689 (N_25689,N_25377,N_25253);
nor U25690 (N_25690,N_25425,N_25302);
and U25691 (N_25691,N_25465,N_25286);
and U25692 (N_25692,N_25376,N_25111);
nand U25693 (N_25693,N_25256,N_25042);
and U25694 (N_25694,N_25043,N_25157);
xnor U25695 (N_25695,N_25148,N_25379);
xnor U25696 (N_25696,N_25117,N_25269);
nand U25697 (N_25697,N_25065,N_25018);
nor U25698 (N_25698,N_25058,N_25200);
nor U25699 (N_25699,N_25478,N_25229);
nor U25700 (N_25700,N_25023,N_25347);
xnor U25701 (N_25701,N_25190,N_25171);
and U25702 (N_25702,N_25027,N_25261);
nor U25703 (N_25703,N_25274,N_25221);
or U25704 (N_25704,N_25034,N_25272);
and U25705 (N_25705,N_25224,N_25084);
nor U25706 (N_25706,N_25370,N_25491);
xor U25707 (N_25707,N_25481,N_25428);
nor U25708 (N_25708,N_25234,N_25346);
xnor U25709 (N_25709,N_25335,N_25480);
nand U25710 (N_25710,N_25373,N_25355);
and U25711 (N_25711,N_25282,N_25466);
xor U25712 (N_25712,N_25292,N_25400);
and U25713 (N_25713,N_25049,N_25409);
or U25714 (N_25714,N_25477,N_25112);
or U25715 (N_25715,N_25032,N_25113);
xor U25716 (N_25716,N_25301,N_25431);
and U25717 (N_25717,N_25216,N_25483);
and U25718 (N_25718,N_25306,N_25374);
nor U25719 (N_25719,N_25191,N_25330);
nand U25720 (N_25720,N_25445,N_25143);
or U25721 (N_25721,N_25006,N_25205);
and U25722 (N_25722,N_25003,N_25020);
nor U25723 (N_25723,N_25265,N_25238);
or U25724 (N_25724,N_25249,N_25467);
and U25725 (N_25725,N_25040,N_25014);
or U25726 (N_25726,N_25314,N_25093);
nor U25727 (N_25727,N_25484,N_25433);
nand U25728 (N_25728,N_25035,N_25215);
nor U25729 (N_25729,N_25017,N_25062);
or U25730 (N_25730,N_25210,N_25021);
or U25731 (N_25731,N_25460,N_25442);
nor U25732 (N_25732,N_25266,N_25243);
xor U25733 (N_25733,N_25416,N_25007);
and U25734 (N_25734,N_25367,N_25418);
nor U25735 (N_25735,N_25495,N_25375);
nand U25736 (N_25736,N_25344,N_25124);
nor U25737 (N_25737,N_25033,N_25462);
and U25738 (N_25738,N_25169,N_25319);
nand U25739 (N_25739,N_25313,N_25408);
and U25740 (N_25740,N_25432,N_25066);
nor U25741 (N_25741,N_25015,N_25412);
and U25742 (N_25742,N_25498,N_25250);
xor U25743 (N_25743,N_25461,N_25090);
nand U25744 (N_25744,N_25303,N_25013);
or U25745 (N_25745,N_25315,N_25128);
xnor U25746 (N_25746,N_25394,N_25103);
or U25747 (N_25747,N_25345,N_25324);
and U25748 (N_25748,N_25102,N_25050);
and U25749 (N_25749,N_25107,N_25194);
nand U25750 (N_25750,N_25068,N_25449);
or U25751 (N_25751,N_25074,N_25020);
nand U25752 (N_25752,N_25056,N_25197);
nand U25753 (N_25753,N_25384,N_25486);
nor U25754 (N_25754,N_25434,N_25404);
or U25755 (N_25755,N_25056,N_25370);
or U25756 (N_25756,N_25039,N_25030);
xnor U25757 (N_25757,N_25386,N_25002);
nor U25758 (N_25758,N_25292,N_25282);
xnor U25759 (N_25759,N_25148,N_25463);
or U25760 (N_25760,N_25118,N_25079);
nand U25761 (N_25761,N_25421,N_25426);
nor U25762 (N_25762,N_25116,N_25435);
and U25763 (N_25763,N_25493,N_25119);
or U25764 (N_25764,N_25367,N_25436);
nor U25765 (N_25765,N_25204,N_25251);
xor U25766 (N_25766,N_25482,N_25162);
xnor U25767 (N_25767,N_25443,N_25481);
xor U25768 (N_25768,N_25004,N_25233);
nand U25769 (N_25769,N_25333,N_25341);
and U25770 (N_25770,N_25043,N_25212);
and U25771 (N_25771,N_25015,N_25439);
nand U25772 (N_25772,N_25159,N_25155);
or U25773 (N_25773,N_25141,N_25454);
or U25774 (N_25774,N_25159,N_25038);
xnor U25775 (N_25775,N_25191,N_25160);
and U25776 (N_25776,N_25144,N_25071);
nand U25777 (N_25777,N_25426,N_25287);
nor U25778 (N_25778,N_25174,N_25015);
and U25779 (N_25779,N_25228,N_25482);
xnor U25780 (N_25780,N_25459,N_25106);
nor U25781 (N_25781,N_25406,N_25087);
or U25782 (N_25782,N_25141,N_25106);
nor U25783 (N_25783,N_25441,N_25182);
or U25784 (N_25784,N_25452,N_25220);
and U25785 (N_25785,N_25438,N_25038);
nand U25786 (N_25786,N_25412,N_25145);
or U25787 (N_25787,N_25462,N_25463);
nand U25788 (N_25788,N_25195,N_25225);
nand U25789 (N_25789,N_25223,N_25204);
xor U25790 (N_25790,N_25386,N_25496);
nor U25791 (N_25791,N_25206,N_25018);
or U25792 (N_25792,N_25086,N_25457);
nand U25793 (N_25793,N_25385,N_25325);
and U25794 (N_25794,N_25390,N_25446);
and U25795 (N_25795,N_25143,N_25396);
nand U25796 (N_25796,N_25193,N_25404);
or U25797 (N_25797,N_25147,N_25025);
nand U25798 (N_25798,N_25147,N_25269);
and U25799 (N_25799,N_25014,N_25192);
nand U25800 (N_25800,N_25010,N_25211);
nor U25801 (N_25801,N_25187,N_25450);
nand U25802 (N_25802,N_25330,N_25478);
or U25803 (N_25803,N_25174,N_25292);
nor U25804 (N_25804,N_25184,N_25414);
and U25805 (N_25805,N_25146,N_25256);
nand U25806 (N_25806,N_25137,N_25050);
nor U25807 (N_25807,N_25404,N_25366);
xor U25808 (N_25808,N_25240,N_25154);
and U25809 (N_25809,N_25459,N_25029);
xnor U25810 (N_25810,N_25129,N_25219);
xor U25811 (N_25811,N_25267,N_25047);
xnor U25812 (N_25812,N_25322,N_25019);
xnor U25813 (N_25813,N_25158,N_25026);
and U25814 (N_25814,N_25132,N_25210);
xor U25815 (N_25815,N_25482,N_25252);
nand U25816 (N_25816,N_25063,N_25456);
nand U25817 (N_25817,N_25242,N_25216);
and U25818 (N_25818,N_25430,N_25470);
xor U25819 (N_25819,N_25491,N_25441);
xor U25820 (N_25820,N_25116,N_25108);
xor U25821 (N_25821,N_25032,N_25109);
and U25822 (N_25822,N_25227,N_25372);
nand U25823 (N_25823,N_25083,N_25213);
xor U25824 (N_25824,N_25252,N_25221);
or U25825 (N_25825,N_25099,N_25146);
xnor U25826 (N_25826,N_25355,N_25356);
or U25827 (N_25827,N_25415,N_25311);
or U25828 (N_25828,N_25428,N_25194);
or U25829 (N_25829,N_25366,N_25215);
and U25830 (N_25830,N_25322,N_25293);
nor U25831 (N_25831,N_25358,N_25369);
and U25832 (N_25832,N_25130,N_25002);
nor U25833 (N_25833,N_25199,N_25172);
nor U25834 (N_25834,N_25095,N_25079);
and U25835 (N_25835,N_25191,N_25127);
or U25836 (N_25836,N_25185,N_25246);
nand U25837 (N_25837,N_25001,N_25377);
nand U25838 (N_25838,N_25460,N_25432);
and U25839 (N_25839,N_25467,N_25406);
or U25840 (N_25840,N_25182,N_25064);
or U25841 (N_25841,N_25422,N_25008);
and U25842 (N_25842,N_25076,N_25185);
nor U25843 (N_25843,N_25449,N_25127);
nor U25844 (N_25844,N_25383,N_25017);
or U25845 (N_25845,N_25053,N_25402);
and U25846 (N_25846,N_25026,N_25369);
nand U25847 (N_25847,N_25444,N_25274);
or U25848 (N_25848,N_25453,N_25176);
xnor U25849 (N_25849,N_25166,N_25370);
nand U25850 (N_25850,N_25125,N_25202);
nand U25851 (N_25851,N_25406,N_25439);
and U25852 (N_25852,N_25246,N_25058);
nor U25853 (N_25853,N_25179,N_25158);
or U25854 (N_25854,N_25215,N_25272);
nor U25855 (N_25855,N_25461,N_25367);
xor U25856 (N_25856,N_25103,N_25306);
and U25857 (N_25857,N_25432,N_25213);
xnor U25858 (N_25858,N_25012,N_25469);
nand U25859 (N_25859,N_25374,N_25076);
and U25860 (N_25860,N_25475,N_25314);
xor U25861 (N_25861,N_25002,N_25302);
nor U25862 (N_25862,N_25474,N_25024);
or U25863 (N_25863,N_25217,N_25035);
or U25864 (N_25864,N_25427,N_25137);
and U25865 (N_25865,N_25404,N_25176);
nand U25866 (N_25866,N_25295,N_25438);
nand U25867 (N_25867,N_25112,N_25030);
nand U25868 (N_25868,N_25024,N_25343);
nor U25869 (N_25869,N_25056,N_25297);
and U25870 (N_25870,N_25398,N_25220);
xnor U25871 (N_25871,N_25344,N_25135);
nand U25872 (N_25872,N_25120,N_25279);
xor U25873 (N_25873,N_25465,N_25387);
nor U25874 (N_25874,N_25179,N_25043);
xor U25875 (N_25875,N_25079,N_25212);
or U25876 (N_25876,N_25121,N_25204);
nor U25877 (N_25877,N_25445,N_25346);
or U25878 (N_25878,N_25230,N_25174);
nor U25879 (N_25879,N_25285,N_25125);
or U25880 (N_25880,N_25391,N_25400);
or U25881 (N_25881,N_25140,N_25153);
xnor U25882 (N_25882,N_25226,N_25153);
xnor U25883 (N_25883,N_25077,N_25263);
nor U25884 (N_25884,N_25169,N_25087);
xnor U25885 (N_25885,N_25067,N_25291);
nand U25886 (N_25886,N_25116,N_25395);
nand U25887 (N_25887,N_25099,N_25283);
nand U25888 (N_25888,N_25494,N_25335);
nor U25889 (N_25889,N_25450,N_25244);
or U25890 (N_25890,N_25257,N_25316);
nor U25891 (N_25891,N_25405,N_25498);
or U25892 (N_25892,N_25083,N_25245);
xor U25893 (N_25893,N_25016,N_25048);
xnor U25894 (N_25894,N_25171,N_25165);
and U25895 (N_25895,N_25360,N_25020);
nor U25896 (N_25896,N_25020,N_25131);
xor U25897 (N_25897,N_25390,N_25337);
nor U25898 (N_25898,N_25449,N_25407);
xnor U25899 (N_25899,N_25091,N_25441);
nor U25900 (N_25900,N_25470,N_25085);
or U25901 (N_25901,N_25383,N_25371);
nor U25902 (N_25902,N_25418,N_25147);
or U25903 (N_25903,N_25235,N_25099);
or U25904 (N_25904,N_25433,N_25282);
nand U25905 (N_25905,N_25469,N_25090);
nor U25906 (N_25906,N_25324,N_25121);
nor U25907 (N_25907,N_25491,N_25220);
nor U25908 (N_25908,N_25394,N_25499);
nor U25909 (N_25909,N_25378,N_25448);
nand U25910 (N_25910,N_25319,N_25356);
or U25911 (N_25911,N_25242,N_25062);
nand U25912 (N_25912,N_25388,N_25183);
nand U25913 (N_25913,N_25093,N_25486);
nor U25914 (N_25914,N_25361,N_25030);
nor U25915 (N_25915,N_25005,N_25000);
nand U25916 (N_25916,N_25042,N_25062);
xor U25917 (N_25917,N_25414,N_25445);
and U25918 (N_25918,N_25427,N_25227);
or U25919 (N_25919,N_25259,N_25493);
nand U25920 (N_25920,N_25004,N_25245);
and U25921 (N_25921,N_25160,N_25129);
and U25922 (N_25922,N_25324,N_25307);
and U25923 (N_25923,N_25049,N_25419);
and U25924 (N_25924,N_25361,N_25059);
nand U25925 (N_25925,N_25411,N_25497);
and U25926 (N_25926,N_25093,N_25006);
and U25927 (N_25927,N_25384,N_25392);
nand U25928 (N_25928,N_25379,N_25158);
and U25929 (N_25929,N_25066,N_25202);
and U25930 (N_25930,N_25242,N_25269);
nand U25931 (N_25931,N_25160,N_25248);
nor U25932 (N_25932,N_25050,N_25150);
or U25933 (N_25933,N_25012,N_25458);
nor U25934 (N_25934,N_25024,N_25266);
nor U25935 (N_25935,N_25463,N_25472);
and U25936 (N_25936,N_25082,N_25093);
nand U25937 (N_25937,N_25206,N_25493);
nor U25938 (N_25938,N_25262,N_25148);
and U25939 (N_25939,N_25399,N_25238);
and U25940 (N_25940,N_25236,N_25417);
or U25941 (N_25941,N_25166,N_25484);
or U25942 (N_25942,N_25102,N_25064);
or U25943 (N_25943,N_25442,N_25324);
or U25944 (N_25944,N_25381,N_25098);
xor U25945 (N_25945,N_25483,N_25176);
nor U25946 (N_25946,N_25379,N_25342);
or U25947 (N_25947,N_25296,N_25062);
xor U25948 (N_25948,N_25462,N_25207);
nand U25949 (N_25949,N_25272,N_25117);
and U25950 (N_25950,N_25043,N_25084);
or U25951 (N_25951,N_25481,N_25183);
nand U25952 (N_25952,N_25118,N_25115);
nand U25953 (N_25953,N_25112,N_25222);
nor U25954 (N_25954,N_25206,N_25335);
and U25955 (N_25955,N_25317,N_25263);
nand U25956 (N_25956,N_25485,N_25256);
nor U25957 (N_25957,N_25348,N_25454);
and U25958 (N_25958,N_25294,N_25433);
xnor U25959 (N_25959,N_25046,N_25203);
and U25960 (N_25960,N_25027,N_25421);
and U25961 (N_25961,N_25472,N_25222);
or U25962 (N_25962,N_25412,N_25259);
nand U25963 (N_25963,N_25005,N_25069);
xor U25964 (N_25964,N_25364,N_25053);
nand U25965 (N_25965,N_25304,N_25001);
and U25966 (N_25966,N_25148,N_25246);
nor U25967 (N_25967,N_25407,N_25382);
nor U25968 (N_25968,N_25488,N_25098);
and U25969 (N_25969,N_25263,N_25468);
or U25970 (N_25970,N_25449,N_25382);
xnor U25971 (N_25971,N_25094,N_25378);
nand U25972 (N_25972,N_25420,N_25133);
xor U25973 (N_25973,N_25190,N_25342);
nand U25974 (N_25974,N_25331,N_25466);
nor U25975 (N_25975,N_25180,N_25381);
xnor U25976 (N_25976,N_25393,N_25397);
or U25977 (N_25977,N_25292,N_25266);
nand U25978 (N_25978,N_25287,N_25411);
nand U25979 (N_25979,N_25139,N_25205);
nor U25980 (N_25980,N_25041,N_25271);
and U25981 (N_25981,N_25404,N_25388);
nand U25982 (N_25982,N_25490,N_25051);
xor U25983 (N_25983,N_25331,N_25126);
xor U25984 (N_25984,N_25027,N_25406);
xor U25985 (N_25985,N_25060,N_25005);
or U25986 (N_25986,N_25441,N_25296);
nor U25987 (N_25987,N_25443,N_25385);
and U25988 (N_25988,N_25438,N_25363);
and U25989 (N_25989,N_25188,N_25098);
or U25990 (N_25990,N_25192,N_25359);
nor U25991 (N_25991,N_25174,N_25441);
nand U25992 (N_25992,N_25427,N_25336);
and U25993 (N_25993,N_25464,N_25190);
xor U25994 (N_25994,N_25078,N_25310);
nor U25995 (N_25995,N_25043,N_25422);
nand U25996 (N_25996,N_25133,N_25314);
nor U25997 (N_25997,N_25492,N_25209);
or U25998 (N_25998,N_25383,N_25288);
and U25999 (N_25999,N_25016,N_25287);
or U26000 (N_26000,N_25600,N_25908);
or U26001 (N_26001,N_25892,N_25794);
nand U26002 (N_26002,N_25901,N_25996);
or U26003 (N_26003,N_25700,N_25648);
nand U26004 (N_26004,N_25880,N_25638);
and U26005 (N_26005,N_25503,N_25894);
or U26006 (N_26006,N_25768,N_25691);
nand U26007 (N_26007,N_25599,N_25866);
xor U26008 (N_26008,N_25909,N_25893);
or U26009 (N_26009,N_25564,N_25764);
or U26010 (N_26010,N_25929,N_25834);
xnor U26011 (N_26011,N_25873,N_25955);
nor U26012 (N_26012,N_25651,N_25591);
nor U26013 (N_26013,N_25555,N_25655);
and U26014 (N_26014,N_25505,N_25823);
nor U26015 (N_26015,N_25731,N_25981);
xor U26016 (N_26016,N_25742,N_25608);
nor U26017 (N_26017,N_25515,N_25863);
or U26018 (N_26018,N_25728,N_25628);
and U26019 (N_26019,N_25560,N_25891);
and U26020 (N_26020,N_25524,N_25705);
xor U26021 (N_26021,N_25766,N_25641);
nand U26022 (N_26022,N_25843,N_25623);
xor U26023 (N_26023,N_25669,N_25750);
nor U26024 (N_26024,N_25722,N_25676);
and U26025 (N_26025,N_25601,N_25983);
nand U26026 (N_26026,N_25551,N_25952);
and U26027 (N_26027,N_25542,N_25825);
nand U26028 (N_26028,N_25785,N_25851);
or U26029 (N_26029,N_25887,N_25947);
nor U26030 (N_26030,N_25788,N_25985);
xnor U26031 (N_26031,N_25737,N_25609);
nand U26032 (N_26032,N_25906,N_25500);
nor U26033 (N_26033,N_25805,N_25590);
or U26034 (N_26034,N_25864,N_25614);
and U26035 (N_26035,N_25944,N_25718);
nor U26036 (N_26036,N_25632,N_25663);
nand U26037 (N_26037,N_25882,N_25987);
xor U26038 (N_26038,N_25808,N_25773);
xor U26039 (N_26039,N_25890,N_25652);
and U26040 (N_26040,N_25620,N_25568);
and U26041 (N_26041,N_25937,N_25791);
nand U26042 (N_26042,N_25888,N_25814);
xor U26043 (N_26043,N_25525,N_25685);
nand U26044 (N_26044,N_25790,N_25535);
or U26045 (N_26045,N_25978,N_25656);
nor U26046 (N_26046,N_25506,N_25980);
or U26047 (N_26047,N_25842,N_25635);
nor U26048 (N_26048,N_25964,N_25803);
nand U26049 (N_26049,N_25777,N_25917);
nand U26050 (N_26050,N_25537,N_25580);
and U26051 (N_26051,N_25670,N_25789);
nand U26052 (N_26052,N_25876,N_25857);
xnor U26053 (N_26053,N_25820,N_25684);
xnor U26054 (N_26054,N_25567,N_25925);
xnor U26055 (N_26055,N_25569,N_25703);
xor U26056 (N_26056,N_25819,N_25693);
or U26057 (N_26057,N_25778,N_25885);
nand U26058 (N_26058,N_25799,N_25786);
nor U26059 (N_26059,N_25714,N_25593);
or U26060 (N_26060,N_25715,N_25853);
and U26061 (N_26061,N_25833,N_25698);
nand U26062 (N_26062,N_25939,N_25727);
xor U26063 (N_26063,N_25962,N_25840);
xnor U26064 (N_26064,N_25668,N_25918);
nand U26065 (N_26065,N_25531,N_25674);
xnor U26066 (N_26066,N_25919,N_25709);
or U26067 (N_26067,N_25527,N_25683);
or U26068 (N_26068,N_25874,N_25994);
nor U26069 (N_26069,N_25639,N_25875);
and U26070 (N_26070,N_25877,N_25736);
xor U26071 (N_26071,N_25854,N_25837);
or U26072 (N_26072,N_25859,N_25561);
nor U26073 (N_26073,N_25538,N_25606);
nand U26074 (N_26074,N_25659,N_25975);
xor U26075 (N_26075,N_25924,N_25589);
and U26076 (N_26076,N_25896,N_25692);
xor U26077 (N_26077,N_25920,N_25749);
nor U26078 (N_26078,N_25634,N_25508);
and U26079 (N_26079,N_25578,N_25583);
nand U26080 (N_26080,N_25534,N_25966);
xnor U26081 (N_26081,N_25811,N_25661);
nor U26082 (N_26082,N_25815,N_25526);
or U26083 (N_26083,N_25626,N_25690);
xnor U26084 (N_26084,N_25686,N_25549);
nand U26085 (N_26085,N_25809,N_25587);
nor U26086 (N_26086,N_25940,N_25830);
and U26087 (N_26087,N_25780,N_25642);
and U26088 (N_26088,N_25543,N_25867);
xnor U26089 (N_26089,N_25563,N_25558);
nor U26090 (N_26090,N_25774,N_25984);
xor U26091 (N_26091,N_25776,N_25598);
and U26092 (N_26092,N_25817,N_25566);
nor U26093 (N_26093,N_25574,N_25895);
nand U26094 (N_26094,N_25979,N_25657);
nand U26095 (N_26095,N_25592,N_25547);
nor U26096 (N_26096,N_25935,N_25724);
nand U26097 (N_26097,N_25701,N_25681);
nand U26098 (N_26098,N_25629,N_25914);
and U26099 (N_26099,N_25577,N_25695);
nand U26100 (N_26100,N_25689,N_25782);
nand U26101 (N_26101,N_25904,N_25511);
nand U26102 (N_26102,N_25710,N_25730);
or U26103 (N_26103,N_25713,N_25631);
xnor U26104 (N_26104,N_25579,N_25910);
nor U26105 (N_26105,N_25618,N_25998);
nand U26106 (N_26106,N_25946,N_25930);
and U26107 (N_26107,N_25702,N_25848);
and U26108 (N_26108,N_25586,N_25872);
nor U26109 (N_26109,N_25771,N_25793);
and U26110 (N_26110,N_25800,N_25868);
nand U26111 (N_26111,N_25915,N_25550);
or U26112 (N_26112,N_25576,N_25616);
xnor U26113 (N_26113,N_25509,N_25959);
or U26114 (N_26114,N_25662,N_25565);
and U26115 (N_26115,N_25796,N_25716);
nor U26116 (N_26116,N_25798,N_25826);
xor U26117 (N_26117,N_25779,N_25839);
xor U26118 (N_26118,N_25832,N_25957);
or U26119 (N_26119,N_25625,N_25660);
nand U26120 (N_26120,N_25529,N_25951);
and U26121 (N_26121,N_25611,N_25871);
and U26122 (N_26122,N_25516,N_25643);
xor U26123 (N_26123,N_25640,N_25938);
and U26124 (N_26124,N_25645,N_25767);
nand U26125 (N_26125,N_25835,N_25688);
xnor U26126 (N_26126,N_25649,N_25769);
or U26127 (N_26127,N_25824,N_25934);
or U26128 (N_26128,N_25741,N_25729);
and U26129 (N_26129,N_25781,N_25630);
or U26130 (N_26130,N_25671,N_25562);
xor U26131 (N_26131,N_25943,N_25510);
xor U26132 (N_26132,N_25637,N_25816);
nand U26133 (N_26133,N_25760,N_25536);
and U26134 (N_26134,N_25926,N_25812);
nor U26135 (N_26135,N_25968,N_25912);
xnor U26136 (N_26136,N_25666,N_25810);
or U26137 (N_26137,N_25725,N_25995);
or U26138 (N_26138,N_25723,N_25818);
and U26139 (N_26139,N_25928,N_25763);
nor U26140 (N_26140,N_25862,N_25707);
xnor U26141 (N_26141,N_25949,N_25664);
nand U26142 (N_26142,N_25673,N_25879);
xnor U26143 (N_26143,N_25617,N_25739);
xor U26144 (N_26144,N_25588,N_25612);
nor U26145 (N_26145,N_25519,N_25932);
xor U26146 (N_26146,N_25687,N_25855);
nand U26147 (N_26147,N_25581,N_25502);
nand U26148 (N_26148,N_25988,N_25712);
or U26149 (N_26149,N_25953,N_25604);
and U26150 (N_26150,N_25927,N_25594);
or U26151 (N_26151,N_25976,N_25522);
nand U26152 (N_26152,N_25532,N_25615);
or U26153 (N_26153,N_25967,N_25571);
xor U26154 (N_26154,N_25677,N_25748);
nand U26155 (N_26155,N_25554,N_25992);
or U26156 (N_26156,N_25807,N_25784);
or U26157 (N_26157,N_25762,N_25504);
and U26158 (N_26158,N_25921,N_25514);
xnor U26159 (N_26159,N_25758,N_25878);
and U26160 (N_26160,N_25679,N_25933);
or U26161 (N_26161,N_25883,N_25720);
nor U26162 (N_26162,N_25989,N_25675);
and U26163 (N_26163,N_25726,N_25732);
nand U26164 (N_26164,N_25621,N_25694);
nor U26165 (N_26165,N_25956,N_25546);
nor U26166 (N_26166,N_25597,N_25821);
nor U26167 (N_26167,N_25922,N_25570);
or U26168 (N_26168,N_25958,N_25772);
nor U26169 (N_26169,N_25977,N_25861);
nand U26170 (N_26170,N_25665,N_25636);
xor U26171 (N_26171,N_25556,N_25521);
and U26172 (N_26172,N_25745,N_25624);
xor U26173 (N_26173,N_25738,N_25838);
nor U26174 (N_26174,N_25552,N_25595);
and U26175 (N_26175,N_25787,N_25619);
or U26176 (N_26176,N_25517,N_25813);
or U26177 (N_26177,N_25540,N_25513);
or U26178 (N_26178,N_25865,N_25905);
and U26179 (N_26179,N_25942,N_25870);
nand U26180 (N_26180,N_25801,N_25582);
or U26181 (N_26181,N_25858,N_25783);
or U26182 (N_26182,N_25733,N_25841);
xnor U26183 (N_26183,N_25969,N_25545);
xnor U26184 (N_26184,N_25847,N_25548);
and U26185 (N_26185,N_25907,N_25539);
nor U26186 (N_26186,N_25795,N_25973);
nand U26187 (N_26187,N_25775,N_25916);
and U26188 (N_26188,N_25607,N_25913);
xnor U26189 (N_26189,N_25849,N_25902);
nand U26190 (N_26190,N_25881,N_25530);
nand U26191 (N_26191,N_25734,N_25610);
nand U26192 (N_26192,N_25804,N_25644);
nor U26193 (N_26193,N_25697,N_25982);
or U26194 (N_26194,N_25633,N_25706);
or U26195 (N_26195,N_25936,N_25584);
or U26196 (N_26196,N_25735,N_25757);
or U26197 (N_26197,N_25699,N_25856);
xor U26198 (N_26198,N_25654,N_25553);
xor U26199 (N_26199,N_25899,N_25869);
or U26200 (N_26200,N_25802,N_25523);
nor U26201 (N_26201,N_25828,N_25948);
nand U26202 (N_26202,N_25647,N_25603);
nand U26203 (N_26203,N_25528,N_25754);
and U26204 (N_26204,N_25708,N_25667);
or U26205 (N_26205,N_25605,N_25646);
or U26206 (N_26206,N_25831,N_25696);
nor U26207 (N_26207,N_25993,N_25575);
nand U26208 (N_26208,N_25622,N_25974);
nor U26209 (N_26209,N_25756,N_25886);
nand U26210 (N_26210,N_25682,N_25931);
nor U26211 (N_26211,N_25596,N_25844);
xnor U26212 (N_26212,N_25761,N_25573);
or U26213 (N_26213,N_25518,N_25963);
and U26214 (N_26214,N_25965,N_25672);
nor U26215 (N_26215,N_25743,N_25752);
and U26216 (N_26216,N_25845,N_25827);
nor U26217 (N_26217,N_25884,N_25889);
nor U26218 (N_26218,N_25900,N_25711);
or U26219 (N_26219,N_25923,N_25755);
or U26220 (N_26220,N_25759,N_25746);
and U26221 (N_26221,N_25991,N_25602);
or U26222 (N_26222,N_25897,N_25770);
xor U26223 (N_26223,N_25860,N_25613);
xnor U26224 (N_26224,N_25740,N_25544);
xor U26225 (N_26225,N_25751,N_25986);
and U26226 (N_26226,N_25747,N_25792);
xnor U26227 (N_26227,N_25717,N_25627);
nor U26228 (N_26228,N_25572,N_25678);
nor U26229 (N_26229,N_25520,N_25765);
nor U26230 (N_26230,N_25954,N_25971);
and U26231 (N_26231,N_25806,N_25846);
nor U26232 (N_26232,N_25970,N_25950);
or U26233 (N_26233,N_25945,N_25990);
or U26234 (N_26234,N_25960,N_25797);
or U26235 (N_26235,N_25680,N_25822);
xor U26236 (N_26236,N_25650,N_25507);
nand U26237 (N_26237,N_25997,N_25829);
and U26238 (N_26238,N_25852,N_25850);
and U26239 (N_26239,N_25999,N_25898);
xor U26240 (N_26240,N_25961,N_25559);
nor U26241 (N_26241,N_25541,N_25903);
xnor U26242 (N_26242,N_25744,N_25972);
or U26243 (N_26243,N_25658,N_25585);
or U26244 (N_26244,N_25512,N_25719);
or U26245 (N_26245,N_25911,N_25836);
xnor U26246 (N_26246,N_25753,N_25557);
or U26247 (N_26247,N_25501,N_25941);
nand U26248 (N_26248,N_25533,N_25721);
xnor U26249 (N_26249,N_25704,N_25653);
or U26250 (N_26250,N_25770,N_25787);
nor U26251 (N_26251,N_25900,N_25654);
nand U26252 (N_26252,N_25740,N_25745);
and U26253 (N_26253,N_25958,N_25923);
or U26254 (N_26254,N_25582,N_25699);
or U26255 (N_26255,N_25839,N_25897);
xnor U26256 (N_26256,N_25866,N_25543);
nor U26257 (N_26257,N_25554,N_25514);
and U26258 (N_26258,N_25945,N_25756);
and U26259 (N_26259,N_25756,N_25866);
and U26260 (N_26260,N_25647,N_25916);
nand U26261 (N_26261,N_25955,N_25567);
nand U26262 (N_26262,N_25657,N_25995);
xor U26263 (N_26263,N_25666,N_25771);
or U26264 (N_26264,N_25765,N_25766);
xnor U26265 (N_26265,N_25668,N_25597);
nor U26266 (N_26266,N_25979,N_25839);
or U26267 (N_26267,N_25681,N_25953);
xnor U26268 (N_26268,N_25935,N_25642);
or U26269 (N_26269,N_25966,N_25573);
xnor U26270 (N_26270,N_25527,N_25682);
nand U26271 (N_26271,N_25966,N_25835);
and U26272 (N_26272,N_25624,N_25622);
and U26273 (N_26273,N_25997,N_25652);
nor U26274 (N_26274,N_25619,N_25735);
nor U26275 (N_26275,N_25609,N_25797);
and U26276 (N_26276,N_25623,N_25624);
nor U26277 (N_26277,N_25942,N_25874);
or U26278 (N_26278,N_25555,N_25800);
and U26279 (N_26279,N_25994,N_25989);
or U26280 (N_26280,N_25597,N_25586);
and U26281 (N_26281,N_25986,N_25667);
nor U26282 (N_26282,N_25836,N_25758);
and U26283 (N_26283,N_25520,N_25742);
xor U26284 (N_26284,N_25748,N_25819);
nor U26285 (N_26285,N_25504,N_25809);
xnor U26286 (N_26286,N_25567,N_25758);
xnor U26287 (N_26287,N_25848,N_25968);
nand U26288 (N_26288,N_25541,N_25949);
or U26289 (N_26289,N_25642,N_25548);
xnor U26290 (N_26290,N_25992,N_25622);
nor U26291 (N_26291,N_25763,N_25868);
or U26292 (N_26292,N_25779,N_25894);
or U26293 (N_26293,N_25978,N_25792);
or U26294 (N_26294,N_25943,N_25979);
and U26295 (N_26295,N_25577,N_25694);
and U26296 (N_26296,N_25568,N_25981);
and U26297 (N_26297,N_25757,N_25677);
nor U26298 (N_26298,N_25516,N_25929);
nor U26299 (N_26299,N_25807,N_25654);
xnor U26300 (N_26300,N_25534,N_25721);
nand U26301 (N_26301,N_25755,N_25561);
xor U26302 (N_26302,N_25822,N_25951);
nor U26303 (N_26303,N_25534,N_25686);
or U26304 (N_26304,N_25723,N_25821);
nor U26305 (N_26305,N_25909,N_25748);
nand U26306 (N_26306,N_25611,N_25695);
or U26307 (N_26307,N_25760,N_25568);
or U26308 (N_26308,N_25947,N_25586);
xnor U26309 (N_26309,N_25639,N_25882);
and U26310 (N_26310,N_25735,N_25736);
nor U26311 (N_26311,N_25670,N_25780);
nand U26312 (N_26312,N_25877,N_25976);
nand U26313 (N_26313,N_25798,N_25658);
xnor U26314 (N_26314,N_25722,N_25692);
or U26315 (N_26315,N_25734,N_25880);
nor U26316 (N_26316,N_25975,N_25539);
or U26317 (N_26317,N_25812,N_25726);
nor U26318 (N_26318,N_25860,N_25735);
and U26319 (N_26319,N_25756,N_25589);
and U26320 (N_26320,N_25870,N_25925);
nor U26321 (N_26321,N_25893,N_25706);
nor U26322 (N_26322,N_25734,N_25748);
or U26323 (N_26323,N_25984,N_25908);
and U26324 (N_26324,N_25587,N_25658);
nand U26325 (N_26325,N_25601,N_25642);
or U26326 (N_26326,N_25626,N_25679);
nand U26327 (N_26327,N_25818,N_25900);
nand U26328 (N_26328,N_25553,N_25958);
or U26329 (N_26329,N_25758,N_25626);
nand U26330 (N_26330,N_25647,N_25772);
or U26331 (N_26331,N_25844,N_25526);
or U26332 (N_26332,N_25673,N_25509);
and U26333 (N_26333,N_25527,N_25891);
and U26334 (N_26334,N_25901,N_25552);
nor U26335 (N_26335,N_25577,N_25654);
nor U26336 (N_26336,N_25955,N_25859);
nand U26337 (N_26337,N_25829,N_25709);
or U26338 (N_26338,N_25582,N_25888);
nor U26339 (N_26339,N_25822,N_25914);
nand U26340 (N_26340,N_25850,N_25593);
nand U26341 (N_26341,N_25506,N_25526);
and U26342 (N_26342,N_25532,N_25889);
nor U26343 (N_26343,N_25699,N_25934);
nand U26344 (N_26344,N_25571,N_25548);
nand U26345 (N_26345,N_25891,N_25996);
xnor U26346 (N_26346,N_25966,N_25985);
xor U26347 (N_26347,N_25784,N_25823);
nor U26348 (N_26348,N_25902,N_25801);
or U26349 (N_26349,N_25607,N_25853);
or U26350 (N_26350,N_25785,N_25598);
nor U26351 (N_26351,N_25510,N_25999);
and U26352 (N_26352,N_25865,N_25504);
nand U26353 (N_26353,N_25937,N_25517);
nand U26354 (N_26354,N_25602,N_25635);
and U26355 (N_26355,N_25639,N_25711);
nand U26356 (N_26356,N_25515,N_25640);
nor U26357 (N_26357,N_25553,N_25532);
nor U26358 (N_26358,N_25861,N_25974);
nand U26359 (N_26359,N_25775,N_25573);
nor U26360 (N_26360,N_25980,N_25750);
nand U26361 (N_26361,N_25764,N_25674);
nor U26362 (N_26362,N_25518,N_25547);
xnor U26363 (N_26363,N_25915,N_25981);
xnor U26364 (N_26364,N_25541,N_25951);
and U26365 (N_26365,N_25946,N_25972);
nor U26366 (N_26366,N_25948,N_25837);
xor U26367 (N_26367,N_25640,N_25873);
nor U26368 (N_26368,N_25905,N_25887);
or U26369 (N_26369,N_25542,N_25516);
xor U26370 (N_26370,N_25688,N_25658);
or U26371 (N_26371,N_25555,N_25987);
nand U26372 (N_26372,N_25659,N_25710);
xor U26373 (N_26373,N_25858,N_25727);
xor U26374 (N_26374,N_25724,N_25847);
nand U26375 (N_26375,N_25867,N_25639);
xnor U26376 (N_26376,N_25685,N_25861);
or U26377 (N_26377,N_25991,N_25935);
nor U26378 (N_26378,N_25518,N_25759);
nand U26379 (N_26379,N_25999,N_25839);
or U26380 (N_26380,N_25696,N_25522);
nor U26381 (N_26381,N_25915,N_25522);
xor U26382 (N_26382,N_25502,N_25603);
and U26383 (N_26383,N_25540,N_25795);
xor U26384 (N_26384,N_25936,N_25738);
nor U26385 (N_26385,N_25943,N_25630);
or U26386 (N_26386,N_25901,N_25979);
and U26387 (N_26387,N_25506,N_25546);
nand U26388 (N_26388,N_25797,N_25752);
xor U26389 (N_26389,N_25539,N_25954);
xor U26390 (N_26390,N_25957,N_25540);
nor U26391 (N_26391,N_25961,N_25706);
nor U26392 (N_26392,N_25856,N_25512);
and U26393 (N_26393,N_25592,N_25673);
or U26394 (N_26394,N_25826,N_25639);
and U26395 (N_26395,N_25905,N_25969);
nor U26396 (N_26396,N_25668,N_25907);
nand U26397 (N_26397,N_25683,N_25826);
or U26398 (N_26398,N_25996,N_25871);
nand U26399 (N_26399,N_25796,N_25531);
nand U26400 (N_26400,N_25957,N_25639);
nor U26401 (N_26401,N_25504,N_25986);
or U26402 (N_26402,N_25521,N_25628);
and U26403 (N_26403,N_25973,N_25693);
or U26404 (N_26404,N_25687,N_25848);
and U26405 (N_26405,N_25843,N_25745);
nand U26406 (N_26406,N_25862,N_25937);
and U26407 (N_26407,N_25686,N_25841);
or U26408 (N_26408,N_25831,N_25825);
xnor U26409 (N_26409,N_25576,N_25916);
xor U26410 (N_26410,N_25897,N_25648);
nand U26411 (N_26411,N_25870,N_25525);
xnor U26412 (N_26412,N_25741,N_25519);
nand U26413 (N_26413,N_25709,N_25555);
nor U26414 (N_26414,N_25710,N_25920);
xnor U26415 (N_26415,N_25820,N_25852);
or U26416 (N_26416,N_25509,N_25710);
and U26417 (N_26417,N_25867,N_25653);
xor U26418 (N_26418,N_25927,N_25931);
or U26419 (N_26419,N_25875,N_25950);
nand U26420 (N_26420,N_25584,N_25726);
and U26421 (N_26421,N_25947,N_25750);
xnor U26422 (N_26422,N_25916,N_25535);
nand U26423 (N_26423,N_25722,N_25912);
xor U26424 (N_26424,N_25582,N_25637);
xnor U26425 (N_26425,N_25904,N_25751);
nor U26426 (N_26426,N_25955,N_25756);
nand U26427 (N_26427,N_25880,N_25961);
nor U26428 (N_26428,N_25626,N_25503);
xnor U26429 (N_26429,N_25624,N_25687);
xor U26430 (N_26430,N_25775,N_25823);
nand U26431 (N_26431,N_25968,N_25923);
nand U26432 (N_26432,N_25538,N_25714);
and U26433 (N_26433,N_25930,N_25580);
xor U26434 (N_26434,N_25804,N_25735);
and U26435 (N_26435,N_25785,N_25651);
and U26436 (N_26436,N_25572,N_25795);
nand U26437 (N_26437,N_25843,N_25930);
or U26438 (N_26438,N_25565,N_25879);
xor U26439 (N_26439,N_25628,N_25759);
xnor U26440 (N_26440,N_25625,N_25553);
nor U26441 (N_26441,N_25927,N_25620);
or U26442 (N_26442,N_25891,N_25553);
xor U26443 (N_26443,N_25995,N_25716);
nor U26444 (N_26444,N_25972,N_25598);
nor U26445 (N_26445,N_25836,N_25614);
xor U26446 (N_26446,N_25970,N_25945);
and U26447 (N_26447,N_25583,N_25620);
xor U26448 (N_26448,N_25549,N_25985);
xor U26449 (N_26449,N_25981,N_25838);
or U26450 (N_26450,N_25578,N_25850);
xor U26451 (N_26451,N_25855,N_25591);
nor U26452 (N_26452,N_25689,N_25884);
nand U26453 (N_26453,N_25944,N_25605);
xor U26454 (N_26454,N_25700,N_25551);
xnor U26455 (N_26455,N_25889,N_25795);
nand U26456 (N_26456,N_25668,N_25655);
nand U26457 (N_26457,N_25705,N_25587);
and U26458 (N_26458,N_25742,N_25665);
nor U26459 (N_26459,N_25891,N_25967);
nand U26460 (N_26460,N_25743,N_25802);
xnor U26461 (N_26461,N_25755,N_25645);
nand U26462 (N_26462,N_25993,N_25671);
nor U26463 (N_26463,N_25726,N_25521);
nand U26464 (N_26464,N_25946,N_25919);
and U26465 (N_26465,N_25954,N_25660);
or U26466 (N_26466,N_25569,N_25668);
nand U26467 (N_26467,N_25820,N_25842);
and U26468 (N_26468,N_25659,N_25592);
nor U26469 (N_26469,N_25606,N_25910);
and U26470 (N_26470,N_25900,N_25525);
nand U26471 (N_26471,N_25824,N_25926);
nand U26472 (N_26472,N_25837,N_25805);
xnor U26473 (N_26473,N_25773,N_25715);
and U26474 (N_26474,N_25537,N_25835);
or U26475 (N_26475,N_25732,N_25652);
and U26476 (N_26476,N_25969,N_25659);
and U26477 (N_26477,N_25874,N_25811);
and U26478 (N_26478,N_25817,N_25747);
nor U26479 (N_26479,N_25824,N_25938);
and U26480 (N_26480,N_25901,N_25962);
xnor U26481 (N_26481,N_25865,N_25852);
nand U26482 (N_26482,N_25642,N_25537);
or U26483 (N_26483,N_25748,N_25792);
nor U26484 (N_26484,N_25717,N_25812);
nand U26485 (N_26485,N_25938,N_25794);
nand U26486 (N_26486,N_25891,N_25951);
or U26487 (N_26487,N_25519,N_25603);
nor U26488 (N_26488,N_25787,N_25968);
nor U26489 (N_26489,N_25866,N_25783);
xor U26490 (N_26490,N_25978,N_25816);
xor U26491 (N_26491,N_25703,N_25617);
and U26492 (N_26492,N_25582,N_25721);
and U26493 (N_26493,N_25975,N_25749);
nor U26494 (N_26494,N_25978,N_25961);
nand U26495 (N_26495,N_25976,N_25518);
xor U26496 (N_26496,N_25693,N_25781);
xnor U26497 (N_26497,N_25514,N_25750);
xnor U26498 (N_26498,N_25704,N_25613);
or U26499 (N_26499,N_25604,N_25590);
nor U26500 (N_26500,N_26067,N_26258);
nor U26501 (N_26501,N_26068,N_26119);
xnor U26502 (N_26502,N_26193,N_26399);
nand U26503 (N_26503,N_26183,N_26162);
or U26504 (N_26504,N_26489,N_26314);
nand U26505 (N_26505,N_26156,N_26495);
and U26506 (N_26506,N_26187,N_26407);
xor U26507 (N_26507,N_26313,N_26262);
or U26508 (N_26508,N_26134,N_26225);
nor U26509 (N_26509,N_26369,N_26202);
nand U26510 (N_26510,N_26390,N_26205);
and U26511 (N_26511,N_26397,N_26159);
and U26512 (N_26512,N_26403,N_26084);
xor U26513 (N_26513,N_26124,N_26411);
nand U26514 (N_26514,N_26113,N_26158);
xnor U26515 (N_26515,N_26039,N_26227);
nor U26516 (N_26516,N_26102,N_26022);
and U26517 (N_26517,N_26412,N_26080);
nand U26518 (N_26518,N_26016,N_26437);
nand U26519 (N_26519,N_26085,N_26035);
or U26520 (N_26520,N_26107,N_26059);
nor U26521 (N_26521,N_26378,N_26062);
or U26522 (N_26522,N_26027,N_26430);
nand U26523 (N_26523,N_26478,N_26337);
xor U26524 (N_26524,N_26402,N_26295);
nand U26525 (N_26525,N_26329,N_26150);
xnor U26526 (N_26526,N_26223,N_26045);
xnor U26527 (N_26527,N_26398,N_26484);
nor U26528 (N_26528,N_26154,N_26466);
nor U26529 (N_26529,N_26194,N_26093);
or U26530 (N_26530,N_26289,N_26488);
nand U26531 (N_26531,N_26429,N_26191);
or U26532 (N_26532,N_26286,N_26151);
or U26533 (N_26533,N_26356,N_26438);
and U26534 (N_26534,N_26136,N_26307);
or U26535 (N_26535,N_26335,N_26100);
and U26536 (N_26536,N_26155,N_26074);
xor U26537 (N_26537,N_26097,N_26081);
xnor U26538 (N_26538,N_26011,N_26481);
and U26539 (N_26539,N_26005,N_26052);
nand U26540 (N_26540,N_26334,N_26228);
and U26541 (N_26541,N_26216,N_26328);
xnor U26542 (N_26542,N_26239,N_26254);
or U26543 (N_26543,N_26196,N_26463);
and U26544 (N_26544,N_26199,N_26259);
nand U26545 (N_26545,N_26304,N_26315);
and U26546 (N_26546,N_26070,N_26298);
and U26547 (N_26547,N_26171,N_26336);
nand U26548 (N_26548,N_26123,N_26387);
nor U26549 (N_26549,N_26371,N_26230);
nand U26550 (N_26550,N_26181,N_26401);
nor U26551 (N_26551,N_26445,N_26391);
and U26552 (N_26552,N_26203,N_26414);
nor U26553 (N_26553,N_26043,N_26053);
nor U26554 (N_26554,N_26094,N_26343);
nor U26555 (N_26555,N_26498,N_26008);
nor U26556 (N_26556,N_26088,N_26153);
and U26557 (N_26557,N_26330,N_26038);
xor U26558 (N_26558,N_26244,N_26044);
nand U26559 (N_26559,N_26101,N_26376);
nand U26560 (N_26560,N_26243,N_26490);
nand U26561 (N_26561,N_26121,N_26108);
or U26562 (N_26562,N_26198,N_26423);
nor U26563 (N_26563,N_26461,N_26130);
xor U26564 (N_26564,N_26160,N_26413);
and U26565 (N_26565,N_26351,N_26055);
nor U26566 (N_26566,N_26362,N_26098);
xor U26567 (N_26567,N_26241,N_26152);
or U26568 (N_26568,N_26260,N_26006);
nor U26569 (N_26569,N_26116,N_26273);
and U26570 (N_26570,N_26275,N_26341);
nand U26571 (N_26571,N_26057,N_26457);
or U26572 (N_26572,N_26188,N_26071);
nand U26573 (N_26573,N_26109,N_26179);
xor U26574 (N_26574,N_26416,N_26197);
nor U26575 (N_26575,N_26344,N_26050);
xor U26576 (N_26576,N_26157,N_26104);
or U26577 (N_26577,N_26034,N_26382);
or U26578 (N_26578,N_26049,N_26432);
nor U26579 (N_26579,N_26308,N_26082);
and U26580 (N_26580,N_26316,N_26089);
xor U26581 (N_26581,N_26069,N_26221);
and U26582 (N_26582,N_26238,N_26345);
and U26583 (N_26583,N_26213,N_26168);
nand U26584 (N_26584,N_26173,N_26145);
xnor U26585 (N_26585,N_26302,N_26299);
nor U26586 (N_26586,N_26246,N_26122);
and U26587 (N_26587,N_26083,N_26493);
and U26588 (N_26588,N_26452,N_26185);
xor U26589 (N_26589,N_26415,N_26340);
nand U26590 (N_26590,N_26066,N_26318);
or U26591 (N_26591,N_26296,N_26087);
xor U26592 (N_26592,N_26443,N_26353);
xnor U26593 (N_26593,N_26475,N_26032);
xor U26594 (N_26594,N_26499,N_26367);
xor U26595 (N_26595,N_26078,N_26110);
nand U26596 (N_26596,N_26224,N_26287);
nand U26597 (N_26597,N_26480,N_26099);
nand U26598 (N_26598,N_26249,N_26169);
and U26599 (N_26599,N_26389,N_26264);
xor U26600 (N_26600,N_26209,N_26294);
xnor U26601 (N_26601,N_26192,N_26352);
xor U26602 (N_26602,N_26469,N_26141);
and U26603 (N_26603,N_26211,N_26126);
and U26604 (N_26604,N_26031,N_26494);
and U26605 (N_26605,N_26139,N_26460);
xor U26606 (N_26606,N_26327,N_26447);
xor U26607 (N_26607,N_26132,N_26040);
and U26608 (N_26608,N_26002,N_26024);
nand U26609 (N_26609,N_26060,N_26394);
xnor U26610 (N_26610,N_26048,N_26143);
nor U26611 (N_26611,N_26346,N_26233);
nand U26612 (N_26612,N_26491,N_26410);
nand U26613 (N_26613,N_26496,N_26456);
or U26614 (N_26614,N_26373,N_26189);
or U26615 (N_26615,N_26476,N_26127);
nand U26616 (N_26616,N_26058,N_26009);
nor U26617 (N_26617,N_26013,N_26279);
nor U26618 (N_26618,N_26242,N_26272);
nand U26619 (N_26619,N_26231,N_26112);
and U26620 (N_26620,N_26129,N_26486);
xor U26621 (N_26621,N_26095,N_26366);
xnor U26622 (N_26622,N_26365,N_26148);
or U26623 (N_26623,N_26020,N_26061);
and U26624 (N_26624,N_26106,N_26255);
or U26625 (N_26625,N_26265,N_26218);
nand U26626 (N_26626,N_26170,N_26103);
nand U26627 (N_26627,N_26408,N_26096);
and U26628 (N_26628,N_26207,N_26282);
and U26629 (N_26629,N_26146,N_26424);
or U26630 (N_26630,N_26404,N_26140);
xor U26631 (N_26631,N_26485,N_26444);
or U26632 (N_26632,N_26248,N_26277);
and U26633 (N_26633,N_26470,N_26386);
or U26634 (N_26634,N_26453,N_26442);
and U26635 (N_26635,N_26274,N_26174);
nor U26636 (N_26636,N_26464,N_26291);
or U26637 (N_26637,N_26208,N_26014);
xor U26638 (N_26638,N_26131,N_26120);
nand U26639 (N_26639,N_26090,N_26497);
nand U26640 (N_26640,N_26036,N_26252);
xnor U26641 (N_26641,N_26017,N_26332);
nor U26642 (N_26642,N_26065,N_26285);
nand U26643 (N_26643,N_26138,N_26271);
nor U26644 (N_26644,N_26263,N_26492);
nor U26645 (N_26645,N_26392,N_26165);
nor U26646 (N_26646,N_26214,N_26030);
nand U26647 (N_26647,N_26210,N_26217);
nor U26648 (N_26648,N_26405,N_26305);
nor U26649 (N_26649,N_26306,N_26280);
xnor U26650 (N_26650,N_26025,N_26235);
nand U26651 (N_26651,N_26163,N_26473);
or U26652 (N_26652,N_26135,N_26482);
xnor U26653 (N_26653,N_26114,N_26317);
or U26654 (N_26654,N_26003,N_26180);
or U26655 (N_26655,N_26293,N_26363);
nand U26656 (N_26656,N_26086,N_26439);
and U26657 (N_26657,N_26417,N_26381);
nor U26658 (N_26658,N_26245,N_26322);
nor U26659 (N_26659,N_26076,N_26257);
or U26660 (N_26660,N_26396,N_26177);
nand U26661 (N_26661,N_26161,N_26418);
or U26662 (N_26662,N_26425,N_26250);
nand U26663 (N_26663,N_26350,N_26237);
xnor U26664 (N_26664,N_26338,N_26467);
xor U26665 (N_26665,N_26459,N_26182);
xnor U26666 (N_26666,N_26310,N_26427);
nor U26667 (N_26667,N_26281,N_26440);
xnor U26668 (N_26668,N_26247,N_26283);
nand U26669 (N_26669,N_26000,N_26349);
nand U26670 (N_26670,N_26270,N_26200);
nor U26671 (N_26671,N_26276,N_26474);
nand U26672 (N_26672,N_26320,N_26487);
nand U26673 (N_26673,N_26311,N_26001);
xnor U26674 (N_26674,N_26023,N_26364);
and U26675 (N_26675,N_26374,N_26454);
xor U26676 (N_26676,N_26021,N_26063);
or U26677 (N_26677,N_26325,N_26465);
nor U26678 (N_26678,N_26400,N_26184);
nor U26679 (N_26679,N_26377,N_26303);
nor U26680 (N_26680,N_26347,N_26360);
xor U26681 (N_26681,N_26175,N_26166);
xnor U26682 (N_26682,N_26072,N_26133);
xnor U26683 (N_26683,N_26051,N_26395);
and U26684 (N_26684,N_26015,N_26357);
nand U26685 (N_26685,N_26167,N_26393);
and U26686 (N_26686,N_26268,N_26370);
and U26687 (N_26687,N_26288,N_26240);
nor U26688 (N_26688,N_26018,N_26117);
xor U26689 (N_26689,N_26358,N_26149);
or U26690 (N_26690,N_26075,N_26375);
and U26691 (N_26691,N_26222,N_26385);
nand U26692 (N_26692,N_26331,N_26436);
and U26693 (N_26693,N_26128,N_26256);
nor U26694 (N_26694,N_26409,N_26195);
or U26695 (N_26695,N_26301,N_26007);
and U26696 (N_26696,N_26348,N_26118);
or U26697 (N_26697,N_26319,N_26219);
xor U26698 (N_26698,N_26321,N_26064);
and U26699 (N_26699,N_26426,N_26462);
and U26700 (N_26700,N_26041,N_26446);
and U26701 (N_26701,N_26278,N_26326);
xor U26702 (N_26702,N_26012,N_26312);
nand U26703 (N_26703,N_26309,N_26226);
and U26704 (N_26704,N_26419,N_26029);
nand U26705 (N_26705,N_26212,N_26284);
nor U26706 (N_26706,N_26379,N_26354);
nand U26707 (N_26707,N_26054,N_26267);
or U26708 (N_26708,N_26144,N_26406);
xor U26709 (N_26709,N_26042,N_26033);
or U26710 (N_26710,N_26434,N_26215);
or U26711 (N_26711,N_26232,N_26186);
nor U26712 (N_26712,N_26201,N_26046);
xnor U26713 (N_26713,N_26028,N_26142);
xnor U26714 (N_26714,N_26111,N_26251);
or U26715 (N_26715,N_26172,N_26483);
nand U26716 (N_26716,N_26448,N_26026);
xor U26717 (N_26717,N_26269,N_26450);
nand U26718 (N_26718,N_26220,N_26384);
or U26719 (N_26719,N_26458,N_26164);
and U26720 (N_26720,N_26324,N_26455);
or U26721 (N_26721,N_26204,N_26056);
xor U26722 (N_26722,N_26297,N_26004);
xor U26723 (N_26723,N_26372,N_26253);
and U26724 (N_26724,N_26236,N_26125);
or U26725 (N_26725,N_26092,N_26229);
and U26726 (N_26726,N_26323,N_26290);
xnor U26727 (N_26727,N_26388,N_26435);
and U26728 (N_26728,N_26368,N_26451);
nand U26729 (N_26729,N_26234,N_26355);
nor U26730 (N_26730,N_26359,N_26342);
or U26731 (N_26731,N_26091,N_26422);
and U26732 (N_26732,N_26176,N_26206);
xnor U26733 (N_26733,N_26178,N_26380);
xnor U26734 (N_26734,N_26472,N_26105);
nor U26735 (N_26735,N_26266,N_26421);
nor U26736 (N_26736,N_26037,N_26339);
and U26737 (N_26737,N_26449,N_26477);
or U26738 (N_26738,N_26115,N_26019);
nand U26739 (N_26739,N_26433,N_26190);
nand U26740 (N_26740,N_26010,N_26420);
xnor U26741 (N_26741,N_26383,N_26047);
nor U26742 (N_26742,N_26147,N_26471);
nand U26743 (N_26743,N_26073,N_26441);
and U26744 (N_26744,N_26468,N_26361);
nor U26745 (N_26745,N_26261,N_26479);
and U26746 (N_26746,N_26300,N_26077);
or U26747 (N_26747,N_26333,N_26079);
xnor U26748 (N_26748,N_26137,N_26431);
and U26749 (N_26749,N_26428,N_26292);
or U26750 (N_26750,N_26316,N_26234);
or U26751 (N_26751,N_26267,N_26019);
xnor U26752 (N_26752,N_26217,N_26410);
nand U26753 (N_26753,N_26461,N_26091);
xor U26754 (N_26754,N_26086,N_26252);
or U26755 (N_26755,N_26201,N_26404);
nand U26756 (N_26756,N_26266,N_26357);
xnor U26757 (N_26757,N_26049,N_26243);
or U26758 (N_26758,N_26231,N_26090);
nor U26759 (N_26759,N_26478,N_26292);
and U26760 (N_26760,N_26279,N_26198);
nor U26761 (N_26761,N_26407,N_26167);
nand U26762 (N_26762,N_26437,N_26317);
nand U26763 (N_26763,N_26123,N_26161);
xnor U26764 (N_26764,N_26264,N_26107);
or U26765 (N_26765,N_26131,N_26051);
nor U26766 (N_26766,N_26313,N_26312);
xnor U26767 (N_26767,N_26165,N_26434);
nand U26768 (N_26768,N_26314,N_26089);
nand U26769 (N_26769,N_26311,N_26120);
nor U26770 (N_26770,N_26006,N_26000);
nand U26771 (N_26771,N_26325,N_26093);
nor U26772 (N_26772,N_26230,N_26370);
nand U26773 (N_26773,N_26294,N_26076);
and U26774 (N_26774,N_26226,N_26148);
xnor U26775 (N_26775,N_26285,N_26371);
and U26776 (N_26776,N_26468,N_26480);
and U26777 (N_26777,N_26097,N_26186);
nor U26778 (N_26778,N_26080,N_26131);
xor U26779 (N_26779,N_26235,N_26177);
nor U26780 (N_26780,N_26317,N_26350);
and U26781 (N_26781,N_26464,N_26310);
or U26782 (N_26782,N_26461,N_26354);
and U26783 (N_26783,N_26485,N_26002);
or U26784 (N_26784,N_26021,N_26163);
nor U26785 (N_26785,N_26140,N_26305);
nand U26786 (N_26786,N_26454,N_26423);
and U26787 (N_26787,N_26062,N_26074);
nor U26788 (N_26788,N_26469,N_26326);
and U26789 (N_26789,N_26241,N_26388);
nor U26790 (N_26790,N_26463,N_26452);
and U26791 (N_26791,N_26199,N_26486);
nor U26792 (N_26792,N_26319,N_26131);
and U26793 (N_26793,N_26217,N_26483);
xnor U26794 (N_26794,N_26398,N_26423);
nor U26795 (N_26795,N_26405,N_26176);
nor U26796 (N_26796,N_26051,N_26210);
and U26797 (N_26797,N_26393,N_26065);
or U26798 (N_26798,N_26176,N_26358);
xnor U26799 (N_26799,N_26467,N_26134);
or U26800 (N_26800,N_26020,N_26415);
and U26801 (N_26801,N_26252,N_26367);
or U26802 (N_26802,N_26316,N_26166);
or U26803 (N_26803,N_26204,N_26193);
xnor U26804 (N_26804,N_26117,N_26476);
or U26805 (N_26805,N_26067,N_26409);
or U26806 (N_26806,N_26387,N_26155);
nor U26807 (N_26807,N_26235,N_26425);
or U26808 (N_26808,N_26294,N_26062);
nor U26809 (N_26809,N_26396,N_26275);
nor U26810 (N_26810,N_26498,N_26259);
nand U26811 (N_26811,N_26419,N_26119);
or U26812 (N_26812,N_26483,N_26397);
nor U26813 (N_26813,N_26410,N_26411);
xor U26814 (N_26814,N_26258,N_26122);
or U26815 (N_26815,N_26360,N_26468);
nand U26816 (N_26816,N_26152,N_26201);
and U26817 (N_26817,N_26405,N_26424);
nor U26818 (N_26818,N_26014,N_26080);
and U26819 (N_26819,N_26398,N_26107);
xnor U26820 (N_26820,N_26301,N_26178);
nor U26821 (N_26821,N_26498,N_26077);
nor U26822 (N_26822,N_26449,N_26065);
or U26823 (N_26823,N_26167,N_26106);
nand U26824 (N_26824,N_26481,N_26272);
or U26825 (N_26825,N_26417,N_26491);
or U26826 (N_26826,N_26087,N_26237);
xor U26827 (N_26827,N_26027,N_26473);
xor U26828 (N_26828,N_26429,N_26483);
nor U26829 (N_26829,N_26203,N_26286);
and U26830 (N_26830,N_26202,N_26235);
nand U26831 (N_26831,N_26020,N_26195);
nor U26832 (N_26832,N_26213,N_26183);
nand U26833 (N_26833,N_26058,N_26407);
and U26834 (N_26834,N_26040,N_26033);
nand U26835 (N_26835,N_26277,N_26249);
and U26836 (N_26836,N_26188,N_26147);
xor U26837 (N_26837,N_26293,N_26238);
and U26838 (N_26838,N_26211,N_26493);
and U26839 (N_26839,N_26483,N_26492);
or U26840 (N_26840,N_26289,N_26262);
nor U26841 (N_26841,N_26257,N_26229);
or U26842 (N_26842,N_26493,N_26023);
nor U26843 (N_26843,N_26078,N_26021);
or U26844 (N_26844,N_26152,N_26125);
and U26845 (N_26845,N_26253,N_26055);
or U26846 (N_26846,N_26249,N_26354);
and U26847 (N_26847,N_26188,N_26438);
nand U26848 (N_26848,N_26048,N_26466);
and U26849 (N_26849,N_26181,N_26143);
xor U26850 (N_26850,N_26257,N_26353);
xor U26851 (N_26851,N_26319,N_26203);
nor U26852 (N_26852,N_26268,N_26026);
nor U26853 (N_26853,N_26351,N_26158);
nand U26854 (N_26854,N_26453,N_26460);
and U26855 (N_26855,N_26496,N_26403);
xnor U26856 (N_26856,N_26369,N_26007);
or U26857 (N_26857,N_26091,N_26075);
or U26858 (N_26858,N_26005,N_26231);
and U26859 (N_26859,N_26479,N_26225);
and U26860 (N_26860,N_26131,N_26086);
nor U26861 (N_26861,N_26327,N_26255);
xnor U26862 (N_26862,N_26028,N_26104);
nor U26863 (N_26863,N_26176,N_26242);
and U26864 (N_26864,N_26293,N_26017);
nand U26865 (N_26865,N_26163,N_26047);
nor U26866 (N_26866,N_26120,N_26342);
xor U26867 (N_26867,N_26308,N_26075);
nor U26868 (N_26868,N_26201,N_26486);
xnor U26869 (N_26869,N_26031,N_26390);
and U26870 (N_26870,N_26046,N_26156);
and U26871 (N_26871,N_26159,N_26270);
or U26872 (N_26872,N_26358,N_26365);
xnor U26873 (N_26873,N_26474,N_26345);
nor U26874 (N_26874,N_26225,N_26403);
or U26875 (N_26875,N_26357,N_26174);
and U26876 (N_26876,N_26323,N_26082);
nor U26877 (N_26877,N_26497,N_26266);
or U26878 (N_26878,N_26164,N_26269);
and U26879 (N_26879,N_26182,N_26093);
and U26880 (N_26880,N_26377,N_26404);
and U26881 (N_26881,N_26143,N_26001);
and U26882 (N_26882,N_26112,N_26032);
and U26883 (N_26883,N_26198,N_26159);
nor U26884 (N_26884,N_26117,N_26248);
xor U26885 (N_26885,N_26298,N_26377);
or U26886 (N_26886,N_26182,N_26211);
nand U26887 (N_26887,N_26239,N_26247);
and U26888 (N_26888,N_26170,N_26136);
nand U26889 (N_26889,N_26344,N_26399);
xnor U26890 (N_26890,N_26278,N_26447);
nor U26891 (N_26891,N_26281,N_26413);
nand U26892 (N_26892,N_26184,N_26011);
nor U26893 (N_26893,N_26419,N_26426);
nand U26894 (N_26894,N_26207,N_26389);
and U26895 (N_26895,N_26121,N_26148);
xor U26896 (N_26896,N_26159,N_26022);
nand U26897 (N_26897,N_26245,N_26407);
nand U26898 (N_26898,N_26141,N_26198);
and U26899 (N_26899,N_26015,N_26212);
nand U26900 (N_26900,N_26158,N_26044);
and U26901 (N_26901,N_26170,N_26216);
nand U26902 (N_26902,N_26016,N_26359);
xnor U26903 (N_26903,N_26068,N_26220);
xor U26904 (N_26904,N_26117,N_26228);
or U26905 (N_26905,N_26498,N_26020);
nand U26906 (N_26906,N_26136,N_26138);
or U26907 (N_26907,N_26121,N_26016);
nand U26908 (N_26908,N_26209,N_26361);
or U26909 (N_26909,N_26278,N_26392);
or U26910 (N_26910,N_26395,N_26037);
or U26911 (N_26911,N_26390,N_26440);
or U26912 (N_26912,N_26335,N_26446);
or U26913 (N_26913,N_26393,N_26027);
nor U26914 (N_26914,N_26263,N_26430);
nand U26915 (N_26915,N_26237,N_26261);
or U26916 (N_26916,N_26462,N_26049);
nand U26917 (N_26917,N_26144,N_26180);
nor U26918 (N_26918,N_26384,N_26192);
nand U26919 (N_26919,N_26297,N_26278);
and U26920 (N_26920,N_26264,N_26306);
and U26921 (N_26921,N_26390,N_26358);
or U26922 (N_26922,N_26154,N_26264);
xnor U26923 (N_26923,N_26332,N_26324);
xnor U26924 (N_26924,N_26036,N_26128);
and U26925 (N_26925,N_26142,N_26284);
and U26926 (N_26926,N_26456,N_26035);
or U26927 (N_26927,N_26302,N_26041);
or U26928 (N_26928,N_26240,N_26479);
and U26929 (N_26929,N_26396,N_26020);
xor U26930 (N_26930,N_26087,N_26439);
nor U26931 (N_26931,N_26401,N_26429);
xnor U26932 (N_26932,N_26168,N_26214);
nor U26933 (N_26933,N_26300,N_26277);
nand U26934 (N_26934,N_26461,N_26459);
nand U26935 (N_26935,N_26382,N_26036);
xnor U26936 (N_26936,N_26240,N_26011);
xor U26937 (N_26937,N_26312,N_26383);
or U26938 (N_26938,N_26271,N_26044);
nor U26939 (N_26939,N_26139,N_26142);
and U26940 (N_26940,N_26091,N_26385);
nand U26941 (N_26941,N_26420,N_26272);
nor U26942 (N_26942,N_26146,N_26202);
xor U26943 (N_26943,N_26477,N_26380);
and U26944 (N_26944,N_26154,N_26487);
nand U26945 (N_26945,N_26197,N_26163);
or U26946 (N_26946,N_26110,N_26096);
xor U26947 (N_26947,N_26303,N_26157);
xor U26948 (N_26948,N_26300,N_26327);
and U26949 (N_26949,N_26022,N_26488);
nand U26950 (N_26950,N_26131,N_26007);
xnor U26951 (N_26951,N_26305,N_26271);
or U26952 (N_26952,N_26314,N_26054);
and U26953 (N_26953,N_26226,N_26185);
nand U26954 (N_26954,N_26413,N_26319);
or U26955 (N_26955,N_26395,N_26458);
and U26956 (N_26956,N_26469,N_26242);
nor U26957 (N_26957,N_26484,N_26252);
nor U26958 (N_26958,N_26117,N_26058);
and U26959 (N_26959,N_26430,N_26472);
and U26960 (N_26960,N_26169,N_26190);
nor U26961 (N_26961,N_26074,N_26032);
nor U26962 (N_26962,N_26392,N_26050);
nor U26963 (N_26963,N_26294,N_26428);
or U26964 (N_26964,N_26131,N_26134);
nand U26965 (N_26965,N_26342,N_26157);
and U26966 (N_26966,N_26487,N_26174);
or U26967 (N_26967,N_26450,N_26345);
or U26968 (N_26968,N_26209,N_26138);
and U26969 (N_26969,N_26448,N_26199);
nand U26970 (N_26970,N_26308,N_26257);
nor U26971 (N_26971,N_26487,N_26162);
nor U26972 (N_26972,N_26243,N_26322);
nor U26973 (N_26973,N_26238,N_26378);
or U26974 (N_26974,N_26238,N_26219);
or U26975 (N_26975,N_26176,N_26245);
xor U26976 (N_26976,N_26220,N_26471);
or U26977 (N_26977,N_26120,N_26072);
nand U26978 (N_26978,N_26387,N_26255);
and U26979 (N_26979,N_26423,N_26292);
xnor U26980 (N_26980,N_26421,N_26320);
xnor U26981 (N_26981,N_26069,N_26204);
nor U26982 (N_26982,N_26430,N_26096);
or U26983 (N_26983,N_26024,N_26482);
and U26984 (N_26984,N_26012,N_26313);
xnor U26985 (N_26985,N_26251,N_26320);
nand U26986 (N_26986,N_26424,N_26095);
nor U26987 (N_26987,N_26252,N_26394);
nand U26988 (N_26988,N_26465,N_26285);
nor U26989 (N_26989,N_26146,N_26484);
nor U26990 (N_26990,N_26205,N_26164);
xnor U26991 (N_26991,N_26181,N_26031);
nand U26992 (N_26992,N_26274,N_26166);
or U26993 (N_26993,N_26175,N_26195);
nor U26994 (N_26994,N_26005,N_26478);
nand U26995 (N_26995,N_26161,N_26107);
or U26996 (N_26996,N_26373,N_26207);
nand U26997 (N_26997,N_26310,N_26433);
nand U26998 (N_26998,N_26183,N_26125);
xor U26999 (N_26999,N_26355,N_26177);
nor U27000 (N_27000,N_26959,N_26571);
or U27001 (N_27001,N_26615,N_26549);
nand U27002 (N_27002,N_26568,N_26869);
nand U27003 (N_27003,N_26920,N_26552);
and U27004 (N_27004,N_26616,N_26888);
and U27005 (N_27005,N_26767,N_26508);
nor U27006 (N_27006,N_26621,N_26627);
xor U27007 (N_27007,N_26978,N_26611);
and U27008 (N_27008,N_26737,N_26749);
nand U27009 (N_27009,N_26642,N_26729);
nor U27010 (N_27010,N_26591,N_26822);
nor U27011 (N_27011,N_26646,N_26525);
nand U27012 (N_27012,N_26899,N_26894);
nor U27013 (N_27013,N_26847,N_26764);
or U27014 (N_27014,N_26942,N_26871);
nor U27015 (N_27015,N_26779,N_26861);
and U27016 (N_27016,N_26517,N_26747);
nor U27017 (N_27017,N_26579,N_26628);
nand U27018 (N_27018,N_26909,N_26710);
nor U27019 (N_27019,N_26940,N_26809);
or U27020 (N_27020,N_26643,N_26509);
nor U27021 (N_27021,N_26902,N_26532);
nor U27022 (N_27022,N_26863,N_26974);
nand U27023 (N_27023,N_26752,N_26722);
or U27024 (N_27024,N_26703,N_26964);
and U27025 (N_27025,N_26740,N_26651);
nor U27026 (N_27026,N_26711,N_26501);
nor U27027 (N_27027,N_26785,N_26801);
nand U27028 (N_27028,N_26707,N_26852);
or U27029 (N_27029,N_26626,N_26728);
and U27030 (N_27030,N_26715,N_26953);
and U27031 (N_27031,N_26991,N_26682);
nor U27032 (N_27032,N_26613,N_26606);
and U27033 (N_27033,N_26693,N_26792);
nand U27034 (N_27034,N_26567,N_26815);
and U27035 (N_27035,N_26622,N_26936);
nor U27036 (N_27036,N_26690,N_26840);
nand U27037 (N_27037,N_26855,N_26835);
xor U27038 (N_27038,N_26604,N_26772);
and U27039 (N_27039,N_26761,N_26521);
or U27040 (N_27040,N_26979,N_26506);
nor U27041 (N_27041,N_26988,N_26585);
or U27042 (N_27042,N_26935,N_26813);
nor U27043 (N_27043,N_26955,N_26857);
and U27044 (N_27044,N_26745,N_26912);
nand U27045 (N_27045,N_26897,N_26851);
or U27046 (N_27046,N_26967,N_26803);
xor U27047 (N_27047,N_26791,N_26562);
nor U27048 (N_27048,N_26575,N_26763);
nand U27049 (N_27049,N_26721,N_26687);
or U27050 (N_27050,N_26723,N_26545);
and U27051 (N_27051,N_26588,N_26757);
nand U27052 (N_27052,N_26896,N_26544);
or U27053 (N_27053,N_26529,N_26697);
nand U27054 (N_27054,N_26724,N_26793);
nor U27055 (N_27055,N_26584,N_26742);
xnor U27056 (N_27056,N_26702,N_26865);
nor U27057 (N_27057,N_26760,N_26895);
nor U27058 (N_27058,N_26636,N_26586);
nor U27059 (N_27059,N_26524,N_26790);
nor U27060 (N_27060,N_26546,N_26777);
and U27061 (N_27061,N_26582,N_26531);
nor U27062 (N_27062,N_26716,N_26713);
nor U27063 (N_27063,N_26797,N_26883);
and U27064 (N_27064,N_26679,N_26598);
nor U27065 (N_27065,N_26886,N_26539);
and U27066 (N_27066,N_26836,N_26918);
nor U27067 (N_27067,N_26898,N_26831);
and U27068 (N_27068,N_26589,N_26877);
or U27069 (N_27069,N_26830,N_26692);
or U27070 (N_27070,N_26624,N_26948);
or U27071 (N_27071,N_26971,N_26945);
and U27072 (N_27072,N_26558,N_26655);
xor U27073 (N_27073,N_26563,N_26890);
xor U27074 (N_27074,N_26972,N_26727);
xor U27075 (N_27075,N_26609,N_26607);
and U27076 (N_27076,N_26518,N_26720);
xor U27077 (N_27077,N_26812,N_26786);
nand U27078 (N_27078,N_26778,N_26961);
xnor U27079 (N_27079,N_26774,N_26572);
and U27080 (N_27080,N_26640,N_26676);
xor U27081 (N_27081,N_26998,N_26997);
or U27082 (N_27082,N_26800,N_26580);
nand U27083 (N_27083,N_26866,N_26798);
and U27084 (N_27084,N_26783,N_26770);
xnor U27085 (N_27085,N_26838,N_26956);
and U27086 (N_27086,N_26769,N_26969);
and U27087 (N_27087,N_26629,N_26817);
or U27088 (N_27088,N_26516,N_26893);
or U27089 (N_27089,N_26931,N_26534);
or U27090 (N_27090,N_26736,N_26592);
nor U27091 (N_27091,N_26553,N_26947);
and U27092 (N_27092,N_26590,N_26503);
nor U27093 (N_27093,N_26650,N_26827);
or U27094 (N_27094,N_26686,N_26677);
nand U27095 (N_27095,N_26977,N_26984);
nand U27096 (N_27096,N_26891,N_26907);
and U27097 (N_27097,N_26818,N_26708);
nand U27098 (N_27098,N_26905,N_26704);
or U27099 (N_27099,N_26867,N_26758);
nor U27100 (N_27100,N_26914,N_26528);
xnor U27101 (N_27101,N_26773,N_26673);
or U27102 (N_27102,N_26751,N_26725);
or U27103 (N_27103,N_26862,N_26832);
nor U27104 (N_27104,N_26846,N_26929);
and U27105 (N_27105,N_26637,N_26879);
xor U27106 (N_27106,N_26928,N_26634);
nor U27107 (N_27107,N_26685,N_26689);
or U27108 (N_27108,N_26939,N_26917);
and U27109 (N_27109,N_26927,N_26638);
and U27110 (N_27110,N_26806,N_26631);
and U27111 (N_27111,N_26674,N_26536);
nor U27112 (N_27112,N_26548,N_26941);
and U27113 (N_27113,N_26874,N_26739);
or U27114 (N_27114,N_26816,N_26995);
xor U27115 (N_27115,N_26668,N_26933);
xnor U27116 (N_27116,N_26714,N_26765);
xor U27117 (N_27117,N_26841,N_26973);
and U27118 (N_27118,N_26581,N_26908);
xnor U27119 (N_27119,N_26523,N_26963);
nand U27120 (N_27120,N_26738,N_26987);
or U27121 (N_27121,N_26660,N_26976);
xor U27122 (N_27122,N_26576,N_26578);
xnor U27123 (N_27123,N_26620,N_26916);
xnor U27124 (N_27124,N_26966,N_26930);
xnor U27125 (N_27125,N_26949,N_26656);
and U27126 (N_27126,N_26648,N_26990);
nand U27127 (N_27127,N_26989,N_26537);
and U27128 (N_27128,N_26502,N_26970);
nor U27129 (N_27129,N_26639,N_26641);
nor U27130 (N_27130,N_26698,N_26645);
xnor U27131 (N_27131,N_26670,N_26975);
xnor U27132 (N_27132,N_26882,N_26848);
nor U27133 (N_27133,N_26864,N_26925);
and U27134 (N_27134,N_26850,N_26810);
nand U27135 (N_27135,N_26605,N_26860);
nor U27136 (N_27136,N_26768,N_26780);
and U27137 (N_27137,N_26943,N_26644);
and U27138 (N_27138,N_26533,N_26664);
or U27139 (N_27139,N_26981,N_26735);
or U27140 (N_27140,N_26659,N_26718);
nor U27141 (N_27141,N_26633,N_26610);
nand U27142 (N_27142,N_26922,N_26535);
or U27143 (N_27143,N_26530,N_26824);
xor U27144 (N_27144,N_26665,N_26919);
nand U27145 (N_27145,N_26577,N_26510);
or U27146 (N_27146,N_26802,N_26599);
nor U27147 (N_27147,N_26960,N_26678);
xnor U27148 (N_27148,N_26903,N_26782);
nor U27149 (N_27149,N_26873,N_26712);
nor U27150 (N_27150,N_26829,N_26954);
nor U27151 (N_27151,N_26808,N_26926);
nand U27152 (N_27152,N_26547,N_26667);
xnor U27153 (N_27153,N_26881,N_26666);
nor U27154 (N_27154,N_26889,N_26837);
or U27155 (N_27155,N_26618,N_26635);
and U27156 (N_27156,N_26849,N_26968);
xor U27157 (N_27157,N_26819,N_26733);
nor U27158 (N_27158,N_26781,N_26619);
xnor U27159 (N_27159,N_26787,N_26680);
or U27160 (N_27160,N_26853,N_26684);
or U27161 (N_27161,N_26617,N_26843);
nor U27162 (N_27162,N_26595,N_26858);
nand U27163 (N_27163,N_26557,N_26825);
xor U27164 (N_27164,N_26993,N_26694);
or U27165 (N_27165,N_26662,N_26750);
or U27166 (N_27166,N_26504,N_26992);
nand U27167 (N_27167,N_26944,N_26833);
xor U27168 (N_27168,N_26505,N_26614);
and U27169 (N_27169,N_26910,N_26520);
nand U27170 (N_27170,N_26965,N_26734);
nor U27171 (N_27171,N_26705,N_26878);
nand U27172 (N_27172,N_26934,N_26744);
nand U27173 (N_27173,N_26755,N_26700);
and U27174 (N_27174,N_26647,N_26804);
and U27175 (N_27175,N_26880,N_26796);
nor U27176 (N_27176,N_26859,N_26982);
or U27177 (N_27177,N_26538,N_26741);
nor U27178 (N_27178,N_26514,N_26526);
xnor U27179 (N_27179,N_26911,N_26746);
and U27180 (N_27180,N_26658,N_26856);
and U27181 (N_27181,N_26554,N_26559);
nand U27182 (N_27182,N_26784,N_26766);
nand U27183 (N_27183,N_26630,N_26826);
xor U27184 (N_27184,N_26834,N_26892);
nand U27185 (N_27185,N_26994,N_26950);
or U27186 (N_27186,N_26701,N_26719);
or U27187 (N_27187,N_26985,N_26543);
xnor U27188 (N_27188,N_26748,N_26717);
nand U27189 (N_27189,N_26593,N_26795);
xor U27190 (N_27190,N_26952,N_26583);
nand U27191 (N_27191,N_26519,N_26671);
nand U27192 (N_27192,N_26632,N_26601);
and U27193 (N_27193,N_26602,N_26675);
nor U27194 (N_27194,N_26625,N_26962);
nand U27195 (N_27195,N_26937,N_26654);
nor U27196 (N_27196,N_26730,N_26566);
and U27197 (N_27197,N_26870,N_26921);
nand U27198 (N_27198,N_26726,N_26569);
xor U27199 (N_27199,N_26805,N_26603);
nand U27200 (N_27200,N_26570,N_26688);
xnor U27201 (N_27201,N_26556,N_26564);
nand U27202 (N_27202,N_26683,N_26600);
nor U27203 (N_27203,N_26799,N_26854);
xor U27204 (N_27204,N_26555,N_26649);
xnor U27205 (N_27205,N_26884,N_26958);
xor U27206 (N_27206,N_26901,N_26923);
nand U27207 (N_27207,N_26731,N_26663);
xnor U27208 (N_27208,N_26946,N_26999);
nor U27209 (N_27209,N_26596,N_26913);
xnor U27210 (N_27210,N_26762,N_26756);
or U27211 (N_27211,N_26844,N_26672);
or U27212 (N_27212,N_26587,N_26608);
or U27213 (N_27213,N_26820,N_26868);
nand U27214 (N_27214,N_26828,N_26681);
or U27215 (N_27215,N_26527,N_26821);
nand U27216 (N_27216,N_26876,N_26561);
or U27217 (N_27217,N_26807,N_26696);
nor U27218 (N_27218,N_26906,N_26904);
or U27219 (N_27219,N_26823,N_26938);
nand U27220 (N_27220,N_26932,N_26951);
xnor U27221 (N_27221,N_26789,N_26842);
and U27222 (N_27222,N_26661,N_26565);
or U27223 (N_27223,N_26743,N_26597);
xor U27224 (N_27224,N_26507,N_26753);
nand U27225 (N_27225,N_26657,N_26788);
and U27226 (N_27226,N_26560,N_26706);
nand U27227 (N_27227,N_26653,N_26915);
nor U27228 (N_27228,N_26875,N_26542);
and U27229 (N_27229,N_26980,N_26709);
or U27230 (N_27230,N_26594,N_26691);
and U27231 (N_27231,N_26983,N_26986);
nand U27232 (N_27232,N_26652,N_26515);
xor U27233 (N_27233,N_26695,N_26924);
nor U27234 (N_27234,N_26512,N_26574);
nor U27235 (N_27235,N_26754,N_26541);
nand U27236 (N_27236,N_26845,N_26872);
xor U27237 (N_27237,N_26540,N_26771);
nor U27238 (N_27238,N_26794,N_26612);
or U27239 (N_27239,N_26814,N_26511);
nand U27240 (N_27240,N_26887,N_26573);
or U27241 (N_27241,N_26550,N_26623);
nor U27242 (N_27242,N_26513,N_26900);
or U27243 (N_27243,N_26551,N_26759);
nor U27244 (N_27244,N_26775,N_26522);
xor U27245 (N_27245,N_26669,N_26957);
nand U27246 (N_27246,N_26500,N_26811);
or U27247 (N_27247,N_26839,N_26996);
nor U27248 (N_27248,N_26885,N_26776);
nand U27249 (N_27249,N_26732,N_26699);
or U27250 (N_27250,N_26870,N_26662);
xor U27251 (N_27251,N_26747,N_26823);
xnor U27252 (N_27252,N_26626,N_26836);
nor U27253 (N_27253,N_26856,N_26605);
nor U27254 (N_27254,N_26957,N_26573);
or U27255 (N_27255,N_26935,N_26966);
xor U27256 (N_27256,N_26951,N_26834);
and U27257 (N_27257,N_26590,N_26723);
xor U27258 (N_27258,N_26779,N_26961);
or U27259 (N_27259,N_26580,N_26629);
xnor U27260 (N_27260,N_26970,N_26934);
or U27261 (N_27261,N_26743,N_26673);
nor U27262 (N_27262,N_26892,N_26991);
or U27263 (N_27263,N_26928,N_26710);
nor U27264 (N_27264,N_26660,N_26771);
nand U27265 (N_27265,N_26842,N_26510);
nand U27266 (N_27266,N_26686,N_26826);
or U27267 (N_27267,N_26612,N_26523);
nand U27268 (N_27268,N_26964,N_26705);
or U27269 (N_27269,N_26869,N_26648);
xnor U27270 (N_27270,N_26741,N_26675);
and U27271 (N_27271,N_26547,N_26931);
xor U27272 (N_27272,N_26856,N_26912);
and U27273 (N_27273,N_26733,N_26708);
nand U27274 (N_27274,N_26795,N_26560);
nor U27275 (N_27275,N_26651,N_26535);
xor U27276 (N_27276,N_26827,N_26632);
and U27277 (N_27277,N_26846,N_26789);
and U27278 (N_27278,N_26748,N_26826);
nand U27279 (N_27279,N_26820,N_26610);
or U27280 (N_27280,N_26827,N_26862);
and U27281 (N_27281,N_26657,N_26964);
xnor U27282 (N_27282,N_26780,N_26996);
nor U27283 (N_27283,N_26807,N_26915);
nand U27284 (N_27284,N_26674,N_26682);
xnor U27285 (N_27285,N_26794,N_26712);
nand U27286 (N_27286,N_26643,N_26583);
nand U27287 (N_27287,N_26932,N_26571);
xor U27288 (N_27288,N_26643,N_26580);
nand U27289 (N_27289,N_26836,N_26816);
and U27290 (N_27290,N_26602,N_26927);
xnor U27291 (N_27291,N_26575,N_26835);
nor U27292 (N_27292,N_26885,N_26894);
nor U27293 (N_27293,N_26518,N_26588);
or U27294 (N_27294,N_26899,N_26696);
nor U27295 (N_27295,N_26907,N_26556);
and U27296 (N_27296,N_26971,N_26844);
and U27297 (N_27297,N_26844,N_26656);
xor U27298 (N_27298,N_26522,N_26518);
or U27299 (N_27299,N_26793,N_26786);
nand U27300 (N_27300,N_26516,N_26684);
nand U27301 (N_27301,N_26537,N_26781);
or U27302 (N_27302,N_26697,N_26734);
xnor U27303 (N_27303,N_26570,N_26919);
nand U27304 (N_27304,N_26897,N_26871);
or U27305 (N_27305,N_26519,N_26765);
and U27306 (N_27306,N_26992,N_26661);
nor U27307 (N_27307,N_26671,N_26597);
nor U27308 (N_27308,N_26868,N_26874);
nand U27309 (N_27309,N_26758,N_26912);
nor U27310 (N_27310,N_26828,N_26931);
nor U27311 (N_27311,N_26973,N_26844);
nor U27312 (N_27312,N_26667,N_26652);
xor U27313 (N_27313,N_26776,N_26954);
nand U27314 (N_27314,N_26921,N_26565);
xnor U27315 (N_27315,N_26695,N_26936);
nand U27316 (N_27316,N_26917,N_26988);
xnor U27317 (N_27317,N_26977,N_26970);
nor U27318 (N_27318,N_26599,N_26513);
or U27319 (N_27319,N_26715,N_26998);
xnor U27320 (N_27320,N_26627,N_26997);
nor U27321 (N_27321,N_26981,N_26508);
nand U27322 (N_27322,N_26689,N_26553);
or U27323 (N_27323,N_26811,N_26833);
nor U27324 (N_27324,N_26536,N_26604);
and U27325 (N_27325,N_26588,N_26880);
or U27326 (N_27326,N_26854,N_26607);
or U27327 (N_27327,N_26509,N_26554);
xor U27328 (N_27328,N_26630,N_26624);
nand U27329 (N_27329,N_26577,N_26545);
nand U27330 (N_27330,N_26532,N_26949);
nor U27331 (N_27331,N_26609,N_26664);
nor U27332 (N_27332,N_26603,N_26717);
or U27333 (N_27333,N_26850,N_26731);
or U27334 (N_27334,N_26643,N_26590);
or U27335 (N_27335,N_26545,N_26694);
or U27336 (N_27336,N_26937,N_26979);
nand U27337 (N_27337,N_26627,N_26977);
and U27338 (N_27338,N_26555,N_26821);
xnor U27339 (N_27339,N_26817,N_26973);
and U27340 (N_27340,N_26948,N_26564);
xor U27341 (N_27341,N_26671,N_26629);
or U27342 (N_27342,N_26889,N_26697);
and U27343 (N_27343,N_26521,N_26792);
xnor U27344 (N_27344,N_26666,N_26985);
and U27345 (N_27345,N_26809,N_26826);
nor U27346 (N_27346,N_26944,N_26509);
nand U27347 (N_27347,N_26565,N_26647);
xnor U27348 (N_27348,N_26889,N_26571);
and U27349 (N_27349,N_26987,N_26942);
or U27350 (N_27350,N_26521,N_26690);
xnor U27351 (N_27351,N_26789,N_26803);
or U27352 (N_27352,N_26950,N_26510);
nor U27353 (N_27353,N_26657,N_26806);
or U27354 (N_27354,N_26762,N_26675);
xnor U27355 (N_27355,N_26830,N_26737);
nor U27356 (N_27356,N_26883,N_26935);
nor U27357 (N_27357,N_26898,N_26815);
and U27358 (N_27358,N_26859,N_26848);
or U27359 (N_27359,N_26664,N_26765);
and U27360 (N_27360,N_26766,N_26817);
nand U27361 (N_27361,N_26683,N_26656);
xor U27362 (N_27362,N_26731,N_26685);
and U27363 (N_27363,N_26956,N_26775);
nor U27364 (N_27364,N_26923,N_26818);
and U27365 (N_27365,N_26673,N_26818);
or U27366 (N_27366,N_26750,N_26609);
nor U27367 (N_27367,N_26533,N_26809);
or U27368 (N_27368,N_26791,N_26805);
or U27369 (N_27369,N_26586,N_26697);
and U27370 (N_27370,N_26815,N_26606);
and U27371 (N_27371,N_26763,N_26706);
nor U27372 (N_27372,N_26979,N_26745);
nand U27373 (N_27373,N_26516,N_26610);
nor U27374 (N_27374,N_26696,N_26783);
or U27375 (N_27375,N_26726,N_26754);
and U27376 (N_27376,N_26872,N_26950);
nor U27377 (N_27377,N_26952,N_26690);
xnor U27378 (N_27378,N_26758,N_26898);
and U27379 (N_27379,N_26844,N_26993);
nand U27380 (N_27380,N_26702,N_26931);
or U27381 (N_27381,N_26764,N_26594);
nor U27382 (N_27382,N_26635,N_26960);
nand U27383 (N_27383,N_26978,N_26933);
xnor U27384 (N_27384,N_26970,N_26943);
nand U27385 (N_27385,N_26767,N_26941);
xor U27386 (N_27386,N_26913,N_26590);
xnor U27387 (N_27387,N_26548,N_26605);
or U27388 (N_27388,N_26836,N_26762);
nand U27389 (N_27389,N_26968,N_26648);
xor U27390 (N_27390,N_26749,N_26542);
or U27391 (N_27391,N_26690,N_26522);
nor U27392 (N_27392,N_26975,N_26875);
xnor U27393 (N_27393,N_26847,N_26766);
nand U27394 (N_27394,N_26838,N_26543);
or U27395 (N_27395,N_26614,N_26694);
and U27396 (N_27396,N_26638,N_26866);
nand U27397 (N_27397,N_26581,N_26871);
nand U27398 (N_27398,N_26891,N_26797);
nor U27399 (N_27399,N_26692,N_26879);
nand U27400 (N_27400,N_26506,N_26595);
or U27401 (N_27401,N_26618,N_26800);
or U27402 (N_27402,N_26625,N_26811);
and U27403 (N_27403,N_26875,N_26659);
nand U27404 (N_27404,N_26649,N_26757);
nor U27405 (N_27405,N_26810,N_26816);
and U27406 (N_27406,N_26687,N_26873);
nor U27407 (N_27407,N_26563,N_26661);
and U27408 (N_27408,N_26690,N_26987);
xnor U27409 (N_27409,N_26770,N_26700);
xnor U27410 (N_27410,N_26532,N_26728);
or U27411 (N_27411,N_26959,N_26652);
and U27412 (N_27412,N_26928,N_26851);
or U27413 (N_27413,N_26644,N_26858);
nor U27414 (N_27414,N_26820,N_26701);
or U27415 (N_27415,N_26851,N_26741);
nand U27416 (N_27416,N_26731,N_26772);
xor U27417 (N_27417,N_26535,N_26795);
and U27418 (N_27418,N_26745,N_26540);
nand U27419 (N_27419,N_26835,N_26767);
or U27420 (N_27420,N_26609,N_26753);
nor U27421 (N_27421,N_26694,N_26623);
and U27422 (N_27422,N_26605,N_26627);
nand U27423 (N_27423,N_26726,N_26983);
or U27424 (N_27424,N_26866,N_26710);
or U27425 (N_27425,N_26829,N_26836);
or U27426 (N_27426,N_26575,N_26756);
nor U27427 (N_27427,N_26998,N_26854);
nor U27428 (N_27428,N_26911,N_26689);
nand U27429 (N_27429,N_26682,N_26515);
and U27430 (N_27430,N_26632,N_26838);
or U27431 (N_27431,N_26854,N_26742);
nor U27432 (N_27432,N_26791,N_26660);
nor U27433 (N_27433,N_26973,N_26815);
nor U27434 (N_27434,N_26688,N_26524);
or U27435 (N_27435,N_26601,N_26778);
nand U27436 (N_27436,N_26997,N_26729);
or U27437 (N_27437,N_26687,N_26632);
or U27438 (N_27438,N_26815,N_26894);
xor U27439 (N_27439,N_26731,N_26630);
and U27440 (N_27440,N_26672,N_26979);
nand U27441 (N_27441,N_26748,N_26633);
xor U27442 (N_27442,N_26781,N_26933);
nor U27443 (N_27443,N_26967,N_26869);
or U27444 (N_27444,N_26908,N_26586);
nor U27445 (N_27445,N_26955,N_26547);
nor U27446 (N_27446,N_26814,N_26724);
and U27447 (N_27447,N_26524,N_26716);
nand U27448 (N_27448,N_26936,N_26952);
and U27449 (N_27449,N_26726,N_26962);
or U27450 (N_27450,N_26797,N_26998);
or U27451 (N_27451,N_26955,N_26818);
and U27452 (N_27452,N_26967,N_26899);
or U27453 (N_27453,N_26908,N_26642);
nor U27454 (N_27454,N_26759,N_26915);
nand U27455 (N_27455,N_26563,N_26916);
and U27456 (N_27456,N_26635,N_26781);
nand U27457 (N_27457,N_26634,N_26536);
and U27458 (N_27458,N_26930,N_26521);
and U27459 (N_27459,N_26843,N_26558);
nand U27460 (N_27460,N_26721,N_26872);
and U27461 (N_27461,N_26858,N_26660);
xor U27462 (N_27462,N_26849,N_26543);
and U27463 (N_27463,N_26836,N_26616);
or U27464 (N_27464,N_26742,N_26976);
or U27465 (N_27465,N_26818,N_26860);
nand U27466 (N_27466,N_26729,N_26722);
nand U27467 (N_27467,N_26526,N_26584);
nor U27468 (N_27468,N_26548,N_26922);
or U27469 (N_27469,N_26653,N_26815);
xor U27470 (N_27470,N_26614,N_26718);
and U27471 (N_27471,N_26646,N_26814);
nor U27472 (N_27472,N_26679,N_26774);
xnor U27473 (N_27473,N_26997,N_26935);
nand U27474 (N_27474,N_26540,N_26895);
or U27475 (N_27475,N_26743,N_26807);
xor U27476 (N_27476,N_26602,N_26611);
or U27477 (N_27477,N_26955,N_26746);
xnor U27478 (N_27478,N_26817,N_26805);
nand U27479 (N_27479,N_26711,N_26897);
nand U27480 (N_27480,N_26526,N_26850);
and U27481 (N_27481,N_26742,N_26683);
xnor U27482 (N_27482,N_26670,N_26708);
and U27483 (N_27483,N_26749,N_26639);
nor U27484 (N_27484,N_26820,N_26595);
nand U27485 (N_27485,N_26999,N_26524);
and U27486 (N_27486,N_26597,N_26850);
or U27487 (N_27487,N_26840,N_26740);
nand U27488 (N_27488,N_26673,N_26844);
or U27489 (N_27489,N_26806,N_26982);
nand U27490 (N_27490,N_26945,N_26762);
xor U27491 (N_27491,N_26958,N_26633);
nand U27492 (N_27492,N_26645,N_26953);
xor U27493 (N_27493,N_26650,N_26528);
nand U27494 (N_27494,N_26818,N_26814);
xnor U27495 (N_27495,N_26774,N_26839);
or U27496 (N_27496,N_26512,N_26812);
and U27497 (N_27497,N_26561,N_26813);
xor U27498 (N_27498,N_26583,N_26939);
or U27499 (N_27499,N_26651,N_26884);
and U27500 (N_27500,N_27394,N_27254);
nand U27501 (N_27501,N_27398,N_27061);
and U27502 (N_27502,N_27341,N_27369);
or U27503 (N_27503,N_27024,N_27452);
and U27504 (N_27504,N_27118,N_27349);
or U27505 (N_27505,N_27071,N_27330);
nor U27506 (N_27506,N_27206,N_27337);
xor U27507 (N_27507,N_27161,N_27142);
nor U27508 (N_27508,N_27209,N_27011);
and U27509 (N_27509,N_27256,N_27151);
xnor U27510 (N_27510,N_27252,N_27305);
xnor U27511 (N_27511,N_27304,N_27019);
nor U27512 (N_27512,N_27469,N_27180);
and U27513 (N_27513,N_27390,N_27288);
and U27514 (N_27514,N_27395,N_27350);
and U27515 (N_27515,N_27086,N_27445);
and U27516 (N_27516,N_27447,N_27217);
xnor U27517 (N_27517,N_27176,N_27268);
nor U27518 (N_27518,N_27257,N_27426);
nor U27519 (N_27519,N_27290,N_27249);
or U27520 (N_27520,N_27476,N_27236);
or U27521 (N_27521,N_27121,N_27187);
and U27522 (N_27522,N_27382,N_27001);
nor U27523 (N_27523,N_27059,N_27432);
nor U27524 (N_27524,N_27181,N_27040);
nand U27525 (N_27525,N_27296,N_27072);
nor U27526 (N_27526,N_27427,N_27492);
nor U27527 (N_27527,N_27074,N_27352);
nor U27528 (N_27528,N_27013,N_27131);
nor U27529 (N_27529,N_27092,N_27077);
nand U27530 (N_27530,N_27424,N_27220);
or U27531 (N_27531,N_27091,N_27234);
nand U27532 (N_27532,N_27282,N_27250);
or U27533 (N_27533,N_27251,N_27497);
xnor U27534 (N_27534,N_27300,N_27479);
and U27535 (N_27535,N_27309,N_27088);
and U27536 (N_27536,N_27443,N_27458);
or U27537 (N_27537,N_27124,N_27127);
xnor U27538 (N_27538,N_27007,N_27293);
nor U27539 (N_27539,N_27351,N_27302);
xnor U27540 (N_27540,N_27402,N_27363);
nor U27541 (N_27541,N_27025,N_27437);
and U27542 (N_27542,N_27055,N_27473);
nand U27543 (N_27543,N_27267,N_27143);
xor U27544 (N_27544,N_27283,N_27232);
nand U27545 (N_27545,N_27237,N_27372);
or U27546 (N_27546,N_27201,N_27393);
nand U27547 (N_27547,N_27397,N_27155);
xnor U27548 (N_27548,N_27245,N_27406);
nor U27549 (N_27549,N_27488,N_27020);
nand U27550 (N_27550,N_27174,N_27238);
nor U27551 (N_27551,N_27422,N_27491);
and U27552 (N_27552,N_27333,N_27311);
nor U27553 (N_27553,N_27212,N_27216);
nand U27554 (N_27554,N_27291,N_27226);
and U27555 (N_27555,N_27178,N_27042);
nand U27556 (N_27556,N_27389,N_27494);
xor U27557 (N_27557,N_27010,N_27002);
xor U27558 (N_27558,N_27246,N_27213);
or U27559 (N_27559,N_27258,N_27281);
xnor U27560 (N_27560,N_27158,N_27459);
nand U27561 (N_27561,N_27248,N_27436);
and U27562 (N_27562,N_27493,N_27327);
nor U27563 (N_27563,N_27353,N_27414);
xnor U27564 (N_27564,N_27123,N_27218);
xnor U27565 (N_27565,N_27457,N_27316);
and U27566 (N_27566,N_27243,N_27312);
or U27567 (N_27567,N_27244,N_27358);
or U27568 (N_27568,N_27100,N_27102);
and U27569 (N_27569,N_27381,N_27044);
or U27570 (N_27570,N_27418,N_27294);
and U27571 (N_27571,N_27379,N_27346);
nand U27572 (N_27572,N_27191,N_27292);
xor U27573 (N_27573,N_27079,N_27430);
and U27574 (N_27574,N_27221,N_27108);
and U27575 (N_27575,N_27183,N_27451);
and U27576 (N_27576,N_27377,N_27429);
nor U27577 (N_27577,N_27462,N_27223);
and U27578 (N_27578,N_27057,N_27295);
and U27579 (N_27579,N_27126,N_27310);
nor U27580 (N_27580,N_27075,N_27365);
xnor U27581 (N_27581,N_27166,N_27169);
xnor U27582 (N_27582,N_27374,N_27313);
and U27583 (N_27583,N_27134,N_27415);
or U27584 (N_27584,N_27208,N_27242);
and U27585 (N_27585,N_27081,N_27043);
xor U27586 (N_27586,N_27205,N_27317);
and U27587 (N_27587,N_27391,N_27315);
nand U27588 (N_27588,N_27229,N_27064);
nor U27589 (N_27589,N_27222,N_27483);
and U27590 (N_27590,N_27210,N_27356);
nand U27591 (N_27591,N_27199,N_27320);
nor U27592 (N_27592,N_27386,N_27160);
xor U27593 (N_27593,N_27195,N_27113);
xnor U27594 (N_27594,N_27371,N_27400);
nor U27595 (N_27595,N_27408,N_27261);
nand U27596 (N_27596,N_27095,N_27197);
nor U27597 (N_27597,N_27224,N_27388);
and U27598 (N_27598,N_27384,N_27110);
and U27599 (N_27599,N_27307,N_27101);
xor U27600 (N_27600,N_27182,N_27004);
nand U27601 (N_27601,N_27287,N_27136);
nand U27602 (N_27602,N_27423,N_27046);
xor U27603 (N_27603,N_27050,N_27318);
nor U27604 (N_27604,N_27409,N_27319);
or U27605 (N_27605,N_27485,N_27284);
xnor U27606 (N_27606,N_27023,N_27495);
xor U27607 (N_27607,N_27240,N_27165);
or U27608 (N_27608,N_27027,N_27198);
nor U27609 (N_27609,N_27119,N_27419);
or U27610 (N_27610,N_27093,N_27135);
and U27611 (N_27611,N_27463,N_27339);
or U27612 (N_27612,N_27401,N_27157);
or U27613 (N_27613,N_27475,N_27247);
or U27614 (N_27614,N_27367,N_27303);
nand U27615 (N_27615,N_27299,N_27331);
and U27616 (N_27616,N_27440,N_27122);
or U27617 (N_27617,N_27233,N_27227);
nand U27618 (N_27618,N_27487,N_27308);
or U27619 (N_27619,N_27029,N_27453);
or U27620 (N_27620,N_27163,N_27450);
xor U27621 (N_27621,N_27144,N_27276);
and U27622 (N_27622,N_27175,N_27104);
xnor U27623 (N_27623,N_27412,N_27006);
nand U27624 (N_27624,N_27364,N_27321);
and U27625 (N_27625,N_27411,N_27008);
nand U27626 (N_27626,N_27038,N_27439);
and U27627 (N_27627,N_27060,N_27026);
nand U27628 (N_27628,N_27062,N_27015);
or U27629 (N_27629,N_27273,N_27404);
and U27630 (N_27630,N_27066,N_27152);
nor U27631 (N_27631,N_27137,N_27156);
nor U27632 (N_27632,N_27428,N_27239);
nand U27633 (N_27633,N_27482,N_27489);
and U27634 (N_27634,N_27005,N_27380);
nor U27635 (N_27635,N_27410,N_27076);
or U27636 (N_27636,N_27065,N_27354);
and U27637 (N_27637,N_27202,N_27070);
nor U27638 (N_27638,N_27200,N_27097);
or U27639 (N_27639,N_27347,N_27470);
nor U27640 (N_27640,N_27107,N_27396);
xnor U27641 (N_27641,N_27499,N_27052);
nor U27642 (N_27642,N_27279,N_27405);
and U27643 (N_27643,N_27150,N_27326);
xor U27644 (N_27644,N_27269,N_27085);
or U27645 (N_27645,N_27253,N_27037);
xnor U27646 (N_27646,N_27480,N_27344);
nand U27647 (N_27647,N_27285,N_27056);
and U27648 (N_27648,N_27460,N_27231);
nand U27649 (N_27649,N_27045,N_27106);
xnor U27650 (N_27650,N_27022,N_27036);
or U27651 (N_27651,N_27177,N_27105);
nand U27652 (N_27652,N_27474,N_27498);
xnor U27653 (N_27653,N_27111,N_27442);
and U27654 (N_27654,N_27449,N_27096);
xnor U27655 (N_27655,N_27342,N_27266);
and U27656 (N_27656,N_27324,N_27017);
nor U27657 (N_27657,N_27031,N_27129);
xnor U27658 (N_27658,N_27009,N_27345);
xor U27659 (N_27659,N_27435,N_27145);
and U27660 (N_27660,N_27286,N_27306);
nand U27661 (N_27661,N_27271,N_27454);
and U27662 (N_27662,N_27047,N_27467);
xnor U27663 (N_27663,N_27033,N_27069);
nor U27664 (N_27664,N_27048,N_27378);
or U27665 (N_27665,N_27193,N_27192);
nor U27666 (N_27666,N_27018,N_27496);
and U27667 (N_27667,N_27301,N_27416);
or U27668 (N_27668,N_27032,N_27051);
nor U27669 (N_27669,N_27203,N_27194);
nand U27670 (N_27670,N_27265,N_27263);
nand U27671 (N_27671,N_27366,N_27219);
or U27672 (N_27672,N_27444,N_27434);
nor U27673 (N_27673,N_27000,N_27099);
nand U27674 (N_27674,N_27185,N_27385);
and U27675 (N_27675,N_27413,N_27146);
or U27676 (N_27676,N_27448,N_27370);
and U27677 (N_27677,N_27215,N_27139);
or U27678 (N_27678,N_27278,N_27103);
and U27679 (N_27679,N_27360,N_27259);
and U27680 (N_27680,N_27357,N_27468);
xor U27681 (N_27681,N_27179,N_27204);
xnor U27682 (N_27682,N_27117,N_27417);
or U27683 (N_27683,N_27115,N_27164);
and U27684 (N_27684,N_27338,N_27477);
xnor U27685 (N_27685,N_27264,N_27186);
or U27686 (N_27686,N_27325,N_27464);
and U27687 (N_27687,N_27270,N_27132);
or U27688 (N_27688,N_27171,N_27128);
or U27689 (N_27689,N_27335,N_27478);
nor U27690 (N_27690,N_27328,N_27109);
xor U27691 (N_27691,N_27016,N_27277);
nand U27692 (N_27692,N_27188,N_27012);
nand U27693 (N_27693,N_27272,N_27087);
nand U27694 (N_27694,N_27438,N_27420);
nor U27695 (N_27695,N_27207,N_27073);
xnor U27696 (N_27696,N_27130,N_27159);
and U27697 (N_27697,N_27433,N_27230);
or U27698 (N_27698,N_27116,N_27035);
and U27699 (N_27699,N_27082,N_27446);
or U27700 (N_27700,N_27089,N_27332);
and U27701 (N_27701,N_27068,N_27336);
and U27702 (N_27702,N_27375,N_27228);
xor U27703 (N_27703,N_27484,N_27399);
and U27704 (N_27704,N_27297,N_27425);
nand U27705 (N_27705,N_27274,N_27211);
xnor U27706 (N_27706,N_27376,N_27141);
nor U27707 (N_27707,N_27368,N_27235);
nor U27708 (N_27708,N_27334,N_27340);
xor U27709 (N_27709,N_27214,N_27080);
nor U27710 (N_27710,N_27098,N_27361);
or U27711 (N_27711,N_27472,N_27063);
nand U27712 (N_27712,N_27456,N_27486);
nand U27713 (N_27713,N_27275,N_27153);
xor U27714 (N_27714,N_27348,N_27373);
nor U27715 (N_27715,N_27162,N_27041);
nor U27716 (N_27716,N_27125,N_27289);
or U27717 (N_27717,N_27021,N_27039);
nand U27718 (N_27718,N_27329,N_27090);
nand U27719 (N_27719,N_27461,N_27225);
and U27720 (N_27720,N_27314,N_27189);
nor U27721 (N_27721,N_27322,N_27260);
xor U27722 (N_27722,N_27058,N_27421);
and U27723 (N_27723,N_27078,N_27392);
and U27724 (N_27724,N_27481,N_27034);
or U27725 (N_27725,N_27030,N_27383);
or U27726 (N_27726,N_27407,N_27184);
or U27727 (N_27727,N_27148,N_27465);
and U27728 (N_27728,N_27343,N_27147);
and U27729 (N_27729,N_27359,N_27431);
or U27730 (N_27730,N_27094,N_27262);
nor U27731 (N_27731,N_27466,N_27355);
and U27732 (N_27732,N_27003,N_27170);
and U27733 (N_27733,N_27323,N_27133);
nor U27734 (N_27734,N_27387,N_27471);
and U27735 (N_27735,N_27083,N_27172);
and U27736 (N_27736,N_27138,N_27255);
nor U27737 (N_27737,N_27455,N_27190);
nor U27738 (N_27738,N_27114,N_27120);
xor U27739 (N_27739,N_27140,N_27084);
or U27740 (N_27740,N_27168,N_27154);
nand U27741 (N_27741,N_27173,N_27053);
nor U27742 (N_27742,N_27149,N_27028);
xor U27743 (N_27743,N_27241,N_27196);
nand U27744 (N_27744,N_27403,N_27298);
xnor U27745 (N_27745,N_27167,N_27067);
or U27746 (N_27746,N_27280,N_27441);
and U27747 (N_27747,N_27362,N_27014);
nand U27748 (N_27748,N_27054,N_27049);
nand U27749 (N_27749,N_27112,N_27490);
or U27750 (N_27750,N_27314,N_27069);
nand U27751 (N_27751,N_27411,N_27106);
or U27752 (N_27752,N_27458,N_27065);
nand U27753 (N_27753,N_27268,N_27427);
or U27754 (N_27754,N_27230,N_27137);
nand U27755 (N_27755,N_27403,N_27055);
nor U27756 (N_27756,N_27104,N_27112);
or U27757 (N_27757,N_27364,N_27492);
and U27758 (N_27758,N_27162,N_27103);
or U27759 (N_27759,N_27384,N_27074);
nand U27760 (N_27760,N_27372,N_27111);
or U27761 (N_27761,N_27330,N_27303);
nand U27762 (N_27762,N_27430,N_27467);
or U27763 (N_27763,N_27197,N_27200);
xor U27764 (N_27764,N_27017,N_27498);
and U27765 (N_27765,N_27406,N_27014);
nor U27766 (N_27766,N_27079,N_27166);
or U27767 (N_27767,N_27073,N_27165);
nor U27768 (N_27768,N_27113,N_27030);
nand U27769 (N_27769,N_27413,N_27448);
and U27770 (N_27770,N_27189,N_27113);
nand U27771 (N_27771,N_27309,N_27174);
nand U27772 (N_27772,N_27204,N_27060);
nor U27773 (N_27773,N_27470,N_27415);
or U27774 (N_27774,N_27138,N_27166);
nor U27775 (N_27775,N_27437,N_27348);
or U27776 (N_27776,N_27325,N_27115);
nor U27777 (N_27777,N_27273,N_27161);
or U27778 (N_27778,N_27208,N_27436);
or U27779 (N_27779,N_27376,N_27373);
or U27780 (N_27780,N_27240,N_27035);
or U27781 (N_27781,N_27227,N_27376);
xor U27782 (N_27782,N_27192,N_27070);
nand U27783 (N_27783,N_27433,N_27292);
and U27784 (N_27784,N_27144,N_27352);
xnor U27785 (N_27785,N_27419,N_27422);
nor U27786 (N_27786,N_27081,N_27430);
and U27787 (N_27787,N_27306,N_27315);
xor U27788 (N_27788,N_27117,N_27238);
nand U27789 (N_27789,N_27408,N_27105);
nor U27790 (N_27790,N_27284,N_27467);
or U27791 (N_27791,N_27095,N_27421);
and U27792 (N_27792,N_27357,N_27250);
nand U27793 (N_27793,N_27211,N_27487);
or U27794 (N_27794,N_27103,N_27378);
and U27795 (N_27795,N_27363,N_27376);
xor U27796 (N_27796,N_27154,N_27018);
nor U27797 (N_27797,N_27155,N_27437);
nand U27798 (N_27798,N_27467,N_27031);
and U27799 (N_27799,N_27473,N_27436);
and U27800 (N_27800,N_27446,N_27003);
and U27801 (N_27801,N_27387,N_27099);
nand U27802 (N_27802,N_27386,N_27105);
and U27803 (N_27803,N_27032,N_27445);
and U27804 (N_27804,N_27278,N_27148);
nor U27805 (N_27805,N_27480,N_27277);
xnor U27806 (N_27806,N_27342,N_27041);
nand U27807 (N_27807,N_27476,N_27098);
nand U27808 (N_27808,N_27229,N_27012);
nand U27809 (N_27809,N_27292,N_27480);
nor U27810 (N_27810,N_27154,N_27099);
or U27811 (N_27811,N_27045,N_27016);
xnor U27812 (N_27812,N_27088,N_27430);
or U27813 (N_27813,N_27429,N_27352);
nand U27814 (N_27814,N_27187,N_27044);
or U27815 (N_27815,N_27491,N_27052);
or U27816 (N_27816,N_27141,N_27469);
xnor U27817 (N_27817,N_27002,N_27345);
nor U27818 (N_27818,N_27067,N_27433);
nand U27819 (N_27819,N_27488,N_27201);
nor U27820 (N_27820,N_27440,N_27194);
and U27821 (N_27821,N_27050,N_27280);
nand U27822 (N_27822,N_27497,N_27074);
or U27823 (N_27823,N_27244,N_27483);
xnor U27824 (N_27824,N_27309,N_27220);
nor U27825 (N_27825,N_27292,N_27346);
xor U27826 (N_27826,N_27060,N_27281);
and U27827 (N_27827,N_27048,N_27415);
nor U27828 (N_27828,N_27012,N_27038);
nor U27829 (N_27829,N_27340,N_27331);
xnor U27830 (N_27830,N_27207,N_27164);
nor U27831 (N_27831,N_27154,N_27256);
xor U27832 (N_27832,N_27309,N_27107);
or U27833 (N_27833,N_27304,N_27008);
and U27834 (N_27834,N_27050,N_27188);
xnor U27835 (N_27835,N_27407,N_27263);
or U27836 (N_27836,N_27336,N_27349);
nor U27837 (N_27837,N_27346,N_27136);
nand U27838 (N_27838,N_27010,N_27213);
xnor U27839 (N_27839,N_27497,N_27441);
and U27840 (N_27840,N_27119,N_27070);
nor U27841 (N_27841,N_27376,N_27269);
nor U27842 (N_27842,N_27429,N_27169);
nor U27843 (N_27843,N_27381,N_27054);
xor U27844 (N_27844,N_27416,N_27319);
nor U27845 (N_27845,N_27437,N_27139);
nand U27846 (N_27846,N_27261,N_27394);
and U27847 (N_27847,N_27193,N_27423);
and U27848 (N_27848,N_27323,N_27068);
nor U27849 (N_27849,N_27389,N_27099);
and U27850 (N_27850,N_27281,N_27205);
or U27851 (N_27851,N_27047,N_27249);
nor U27852 (N_27852,N_27238,N_27334);
xor U27853 (N_27853,N_27145,N_27027);
or U27854 (N_27854,N_27024,N_27119);
and U27855 (N_27855,N_27404,N_27368);
and U27856 (N_27856,N_27213,N_27493);
nor U27857 (N_27857,N_27461,N_27470);
nor U27858 (N_27858,N_27325,N_27226);
xnor U27859 (N_27859,N_27104,N_27436);
xor U27860 (N_27860,N_27408,N_27445);
and U27861 (N_27861,N_27433,N_27380);
and U27862 (N_27862,N_27433,N_27478);
xnor U27863 (N_27863,N_27063,N_27212);
nor U27864 (N_27864,N_27338,N_27054);
nand U27865 (N_27865,N_27008,N_27005);
nor U27866 (N_27866,N_27398,N_27199);
and U27867 (N_27867,N_27042,N_27327);
xor U27868 (N_27868,N_27435,N_27442);
nand U27869 (N_27869,N_27160,N_27120);
nand U27870 (N_27870,N_27492,N_27395);
xnor U27871 (N_27871,N_27453,N_27381);
xnor U27872 (N_27872,N_27455,N_27175);
nor U27873 (N_27873,N_27214,N_27348);
or U27874 (N_27874,N_27249,N_27206);
and U27875 (N_27875,N_27147,N_27152);
nor U27876 (N_27876,N_27419,N_27042);
or U27877 (N_27877,N_27173,N_27122);
or U27878 (N_27878,N_27182,N_27019);
and U27879 (N_27879,N_27213,N_27309);
xnor U27880 (N_27880,N_27107,N_27271);
nor U27881 (N_27881,N_27221,N_27148);
xor U27882 (N_27882,N_27422,N_27204);
and U27883 (N_27883,N_27438,N_27201);
xor U27884 (N_27884,N_27383,N_27097);
or U27885 (N_27885,N_27343,N_27470);
and U27886 (N_27886,N_27403,N_27139);
or U27887 (N_27887,N_27244,N_27350);
nand U27888 (N_27888,N_27480,N_27346);
nor U27889 (N_27889,N_27076,N_27367);
and U27890 (N_27890,N_27424,N_27412);
or U27891 (N_27891,N_27386,N_27115);
nand U27892 (N_27892,N_27263,N_27460);
xnor U27893 (N_27893,N_27065,N_27479);
nand U27894 (N_27894,N_27149,N_27078);
or U27895 (N_27895,N_27406,N_27065);
nand U27896 (N_27896,N_27116,N_27352);
nor U27897 (N_27897,N_27082,N_27292);
nand U27898 (N_27898,N_27468,N_27270);
and U27899 (N_27899,N_27415,N_27055);
xnor U27900 (N_27900,N_27112,N_27124);
or U27901 (N_27901,N_27067,N_27088);
nand U27902 (N_27902,N_27474,N_27166);
nor U27903 (N_27903,N_27328,N_27007);
or U27904 (N_27904,N_27371,N_27487);
xor U27905 (N_27905,N_27278,N_27280);
and U27906 (N_27906,N_27479,N_27254);
and U27907 (N_27907,N_27493,N_27153);
and U27908 (N_27908,N_27152,N_27091);
xor U27909 (N_27909,N_27256,N_27456);
xor U27910 (N_27910,N_27479,N_27218);
nor U27911 (N_27911,N_27250,N_27050);
or U27912 (N_27912,N_27343,N_27400);
xnor U27913 (N_27913,N_27428,N_27269);
nor U27914 (N_27914,N_27439,N_27133);
and U27915 (N_27915,N_27122,N_27451);
xor U27916 (N_27916,N_27199,N_27015);
nor U27917 (N_27917,N_27182,N_27370);
and U27918 (N_27918,N_27308,N_27033);
or U27919 (N_27919,N_27061,N_27308);
and U27920 (N_27920,N_27094,N_27499);
xor U27921 (N_27921,N_27136,N_27443);
or U27922 (N_27922,N_27360,N_27010);
nor U27923 (N_27923,N_27387,N_27458);
and U27924 (N_27924,N_27304,N_27404);
nor U27925 (N_27925,N_27093,N_27398);
xor U27926 (N_27926,N_27296,N_27025);
or U27927 (N_27927,N_27395,N_27072);
and U27928 (N_27928,N_27365,N_27342);
nor U27929 (N_27929,N_27097,N_27406);
xnor U27930 (N_27930,N_27091,N_27252);
xor U27931 (N_27931,N_27136,N_27378);
nor U27932 (N_27932,N_27190,N_27481);
nor U27933 (N_27933,N_27351,N_27062);
or U27934 (N_27934,N_27107,N_27240);
or U27935 (N_27935,N_27396,N_27253);
nand U27936 (N_27936,N_27272,N_27432);
nor U27937 (N_27937,N_27121,N_27310);
or U27938 (N_27938,N_27218,N_27332);
and U27939 (N_27939,N_27222,N_27374);
xor U27940 (N_27940,N_27148,N_27285);
and U27941 (N_27941,N_27255,N_27050);
or U27942 (N_27942,N_27383,N_27079);
and U27943 (N_27943,N_27072,N_27289);
nand U27944 (N_27944,N_27460,N_27211);
nand U27945 (N_27945,N_27194,N_27004);
nor U27946 (N_27946,N_27164,N_27348);
xor U27947 (N_27947,N_27447,N_27024);
or U27948 (N_27948,N_27254,N_27478);
nor U27949 (N_27949,N_27066,N_27493);
xor U27950 (N_27950,N_27158,N_27099);
nor U27951 (N_27951,N_27114,N_27401);
and U27952 (N_27952,N_27211,N_27235);
and U27953 (N_27953,N_27192,N_27075);
nand U27954 (N_27954,N_27121,N_27188);
nor U27955 (N_27955,N_27356,N_27024);
nor U27956 (N_27956,N_27080,N_27250);
nand U27957 (N_27957,N_27255,N_27471);
nor U27958 (N_27958,N_27103,N_27392);
nor U27959 (N_27959,N_27161,N_27187);
xor U27960 (N_27960,N_27403,N_27135);
nor U27961 (N_27961,N_27270,N_27014);
nand U27962 (N_27962,N_27261,N_27165);
or U27963 (N_27963,N_27404,N_27347);
xnor U27964 (N_27964,N_27404,N_27172);
nor U27965 (N_27965,N_27477,N_27403);
and U27966 (N_27966,N_27060,N_27383);
and U27967 (N_27967,N_27244,N_27471);
nor U27968 (N_27968,N_27486,N_27428);
xnor U27969 (N_27969,N_27462,N_27352);
nand U27970 (N_27970,N_27041,N_27147);
nor U27971 (N_27971,N_27028,N_27196);
nor U27972 (N_27972,N_27026,N_27409);
xor U27973 (N_27973,N_27139,N_27052);
or U27974 (N_27974,N_27248,N_27378);
nand U27975 (N_27975,N_27197,N_27213);
xnor U27976 (N_27976,N_27014,N_27360);
xor U27977 (N_27977,N_27304,N_27261);
or U27978 (N_27978,N_27104,N_27156);
or U27979 (N_27979,N_27090,N_27323);
nor U27980 (N_27980,N_27347,N_27065);
or U27981 (N_27981,N_27301,N_27052);
or U27982 (N_27982,N_27292,N_27112);
nand U27983 (N_27983,N_27199,N_27343);
xor U27984 (N_27984,N_27090,N_27317);
xor U27985 (N_27985,N_27060,N_27443);
nor U27986 (N_27986,N_27083,N_27110);
and U27987 (N_27987,N_27336,N_27180);
and U27988 (N_27988,N_27035,N_27251);
and U27989 (N_27989,N_27267,N_27318);
or U27990 (N_27990,N_27415,N_27195);
xnor U27991 (N_27991,N_27199,N_27149);
or U27992 (N_27992,N_27212,N_27100);
nand U27993 (N_27993,N_27038,N_27473);
nand U27994 (N_27994,N_27434,N_27213);
or U27995 (N_27995,N_27007,N_27381);
or U27996 (N_27996,N_27251,N_27412);
and U27997 (N_27997,N_27104,N_27181);
nand U27998 (N_27998,N_27037,N_27373);
xnor U27999 (N_27999,N_27034,N_27118);
nor U28000 (N_28000,N_27944,N_27751);
xor U28001 (N_28001,N_27572,N_27966);
nor U28002 (N_28002,N_27673,N_27921);
or U28003 (N_28003,N_27747,N_27840);
nor U28004 (N_28004,N_27817,N_27524);
or U28005 (N_28005,N_27909,N_27919);
nor U28006 (N_28006,N_27641,N_27976);
and U28007 (N_28007,N_27750,N_27502);
or U28008 (N_28008,N_27813,N_27748);
and U28009 (N_28009,N_27636,N_27684);
nor U28010 (N_28010,N_27903,N_27827);
and U28011 (N_28011,N_27836,N_27563);
or U28012 (N_28012,N_27870,N_27842);
or U28013 (N_28013,N_27878,N_27717);
xor U28014 (N_28014,N_27759,N_27805);
or U28015 (N_28015,N_27676,N_27807);
and U28016 (N_28016,N_27999,N_27943);
or U28017 (N_28017,N_27588,N_27810);
xnor U28018 (N_28018,N_27961,N_27783);
or U28019 (N_28019,N_27512,N_27906);
and U28020 (N_28020,N_27890,N_27616);
and U28021 (N_28021,N_27733,N_27874);
xor U28022 (N_28022,N_27738,N_27682);
xor U28023 (N_28023,N_27631,N_27758);
or U28024 (N_28024,N_27736,N_27774);
and U28025 (N_28025,N_27649,N_27568);
or U28026 (N_28026,N_27958,N_27861);
nor U28027 (N_28027,N_27669,N_27674);
or U28028 (N_28028,N_27993,N_27691);
nand U28029 (N_28029,N_27938,N_27911);
xnor U28030 (N_28030,N_27700,N_27784);
xor U28031 (N_28031,N_27963,N_27528);
nand U28032 (N_28032,N_27642,N_27735);
or U28033 (N_28033,N_27865,N_27532);
nor U28034 (N_28034,N_27744,N_27816);
and U28035 (N_28035,N_27896,N_27908);
or U28036 (N_28036,N_27686,N_27949);
and U28037 (N_28037,N_27771,N_27763);
or U28038 (N_28038,N_27651,N_27811);
and U28039 (N_28039,N_27534,N_27786);
nor U28040 (N_28040,N_27756,N_27897);
or U28041 (N_28041,N_27607,N_27606);
nand U28042 (N_28042,N_27787,N_27598);
or U28043 (N_28043,N_27515,N_27710);
or U28044 (N_28044,N_27561,N_27765);
xor U28045 (N_28045,N_27715,N_27675);
nor U28046 (N_28046,N_27581,N_27677);
nor U28047 (N_28047,N_27804,N_27867);
and U28048 (N_28048,N_27950,N_27752);
or U28049 (N_28049,N_27764,N_27955);
nor U28050 (N_28050,N_27998,N_27977);
xor U28051 (N_28051,N_27728,N_27894);
or U28052 (N_28052,N_27547,N_27799);
nor U28053 (N_28053,N_27823,N_27514);
or U28054 (N_28054,N_27671,N_27615);
xor U28055 (N_28055,N_27688,N_27910);
or U28056 (N_28056,N_27645,N_27806);
xor U28057 (N_28057,N_27725,N_27790);
nor U28058 (N_28058,N_27826,N_27838);
and U28059 (N_28059,N_27730,N_27656);
and U28060 (N_28060,N_27685,N_27754);
or U28061 (N_28061,N_27757,N_27780);
or U28062 (N_28062,N_27926,N_27550);
or U28063 (N_28063,N_27599,N_27832);
or U28064 (N_28064,N_27791,N_27925);
xnor U28065 (N_28065,N_27716,N_27628);
nor U28066 (N_28066,N_27558,N_27866);
or U28067 (N_28067,N_27985,N_27626);
or U28068 (N_28068,N_27907,N_27658);
or U28069 (N_28069,N_27697,N_27883);
nand U28070 (N_28070,N_27574,N_27970);
or U28071 (N_28071,N_27851,N_27794);
nor U28072 (N_28072,N_27683,N_27647);
nor U28073 (N_28073,N_27644,N_27973);
and U28074 (N_28074,N_27650,N_27583);
nand U28075 (N_28075,N_27538,N_27672);
xnor U28076 (N_28076,N_27662,N_27916);
or U28077 (N_28077,N_27777,N_27749);
or U28078 (N_28078,N_27539,N_27990);
xnor U28079 (N_28079,N_27796,N_27664);
and U28080 (N_28080,N_27601,N_27776);
or U28081 (N_28081,N_27580,N_27872);
or U28082 (N_28082,N_27726,N_27869);
or U28083 (N_28083,N_27595,N_27564);
or U28084 (N_28084,N_27881,N_27629);
xnor U28085 (N_28085,N_27828,N_27948);
nor U28086 (N_28086,N_27830,N_27873);
or U28087 (N_28087,N_27613,N_27722);
nand U28088 (N_28088,N_27905,N_27510);
nor U28089 (N_28089,N_27996,N_27737);
xor U28090 (N_28090,N_27923,N_27654);
or U28091 (N_28091,N_27969,N_27850);
or U28092 (N_28092,N_27960,N_27552);
nor U28093 (N_28093,N_27681,N_27541);
or U28094 (N_28094,N_27693,N_27505);
and U28095 (N_28095,N_27600,N_27788);
nand U28096 (N_28096,N_27935,N_27729);
nor U28097 (N_28097,N_27959,N_27648);
xnor U28098 (N_28098,N_27618,N_27871);
nand U28099 (N_28099,N_27741,N_27770);
nand U28100 (N_28100,N_27971,N_27530);
and U28101 (N_28101,N_27667,N_27980);
and U28102 (N_28102,N_27690,N_27655);
and U28103 (N_28103,N_27540,N_27834);
or U28104 (N_28104,N_27582,N_27608);
nor U28105 (N_28105,N_27900,N_27974);
xnor U28106 (N_28106,N_27824,N_27852);
nor U28107 (N_28107,N_27553,N_27500);
nor U28108 (N_28108,N_27863,N_27934);
xor U28109 (N_28109,N_27868,N_27507);
and U28110 (N_28110,N_27696,N_27732);
or U28111 (N_28111,N_27533,N_27857);
or U28112 (N_28112,N_27860,N_27835);
xnor U28113 (N_28113,N_27609,N_27979);
nand U28114 (N_28114,N_27933,N_27593);
nand U28115 (N_28115,N_27854,N_27922);
and U28116 (N_28116,N_27594,N_27603);
and U28117 (N_28117,N_27818,N_27635);
nor U28118 (N_28118,N_27508,N_27767);
nor U28119 (N_28119,N_27839,N_27537);
or U28120 (N_28120,N_27724,N_27841);
nand U28121 (N_28121,N_27779,N_27521);
xnor U28122 (N_28122,N_27978,N_27984);
xnor U28123 (N_28123,N_27927,N_27556);
or U28124 (N_28124,N_27638,N_27701);
or U28125 (N_28125,N_27511,N_27740);
and U28126 (N_28126,N_27578,N_27800);
or U28127 (N_28127,N_27972,N_27663);
and U28128 (N_28128,N_27571,N_27987);
nand U28129 (N_28129,N_27619,N_27542);
or U28130 (N_28130,N_27584,N_27962);
or U28131 (N_28131,N_27821,N_27940);
xnor U28132 (N_28132,N_27742,N_27589);
nand U28133 (N_28133,N_27659,N_27723);
nor U28134 (N_28134,N_27592,N_27525);
and U28135 (N_28135,N_27875,N_27936);
and U28136 (N_28136,N_27731,N_27930);
or U28137 (N_28137,N_27829,N_27951);
and U28138 (N_28138,N_27893,N_27775);
nand U28139 (N_28139,N_27657,N_27965);
or U28140 (N_28140,N_27988,N_27891);
and U28141 (N_28141,N_27781,N_27877);
xnor U28142 (N_28142,N_27745,N_27699);
nor U28143 (N_28143,N_27803,N_27762);
xor U28144 (N_28144,N_27720,N_27882);
nor U28145 (N_28145,N_27705,N_27565);
or U28146 (N_28146,N_27646,N_27831);
nand U28147 (N_28147,N_27702,N_27822);
nor U28148 (N_28148,N_27622,N_27789);
nor U28149 (N_28149,N_27653,N_27562);
and U28150 (N_28150,N_27739,N_27637);
nand U28151 (N_28151,N_27549,N_27579);
xnor U28152 (N_28152,N_27769,N_27630);
xor U28153 (N_28153,N_27687,N_27727);
and U28154 (N_28154,N_27880,N_27527);
and U28155 (N_28155,N_27522,N_27825);
nor U28156 (N_28156,N_27848,N_27627);
and U28157 (N_28157,N_27798,N_27819);
and U28158 (N_28158,N_27518,N_27709);
nor U28159 (N_28159,N_27519,N_27661);
nor U28160 (N_28160,N_27914,N_27912);
or U28161 (N_28161,N_27853,N_27597);
nand U28162 (N_28162,N_27753,N_27809);
xnor U28163 (N_28163,N_27557,N_27703);
nor U28164 (N_28164,N_27560,N_27576);
xnor U28165 (N_28165,N_27634,N_27801);
nand U28166 (N_28166,N_27529,N_27611);
xnor U28167 (N_28167,N_27523,N_27968);
nand U28168 (N_28168,N_27617,N_27610);
nor U28169 (N_28169,N_27773,N_27888);
nor U28170 (N_28170,N_27548,N_27591);
nor U28171 (N_28171,N_27778,N_27820);
or U28172 (N_28172,N_27516,N_27504);
nor U28173 (N_28173,N_27555,N_27939);
xnor U28174 (N_28174,N_27713,N_27666);
xor U28175 (N_28175,N_27721,N_27678);
and U28176 (N_28176,N_27889,N_27743);
and U28177 (N_28177,N_27692,N_27604);
or U28178 (N_28178,N_27833,N_27639);
nor U28179 (N_28179,N_27680,N_27625);
nor U28180 (N_28180,N_27975,N_27567);
nand U28181 (N_28181,N_27632,N_27846);
and U28182 (N_28182,N_27668,N_27714);
xor U28183 (N_28183,N_27768,N_27952);
xor U28184 (N_28184,N_27670,N_27795);
or U28185 (N_28185,N_27620,N_27808);
nand U28186 (N_28186,N_27577,N_27859);
xnor U28187 (N_28187,N_27652,N_27506);
nor U28188 (N_28188,N_27526,N_27785);
nor U28189 (N_28189,N_27815,N_27901);
and U28190 (N_28190,N_27719,N_27928);
xnor U28191 (N_28191,N_27876,N_27694);
or U28192 (N_28192,N_27981,N_27802);
xor U28193 (N_28193,N_27904,N_27941);
and U28194 (N_28194,N_27986,N_27953);
nor U28195 (N_28195,N_27706,N_27918);
nor U28196 (N_28196,N_27689,N_27913);
nor U28197 (N_28197,N_27760,N_27793);
or U28198 (N_28198,N_27551,N_27543);
nand U28199 (N_28199,N_27660,N_27612);
and U28200 (N_28200,N_27711,N_27708);
and U28201 (N_28201,N_27575,N_27898);
nand U28202 (N_28202,N_27957,N_27665);
xor U28203 (N_28203,N_27895,N_27569);
nand U28204 (N_28204,N_27994,N_27915);
or U28205 (N_28205,N_27982,N_27503);
nand U28206 (N_28206,N_27899,N_27746);
and U28207 (N_28207,N_27812,N_27992);
nor U28208 (N_28208,N_27761,N_27573);
or U28209 (N_28209,N_27707,N_27566);
or U28210 (N_28210,N_27864,N_27570);
nand U28211 (N_28211,N_27704,N_27590);
nand U28212 (N_28212,N_27633,N_27643);
nand U28213 (N_28213,N_27929,N_27640);
nor U28214 (N_28214,N_27837,N_27695);
nor U28215 (N_28215,N_27856,N_27847);
or U28216 (N_28216,N_27967,N_27879);
or U28217 (N_28217,N_27614,N_27862);
nor U28218 (N_28218,N_27843,N_27983);
and U28219 (N_28219,N_27559,N_27845);
and U28220 (N_28220,N_27931,N_27991);
xnor U28221 (N_28221,N_27509,N_27887);
or U28222 (N_28222,N_27792,N_27964);
and U28223 (N_28223,N_27585,N_27814);
or U28224 (N_28224,N_27849,N_27956);
or U28225 (N_28225,N_27892,N_27995);
xor U28226 (N_28226,N_27698,N_27587);
xnor U28227 (N_28227,N_27536,N_27954);
and U28228 (N_28228,N_27924,N_27885);
nand U28229 (N_28229,N_27718,N_27520);
or U28230 (N_28230,N_27884,N_27679);
or U28231 (N_28231,N_27531,N_27844);
or U28232 (N_28232,N_27917,N_27755);
xor U28233 (N_28233,N_27517,N_27947);
and U28234 (N_28234,N_27946,N_27712);
xnor U28235 (N_28235,N_27886,N_27932);
nand U28236 (N_28236,N_27937,N_27782);
or U28237 (N_28237,N_27546,N_27772);
or U28238 (N_28238,N_27989,N_27586);
nor U28239 (N_28239,N_27766,N_27855);
nand U28240 (N_28240,N_27734,N_27605);
or U28241 (N_28241,N_27602,N_27920);
nand U28242 (N_28242,N_27997,N_27858);
and U28243 (N_28243,N_27945,N_27621);
and U28244 (N_28244,N_27902,N_27513);
and U28245 (N_28245,N_27535,N_27797);
or U28246 (N_28246,N_27501,N_27596);
and U28247 (N_28247,N_27942,N_27624);
and U28248 (N_28248,N_27545,N_27623);
xor U28249 (N_28249,N_27554,N_27544);
and U28250 (N_28250,N_27621,N_27641);
nand U28251 (N_28251,N_27898,N_27877);
nand U28252 (N_28252,N_27639,N_27610);
nand U28253 (N_28253,N_27704,N_27644);
and U28254 (N_28254,N_27508,N_27539);
or U28255 (N_28255,N_27572,N_27839);
nor U28256 (N_28256,N_27636,N_27748);
or U28257 (N_28257,N_27502,N_27732);
nor U28258 (N_28258,N_27851,N_27610);
nand U28259 (N_28259,N_27955,N_27754);
nor U28260 (N_28260,N_27567,N_27742);
and U28261 (N_28261,N_27612,N_27695);
or U28262 (N_28262,N_27905,N_27799);
nand U28263 (N_28263,N_27853,N_27997);
and U28264 (N_28264,N_27543,N_27559);
xnor U28265 (N_28265,N_27895,N_27949);
nor U28266 (N_28266,N_27615,N_27620);
or U28267 (N_28267,N_27652,N_27695);
and U28268 (N_28268,N_27927,N_27960);
nand U28269 (N_28269,N_27557,N_27807);
nor U28270 (N_28270,N_27947,N_27516);
and U28271 (N_28271,N_27842,N_27578);
or U28272 (N_28272,N_27812,N_27533);
nand U28273 (N_28273,N_27718,N_27965);
xor U28274 (N_28274,N_27702,N_27547);
nand U28275 (N_28275,N_27871,N_27866);
xnor U28276 (N_28276,N_27868,N_27947);
nand U28277 (N_28277,N_27511,N_27895);
nand U28278 (N_28278,N_27548,N_27941);
xnor U28279 (N_28279,N_27795,N_27889);
and U28280 (N_28280,N_27893,N_27784);
nor U28281 (N_28281,N_27981,N_27739);
nor U28282 (N_28282,N_27983,N_27954);
nor U28283 (N_28283,N_27609,N_27520);
xor U28284 (N_28284,N_27721,N_27914);
nor U28285 (N_28285,N_27833,N_27869);
nor U28286 (N_28286,N_27916,N_27961);
xor U28287 (N_28287,N_27652,N_27790);
or U28288 (N_28288,N_27912,N_27910);
and U28289 (N_28289,N_27780,N_27882);
nand U28290 (N_28290,N_27615,N_27976);
xnor U28291 (N_28291,N_27976,N_27816);
nand U28292 (N_28292,N_27783,N_27650);
and U28293 (N_28293,N_27858,N_27804);
nor U28294 (N_28294,N_27740,N_27640);
nand U28295 (N_28295,N_27832,N_27990);
nor U28296 (N_28296,N_27815,N_27756);
nor U28297 (N_28297,N_27901,N_27763);
nor U28298 (N_28298,N_27756,N_27726);
and U28299 (N_28299,N_27716,N_27999);
or U28300 (N_28300,N_27510,N_27653);
and U28301 (N_28301,N_27955,N_27887);
and U28302 (N_28302,N_27862,N_27601);
and U28303 (N_28303,N_27936,N_27852);
or U28304 (N_28304,N_27881,N_27750);
or U28305 (N_28305,N_27940,N_27611);
xor U28306 (N_28306,N_27890,N_27948);
nor U28307 (N_28307,N_27504,N_27907);
nand U28308 (N_28308,N_27978,N_27746);
xor U28309 (N_28309,N_27795,N_27959);
or U28310 (N_28310,N_27553,N_27550);
xor U28311 (N_28311,N_27576,N_27745);
nor U28312 (N_28312,N_27589,N_27735);
or U28313 (N_28313,N_27770,N_27521);
nand U28314 (N_28314,N_27836,N_27670);
nor U28315 (N_28315,N_27546,N_27693);
nor U28316 (N_28316,N_27553,N_27808);
and U28317 (N_28317,N_27775,N_27567);
xor U28318 (N_28318,N_27511,N_27760);
and U28319 (N_28319,N_27867,N_27786);
xor U28320 (N_28320,N_27546,N_27655);
nand U28321 (N_28321,N_27947,N_27688);
or U28322 (N_28322,N_27800,N_27614);
or U28323 (N_28323,N_27679,N_27771);
and U28324 (N_28324,N_27758,N_27932);
and U28325 (N_28325,N_27893,N_27937);
or U28326 (N_28326,N_27596,N_27580);
or U28327 (N_28327,N_27661,N_27567);
and U28328 (N_28328,N_27673,N_27679);
nand U28329 (N_28329,N_27928,N_27573);
xor U28330 (N_28330,N_27541,N_27803);
and U28331 (N_28331,N_27946,N_27985);
or U28332 (N_28332,N_27785,N_27851);
or U28333 (N_28333,N_27592,N_27581);
and U28334 (N_28334,N_27739,N_27724);
nor U28335 (N_28335,N_27793,N_27566);
nor U28336 (N_28336,N_27722,N_27887);
xnor U28337 (N_28337,N_27728,N_27799);
or U28338 (N_28338,N_27930,N_27699);
nand U28339 (N_28339,N_27954,N_27799);
or U28340 (N_28340,N_27706,N_27932);
nand U28341 (N_28341,N_27545,N_27691);
nor U28342 (N_28342,N_27842,N_27929);
xnor U28343 (N_28343,N_27798,N_27584);
nor U28344 (N_28344,N_27976,N_27643);
and U28345 (N_28345,N_27803,N_27729);
or U28346 (N_28346,N_27967,N_27620);
or U28347 (N_28347,N_27816,N_27884);
nand U28348 (N_28348,N_27580,N_27855);
or U28349 (N_28349,N_27571,N_27817);
nor U28350 (N_28350,N_27923,N_27985);
and U28351 (N_28351,N_27590,N_27641);
nand U28352 (N_28352,N_27702,N_27634);
xor U28353 (N_28353,N_27761,N_27636);
and U28354 (N_28354,N_27545,N_27749);
nand U28355 (N_28355,N_27854,N_27725);
xor U28356 (N_28356,N_27943,N_27676);
xor U28357 (N_28357,N_27771,N_27815);
xnor U28358 (N_28358,N_27845,N_27595);
nor U28359 (N_28359,N_27789,N_27733);
and U28360 (N_28360,N_27773,N_27649);
nand U28361 (N_28361,N_27690,N_27590);
nand U28362 (N_28362,N_27681,N_27565);
xnor U28363 (N_28363,N_27956,N_27804);
nor U28364 (N_28364,N_27659,N_27699);
or U28365 (N_28365,N_27737,N_27509);
xor U28366 (N_28366,N_27682,N_27980);
nor U28367 (N_28367,N_27733,N_27825);
nand U28368 (N_28368,N_27952,N_27755);
nand U28369 (N_28369,N_27681,N_27659);
nor U28370 (N_28370,N_27794,N_27797);
or U28371 (N_28371,N_27818,N_27725);
nor U28372 (N_28372,N_27527,N_27864);
nand U28373 (N_28373,N_27832,N_27955);
or U28374 (N_28374,N_27839,N_27814);
or U28375 (N_28375,N_27670,N_27699);
nand U28376 (N_28376,N_27945,N_27635);
and U28377 (N_28377,N_27783,N_27511);
or U28378 (N_28378,N_27547,N_27633);
xor U28379 (N_28379,N_27750,N_27736);
nor U28380 (N_28380,N_27949,N_27625);
nand U28381 (N_28381,N_27758,N_27616);
nand U28382 (N_28382,N_27591,N_27931);
nand U28383 (N_28383,N_27718,N_27684);
nor U28384 (N_28384,N_27850,N_27908);
xor U28385 (N_28385,N_27810,N_27717);
or U28386 (N_28386,N_27653,N_27535);
or U28387 (N_28387,N_27986,N_27686);
xnor U28388 (N_28388,N_27853,N_27959);
and U28389 (N_28389,N_27966,N_27756);
nor U28390 (N_28390,N_27522,N_27701);
or U28391 (N_28391,N_27723,N_27631);
nor U28392 (N_28392,N_27527,N_27583);
nand U28393 (N_28393,N_27837,N_27550);
or U28394 (N_28394,N_27881,N_27850);
xor U28395 (N_28395,N_27519,N_27967);
and U28396 (N_28396,N_27814,N_27979);
xor U28397 (N_28397,N_27641,N_27656);
nand U28398 (N_28398,N_27705,N_27560);
xnor U28399 (N_28399,N_27721,N_27748);
xnor U28400 (N_28400,N_27847,N_27806);
and U28401 (N_28401,N_27982,N_27549);
nor U28402 (N_28402,N_27736,N_27747);
xnor U28403 (N_28403,N_27857,N_27625);
nand U28404 (N_28404,N_27787,N_27680);
xor U28405 (N_28405,N_27690,N_27721);
and U28406 (N_28406,N_27981,N_27594);
or U28407 (N_28407,N_27892,N_27664);
and U28408 (N_28408,N_27517,N_27502);
nor U28409 (N_28409,N_27954,N_27679);
xor U28410 (N_28410,N_27667,N_27885);
or U28411 (N_28411,N_27570,N_27811);
xor U28412 (N_28412,N_27824,N_27836);
or U28413 (N_28413,N_27949,N_27748);
or U28414 (N_28414,N_27751,N_27639);
nand U28415 (N_28415,N_27983,N_27962);
nor U28416 (N_28416,N_27699,N_27801);
xnor U28417 (N_28417,N_27800,N_27598);
xnor U28418 (N_28418,N_27814,N_27685);
nand U28419 (N_28419,N_27597,N_27814);
or U28420 (N_28420,N_27720,N_27895);
nor U28421 (N_28421,N_27809,N_27680);
and U28422 (N_28422,N_27730,N_27738);
xor U28423 (N_28423,N_27874,N_27628);
or U28424 (N_28424,N_27977,N_27875);
or U28425 (N_28425,N_27705,N_27629);
or U28426 (N_28426,N_27974,N_27512);
and U28427 (N_28427,N_27522,N_27535);
nor U28428 (N_28428,N_27625,N_27667);
nand U28429 (N_28429,N_27686,N_27669);
nand U28430 (N_28430,N_27941,N_27902);
and U28431 (N_28431,N_27569,N_27887);
nor U28432 (N_28432,N_27583,N_27965);
or U28433 (N_28433,N_27572,N_27790);
nor U28434 (N_28434,N_27791,N_27958);
nand U28435 (N_28435,N_27696,N_27609);
nor U28436 (N_28436,N_27787,N_27876);
nand U28437 (N_28437,N_27915,N_27614);
nor U28438 (N_28438,N_27950,N_27562);
nand U28439 (N_28439,N_27940,N_27630);
nand U28440 (N_28440,N_27538,N_27855);
and U28441 (N_28441,N_27856,N_27541);
and U28442 (N_28442,N_27878,N_27679);
nor U28443 (N_28443,N_27797,N_27911);
and U28444 (N_28444,N_27692,N_27711);
and U28445 (N_28445,N_27754,N_27861);
and U28446 (N_28446,N_27996,N_27809);
xnor U28447 (N_28447,N_27878,N_27732);
xor U28448 (N_28448,N_27706,N_27894);
nor U28449 (N_28449,N_27664,N_27989);
nand U28450 (N_28450,N_27805,N_27588);
or U28451 (N_28451,N_27843,N_27851);
or U28452 (N_28452,N_27803,N_27515);
xor U28453 (N_28453,N_27738,N_27903);
xnor U28454 (N_28454,N_27508,N_27777);
and U28455 (N_28455,N_27869,N_27762);
nor U28456 (N_28456,N_27853,N_27690);
and U28457 (N_28457,N_27551,N_27726);
or U28458 (N_28458,N_27664,N_27510);
and U28459 (N_28459,N_27915,N_27533);
nor U28460 (N_28460,N_27510,N_27698);
xor U28461 (N_28461,N_27825,N_27878);
and U28462 (N_28462,N_27779,N_27763);
or U28463 (N_28463,N_27816,N_27579);
xnor U28464 (N_28464,N_27872,N_27893);
and U28465 (N_28465,N_27815,N_27633);
and U28466 (N_28466,N_27854,N_27794);
xor U28467 (N_28467,N_27699,N_27725);
and U28468 (N_28468,N_27758,N_27571);
and U28469 (N_28469,N_27635,N_27800);
xnor U28470 (N_28470,N_27726,N_27712);
nor U28471 (N_28471,N_27662,N_27976);
xor U28472 (N_28472,N_27922,N_27631);
nor U28473 (N_28473,N_27531,N_27591);
and U28474 (N_28474,N_27511,N_27891);
nor U28475 (N_28475,N_27884,N_27841);
xor U28476 (N_28476,N_27706,N_27518);
and U28477 (N_28477,N_27685,N_27693);
nand U28478 (N_28478,N_27691,N_27628);
xor U28479 (N_28479,N_27859,N_27576);
nand U28480 (N_28480,N_27797,N_27713);
nor U28481 (N_28481,N_27793,N_27922);
and U28482 (N_28482,N_27958,N_27792);
nor U28483 (N_28483,N_27521,N_27665);
xnor U28484 (N_28484,N_27980,N_27854);
and U28485 (N_28485,N_27750,N_27611);
and U28486 (N_28486,N_27540,N_27644);
xor U28487 (N_28487,N_27603,N_27591);
or U28488 (N_28488,N_27803,N_27681);
nor U28489 (N_28489,N_27815,N_27559);
xnor U28490 (N_28490,N_27698,N_27771);
or U28491 (N_28491,N_27599,N_27754);
or U28492 (N_28492,N_27572,N_27994);
and U28493 (N_28493,N_27935,N_27878);
or U28494 (N_28494,N_27828,N_27895);
and U28495 (N_28495,N_27931,N_27559);
or U28496 (N_28496,N_27601,N_27615);
nor U28497 (N_28497,N_27604,N_27992);
nand U28498 (N_28498,N_27912,N_27502);
and U28499 (N_28499,N_27783,N_27587);
or U28500 (N_28500,N_28239,N_28455);
nor U28501 (N_28501,N_28301,N_28438);
nor U28502 (N_28502,N_28136,N_28374);
nor U28503 (N_28503,N_28055,N_28447);
nor U28504 (N_28504,N_28352,N_28103);
nand U28505 (N_28505,N_28470,N_28068);
nand U28506 (N_28506,N_28014,N_28430);
and U28507 (N_28507,N_28403,N_28385);
nor U28508 (N_28508,N_28332,N_28356);
xnor U28509 (N_28509,N_28324,N_28446);
and U28510 (N_28510,N_28180,N_28183);
or U28511 (N_28511,N_28229,N_28241);
nand U28512 (N_28512,N_28484,N_28432);
nor U28513 (N_28513,N_28348,N_28359);
or U28514 (N_28514,N_28380,N_28145);
or U28515 (N_28515,N_28207,N_28233);
or U28516 (N_28516,N_28031,N_28066);
xnor U28517 (N_28517,N_28421,N_28046);
nand U28518 (N_28518,N_28429,N_28108);
xor U28519 (N_28519,N_28431,N_28354);
nand U28520 (N_28520,N_28258,N_28069);
xor U28521 (N_28521,N_28246,N_28290);
and U28522 (N_28522,N_28110,N_28237);
or U28523 (N_28523,N_28276,N_28414);
nand U28524 (N_28524,N_28130,N_28363);
nand U28525 (N_28525,N_28027,N_28309);
nor U28526 (N_28526,N_28169,N_28373);
nor U28527 (N_28527,N_28372,N_28342);
and U28528 (N_28528,N_28409,N_28123);
and U28529 (N_28529,N_28305,N_28405);
nor U28530 (N_28530,N_28023,N_28201);
nor U28531 (N_28531,N_28057,N_28115);
nand U28532 (N_28532,N_28378,N_28442);
or U28533 (N_28533,N_28050,N_28102);
or U28534 (N_28534,N_28141,N_28077);
or U28535 (N_28535,N_28216,N_28091);
and U28536 (N_28536,N_28061,N_28079);
or U28537 (N_28537,N_28310,N_28037);
nand U28538 (N_28538,N_28010,N_28499);
xor U28539 (N_28539,N_28347,N_28304);
and U28540 (N_28540,N_28049,N_28357);
and U28541 (N_28541,N_28179,N_28181);
nor U28542 (N_28542,N_28424,N_28479);
or U28543 (N_28543,N_28029,N_28004);
and U28544 (N_28544,N_28149,N_28428);
and U28545 (N_28545,N_28056,N_28298);
nand U28546 (N_28546,N_28096,N_28367);
xor U28547 (N_28547,N_28411,N_28022);
or U28548 (N_28548,N_28376,N_28393);
xor U28549 (N_28549,N_28427,N_28158);
and U28550 (N_28550,N_28370,N_28016);
or U28551 (N_28551,N_28351,N_28089);
xnor U28552 (N_28552,N_28490,N_28238);
or U28553 (N_28553,N_28331,N_28090);
nor U28554 (N_28554,N_28398,N_28203);
xnor U28555 (N_28555,N_28418,N_28340);
nand U28556 (N_28556,N_28255,N_28106);
and U28557 (N_28557,N_28457,N_28163);
xnor U28558 (N_28558,N_28485,N_28150);
xor U28559 (N_28559,N_28425,N_28140);
nand U28560 (N_28560,N_28307,N_28086);
nand U28561 (N_28561,N_28226,N_28338);
nor U28562 (N_28562,N_28256,N_28253);
and U28563 (N_28563,N_28325,N_28048);
or U28564 (N_28564,N_28058,N_28282);
xor U28565 (N_28565,N_28406,N_28467);
or U28566 (N_28566,N_28222,N_28283);
and U28567 (N_28567,N_28420,N_28146);
or U28568 (N_28568,N_28364,N_28084);
xor U28569 (N_28569,N_28394,N_28192);
nand U28570 (N_28570,N_28471,N_28085);
xnor U28571 (N_28571,N_28137,N_28041);
nand U28572 (N_28572,N_28133,N_28371);
or U28573 (N_28573,N_28337,N_28087);
nor U28574 (N_28574,N_28320,N_28458);
and U28575 (N_28575,N_28111,N_28007);
or U28576 (N_28576,N_28142,N_28333);
nand U28577 (N_28577,N_28412,N_28443);
nor U28578 (N_28578,N_28289,N_28186);
and U28579 (N_28579,N_28065,N_28159);
xnor U28580 (N_28580,N_28161,N_28097);
nand U28581 (N_28581,N_28071,N_28475);
nor U28582 (N_28582,N_28248,N_28217);
nor U28583 (N_28583,N_28189,N_28230);
nand U28584 (N_28584,N_28358,N_28225);
nand U28585 (N_28585,N_28040,N_28188);
or U28586 (N_28586,N_28441,N_28059);
nand U28587 (N_28587,N_28117,N_28134);
or U28588 (N_28588,N_28195,N_28033);
or U28589 (N_28589,N_28461,N_28328);
xnor U28590 (N_28590,N_28051,N_28015);
nand U28591 (N_28591,N_28082,N_28402);
xnor U28592 (N_28592,N_28361,N_28463);
xnor U28593 (N_28593,N_28291,N_28384);
nor U28594 (N_28594,N_28062,N_28336);
or U28595 (N_28595,N_28480,N_28350);
xor U28596 (N_28596,N_28001,N_28468);
xnor U28597 (N_28597,N_28210,N_28262);
or U28598 (N_28598,N_28275,N_28220);
nor U28599 (N_28599,N_28388,N_28121);
and U28600 (N_28600,N_28245,N_28172);
nand U28601 (N_28601,N_28284,N_28139);
and U28602 (N_28602,N_28026,N_28176);
or U28603 (N_28603,N_28017,N_28240);
nor U28604 (N_28604,N_28083,N_28346);
xnor U28605 (N_28605,N_28072,N_28138);
nor U28606 (N_28606,N_28032,N_28379);
or U28607 (N_28607,N_28482,N_28494);
and U28608 (N_28608,N_28391,N_28327);
nor U28609 (N_28609,N_28153,N_28131);
and U28610 (N_28610,N_28098,N_28362);
nor U28611 (N_28611,N_28168,N_28036);
xor U28612 (N_28612,N_28144,N_28116);
nor U28613 (N_28613,N_28281,N_28043);
nand U28614 (N_28614,N_28316,N_28143);
and U28615 (N_28615,N_28413,N_28382);
nor U28616 (N_28616,N_28278,N_28236);
or U28617 (N_28617,N_28473,N_28157);
nor U28618 (N_28618,N_28193,N_28219);
or U28619 (N_28619,N_28392,N_28271);
or U28620 (N_28620,N_28326,N_28250);
or U28621 (N_28621,N_28293,N_28148);
xor U28622 (N_28622,N_28400,N_28389);
or U28623 (N_28623,N_28197,N_28269);
or U28624 (N_28624,N_28063,N_28481);
nand U28625 (N_28625,N_28273,N_28488);
xor U28626 (N_28626,N_28487,N_28218);
nor U28627 (N_28627,N_28060,N_28044);
nand U28628 (N_28628,N_28349,N_28295);
or U28629 (N_28629,N_28317,N_28297);
and U28630 (N_28630,N_28177,N_28194);
or U28631 (N_28631,N_28377,N_28156);
nor U28632 (N_28632,N_28170,N_28109);
nor U28633 (N_28633,N_28094,N_28296);
or U28634 (N_28634,N_28025,N_28306);
xor U28635 (N_28635,N_28073,N_28011);
and U28636 (N_28636,N_28452,N_28280);
and U28637 (N_28637,N_28341,N_28088);
nand U28638 (N_28638,N_28323,N_28020);
or U28639 (N_28639,N_28205,N_28100);
nand U28640 (N_28640,N_28249,N_28232);
xnor U28641 (N_28641,N_28243,N_28019);
xor U28642 (N_28642,N_28129,N_28311);
nor U28643 (N_28643,N_28434,N_28000);
or U28644 (N_28644,N_28167,N_28439);
or U28645 (N_28645,N_28302,N_28396);
or U28646 (N_28646,N_28437,N_28335);
or U28647 (N_28647,N_28303,N_28469);
nand U28648 (N_28648,N_28399,N_28199);
nor U28649 (N_28649,N_28417,N_28407);
xor U28650 (N_28650,N_28215,N_28206);
or U28651 (N_28651,N_28006,N_28375);
xor U28652 (N_28652,N_28074,N_28449);
and U28653 (N_28653,N_28070,N_28478);
nand U28654 (N_28654,N_28265,N_28477);
or U28655 (N_28655,N_28314,N_28279);
nand U28656 (N_28656,N_28254,N_28005);
or U28657 (N_28657,N_28268,N_28285);
and U28658 (N_28658,N_28292,N_28287);
or U28659 (N_28659,N_28208,N_28496);
xnor U28660 (N_28660,N_28120,N_28360);
and U28661 (N_28661,N_28410,N_28235);
and U28662 (N_28662,N_28196,N_28453);
xor U28663 (N_28663,N_28259,N_28223);
and U28664 (N_28664,N_28459,N_28112);
nand U28665 (N_28665,N_28113,N_28247);
or U28666 (N_28666,N_28118,N_28387);
and U28667 (N_28667,N_28415,N_28002);
nor U28668 (N_28668,N_28288,N_28200);
or U28669 (N_28669,N_28003,N_28132);
xnor U28670 (N_28670,N_28191,N_28404);
or U28671 (N_28671,N_28178,N_28125);
and U28672 (N_28672,N_28093,N_28152);
nor U28673 (N_28673,N_28164,N_28483);
and U28674 (N_28674,N_28454,N_28300);
nand U28675 (N_28675,N_28187,N_28234);
nor U28676 (N_28676,N_28464,N_28299);
xor U28677 (N_28677,N_28104,N_28209);
nor U28678 (N_28678,N_28095,N_28105);
and U28679 (N_28679,N_28313,N_28173);
xor U28680 (N_28680,N_28476,N_28128);
and U28681 (N_28681,N_28368,N_28277);
or U28682 (N_28682,N_28423,N_28486);
and U28683 (N_28683,N_28008,N_28166);
nor U28684 (N_28684,N_28426,N_28204);
xnor U28685 (N_28685,N_28076,N_28224);
nor U28686 (N_28686,N_28127,N_28244);
or U28687 (N_28687,N_28024,N_28039);
xor U28688 (N_28688,N_28472,N_28184);
and U28689 (N_28689,N_28312,N_28242);
and U28690 (N_28690,N_28462,N_28042);
xnor U28691 (N_28691,N_28264,N_28135);
and U28692 (N_28692,N_28053,N_28498);
or U28693 (N_28693,N_28344,N_28185);
nand U28694 (N_28694,N_28445,N_28272);
nand U28695 (N_28695,N_28274,N_28101);
and U28696 (N_28696,N_28345,N_28366);
and U28697 (N_28697,N_28260,N_28221);
or U28698 (N_28698,N_28021,N_28081);
nand U28699 (N_28699,N_28013,N_28365);
nand U28700 (N_28700,N_28497,N_28329);
nand U28701 (N_28701,N_28495,N_28444);
xor U28702 (N_28702,N_28492,N_28231);
or U28703 (N_28703,N_28251,N_28450);
nor U28704 (N_28704,N_28092,N_28381);
nand U28705 (N_28705,N_28182,N_28227);
and U28706 (N_28706,N_28212,N_28343);
xor U28707 (N_28707,N_28319,N_28416);
nand U28708 (N_28708,N_28321,N_28047);
or U28709 (N_28709,N_28114,N_28465);
and U28710 (N_28710,N_28160,N_28355);
nand U28711 (N_28711,N_28322,N_28162);
and U28712 (N_28712,N_28334,N_28436);
or U28713 (N_28713,N_28460,N_28390);
xor U28714 (N_28714,N_28211,N_28466);
or U28715 (N_28715,N_28214,N_28294);
and U28716 (N_28716,N_28151,N_28052);
xnor U28717 (N_28717,N_28315,N_28395);
or U28718 (N_28718,N_28228,N_28080);
nand U28719 (N_28719,N_28018,N_28078);
nand U28720 (N_28720,N_28067,N_28165);
and U28721 (N_28721,N_28034,N_28154);
nor U28722 (N_28722,N_28408,N_28038);
and U28723 (N_28723,N_28419,N_28339);
xnor U28724 (N_28724,N_28383,N_28126);
or U28725 (N_28725,N_28122,N_28286);
xnor U28726 (N_28726,N_28012,N_28124);
nand U28727 (N_28727,N_28318,N_28107);
or U28728 (N_28728,N_28030,N_28213);
or U28729 (N_28729,N_28252,N_28035);
nand U28730 (N_28730,N_28451,N_28147);
and U28731 (N_28731,N_28330,N_28491);
and U28732 (N_28732,N_28353,N_28456);
xor U28733 (N_28733,N_28489,N_28075);
nor U28734 (N_28734,N_28422,N_28270);
and U28735 (N_28735,N_28155,N_28190);
or U28736 (N_28736,N_28267,N_28202);
xor U28737 (N_28737,N_28064,N_28263);
or U28738 (N_28738,N_28198,N_28257);
and U28739 (N_28739,N_28435,N_28433);
or U28740 (N_28740,N_28493,N_28175);
nand U28741 (N_28741,N_28045,N_28054);
or U28742 (N_28742,N_28474,N_28174);
or U28743 (N_28743,N_28369,N_28028);
and U28744 (N_28744,N_28266,N_28261);
xnor U28745 (N_28745,N_28386,N_28308);
nand U28746 (N_28746,N_28119,N_28448);
nor U28747 (N_28747,N_28401,N_28099);
or U28748 (N_28748,N_28171,N_28440);
nand U28749 (N_28749,N_28009,N_28397);
and U28750 (N_28750,N_28386,N_28146);
or U28751 (N_28751,N_28409,N_28469);
nand U28752 (N_28752,N_28047,N_28002);
or U28753 (N_28753,N_28060,N_28012);
nand U28754 (N_28754,N_28020,N_28294);
or U28755 (N_28755,N_28042,N_28257);
and U28756 (N_28756,N_28117,N_28196);
xnor U28757 (N_28757,N_28052,N_28427);
nor U28758 (N_28758,N_28336,N_28453);
and U28759 (N_28759,N_28104,N_28030);
nor U28760 (N_28760,N_28270,N_28315);
xnor U28761 (N_28761,N_28337,N_28430);
and U28762 (N_28762,N_28388,N_28421);
xor U28763 (N_28763,N_28095,N_28047);
nor U28764 (N_28764,N_28387,N_28317);
or U28765 (N_28765,N_28444,N_28359);
xor U28766 (N_28766,N_28056,N_28213);
or U28767 (N_28767,N_28429,N_28140);
and U28768 (N_28768,N_28136,N_28431);
nand U28769 (N_28769,N_28238,N_28095);
nand U28770 (N_28770,N_28330,N_28105);
nor U28771 (N_28771,N_28078,N_28004);
nor U28772 (N_28772,N_28486,N_28086);
xor U28773 (N_28773,N_28127,N_28459);
and U28774 (N_28774,N_28298,N_28441);
nand U28775 (N_28775,N_28009,N_28432);
or U28776 (N_28776,N_28438,N_28113);
nor U28777 (N_28777,N_28193,N_28317);
nor U28778 (N_28778,N_28205,N_28077);
and U28779 (N_28779,N_28391,N_28237);
xor U28780 (N_28780,N_28282,N_28385);
nor U28781 (N_28781,N_28008,N_28124);
xor U28782 (N_28782,N_28255,N_28254);
nor U28783 (N_28783,N_28438,N_28117);
nand U28784 (N_28784,N_28143,N_28179);
nor U28785 (N_28785,N_28009,N_28359);
nand U28786 (N_28786,N_28347,N_28058);
nand U28787 (N_28787,N_28051,N_28489);
xor U28788 (N_28788,N_28448,N_28209);
and U28789 (N_28789,N_28013,N_28125);
xnor U28790 (N_28790,N_28418,N_28380);
nor U28791 (N_28791,N_28107,N_28454);
and U28792 (N_28792,N_28347,N_28052);
or U28793 (N_28793,N_28078,N_28061);
nand U28794 (N_28794,N_28035,N_28199);
or U28795 (N_28795,N_28245,N_28341);
nor U28796 (N_28796,N_28307,N_28277);
and U28797 (N_28797,N_28359,N_28406);
xor U28798 (N_28798,N_28005,N_28392);
or U28799 (N_28799,N_28069,N_28383);
nand U28800 (N_28800,N_28462,N_28248);
and U28801 (N_28801,N_28485,N_28311);
nand U28802 (N_28802,N_28428,N_28440);
nor U28803 (N_28803,N_28488,N_28145);
and U28804 (N_28804,N_28231,N_28334);
nand U28805 (N_28805,N_28100,N_28275);
or U28806 (N_28806,N_28185,N_28368);
xor U28807 (N_28807,N_28497,N_28259);
xor U28808 (N_28808,N_28408,N_28279);
nand U28809 (N_28809,N_28324,N_28185);
nor U28810 (N_28810,N_28290,N_28447);
nor U28811 (N_28811,N_28093,N_28210);
or U28812 (N_28812,N_28165,N_28480);
xor U28813 (N_28813,N_28045,N_28337);
nand U28814 (N_28814,N_28015,N_28004);
xnor U28815 (N_28815,N_28075,N_28116);
nor U28816 (N_28816,N_28045,N_28412);
xor U28817 (N_28817,N_28319,N_28056);
xor U28818 (N_28818,N_28488,N_28307);
and U28819 (N_28819,N_28411,N_28350);
nand U28820 (N_28820,N_28356,N_28293);
xor U28821 (N_28821,N_28392,N_28048);
and U28822 (N_28822,N_28204,N_28269);
and U28823 (N_28823,N_28187,N_28494);
or U28824 (N_28824,N_28290,N_28180);
xnor U28825 (N_28825,N_28359,N_28365);
nor U28826 (N_28826,N_28337,N_28413);
or U28827 (N_28827,N_28335,N_28050);
xnor U28828 (N_28828,N_28037,N_28465);
or U28829 (N_28829,N_28433,N_28214);
nand U28830 (N_28830,N_28269,N_28483);
or U28831 (N_28831,N_28060,N_28399);
nor U28832 (N_28832,N_28439,N_28077);
xor U28833 (N_28833,N_28417,N_28349);
nand U28834 (N_28834,N_28465,N_28440);
nand U28835 (N_28835,N_28064,N_28342);
and U28836 (N_28836,N_28348,N_28012);
xor U28837 (N_28837,N_28108,N_28459);
nand U28838 (N_28838,N_28159,N_28246);
and U28839 (N_28839,N_28067,N_28219);
or U28840 (N_28840,N_28375,N_28422);
and U28841 (N_28841,N_28402,N_28086);
or U28842 (N_28842,N_28167,N_28133);
nor U28843 (N_28843,N_28314,N_28447);
or U28844 (N_28844,N_28031,N_28304);
nand U28845 (N_28845,N_28318,N_28384);
or U28846 (N_28846,N_28400,N_28382);
xor U28847 (N_28847,N_28164,N_28023);
xnor U28848 (N_28848,N_28304,N_28177);
and U28849 (N_28849,N_28453,N_28162);
nand U28850 (N_28850,N_28370,N_28436);
and U28851 (N_28851,N_28263,N_28254);
nand U28852 (N_28852,N_28453,N_28224);
or U28853 (N_28853,N_28031,N_28098);
or U28854 (N_28854,N_28168,N_28043);
xor U28855 (N_28855,N_28496,N_28060);
nor U28856 (N_28856,N_28169,N_28464);
nand U28857 (N_28857,N_28280,N_28063);
nand U28858 (N_28858,N_28409,N_28242);
nand U28859 (N_28859,N_28259,N_28171);
nand U28860 (N_28860,N_28490,N_28284);
xor U28861 (N_28861,N_28123,N_28190);
and U28862 (N_28862,N_28089,N_28426);
or U28863 (N_28863,N_28497,N_28327);
nand U28864 (N_28864,N_28427,N_28262);
nand U28865 (N_28865,N_28109,N_28038);
and U28866 (N_28866,N_28323,N_28465);
nor U28867 (N_28867,N_28457,N_28425);
and U28868 (N_28868,N_28351,N_28227);
or U28869 (N_28869,N_28049,N_28365);
and U28870 (N_28870,N_28376,N_28108);
xor U28871 (N_28871,N_28360,N_28435);
xor U28872 (N_28872,N_28119,N_28141);
or U28873 (N_28873,N_28385,N_28241);
nand U28874 (N_28874,N_28086,N_28427);
and U28875 (N_28875,N_28393,N_28054);
and U28876 (N_28876,N_28190,N_28284);
or U28877 (N_28877,N_28025,N_28214);
nor U28878 (N_28878,N_28492,N_28335);
or U28879 (N_28879,N_28364,N_28070);
xnor U28880 (N_28880,N_28062,N_28464);
or U28881 (N_28881,N_28357,N_28356);
and U28882 (N_28882,N_28408,N_28369);
and U28883 (N_28883,N_28220,N_28397);
and U28884 (N_28884,N_28443,N_28320);
or U28885 (N_28885,N_28207,N_28032);
nand U28886 (N_28886,N_28316,N_28252);
nand U28887 (N_28887,N_28004,N_28482);
and U28888 (N_28888,N_28251,N_28173);
and U28889 (N_28889,N_28067,N_28373);
nor U28890 (N_28890,N_28167,N_28455);
nor U28891 (N_28891,N_28323,N_28492);
and U28892 (N_28892,N_28227,N_28488);
or U28893 (N_28893,N_28078,N_28102);
nor U28894 (N_28894,N_28183,N_28482);
and U28895 (N_28895,N_28362,N_28037);
nor U28896 (N_28896,N_28208,N_28196);
nor U28897 (N_28897,N_28022,N_28238);
xor U28898 (N_28898,N_28419,N_28031);
xnor U28899 (N_28899,N_28130,N_28313);
nor U28900 (N_28900,N_28119,N_28162);
xor U28901 (N_28901,N_28008,N_28284);
nor U28902 (N_28902,N_28126,N_28199);
or U28903 (N_28903,N_28391,N_28269);
nor U28904 (N_28904,N_28104,N_28254);
nor U28905 (N_28905,N_28262,N_28106);
nand U28906 (N_28906,N_28207,N_28215);
nand U28907 (N_28907,N_28418,N_28092);
and U28908 (N_28908,N_28141,N_28302);
xnor U28909 (N_28909,N_28006,N_28286);
nor U28910 (N_28910,N_28024,N_28102);
xnor U28911 (N_28911,N_28252,N_28056);
and U28912 (N_28912,N_28155,N_28498);
nand U28913 (N_28913,N_28391,N_28159);
or U28914 (N_28914,N_28198,N_28124);
and U28915 (N_28915,N_28181,N_28363);
xor U28916 (N_28916,N_28292,N_28320);
and U28917 (N_28917,N_28182,N_28143);
nand U28918 (N_28918,N_28421,N_28448);
nor U28919 (N_28919,N_28138,N_28411);
or U28920 (N_28920,N_28129,N_28093);
and U28921 (N_28921,N_28092,N_28172);
nand U28922 (N_28922,N_28049,N_28325);
nor U28923 (N_28923,N_28446,N_28358);
xnor U28924 (N_28924,N_28442,N_28203);
nor U28925 (N_28925,N_28173,N_28435);
or U28926 (N_28926,N_28474,N_28259);
nand U28927 (N_28927,N_28153,N_28298);
or U28928 (N_28928,N_28267,N_28205);
or U28929 (N_28929,N_28467,N_28122);
or U28930 (N_28930,N_28386,N_28258);
xnor U28931 (N_28931,N_28000,N_28225);
or U28932 (N_28932,N_28279,N_28151);
nor U28933 (N_28933,N_28290,N_28401);
or U28934 (N_28934,N_28393,N_28447);
and U28935 (N_28935,N_28260,N_28263);
nand U28936 (N_28936,N_28189,N_28281);
nor U28937 (N_28937,N_28091,N_28262);
or U28938 (N_28938,N_28206,N_28279);
xnor U28939 (N_28939,N_28333,N_28442);
nand U28940 (N_28940,N_28350,N_28475);
nand U28941 (N_28941,N_28242,N_28362);
and U28942 (N_28942,N_28376,N_28298);
and U28943 (N_28943,N_28385,N_28375);
and U28944 (N_28944,N_28281,N_28039);
nand U28945 (N_28945,N_28457,N_28237);
or U28946 (N_28946,N_28182,N_28429);
nor U28947 (N_28947,N_28349,N_28488);
nand U28948 (N_28948,N_28169,N_28002);
or U28949 (N_28949,N_28329,N_28352);
or U28950 (N_28950,N_28480,N_28241);
or U28951 (N_28951,N_28386,N_28032);
nor U28952 (N_28952,N_28332,N_28284);
and U28953 (N_28953,N_28108,N_28221);
and U28954 (N_28954,N_28336,N_28189);
nand U28955 (N_28955,N_28288,N_28015);
nand U28956 (N_28956,N_28392,N_28267);
or U28957 (N_28957,N_28275,N_28176);
xnor U28958 (N_28958,N_28138,N_28225);
nor U28959 (N_28959,N_28208,N_28065);
xnor U28960 (N_28960,N_28125,N_28102);
nor U28961 (N_28961,N_28112,N_28430);
nand U28962 (N_28962,N_28138,N_28359);
nand U28963 (N_28963,N_28416,N_28236);
nor U28964 (N_28964,N_28066,N_28380);
nand U28965 (N_28965,N_28113,N_28454);
and U28966 (N_28966,N_28106,N_28128);
nand U28967 (N_28967,N_28184,N_28231);
xor U28968 (N_28968,N_28148,N_28085);
and U28969 (N_28969,N_28365,N_28441);
and U28970 (N_28970,N_28380,N_28071);
xnor U28971 (N_28971,N_28253,N_28059);
and U28972 (N_28972,N_28322,N_28319);
nand U28973 (N_28973,N_28240,N_28499);
and U28974 (N_28974,N_28017,N_28421);
or U28975 (N_28975,N_28296,N_28293);
and U28976 (N_28976,N_28211,N_28365);
and U28977 (N_28977,N_28332,N_28450);
xor U28978 (N_28978,N_28015,N_28192);
and U28979 (N_28979,N_28218,N_28461);
xnor U28980 (N_28980,N_28342,N_28410);
nand U28981 (N_28981,N_28289,N_28338);
or U28982 (N_28982,N_28351,N_28141);
nand U28983 (N_28983,N_28411,N_28178);
nand U28984 (N_28984,N_28092,N_28440);
nand U28985 (N_28985,N_28159,N_28204);
or U28986 (N_28986,N_28429,N_28313);
nor U28987 (N_28987,N_28293,N_28341);
nand U28988 (N_28988,N_28401,N_28420);
xnor U28989 (N_28989,N_28016,N_28135);
or U28990 (N_28990,N_28345,N_28028);
nand U28991 (N_28991,N_28087,N_28059);
nor U28992 (N_28992,N_28336,N_28092);
nand U28993 (N_28993,N_28464,N_28383);
or U28994 (N_28994,N_28250,N_28343);
nor U28995 (N_28995,N_28282,N_28026);
or U28996 (N_28996,N_28357,N_28069);
or U28997 (N_28997,N_28051,N_28182);
and U28998 (N_28998,N_28129,N_28080);
nand U28999 (N_28999,N_28153,N_28221);
nand U29000 (N_29000,N_28954,N_28810);
nor U29001 (N_29001,N_28703,N_28501);
nand U29002 (N_29002,N_28879,N_28798);
xnor U29003 (N_29003,N_28952,N_28697);
nand U29004 (N_29004,N_28995,N_28631);
xor U29005 (N_29005,N_28532,N_28706);
xor U29006 (N_29006,N_28669,N_28593);
nor U29007 (N_29007,N_28909,N_28989);
or U29008 (N_29008,N_28639,N_28524);
xor U29009 (N_29009,N_28663,N_28903);
xnor U29010 (N_29010,N_28745,N_28737);
and U29011 (N_29011,N_28727,N_28950);
or U29012 (N_29012,N_28625,N_28980);
xor U29013 (N_29013,N_28585,N_28734);
xor U29014 (N_29014,N_28702,N_28761);
and U29015 (N_29015,N_28534,N_28785);
or U29016 (N_29016,N_28672,N_28851);
nand U29017 (N_29017,N_28620,N_28649);
nor U29018 (N_29018,N_28956,N_28522);
xnor U29019 (N_29019,N_28997,N_28555);
nand U29020 (N_29020,N_28875,N_28780);
xor U29021 (N_29021,N_28644,N_28862);
nand U29022 (N_29022,N_28874,N_28882);
or U29023 (N_29023,N_28544,N_28947);
nor U29024 (N_29024,N_28513,N_28925);
nor U29025 (N_29025,N_28633,N_28720);
xor U29026 (N_29026,N_28955,N_28677);
or U29027 (N_29027,N_28622,N_28987);
nand U29028 (N_29028,N_28948,N_28923);
and U29029 (N_29029,N_28542,N_28628);
xor U29030 (N_29030,N_28578,N_28605);
or U29031 (N_29031,N_28968,N_28523);
or U29032 (N_29032,N_28796,N_28673);
and U29033 (N_29033,N_28566,N_28732);
and U29034 (N_29034,N_28920,N_28864);
and U29035 (N_29035,N_28717,N_28951);
xnor U29036 (N_29036,N_28609,N_28567);
or U29037 (N_29037,N_28801,N_28881);
and U29038 (N_29038,N_28743,N_28825);
nand U29039 (N_29039,N_28809,N_28763);
or U29040 (N_29040,N_28531,N_28661);
or U29041 (N_29041,N_28539,N_28787);
nand U29042 (N_29042,N_28993,N_28502);
xor U29043 (N_29043,N_28844,N_28507);
xnor U29044 (N_29044,N_28814,N_28772);
and U29045 (N_29045,N_28797,N_28510);
nand U29046 (N_29046,N_28969,N_28617);
xor U29047 (N_29047,N_28754,N_28937);
xor U29048 (N_29048,N_28944,N_28515);
xnor U29049 (N_29049,N_28921,N_28652);
xor U29050 (N_29050,N_28843,N_28610);
xor U29051 (N_29051,N_28592,N_28675);
or U29052 (N_29052,N_28867,N_28831);
and U29053 (N_29053,N_28876,N_28670);
nor U29054 (N_29054,N_28816,N_28688);
xor U29055 (N_29055,N_28884,N_28840);
nand U29056 (N_29056,N_28758,N_28919);
nand U29057 (N_29057,N_28779,N_28619);
and U29058 (N_29058,N_28671,N_28521);
nand U29059 (N_29059,N_28709,N_28792);
or U29060 (N_29060,N_28505,N_28654);
xnor U29061 (N_29061,N_28568,N_28963);
nor U29062 (N_29062,N_28961,N_28943);
xor U29063 (N_29063,N_28612,N_28976);
nand U29064 (N_29064,N_28865,N_28778);
nor U29065 (N_29065,N_28829,N_28794);
xnor U29066 (N_29066,N_28646,N_28777);
nor U29067 (N_29067,N_28516,N_28888);
nand U29068 (N_29068,N_28603,N_28967);
nand U29069 (N_29069,N_28514,N_28551);
xnor U29070 (N_29070,N_28626,N_28711);
xor U29071 (N_29071,N_28791,N_28540);
and U29072 (N_29072,N_28695,N_28966);
or U29073 (N_29073,N_28666,N_28852);
nand U29074 (N_29074,N_28554,N_28580);
or U29075 (N_29075,N_28965,N_28811);
and U29076 (N_29076,N_28726,N_28691);
nor U29077 (N_29077,N_28945,N_28953);
and U29078 (N_29078,N_28984,N_28665);
or U29079 (N_29079,N_28596,N_28978);
nor U29080 (N_29080,N_28880,N_28667);
or U29081 (N_29081,N_28579,N_28838);
nand U29082 (N_29082,N_28598,N_28597);
nand U29083 (N_29083,N_28729,N_28648);
nor U29084 (N_29084,N_28616,N_28550);
nor U29085 (N_29085,N_28537,N_28922);
or U29086 (N_29086,N_28813,N_28519);
xnor U29087 (N_29087,N_28916,N_28553);
or U29088 (N_29088,N_28636,N_28569);
and U29089 (N_29089,N_28680,N_28728);
nand U29090 (N_29090,N_28664,N_28698);
and U29091 (N_29091,N_28802,N_28645);
nand U29092 (N_29092,N_28915,N_28640);
nand U29093 (N_29093,N_28520,N_28736);
or U29094 (N_29094,N_28863,N_28681);
and U29095 (N_29095,N_28694,N_28872);
and U29096 (N_29096,N_28774,N_28700);
and U29097 (N_29097,N_28739,N_28990);
nand U29098 (N_29098,N_28708,N_28715);
nand U29099 (N_29099,N_28582,N_28552);
and U29100 (N_29100,N_28946,N_28756);
or U29101 (N_29101,N_28602,N_28722);
nand U29102 (N_29102,N_28861,N_28784);
nand U29103 (N_29103,N_28575,N_28588);
and U29104 (N_29104,N_28559,N_28577);
nand U29105 (N_29105,N_28599,N_28614);
nor U29106 (N_29106,N_28674,N_28767);
or U29107 (N_29107,N_28890,N_28939);
nand U29108 (N_29108,N_28892,N_28590);
xor U29109 (N_29109,N_28750,N_28526);
or U29110 (N_29110,N_28710,N_28854);
nor U29111 (N_29111,N_28918,N_28871);
nor U29112 (N_29112,N_28988,N_28981);
or U29113 (N_29113,N_28701,N_28632);
xor U29114 (N_29114,N_28886,N_28819);
nand U29115 (N_29115,N_28817,N_28613);
and U29116 (N_29116,N_28744,N_28634);
xnor U29117 (N_29117,N_28781,N_28934);
xor U29118 (N_29118,N_28713,N_28860);
nand U29119 (N_29119,N_28856,N_28752);
xnor U29120 (N_29120,N_28933,N_28841);
xor U29121 (N_29121,N_28977,N_28790);
nand U29122 (N_29122,N_28679,N_28740);
nand U29123 (N_29123,N_28926,N_28941);
nand U29124 (N_29124,N_28583,N_28912);
nor U29125 (N_29125,N_28776,N_28799);
xnor U29126 (N_29126,N_28848,N_28741);
or U29127 (N_29127,N_28812,N_28857);
nand U29128 (N_29128,N_28899,N_28572);
and U29129 (N_29129,N_28601,N_28647);
or U29130 (N_29130,N_28508,N_28627);
and U29131 (N_29131,N_28716,N_28747);
nor U29132 (N_29132,N_28623,N_28742);
nand U29133 (N_29133,N_28653,N_28564);
nand U29134 (N_29134,N_28571,N_28746);
xnor U29135 (N_29135,N_28974,N_28805);
xnor U29136 (N_29136,N_28635,N_28725);
or U29137 (N_29137,N_28996,N_28705);
and U29138 (N_29138,N_28604,N_28975);
and U29139 (N_29139,N_28712,N_28998);
nor U29140 (N_29140,N_28558,N_28942);
or U29141 (N_29141,N_28893,N_28718);
and U29142 (N_29142,N_28894,N_28979);
nand U29143 (N_29143,N_28581,N_28846);
nor U29144 (N_29144,N_28775,N_28594);
xor U29145 (N_29145,N_28803,N_28731);
xor U29146 (N_29146,N_28949,N_28693);
and U29147 (N_29147,N_28656,N_28659);
nand U29148 (N_29148,N_28906,N_28958);
nor U29149 (N_29149,N_28897,N_28618);
and U29150 (N_29150,N_28836,N_28655);
nor U29151 (N_29151,N_28684,N_28985);
or U29152 (N_29152,N_28962,N_28678);
nor U29153 (N_29153,N_28707,N_28765);
or U29154 (N_29154,N_28541,N_28807);
nor U29155 (N_29155,N_28512,N_28904);
nor U29156 (N_29156,N_28660,N_28895);
nand U29157 (N_29157,N_28847,N_28690);
and U29158 (N_29158,N_28549,N_28692);
or U29159 (N_29159,N_28587,N_28629);
nor U29160 (N_29160,N_28859,N_28808);
xnor U29161 (N_29161,N_28839,N_28509);
xnor U29162 (N_29162,N_28749,N_28986);
and U29163 (N_29163,N_28891,N_28905);
nand U29164 (N_29164,N_28833,N_28611);
nor U29165 (N_29165,N_28768,N_28651);
or U29166 (N_29166,N_28608,N_28931);
xor U29167 (N_29167,N_28547,N_28806);
xor U29168 (N_29168,N_28957,N_28858);
xnor U29169 (N_29169,N_28936,N_28615);
and U29170 (N_29170,N_28548,N_28907);
and U29171 (N_29171,N_28910,N_28866);
and U29172 (N_29172,N_28911,N_28832);
xnor U29173 (N_29173,N_28517,N_28557);
nor U29174 (N_29174,N_28714,N_28855);
nand U29175 (N_29175,N_28721,N_28759);
nor U29176 (N_29176,N_28992,N_28538);
nand U29177 (N_29177,N_28683,N_28589);
xnor U29178 (N_29178,N_28535,N_28641);
and U29179 (N_29179,N_28826,N_28586);
nor U29180 (N_29180,N_28972,N_28887);
nor U29181 (N_29181,N_28823,N_28917);
xnor U29182 (N_29182,N_28773,N_28771);
or U29183 (N_29183,N_28543,N_28643);
xor U29184 (N_29184,N_28835,N_28927);
nand U29185 (N_29185,N_28682,N_28769);
nand U29186 (N_29186,N_28699,N_28650);
nor U29187 (N_29187,N_28970,N_28511);
or U29188 (N_29188,N_28533,N_28686);
nor U29189 (N_29189,N_28815,N_28658);
nand U29190 (N_29190,N_28935,N_28563);
xor U29191 (N_29191,N_28766,N_28999);
xnor U29192 (N_29192,N_28556,N_28574);
and U29193 (N_29193,N_28770,N_28696);
xor U29194 (N_29194,N_28724,N_28637);
or U29195 (N_29195,N_28687,N_28914);
or U29196 (N_29196,N_28793,N_28624);
nand U29197 (N_29197,N_28527,N_28530);
or U29198 (N_29198,N_28896,N_28940);
nor U29199 (N_29199,N_28938,N_28877);
nor U29200 (N_29200,N_28570,N_28735);
or U29201 (N_29201,N_28573,N_28500);
or U29202 (N_29202,N_28902,N_28748);
or U29203 (N_29203,N_28783,N_28506);
nor U29204 (N_29204,N_28719,N_28821);
nor U29205 (N_29205,N_28837,N_28789);
nor U29206 (N_29206,N_28845,N_28730);
and U29207 (N_29207,N_28788,N_28900);
nand U29208 (N_29208,N_28536,N_28878);
xnor U29209 (N_29209,N_28529,N_28804);
xor U29210 (N_29210,N_28822,N_28924);
xnor U29211 (N_29211,N_28930,N_28868);
nor U29212 (N_29212,N_28869,N_28503);
nor U29213 (N_29213,N_28800,N_28982);
nor U29214 (N_29214,N_28971,N_28818);
nand U29215 (N_29215,N_28753,N_28662);
xor U29216 (N_29216,N_28546,N_28638);
or U29217 (N_29217,N_28853,N_28689);
and U29218 (N_29218,N_28668,N_28723);
xnor U29219 (N_29219,N_28883,N_28782);
xor U29220 (N_29220,N_28762,N_28828);
and U29221 (N_29221,N_28561,N_28525);
nand U29222 (N_29222,N_28960,N_28606);
or U29223 (N_29223,N_28600,N_28760);
xnor U29224 (N_29224,N_28994,N_28764);
xor U29225 (N_29225,N_28834,N_28560);
nand U29226 (N_29226,N_28751,N_28518);
or U29227 (N_29227,N_28545,N_28959);
nand U29228 (N_29228,N_28820,N_28908);
nand U29229 (N_29229,N_28786,N_28591);
or U29230 (N_29230,N_28584,N_28504);
or U29231 (N_29231,N_28704,N_28929);
nor U29232 (N_29232,N_28913,N_28576);
xor U29233 (N_29233,N_28738,N_28973);
nor U29234 (N_29234,N_28873,N_28932);
nor U29235 (N_29235,N_28898,N_28901);
or U29236 (N_29236,N_28983,N_28757);
and U29237 (N_29237,N_28621,N_28850);
nor U29238 (N_29238,N_28676,N_28885);
xnor U29239 (N_29239,N_28928,N_28607);
xnor U29240 (N_29240,N_28889,N_28849);
nor U29241 (N_29241,N_28657,N_28685);
nor U29242 (N_29242,N_28830,N_28642);
xor U29243 (N_29243,N_28795,N_28870);
nor U29244 (N_29244,N_28755,N_28824);
xnor U29245 (N_29245,N_28991,N_28562);
nor U29246 (N_29246,N_28827,N_28630);
nor U29247 (N_29247,N_28733,N_28964);
xor U29248 (N_29248,N_28595,N_28565);
or U29249 (N_29249,N_28842,N_28528);
or U29250 (N_29250,N_28711,N_28973);
xor U29251 (N_29251,N_28705,N_28589);
nand U29252 (N_29252,N_28734,N_28833);
nor U29253 (N_29253,N_28809,N_28944);
and U29254 (N_29254,N_28593,N_28662);
nand U29255 (N_29255,N_28960,N_28902);
nand U29256 (N_29256,N_28824,N_28629);
and U29257 (N_29257,N_28979,N_28777);
or U29258 (N_29258,N_28874,N_28741);
xor U29259 (N_29259,N_28553,N_28779);
xor U29260 (N_29260,N_28966,N_28558);
or U29261 (N_29261,N_28571,N_28818);
and U29262 (N_29262,N_28646,N_28700);
xnor U29263 (N_29263,N_28504,N_28691);
xnor U29264 (N_29264,N_28826,N_28759);
nand U29265 (N_29265,N_28926,N_28901);
nand U29266 (N_29266,N_28905,N_28979);
nand U29267 (N_29267,N_28700,N_28948);
nor U29268 (N_29268,N_28555,N_28721);
and U29269 (N_29269,N_28919,N_28665);
nand U29270 (N_29270,N_28926,N_28679);
nor U29271 (N_29271,N_28672,N_28832);
nor U29272 (N_29272,N_28794,N_28924);
nand U29273 (N_29273,N_28510,N_28549);
nor U29274 (N_29274,N_28507,N_28860);
and U29275 (N_29275,N_28584,N_28804);
or U29276 (N_29276,N_28917,N_28583);
nand U29277 (N_29277,N_28509,N_28798);
nor U29278 (N_29278,N_28576,N_28725);
or U29279 (N_29279,N_28955,N_28556);
and U29280 (N_29280,N_28570,N_28752);
or U29281 (N_29281,N_28944,N_28614);
nand U29282 (N_29282,N_28682,N_28685);
nand U29283 (N_29283,N_28993,N_28602);
xor U29284 (N_29284,N_28958,N_28642);
xnor U29285 (N_29285,N_28784,N_28523);
nor U29286 (N_29286,N_28567,N_28806);
nand U29287 (N_29287,N_28829,N_28720);
nor U29288 (N_29288,N_28679,N_28617);
nor U29289 (N_29289,N_28947,N_28876);
xor U29290 (N_29290,N_28788,N_28846);
nand U29291 (N_29291,N_28738,N_28734);
and U29292 (N_29292,N_28988,N_28546);
nor U29293 (N_29293,N_28971,N_28751);
or U29294 (N_29294,N_28662,N_28555);
or U29295 (N_29295,N_28706,N_28939);
or U29296 (N_29296,N_28540,N_28502);
and U29297 (N_29297,N_28840,N_28901);
or U29298 (N_29298,N_28585,N_28868);
nand U29299 (N_29299,N_28999,N_28819);
xnor U29300 (N_29300,N_28572,N_28970);
nand U29301 (N_29301,N_28932,N_28862);
nor U29302 (N_29302,N_28553,N_28811);
or U29303 (N_29303,N_28685,N_28951);
nand U29304 (N_29304,N_28623,N_28561);
xnor U29305 (N_29305,N_28516,N_28751);
or U29306 (N_29306,N_28950,N_28520);
xnor U29307 (N_29307,N_28953,N_28952);
nand U29308 (N_29308,N_28952,N_28647);
or U29309 (N_29309,N_28875,N_28854);
nand U29310 (N_29310,N_28780,N_28624);
or U29311 (N_29311,N_28853,N_28701);
or U29312 (N_29312,N_28669,N_28703);
or U29313 (N_29313,N_28519,N_28557);
or U29314 (N_29314,N_28663,N_28826);
nor U29315 (N_29315,N_28891,N_28908);
nor U29316 (N_29316,N_28635,N_28839);
xor U29317 (N_29317,N_28977,N_28555);
nor U29318 (N_29318,N_28653,N_28562);
or U29319 (N_29319,N_28738,N_28757);
nor U29320 (N_29320,N_28573,N_28899);
xor U29321 (N_29321,N_28569,N_28616);
nor U29322 (N_29322,N_28947,N_28887);
xnor U29323 (N_29323,N_28983,N_28513);
and U29324 (N_29324,N_28894,N_28825);
xor U29325 (N_29325,N_28979,N_28573);
nor U29326 (N_29326,N_28640,N_28505);
nor U29327 (N_29327,N_28743,N_28991);
nor U29328 (N_29328,N_28580,N_28662);
or U29329 (N_29329,N_28770,N_28719);
and U29330 (N_29330,N_28675,N_28536);
xnor U29331 (N_29331,N_28804,N_28701);
and U29332 (N_29332,N_28951,N_28867);
and U29333 (N_29333,N_28923,N_28745);
or U29334 (N_29334,N_28826,N_28735);
and U29335 (N_29335,N_28553,N_28841);
and U29336 (N_29336,N_28793,N_28607);
or U29337 (N_29337,N_28633,N_28858);
xor U29338 (N_29338,N_28700,N_28529);
nor U29339 (N_29339,N_28997,N_28584);
and U29340 (N_29340,N_28743,N_28900);
and U29341 (N_29341,N_28587,N_28689);
nor U29342 (N_29342,N_28852,N_28812);
nand U29343 (N_29343,N_28913,N_28615);
or U29344 (N_29344,N_28626,N_28755);
and U29345 (N_29345,N_28674,N_28512);
nor U29346 (N_29346,N_28838,N_28960);
xor U29347 (N_29347,N_28557,N_28524);
xnor U29348 (N_29348,N_28783,N_28879);
xor U29349 (N_29349,N_28949,N_28729);
and U29350 (N_29350,N_28519,N_28570);
xor U29351 (N_29351,N_28732,N_28540);
nor U29352 (N_29352,N_28932,N_28620);
and U29353 (N_29353,N_28886,N_28996);
and U29354 (N_29354,N_28935,N_28802);
and U29355 (N_29355,N_28832,N_28527);
xor U29356 (N_29356,N_28553,N_28702);
nand U29357 (N_29357,N_28625,N_28521);
and U29358 (N_29358,N_28614,N_28876);
or U29359 (N_29359,N_28519,N_28805);
nand U29360 (N_29360,N_28699,N_28669);
xor U29361 (N_29361,N_28894,N_28804);
nand U29362 (N_29362,N_28935,N_28960);
nor U29363 (N_29363,N_28581,N_28745);
nor U29364 (N_29364,N_28782,N_28587);
and U29365 (N_29365,N_28654,N_28786);
xnor U29366 (N_29366,N_28904,N_28635);
nand U29367 (N_29367,N_28956,N_28507);
and U29368 (N_29368,N_28652,N_28845);
xnor U29369 (N_29369,N_28609,N_28910);
nor U29370 (N_29370,N_28552,N_28916);
and U29371 (N_29371,N_28503,N_28541);
nand U29372 (N_29372,N_28906,N_28713);
nand U29373 (N_29373,N_28814,N_28890);
and U29374 (N_29374,N_28576,N_28867);
and U29375 (N_29375,N_28799,N_28584);
and U29376 (N_29376,N_28820,N_28629);
xor U29377 (N_29377,N_28951,N_28648);
or U29378 (N_29378,N_28875,N_28540);
nor U29379 (N_29379,N_28850,N_28974);
nor U29380 (N_29380,N_28651,N_28724);
nand U29381 (N_29381,N_28624,N_28834);
and U29382 (N_29382,N_28651,N_28992);
nor U29383 (N_29383,N_28800,N_28673);
xnor U29384 (N_29384,N_28580,N_28762);
or U29385 (N_29385,N_28646,N_28624);
xnor U29386 (N_29386,N_28859,N_28551);
xnor U29387 (N_29387,N_28687,N_28867);
nand U29388 (N_29388,N_28699,N_28829);
nand U29389 (N_29389,N_28683,N_28765);
and U29390 (N_29390,N_28905,N_28984);
and U29391 (N_29391,N_28564,N_28931);
nor U29392 (N_29392,N_28954,N_28647);
or U29393 (N_29393,N_28715,N_28515);
or U29394 (N_29394,N_28763,N_28792);
or U29395 (N_29395,N_28809,N_28908);
and U29396 (N_29396,N_28944,N_28631);
nand U29397 (N_29397,N_28754,N_28839);
nor U29398 (N_29398,N_28507,N_28629);
xor U29399 (N_29399,N_28940,N_28979);
and U29400 (N_29400,N_28606,N_28944);
xnor U29401 (N_29401,N_28622,N_28998);
nor U29402 (N_29402,N_28538,N_28956);
or U29403 (N_29403,N_28969,N_28997);
xor U29404 (N_29404,N_28805,N_28698);
xor U29405 (N_29405,N_28813,N_28863);
nand U29406 (N_29406,N_28626,N_28874);
and U29407 (N_29407,N_28832,N_28809);
nor U29408 (N_29408,N_28823,N_28974);
xnor U29409 (N_29409,N_28710,N_28895);
nand U29410 (N_29410,N_28541,N_28545);
or U29411 (N_29411,N_28859,N_28887);
nor U29412 (N_29412,N_28686,N_28999);
or U29413 (N_29413,N_28963,N_28844);
or U29414 (N_29414,N_28663,N_28511);
xor U29415 (N_29415,N_28611,N_28862);
and U29416 (N_29416,N_28650,N_28672);
and U29417 (N_29417,N_28898,N_28518);
or U29418 (N_29418,N_28979,N_28600);
and U29419 (N_29419,N_28836,N_28912);
nand U29420 (N_29420,N_28775,N_28821);
xor U29421 (N_29421,N_28850,N_28717);
and U29422 (N_29422,N_28670,N_28588);
nand U29423 (N_29423,N_28666,N_28715);
xnor U29424 (N_29424,N_28855,N_28804);
nand U29425 (N_29425,N_28703,N_28848);
xor U29426 (N_29426,N_28863,N_28579);
nor U29427 (N_29427,N_28605,N_28614);
xnor U29428 (N_29428,N_28691,N_28737);
nand U29429 (N_29429,N_28574,N_28613);
nor U29430 (N_29430,N_28990,N_28647);
and U29431 (N_29431,N_28959,N_28609);
or U29432 (N_29432,N_28903,N_28908);
nand U29433 (N_29433,N_28885,N_28613);
nand U29434 (N_29434,N_28906,N_28853);
and U29435 (N_29435,N_28737,N_28754);
xor U29436 (N_29436,N_28975,N_28816);
nand U29437 (N_29437,N_28767,N_28796);
nor U29438 (N_29438,N_28564,N_28510);
nand U29439 (N_29439,N_28502,N_28560);
and U29440 (N_29440,N_28683,N_28561);
xor U29441 (N_29441,N_28621,N_28513);
xnor U29442 (N_29442,N_28633,N_28716);
nand U29443 (N_29443,N_28988,N_28915);
or U29444 (N_29444,N_28658,N_28821);
nand U29445 (N_29445,N_28765,N_28708);
or U29446 (N_29446,N_28503,N_28883);
nor U29447 (N_29447,N_28607,N_28760);
nor U29448 (N_29448,N_28813,N_28935);
nand U29449 (N_29449,N_28719,N_28795);
nand U29450 (N_29450,N_28856,N_28892);
nor U29451 (N_29451,N_28859,N_28511);
nor U29452 (N_29452,N_28628,N_28864);
xor U29453 (N_29453,N_28947,N_28714);
and U29454 (N_29454,N_28691,N_28940);
and U29455 (N_29455,N_28725,N_28809);
xnor U29456 (N_29456,N_28795,N_28559);
and U29457 (N_29457,N_28771,N_28990);
nor U29458 (N_29458,N_28751,N_28935);
nor U29459 (N_29459,N_28806,N_28972);
or U29460 (N_29460,N_28706,N_28858);
and U29461 (N_29461,N_28582,N_28551);
xor U29462 (N_29462,N_28977,N_28657);
nor U29463 (N_29463,N_28717,N_28995);
or U29464 (N_29464,N_28555,N_28785);
and U29465 (N_29465,N_28882,N_28934);
nand U29466 (N_29466,N_28853,N_28758);
nand U29467 (N_29467,N_28817,N_28750);
nand U29468 (N_29468,N_28724,N_28716);
nand U29469 (N_29469,N_28969,N_28853);
nand U29470 (N_29470,N_28762,N_28703);
or U29471 (N_29471,N_28973,N_28507);
and U29472 (N_29472,N_28658,N_28625);
and U29473 (N_29473,N_28903,N_28645);
and U29474 (N_29474,N_28833,N_28985);
or U29475 (N_29475,N_28648,N_28904);
xnor U29476 (N_29476,N_28837,N_28936);
nor U29477 (N_29477,N_28561,N_28965);
nor U29478 (N_29478,N_28632,N_28950);
and U29479 (N_29479,N_28923,N_28872);
and U29480 (N_29480,N_28954,N_28982);
xor U29481 (N_29481,N_28918,N_28922);
nand U29482 (N_29482,N_28691,N_28646);
and U29483 (N_29483,N_28670,N_28822);
nand U29484 (N_29484,N_28817,N_28871);
nor U29485 (N_29485,N_28820,N_28535);
and U29486 (N_29486,N_28952,N_28658);
nor U29487 (N_29487,N_28512,N_28945);
or U29488 (N_29488,N_28545,N_28792);
nand U29489 (N_29489,N_28889,N_28804);
nor U29490 (N_29490,N_28605,N_28856);
nand U29491 (N_29491,N_28673,N_28553);
nand U29492 (N_29492,N_28531,N_28852);
and U29493 (N_29493,N_28514,N_28704);
and U29494 (N_29494,N_28793,N_28680);
xnor U29495 (N_29495,N_28708,N_28760);
nor U29496 (N_29496,N_28782,N_28529);
nor U29497 (N_29497,N_28604,N_28597);
and U29498 (N_29498,N_28834,N_28889);
xor U29499 (N_29499,N_28647,N_28627);
or U29500 (N_29500,N_29140,N_29001);
nor U29501 (N_29501,N_29341,N_29136);
nand U29502 (N_29502,N_29375,N_29233);
xor U29503 (N_29503,N_29003,N_29293);
xnor U29504 (N_29504,N_29403,N_29456);
or U29505 (N_29505,N_29334,N_29498);
xnor U29506 (N_29506,N_29129,N_29213);
and U29507 (N_29507,N_29193,N_29066);
nor U29508 (N_29508,N_29306,N_29261);
or U29509 (N_29509,N_29362,N_29472);
or U29510 (N_29510,N_29385,N_29407);
nand U29511 (N_29511,N_29423,N_29182);
and U29512 (N_29512,N_29022,N_29455);
nor U29513 (N_29513,N_29286,N_29234);
nor U29514 (N_29514,N_29322,N_29390);
nand U29515 (N_29515,N_29368,N_29007);
nand U29516 (N_29516,N_29454,N_29283);
nand U29517 (N_29517,N_29161,N_29394);
and U29518 (N_29518,N_29443,N_29358);
nand U29519 (N_29519,N_29133,N_29298);
xnor U29520 (N_29520,N_29014,N_29131);
and U29521 (N_29521,N_29370,N_29388);
nand U29522 (N_29522,N_29119,N_29231);
and U29523 (N_29523,N_29300,N_29053);
nand U29524 (N_29524,N_29065,N_29484);
nor U29525 (N_29525,N_29093,N_29100);
and U29526 (N_29526,N_29062,N_29452);
nand U29527 (N_29527,N_29255,N_29372);
nand U29528 (N_29528,N_29139,N_29171);
or U29529 (N_29529,N_29052,N_29378);
or U29530 (N_29530,N_29288,N_29451);
and U29531 (N_29531,N_29246,N_29265);
nand U29532 (N_29532,N_29128,N_29389);
and U29533 (N_29533,N_29118,N_29312);
nor U29534 (N_29534,N_29252,N_29153);
nor U29535 (N_29535,N_29294,N_29225);
or U29536 (N_29536,N_29228,N_29215);
and U29537 (N_29537,N_29026,N_29258);
and U29538 (N_29538,N_29301,N_29488);
and U29539 (N_29539,N_29430,N_29256);
nor U29540 (N_29540,N_29167,N_29168);
or U29541 (N_29541,N_29427,N_29130);
or U29542 (N_29542,N_29369,N_29108);
nor U29543 (N_29543,N_29303,N_29075);
xnor U29544 (N_29544,N_29480,N_29479);
and U29545 (N_29545,N_29307,N_29146);
nor U29546 (N_29546,N_29400,N_29410);
and U29547 (N_29547,N_29332,N_29360);
nand U29548 (N_29548,N_29338,N_29240);
and U29549 (N_29549,N_29490,N_29132);
nor U29550 (N_29550,N_29395,N_29470);
or U29551 (N_29551,N_29273,N_29393);
nor U29552 (N_29552,N_29422,N_29416);
xnor U29553 (N_29553,N_29379,N_29235);
or U29554 (N_29554,N_29481,N_29012);
xnor U29555 (N_29555,N_29150,N_29177);
nand U29556 (N_29556,N_29381,N_29382);
and U29557 (N_29557,N_29267,N_29105);
nand U29558 (N_29558,N_29000,N_29324);
nand U29559 (N_29559,N_29323,N_29259);
and U29560 (N_29560,N_29226,N_29116);
and U29561 (N_29561,N_29084,N_29495);
or U29562 (N_29562,N_29325,N_29436);
xor U29563 (N_29563,N_29019,N_29018);
nor U29564 (N_29564,N_29309,N_29371);
and U29565 (N_29565,N_29328,N_29232);
or U29566 (N_29566,N_29173,N_29194);
and U29567 (N_29567,N_29056,N_29290);
xnor U29568 (N_29568,N_29098,N_29185);
and U29569 (N_29569,N_29079,N_29406);
xor U29570 (N_29570,N_29396,N_29186);
and U29571 (N_29571,N_29411,N_29178);
nor U29572 (N_29572,N_29155,N_29159);
and U29573 (N_29573,N_29114,N_29188);
nand U29574 (N_29574,N_29230,N_29376);
nand U29575 (N_29575,N_29117,N_29103);
nand U29576 (N_29576,N_29333,N_29189);
or U29577 (N_29577,N_29318,N_29450);
nor U29578 (N_29578,N_29096,N_29074);
or U29579 (N_29579,N_29275,N_29043);
nand U29580 (N_29580,N_29086,N_29200);
nor U29581 (N_29581,N_29239,N_29420);
or U29582 (N_29582,N_29070,N_29336);
or U29583 (N_29583,N_29181,N_29434);
and U29584 (N_29584,N_29424,N_29278);
nor U29585 (N_29585,N_29138,N_29072);
nand U29586 (N_29586,N_29080,N_29467);
and U29587 (N_29587,N_29216,N_29064);
nand U29588 (N_29588,N_29426,N_29435);
nor U29589 (N_29589,N_29489,N_29099);
xnor U29590 (N_29590,N_29089,N_29404);
xnor U29591 (N_29591,N_29243,N_29224);
xor U29592 (N_29592,N_29059,N_29359);
nor U29593 (N_29593,N_29269,N_29366);
nand U29594 (N_29594,N_29297,N_29095);
or U29595 (N_29595,N_29184,N_29448);
xnor U29596 (N_29596,N_29190,N_29260);
or U29597 (N_29597,N_29331,N_29041);
nor U29598 (N_29598,N_29262,N_29046);
or U29599 (N_29599,N_29081,N_29061);
and U29600 (N_29600,N_29463,N_29345);
or U29601 (N_29601,N_29045,N_29044);
xor U29602 (N_29602,N_29398,N_29414);
nor U29603 (N_29603,N_29157,N_29326);
and U29604 (N_29604,N_29485,N_29029);
nand U29605 (N_29605,N_29214,N_29280);
nor U29606 (N_29606,N_29152,N_29329);
nand U29607 (N_29607,N_29316,N_29060);
and U29608 (N_29608,N_29342,N_29164);
or U29609 (N_29609,N_29154,N_29284);
or U29610 (N_29610,N_29433,N_29349);
and U29611 (N_29611,N_29282,N_29471);
xnor U29612 (N_29612,N_29363,N_29257);
nor U29613 (N_29613,N_29149,N_29040);
and U29614 (N_29614,N_29109,N_29276);
nand U29615 (N_29615,N_29289,N_29440);
and U29616 (N_29616,N_29198,N_29077);
nand U29617 (N_29617,N_29206,N_29391);
nand U29618 (N_29618,N_29314,N_29175);
nand U29619 (N_29619,N_29217,N_29272);
xnor U29620 (N_29620,N_29346,N_29110);
and U29621 (N_29621,N_29068,N_29374);
xnor U29622 (N_29622,N_29067,N_29285);
or U29623 (N_29623,N_29158,N_29383);
xnor U29624 (N_29624,N_29445,N_29247);
or U29625 (N_29625,N_29348,N_29042);
and U29626 (N_29626,N_29361,N_29104);
and U29627 (N_29627,N_29458,N_29351);
or U29628 (N_29628,N_29251,N_29137);
nor U29629 (N_29629,N_29340,N_29085);
xor U29630 (N_29630,N_29250,N_29073);
and U29631 (N_29631,N_29237,N_29486);
nand U29632 (N_29632,N_29076,N_29199);
xnor U29633 (N_29633,N_29499,N_29475);
and U29634 (N_29634,N_29094,N_29425);
and U29635 (N_29635,N_29305,N_29187);
nand U29636 (N_29636,N_29446,N_29170);
nor U29637 (N_29637,N_29134,N_29373);
nand U29638 (N_29638,N_29429,N_29428);
nor U29639 (N_29639,N_29493,N_29017);
xor U29640 (N_29640,N_29219,N_29156);
and U29641 (N_29641,N_29277,N_29263);
nor U29642 (N_29642,N_29179,N_29028);
or U29643 (N_29643,N_29270,N_29241);
xor U29644 (N_29644,N_29048,N_29264);
nand U29645 (N_29645,N_29352,N_29102);
nor U29646 (N_29646,N_29036,N_29160);
or U29647 (N_29647,N_29421,N_29412);
nor U29648 (N_29648,N_29476,N_29483);
and U29649 (N_29649,N_29354,N_29055);
or U29650 (N_29650,N_29032,N_29191);
or U29651 (N_29651,N_29350,N_29165);
xor U29652 (N_29652,N_29208,N_29419);
and U29653 (N_29653,N_29209,N_29169);
and U29654 (N_29654,N_29405,N_29365);
or U29655 (N_29655,N_29266,N_29002);
nand U29656 (N_29656,N_29166,N_29296);
and U29657 (N_29657,N_29466,N_29311);
or U29658 (N_29658,N_29218,N_29111);
nor U29659 (N_29659,N_29092,N_29386);
or U29660 (N_29660,N_29457,N_29431);
and U29661 (N_29661,N_29008,N_29088);
nor U29662 (N_29662,N_29050,N_29281);
and U29663 (N_29663,N_29313,N_29006);
xor U29664 (N_29664,N_29172,N_29473);
nand U29665 (N_29665,N_29027,N_29401);
xor U29666 (N_29666,N_29229,N_29034);
and U29667 (N_29667,N_29245,N_29364);
xnor U29668 (N_29668,N_29024,N_29151);
nor U29669 (N_29669,N_29207,N_29377);
or U29670 (N_29670,N_29020,N_29091);
nand U29671 (N_29671,N_29437,N_29121);
or U29672 (N_29672,N_29384,N_29078);
or U29673 (N_29673,N_29087,N_29183);
or U29674 (N_29674,N_29248,N_29442);
or U29675 (N_29675,N_29477,N_29063);
xor U29676 (N_29676,N_29271,N_29347);
and U29677 (N_29677,N_29005,N_29465);
or U29678 (N_29678,N_29071,N_29144);
nand U29679 (N_29679,N_29126,N_29037);
or U29680 (N_29680,N_29021,N_29195);
or U29681 (N_29681,N_29143,N_29176);
nor U29682 (N_29682,N_29492,N_29353);
or U29683 (N_29683,N_29025,N_29106);
nand U29684 (N_29684,N_29221,N_29462);
and U29685 (N_29685,N_29212,N_29009);
nor U29686 (N_29686,N_29013,N_29120);
nor U29687 (N_29687,N_29344,N_29315);
and U29688 (N_29688,N_29474,N_29011);
xnor U29689 (N_29689,N_29201,N_29447);
and U29690 (N_29690,N_29279,N_29337);
nor U29691 (N_29691,N_29469,N_29295);
and U29692 (N_29692,N_29030,N_29090);
nand U29693 (N_29693,N_29461,N_29408);
nor U29694 (N_29694,N_29380,N_29418);
xor U29695 (N_29695,N_29222,N_29432);
nor U29696 (N_29696,N_29319,N_29339);
and U29697 (N_29697,N_29453,N_29039);
nand U29698 (N_29698,N_29491,N_29254);
or U29699 (N_29699,N_29327,N_29335);
xnor U29700 (N_29700,N_29197,N_29417);
and U29701 (N_29701,N_29127,N_29253);
and U29702 (N_29702,N_29497,N_29141);
or U29703 (N_29703,N_29399,N_29274);
and U29704 (N_29704,N_29242,N_29478);
and U29705 (N_29705,N_29082,N_29115);
nor U29706 (N_29706,N_29460,N_29268);
nor U29707 (N_29707,N_29392,N_29023);
xnor U29708 (N_29708,N_29049,N_29449);
and U29709 (N_29709,N_29205,N_29220);
and U29710 (N_29710,N_29145,N_29125);
xnor U29711 (N_29711,N_29202,N_29142);
xnor U29712 (N_29712,N_29054,N_29482);
xor U29713 (N_29713,N_29464,N_29174);
or U29714 (N_29714,N_29236,N_29097);
xor U29715 (N_29715,N_29387,N_29238);
nor U29716 (N_29716,N_29180,N_29192);
and U29717 (N_29717,N_29163,N_29302);
or U29718 (N_29718,N_29402,N_29494);
nor U29719 (N_29719,N_29101,N_29162);
and U29720 (N_29720,N_29122,N_29304);
and U29721 (N_29721,N_29148,N_29038);
nand U29722 (N_29722,N_29147,N_29413);
or U29723 (N_29723,N_29468,N_29310);
or U29724 (N_29724,N_29397,N_29069);
xnor U29725 (N_29725,N_29496,N_29010);
and U29726 (N_29726,N_29244,N_29107);
or U29727 (N_29727,N_29343,N_29223);
nor U29728 (N_29728,N_29015,N_29033);
xor U29729 (N_29729,N_29057,N_29367);
nor U29730 (N_29730,N_29459,N_29320);
nand U29731 (N_29731,N_29196,N_29356);
and U29732 (N_29732,N_29355,N_29083);
and U29733 (N_29733,N_29249,N_29287);
nand U29734 (N_29734,N_29210,N_29438);
or U29735 (N_29735,N_29439,N_29047);
nor U29736 (N_29736,N_29357,N_29444);
and U29737 (N_29737,N_29035,N_29123);
or U29738 (N_29738,N_29415,N_29227);
and U29739 (N_29739,N_29051,N_29211);
and U29740 (N_29740,N_29330,N_29203);
nor U29741 (N_29741,N_29291,N_29016);
and U29742 (N_29742,N_29292,N_29204);
or U29743 (N_29743,N_29409,N_29487);
nor U29744 (N_29744,N_29112,N_29317);
nand U29745 (N_29745,N_29058,N_29321);
or U29746 (N_29746,N_29124,N_29113);
xnor U29747 (N_29747,N_29308,N_29135);
nor U29748 (N_29748,N_29004,N_29031);
and U29749 (N_29749,N_29441,N_29299);
nand U29750 (N_29750,N_29206,N_29290);
or U29751 (N_29751,N_29289,N_29068);
or U29752 (N_29752,N_29263,N_29049);
nor U29753 (N_29753,N_29261,N_29332);
nand U29754 (N_29754,N_29443,N_29451);
and U29755 (N_29755,N_29151,N_29085);
or U29756 (N_29756,N_29261,N_29293);
and U29757 (N_29757,N_29357,N_29347);
xor U29758 (N_29758,N_29339,N_29446);
xor U29759 (N_29759,N_29243,N_29303);
nand U29760 (N_29760,N_29307,N_29293);
xor U29761 (N_29761,N_29010,N_29431);
nor U29762 (N_29762,N_29441,N_29022);
nand U29763 (N_29763,N_29142,N_29264);
or U29764 (N_29764,N_29112,N_29332);
xnor U29765 (N_29765,N_29243,N_29327);
xnor U29766 (N_29766,N_29020,N_29072);
nand U29767 (N_29767,N_29364,N_29131);
xnor U29768 (N_29768,N_29080,N_29060);
xor U29769 (N_29769,N_29239,N_29181);
or U29770 (N_29770,N_29084,N_29422);
or U29771 (N_29771,N_29395,N_29054);
and U29772 (N_29772,N_29089,N_29027);
nor U29773 (N_29773,N_29265,N_29352);
and U29774 (N_29774,N_29065,N_29101);
xor U29775 (N_29775,N_29358,N_29252);
and U29776 (N_29776,N_29362,N_29231);
or U29777 (N_29777,N_29456,N_29173);
nand U29778 (N_29778,N_29382,N_29207);
nor U29779 (N_29779,N_29117,N_29359);
nand U29780 (N_29780,N_29104,N_29156);
nor U29781 (N_29781,N_29457,N_29241);
or U29782 (N_29782,N_29478,N_29338);
and U29783 (N_29783,N_29361,N_29373);
and U29784 (N_29784,N_29173,N_29202);
nand U29785 (N_29785,N_29446,N_29350);
nor U29786 (N_29786,N_29056,N_29340);
and U29787 (N_29787,N_29332,N_29036);
nand U29788 (N_29788,N_29412,N_29175);
or U29789 (N_29789,N_29095,N_29078);
nor U29790 (N_29790,N_29012,N_29377);
nand U29791 (N_29791,N_29475,N_29381);
and U29792 (N_29792,N_29330,N_29461);
nand U29793 (N_29793,N_29297,N_29467);
or U29794 (N_29794,N_29035,N_29225);
nand U29795 (N_29795,N_29267,N_29238);
nand U29796 (N_29796,N_29219,N_29492);
xnor U29797 (N_29797,N_29014,N_29160);
and U29798 (N_29798,N_29219,N_29079);
xor U29799 (N_29799,N_29420,N_29373);
or U29800 (N_29800,N_29289,N_29305);
nor U29801 (N_29801,N_29044,N_29453);
xnor U29802 (N_29802,N_29256,N_29384);
and U29803 (N_29803,N_29412,N_29234);
nor U29804 (N_29804,N_29454,N_29233);
and U29805 (N_29805,N_29371,N_29314);
and U29806 (N_29806,N_29340,N_29183);
xor U29807 (N_29807,N_29477,N_29114);
nand U29808 (N_29808,N_29030,N_29024);
nand U29809 (N_29809,N_29005,N_29463);
nand U29810 (N_29810,N_29036,N_29100);
nor U29811 (N_29811,N_29218,N_29153);
and U29812 (N_29812,N_29023,N_29340);
nand U29813 (N_29813,N_29102,N_29170);
nor U29814 (N_29814,N_29212,N_29306);
xor U29815 (N_29815,N_29232,N_29355);
xor U29816 (N_29816,N_29077,N_29052);
xnor U29817 (N_29817,N_29175,N_29453);
or U29818 (N_29818,N_29342,N_29269);
or U29819 (N_29819,N_29210,N_29218);
nor U29820 (N_29820,N_29088,N_29152);
xor U29821 (N_29821,N_29356,N_29033);
or U29822 (N_29822,N_29066,N_29441);
or U29823 (N_29823,N_29328,N_29015);
nand U29824 (N_29824,N_29204,N_29105);
or U29825 (N_29825,N_29469,N_29044);
xnor U29826 (N_29826,N_29340,N_29052);
xnor U29827 (N_29827,N_29065,N_29050);
nor U29828 (N_29828,N_29248,N_29450);
nor U29829 (N_29829,N_29243,N_29006);
nor U29830 (N_29830,N_29377,N_29147);
and U29831 (N_29831,N_29108,N_29281);
or U29832 (N_29832,N_29096,N_29109);
nor U29833 (N_29833,N_29382,N_29054);
nor U29834 (N_29834,N_29016,N_29112);
nand U29835 (N_29835,N_29084,N_29114);
xnor U29836 (N_29836,N_29292,N_29138);
nand U29837 (N_29837,N_29108,N_29312);
nand U29838 (N_29838,N_29117,N_29459);
or U29839 (N_29839,N_29102,N_29069);
or U29840 (N_29840,N_29004,N_29471);
nor U29841 (N_29841,N_29155,N_29402);
xor U29842 (N_29842,N_29275,N_29111);
and U29843 (N_29843,N_29376,N_29359);
and U29844 (N_29844,N_29200,N_29133);
nor U29845 (N_29845,N_29048,N_29141);
and U29846 (N_29846,N_29058,N_29161);
nor U29847 (N_29847,N_29305,N_29369);
nor U29848 (N_29848,N_29403,N_29378);
and U29849 (N_29849,N_29411,N_29436);
and U29850 (N_29850,N_29300,N_29387);
and U29851 (N_29851,N_29148,N_29104);
or U29852 (N_29852,N_29396,N_29286);
or U29853 (N_29853,N_29285,N_29186);
and U29854 (N_29854,N_29304,N_29272);
xor U29855 (N_29855,N_29038,N_29412);
or U29856 (N_29856,N_29089,N_29038);
or U29857 (N_29857,N_29459,N_29172);
xor U29858 (N_29858,N_29060,N_29365);
and U29859 (N_29859,N_29343,N_29485);
or U29860 (N_29860,N_29221,N_29274);
nor U29861 (N_29861,N_29391,N_29483);
and U29862 (N_29862,N_29427,N_29206);
nor U29863 (N_29863,N_29037,N_29208);
xor U29864 (N_29864,N_29068,N_29444);
xnor U29865 (N_29865,N_29049,N_29305);
nor U29866 (N_29866,N_29311,N_29359);
and U29867 (N_29867,N_29342,N_29327);
nor U29868 (N_29868,N_29484,N_29191);
nor U29869 (N_29869,N_29427,N_29399);
xor U29870 (N_29870,N_29049,N_29346);
nor U29871 (N_29871,N_29061,N_29477);
or U29872 (N_29872,N_29445,N_29115);
and U29873 (N_29873,N_29285,N_29393);
and U29874 (N_29874,N_29353,N_29469);
and U29875 (N_29875,N_29300,N_29196);
nor U29876 (N_29876,N_29286,N_29388);
nor U29877 (N_29877,N_29205,N_29204);
nor U29878 (N_29878,N_29347,N_29317);
and U29879 (N_29879,N_29123,N_29436);
xnor U29880 (N_29880,N_29205,N_29461);
xor U29881 (N_29881,N_29397,N_29135);
nor U29882 (N_29882,N_29113,N_29175);
nor U29883 (N_29883,N_29311,N_29102);
xor U29884 (N_29884,N_29133,N_29093);
or U29885 (N_29885,N_29017,N_29426);
nor U29886 (N_29886,N_29021,N_29361);
nand U29887 (N_29887,N_29300,N_29212);
nor U29888 (N_29888,N_29498,N_29149);
nor U29889 (N_29889,N_29051,N_29150);
xnor U29890 (N_29890,N_29249,N_29198);
or U29891 (N_29891,N_29265,N_29262);
nor U29892 (N_29892,N_29274,N_29047);
xnor U29893 (N_29893,N_29154,N_29226);
nor U29894 (N_29894,N_29178,N_29234);
or U29895 (N_29895,N_29406,N_29060);
nand U29896 (N_29896,N_29262,N_29014);
nor U29897 (N_29897,N_29395,N_29401);
or U29898 (N_29898,N_29494,N_29268);
and U29899 (N_29899,N_29039,N_29321);
or U29900 (N_29900,N_29220,N_29273);
and U29901 (N_29901,N_29057,N_29261);
xnor U29902 (N_29902,N_29001,N_29127);
and U29903 (N_29903,N_29304,N_29395);
nand U29904 (N_29904,N_29411,N_29306);
nor U29905 (N_29905,N_29124,N_29375);
and U29906 (N_29906,N_29083,N_29164);
nor U29907 (N_29907,N_29137,N_29209);
nand U29908 (N_29908,N_29059,N_29456);
nand U29909 (N_29909,N_29491,N_29175);
xnor U29910 (N_29910,N_29234,N_29334);
nor U29911 (N_29911,N_29476,N_29337);
xnor U29912 (N_29912,N_29332,N_29162);
nor U29913 (N_29913,N_29368,N_29499);
nand U29914 (N_29914,N_29416,N_29045);
nor U29915 (N_29915,N_29304,N_29283);
nor U29916 (N_29916,N_29072,N_29198);
xnor U29917 (N_29917,N_29432,N_29164);
and U29918 (N_29918,N_29463,N_29021);
and U29919 (N_29919,N_29027,N_29271);
xor U29920 (N_29920,N_29074,N_29198);
and U29921 (N_29921,N_29044,N_29317);
and U29922 (N_29922,N_29446,N_29319);
and U29923 (N_29923,N_29228,N_29065);
and U29924 (N_29924,N_29428,N_29198);
and U29925 (N_29925,N_29041,N_29116);
nand U29926 (N_29926,N_29244,N_29111);
and U29927 (N_29927,N_29131,N_29182);
nor U29928 (N_29928,N_29114,N_29015);
and U29929 (N_29929,N_29089,N_29361);
and U29930 (N_29930,N_29492,N_29068);
and U29931 (N_29931,N_29091,N_29224);
or U29932 (N_29932,N_29471,N_29120);
or U29933 (N_29933,N_29134,N_29362);
or U29934 (N_29934,N_29102,N_29049);
and U29935 (N_29935,N_29193,N_29077);
and U29936 (N_29936,N_29288,N_29487);
and U29937 (N_29937,N_29069,N_29477);
nand U29938 (N_29938,N_29000,N_29378);
and U29939 (N_29939,N_29170,N_29361);
nand U29940 (N_29940,N_29481,N_29406);
xnor U29941 (N_29941,N_29151,N_29051);
or U29942 (N_29942,N_29463,N_29161);
nand U29943 (N_29943,N_29307,N_29338);
and U29944 (N_29944,N_29357,N_29160);
and U29945 (N_29945,N_29134,N_29273);
nor U29946 (N_29946,N_29064,N_29386);
nand U29947 (N_29947,N_29344,N_29288);
or U29948 (N_29948,N_29042,N_29073);
and U29949 (N_29949,N_29292,N_29305);
or U29950 (N_29950,N_29062,N_29408);
nor U29951 (N_29951,N_29189,N_29159);
nand U29952 (N_29952,N_29389,N_29156);
nor U29953 (N_29953,N_29237,N_29089);
xor U29954 (N_29954,N_29062,N_29085);
or U29955 (N_29955,N_29431,N_29425);
nand U29956 (N_29956,N_29358,N_29102);
or U29957 (N_29957,N_29168,N_29411);
and U29958 (N_29958,N_29086,N_29106);
nand U29959 (N_29959,N_29151,N_29073);
or U29960 (N_29960,N_29076,N_29447);
xor U29961 (N_29961,N_29237,N_29298);
or U29962 (N_29962,N_29018,N_29130);
nor U29963 (N_29963,N_29016,N_29445);
nand U29964 (N_29964,N_29061,N_29402);
or U29965 (N_29965,N_29020,N_29302);
nor U29966 (N_29966,N_29487,N_29166);
nand U29967 (N_29967,N_29413,N_29090);
or U29968 (N_29968,N_29284,N_29229);
or U29969 (N_29969,N_29154,N_29242);
nand U29970 (N_29970,N_29283,N_29099);
nor U29971 (N_29971,N_29292,N_29387);
or U29972 (N_29972,N_29226,N_29206);
nor U29973 (N_29973,N_29311,N_29443);
xor U29974 (N_29974,N_29146,N_29026);
and U29975 (N_29975,N_29339,N_29035);
and U29976 (N_29976,N_29082,N_29422);
nand U29977 (N_29977,N_29391,N_29035);
nand U29978 (N_29978,N_29353,N_29016);
nand U29979 (N_29979,N_29494,N_29393);
or U29980 (N_29980,N_29445,N_29051);
nor U29981 (N_29981,N_29367,N_29074);
and U29982 (N_29982,N_29103,N_29414);
nand U29983 (N_29983,N_29406,N_29280);
nor U29984 (N_29984,N_29204,N_29303);
nand U29985 (N_29985,N_29274,N_29406);
nor U29986 (N_29986,N_29389,N_29086);
and U29987 (N_29987,N_29050,N_29449);
xor U29988 (N_29988,N_29197,N_29173);
xor U29989 (N_29989,N_29482,N_29323);
nor U29990 (N_29990,N_29014,N_29052);
xor U29991 (N_29991,N_29218,N_29278);
xnor U29992 (N_29992,N_29084,N_29135);
or U29993 (N_29993,N_29476,N_29022);
or U29994 (N_29994,N_29322,N_29336);
xnor U29995 (N_29995,N_29459,N_29072);
xor U29996 (N_29996,N_29304,N_29113);
or U29997 (N_29997,N_29012,N_29301);
or U29998 (N_29998,N_29114,N_29017);
and U29999 (N_29999,N_29002,N_29440);
or U30000 (N_30000,N_29760,N_29691);
and U30001 (N_30001,N_29692,N_29716);
or U30002 (N_30002,N_29801,N_29891);
or U30003 (N_30003,N_29941,N_29738);
and U30004 (N_30004,N_29638,N_29615);
or U30005 (N_30005,N_29773,N_29748);
nand U30006 (N_30006,N_29988,N_29602);
nor U30007 (N_30007,N_29528,N_29839);
and U30008 (N_30008,N_29882,N_29531);
xor U30009 (N_30009,N_29996,N_29858);
or U30010 (N_30010,N_29823,N_29969);
xor U30011 (N_30011,N_29681,N_29919);
xor U30012 (N_30012,N_29982,N_29902);
nand U30013 (N_30013,N_29943,N_29699);
nand U30014 (N_30014,N_29763,N_29893);
xor U30015 (N_30015,N_29625,N_29974);
nand U30016 (N_30016,N_29875,N_29755);
and U30017 (N_30017,N_29872,N_29605);
and U30018 (N_30018,N_29607,N_29568);
nand U30019 (N_30019,N_29684,N_29787);
xnor U30020 (N_30020,N_29851,N_29733);
nand U30021 (N_30021,N_29689,N_29912);
nand U30022 (N_30022,N_29965,N_29961);
or U30023 (N_30023,N_29778,N_29598);
nor U30024 (N_30024,N_29546,N_29599);
and U30025 (N_30025,N_29987,N_29523);
xnor U30026 (N_30026,N_29509,N_29795);
or U30027 (N_30027,N_29620,N_29517);
and U30028 (N_30028,N_29832,N_29890);
nor U30029 (N_30029,N_29928,N_29861);
and U30030 (N_30030,N_29767,N_29967);
and U30031 (N_30031,N_29871,N_29572);
nor U30032 (N_30032,N_29925,N_29538);
nor U30033 (N_30033,N_29551,N_29588);
xnor U30034 (N_30034,N_29918,N_29934);
or U30035 (N_30035,N_29597,N_29563);
or U30036 (N_30036,N_29808,N_29734);
and U30037 (N_30037,N_29603,N_29537);
xor U30038 (N_30038,N_29993,N_29533);
or U30039 (N_30039,N_29582,N_29897);
or U30040 (N_30040,N_29717,N_29975);
xnor U30041 (N_30041,N_29885,N_29736);
or U30042 (N_30042,N_29707,N_29990);
xnor U30043 (N_30043,N_29814,N_29848);
and U30044 (N_30044,N_29650,N_29953);
and U30045 (N_30045,N_29589,N_29973);
xor U30046 (N_30046,N_29878,N_29593);
xor U30047 (N_30047,N_29504,N_29566);
nand U30048 (N_30048,N_29571,N_29962);
and U30049 (N_30049,N_29892,N_29732);
nor U30050 (N_30050,N_29741,N_29570);
nand U30051 (N_30051,N_29718,N_29849);
nor U30052 (N_30052,N_29610,N_29830);
xnor U30053 (N_30053,N_29989,N_29527);
nand U30054 (N_30054,N_29754,N_29797);
nor U30055 (N_30055,N_29560,N_29781);
xnor U30056 (N_30056,N_29826,N_29735);
and U30057 (N_30057,N_29894,N_29581);
and U30058 (N_30058,N_29929,N_29578);
and U30059 (N_30059,N_29654,N_29970);
or U30060 (N_30060,N_29617,N_29668);
and U30061 (N_30061,N_29793,N_29909);
and U30062 (N_30062,N_29661,N_29824);
nand U30063 (N_30063,N_29916,N_29591);
and U30064 (N_30064,N_29514,N_29626);
and U30065 (N_30065,N_29653,N_29991);
nor U30066 (N_30066,N_29583,N_29715);
and U30067 (N_30067,N_29776,N_29536);
xor U30068 (N_30068,N_29652,N_29587);
or U30069 (N_30069,N_29696,N_29519);
xor U30070 (N_30070,N_29633,N_29976);
and U30071 (N_30071,N_29868,N_29992);
nand U30072 (N_30072,N_29812,N_29827);
or U30073 (N_30073,N_29769,N_29933);
xor U30074 (N_30074,N_29917,N_29765);
nor U30075 (N_30075,N_29695,N_29980);
or U30076 (N_30076,N_29694,N_29543);
nand U30077 (N_30077,N_29883,N_29835);
nand U30078 (N_30078,N_29688,N_29983);
and U30079 (N_30079,N_29792,N_29977);
nand U30080 (N_30080,N_29512,N_29511);
and U30081 (N_30081,N_29687,N_29667);
and U30082 (N_30082,N_29880,N_29922);
nand U30083 (N_30083,N_29942,N_29771);
and U30084 (N_30084,N_29518,N_29960);
and U30085 (N_30085,N_29567,N_29646);
nor U30086 (N_30086,N_29639,N_29714);
or U30087 (N_30087,N_29746,N_29674);
and U30088 (N_30088,N_29539,N_29958);
xor U30089 (N_30089,N_29817,N_29540);
nor U30090 (N_30090,N_29936,N_29752);
or U30091 (N_30091,N_29630,N_29606);
nand U30092 (N_30092,N_29998,N_29595);
nand U30093 (N_30093,N_29686,N_29800);
or U30094 (N_30094,N_29818,N_29678);
or U30095 (N_30095,N_29949,N_29784);
xnor U30096 (N_30096,N_29986,N_29863);
or U30097 (N_30097,N_29621,N_29867);
nor U30098 (N_30098,N_29618,N_29683);
nand U30099 (N_30099,N_29864,N_29997);
nand U30100 (N_30100,N_29665,N_29641);
xnor U30101 (N_30101,N_29939,N_29899);
and U30102 (N_30102,N_29901,N_29904);
xor U30103 (N_30103,N_29815,N_29783);
nor U30104 (N_30104,N_29500,N_29915);
xnor U30105 (N_30105,N_29505,N_29666);
and U30106 (N_30106,N_29931,N_29676);
or U30107 (N_30107,N_29802,N_29833);
nor U30108 (N_30108,N_29999,N_29542);
xor U30109 (N_30109,N_29657,N_29644);
nand U30110 (N_30110,N_29836,N_29782);
nor U30111 (N_30111,N_29921,N_29898);
and U30112 (N_30112,N_29722,N_29723);
or U30113 (N_30113,N_29645,N_29766);
xnor U30114 (N_30114,N_29556,N_29558);
nor U30115 (N_30115,N_29649,N_29825);
nand U30116 (N_30116,N_29959,N_29788);
or U30117 (N_30117,N_29865,N_29955);
xnor U30118 (N_30118,N_29946,N_29576);
and U30119 (N_30119,N_29614,N_29786);
nor U30120 (N_30120,N_29554,N_29747);
or U30121 (N_30121,N_29724,N_29907);
nand U30122 (N_30122,N_29790,N_29577);
or U30123 (N_30123,N_29995,N_29524);
nor U30124 (N_30124,N_29662,N_29697);
and U30125 (N_30125,N_29937,N_29503);
and U30126 (N_30126,N_29711,N_29940);
or U30127 (N_30127,N_29643,N_29580);
or U30128 (N_30128,N_29777,N_29561);
xnor U30129 (N_30129,N_29804,N_29710);
nor U30130 (N_30130,N_29908,N_29809);
nand U30131 (N_30131,N_29856,N_29612);
nand U30132 (N_30132,N_29900,N_29821);
and U30133 (N_30133,N_29544,N_29964);
or U30134 (N_30134,N_29552,N_29770);
xor U30135 (N_30135,N_29834,N_29966);
xnor U30136 (N_30136,N_29515,N_29660);
and U30137 (N_30137,N_29706,N_29506);
or U30138 (N_30138,N_29669,N_29664);
or U30139 (N_30139,N_29640,N_29742);
nor U30140 (N_30140,N_29859,N_29642);
nand U30141 (N_30141,N_29550,N_29564);
xor U30142 (N_30142,N_29535,N_29870);
and U30143 (N_30143,N_29957,N_29753);
nor U30144 (N_30144,N_29651,N_29762);
xor U30145 (N_30145,N_29829,N_29682);
xnor U30146 (N_30146,N_29884,N_29726);
nor U30147 (N_30147,N_29629,N_29616);
or U30148 (N_30148,N_29575,N_29844);
or U30149 (N_30149,N_29927,N_29796);
nand U30150 (N_30150,N_29545,N_29850);
or U30151 (N_30151,N_29789,N_29948);
nor U30152 (N_30152,N_29979,N_29613);
xor U30153 (N_30153,N_29702,N_29843);
nor U30154 (N_30154,N_29530,N_29520);
or U30155 (N_30155,N_29635,N_29888);
xor U30156 (N_30156,N_29985,N_29529);
nor U30157 (N_30157,N_29508,N_29584);
nand U30158 (N_30158,N_29585,N_29764);
nor U30159 (N_30159,N_29775,N_29785);
and U30160 (N_30160,N_29932,N_29952);
and U30161 (N_30161,N_29590,N_29648);
and U30162 (N_30162,N_29994,N_29659);
and U30163 (N_30163,N_29586,N_29761);
and U30164 (N_30164,N_29920,N_29751);
and U30165 (N_30165,N_29728,N_29956);
and U30166 (N_30166,N_29548,N_29963);
or U30167 (N_30167,N_29604,N_29935);
nor U30168 (N_30168,N_29516,N_29816);
nand U30169 (N_30169,N_29675,N_29737);
or U30170 (N_30170,N_29914,N_29522);
nand U30171 (N_30171,N_29806,N_29779);
and U30172 (N_30172,N_29938,N_29820);
nor U30173 (N_30173,N_29525,N_29739);
nand U30174 (N_30174,N_29947,N_29768);
nor U30175 (N_30175,N_29709,N_29951);
xnor U30176 (N_30176,N_29670,N_29805);
or U30177 (N_30177,N_29549,N_29831);
xor U30178 (N_30178,N_29950,N_29624);
xnor U30179 (N_30179,N_29924,N_29611);
or U30180 (N_30180,N_29592,N_29693);
nor U30181 (N_30181,N_29877,N_29690);
nand U30182 (N_30182,N_29876,N_29534);
xnor U30183 (N_30183,N_29730,N_29622);
or U30184 (N_30184,N_29559,N_29807);
nor U30185 (N_30185,N_29672,N_29923);
nor U30186 (N_30186,N_29757,N_29698);
and U30187 (N_30187,N_29944,N_29532);
or U30188 (N_30188,N_29842,N_29813);
and U30189 (N_30189,N_29526,N_29634);
nor U30190 (N_30190,N_29811,N_29886);
nand U30191 (N_30191,N_29862,N_29565);
or U30192 (N_30192,N_29743,N_29846);
nor U30193 (N_30193,N_29853,N_29573);
and U30194 (N_30194,N_29700,N_29896);
nand U30195 (N_30195,N_29708,N_29874);
nand U30196 (N_30196,N_29873,N_29838);
or U30197 (N_30197,N_29574,N_29895);
nand U30198 (N_30198,N_29841,N_29889);
and U30199 (N_30199,N_29745,N_29930);
or U30200 (N_30200,N_29758,N_29673);
nor U30201 (N_30201,N_29855,N_29513);
nor U30202 (N_30202,N_29507,N_29647);
nor U30203 (N_30203,N_29596,N_29803);
nand U30204 (N_30204,N_29601,N_29954);
xnor U30205 (N_30205,N_29866,N_29852);
xnor U30206 (N_30206,N_29671,N_29677);
or U30207 (N_30207,N_29911,N_29981);
and U30208 (N_30208,N_29719,N_29984);
xnor U30209 (N_30209,N_29562,N_29740);
xor U30210 (N_30210,N_29972,N_29600);
and U30211 (N_30211,N_29854,N_29663);
xor U30212 (N_30212,N_29685,N_29627);
nand U30213 (N_30213,N_29623,N_29679);
and U30214 (N_30214,N_29656,N_29869);
or U30215 (N_30215,N_29791,N_29501);
xor U30216 (N_30216,N_29720,N_29798);
xnor U30217 (N_30217,N_29705,N_29594);
nand U30218 (N_30218,N_29968,N_29541);
nor U30219 (N_30219,N_29701,N_29799);
xor U30220 (N_30220,N_29502,N_29780);
nor U30221 (N_30221,N_29636,N_29978);
or U30222 (N_30222,N_29905,N_29727);
and U30223 (N_30223,N_29712,N_29756);
nor U30224 (N_30224,N_29658,N_29631);
or U30225 (N_30225,N_29655,N_29608);
and U30226 (N_30226,N_29731,N_29774);
nor U30227 (N_30227,N_29680,N_29819);
and U30228 (N_30228,N_29750,N_29510);
nor U30229 (N_30229,N_29794,N_29632);
nand U30230 (N_30230,N_29713,N_29637);
nor U30231 (N_30231,N_29860,N_29971);
nor U30232 (N_30232,N_29569,N_29879);
and U30233 (N_30233,N_29845,N_29619);
xnor U30234 (N_30234,N_29926,N_29945);
nand U30235 (N_30235,N_29557,N_29759);
xor U30236 (N_30236,N_29521,N_29721);
and U30237 (N_30237,N_29628,N_29725);
or U30238 (N_30238,N_29744,N_29772);
or U30239 (N_30239,N_29609,N_29857);
or U30240 (N_30240,N_29903,N_29703);
nor U30241 (N_30241,N_29837,N_29840);
and U30242 (N_30242,N_29906,N_29887);
and U30243 (N_30243,N_29749,N_29828);
or U30244 (N_30244,N_29704,N_29910);
and U30245 (N_30245,N_29822,N_29555);
nor U30246 (N_30246,N_29729,N_29547);
or U30247 (N_30247,N_29913,N_29810);
and U30248 (N_30248,N_29579,N_29847);
nor U30249 (N_30249,N_29553,N_29881);
nand U30250 (N_30250,N_29645,N_29588);
nor U30251 (N_30251,N_29779,N_29841);
and U30252 (N_30252,N_29900,N_29667);
and U30253 (N_30253,N_29775,N_29928);
xor U30254 (N_30254,N_29765,N_29507);
nor U30255 (N_30255,N_29972,N_29654);
nand U30256 (N_30256,N_29858,N_29706);
nor U30257 (N_30257,N_29913,N_29624);
xor U30258 (N_30258,N_29594,N_29831);
nor U30259 (N_30259,N_29560,N_29710);
nor U30260 (N_30260,N_29587,N_29730);
and U30261 (N_30261,N_29690,N_29516);
nor U30262 (N_30262,N_29919,N_29753);
xor U30263 (N_30263,N_29550,N_29809);
xor U30264 (N_30264,N_29510,N_29620);
nor U30265 (N_30265,N_29989,N_29983);
or U30266 (N_30266,N_29921,N_29674);
xnor U30267 (N_30267,N_29584,N_29501);
nor U30268 (N_30268,N_29811,N_29527);
and U30269 (N_30269,N_29650,N_29739);
xor U30270 (N_30270,N_29813,N_29834);
and U30271 (N_30271,N_29739,N_29952);
or U30272 (N_30272,N_29635,N_29742);
and U30273 (N_30273,N_29520,N_29719);
and U30274 (N_30274,N_29594,N_29573);
or U30275 (N_30275,N_29690,N_29853);
xnor U30276 (N_30276,N_29527,N_29792);
nor U30277 (N_30277,N_29964,N_29723);
nor U30278 (N_30278,N_29731,N_29889);
nand U30279 (N_30279,N_29591,N_29778);
or U30280 (N_30280,N_29899,N_29880);
nor U30281 (N_30281,N_29893,N_29949);
xor U30282 (N_30282,N_29943,N_29876);
nand U30283 (N_30283,N_29630,N_29830);
or U30284 (N_30284,N_29747,N_29782);
nor U30285 (N_30285,N_29877,N_29735);
xnor U30286 (N_30286,N_29736,N_29800);
xnor U30287 (N_30287,N_29853,N_29729);
and U30288 (N_30288,N_29522,N_29549);
nor U30289 (N_30289,N_29769,N_29711);
nand U30290 (N_30290,N_29516,N_29812);
and U30291 (N_30291,N_29986,N_29928);
nand U30292 (N_30292,N_29630,N_29664);
xor U30293 (N_30293,N_29841,N_29859);
or U30294 (N_30294,N_29598,N_29642);
and U30295 (N_30295,N_29768,N_29652);
nand U30296 (N_30296,N_29661,N_29615);
or U30297 (N_30297,N_29764,N_29852);
and U30298 (N_30298,N_29811,N_29723);
or U30299 (N_30299,N_29872,N_29700);
and U30300 (N_30300,N_29523,N_29625);
xnor U30301 (N_30301,N_29532,N_29561);
or U30302 (N_30302,N_29632,N_29842);
nand U30303 (N_30303,N_29735,N_29535);
xor U30304 (N_30304,N_29983,N_29930);
xnor U30305 (N_30305,N_29676,N_29845);
and U30306 (N_30306,N_29504,N_29890);
or U30307 (N_30307,N_29509,N_29546);
xnor U30308 (N_30308,N_29911,N_29861);
nor U30309 (N_30309,N_29660,N_29597);
nand U30310 (N_30310,N_29776,N_29963);
and U30311 (N_30311,N_29845,N_29888);
xor U30312 (N_30312,N_29954,N_29593);
xnor U30313 (N_30313,N_29917,N_29864);
or U30314 (N_30314,N_29677,N_29604);
or U30315 (N_30315,N_29936,N_29724);
nor U30316 (N_30316,N_29517,N_29751);
or U30317 (N_30317,N_29915,N_29685);
and U30318 (N_30318,N_29941,N_29622);
nand U30319 (N_30319,N_29906,N_29570);
nand U30320 (N_30320,N_29613,N_29524);
nor U30321 (N_30321,N_29770,N_29899);
and U30322 (N_30322,N_29554,N_29982);
and U30323 (N_30323,N_29800,N_29695);
nor U30324 (N_30324,N_29777,N_29876);
or U30325 (N_30325,N_29874,N_29782);
xor U30326 (N_30326,N_29506,N_29510);
or U30327 (N_30327,N_29843,N_29972);
and U30328 (N_30328,N_29875,N_29657);
nand U30329 (N_30329,N_29507,N_29919);
or U30330 (N_30330,N_29645,N_29587);
nand U30331 (N_30331,N_29803,N_29550);
nand U30332 (N_30332,N_29526,N_29754);
or U30333 (N_30333,N_29767,N_29569);
xor U30334 (N_30334,N_29705,N_29838);
nand U30335 (N_30335,N_29622,N_29951);
xor U30336 (N_30336,N_29909,N_29957);
and U30337 (N_30337,N_29853,N_29939);
xor U30338 (N_30338,N_29802,N_29644);
nor U30339 (N_30339,N_29655,N_29582);
nand U30340 (N_30340,N_29902,N_29784);
nor U30341 (N_30341,N_29947,N_29679);
xor U30342 (N_30342,N_29823,N_29773);
xor U30343 (N_30343,N_29793,N_29804);
or U30344 (N_30344,N_29684,N_29594);
xnor U30345 (N_30345,N_29576,N_29506);
and U30346 (N_30346,N_29851,N_29907);
nand U30347 (N_30347,N_29962,N_29500);
or U30348 (N_30348,N_29690,N_29604);
or U30349 (N_30349,N_29963,N_29553);
nor U30350 (N_30350,N_29755,N_29792);
and U30351 (N_30351,N_29610,N_29529);
nor U30352 (N_30352,N_29920,N_29790);
xnor U30353 (N_30353,N_29824,N_29809);
and U30354 (N_30354,N_29762,N_29728);
or U30355 (N_30355,N_29761,N_29752);
nor U30356 (N_30356,N_29610,N_29667);
or U30357 (N_30357,N_29919,N_29703);
and U30358 (N_30358,N_29827,N_29855);
xnor U30359 (N_30359,N_29516,N_29601);
nor U30360 (N_30360,N_29645,N_29583);
nand U30361 (N_30361,N_29975,N_29553);
and U30362 (N_30362,N_29749,N_29531);
nor U30363 (N_30363,N_29807,N_29521);
and U30364 (N_30364,N_29720,N_29577);
and U30365 (N_30365,N_29584,N_29896);
nand U30366 (N_30366,N_29701,N_29955);
xor U30367 (N_30367,N_29861,N_29686);
and U30368 (N_30368,N_29904,N_29810);
or U30369 (N_30369,N_29656,N_29951);
xnor U30370 (N_30370,N_29810,N_29949);
or U30371 (N_30371,N_29861,N_29510);
or U30372 (N_30372,N_29782,N_29690);
nand U30373 (N_30373,N_29667,N_29503);
nor U30374 (N_30374,N_29686,N_29602);
nor U30375 (N_30375,N_29573,N_29778);
nor U30376 (N_30376,N_29777,N_29836);
nor U30377 (N_30377,N_29786,N_29793);
and U30378 (N_30378,N_29506,N_29507);
or U30379 (N_30379,N_29691,N_29907);
xor U30380 (N_30380,N_29563,N_29877);
or U30381 (N_30381,N_29939,N_29766);
xnor U30382 (N_30382,N_29567,N_29671);
and U30383 (N_30383,N_29790,N_29815);
and U30384 (N_30384,N_29505,N_29806);
nor U30385 (N_30385,N_29864,N_29541);
or U30386 (N_30386,N_29894,N_29604);
nor U30387 (N_30387,N_29846,N_29799);
xnor U30388 (N_30388,N_29837,N_29522);
or U30389 (N_30389,N_29953,N_29811);
xnor U30390 (N_30390,N_29662,N_29638);
or U30391 (N_30391,N_29976,N_29828);
or U30392 (N_30392,N_29705,N_29970);
and U30393 (N_30393,N_29944,N_29789);
nand U30394 (N_30394,N_29615,N_29512);
nor U30395 (N_30395,N_29978,N_29857);
or U30396 (N_30396,N_29574,N_29596);
or U30397 (N_30397,N_29999,N_29730);
and U30398 (N_30398,N_29603,N_29637);
xnor U30399 (N_30399,N_29509,N_29908);
nor U30400 (N_30400,N_29970,N_29741);
nand U30401 (N_30401,N_29582,N_29760);
nand U30402 (N_30402,N_29640,N_29747);
xor U30403 (N_30403,N_29626,N_29727);
nor U30404 (N_30404,N_29653,N_29680);
or U30405 (N_30405,N_29966,N_29590);
nor U30406 (N_30406,N_29584,N_29801);
and U30407 (N_30407,N_29518,N_29612);
xnor U30408 (N_30408,N_29677,N_29519);
or U30409 (N_30409,N_29957,N_29959);
and U30410 (N_30410,N_29984,N_29758);
and U30411 (N_30411,N_29786,N_29735);
and U30412 (N_30412,N_29583,N_29535);
xor U30413 (N_30413,N_29565,N_29942);
xor U30414 (N_30414,N_29695,N_29545);
nor U30415 (N_30415,N_29983,N_29610);
or U30416 (N_30416,N_29868,N_29697);
and U30417 (N_30417,N_29734,N_29527);
xor U30418 (N_30418,N_29652,N_29658);
xor U30419 (N_30419,N_29706,N_29965);
and U30420 (N_30420,N_29513,N_29552);
and U30421 (N_30421,N_29944,N_29651);
nand U30422 (N_30422,N_29527,N_29622);
and U30423 (N_30423,N_29731,N_29802);
nor U30424 (N_30424,N_29885,N_29841);
or U30425 (N_30425,N_29634,N_29705);
nand U30426 (N_30426,N_29920,N_29876);
and U30427 (N_30427,N_29788,N_29533);
nand U30428 (N_30428,N_29977,N_29935);
or U30429 (N_30429,N_29815,N_29748);
nand U30430 (N_30430,N_29551,N_29972);
and U30431 (N_30431,N_29807,N_29563);
xnor U30432 (N_30432,N_29874,N_29912);
and U30433 (N_30433,N_29970,N_29800);
and U30434 (N_30434,N_29862,N_29733);
nand U30435 (N_30435,N_29594,N_29682);
nor U30436 (N_30436,N_29922,N_29830);
nand U30437 (N_30437,N_29687,N_29924);
xor U30438 (N_30438,N_29782,N_29611);
xnor U30439 (N_30439,N_29676,N_29628);
nand U30440 (N_30440,N_29789,N_29624);
and U30441 (N_30441,N_29686,N_29891);
xnor U30442 (N_30442,N_29806,N_29576);
xor U30443 (N_30443,N_29736,N_29549);
or U30444 (N_30444,N_29790,N_29781);
xnor U30445 (N_30445,N_29738,N_29515);
or U30446 (N_30446,N_29629,N_29965);
and U30447 (N_30447,N_29734,N_29925);
or U30448 (N_30448,N_29502,N_29530);
and U30449 (N_30449,N_29666,N_29545);
and U30450 (N_30450,N_29757,N_29925);
or U30451 (N_30451,N_29853,N_29552);
and U30452 (N_30452,N_29842,N_29859);
or U30453 (N_30453,N_29574,N_29881);
or U30454 (N_30454,N_29784,N_29950);
and U30455 (N_30455,N_29533,N_29933);
nand U30456 (N_30456,N_29588,N_29684);
or U30457 (N_30457,N_29560,N_29615);
nor U30458 (N_30458,N_29658,N_29951);
xor U30459 (N_30459,N_29714,N_29588);
nand U30460 (N_30460,N_29768,N_29599);
and U30461 (N_30461,N_29959,N_29944);
nor U30462 (N_30462,N_29871,N_29635);
nand U30463 (N_30463,N_29510,N_29758);
and U30464 (N_30464,N_29949,N_29785);
and U30465 (N_30465,N_29986,N_29635);
xor U30466 (N_30466,N_29648,N_29905);
nand U30467 (N_30467,N_29897,N_29525);
or U30468 (N_30468,N_29511,N_29961);
nor U30469 (N_30469,N_29648,N_29986);
nor U30470 (N_30470,N_29579,N_29825);
xnor U30471 (N_30471,N_29585,N_29853);
or U30472 (N_30472,N_29508,N_29513);
or U30473 (N_30473,N_29542,N_29886);
xnor U30474 (N_30474,N_29664,N_29624);
nand U30475 (N_30475,N_29835,N_29980);
nand U30476 (N_30476,N_29659,N_29957);
or U30477 (N_30477,N_29883,N_29700);
xnor U30478 (N_30478,N_29503,N_29579);
or U30479 (N_30479,N_29882,N_29888);
nor U30480 (N_30480,N_29994,N_29857);
and U30481 (N_30481,N_29947,N_29907);
and U30482 (N_30482,N_29873,N_29842);
xnor U30483 (N_30483,N_29601,N_29834);
xor U30484 (N_30484,N_29757,N_29929);
nor U30485 (N_30485,N_29804,N_29694);
or U30486 (N_30486,N_29922,N_29531);
xor U30487 (N_30487,N_29870,N_29911);
xor U30488 (N_30488,N_29614,N_29879);
nand U30489 (N_30489,N_29723,N_29627);
nand U30490 (N_30490,N_29521,N_29815);
and U30491 (N_30491,N_29530,N_29938);
xnor U30492 (N_30492,N_29871,N_29673);
and U30493 (N_30493,N_29547,N_29905);
and U30494 (N_30494,N_29963,N_29822);
nor U30495 (N_30495,N_29970,N_29644);
or U30496 (N_30496,N_29951,N_29698);
and U30497 (N_30497,N_29546,N_29592);
or U30498 (N_30498,N_29937,N_29777);
nand U30499 (N_30499,N_29630,N_29711);
nor U30500 (N_30500,N_30023,N_30125);
or U30501 (N_30501,N_30068,N_30117);
or U30502 (N_30502,N_30083,N_30206);
nor U30503 (N_30503,N_30097,N_30468);
xor U30504 (N_30504,N_30153,N_30178);
xnor U30505 (N_30505,N_30240,N_30357);
and U30506 (N_30506,N_30067,N_30127);
and U30507 (N_30507,N_30166,N_30218);
nor U30508 (N_30508,N_30364,N_30103);
nand U30509 (N_30509,N_30078,N_30350);
xor U30510 (N_30510,N_30219,N_30325);
or U30511 (N_30511,N_30099,N_30165);
and U30512 (N_30512,N_30048,N_30447);
xor U30513 (N_30513,N_30060,N_30381);
and U30514 (N_30514,N_30435,N_30116);
nor U30515 (N_30515,N_30294,N_30304);
nor U30516 (N_30516,N_30188,N_30184);
nand U30517 (N_30517,N_30226,N_30293);
xor U30518 (N_30518,N_30448,N_30192);
nor U30519 (N_30519,N_30222,N_30253);
nor U30520 (N_30520,N_30079,N_30285);
or U30521 (N_30521,N_30174,N_30400);
nand U30522 (N_30522,N_30171,N_30076);
and U30523 (N_30523,N_30202,N_30061);
and U30524 (N_30524,N_30105,N_30254);
nand U30525 (N_30525,N_30035,N_30498);
xor U30526 (N_30526,N_30248,N_30157);
nor U30527 (N_30527,N_30493,N_30322);
or U30528 (N_30528,N_30112,N_30172);
xor U30529 (N_30529,N_30471,N_30451);
or U30530 (N_30530,N_30241,N_30394);
and U30531 (N_30531,N_30045,N_30413);
xor U30532 (N_30532,N_30311,N_30225);
nand U30533 (N_30533,N_30091,N_30303);
xnor U30534 (N_30534,N_30147,N_30146);
or U30535 (N_30535,N_30429,N_30314);
nand U30536 (N_30536,N_30133,N_30000);
or U30537 (N_30537,N_30194,N_30280);
nand U30538 (N_30538,N_30109,N_30110);
or U30539 (N_30539,N_30211,N_30197);
nand U30540 (N_30540,N_30030,N_30047);
nor U30541 (N_30541,N_30255,N_30385);
and U30542 (N_30542,N_30088,N_30329);
xnor U30543 (N_30543,N_30302,N_30195);
xnor U30544 (N_30544,N_30463,N_30049);
nand U30545 (N_30545,N_30081,N_30472);
and U30546 (N_30546,N_30270,N_30115);
xor U30547 (N_30547,N_30134,N_30200);
nor U30548 (N_30548,N_30388,N_30331);
xor U30549 (N_30549,N_30425,N_30180);
or U30550 (N_30550,N_30234,N_30063);
nand U30551 (N_30551,N_30274,N_30292);
xnor U30552 (N_30552,N_30397,N_30213);
xnor U30553 (N_30553,N_30461,N_30247);
nor U30554 (N_30554,N_30312,N_30179);
nor U30555 (N_30555,N_30196,N_30299);
nand U30556 (N_30556,N_30443,N_30164);
nand U30557 (N_30557,N_30428,N_30422);
or U30558 (N_30558,N_30283,N_30220);
nand U30559 (N_30559,N_30243,N_30017);
and U30560 (N_30560,N_30469,N_30440);
nand U30561 (N_30561,N_30136,N_30279);
xnor U30562 (N_30562,N_30345,N_30052);
xor U30563 (N_30563,N_30137,N_30305);
xor U30564 (N_30564,N_30129,N_30170);
nand U30565 (N_30565,N_30453,N_30346);
nand U30566 (N_30566,N_30231,N_30260);
nor U30567 (N_30567,N_30177,N_30439);
nand U30568 (N_30568,N_30215,N_30198);
xor U30569 (N_30569,N_30221,N_30335);
or U30570 (N_30570,N_30431,N_30114);
and U30571 (N_30571,N_30239,N_30058);
or U30572 (N_30572,N_30277,N_30075);
xnor U30573 (N_30573,N_30475,N_30173);
nand U30574 (N_30574,N_30444,N_30118);
nand U30575 (N_30575,N_30155,N_30056);
nand U30576 (N_30576,N_30190,N_30022);
nor U30577 (N_30577,N_30094,N_30089);
xnor U30578 (N_30578,N_30119,N_30427);
and U30579 (N_30579,N_30009,N_30405);
nor U30580 (N_30580,N_30046,N_30347);
or U30581 (N_30581,N_30135,N_30418);
nand U30582 (N_30582,N_30499,N_30483);
nor U30583 (N_30583,N_30482,N_30455);
nand U30584 (N_30584,N_30430,N_30488);
xnor U30585 (N_30585,N_30167,N_30041);
xor U30586 (N_30586,N_30309,N_30408);
and U30587 (N_30587,N_30460,N_30417);
and U30588 (N_30588,N_30301,N_30066);
and U30589 (N_30589,N_30378,N_30182);
or U30590 (N_30590,N_30007,N_30396);
or U30591 (N_30591,N_30039,N_30323);
xor U30592 (N_30592,N_30474,N_30193);
xor U30593 (N_30593,N_30491,N_30233);
or U30594 (N_30594,N_30002,N_30020);
nand U30595 (N_30595,N_30450,N_30242);
xnor U30596 (N_30596,N_30128,N_30420);
or U30597 (N_30597,N_30281,N_30106);
nor U30598 (N_30598,N_30399,N_30296);
or U30599 (N_30599,N_30236,N_30126);
and U30600 (N_30600,N_30393,N_30466);
nand U30601 (N_30601,N_30087,N_30070);
and U30602 (N_30602,N_30496,N_30336);
nor U30603 (N_30603,N_30288,N_30175);
nand U30604 (N_30604,N_30203,N_30481);
and U30605 (N_30605,N_30262,N_30452);
nand U30606 (N_30606,N_30354,N_30057);
nor U30607 (N_30607,N_30343,N_30423);
and U30608 (N_30608,N_30064,N_30355);
and U30609 (N_30609,N_30290,N_30478);
nand U30610 (N_30610,N_30214,N_30001);
xor U30611 (N_30611,N_30289,N_30217);
and U30612 (N_30612,N_30228,N_30208);
or U30613 (N_30613,N_30404,N_30362);
or U30614 (N_30614,N_30424,N_30264);
nor U30615 (N_30615,N_30025,N_30433);
xor U30616 (N_30616,N_30123,N_30005);
nand U30617 (N_30617,N_30207,N_30216);
xnor U30618 (N_30618,N_30010,N_30286);
xor U30619 (N_30619,N_30391,N_30374);
or U30620 (N_30620,N_30145,N_30326);
and U30621 (N_30621,N_30080,N_30138);
nor U30622 (N_30622,N_30386,N_30011);
xor U30623 (N_30623,N_30340,N_30232);
or U30624 (N_30624,N_30419,N_30142);
or U30625 (N_30625,N_30490,N_30051);
nand U30626 (N_30626,N_30016,N_30053);
nand U30627 (N_30627,N_30449,N_30410);
nor U30628 (N_30628,N_30229,N_30363);
or U30629 (N_30629,N_30409,N_30436);
nor U30630 (N_30630,N_30244,N_30084);
and U30631 (N_30631,N_30278,N_30210);
nand U30632 (N_30632,N_30122,N_30392);
and U30633 (N_30633,N_30008,N_30238);
xor U30634 (N_30634,N_30367,N_30470);
and U30635 (N_30635,N_30096,N_30037);
xor U30636 (N_30636,N_30403,N_30162);
or U30637 (N_30637,N_30344,N_30199);
nand U30638 (N_30638,N_30159,N_30237);
xor U30639 (N_30639,N_30090,N_30402);
xnor U30640 (N_30640,N_30334,N_30100);
nor U30641 (N_30641,N_30212,N_30019);
or U30642 (N_30642,N_30446,N_30298);
or U30643 (N_30643,N_30065,N_30265);
or U30644 (N_30644,N_30026,N_30258);
and U30645 (N_30645,N_30489,N_30456);
nor U30646 (N_30646,N_30328,N_30181);
xor U30647 (N_30647,N_30072,N_30168);
or U30648 (N_30648,N_30102,N_30327);
nand U30649 (N_30649,N_30441,N_30291);
xor U30650 (N_30650,N_30121,N_30191);
xor U30651 (N_30651,N_30415,N_30406);
nor U30652 (N_30652,N_30003,N_30158);
nand U30653 (N_30653,N_30380,N_30261);
nor U30654 (N_30654,N_30006,N_30412);
nand U30655 (N_30655,N_30376,N_30401);
xnor U30656 (N_30656,N_30368,N_30031);
xnor U30657 (N_30657,N_30004,N_30313);
nand U30658 (N_30658,N_30223,N_30148);
or U30659 (N_30659,N_30377,N_30477);
and U30660 (N_30660,N_30205,N_30356);
and U30661 (N_30661,N_30484,N_30479);
nand U30662 (N_30662,N_30390,N_30111);
nor U30663 (N_30663,N_30445,N_30324);
or U30664 (N_30664,N_30032,N_30055);
or U30665 (N_30665,N_30485,N_30308);
nand U30666 (N_30666,N_30082,N_30276);
nor U30667 (N_30667,N_30021,N_30338);
and U30668 (N_30668,N_30272,N_30250);
and U30669 (N_30669,N_30271,N_30073);
or U30670 (N_30670,N_30341,N_30152);
nor U30671 (N_30671,N_30266,N_30014);
and U30672 (N_30672,N_30373,N_30269);
xor U30673 (N_30673,N_30342,N_30370);
nand U30674 (N_30674,N_30186,N_30071);
or U30675 (N_30675,N_30108,N_30131);
and U30676 (N_30676,N_30185,N_30092);
or U30677 (N_30677,N_30337,N_30124);
and U30678 (N_30678,N_30132,N_30379);
nor U30679 (N_30679,N_30365,N_30414);
xnor U30680 (N_30680,N_30263,N_30044);
nor U30681 (N_30681,N_30437,N_30140);
nand U30682 (N_30682,N_30306,N_30421);
xor U30683 (N_30683,N_30361,N_30224);
and U30684 (N_30684,N_30150,N_30204);
xnor U30685 (N_30685,N_30040,N_30351);
nor U30686 (N_30686,N_30467,N_30256);
nor U30687 (N_30687,N_30395,N_30487);
nand U30688 (N_30688,N_30387,N_30230);
and U30689 (N_30689,N_30473,N_30348);
or U30690 (N_30690,N_30149,N_30257);
or U30691 (N_30691,N_30369,N_30201);
nand U30692 (N_30692,N_30161,N_30321);
nand U30693 (N_30693,N_30320,N_30176);
nor U30694 (N_30694,N_30457,N_30015);
nand U30695 (N_30695,N_30013,N_30163);
and U30696 (N_30696,N_30101,N_30295);
nor U30697 (N_30697,N_30034,N_30120);
and U30698 (N_30698,N_30438,N_30315);
nand U30699 (N_30699,N_30077,N_30416);
xor U30700 (N_30700,N_30411,N_30426);
nor U30701 (N_30701,N_30383,N_30209);
xnor U30702 (N_30702,N_30036,N_30476);
nand U30703 (N_30703,N_30113,N_30442);
xnor U30704 (N_30704,N_30458,N_30360);
and U30705 (N_30705,N_30027,N_30495);
nand U30706 (N_30706,N_30375,N_30454);
and U30707 (N_30707,N_30038,N_30389);
nor U30708 (N_30708,N_30259,N_30282);
nand U30709 (N_30709,N_30330,N_30059);
xor U30710 (N_30710,N_30307,N_30024);
nor U30711 (N_30711,N_30434,N_30332);
nor U30712 (N_30712,N_30251,N_30085);
and U30713 (N_30713,N_30143,N_30384);
xnor U30714 (N_30714,N_30086,N_30486);
or U30715 (N_30715,N_30012,N_30156);
nand U30716 (N_30716,N_30069,N_30382);
nand U30717 (N_30717,N_30339,N_30359);
and U30718 (N_30718,N_30492,N_30141);
or U30719 (N_30719,N_30317,N_30300);
nand U30720 (N_30720,N_30107,N_30462);
nor U30721 (N_30721,N_30054,N_30316);
or U30722 (N_30722,N_30358,N_30227);
nor U30723 (N_30723,N_30353,N_30028);
or U30724 (N_30724,N_30183,N_30249);
xor U30725 (N_30725,N_30095,N_30189);
xnor U30726 (N_30726,N_30187,N_30480);
nor U30727 (N_30727,N_30284,N_30352);
nor U30728 (N_30728,N_30318,N_30297);
nand U30729 (N_30729,N_30151,N_30093);
xnor U30730 (N_30730,N_30130,N_30235);
or U30731 (N_30731,N_30372,N_30018);
xnor U30732 (N_30732,N_30074,N_30459);
nor U30733 (N_30733,N_30154,N_30287);
nand U30734 (N_30734,N_30245,N_30349);
xor U30735 (N_30735,N_30139,N_30465);
nor U30736 (N_30736,N_30371,N_30319);
nand U30737 (N_30737,N_30144,N_30333);
nor U30738 (N_30738,N_30407,N_30494);
and U30739 (N_30739,N_30042,N_30043);
xnor U30740 (N_30740,N_30497,N_30252);
or U30741 (N_30741,N_30029,N_30268);
and U30742 (N_30742,N_30098,N_30104);
nand U30743 (N_30743,N_30169,N_30033);
or U30744 (N_30744,N_30398,N_30050);
or U30745 (N_30745,N_30366,N_30062);
or U30746 (N_30746,N_30275,N_30160);
or U30747 (N_30747,N_30267,N_30246);
and U30748 (N_30748,N_30310,N_30464);
nand U30749 (N_30749,N_30273,N_30432);
nor U30750 (N_30750,N_30046,N_30018);
nand U30751 (N_30751,N_30376,N_30144);
nor U30752 (N_30752,N_30140,N_30419);
and U30753 (N_30753,N_30446,N_30092);
and U30754 (N_30754,N_30010,N_30004);
or U30755 (N_30755,N_30482,N_30068);
nand U30756 (N_30756,N_30049,N_30142);
and U30757 (N_30757,N_30431,N_30408);
and U30758 (N_30758,N_30229,N_30187);
nand U30759 (N_30759,N_30092,N_30479);
nor U30760 (N_30760,N_30495,N_30353);
nand U30761 (N_30761,N_30137,N_30220);
and U30762 (N_30762,N_30419,N_30315);
or U30763 (N_30763,N_30134,N_30477);
nor U30764 (N_30764,N_30409,N_30204);
nor U30765 (N_30765,N_30230,N_30340);
and U30766 (N_30766,N_30485,N_30362);
nand U30767 (N_30767,N_30440,N_30229);
or U30768 (N_30768,N_30462,N_30392);
nand U30769 (N_30769,N_30314,N_30294);
xor U30770 (N_30770,N_30360,N_30289);
xnor U30771 (N_30771,N_30315,N_30420);
or U30772 (N_30772,N_30276,N_30124);
or U30773 (N_30773,N_30080,N_30432);
or U30774 (N_30774,N_30375,N_30084);
or U30775 (N_30775,N_30170,N_30194);
xnor U30776 (N_30776,N_30239,N_30019);
and U30777 (N_30777,N_30143,N_30080);
nor U30778 (N_30778,N_30059,N_30466);
or U30779 (N_30779,N_30280,N_30424);
or U30780 (N_30780,N_30215,N_30498);
nor U30781 (N_30781,N_30197,N_30158);
nor U30782 (N_30782,N_30356,N_30392);
nor U30783 (N_30783,N_30180,N_30314);
nand U30784 (N_30784,N_30166,N_30145);
and U30785 (N_30785,N_30487,N_30126);
or U30786 (N_30786,N_30461,N_30480);
nand U30787 (N_30787,N_30134,N_30102);
nand U30788 (N_30788,N_30068,N_30426);
and U30789 (N_30789,N_30009,N_30234);
nor U30790 (N_30790,N_30219,N_30048);
nor U30791 (N_30791,N_30445,N_30433);
or U30792 (N_30792,N_30260,N_30365);
nor U30793 (N_30793,N_30196,N_30123);
or U30794 (N_30794,N_30061,N_30425);
and U30795 (N_30795,N_30414,N_30041);
or U30796 (N_30796,N_30111,N_30426);
xnor U30797 (N_30797,N_30116,N_30484);
nor U30798 (N_30798,N_30491,N_30420);
xnor U30799 (N_30799,N_30201,N_30489);
nand U30800 (N_30800,N_30094,N_30109);
xnor U30801 (N_30801,N_30267,N_30090);
and U30802 (N_30802,N_30027,N_30447);
nand U30803 (N_30803,N_30417,N_30412);
or U30804 (N_30804,N_30368,N_30170);
xor U30805 (N_30805,N_30415,N_30489);
or U30806 (N_30806,N_30118,N_30386);
nand U30807 (N_30807,N_30111,N_30424);
nor U30808 (N_30808,N_30080,N_30258);
nand U30809 (N_30809,N_30474,N_30168);
nand U30810 (N_30810,N_30077,N_30166);
nand U30811 (N_30811,N_30219,N_30370);
or U30812 (N_30812,N_30239,N_30105);
nor U30813 (N_30813,N_30032,N_30200);
xnor U30814 (N_30814,N_30074,N_30333);
nand U30815 (N_30815,N_30324,N_30102);
nor U30816 (N_30816,N_30064,N_30249);
nor U30817 (N_30817,N_30225,N_30272);
or U30818 (N_30818,N_30217,N_30365);
nor U30819 (N_30819,N_30120,N_30243);
or U30820 (N_30820,N_30044,N_30485);
or U30821 (N_30821,N_30038,N_30416);
nor U30822 (N_30822,N_30368,N_30356);
or U30823 (N_30823,N_30446,N_30269);
or U30824 (N_30824,N_30467,N_30289);
or U30825 (N_30825,N_30138,N_30415);
nand U30826 (N_30826,N_30418,N_30146);
and U30827 (N_30827,N_30190,N_30313);
and U30828 (N_30828,N_30143,N_30125);
xor U30829 (N_30829,N_30078,N_30198);
xnor U30830 (N_30830,N_30124,N_30449);
nor U30831 (N_30831,N_30352,N_30406);
nand U30832 (N_30832,N_30395,N_30303);
and U30833 (N_30833,N_30298,N_30474);
and U30834 (N_30834,N_30147,N_30070);
nor U30835 (N_30835,N_30415,N_30236);
nor U30836 (N_30836,N_30262,N_30332);
and U30837 (N_30837,N_30482,N_30400);
xnor U30838 (N_30838,N_30037,N_30372);
and U30839 (N_30839,N_30316,N_30223);
nand U30840 (N_30840,N_30177,N_30028);
or U30841 (N_30841,N_30376,N_30406);
and U30842 (N_30842,N_30404,N_30175);
and U30843 (N_30843,N_30390,N_30120);
nor U30844 (N_30844,N_30029,N_30312);
xor U30845 (N_30845,N_30386,N_30125);
or U30846 (N_30846,N_30299,N_30336);
and U30847 (N_30847,N_30100,N_30336);
or U30848 (N_30848,N_30218,N_30241);
nand U30849 (N_30849,N_30193,N_30147);
and U30850 (N_30850,N_30432,N_30279);
and U30851 (N_30851,N_30405,N_30096);
xnor U30852 (N_30852,N_30000,N_30450);
nand U30853 (N_30853,N_30339,N_30401);
xor U30854 (N_30854,N_30056,N_30141);
and U30855 (N_30855,N_30313,N_30371);
xnor U30856 (N_30856,N_30358,N_30131);
xor U30857 (N_30857,N_30123,N_30212);
or U30858 (N_30858,N_30104,N_30473);
or U30859 (N_30859,N_30250,N_30144);
xnor U30860 (N_30860,N_30275,N_30101);
or U30861 (N_30861,N_30028,N_30465);
or U30862 (N_30862,N_30147,N_30067);
nor U30863 (N_30863,N_30403,N_30077);
nor U30864 (N_30864,N_30268,N_30283);
and U30865 (N_30865,N_30059,N_30290);
or U30866 (N_30866,N_30137,N_30067);
or U30867 (N_30867,N_30224,N_30487);
nor U30868 (N_30868,N_30398,N_30058);
or U30869 (N_30869,N_30321,N_30001);
nor U30870 (N_30870,N_30097,N_30113);
or U30871 (N_30871,N_30056,N_30320);
or U30872 (N_30872,N_30058,N_30061);
and U30873 (N_30873,N_30296,N_30321);
nand U30874 (N_30874,N_30351,N_30098);
xor U30875 (N_30875,N_30420,N_30058);
or U30876 (N_30876,N_30160,N_30488);
nand U30877 (N_30877,N_30418,N_30181);
and U30878 (N_30878,N_30295,N_30141);
and U30879 (N_30879,N_30080,N_30074);
nor U30880 (N_30880,N_30087,N_30080);
or U30881 (N_30881,N_30432,N_30475);
nor U30882 (N_30882,N_30439,N_30069);
or U30883 (N_30883,N_30305,N_30412);
or U30884 (N_30884,N_30247,N_30391);
or U30885 (N_30885,N_30161,N_30287);
and U30886 (N_30886,N_30405,N_30396);
xnor U30887 (N_30887,N_30118,N_30060);
xnor U30888 (N_30888,N_30492,N_30476);
and U30889 (N_30889,N_30001,N_30016);
and U30890 (N_30890,N_30455,N_30033);
nand U30891 (N_30891,N_30381,N_30258);
nand U30892 (N_30892,N_30419,N_30234);
nand U30893 (N_30893,N_30046,N_30095);
or U30894 (N_30894,N_30273,N_30139);
xnor U30895 (N_30895,N_30064,N_30018);
and U30896 (N_30896,N_30061,N_30246);
or U30897 (N_30897,N_30342,N_30361);
and U30898 (N_30898,N_30125,N_30220);
nor U30899 (N_30899,N_30321,N_30049);
xnor U30900 (N_30900,N_30381,N_30292);
or U30901 (N_30901,N_30461,N_30146);
nand U30902 (N_30902,N_30071,N_30369);
and U30903 (N_30903,N_30376,N_30075);
and U30904 (N_30904,N_30392,N_30413);
nor U30905 (N_30905,N_30165,N_30460);
nor U30906 (N_30906,N_30274,N_30335);
or U30907 (N_30907,N_30080,N_30342);
and U30908 (N_30908,N_30165,N_30390);
nand U30909 (N_30909,N_30076,N_30005);
and U30910 (N_30910,N_30497,N_30016);
xnor U30911 (N_30911,N_30353,N_30151);
xor U30912 (N_30912,N_30134,N_30450);
nand U30913 (N_30913,N_30448,N_30402);
xor U30914 (N_30914,N_30182,N_30178);
or U30915 (N_30915,N_30252,N_30350);
and U30916 (N_30916,N_30011,N_30298);
xnor U30917 (N_30917,N_30283,N_30346);
nand U30918 (N_30918,N_30442,N_30235);
xor U30919 (N_30919,N_30374,N_30380);
nor U30920 (N_30920,N_30159,N_30429);
xor U30921 (N_30921,N_30341,N_30241);
or U30922 (N_30922,N_30482,N_30221);
and U30923 (N_30923,N_30203,N_30179);
or U30924 (N_30924,N_30350,N_30420);
or U30925 (N_30925,N_30333,N_30130);
and U30926 (N_30926,N_30465,N_30106);
nand U30927 (N_30927,N_30396,N_30044);
and U30928 (N_30928,N_30235,N_30369);
nand U30929 (N_30929,N_30164,N_30158);
xor U30930 (N_30930,N_30376,N_30425);
xor U30931 (N_30931,N_30350,N_30207);
and U30932 (N_30932,N_30044,N_30478);
and U30933 (N_30933,N_30000,N_30258);
nor U30934 (N_30934,N_30006,N_30335);
nor U30935 (N_30935,N_30214,N_30457);
xor U30936 (N_30936,N_30479,N_30290);
or U30937 (N_30937,N_30461,N_30285);
nand U30938 (N_30938,N_30378,N_30320);
xor U30939 (N_30939,N_30069,N_30118);
nand U30940 (N_30940,N_30128,N_30091);
or U30941 (N_30941,N_30068,N_30299);
or U30942 (N_30942,N_30032,N_30480);
nand U30943 (N_30943,N_30231,N_30272);
or U30944 (N_30944,N_30020,N_30313);
or U30945 (N_30945,N_30229,N_30278);
nor U30946 (N_30946,N_30489,N_30317);
and U30947 (N_30947,N_30037,N_30487);
xnor U30948 (N_30948,N_30081,N_30302);
nand U30949 (N_30949,N_30340,N_30219);
or U30950 (N_30950,N_30496,N_30053);
nor U30951 (N_30951,N_30372,N_30216);
or U30952 (N_30952,N_30479,N_30283);
nand U30953 (N_30953,N_30181,N_30260);
xor U30954 (N_30954,N_30436,N_30011);
nor U30955 (N_30955,N_30229,N_30315);
and U30956 (N_30956,N_30017,N_30132);
xnor U30957 (N_30957,N_30291,N_30089);
nand U30958 (N_30958,N_30169,N_30268);
nor U30959 (N_30959,N_30352,N_30264);
or U30960 (N_30960,N_30274,N_30394);
and U30961 (N_30961,N_30281,N_30374);
and U30962 (N_30962,N_30289,N_30059);
nor U30963 (N_30963,N_30172,N_30367);
or U30964 (N_30964,N_30359,N_30079);
nand U30965 (N_30965,N_30146,N_30426);
nand U30966 (N_30966,N_30184,N_30498);
nand U30967 (N_30967,N_30147,N_30448);
nor U30968 (N_30968,N_30050,N_30441);
or U30969 (N_30969,N_30455,N_30495);
nand U30970 (N_30970,N_30340,N_30387);
and U30971 (N_30971,N_30050,N_30285);
and U30972 (N_30972,N_30467,N_30051);
nor U30973 (N_30973,N_30295,N_30149);
xor U30974 (N_30974,N_30405,N_30414);
xnor U30975 (N_30975,N_30110,N_30117);
xor U30976 (N_30976,N_30383,N_30180);
or U30977 (N_30977,N_30026,N_30141);
nand U30978 (N_30978,N_30420,N_30408);
and U30979 (N_30979,N_30389,N_30069);
and U30980 (N_30980,N_30114,N_30029);
and U30981 (N_30981,N_30340,N_30339);
or U30982 (N_30982,N_30266,N_30013);
nand U30983 (N_30983,N_30089,N_30306);
nand U30984 (N_30984,N_30433,N_30230);
nor U30985 (N_30985,N_30039,N_30388);
xnor U30986 (N_30986,N_30319,N_30242);
or U30987 (N_30987,N_30025,N_30357);
xnor U30988 (N_30988,N_30025,N_30008);
nand U30989 (N_30989,N_30105,N_30307);
nor U30990 (N_30990,N_30046,N_30202);
xor U30991 (N_30991,N_30160,N_30087);
or U30992 (N_30992,N_30321,N_30261);
nand U30993 (N_30993,N_30033,N_30372);
nor U30994 (N_30994,N_30221,N_30077);
nand U30995 (N_30995,N_30010,N_30084);
and U30996 (N_30996,N_30274,N_30023);
nor U30997 (N_30997,N_30381,N_30281);
and U30998 (N_30998,N_30209,N_30115);
or U30999 (N_30999,N_30051,N_30182);
or U31000 (N_31000,N_30628,N_30600);
or U31001 (N_31001,N_30556,N_30551);
nor U31002 (N_31002,N_30879,N_30648);
nand U31003 (N_31003,N_30580,N_30785);
nor U31004 (N_31004,N_30905,N_30805);
xor U31005 (N_31005,N_30882,N_30668);
nor U31006 (N_31006,N_30962,N_30776);
or U31007 (N_31007,N_30566,N_30778);
nor U31008 (N_31008,N_30663,N_30715);
xor U31009 (N_31009,N_30756,N_30500);
or U31010 (N_31010,N_30986,N_30901);
and U31011 (N_31011,N_30814,N_30892);
nand U31012 (N_31012,N_30997,N_30545);
or U31013 (N_31013,N_30976,N_30810);
and U31014 (N_31014,N_30559,N_30771);
nor U31015 (N_31015,N_30590,N_30994);
or U31016 (N_31016,N_30624,N_30841);
nor U31017 (N_31017,N_30666,N_30627);
nand U31018 (N_31018,N_30846,N_30916);
nor U31019 (N_31019,N_30652,N_30938);
or U31020 (N_31020,N_30709,N_30923);
nand U31021 (N_31021,N_30594,N_30554);
nor U31022 (N_31022,N_30745,N_30830);
or U31023 (N_31023,N_30679,N_30815);
xor U31024 (N_31024,N_30525,N_30966);
or U31025 (N_31025,N_30783,N_30767);
and U31026 (N_31026,N_30929,N_30739);
or U31027 (N_31027,N_30670,N_30937);
nand U31028 (N_31028,N_30544,N_30788);
nor U31029 (N_31029,N_30769,N_30773);
nor U31030 (N_31030,N_30957,N_30607);
xnor U31031 (N_31031,N_30692,N_30862);
xnor U31032 (N_31032,N_30506,N_30516);
or U31033 (N_31033,N_30729,N_30738);
nor U31034 (N_31034,N_30806,N_30874);
nor U31035 (N_31035,N_30755,N_30602);
or U31036 (N_31036,N_30890,N_30943);
nand U31037 (N_31037,N_30936,N_30680);
xor U31038 (N_31038,N_30939,N_30548);
nand U31039 (N_31039,N_30909,N_30694);
nor U31040 (N_31040,N_30996,N_30904);
xnor U31041 (N_31041,N_30768,N_30780);
nand U31042 (N_31042,N_30542,N_30575);
nand U31043 (N_31043,N_30722,N_30796);
and U31044 (N_31044,N_30610,N_30884);
or U31045 (N_31045,N_30565,N_30880);
or U31046 (N_31046,N_30951,N_30711);
nand U31047 (N_31047,N_30681,N_30959);
and U31048 (N_31048,N_30707,N_30800);
nand U31049 (N_31049,N_30868,N_30691);
nor U31050 (N_31050,N_30592,N_30665);
xor U31051 (N_31051,N_30917,N_30688);
nand U31052 (N_31052,N_30974,N_30553);
and U31053 (N_31053,N_30913,N_30889);
nand U31054 (N_31054,N_30759,N_30945);
xnor U31055 (N_31055,N_30644,N_30664);
xnor U31056 (N_31056,N_30865,N_30730);
xor U31057 (N_31057,N_30657,N_30898);
xor U31058 (N_31058,N_30908,N_30712);
nor U31059 (N_31059,N_30561,N_30522);
nor U31060 (N_31060,N_30779,N_30503);
and U31061 (N_31061,N_30514,N_30507);
nand U31062 (N_31062,N_30878,N_30741);
and U31063 (N_31063,N_30870,N_30971);
nand U31064 (N_31064,N_30751,N_30579);
and U31065 (N_31065,N_30912,N_30930);
and U31066 (N_31066,N_30911,N_30601);
xnor U31067 (N_31067,N_30984,N_30724);
nor U31068 (N_31068,N_30761,N_30988);
or U31069 (N_31069,N_30574,N_30940);
and U31070 (N_31070,N_30825,N_30813);
xor U31071 (N_31071,N_30550,N_30696);
or U31072 (N_31072,N_30686,N_30701);
xnor U31073 (N_31073,N_30535,N_30989);
nand U31074 (N_31074,N_30802,N_30650);
nor U31075 (N_31075,N_30669,N_30833);
nor U31076 (N_31076,N_30826,N_30999);
nand U31077 (N_31077,N_30505,N_30546);
or U31078 (N_31078,N_30533,N_30791);
nor U31079 (N_31079,N_30706,N_30671);
xor U31080 (N_31080,N_30736,N_30599);
nor U31081 (N_31081,N_30964,N_30570);
xnor U31082 (N_31082,N_30513,N_30555);
and U31083 (N_31083,N_30534,N_30972);
nor U31084 (N_31084,N_30772,N_30797);
or U31085 (N_31085,N_30812,N_30893);
xnor U31086 (N_31086,N_30655,N_30817);
nand U31087 (N_31087,N_30743,N_30941);
nor U31088 (N_31088,N_30683,N_30987);
or U31089 (N_31089,N_30876,N_30928);
nand U31090 (N_31090,N_30511,N_30858);
or U31091 (N_31091,N_30867,N_30883);
nand U31092 (N_31092,N_30907,N_30922);
and U31093 (N_31093,N_30843,N_30848);
nor U31094 (N_31094,N_30558,N_30992);
nand U31095 (N_31095,N_30895,N_30524);
nand U31096 (N_31096,N_30869,N_30568);
nand U31097 (N_31097,N_30864,N_30571);
or U31098 (N_31098,N_30623,N_30527);
and U31099 (N_31099,N_30539,N_30781);
and U31100 (N_31100,N_30541,N_30614);
nand U31101 (N_31101,N_30836,N_30667);
nand U31102 (N_31102,N_30630,N_30721);
nor U31103 (N_31103,N_30762,N_30727);
xor U31104 (N_31104,N_30888,N_30676);
or U31105 (N_31105,N_30983,N_30713);
and U31106 (N_31106,N_30645,N_30801);
nor U31107 (N_31107,N_30637,N_30685);
xor U31108 (N_31108,N_30958,N_30920);
and U31109 (N_31109,N_30654,N_30563);
and U31110 (N_31110,N_30823,N_30749);
nand U31111 (N_31111,N_30529,N_30746);
xor U31112 (N_31112,N_30946,N_30793);
xor U31113 (N_31113,N_30723,N_30961);
nand U31114 (N_31114,N_30857,N_30789);
nand U31115 (N_31115,N_30734,N_30673);
nand U31116 (N_31116,N_30642,N_30786);
or U31117 (N_31117,N_30595,N_30611);
xor U31118 (N_31118,N_30641,N_30822);
nand U31119 (N_31119,N_30528,N_30621);
or U31120 (N_31120,N_30872,N_30699);
or U31121 (N_31121,N_30702,N_30687);
nor U31122 (N_31122,N_30803,N_30588);
nand U31123 (N_31123,N_30526,N_30969);
nor U31124 (N_31124,N_30714,N_30859);
xnor U31125 (N_31125,N_30921,N_30863);
nor U31126 (N_31126,N_30717,N_30847);
xnor U31127 (N_31127,N_30952,N_30799);
xor U31128 (N_31128,N_30716,N_30656);
or U31129 (N_31129,N_30586,N_30512);
xnor U31130 (N_31130,N_30998,N_30515);
nand U31131 (N_31131,N_30742,N_30728);
nand U31132 (N_31132,N_30585,N_30617);
nand U31133 (N_31133,N_30619,N_30616);
nor U31134 (N_31134,N_30960,N_30530);
or U31135 (N_31135,N_30861,N_30629);
or U31136 (N_31136,N_30816,N_30675);
nor U31137 (N_31137,N_30837,N_30705);
and U31138 (N_31138,N_30735,N_30918);
and U31139 (N_31139,N_30659,N_30851);
nand U31140 (N_31140,N_30804,N_30564);
xor U31141 (N_31141,N_30933,N_30919);
nand U31142 (N_31142,N_30835,N_30774);
nand U31143 (N_31143,N_30903,N_30626);
xnor U31144 (N_31144,N_30708,N_30661);
and U31145 (N_31145,N_30842,N_30832);
and U31146 (N_31146,N_30733,N_30924);
nand U31147 (N_31147,N_30737,N_30682);
nor U31148 (N_31148,N_30794,N_30598);
nor U31149 (N_31149,N_30583,N_30827);
and U31150 (N_31150,N_30854,N_30609);
nor U31151 (N_31151,N_30632,N_30975);
nor U31152 (N_31152,N_30828,N_30757);
nand U31153 (N_31153,N_30605,N_30981);
and U31154 (N_31154,N_30718,N_30856);
or U31155 (N_31155,N_30567,N_30613);
or U31156 (N_31156,N_30944,N_30660);
nand U31157 (N_31157,N_30636,N_30573);
or U31158 (N_31158,N_30792,N_30519);
and U31159 (N_31159,N_30932,N_30784);
xnor U31160 (N_31160,N_30523,N_30866);
or U31161 (N_31161,N_30543,N_30608);
and U31162 (N_31162,N_30770,N_30521);
and U31163 (N_31163,N_30798,N_30754);
or U31164 (N_31164,N_30578,N_30819);
nor U31165 (N_31165,N_30766,N_30552);
nand U31166 (N_31166,N_30584,N_30719);
or U31167 (N_31167,N_30537,N_30809);
nor U31168 (N_31168,N_30606,N_30993);
nor U31169 (N_31169,N_30820,N_30569);
nor U31170 (N_31170,N_30509,N_30562);
xor U31171 (N_31171,N_30821,N_30593);
nor U31172 (N_31172,N_30710,N_30634);
nor U31173 (N_31173,N_30982,N_30577);
xor U31174 (N_31174,N_30965,N_30517);
nand U31175 (N_31175,N_30560,N_30615);
nand U31176 (N_31176,N_30844,N_30850);
xor U31177 (N_31177,N_30647,N_30576);
xnor U31178 (N_31178,N_30808,N_30956);
xor U31179 (N_31179,N_30980,N_30591);
or U31180 (N_31180,N_30931,N_30536);
and U31181 (N_31181,N_30547,N_30698);
or U31182 (N_31182,N_30587,N_30906);
nor U31183 (N_31183,N_30549,N_30875);
xor U31184 (N_31184,N_30978,N_30845);
or U31185 (N_31185,N_30926,N_30902);
or U31186 (N_31186,N_30697,N_30557);
xnor U31187 (N_31187,N_30760,N_30990);
and U31188 (N_31188,N_30985,N_30855);
or U31189 (N_31189,N_30758,N_30894);
and U31190 (N_31190,N_30777,N_30695);
nor U31191 (N_31191,N_30834,N_30891);
xnor U31192 (N_31192,N_30763,N_30690);
or U31193 (N_31193,N_30635,N_30790);
and U31194 (N_31194,N_30955,N_30925);
nor U31195 (N_31195,N_30995,N_30953);
xor U31196 (N_31196,N_30658,N_30831);
and U31197 (N_31197,N_30887,N_30638);
or U31198 (N_31198,N_30967,N_30947);
nor U31199 (N_31199,N_30674,N_30662);
xor U31200 (N_31200,N_30732,N_30581);
nor U31201 (N_31201,N_30504,N_30753);
nand U31202 (N_31202,N_30508,N_30653);
nor U31203 (N_31203,N_30684,N_30752);
or U31204 (N_31204,N_30818,N_30750);
nand U31205 (N_31205,N_30704,N_30612);
nor U31206 (N_31206,N_30764,N_30622);
xor U31207 (N_31207,N_30775,N_30935);
or U31208 (N_31208,N_30731,N_30838);
or U31209 (N_31209,N_30620,N_30640);
and U31210 (N_31210,N_30703,N_30625);
and U31211 (N_31211,N_30871,N_30782);
nand U31212 (N_31212,N_30839,N_30633);
and U31213 (N_31213,N_30582,N_30852);
or U31214 (N_31214,N_30991,N_30678);
xnor U31215 (N_31215,N_30604,N_30968);
nor U31216 (N_31216,N_30896,N_30914);
xnor U31217 (N_31217,N_30795,N_30881);
nand U31218 (N_31218,N_30725,N_30651);
nor U31219 (N_31219,N_30860,N_30501);
and U31220 (N_31220,N_30572,N_30631);
or U31221 (N_31221,N_30538,N_30700);
and U31222 (N_31222,N_30720,N_30886);
and U31223 (N_31223,N_30693,N_30646);
xnor U31224 (N_31224,N_30531,N_30787);
and U31225 (N_31225,N_30502,N_30596);
and U31226 (N_31226,N_30649,N_30910);
nand U31227 (N_31227,N_30927,N_30589);
and U31228 (N_31228,N_30899,N_30520);
xor U31229 (N_31229,N_30900,N_30950);
and U31230 (N_31230,N_30689,N_30824);
xnor U31231 (N_31231,N_30744,N_30979);
nor U31232 (N_31232,N_30518,N_30540);
nand U31233 (N_31233,N_30807,N_30973);
nand U31234 (N_31234,N_30977,N_30948);
or U31235 (N_31235,N_30726,N_30672);
nand U31236 (N_31236,N_30963,N_30829);
or U31237 (N_31237,N_30934,N_30639);
xnor U31238 (N_31238,N_30949,N_30849);
or U31239 (N_31239,N_30677,N_30915);
nand U31240 (N_31240,N_30740,N_30877);
nor U31241 (N_31241,N_30954,N_30748);
or U31242 (N_31242,N_30532,N_30811);
nor U31243 (N_31243,N_30885,N_30970);
nor U31244 (N_31244,N_30853,N_30942);
or U31245 (N_31245,N_30603,N_30873);
nand U31246 (N_31246,N_30897,N_30840);
or U31247 (N_31247,N_30643,N_30618);
or U31248 (N_31248,N_30510,N_30597);
nand U31249 (N_31249,N_30765,N_30747);
and U31250 (N_31250,N_30591,N_30801);
and U31251 (N_31251,N_30913,N_30968);
nor U31252 (N_31252,N_30791,N_30874);
nand U31253 (N_31253,N_30929,N_30921);
xor U31254 (N_31254,N_30573,N_30796);
or U31255 (N_31255,N_30906,N_30697);
xor U31256 (N_31256,N_30759,N_30669);
and U31257 (N_31257,N_30551,N_30660);
or U31258 (N_31258,N_30737,N_30611);
nor U31259 (N_31259,N_30964,N_30832);
nand U31260 (N_31260,N_30847,N_30710);
nand U31261 (N_31261,N_30757,N_30524);
nor U31262 (N_31262,N_30752,N_30602);
and U31263 (N_31263,N_30770,N_30561);
xnor U31264 (N_31264,N_30983,N_30805);
nand U31265 (N_31265,N_30850,N_30919);
nor U31266 (N_31266,N_30819,N_30902);
and U31267 (N_31267,N_30679,N_30996);
and U31268 (N_31268,N_30807,N_30535);
or U31269 (N_31269,N_30713,N_30752);
nor U31270 (N_31270,N_30500,N_30711);
or U31271 (N_31271,N_30892,N_30761);
and U31272 (N_31272,N_30594,N_30915);
nor U31273 (N_31273,N_30988,N_30823);
xnor U31274 (N_31274,N_30659,N_30995);
xnor U31275 (N_31275,N_30645,N_30911);
and U31276 (N_31276,N_30759,N_30514);
nand U31277 (N_31277,N_30668,N_30862);
xor U31278 (N_31278,N_30881,N_30988);
and U31279 (N_31279,N_30718,N_30573);
nor U31280 (N_31280,N_30806,N_30897);
nor U31281 (N_31281,N_30933,N_30821);
nor U31282 (N_31282,N_30667,N_30877);
nor U31283 (N_31283,N_30992,N_30990);
or U31284 (N_31284,N_30780,N_30800);
nand U31285 (N_31285,N_30805,N_30574);
nand U31286 (N_31286,N_30605,N_30993);
and U31287 (N_31287,N_30943,N_30677);
or U31288 (N_31288,N_30928,N_30702);
nand U31289 (N_31289,N_30813,N_30665);
nor U31290 (N_31290,N_30880,N_30783);
and U31291 (N_31291,N_30521,N_30657);
or U31292 (N_31292,N_30773,N_30543);
xor U31293 (N_31293,N_30742,N_30769);
xor U31294 (N_31294,N_30547,N_30927);
xor U31295 (N_31295,N_30945,N_30733);
or U31296 (N_31296,N_30665,N_30979);
or U31297 (N_31297,N_30942,N_30567);
or U31298 (N_31298,N_30735,N_30705);
nand U31299 (N_31299,N_30545,N_30988);
and U31300 (N_31300,N_30738,N_30502);
xnor U31301 (N_31301,N_30863,N_30855);
xor U31302 (N_31302,N_30692,N_30778);
nand U31303 (N_31303,N_30853,N_30538);
and U31304 (N_31304,N_30552,N_30762);
xor U31305 (N_31305,N_30989,N_30802);
nor U31306 (N_31306,N_30818,N_30894);
or U31307 (N_31307,N_30855,N_30773);
nand U31308 (N_31308,N_30986,N_30930);
or U31309 (N_31309,N_30870,N_30705);
xor U31310 (N_31310,N_30529,N_30779);
or U31311 (N_31311,N_30545,N_30619);
and U31312 (N_31312,N_30994,N_30792);
and U31313 (N_31313,N_30521,N_30846);
nor U31314 (N_31314,N_30809,N_30913);
nor U31315 (N_31315,N_30510,N_30531);
xor U31316 (N_31316,N_30522,N_30785);
nor U31317 (N_31317,N_30844,N_30717);
nor U31318 (N_31318,N_30632,N_30939);
nand U31319 (N_31319,N_30820,N_30915);
and U31320 (N_31320,N_30547,N_30636);
nor U31321 (N_31321,N_30893,N_30947);
nand U31322 (N_31322,N_30983,N_30627);
nand U31323 (N_31323,N_30502,N_30560);
nor U31324 (N_31324,N_30510,N_30800);
nand U31325 (N_31325,N_30930,N_30734);
and U31326 (N_31326,N_30750,N_30888);
or U31327 (N_31327,N_30933,N_30793);
xor U31328 (N_31328,N_30767,N_30754);
nor U31329 (N_31329,N_30854,N_30818);
nor U31330 (N_31330,N_30648,N_30631);
xor U31331 (N_31331,N_30610,N_30835);
and U31332 (N_31332,N_30671,N_30534);
nand U31333 (N_31333,N_30803,N_30736);
xor U31334 (N_31334,N_30541,N_30821);
xnor U31335 (N_31335,N_30858,N_30769);
and U31336 (N_31336,N_30541,N_30514);
and U31337 (N_31337,N_30709,N_30618);
nor U31338 (N_31338,N_30970,N_30735);
nand U31339 (N_31339,N_30867,N_30550);
xor U31340 (N_31340,N_30807,N_30591);
xnor U31341 (N_31341,N_30972,N_30772);
or U31342 (N_31342,N_30983,N_30679);
xnor U31343 (N_31343,N_30972,N_30665);
nor U31344 (N_31344,N_30894,N_30727);
nand U31345 (N_31345,N_30766,N_30734);
or U31346 (N_31346,N_30917,N_30820);
nand U31347 (N_31347,N_30541,N_30693);
xor U31348 (N_31348,N_30987,N_30815);
and U31349 (N_31349,N_30854,N_30707);
or U31350 (N_31350,N_30640,N_30666);
nor U31351 (N_31351,N_30573,N_30974);
or U31352 (N_31352,N_30777,N_30865);
nor U31353 (N_31353,N_30814,N_30713);
nand U31354 (N_31354,N_30538,N_30719);
xnor U31355 (N_31355,N_30525,N_30802);
or U31356 (N_31356,N_30665,N_30732);
xnor U31357 (N_31357,N_30793,N_30944);
xor U31358 (N_31358,N_30836,N_30720);
or U31359 (N_31359,N_30501,N_30641);
nand U31360 (N_31360,N_30882,N_30741);
nor U31361 (N_31361,N_30704,N_30599);
or U31362 (N_31362,N_30913,N_30689);
nand U31363 (N_31363,N_30930,N_30757);
nand U31364 (N_31364,N_30707,N_30999);
nand U31365 (N_31365,N_30683,N_30992);
or U31366 (N_31366,N_30941,N_30880);
xor U31367 (N_31367,N_30928,N_30656);
or U31368 (N_31368,N_30571,N_30815);
nor U31369 (N_31369,N_30613,N_30535);
and U31370 (N_31370,N_30714,N_30945);
nor U31371 (N_31371,N_30509,N_30936);
and U31372 (N_31372,N_30948,N_30683);
nand U31373 (N_31373,N_30778,N_30791);
nor U31374 (N_31374,N_30874,N_30635);
or U31375 (N_31375,N_30641,N_30567);
or U31376 (N_31376,N_30520,N_30950);
xnor U31377 (N_31377,N_30976,N_30835);
nand U31378 (N_31378,N_30573,N_30579);
or U31379 (N_31379,N_30648,N_30526);
or U31380 (N_31380,N_30523,N_30779);
nand U31381 (N_31381,N_30842,N_30755);
xnor U31382 (N_31382,N_30685,N_30535);
xnor U31383 (N_31383,N_30590,N_30588);
or U31384 (N_31384,N_30715,N_30892);
and U31385 (N_31385,N_30986,N_30663);
or U31386 (N_31386,N_30928,N_30826);
nor U31387 (N_31387,N_30597,N_30927);
xor U31388 (N_31388,N_30833,N_30667);
or U31389 (N_31389,N_30786,N_30501);
nand U31390 (N_31390,N_30676,N_30668);
nor U31391 (N_31391,N_30702,N_30626);
xnor U31392 (N_31392,N_30838,N_30904);
and U31393 (N_31393,N_30855,N_30714);
nand U31394 (N_31394,N_30793,N_30923);
and U31395 (N_31395,N_30809,N_30968);
or U31396 (N_31396,N_30640,N_30868);
and U31397 (N_31397,N_30827,N_30999);
xnor U31398 (N_31398,N_30700,N_30620);
or U31399 (N_31399,N_30993,N_30553);
nor U31400 (N_31400,N_30987,N_30874);
nor U31401 (N_31401,N_30516,N_30648);
nand U31402 (N_31402,N_30940,N_30790);
nand U31403 (N_31403,N_30920,N_30548);
xnor U31404 (N_31404,N_30679,N_30966);
and U31405 (N_31405,N_30856,N_30514);
xnor U31406 (N_31406,N_30952,N_30607);
or U31407 (N_31407,N_30978,N_30926);
or U31408 (N_31408,N_30738,N_30706);
nand U31409 (N_31409,N_30964,N_30953);
xnor U31410 (N_31410,N_30627,N_30818);
or U31411 (N_31411,N_30676,N_30651);
and U31412 (N_31412,N_30870,N_30619);
xor U31413 (N_31413,N_30971,N_30543);
xnor U31414 (N_31414,N_30939,N_30734);
nand U31415 (N_31415,N_30772,N_30623);
nand U31416 (N_31416,N_30766,N_30570);
xor U31417 (N_31417,N_30632,N_30781);
xnor U31418 (N_31418,N_30940,N_30910);
and U31419 (N_31419,N_30717,N_30742);
or U31420 (N_31420,N_30512,N_30855);
and U31421 (N_31421,N_30983,N_30601);
xnor U31422 (N_31422,N_30609,N_30689);
and U31423 (N_31423,N_30721,N_30525);
nor U31424 (N_31424,N_30677,N_30592);
nand U31425 (N_31425,N_30652,N_30603);
nand U31426 (N_31426,N_30887,N_30729);
or U31427 (N_31427,N_30950,N_30553);
and U31428 (N_31428,N_30887,N_30648);
or U31429 (N_31429,N_30696,N_30923);
xnor U31430 (N_31430,N_30876,N_30701);
xor U31431 (N_31431,N_30628,N_30578);
or U31432 (N_31432,N_30962,N_30739);
or U31433 (N_31433,N_30603,N_30671);
xor U31434 (N_31434,N_30878,N_30581);
nor U31435 (N_31435,N_30980,N_30806);
nand U31436 (N_31436,N_30772,N_30825);
or U31437 (N_31437,N_30889,N_30650);
or U31438 (N_31438,N_30823,N_30998);
xor U31439 (N_31439,N_30705,N_30920);
xnor U31440 (N_31440,N_30512,N_30983);
nand U31441 (N_31441,N_30500,N_30912);
nand U31442 (N_31442,N_30988,N_30983);
and U31443 (N_31443,N_30864,N_30771);
xnor U31444 (N_31444,N_30918,N_30709);
and U31445 (N_31445,N_30678,N_30739);
nand U31446 (N_31446,N_30890,N_30629);
or U31447 (N_31447,N_30916,N_30646);
nand U31448 (N_31448,N_30766,N_30620);
nand U31449 (N_31449,N_30877,N_30580);
or U31450 (N_31450,N_30651,N_30646);
and U31451 (N_31451,N_30997,N_30827);
and U31452 (N_31452,N_30572,N_30597);
or U31453 (N_31453,N_30816,N_30687);
nand U31454 (N_31454,N_30858,N_30942);
or U31455 (N_31455,N_30543,N_30579);
nor U31456 (N_31456,N_30786,N_30871);
xnor U31457 (N_31457,N_30771,N_30579);
nand U31458 (N_31458,N_30853,N_30909);
or U31459 (N_31459,N_30932,N_30511);
nand U31460 (N_31460,N_30579,N_30502);
or U31461 (N_31461,N_30718,N_30655);
nand U31462 (N_31462,N_30611,N_30544);
xor U31463 (N_31463,N_30734,N_30701);
xnor U31464 (N_31464,N_30981,N_30635);
and U31465 (N_31465,N_30999,N_30858);
or U31466 (N_31466,N_30900,N_30658);
nand U31467 (N_31467,N_30914,N_30893);
nor U31468 (N_31468,N_30630,N_30962);
and U31469 (N_31469,N_30746,N_30904);
nor U31470 (N_31470,N_30915,N_30706);
xor U31471 (N_31471,N_30679,N_30610);
nor U31472 (N_31472,N_30892,N_30952);
nor U31473 (N_31473,N_30949,N_30696);
or U31474 (N_31474,N_30750,N_30788);
and U31475 (N_31475,N_30914,N_30655);
xor U31476 (N_31476,N_30764,N_30870);
or U31477 (N_31477,N_30945,N_30970);
or U31478 (N_31478,N_30643,N_30878);
nand U31479 (N_31479,N_30777,N_30857);
nand U31480 (N_31480,N_30804,N_30754);
nand U31481 (N_31481,N_30562,N_30877);
nand U31482 (N_31482,N_30924,N_30670);
nor U31483 (N_31483,N_30540,N_30994);
xnor U31484 (N_31484,N_30578,N_30642);
or U31485 (N_31485,N_30970,N_30772);
nor U31486 (N_31486,N_30829,N_30649);
xnor U31487 (N_31487,N_30746,N_30689);
nor U31488 (N_31488,N_30604,N_30877);
and U31489 (N_31489,N_30809,N_30707);
xnor U31490 (N_31490,N_30767,N_30852);
nand U31491 (N_31491,N_30626,N_30769);
or U31492 (N_31492,N_30511,N_30957);
nand U31493 (N_31493,N_30913,N_30733);
or U31494 (N_31494,N_30895,N_30542);
and U31495 (N_31495,N_30979,N_30981);
nor U31496 (N_31496,N_30655,N_30552);
nand U31497 (N_31497,N_30682,N_30621);
xnor U31498 (N_31498,N_30892,N_30711);
or U31499 (N_31499,N_30711,N_30803);
xnor U31500 (N_31500,N_31480,N_31058);
nor U31501 (N_31501,N_31191,N_31260);
xnor U31502 (N_31502,N_31493,N_31430);
nor U31503 (N_31503,N_31233,N_31181);
nor U31504 (N_31504,N_31395,N_31294);
nand U31505 (N_31505,N_31164,N_31461);
or U31506 (N_31506,N_31353,N_31485);
nand U31507 (N_31507,N_31162,N_31245);
nand U31508 (N_31508,N_31465,N_31224);
nor U31509 (N_31509,N_31458,N_31014);
and U31510 (N_31510,N_31472,N_31095);
nor U31511 (N_31511,N_31416,N_31086);
nand U31512 (N_31512,N_31109,N_31286);
xnor U31513 (N_31513,N_31230,N_31213);
xor U31514 (N_31514,N_31178,N_31379);
or U31515 (N_31515,N_31141,N_31117);
nor U31516 (N_31516,N_31295,N_31399);
nor U31517 (N_31517,N_31307,N_31049);
nand U31518 (N_31518,N_31115,N_31207);
xor U31519 (N_31519,N_31039,N_31153);
or U31520 (N_31520,N_31124,N_31488);
nand U31521 (N_31521,N_31255,N_31144);
and U31522 (N_31522,N_31275,N_31433);
nand U31523 (N_31523,N_31269,N_31103);
or U31524 (N_31524,N_31177,N_31114);
xor U31525 (N_31525,N_31238,N_31483);
nor U31526 (N_31526,N_31031,N_31234);
xnor U31527 (N_31527,N_31138,N_31427);
nor U31528 (N_31528,N_31360,N_31249);
or U31529 (N_31529,N_31247,N_31273);
and U31530 (N_31530,N_31096,N_31087);
or U31531 (N_31531,N_31385,N_31173);
xor U31532 (N_31532,N_31278,N_31215);
and U31533 (N_31533,N_31121,N_31392);
xor U31534 (N_31534,N_31393,N_31072);
or U31535 (N_31535,N_31217,N_31362);
xor U31536 (N_31536,N_31155,N_31189);
nand U31537 (N_31537,N_31460,N_31139);
and U31538 (N_31538,N_31040,N_31205);
and U31539 (N_31539,N_31146,N_31079);
nor U31540 (N_31540,N_31229,N_31400);
and U31541 (N_31541,N_31467,N_31462);
nor U31542 (N_31542,N_31471,N_31372);
or U31543 (N_31543,N_31339,N_31010);
nand U31544 (N_31544,N_31232,N_31099);
and U31545 (N_31545,N_31332,N_31323);
xor U31546 (N_31546,N_31132,N_31293);
and U31547 (N_31547,N_31347,N_31473);
nor U31548 (N_31548,N_31413,N_31403);
or U31549 (N_31549,N_31280,N_31066);
and U31550 (N_31550,N_31168,N_31478);
nor U31551 (N_31551,N_31365,N_31017);
or U31552 (N_31552,N_31051,N_31348);
nor U31553 (N_31553,N_31450,N_31180);
nor U31554 (N_31554,N_31303,N_31391);
xor U31555 (N_31555,N_31292,N_31226);
and U31556 (N_31556,N_31186,N_31408);
and U31557 (N_31557,N_31006,N_31190);
nor U31558 (N_31558,N_31128,N_31080);
and U31559 (N_31559,N_31404,N_31016);
nand U31560 (N_31560,N_31005,N_31440);
or U31561 (N_31561,N_31169,N_31375);
nand U31562 (N_31562,N_31282,N_31171);
or U31563 (N_31563,N_31491,N_31004);
and U31564 (N_31564,N_31327,N_31383);
or U31565 (N_31565,N_31338,N_31325);
or U31566 (N_31566,N_31075,N_31411);
nor U31567 (N_31567,N_31011,N_31459);
nor U31568 (N_31568,N_31270,N_31432);
and U31569 (N_31569,N_31499,N_31033);
xnor U31570 (N_31570,N_31208,N_31057);
or U31571 (N_31571,N_31291,N_31137);
nor U31572 (N_31572,N_31140,N_31078);
nand U31573 (N_31573,N_31118,N_31160);
nand U31574 (N_31574,N_31065,N_31028);
nor U31575 (N_31575,N_31149,N_31412);
nor U31576 (N_31576,N_31311,N_31134);
and U31577 (N_31577,N_31452,N_31477);
or U31578 (N_31578,N_31243,N_31000);
nor U31579 (N_31579,N_31251,N_31044);
nand U31580 (N_31580,N_31268,N_31464);
and U31581 (N_31581,N_31283,N_31239);
xor U31582 (N_31582,N_31344,N_31402);
xor U31583 (N_31583,N_31236,N_31253);
nor U31584 (N_31584,N_31469,N_31389);
or U31585 (N_31585,N_31201,N_31068);
xnor U31586 (N_31586,N_31007,N_31097);
nor U31587 (N_31587,N_31091,N_31279);
or U31588 (N_31588,N_31377,N_31192);
nor U31589 (N_31589,N_31143,N_31310);
nand U31590 (N_31590,N_31474,N_31210);
nand U31591 (N_31591,N_31159,N_31037);
or U31592 (N_31592,N_31107,N_31198);
xnor U31593 (N_31593,N_31257,N_31074);
nand U31594 (N_31594,N_31104,N_31271);
and U31595 (N_31595,N_31009,N_31034);
and U31596 (N_31596,N_31015,N_31116);
or U31597 (N_31597,N_31076,N_31349);
nor U31598 (N_31598,N_31094,N_31285);
or U31599 (N_31599,N_31359,N_31484);
nand U31600 (N_31600,N_31357,N_31240);
and U31601 (N_31601,N_31219,N_31301);
xnor U31602 (N_31602,N_31148,N_31428);
or U31603 (N_31603,N_31185,N_31417);
and U31604 (N_31604,N_31123,N_31276);
or U31605 (N_31605,N_31422,N_31498);
nand U31606 (N_31606,N_31023,N_31151);
nand U31607 (N_31607,N_31290,N_31130);
nor U31608 (N_31608,N_31437,N_31330);
xnor U31609 (N_31609,N_31366,N_31110);
nor U31610 (N_31610,N_31431,N_31056);
and U31611 (N_31611,N_31263,N_31084);
nor U31612 (N_31612,N_31126,N_31390);
nand U31613 (N_31613,N_31252,N_31166);
nand U31614 (N_31614,N_31421,N_31435);
or U31615 (N_31615,N_31183,N_31259);
nand U31616 (N_31616,N_31083,N_31370);
and U31617 (N_31617,N_31441,N_31463);
and U31618 (N_31618,N_31150,N_31337);
nor U31619 (N_31619,N_31174,N_31256);
xnor U31620 (N_31620,N_31203,N_31012);
and U31621 (N_31621,N_31420,N_31306);
xor U31622 (N_31622,N_31298,N_31053);
nand U31623 (N_31623,N_31482,N_31077);
xnor U31624 (N_31624,N_31088,N_31244);
nor U31625 (N_31625,N_31407,N_31108);
or U31626 (N_31626,N_31093,N_31345);
xnor U31627 (N_31627,N_31127,N_31313);
nor U31628 (N_31628,N_31324,N_31085);
or U31629 (N_31629,N_31106,N_31172);
and U31630 (N_31630,N_31020,N_31001);
and U31631 (N_31631,N_31494,N_31434);
xor U31632 (N_31632,N_31228,N_31456);
xor U31633 (N_31633,N_31328,N_31013);
and U31634 (N_31634,N_31003,N_31351);
nand U31635 (N_31635,N_31312,N_31305);
and U31636 (N_31636,N_31489,N_31200);
and U31637 (N_31637,N_31444,N_31387);
and U31638 (N_31638,N_31061,N_31059);
nor U31639 (N_31639,N_31047,N_31361);
or U31640 (N_31640,N_31487,N_31231);
or U31641 (N_31641,N_31455,N_31424);
and U31642 (N_31642,N_31350,N_31098);
and U31643 (N_31643,N_31025,N_31382);
and U31644 (N_31644,N_31364,N_31336);
nand U31645 (N_31645,N_31157,N_31036);
xor U31646 (N_31646,N_31297,N_31163);
xnor U31647 (N_31647,N_31142,N_31054);
and U31648 (N_31648,N_31202,N_31287);
nor U31649 (N_31649,N_31481,N_31048);
nand U31650 (N_31650,N_31029,N_31131);
nand U31651 (N_31651,N_31439,N_31043);
nor U31652 (N_31652,N_31060,N_31363);
and U31653 (N_31653,N_31340,N_31386);
or U31654 (N_31654,N_31342,N_31175);
and U31655 (N_31655,N_31496,N_31343);
or U31656 (N_31656,N_31414,N_31308);
and U31657 (N_31657,N_31035,N_31062);
or U31658 (N_31658,N_31225,N_31277);
and U31659 (N_31659,N_31199,N_31492);
or U31660 (N_31660,N_31222,N_31398);
nand U31661 (N_31661,N_31064,N_31274);
nor U31662 (N_31662,N_31321,N_31018);
nor U31663 (N_31663,N_31378,N_31329);
and U31664 (N_31664,N_31046,N_31089);
and U31665 (N_31665,N_31438,N_31454);
xnor U31666 (N_31666,N_31267,N_31194);
and U31667 (N_31667,N_31479,N_31211);
and U31668 (N_31668,N_31448,N_31447);
or U31669 (N_31669,N_31248,N_31165);
or U31670 (N_31670,N_31394,N_31376);
xnor U31671 (N_31671,N_31024,N_31355);
xnor U31672 (N_31672,N_31038,N_31170);
and U31673 (N_31673,N_31261,N_31490);
nor U31674 (N_31674,N_31314,N_31442);
and U31675 (N_31675,N_31196,N_31429);
or U31676 (N_31676,N_31242,N_31443);
nor U31677 (N_31677,N_31426,N_31184);
xnor U31678 (N_31678,N_31220,N_31019);
or U31679 (N_31679,N_31216,N_31371);
or U31680 (N_31680,N_31397,N_31021);
and U31681 (N_31681,N_31373,N_31266);
nand U31682 (N_31682,N_31309,N_31002);
and U31683 (N_31683,N_31187,N_31356);
nand U31684 (N_31684,N_31246,N_31026);
nand U31685 (N_31685,N_31179,N_31147);
xor U31686 (N_31686,N_31315,N_31119);
nor U31687 (N_31687,N_31304,N_31195);
and U31688 (N_31688,N_31367,N_31346);
or U31689 (N_31689,N_31453,N_31129);
xnor U31690 (N_31690,N_31334,N_31100);
nor U31691 (N_31691,N_31073,N_31032);
or U31692 (N_31692,N_31204,N_31272);
xor U31693 (N_31693,N_31113,N_31237);
and U31694 (N_31694,N_31125,N_31223);
nor U31695 (N_31695,N_31258,N_31135);
nor U31696 (N_31696,N_31296,N_31476);
nand U31697 (N_31697,N_31102,N_31410);
nor U31698 (N_31698,N_31045,N_31470);
xor U31699 (N_31699,N_31241,N_31111);
and U31700 (N_31700,N_31302,N_31193);
xnor U31701 (N_31701,N_31071,N_31120);
nand U31702 (N_31702,N_31235,N_31406);
nand U31703 (N_31703,N_31380,N_31030);
nor U31704 (N_31704,N_31022,N_31497);
xor U31705 (N_31705,N_31221,N_31449);
or U31706 (N_31706,N_31070,N_31369);
and U31707 (N_31707,N_31212,N_31318);
nor U31708 (N_31708,N_31466,N_31188);
nand U31709 (N_31709,N_31090,N_31358);
and U31710 (N_31710,N_31468,N_31331);
or U31711 (N_31711,N_31105,N_31167);
nand U31712 (N_31712,N_31317,N_31486);
nand U31713 (N_31713,N_31161,N_31320);
xnor U31714 (N_31714,N_31409,N_31457);
or U31715 (N_31715,N_31122,N_31446);
or U31716 (N_31716,N_31423,N_31319);
xnor U31717 (N_31717,N_31069,N_31041);
nor U31718 (N_31718,N_31316,N_31008);
nor U31719 (N_31719,N_31436,N_31055);
nor U31720 (N_31720,N_31067,N_31354);
or U31721 (N_31721,N_31281,N_31152);
and U31722 (N_31722,N_31227,N_31322);
nand U31723 (N_31723,N_31415,N_31451);
or U31724 (N_31724,N_31063,N_31419);
nor U31725 (N_31725,N_31101,N_31042);
or U31726 (N_31726,N_31154,N_31250);
nor U31727 (N_31727,N_31381,N_31475);
nor U31728 (N_31728,N_31418,N_31352);
or U31729 (N_31729,N_31209,N_31288);
nor U31730 (N_31730,N_31197,N_31027);
or U31731 (N_31731,N_31326,N_31092);
nor U31732 (N_31732,N_31052,N_31374);
and U31733 (N_31733,N_31206,N_31289);
nand U31734 (N_31734,N_31341,N_31082);
nand U31735 (N_31735,N_31050,N_31145);
and U31736 (N_31736,N_31405,N_31265);
and U31737 (N_31737,N_31218,N_31158);
nor U31738 (N_31738,N_31262,N_31495);
or U31739 (N_31739,N_31214,N_31299);
nand U31740 (N_31740,N_31136,N_31182);
xor U31741 (N_31741,N_31133,N_31300);
or U31742 (N_31742,N_31112,N_31368);
and U31743 (N_31743,N_31264,N_31425);
nor U31744 (N_31744,N_31445,N_31156);
nor U31745 (N_31745,N_31333,N_31401);
or U31746 (N_31746,N_31388,N_31254);
or U31747 (N_31747,N_31081,N_31284);
or U31748 (N_31748,N_31396,N_31335);
or U31749 (N_31749,N_31176,N_31384);
and U31750 (N_31750,N_31060,N_31087);
xnor U31751 (N_31751,N_31460,N_31432);
nand U31752 (N_31752,N_31019,N_31178);
nand U31753 (N_31753,N_31033,N_31416);
xnor U31754 (N_31754,N_31047,N_31236);
xnor U31755 (N_31755,N_31088,N_31102);
xnor U31756 (N_31756,N_31094,N_31284);
and U31757 (N_31757,N_31286,N_31029);
or U31758 (N_31758,N_31334,N_31144);
nand U31759 (N_31759,N_31156,N_31198);
nor U31760 (N_31760,N_31429,N_31395);
nor U31761 (N_31761,N_31080,N_31065);
and U31762 (N_31762,N_31450,N_31407);
nor U31763 (N_31763,N_31312,N_31075);
nand U31764 (N_31764,N_31444,N_31414);
nor U31765 (N_31765,N_31008,N_31489);
and U31766 (N_31766,N_31357,N_31044);
nand U31767 (N_31767,N_31482,N_31221);
nor U31768 (N_31768,N_31214,N_31275);
nor U31769 (N_31769,N_31040,N_31020);
and U31770 (N_31770,N_31159,N_31225);
nand U31771 (N_31771,N_31498,N_31463);
nand U31772 (N_31772,N_31460,N_31467);
and U31773 (N_31773,N_31092,N_31097);
nor U31774 (N_31774,N_31466,N_31016);
and U31775 (N_31775,N_31493,N_31371);
xor U31776 (N_31776,N_31006,N_31147);
nor U31777 (N_31777,N_31459,N_31074);
nor U31778 (N_31778,N_31245,N_31187);
and U31779 (N_31779,N_31019,N_31363);
nor U31780 (N_31780,N_31058,N_31355);
and U31781 (N_31781,N_31436,N_31227);
xor U31782 (N_31782,N_31173,N_31183);
or U31783 (N_31783,N_31321,N_31403);
nor U31784 (N_31784,N_31005,N_31460);
nand U31785 (N_31785,N_31473,N_31239);
or U31786 (N_31786,N_31241,N_31402);
and U31787 (N_31787,N_31421,N_31164);
xor U31788 (N_31788,N_31278,N_31490);
xor U31789 (N_31789,N_31379,N_31190);
and U31790 (N_31790,N_31307,N_31069);
and U31791 (N_31791,N_31368,N_31306);
xnor U31792 (N_31792,N_31367,N_31022);
nor U31793 (N_31793,N_31427,N_31401);
or U31794 (N_31794,N_31330,N_31109);
xor U31795 (N_31795,N_31120,N_31048);
nand U31796 (N_31796,N_31073,N_31115);
and U31797 (N_31797,N_31146,N_31400);
and U31798 (N_31798,N_31445,N_31462);
nor U31799 (N_31799,N_31471,N_31481);
and U31800 (N_31800,N_31197,N_31412);
nand U31801 (N_31801,N_31040,N_31027);
or U31802 (N_31802,N_31493,N_31359);
nor U31803 (N_31803,N_31013,N_31218);
or U31804 (N_31804,N_31161,N_31471);
xor U31805 (N_31805,N_31439,N_31166);
nor U31806 (N_31806,N_31075,N_31326);
xor U31807 (N_31807,N_31052,N_31010);
xnor U31808 (N_31808,N_31201,N_31258);
and U31809 (N_31809,N_31357,N_31253);
or U31810 (N_31810,N_31072,N_31244);
and U31811 (N_31811,N_31261,N_31177);
or U31812 (N_31812,N_31096,N_31021);
or U31813 (N_31813,N_31358,N_31236);
and U31814 (N_31814,N_31046,N_31083);
nand U31815 (N_31815,N_31162,N_31216);
nor U31816 (N_31816,N_31473,N_31371);
or U31817 (N_31817,N_31234,N_31003);
nand U31818 (N_31818,N_31293,N_31214);
nor U31819 (N_31819,N_31122,N_31296);
and U31820 (N_31820,N_31416,N_31379);
nor U31821 (N_31821,N_31252,N_31398);
or U31822 (N_31822,N_31465,N_31421);
nor U31823 (N_31823,N_31494,N_31478);
xor U31824 (N_31824,N_31275,N_31223);
xor U31825 (N_31825,N_31433,N_31470);
nand U31826 (N_31826,N_31461,N_31150);
nor U31827 (N_31827,N_31353,N_31243);
nand U31828 (N_31828,N_31058,N_31126);
or U31829 (N_31829,N_31493,N_31361);
and U31830 (N_31830,N_31481,N_31391);
nand U31831 (N_31831,N_31456,N_31250);
or U31832 (N_31832,N_31033,N_31372);
and U31833 (N_31833,N_31347,N_31297);
nand U31834 (N_31834,N_31447,N_31397);
and U31835 (N_31835,N_31191,N_31019);
nand U31836 (N_31836,N_31413,N_31276);
nand U31837 (N_31837,N_31253,N_31058);
nand U31838 (N_31838,N_31468,N_31162);
xor U31839 (N_31839,N_31115,N_31466);
or U31840 (N_31840,N_31171,N_31188);
xnor U31841 (N_31841,N_31351,N_31171);
or U31842 (N_31842,N_31029,N_31031);
or U31843 (N_31843,N_31329,N_31115);
or U31844 (N_31844,N_31493,N_31467);
xor U31845 (N_31845,N_31023,N_31428);
nor U31846 (N_31846,N_31446,N_31220);
nor U31847 (N_31847,N_31327,N_31421);
and U31848 (N_31848,N_31233,N_31339);
nor U31849 (N_31849,N_31009,N_31012);
and U31850 (N_31850,N_31192,N_31103);
or U31851 (N_31851,N_31232,N_31046);
nor U31852 (N_31852,N_31351,N_31022);
and U31853 (N_31853,N_31273,N_31067);
and U31854 (N_31854,N_31379,N_31010);
xor U31855 (N_31855,N_31248,N_31250);
nor U31856 (N_31856,N_31393,N_31222);
nand U31857 (N_31857,N_31050,N_31242);
xor U31858 (N_31858,N_31370,N_31146);
xnor U31859 (N_31859,N_31014,N_31020);
nor U31860 (N_31860,N_31399,N_31131);
and U31861 (N_31861,N_31234,N_31257);
or U31862 (N_31862,N_31264,N_31113);
and U31863 (N_31863,N_31423,N_31175);
and U31864 (N_31864,N_31186,N_31007);
xnor U31865 (N_31865,N_31491,N_31411);
xnor U31866 (N_31866,N_31234,N_31055);
nand U31867 (N_31867,N_31123,N_31033);
nor U31868 (N_31868,N_31071,N_31475);
nand U31869 (N_31869,N_31344,N_31132);
or U31870 (N_31870,N_31303,N_31264);
nand U31871 (N_31871,N_31202,N_31264);
or U31872 (N_31872,N_31090,N_31022);
xor U31873 (N_31873,N_31243,N_31229);
xor U31874 (N_31874,N_31091,N_31264);
and U31875 (N_31875,N_31177,N_31069);
xor U31876 (N_31876,N_31035,N_31461);
nand U31877 (N_31877,N_31212,N_31203);
or U31878 (N_31878,N_31354,N_31181);
or U31879 (N_31879,N_31315,N_31006);
or U31880 (N_31880,N_31344,N_31115);
xnor U31881 (N_31881,N_31306,N_31013);
nand U31882 (N_31882,N_31133,N_31196);
xnor U31883 (N_31883,N_31436,N_31382);
nand U31884 (N_31884,N_31201,N_31317);
nor U31885 (N_31885,N_31274,N_31013);
nand U31886 (N_31886,N_31184,N_31247);
xnor U31887 (N_31887,N_31404,N_31174);
xnor U31888 (N_31888,N_31490,N_31418);
nor U31889 (N_31889,N_31178,N_31328);
xor U31890 (N_31890,N_31237,N_31187);
nand U31891 (N_31891,N_31423,N_31072);
xnor U31892 (N_31892,N_31153,N_31064);
nor U31893 (N_31893,N_31224,N_31070);
nor U31894 (N_31894,N_31417,N_31262);
nand U31895 (N_31895,N_31184,N_31491);
nor U31896 (N_31896,N_31452,N_31000);
xor U31897 (N_31897,N_31237,N_31233);
or U31898 (N_31898,N_31156,N_31082);
and U31899 (N_31899,N_31051,N_31430);
nor U31900 (N_31900,N_31161,N_31391);
and U31901 (N_31901,N_31121,N_31099);
or U31902 (N_31902,N_31058,N_31418);
or U31903 (N_31903,N_31182,N_31098);
and U31904 (N_31904,N_31411,N_31138);
xnor U31905 (N_31905,N_31217,N_31131);
and U31906 (N_31906,N_31276,N_31460);
nor U31907 (N_31907,N_31004,N_31440);
and U31908 (N_31908,N_31067,N_31398);
and U31909 (N_31909,N_31322,N_31435);
or U31910 (N_31910,N_31027,N_31112);
xnor U31911 (N_31911,N_31294,N_31224);
and U31912 (N_31912,N_31327,N_31402);
nand U31913 (N_31913,N_31443,N_31379);
and U31914 (N_31914,N_31293,N_31166);
nand U31915 (N_31915,N_31411,N_31139);
nand U31916 (N_31916,N_31013,N_31363);
xnor U31917 (N_31917,N_31025,N_31029);
or U31918 (N_31918,N_31177,N_31051);
or U31919 (N_31919,N_31107,N_31469);
xnor U31920 (N_31920,N_31471,N_31276);
nand U31921 (N_31921,N_31431,N_31024);
or U31922 (N_31922,N_31079,N_31262);
nor U31923 (N_31923,N_31227,N_31361);
nor U31924 (N_31924,N_31132,N_31098);
nor U31925 (N_31925,N_31290,N_31242);
or U31926 (N_31926,N_31250,N_31236);
xnor U31927 (N_31927,N_31257,N_31430);
xnor U31928 (N_31928,N_31224,N_31201);
or U31929 (N_31929,N_31232,N_31005);
nor U31930 (N_31930,N_31402,N_31178);
nor U31931 (N_31931,N_31009,N_31202);
or U31932 (N_31932,N_31327,N_31429);
nand U31933 (N_31933,N_31275,N_31132);
and U31934 (N_31934,N_31262,N_31240);
xnor U31935 (N_31935,N_31428,N_31287);
nand U31936 (N_31936,N_31369,N_31300);
and U31937 (N_31937,N_31049,N_31209);
nor U31938 (N_31938,N_31372,N_31307);
nand U31939 (N_31939,N_31262,N_31473);
nand U31940 (N_31940,N_31089,N_31274);
or U31941 (N_31941,N_31466,N_31105);
or U31942 (N_31942,N_31492,N_31170);
or U31943 (N_31943,N_31012,N_31253);
xor U31944 (N_31944,N_31273,N_31071);
nand U31945 (N_31945,N_31018,N_31056);
xnor U31946 (N_31946,N_31399,N_31380);
or U31947 (N_31947,N_31282,N_31013);
and U31948 (N_31948,N_31132,N_31246);
nor U31949 (N_31949,N_31170,N_31476);
nand U31950 (N_31950,N_31035,N_31047);
nor U31951 (N_31951,N_31019,N_31478);
or U31952 (N_31952,N_31233,N_31156);
and U31953 (N_31953,N_31487,N_31084);
and U31954 (N_31954,N_31446,N_31417);
and U31955 (N_31955,N_31099,N_31220);
nor U31956 (N_31956,N_31313,N_31117);
nor U31957 (N_31957,N_31053,N_31497);
xnor U31958 (N_31958,N_31413,N_31400);
nor U31959 (N_31959,N_31426,N_31450);
and U31960 (N_31960,N_31357,N_31047);
nor U31961 (N_31961,N_31442,N_31311);
nor U31962 (N_31962,N_31006,N_31136);
xnor U31963 (N_31963,N_31373,N_31120);
nand U31964 (N_31964,N_31400,N_31154);
and U31965 (N_31965,N_31056,N_31251);
nand U31966 (N_31966,N_31053,N_31010);
and U31967 (N_31967,N_31292,N_31033);
or U31968 (N_31968,N_31232,N_31089);
nor U31969 (N_31969,N_31291,N_31300);
nand U31970 (N_31970,N_31438,N_31353);
nor U31971 (N_31971,N_31437,N_31022);
or U31972 (N_31972,N_31114,N_31100);
nor U31973 (N_31973,N_31460,N_31080);
nor U31974 (N_31974,N_31030,N_31131);
xor U31975 (N_31975,N_31176,N_31286);
nor U31976 (N_31976,N_31471,N_31178);
nor U31977 (N_31977,N_31227,N_31077);
nor U31978 (N_31978,N_31313,N_31434);
nor U31979 (N_31979,N_31355,N_31310);
nor U31980 (N_31980,N_31082,N_31001);
xnor U31981 (N_31981,N_31220,N_31486);
xor U31982 (N_31982,N_31039,N_31313);
or U31983 (N_31983,N_31284,N_31372);
and U31984 (N_31984,N_31058,N_31375);
or U31985 (N_31985,N_31322,N_31448);
and U31986 (N_31986,N_31399,N_31497);
nor U31987 (N_31987,N_31229,N_31483);
and U31988 (N_31988,N_31142,N_31177);
xnor U31989 (N_31989,N_31071,N_31208);
nor U31990 (N_31990,N_31258,N_31162);
or U31991 (N_31991,N_31276,N_31476);
or U31992 (N_31992,N_31117,N_31453);
nor U31993 (N_31993,N_31231,N_31175);
nand U31994 (N_31994,N_31118,N_31192);
or U31995 (N_31995,N_31103,N_31335);
nand U31996 (N_31996,N_31304,N_31051);
or U31997 (N_31997,N_31245,N_31138);
and U31998 (N_31998,N_31420,N_31427);
xor U31999 (N_31999,N_31198,N_31135);
nand U32000 (N_32000,N_31697,N_31515);
nor U32001 (N_32001,N_31555,N_31758);
and U32002 (N_32002,N_31565,N_31873);
and U32003 (N_32003,N_31943,N_31830);
nor U32004 (N_32004,N_31818,N_31954);
and U32005 (N_32005,N_31920,N_31845);
or U32006 (N_32006,N_31586,N_31611);
and U32007 (N_32007,N_31699,N_31667);
xnor U32008 (N_32008,N_31532,N_31607);
xor U32009 (N_32009,N_31751,N_31548);
xnor U32010 (N_32010,N_31910,N_31942);
xor U32011 (N_32011,N_31575,N_31652);
or U32012 (N_32012,N_31654,N_31746);
and U32013 (N_32013,N_31808,N_31890);
and U32014 (N_32014,N_31940,N_31701);
nor U32015 (N_32015,N_31550,N_31922);
xor U32016 (N_32016,N_31571,N_31535);
nand U32017 (N_32017,N_31825,N_31719);
nand U32018 (N_32018,N_31559,N_31868);
and U32019 (N_32019,N_31681,N_31802);
nand U32020 (N_32020,N_31506,N_31865);
xnor U32021 (N_32021,N_31888,N_31930);
and U32022 (N_32022,N_31627,N_31525);
nor U32023 (N_32023,N_31648,N_31842);
nor U32024 (N_32024,N_31529,N_31848);
xor U32025 (N_32025,N_31821,N_31969);
xor U32026 (N_32026,N_31740,N_31572);
or U32027 (N_32027,N_31588,N_31988);
and U32028 (N_32028,N_31909,N_31584);
and U32029 (N_32029,N_31776,N_31749);
xnor U32030 (N_32030,N_31946,N_31540);
and U32031 (N_32031,N_31747,N_31990);
or U32032 (N_32032,N_31750,N_31502);
nand U32033 (N_32033,N_31963,N_31925);
xnor U32034 (N_32034,N_31763,N_31570);
or U32035 (N_32035,N_31849,N_31884);
nor U32036 (N_32036,N_31709,N_31861);
nand U32037 (N_32037,N_31833,N_31629);
xnor U32038 (N_32038,N_31949,N_31508);
and U32039 (N_32039,N_31926,N_31517);
and U32040 (N_32040,N_31896,N_31616);
and U32041 (N_32041,N_31640,N_31784);
or U32042 (N_32042,N_31753,N_31827);
or U32043 (N_32043,N_31676,N_31564);
and U32044 (N_32044,N_31916,N_31580);
and U32045 (N_32045,N_31579,N_31773);
nor U32046 (N_32046,N_31610,N_31788);
nand U32047 (N_32047,N_31834,N_31992);
nor U32048 (N_32048,N_31671,N_31974);
nor U32049 (N_32049,N_31786,N_31824);
nor U32050 (N_32050,N_31767,N_31505);
and U32051 (N_32051,N_31708,N_31642);
nor U32052 (N_32052,N_31625,N_31686);
nor U32053 (N_32053,N_31677,N_31805);
nor U32054 (N_32054,N_31967,N_31662);
nand U32055 (N_32055,N_31964,N_31975);
or U32056 (N_32056,N_31594,N_31847);
nand U32057 (N_32057,N_31822,N_31986);
and U32058 (N_32058,N_31760,N_31700);
or U32059 (N_32059,N_31601,N_31702);
xnor U32060 (N_32060,N_31578,N_31661);
and U32061 (N_32061,N_31800,N_31630);
and U32062 (N_32062,N_31898,N_31593);
or U32063 (N_32063,N_31595,N_31703);
and U32064 (N_32064,N_31936,N_31774);
or U32065 (N_32065,N_31731,N_31645);
and U32066 (N_32066,N_31779,N_31887);
nor U32067 (N_32067,N_31889,N_31951);
and U32068 (N_32068,N_31966,N_31993);
nand U32069 (N_32069,N_31798,N_31526);
nand U32070 (N_32070,N_31793,N_31810);
and U32071 (N_32071,N_31639,N_31693);
xor U32072 (N_32072,N_31513,N_31866);
xnor U32073 (N_32073,N_31799,N_31835);
or U32074 (N_32074,N_31716,N_31987);
or U32075 (N_32075,N_31807,N_31885);
or U32076 (N_32076,N_31907,N_31553);
or U32077 (N_32077,N_31787,N_31634);
nand U32078 (N_32078,N_31649,N_31734);
xnor U32079 (N_32079,N_31689,N_31694);
xor U32080 (N_32080,N_31696,N_31632);
and U32081 (N_32081,N_31514,N_31770);
xor U32082 (N_32082,N_31547,N_31816);
nand U32083 (N_32083,N_31592,N_31814);
and U32084 (N_32084,N_31950,N_31778);
and U32085 (N_32085,N_31591,N_31935);
nand U32086 (N_32086,N_31981,N_31828);
nand U32087 (N_32087,N_31538,N_31644);
and U32088 (N_32088,N_31599,N_31678);
nand U32089 (N_32089,N_31875,N_31900);
and U32090 (N_32090,N_31809,N_31850);
nand U32091 (N_32091,N_31796,N_31892);
nand U32092 (N_32092,N_31604,N_31903);
or U32093 (N_32093,N_31991,N_31554);
xor U32094 (N_32094,N_31867,N_31569);
or U32095 (N_32095,N_31736,N_31813);
nand U32096 (N_32096,N_31721,N_31820);
or U32097 (N_32097,N_31777,N_31664);
nor U32098 (N_32098,N_31684,N_31621);
xnor U32099 (N_32099,N_31724,N_31541);
nor U32100 (N_32100,N_31706,N_31527);
nand U32101 (N_32101,N_31869,N_31556);
or U32102 (N_32102,N_31979,N_31803);
or U32103 (N_32103,N_31801,N_31836);
nor U32104 (N_32104,N_31831,N_31904);
nor U32105 (N_32105,N_31970,N_31613);
nand U32106 (N_32106,N_31985,N_31536);
nor U32107 (N_32107,N_31782,N_31690);
and U32108 (N_32108,N_31984,N_31918);
xnor U32109 (N_32109,N_31655,N_31618);
nand U32110 (N_32110,N_31815,N_31628);
xnor U32111 (N_32111,N_31609,N_31587);
nand U32112 (N_32112,N_31615,N_31823);
or U32113 (N_32113,N_31728,N_31794);
and U32114 (N_32114,N_31543,N_31668);
xor U32115 (N_32115,N_31840,N_31520);
nor U32116 (N_32116,N_31862,N_31766);
nor U32117 (N_32117,N_31932,N_31860);
and U32118 (N_32118,N_31959,N_31663);
xor U32119 (N_32119,N_31765,N_31600);
and U32120 (N_32120,N_31929,N_31666);
and U32121 (N_32121,N_31509,N_31913);
xnor U32122 (N_32122,N_31960,N_31641);
xor U32123 (N_32123,N_31893,N_31934);
or U32124 (N_32124,N_31881,N_31953);
nor U32125 (N_32125,N_31846,N_31745);
and U32126 (N_32126,N_31501,N_31756);
xor U32127 (N_32127,N_31549,N_31675);
or U32128 (N_32128,N_31635,N_31650);
xnor U32129 (N_32129,N_31646,N_31619);
nor U32130 (N_32130,N_31841,N_31544);
nor U32131 (N_32131,N_31806,N_31658);
or U32132 (N_32132,N_31947,N_31626);
nor U32133 (N_32133,N_31891,N_31722);
or U32134 (N_32134,N_31752,N_31882);
nor U32135 (N_32135,N_31738,N_31853);
xor U32136 (N_32136,N_31519,N_31692);
nand U32137 (N_32137,N_31905,N_31983);
nor U32138 (N_32138,N_31730,N_31605);
xnor U32139 (N_32139,N_31720,N_31817);
nand U32140 (N_32140,N_31617,N_31851);
and U32141 (N_32141,N_31837,N_31704);
or U32142 (N_32142,N_31917,N_31858);
xor U32143 (N_32143,N_31685,N_31945);
or U32144 (N_32144,N_31958,N_31924);
nand U32145 (N_32145,N_31894,N_31608);
xor U32146 (N_32146,N_31856,N_31537);
nand U32147 (N_32147,N_31754,N_31732);
nand U32148 (N_32148,N_31614,N_31557);
xnor U32149 (N_32149,N_31996,N_31741);
and U32150 (N_32150,N_31534,N_31768);
nand U32151 (N_32151,N_31933,N_31524);
or U32152 (N_32152,N_31631,N_31643);
nand U32153 (N_32153,N_31622,N_31672);
and U32154 (N_32154,N_31682,N_31956);
nand U32155 (N_32155,N_31698,N_31997);
or U32156 (N_32156,N_31938,N_31713);
xor U32157 (N_32157,N_31687,N_31819);
or U32158 (N_32158,N_31912,N_31560);
nor U32159 (N_32159,N_31928,N_31546);
nand U32160 (N_32160,N_31665,N_31598);
nor U32161 (N_32161,N_31673,N_31948);
xnor U32162 (N_32162,N_31545,N_31769);
and U32163 (N_32163,N_31757,N_31733);
xor U32164 (N_32164,N_31911,N_31726);
xor U32165 (N_32165,N_31797,N_31574);
or U32166 (N_32166,N_31596,N_31679);
or U32167 (N_32167,N_31968,N_31504);
or U32168 (N_32168,N_31735,N_31651);
nand U32169 (N_32169,N_31590,N_31982);
nor U32170 (N_32170,N_31880,N_31531);
nand U32171 (N_32171,N_31944,N_31670);
nor U32172 (N_32172,N_31879,N_31761);
nor U32173 (N_32173,N_31511,N_31998);
xor U32174 (N_32174,N_31994,N_31759);
and U32175 (N_32175,N_31688,N_31874);
nand U32176 (N_32176,N_31561,N_31727);
or U32177 (N_32177,N_31500,N_31977);
or U32178 (N_32178,N_31962,N_31876);
nand U32179 (N_32179,N_31895,N_31931);
and U32180 (N_32180,N_31582,N_31872);
or U32181 (N_32181,N_31755,N_31707);
nand U32182 (N_32182,N_31542,N_31516);
nand U32183 (N_32183,N_31919,N_31638);
nand U32184 (N_32184,N_31695,N_31973);
nand U32185 (N_32185,N_31999,N_31715);
nor U32186 (N_32186,N_31637,N_31612);
nand U32187 (N_32187,N_31680,N_31980);
nand U32188 (N_32188,N_31705,N_31772);
nor U32189 (N_32189,N_31585,N_31533);
xnor U32190 (N_32190,N_31844,N_31939);
or U32191 (N_32191,N_31583,N_31923);
and U32192 (N_32192,N_31683,N_31781);
nor U32193 (N_32193,N_31915,N_31965);
or U32194 (N_32194,N_31657,N_31804);
or U32195 (N_32195,N_31775,N_31955);
or U32196 (N_32196,N_31937,N_31901);
or U32197 (N_32197,N_31744,N_31624);
and U32198 (N_32198,N_31623,N_31576);
or U32199 (N_32199,N_31512,N_31589);
nand U32200 (N_32200,N_31878,N_31795);
nand U32201 (N_32201,N_31863,N_31660);
xor U32202 (N_32202,N_31636,N_31897);
xnor U32203 (N_32203,N_31886,N_31957);
nor U32204 (N_32204,N_31647,N_31921);
and U32205 (N_32205,N_31762,N_31780);
nand U32206 (N_32206,N_31826,N_31976);
nor U32207 (N_32207,N_31743,N_31839);
xor U32208 (N_32208,N_31523,N_31659);
nand U32209 (N_32209,N_31783,N_31729);
and U32210 (N_32210,N_31854,N_31691);
nor U32211 (N_32211,N_31510,N_31539);
nor U32212 (N_32212,N_31518,N_31972);
or U32213 (N_32213,N_31871,N_31829);
xor U32214 (N_32214,N_31522,N_31567);
xor U32215 (N_32215,N_31718,N_31771);
or U32216 (N_32216,N_31908,N_31902);
and U32217 (N_32217,N_31838,N_31633);
nand U32218 (N_32218,N_31739,N_31785);
nor U32219 (N_32219,N_31852,N_31961);
nand U32220 (N_32220,N_31606,N_31581);
or U32221 (N_32221,N_31717,N_31725);
nor U32222 (N_32222,N_31503,N_31812);
and U32223 (N_32223,N_31530,N_31562);
nor U32224 (N_32224,N_31978,N_31602);
or U32225 (N_32225,N_31528,N_31792);
nor U32226 (N_32226,N_31864,N_31855);
nand U32227 (N_32227,N_31563,N_31711);
nand U32228 (N_32228,N_31952,N_31989);
nor U32229 (N_32229,N_31597,N_31577);
xnor U32230 (N_32230,N_31566,N_31551);
and U32231 (N_32231,N_31789,N_31791);
nand U32232 (N_32232,N_31790,N_31870);
nor U32233 (N_32233,N_31710,N_31906);
nor U32234 (N_32234,N_31832,N_31669);
xor U32235 (N_32235,N_31558,N_31552);
nor U32236 (N_32236,N_31656,N_31674);
nand U32237 (N_32237,N_31603,N_31811);
nor U32238 (N_32238,N_31941,N_31857);
nor U32239 (N_32239,N_31573,N_31620);
and U32240 (N_32240,N_31927,N_31742);
nand U32241 (N_32241,N_31568,N_31899);
nor U32242 (N_32242,N_31877,N_31712);
and U32243 (N_32243,N_31653,N_31748);
nand U32244 (N_32244,N_31843,N_31883);
and U32245 (N_32245,N_31737,N_31764);
xnor U32246 (N_32246,N_31521,N_31971);
nor U32247 (N_32247,N_31995,N_31859);
nor U32248 (N_32248,N_31914,N_31507);
xnor U32249 (N_32249,N_31723,N_31714);
or U32250 (N_32250,N_31957,N_31765);
and U32251 (N_32251,N_31630,N_31829);
nand U32252 (N_32252,N_31993,N_31590);
or U32253 (N_32253,N_31956,N_31710);
or U32254 (N_32254,N_31533,N_31519);
or U32255 (N_32255,N_31590,N_31834);
nor U32256 (N_32256,N_31918,N_31743);
nor U32257 (N_32257,N_31974,N_31648);
nor U32258 (N_32258,N_31602,N_31588);
nand U32259 (N_32259,N_31914,N_31838);
and U32260 (N_32260,N_31643,N_31627);
nand U32261 (N_32261,N_31986,N_31522);
nand U32262 (N_32262,N_31901,N_31593);
xor U32263 (N_32263,N_31836,N_31560);
nor U32264 (N_32264,N_31658,N_31903);
or U32265 (N_32265,N_31617,N_31738);
nor U32266 (N_32266,N_31649,N_31901);
nor U32267 (N_32267,N_31516,N_31540);
or U32268 (N_32268,N_31779,N_31645);
and U32269 (N_32269,N_31887,N_31578);
nand U32270 (N_32270,N_31536,N_31629);
xor U32271 (N_32271,N_31723,N_31509);
nor U32272 (N_32272,N_31886,N_31767);
nor U32273 (N_32273,N_31649,N_31589);
xor U32274 (N_32274,N_31850,N_31773);
or U32275 (N_32275,N_31922,N_31572);
or U32276 (N_32276,N_31730,N_31810);
or U32277 (N_32277,N_31562,N_31792);
and U32278 (N_32278,N_31988,N_31670);
nor U32279 (N_32279,N_31826,N_31937);
nor U32280 (N_32280,N_31962,N_31987);
xor U32281 (N_32281,N_31721,N_31933);
xor U32282 (N_32282,N_31604,N_31992);
nor U32283 (N_32283,N_31817,N_31762);
nand U32284 (N_32284,N_31599,N_31676);
nor U32285 (N_32285,N_31742,N_31814);
and U32286 (N_32286,N_31511,N_31971);
nand U32287 (N_32287,N_31743,N_31563);
nor U32288 (N_32288,N_31954,N_31785);
nor U32289 (N_32289,N_31560,N_31800);
or U32290 (N_32290,N_31983,N_31991);
nand U32291 (N_32291,N_31986,N_31541);
xnor U32292 (N_32292,N_31569,N_31714);
and U32293 (N_32293,N_31842,N_31991);
xor U32294 (N_32294,N_31993,N_31889);
and U32295 (N_32295,N_31646,N_31721);
and U32296 (N_32296,N_31731,N_31704);
or U32297 (N_32297,N_31516,N_31987);
or U32298 (N_32298,N_31932,N_31941);
nand U32299 (N_32299,N_31515,N_31765);
and U32300 (N_32300,N_31857,N_31776);
nand U32301 (N_32301,N_31767,N_31784);
xnor U32302 (N_32302,N_31808,N_31875);
and U32303 (N_32303,N_31995,N_31524);
or U32304 (N_32304,N_31603,N_31791);
or U32305 (N_32305,N_31759,N_31560);
and U32306 (N_32306,N_31725,N_31790);
xnor U32307 (N_32307,N_31979,N_31599);
and U32308 (N_32308,N_31888,N_31517);
xnor U32309 (N_32309,N_31879,N_31575);
nand U32310 (N_32310,N_31829,N_31885);
and U32311 (N_32311,N_31719,N_31518);
nor U32312 (N_32312,N_31715,N_31845);
nor U32313 (N_32313,N_31884,N_31518);
and U32314 (N_32314,N_31576,N_31569);
and U32315 (N_32315,N_31778,N_31712);
nor U32316 (N_32316,N_31970,N_31835);
or U32317 (N_32317,N_31751,N_31515);
nor U32318 (N_32318,N_31926,N_31898);
nor U32319 (N_32319,N_31861,N_31849);
xor U32320 (N_32320,N_31534,N_31575);
nor U32321 (N_32321,N_31587,N_31826);
or U32322 (N_32322,N_31617,N_31849);
nor U32323 (N_32323,N_31896,N_31526);
nor U32324 (N_32324,N_31795,N_31712);
nor U32325 (N_32325,N_31870,N_31822);
nand U32326 (N_32326,N_31700,N_31679);
nand U32327 (N_32327,N_31840,N_31945);
xor U32328 (N_32328,N_31810,N_31744);
or U32329 (N_32329,N_31811,N_31707);
xor U32330 (N_32330,N_31573,N_31924);
xor U32331 (N_32331,N_31521,N_31638);
nand U32332 (N_32332,N_31637,N_31781);
xor U32333 (N_32333,N_31713,N_31721);
nor U32334 (N_32334,N_31586,N_31837);
or U32335 (N_32335,N_31862,N_31984);
or U32336 (N_32336,N_31648,N_31643);
xor U32337 (N_32337,N_31556,N_31939);
xnor U32338 (N_32338,N_31617,N_31615);
or U32339 (N_32339,N_31787,N_31858);
or U32340 (N_32340,N_31669,N_31999);
nor U32341 (N_32341,N_31732,N_31635);
and U32342 (N_32342,N_31793,N_31665);
xor U32343 (N_32343,N_31733,N_31958);
or U32344 (N_32344,N_31911,N_31712);
xor U32345 (N_32345,N_31735,N_31961);
and U32346 (N_32346,N_31616,N_31809);
nor U32347 (N_32347,N_31793,N_31615);
nand U32348 (N_32348,N_31847,N_31624);
nand U32349 (N_32349,N_31503,N_31943);
nor U32350 (N_32350,N_31870,N_31852);
nor U32351 (N_32351,N_31749,N_31930);
and U32352 (N_32352,N_31540,N_31849);
xor U32353 (N_32353,N_31547,N_31871);
or U32354 (N_32354,N_31642,N_31699);
xnor U32355 (N_32355,N_31736,N_31571);
nor U32356 (N_32356,N_31919,N_31711);
or U32357 (N_32357,N_31967,N_31924);
or U32358 (N_32358,N_31660,N_31864);
nand U32359 (N_32359,N_31682,N_31787);
and U32360 (N_32360,N_31804,N_31589);
and U32361 (N_32361,N_31946,N_31854);
and U32362 (N_32362,N_31830,N_31600);
xor U32363 (N_32363,N_31678,N_31830);
xor U32364 (N_32364,N_31799,N_31965);
and U32365 (N_32365,N_31712,N_31924);
xor U32366 (N_32366,N_31706,N_31687);
or U32367 (N_32367,N_31781,N_31531);
or U32368 (N_32368,N_31693,N_31776);
or U32369 (N_32369,N_31660,N_31798);
or U32370 (N_32370,N_31584,N_31892);
and U32371 (N_32371,N_31923,N_31659);
or U32372 (N_32372,N_31955,N_31623);
and U32373 (N_32373,N_31698,N_31542);
and U32374 (N_32374,N_31936,N_31946);
nand U32375 (N_32375,N_31823,N_31757);
xnor U32376 (N_32376,N_31625,N_31682);
nand U32377 (N_32377,N_31775,N_31808);
nor U32378 (N_32378,N_31605,N_31566);
xnor U32379 (N_32379,N_31520,N_31995);
nor U32380 (N_32380,N_31845,N_31900);
and U32381 (N_32381,N_31840,N_31796);
and U32382 (N_32382,N_31921,N_31643);
nand U32383 (N_32383,N_31792,N_31859);
xnor U32384 (N_32384,N_31547,N_31930);
nor U32385 (N_32385,N_31571,N_31780);
and U32386 (N_32386,N_31885,N_31782);
or U32387 (N_32387,N_31778,N_31718);
nand U32388 (N_32388,N_31928,N_31643);
xnor U32389 (N_32389,N_31638,N_31664);
and U32390 (N_32390,N_31617,N_31846);
and U32391 (N_32391,N_31589,N_31794);
xor U32392 (N_32392,N_31835,N_31796);
nor U32393 (N_32393,N_31589,N_31800);
and U32394 (N_32394,N_31767,N_31609);
nor U32395 (N_32395,N_31775,N_31724);
nand U32396 (N_32396,N_31856,N_31760);
and U32397 (N_32397,N_31957,N_31772);
and U32398 (N_32398,N_31507,N_31953);
or U32399 (N_32399,N_31667,N_31735);
or U32400 (N_32400,N_31879,N_31528);
xor U32401 (N_32401,N_31930,N_31536);
nor U32402 (N_32402,N_31817,N_31982);
nand U32403 (N_32403,N_31659,N_31707);
or U32404 (N_32404,N_31821,N_31628);
and U32405 (N_32405,N_31509,N_31696);
and U32406 (N_32406,N_31754,N_31960);
or U32407 (N_32407,N_31659,N_31798);
or U32408 (N_32408,N_31538,N_31961);
nand U32409 (N_32409,N_31523,N_31516);
nand U32410 (N_32410,N_31717,N_31659);
xor U32411 (N_32411,N_31674,N_31891);
nor U32412 (N_32412,N_31612,N_31764);
xnor U32413 (N_32413,N_31870,N_31946);
nand U32414 (N_32414,N_31938,N_31568);
and U32415 (N_32415,N_31751,N_31851);
nand U32416 (N_32416,N_31853,N_31947);
nor U32417 (N_32417,N_31570,N_31520);
and U32418 (N_32418,N_31651,N_31879);
nor U32419 (N_32419,N_31939,N_31717);
or U32420 (N_32420,N_31632,N_31682);
and U32421 (N_32421,N_31910,N_31774);
nand U32422 (N_32422,N_31933,N_31541);
xor U32423 (N_32423,N_31609,N_31622);
nand U32424 (N_32424,N_31996,N_31688);
xnor U32425 (N_32425,N_31516,N_31613);
xor U32426 (N_32426,N_31737,N_31795);
nor U32427 (N_32427,N_31957,N_31971);
or U32428 (N_32428,N_31850,N_31960);
nor U32429 (N_32429,N_31844,N_31613);
nor U32430 (N_32430,N_31679,N_31901);
and U32431 (N_32431,N_31748,N_31787);
xor U32432 (N_32432,N_31970,N_31645);
or U32433 (N_32433,N_31822,N_31525);
nor U32434 (N_32434,N_31739,N_31762);
nor U32435 (N_32435,N_31668,N_31739);
nor U32436 (N_32436,N_31786,N_31992);
nand U32437 (N_32437,N_31973,N_31909);
and U32438 (N_32438,N_31662,N_31844);
and U32439 (N_32439,N_31912,N_31630);
nor U32440 (N_32440,N_31902,N_31761);
or U32441 (N_32441,N_31690,N_31820);
nor U32442 (N_32442,N_31584,N_31874);
or U32443 (N_32443,N_31687,N_31762);
nor U32444 (N_32444,N_31593,N_31684);
xor U32445 (N_32445,N_31951,N_31809);
xor U32446 (N_32446,N_31671,N_31792);
and U32447 (N_32447,N_31893,N_31557);
nor U32448 (N_32448,N_31878,N_31542);
and U32449 (N_32449,N_31619,N_31591);
nor U32450 (N_32450,N_31703,N_31888);
nor U32451 (N_32451,N_31986,N_31774);
xnor U32452 (N_32452,N_31595,N_31793);
or U32453 (N_32453,N_31583,N_31755);
nand U32454 (N_32454,N_31594,N_31750);
xor U32455 (N_32455,N_31859,N_31915);
nor U32456 (N_32456,N_31956,N_31622);
and U32457 (N_32457,N_31785,N_31641);
or U32458 (N_32458,N_31922,N_31682);
nor U32459 (N_32459,N_31839,N_31899);
nand U32460 (N_32460,N_31841,N_31764);
and U32461 (N_32461,N_31567,N_31544);
and U32462 (N_32462,N_31647,N_31639);
and U32463 (N_32463,N_31746,N_31664);
xnor U32464 (N_32464,N_31893,N_31924);
nand U32465 (N_32465,N_31987,N_31809);
nand U32466 (N_32466,N_31754,N_31658);
nand U32467 (N_32467,N_31664,N_31621);
nand U32468 (N_32468,N_31532,N_31662);
xor U32469 (N_32469,N_31928,N_31719);
or U32470 (N_32470,N_31781,N_31771);
nand U32471 (N_32471,N_31590,N_31752);
xnor U32472 (N_32472,N_31586,N_31849);
and U32473 (N_32473,N_31839,N_31762);
xnor U32474 (N_32474,N_31795,N_31970);
and U32475 (N_32475,N_31650,N_31771);
nand U32476 (N_32476,N_31930,N_31843);
nand U32477 (N_32477,N_31933,N_31690);
nor U32478 (N_32478,N_31751,N_31861);
or U32479 (N_32479,N_31518,N_31902);
nand U32480 (N_32480,N_31667,N_31807);
xor U32481 (N_32481,N_31773,N_31728);
nand U32482 (N_32482,N_31600,N_31695);
and U32483 (N_32483,N_31676,N_31644);
nor U32484 (N_32484,N_31579,N_31500);
or U32485 (N_32485,N_31512,N_31936);
and U32486 (N_32486,N_31817,N_31535);
nand U32487 (N_32487,N_31709,N_31611);
and U32488 (N_32488,N_31998,N_31769);
xor U32489 (N_32489,N_31842,N_31746);
nor U32490 (N_32490,N_31689,N_31572);
nand U32491 (N_32491,N_31735,N_31979);
xor U32492 (N_32492,N_31723,N_31923);
or U32493 (N_32493,N_31765,N_31901);
xnor U32494 (N_32494,N_31725,N_31718);
and U32495 (N_32495,N_31778,N_31765);
nor U32496 (N_32496,N_31542,N_31764);
xor U32497 (N_32497,N_31991,N_31922);
or U32498 (N_32498,N_31934,N_31958);
nand U32499 (N_32499,N_31844,N_31969);
nand U32500 (N_32500,N_32209,N_32386);
nand U32501 (N_32501,N_32028,N_32311);
and U32502 (N_32502,N_32148,N_32272);
nand U32503 (N_32503,N_32071,N_32492);
xnor U32504 (N_32504,N_32411,N_32099);
nor U32505 (N_32505,N_32254,N_32076);
or U32506 (N_32506,N_32290,N_32265);
or U32507 (N_32507,N_32193,N_32202);
xor U32508 (N_32508,N_32096,N_32287);
or U32509 (N_32509,N_32298,N_32068);
or U32510 (N_32510,N_32084,N_32266);
nand U32511 (N_32511,N_32032,N_32332);
xor U32512 (N_32512,N_32486,N_32156);
nor U32513 (N_32513,N_32297,N_32334);
xnor U32514 (N_32514,N_32027,N_32374);
xor U32515 (N_32515,N_32181,N_32228);
nor U32516 (N_32516,N_32475,N_32200);
or U32517 (N_32517,N_32196,N_32367);
xnor U32518 (N_32518,N_32155,N_32350);
xor U32519 (N_32519,N_32264,N_32031);
or U32520 (N_32520,N_32442,N_32192);
xnor U32521 (N_32521,N_32410,N_32142);
nor U32522 (N_32522,N_32414,N_32044);
xnor U32523 (N_32523,N_32391,N_32095);
or U32524 (N_32524,N_32303,N_32314);
or U32525 (N_32525,N_32070,N_32212);
or U32526 (N_32526,N_32307,N_32319);
and U32527 (N_32527,N_32333,N_32115);
xnor U32528 (N_32528,N_32432,N_32122);
nor U32529 (N_32529,N_32140,N_32448);
or U32530 (N_32530,N_32178,N_32098);
nand U32531 (N_32531,N_32168,N_32481);
or U32532 (N_32532,N_32129,N_32388);
and U32533 (N_32533,N_32464,N_32474);
xor U32534 (N_32534,N_32006,N_32009);
nand U32535 (N_32535,N_32273,N_32284);
or U32536 (N_32536,N_32083,N_32351);
nand U32537 (N_32537,N_32127,N_32400);
or U32538 (N_32538,N_32439,N_32016);
nand U32539 (N_32539,N_32222,N_32438);
or U32540 (N_32540,N_32053,N_32208);
nand U32541 (N_32541,N_32104,N_32450);
or U32542 (N_32542,N_32288,N_32420);
or U32543 (N_32543,N_32153,N_32326);
xnor U32544 (N_32544,N_32226,N_32357);
and U32545 (N_32545,N_32496,N_32361);
or U32546 (N_32546,N_32130,N_32460);
or U32547 (N_32547,N_32281,N_32433);
nor U32548 (N_32548,N_32154,N_32426);
xnor U32549 (N_32549,N_32413,N_32395);
nor U32550 (N_32550,N_32171,N_32063);
and U32551 (N_32551,N_32493,N_32262);
and U32552 (N_32552,N_32211,N_32416);
and U32553 (N_32553,N_32124,N_32052);
and U32554 (N_32554,N_32335,N_32371);
nand U32555 (N_32555,N_32141,N_32235);
or U32556 (N_32556,N_32424,N_32404);
and U32557 (N_32557,N_32369,N_32091);
xor U32558 (N_32558,N_32189,N_32223);
nand U32559 (N_32559,N_32205,N_32469);
and U32560 (N_32560,N_32406,N_32293);
nand U32561 (N_32561,N_32139,N_32067);
or U32562 (N_32562,N_32112,N_32034);
or U32563 (N_32563,N_32259,N_32373);
xnor U32564 (N_32564,N_32055,N_32106);
nand U32565 (N_32565,N_32147,N_32356);
nor U32566 (N_32566,N_32051,N_32399);
xnor U32567 (N_32567,N_32385,N_32221);
nand U32568 (N_32568,N_32392,N_32118);
or U32569 (N_32569,N_32338,N_32304);
nor U32570 (N_32570,N_32394,N_32283);
nor U32571 (N_32571,N_32230,N_32313);
nand U32572 (N_32572,N_32092,N_32453);
or U32573 (N_32573,N_32479,N_32436);
or U32574 (N_32574,N_32489,N_32383);
nand U32575 (N_32575,N_32049,N_32037);
nor U32576 (N_32576,N_32138,N_32462);
nor U32577 (N_32577,N_32123,N_32372);
or U32578 (N_32578,N_32471,N_32217);
and U32579 (N_32579,N_32105,N_32024);
xor U32580 (N_32580,N_32419,N_32163);
nor U32581 (N_32581,N_32340,N_32275);
nor U32582 (N_32582,N_32476,N_32250);
or U32583 (N_32583,N_32289,N_32446);
nand U32584 (N_32584,N_32403,N_32463);
xor U32585 (N_32585,N_32415,N_32447);
xnor U32586 (N_32586,N_32176,N_32276);
and U32587 (N_32587,N_32038,N_32482);
xnor U32588 (N_32588,N_32239,N_32256);
or U32589 (N_32589,N_32322,N_32498);
nor U32590 (N_32590,N_32429,N_32327);
and U32591 (N_32591,N_32255,N_32260);
nor U32592 (N_32592,N_32454,N_32062);
or U32593 (N_32593,N_32103,N_32491);
nor U32594 (N_32594,N_32179,N_32384);
and U32595 (N_32595,N_32258,N_32337);
nor U32596 (N_32596,N_32309,N_32180);
nand U32597 (N_32597,N_32162,N_32245);
and U32598 (N_32598,N_32146,N_32300);
and U32599 (N_32599,N_32191,N_32198);
and U32600 (N_32600,N_32321,N_32025);
xor U32601 (N_32601,N_32190,N_32261);
and U32602 (N_32602,N_32003,N_32241);
or U32603 (N_32603,N_32020,N_32015);
nor U32604 (N_32604,N_32030,N_32380);
xor U32605 (N_32605,N_32390,N_32008);
xor U32606 (N_32606,N_32472,N_32299);
or U32607 (N_32607,N_32182,N_32434);
or U32608 (N_32608,N_32359,N_32295);
nor U32609 (N_32609,N_32194,N_32381);
and U32610 (N_32610,N_32349,N_32080);
xor U32611 (N_32611,N_32231,N_32086);
nand U32612 (N_32612,N_32488,N_32160);
and U32613 (N_32613,N_32000,N_32011);
nor U32614 (N_32614,N_32277,N_32294);
nor U32615 (N_32615,N_32401,N_32487);
nand U32616 (N_32616,N_32341,N_32477);
and U32617 (N_32617,N_32285,N_32204);
xor U32618 (N_32618,N_32085,N_32268);
xnor U32619 (N_32619,N_32173,N_32207);
and U32620 (N_32620,N_32117,N_32111);
and U32621 (N_32621,N_32210,N_32312);
and U32622 (N_32622,N_32169,N_32177);
xor U32623 (N_32623,N_32377,N_32150);
nand U32624 (N_32624,N_32278,N_32004);
and U32625 (N_32625,N_32119,N_32135);
xor U32626 (N_32626,N_32417,N_32010);
and U32627 (N_32627,N_32232,N_32336);
xnor U32628 (N_32628,N_32056,N_32065);
nor U32629 (N_32629,N_32184,N_32376);
or U32630 (N_32630,N_32305,N_32490);
nand U32631 (N_32631,N_32005,N_32183);
nor U32632 (N_32632,N_32343,N_32286);
or U32633 (N_32633,N_32317,N_32402);
nor U32634 (N_32634,N_32240,N_32218);
and U32635 (N_32635,N_32346,N_32279);
and U32636 (N_32636,N_32257,N_32214);
and U32637 (N_32637,N_32133,N_32165);
or U32638 (N_32638,N_32244,N_32195);
nand U32639 (N_32639,N_32347,N_32363);
nor U32640 (N_32640,N_32220,N_32170);
and U32641 (N_32641,N_32345,N_32012);
and U32642 (N_32642,N_32368,N_32328);
and U32643 (N_32643,N_32048,N_32430);
or U32644 (N_32644,N_32267,N_32074);
xor U32645 (N_32645,N_32451,N_32435);
and U32646 (N_32646,N_32444,N_32301);
xnor U32647 (N_32647,N_32175,N_32078);
or U32648 (N_32648,N_32422,N_32023);
nand U32649 (N_32649,N_32473,N_32470);
or U32650 (N_32650,N_32242,N_32465);
xor U32651 (N_32651,N_32131,N_32229);
nand U32652 (N_32652,N_32249,N_32431);
nand U32653 (N_32653,N_32282,N_32269);
xor U32654 (N_32654,N_32437,N_32354);
xor U32655 (N_32655,N_32029,N_32466);
xnor U32656 (N_32656,N_32246,N_32227);
or U32657 (N_32657,N_32152,N_32039);
nand U32658 (N_32658,N_32019,N_32291);
nand U32659 (N_32659,N_32238,N_32485);
and U32660 (N_32660,N_32398,N_32443);
xnor U32661 (N_32661,N_32233,N_32329);
nor U32662 (N_32662,N_32188,N_32461);
nand U32663 (N_32663,N_32046,N_32126);
nand U32664 (N_32664,N_32405,N_32128);
nand U32665 (N_32665,N_32379,N_32237);
nand U32666 (N_32666,N_32330,N_32325);
nand U32667 (N_32667,N_32088,N_32280);
or U32668 (N_32668,N_32136,N_32108);
and U32669 (N_32669,N_32213,N_32144);
nor U32670 (N_32670,N_32478,N_32166);
xnor U32671 (N_32671,N_32393,N_32263);
nor U32672 (N_32672,N_32035,N_32007);
nand U32673 (N_32673,N_32145,N_32164);
nand U32674 (N_32674,N_32225,N_32236);
xor U32675 (N_32675,N_32054,N_32132);
nor U32676 (N_32676,N_32066,N_32042);
and U32677 (N_32677,N_32089,N_32320);
and U32678 (N_32678,N_32059,N_32362);
or U32679 (N_32679,N_32499,N_32247);
and U32680 (N_32680,N_32026,N_32483);
nor U32681 (N_32681,N_32075,N_32445);
or U32682 (N_32682,N_32014,N_32043);
and U32683 (N_32683,N_32159,N_32370);
or U32684 (N_32684,N_32428,N_32318);
or U32685 (N_32685,N_32073,N_32036);
nor U32686 (N_32686,N_32495,N_32352);
xnor U32687 (N_32687,N_32077,N_32125);
nand U32688 (N_32688,N_32358,N_32100);
xor U32689 (N_32689,N_32167,N_32033);
nor U32690 (N_32690,N_32355,N_32187);
nor U32691 (N_32691,N_32064,N_32151);
xnor U32692 (N_32692,N_32243,N_32107);
nand U32693 (N_32693,N_32081,N_32441);
and U32694 (N_32694,N_32079,N_32018);
nand U32695 (N_32695,N_32480,N_32050);
or U32696 (N_32696,N_32497,N_32093);
xnor U32697 (N_32697,N_32041,N_32484);
xor U32698 (N_32698,N_32094,N_32387);
nor U32699 (N_32699,N_32101,N_32001);
and U32700 (N_32700,N_32186,N_32425);
or U32701 (N_32701,N_32348,N_32324);
nor U32702 (N_32702,N_32114,N_32270);
nand U32703 (N_32703,N_32072,N_32468);
nor U32704 (N_32704,N_32271,N_32360);
and U32705 (N_32705,N_32331,N_32134);
nor U32706 (N_32706,N_32409,N_32344);
xor U32707 (N_32707,N_32274,N_32455);
nor U32708 (N_32708,N_32057,N_32494);
nand U32709 (N_32709,N_32199,N_32161);
or U32710 (N_32710,N_32109,N_32407);
nand U32711 (N_32711,N_32102,N_32292);
nand U32712 (N_32712,N_32197,N_32013);
and U32713 (N_32713,N_32069,N_32060);
nand U32714 (N_32714,N_32158,N_32467);
nand U32715 (N_32715,N_32339,N_32234);
and U32716 (N_32716,N_32206,N_32157);
and U32717 (N_32717,N_32253,N_32408);
or U32718 (N_32718,N_32306,N_32389);
and U32719 (N_32719,N_32087,N_32456);
or U32720 (N_32720,N_32113,N_32397);
xor U32721 (N_32721,N_32047,N_32452);
and U32722 (N_32722,N_32308,N_32045);
and U32723 (N_32723,N_32396,N_32412);
and U32724 (N_32724,N_32017,N_32382);
and U32725 (N_32725,N_32040,N_32224);
nor U32726 (N_32726,N_32310,N_32061);
or U32727 (N_32727,N_32248,N_32219);
nor U32728 (N_32728,N_32058,N_32427);
xnor U32729 (N_32729,N_32143,N_32116);
nor U32730 (N_32730,N_32353,N_32203);
and U32731 (N_32731,N_32201,N_32364);
nand U32732 (N_32732,N_32216,N_32323);
nor U32733 (N_32733,N_32458,N_32366);
nand U32734 (N_32734,N_32090,N_32002);
and U32735 (N_32735,N_32021,N_32149);
xor U32736 (N_32736,N_32185,N_32440);
or U32737 (N_32737,N_32365,N_32449);
xor U32738 (N_32738,N_32423,N_32421);
nor U32739 (N_32739,N_32121,N_32252);
nand U32740 (N_32740,N_32137,N_32110);
and U32741 (N_32741,N_32097,N_32302);
or U32742 (N_32742,N_32316,N_32174);
or U32743 (N_32743,N_32457,N_32315);
nor U32744 (N_32744,N_32375,N_32215);
or U32745 (N_32745,N_32418,N_32296);
xnor U32746 (N_32746,N_32082,N_32378);
or U32747 (N_32747,N_32172,N_32022);
or U32748 (N_32748,N_32251,N_32342);
xor U32749 (N_32749,N_32459,N_32120);
and U32750 (N_32750,N_32431,N_32118);
xnor U32751 (N_32751,N_32224,N_32226);
or U32752 (N_32752,N_32333,N_32191);
and U32753 (N_32753,N_32027,N_32480);
xnor U32754 (N_32754,N_32190,N_32128);
nor U32755 (N_32755,N_32393,N_32405);
and U32756 (N_32756,N_32013,N_32082);
or U32757 (N_32757,N_32449,N_32484);
xnor U32758 (N_32758,N_32228,N_32357);
nor U32759 (N_32759,N_32255,N_32331);
xor U32760 (N_32760,N_32252,N_32013);
and U32761 (N_32761,N_32050,N_32108);
nor U32762 (N_32762,N_32271,N_32133);
nand U32763 (N_32763,N_32469,N_32347);
nor U32764 (N_32764,N_32154,N_32344);
xnor U32765 (N_32765,N_32012,N_32059);
or U32766 (N_32766,N_32325,N_32271);
nand U32767 (N_32767,N_32321,N_32302);
or U32768 (N_32768,N_32186,N_32479);
or U32769 (N_32769,N_32181,N_32345);
nand U32770 (N_32770,N_32402,N_32108);
nor U32771 (N_32771,N_32138,N_32226);
nor U32772 (N_32772,N_32393,N_32350);
and U32773 (N_32773,N_32000,N_32113);
xor U32774 (N_32774,N_32029,N_32290);
nand U32775 (N_32775,N_32101,N_32390);
xor U32776 (N_32776,N_32013,N_32440);
nor U32777 (N_32777,N_32415,N_32463);
and U32778 (N_32778,N_32175,N_32041);
xor U32779 (N_32779,N_32190,N_32249);
or U32780 (N_32780,N_32044,N_32332);
and U32781 (N_32781,N_32369,N_32279);
nor U32782 (N_32782,N_32400,N_32042);
or U32783 (N_32783,N_32162,N_32434);
or U32784 (N_32784,N_32256,N_32416);
and U32785 (N_32785,N_32330,N_32155);
xnor U32786 (N_32786,N_32187,N_32485);
or U32787 (N_32787,N_32495,N_32173);
nor U32788 (N_32788,N_32419,N_32147);
nand U32789 (N_32789,N_32388,N_32449);
nand U32790 (N_32790,N_32443,N_32067);
and U32791 (N_32791,N_32402,N_32182);
or U32792 (N_32792,N_32136,N_32393);
nand U32793 (N_32793,N_32078,N_32428);
xnor U32794 (N_32794,N_32229,N_32056);
nand U32795 (N_32795,N_32243,N_32066);
and U32796 (N_32796,N_32048,N_32338);
nor U32797 (N_32797,N_32262,N_32004);
xnor U32798 (N_32798,N_32431,N_32257);
and U32799 (N_32799,N_32093,N_32377);
or U32800 (N_32800,N_32156,N_32271);
and U32801 (N_32801,N_32464,N_32386);
nand U32802 (N_32802,N_32301,N_32156);
xnor U32803 (N_32803,N_32424,N_32124);
or U32804 (N_32804,N_32039,N_32174);
nand U32805 (N_32805,N_32005,N_32432);
nor U32806 (N_32806,N_32020,N_32144);
or U32807 (N_32807,N_32211,N_32361);
or U32808 (N_32808,N_32421,N_32279);
or U32809 (N_32809,N_32085,N_32471);
or U32810 (N_32810,N_32482,N_32148);
or U32811 (N_32811,N_32192,N_32392);
nand U32812 (N_32812,N_32411,N_32270);
or U32813 (N_32813,N_32080,N_32100);
or U32814 (N_32814,N_32066,N_32115);
and U32815 (N_32815,N_32257,N_32320);
or U32816 (N_32816,N_32326,N_32183);
nand U32817 (N_32817,N_32441,N_32424);
or U32818 (N_32818,N_32498,N_32317);
or U32819 (N_32819,N_32285,N_32484);
and U32820 (N_32820,N_32163,N_32497);
nor U32821 (N_32821,N_32145,N_32139);
nor U32822 (N_32822,N_32201,N_32297);
nor U32823 (N_32823,N_32169,N_32402);
nor U32824 (N_32824,N_32348,N_32251);
nor U32825 (N_32825,N_32197,N_32149);
or U32826 (N_32826,N_32190,N_32286);
nor U32827 (N_32827,N_32085,N_32062);
or U32828 (N_32828,N_32466,N_32223);
and U32829 (N_32829,N_32097,N_32094);
and U32830 (N_32830,N_32158,N_32275);
and U32831 (N_32831,N_32013,N_32245);
nand U32832 (N_32832,N_32291,N_32324);
nand U32833 (N_32833,N_32093,N_32475);
or U32834 (N_32834,N_32484,N_32122);
xor U32835 (N_32835,N_32176,N_32106);
nand U32836 (N_32836,N_32180,N_32218);
nand U32837 (N_32837,N_32366,N_32274);
nor U32838 (N_32838,N_32025,N_32399);
or U32839 (N_32839,N_32021,N_32004);
nor U32840 (N_32840,N_32301,N_32036);
or U32841 (N_32841,N_32203,N_32110);
and U32842 (N_32842,N_32260,N_32212);
and U32843 (N_32843,N_32489,N_32399);
xnor U32844 (N_32844,N_32129,N_32201);
or U32845 (N_32845,N_32319,N_32221);
xor U32846 (N_32846,N_32241,N_32489);
nor U32847 (N_32847,N_32458,N_32474);
xor U32848 (N_32848,N_32014,N_32151);
or U32849 (N_32849,N_32064,N_32378);
and U32850 (N_32850,N_32148,N_32387);
and U32851 (N_32851,N_32182,N_32366);
xnor U32852 (N_32852,N_32276,N_32473);
or U32853 (N_32853,N_32283,N_32216);
nand U32854 (N_32854,N_32299,N_32099);
nor U32855 (N_32855,N_32155,N_32314);
and U32856 (N_32856,N_32442,N_32370);
and U32857 (N_32857,N_32469,N_32491);
or U32858 (N_32858,N_32343,N_32359);
and U32859 (N_32859,N_32117,N_32273);
nor U32860 (N_32860,N_32060,N_32275);
nand U32861 (N_32861,N_32371,N_32315);
or U32862 (N_32862,N_32163,N_32253);
nand U32863 (N_32863,N_32179,N_32020);
and U32864 (N_32864,N_32040,N_32344);
nor U32865 (N_32865,N_32126,N_32384);
nor U32866 (N_32866,N_32272,N_32428);
or U32867 (N_32867,N_32206,N_32066);
or U32868 (N_32868,N_32286,N_32098);
nor U32869 (N_32869,N_32000,N_32371);
and U32870 (N_32870,N_32154,N_32254);
nor U32871 (N_32871,N_32483,N_32404);
nand U32872 (N_32872,N_32174,N_32476);
nand U32873 (N_32873,N_32383,N_32228);
nand U32874 (N_32874,N_32128,N_32010);
or U32875 (N_32875,N_32346,N_32221);
xor U32876 (N_32876,N_32028,N_32485);
or U32877 (N_32877,N_32397,N_32345);
and U32878 (N_32878,N_32010,N_32484);
and U32879 (N_32879,N_32095,N_32189);
nand U32880 (N_32880,N_32469,N_32100);
xnor U32881 (N_32881,N_32438,N_32397);
nand U32882 (N_32882,N_32125,N_32404);
nor U32883 (N_32883,N_32199,N_32440);
and U32884 (N_32884,N_32490,N_32131);
nor U32885 (N_32885,N_32400,N_32448);
and U32886 (N_32886,N_32308,N_32105);
nand U32887 (N_32887,N_32374,N_32260);
xor U32888 (N_32888,N_32152,N_32147);
or U32889 (N_32889,N_32099,N_32169);
and U32890 (N_32890,N_32324,N_32336);
nand U32891 (N_32891,N_32150,N_32119);
nor U32892 (N_32892,N_32423,N_32120);
nand U32893 (N_32893,N_32465,N_32482);
nor U32894 (N_32894,N_32301,N_32327);
and U32895 (N_32895,N_32316,N_32327);
and U32896 (N_32896,N_32252,N_32091);
or U32897 (N_32897,N_32380,N_32001);
and U32898 (N_32898,N_32197,N_32365);
or U32899 (N_32899,N_32367,N_32255);
xnor U32900 (N_32900,N_32432,N_32121);
or U32901 (N_32901,N_32472,N_32159);
and U32902 (N_32902,N_32059,N_32471);
nand U32903 (N_32903,N_32021,N_32431);
and U32904 (N_32904,N_32054,N_32272);
and U32905 (N_32905,N_32017,N_32197);
and U32906 (N_32906,N_32144,N_32312);
xor U32907 (N_32907,N_32339,N_32305);
or U32908 (N_32908,N_32443,N_32422);
nor U32909 (N_32909,N_32039,N_32134);
xnor U32910 (N_32910,N_32061,N_32221);
nor U32911 (N_32911,N_32101,N_32135);
nand U32912 (N_32912,N_32142,N_32415);
or U32913 (N_32913,N_32425,N_32363);
xor U32914 (N_32914,N_32311,N_32018);
xor U32915 (N_32915,N_32332,N_32234);
nand U32916 (N_32916,N_32130,N_32285);
nand U32917 (N_32917,N_32090,N_32489);
nor U32918 (N_32918,N_32445,N_32175);
xor U32919 (N_32919,N_32380,N_32400);
xnor U32920 (N_32920,N_32278,N_32145);
xnor U32921 (N_32921,N_32181,N_32194);
nand U32922 (N_32922,N_32401,N_32310);
nor U32923 (N_32923,N_32079,N_32080);
xor U32924 (N_32924,N_32429,N_32469);
nor U32925 (N_32925,N_32077,N_32263);
or U32926 (N_32926,N_32034,N_32044);
or U32927 (N_32927,N_32373,N_32093);
and U32928 (N_32928,N_32489,N_32208);
xor U32929 (N_32929,N_32383,N_32248);
or U32930 (N_32930,N_32222,N_32100);
nand U32931 (N_32931,N_32127,N_32085);
or U32932 (N_32932,N_32211,N_32489);
or U32933 (N_32933,N_32199,N_32111);
xnor U32934 (N_32934,N_32385,N_32281);
nor U32935 (N_32935,N_32497,N_32466);
or U32936 (N_32936,N_32248,N_32243);
nor U32937 (N_32937,N_32015,N_32461);
nor U32938 (N_32938,N_32156,N_32160);
xnor U32939 (N_32939,N_32342,N_32111);
nand U32940 (N_32940,N_32380,N_32313);
nand U32941 (N_32941,N_32227,N_32350);
nand U32942 (N_32942,N_32480,N_32281);
xor U32943 (N_32943,N_32122,N_32321);
xnor U32944 (N_32944,N_32271,N_32335);
or U32945 (N_32945,N_32480,N_32040);
or U32946 (N_32946,N_32467,N_32237);
or U32947 (N_32947,N_32110,N_32023);
nand U32948 (N_32948,N_32353,N_32175);
or U32949 (N_32949,N_32246,N_32355);
xnor U32950 (N_32950,N_32058,N_32288);
xnor U32951 (N_32951,N_32079,N_32205);
nand U32952 (N_32952,N_32463,N_32165);
nand U32953 (N_32953,N_32207,N_32292);
nor U32954 (N_32954,N_32314,N_32183);
or U32955 (N_32955,N_32065,N_32220);
nor U32956 (N_32956,N_32266,N_32066);
nand U32957 (N_32957,N_32329,N_32135);
and U32958 (N_32958,N_32296,N_32462);
or U32959 (N_32959,N_32102,N_32066);
or U32960 (N_32960,N_32395,N_32308);
nand U32961 (N_32961,N_32455,N_32073);
nor U32962 (N_32962,N_32219,N_32417);
xnor U32963 (N_32963,N_32333,N_32244);
xor U32964 (N_32964,N_32215,N_32420);
xnor U32965 (N_32965,N_32439,N_32301);
nor U32966 (N_32966,N_32217,N_32027);
nor U32967 (N_32967,N_32298,N_32296);
nand U32968 (N_32968,N_32033,N_32142);
nor U32969 (N_32969,N_32494,N_32123);
xor U32970 (N_32970,N_32491,N_32095);
nor U32971 (N_32971,N_32333,N_32215);
nor U32972 (N_32972,N_32367,N_32425);
nand U32973 (N_32973,N_32296,N_32349);
nand U32974 (N_32974,N_32134,N_32187);
nand U32975 (N_32975,N_32058,N_32311);
nor U32976 (N_32976,N_32206,N_32241);
nor U32977 (N_32977,N_32394,N_32429);
nor U32978 (N_32978,N_32164,N_32332);
nand U32979 (N_32979,N_32228,N_32269);
and U32980 (N_32980,N_32182,N_32289);
nor U32981 (N_32981,N_32227,N_32442);
xnor U32982 (N_32982,N_32313,N_32038);
nand U32983 (N_32983,N_32472,N_32311);
nor U32984 (N_32984,N_32220,N_32358);
nor U32985 (N_32985,N_32436,N_32292);
and U32986 (N_32986,N_32008,N_32481);
or U32987 (N_32987,N_32065,N_32235);
nand U32988 (N_32988,N_32461,N_32278);
nor U32989 (N_32989,N_32224,N_32391);
nor U32990 (N_32990,N_32107,N_32354);
xnor U32991 (N_32991,N_32051,N_32059);
nand U32992 (N_32992,N_32473,N_32387);
or U32993 (N_32993,N_32179,N_32446);
and U32994 (N_32994,N_32489,N_32034);
or U32995 (N_32995,N_32046,N_32342);
and U32996 (N_32996,N_32315,N_32100);
and U32997 (N_32997,N_32436,N_32302);
xor U32998 (N_32998,N_32405,N_32003);
or U32999 (N_32999,N_32450,N_32387);
xor U33000 (N_33000,N_32892,N_32832);
nand U33001 (N_33001,N_32682,N_32840);
nor U33002 (N_33002,N_32640,N_32842);
nand U33003 (N_33003,N_32673,N_32802);
nand U33004 (N_33004,N_32618,N_32803);
or U33005 (N_33005,N_32786,N_32548);
nor U33006 (N_33006,N_32895,N_32849);
nor U33007 (N_33007,N_32817,N_32998);
nand U33008 (N_33008,N_32554,N_32760);
or U33009 (N_33009,N_32982,N_32617);
nand U33010 (N_33010,N_32980,N_32899);
and U33011 (N_33011,N_32599,N_32950);
xor U33012 (N_33012,N_32732,N_32806);
and U33013 (N_33013,N_32717,N_32583);
xor U33014 (N_33014,N_32693,N_32742);
and U33015 (N_33015,N_32775,N_32555);
and U33016 (N_33016,N_32983,N_32573);
and U33017 (N_33017,N_32666,N_32518);
nor U33018 (N_33018,N_32795,N_32956);
and U33019 (N_33019,N_32549,N_32722);
or U33020 (N_33020,N_32719,N_32924);
nand U33021 (N_33021,N_32745,N_32592);
or U33022 (N_33022,N_32532,N_32706);
xnor U33023 (N_33023,N_32999,N_32766);
xnor U33024 (N_33024,N_32578,N_32841);
nor U33025 (N_33025,N_32971,N_32597);
nor U33026 (N_33026,N_32923,N_32526);
or U33027 (N_33027,N_32981,N_32522);
xor U33028 (N_33028,N_32900,N_32784);
xnor U33029 (N_33029,N_32995,N_32858);
or U33030 (N_33030,N_32914,N_32725);
or U33031 (N_33031,N_32872,N_32600);
nor U33032 (N_33032,N_32631,N_32728);
or U33033 (N_33033,N_32677,N_32544);
and U33034 (N_33034,N_32959,N_32687);
or U33035 (N_33035,N_32553,N_32712);
or U33036 (N_33036,N_32848,N_32546);
nand U33037 (N_33037,N_32740,N_32884);
and U33038 (N_33038,N_32974,N_32845);
or U33039 (N_33039,N_32965,N_32877);
nand U33040 (N_33040,N_32861,N_32735);
nand U33041 (N_33041,N_32648,N_32608);
or U33042 (N_33042,N_32572,N_32696);
xor U33043 (N_33043,N_32812,N_32870);
or U33044 (N_33044,N_32559,N_32557);
and U33045 (N_33045,N_32616,N_32623);
and U33046 (N_33046,N_32713,N_32844);
nor U33047 (N_33047,N_32621,N_32756);
and U33048 (N_33048,N_32565,N_32826);
nand U33049 (N_33049,N_32500,N_32811);
or U33050 (N_33050,N_32566,N_32523);
or U33051 (N_33051,N_32933,N_32663);
nor U33052 (N_33052,N_32997,N_32765);
or U33053 (N_33053,N_32780,N_32881);
nand U33054 (N_33054,N_32837,N_32516);
nand U33055 (N_33055,N_32750,N_32678);
and U33056 (N_33056,N_32543,N_32751);
xor U33057 (N_33057,N_32643,N_32966);
or U33058 (N_33058,N_32787,N_32568);
and U33059 (N_33059,N_32519,N_32929);
and U33060 (N_33060,N_32530,N_32562);
xor U33061 (N_33061,N_32863,N_32791);
nor U33062 (N_33062,N_32650,N_32962);
or U33063 (N_33063,N_32893,N_32961);
nor U33064 (N_33064,N_32551,N_32550);
xnor U33065 (N_33065,N_32994,N_32828);
xnor U33066 (N_33066,N_32822,N_32627);
or U33067 (N_33067,N_32664,N_32767);
or U33068 (N_33068,N_32778,N_32903);
nor U33069 (N_33069,N_32556,N_32796);
nor U33070 (N_33070,N_32575,N_32936);
nor U33071 (N_33071,N_32584,N_32918);
nor U33072 (N_33072,N_32527,N_32847);
nand U33073 (N_33073,N_32540,N_32976);
nand U33074 (N_33074,N_32957,N_32537);
and U33075 (N_33075,N_32920,N_32862);
nor U33076 (N_33076,N_32602,N_32661);
nor U33077 (N_33077,N_32807,N_32793);
xnor U33078 (N_33078,N_32612,N_32658);
xor U33079 (N_33079,N_32913,N_32619);
nor U33080 (N_33080,N_32911,N_32823);
nor U33081 (N_33081,N_32505,N_32943);
xor U33082 (N_33082,N_32710,N_32590);
nand U33083 (N_33083,N_32581,N_32743);
and U33084 (N_33084,N_32649,N_32529);
xnor U33085 (N_33085,N_32659,N_32637);
xnor U33086 (N_33086,N_32703,N_32656);
nor U33087 (N_33087,N_32738,N_32757);
nor U33088 (N_33088,N_32639,N_32711);
and U33089 (N_33089,N_32718,N_32560);
xor U33090 (N_33090,N_32634,N_32701);
nand U33091 (N_33091,N_32674,N_32759);
or U33092 (N_33092,N_32800,N_32721);
nor U33093 (N_33093,N_32919,N_32978);
nand U33094 (N_33094,N_32908,N_32889);
or U33095 (N_33095,N_32808,N_32968);
nand U33096 (N_33096,N_32577,N_32541);
nand U33097 (N_33097,N_32867,N_32945);
nand U33098 (N_33098,N_32704,N_32922);
or U33099 (N_33099,N_32727,N_32730);
or U33100 (N_33100,N_32790,N_32694);
nand U33101 (N_33101,N_32988,N_32850);
or U33102 (N_33102,N_32932,N_32564);
nor U33103 (N_33103,N_32970,N_32912);
nand U33104 (N_33104,N_32853,N_32883);
or U33105 (N_33105,N_32771,N_32595);
nor U33106 (N_33106,N_32949,N_32671);
nand U33107 (N_33107,N_32657,N_32909);
or U33108 (N_33108,N_32879,N_32801);
xnor U33109 (N_33109,N_32715,N_32773);
nand U33110 (N_33110,N_32944,N_32508);
xor U33111 (N_33111,N_32758,N_32688);
or U33112 (N_33112,N_32977,N_32941);
nand U33113 (N_33113,N_32515,N_32752);
or U33114 (N_33114,N_32938,N_32503);
and U33115 (N_33115,N_32987,N_32927);
xor U33116 (N_33116,N_32521,N_32818);
or U33117 (N_33117,N_32604,N_32825);
xor U33118 (N_33118,N_32967,N_32935);
nor U33119 (N_33119,N_32514,N_32774);
and U33120 (N_33120,N_32902,N_32792);
or U33121 (N_33121,N_32753,N_32940);
nor U33122 (N_33122,N_32964,N_32937);
and U33123 (N_33123,N_32654,N_32824);
or U33124 (N_33124,N_32856,N_32882);
and U33125 (N_33125,N_32552,N_32542);
nand U33126 (N_33126,N_32810,N_32798);
nand U33127 (N_33127,N_32587,N_32630);
nor U33128 (N_33128,N_32680,N_32601);
and U33129 (N_33129,N_32887,N_32520);
nand U33130 (N_33130,N_32628,N_32558);
xnor U33131 (N_33131,N_32839,N_32580);
or U33132 (N_33132,N_32843,N_32814);
nand U33133 (N_33133,N_32763,N_32878);
or U33134 (N_33134,N_32746,N_32985);
or U33135 (N_33135,N_32984,N_32534);
or U33136 (N_33136,N_32739,N_32506);
or U33137 (N_33137,N_32734,N_32524);
xnor U33138 (N_33138,N_32813,N_32741);
nor U33139 (N_33139,N_32579,N_32692);
xor U33140 (N_33140,N_32797,N_32934);
nand U33141 (N_33141,N_32582,N_32799);
xor U33142 (N_33142,N_32836,N_32596);
or U33143 (N_33143,N_32691,N_32954);
nor U33144 (N_33144,N_32653,N_32942);
and U33145 (N_33145,N_32876,N_32831);
and U33146 (N_33146,N_32670,N_32794);
nor U33147 (N_33147,N_32921,N_32915);
or U33148 (N_33148,N_32570,N_32776);
xnor U33149 (N_33149,N_32615,N_32948);
and U33150 (N_33150,N_32834,N_32636);
nand U33151 (N_33151,N_32707,N_32905);
nor U33152 (N_33152,N_32667,N_32598);
xor U33153 (N_33153,N_32672,N_32951);
xor U33154 (N_33154,N_32747,N_32866);
or U33155 (N_33155,N_32737,N_32990);
xnor U33156 (N_33156,N_32655,N_32665);
and U33157 (N_33157,N_32854,N_32733);
nor U33158 (N_33158,N_32857,N_32609);
xnor U33159 (N_33159,N_32629,N_32567);
or U33160 (N_33160,N_32789,N_32859);
nand U33161 (N_33161,N_32864,N_32939);
and U33162 (N_33162,N_32535,N_32642);
nand U33163 (N_33163,N_32716,N_32533);
nand U33164 (N_33164,N_32662,N_32749);
or U33165 (N_33165,N_32809,N_32960);
or U33166 (N_33166,N_32729,N_32901);
xnor U33167 (N_33167,N_32897,N_32586);
nor U33168 (N_33168,N_32865,N_32569);
xor U33169 (N_33169,N_32958,N_32830);
xor U33170 (N_33170,N_32975,N_32547);
or U33171 (N_33171,N_32699,N_32916);
nor U33172 (N_33172,N_32947,N_32821);
or U33173 (N_33173,N_32504,N_32953);
and U33174 (N_33174,N_32772,N_32613);
nor U33175 (N_33175,N_32782,N_32955);
nand U33176 (N_33176,N_32846,N_32539);
or U33177 (N_33177,N_32926,N_32907);
and U33178 (N_33178,N_32898,N_32744);
xor U33179 (N_33179,N_32511,N_32925);
or U33180 (N_33180,N_32835,N_32531);
or U33181 (N_33181,N_32607,N_32788);
nand U33182 (N_33182,N_32886,N_32783);
or U33183 (N_33183,N_32963,N_32819);
xnor U33184 (N_33184,N_32668,N_32512);
and U33185 (N_33185,N_32875,N_32700);
nor U33186 (N_33186,N_32777,N_32633);
or U33187 (N_33187,N_32698,N_32689);
or U33188 (N_33188,N_32779,N_32708);
and U33189 (N_33189,N_32632,N_32611);
and U33190 (N_33190,N_32705,N_32762);
xnor U33191 (N_33191,N_32869,N_32761);
or U33192 (N_33192,N_32873,N_32904);
nand U33193 (N_33193,N_32588,N_32804);
nor U33194 (N_33194,N_32731,N_32880);
or U33195 (N_33195,N_32860,N_32635);
and U33196 (N_33196,N_32686,N_32805);
or U33197 (N_33197,N_32906,N_32685);
nor U33198 (N_33198,N_32679,N_32538);
and U33199 (N_33199,N_32785,N_32501);
and U33200 (N_33200,N_32645,N_32726);
or U33201 (N_33201,N_32972,N_32571);
nand U33202 (N_33202,N_32561,N_32973);
nand U33203 (N_33203,N_32928,N_32626);
nor U33204 (N_33204,N_32991,N_32755);
nor U33205 (N_33205,N_32697,N_32610);
nand U33206 (N_33206,N_32768,N_32720);
or U33207 (N_33207,N_32614,N_32838);
nand U33208 (N_33208,N_32986,N_32690);
nor U33209 (N_33209,N_32695,N_32754);
nor U33210 (N_33210,N_32675,N_32576);
xnor U33211 (N_33211,N_32917,N_32885);
xor U33212 (N_33212,N_32651,N_32709);
xnor U33213 (N_33213,N_32946,N_32574);
xor U33214 (N_33214,N_32868,N_32585);
xor U33215 (N_33215,N_32931,N_32815);
and U33216 (N_33216,N_32769,N_32647);
nand U33217 (N_33217,N_32684,N_32993);
and U33218 (N_33218,N_32545,N_32669);
or U33219 (N_33219,N_32652,N_32992);
nand U33220 (N_33220,N_32827,N_32681);
nor U33221 (N_33221,N_32891,N_32930);
or U33222 (N_33222,N_32702,N_32641);
or U33223 (N_33223,N_32723,N_32676);
and U33224 (N_33224,N_32563,N_32952);
xor U33225 (N_33225,N_32528,N_32624);
or U33226 (N_33226,N_32593,N_32605);
nand U33227 (N_33227,N_32510,N_32736);
and U33228 (N_33228,N_32829,N_32502);
nor U33229 (N_33229,N_32969,N_32591);
and U33230 (N_33230,N_32646,N_32622);
xnor U33231 (N_33231,N_32509,N_32606);
and U33232 (N_33232,N_32890,N_32781);
nor U33233 (N_33233,N_32820,N_32851);
xor U33234 (N_33234,N_32638,N_32888);
and U33235 (N_33235,N_32620,N_32770);
xor U33236 (N_33236,N_32748,N_32644);
xnor U33237 (N_33237,N_32894,N_32816);
nand U33238 (N_33238,N_32896,N_32536);
and U33239 (N_33239,N_32683,N_32855);
nor U33240 (N_33240,N_32625,N_32594);
nand U33241 (N_33241,N_32979,N_32513);
nor U33242 (N_33242,N_32589,N_32603);
or U33243 (N_33243,N_32764,N_32989);
xor U33244 (N_33244,N_32833,N_32724);
nor U33245 (N_33245,N_32507,N_32517);
nor U33246 (N_33246,N_32996,N_32852);
and U33247 (N_33247,N_32910,N_32874);
nor U33248 (N_33248,N_32525,N_32660);
nor U33249 (N_33249,N_32871,N_32714);
and U33250 (N_33250,N_32502,N_32927);
nand U33251 (N_33251,N_32848,N_32894);
nand U33252 (N_33252,N_32677,N_32524);
nand U33253 (N_33253,N_32883,N_32929);
and U33254 (N_33254,N_32610,N_32877);
nand U33255 (N_33255,N_32836,N_32781);
nand U33256 (N_33256,N_32911,N_32897);
nor U33257 (N_33257,N_32869,N_32807);
and U33258 (N_33258,N_32573,N_32913);
nand U33259 (N_33259,N_32617,N_32779);
xor U33260 (N_33260,N_32671,N_32524);
and U33261 (N_33261,N_32555,N_32741);
nor U33262 (N_33262,N_32856,N_32539);
and U33263 (N_33263,N_32896,N_32995);
nor U33264 (N_33264,N_32627,N_32998);
nor U33265 (N_33265,N_32854,N_32844);
and U33266 (N_33266,N_32520,N_32898);
nor U33267 (N_33267,N_32811,N_32914);
nor U33268 (N_33268,N_32556,N_32648);
xnor U33269 (N_33269,N_32545,N_32889);
xor U33270 (N_33270,N_32561,N_32548);
nand U33271 (N_33271,N_32654,N_32679);
nor U33272 (N_33272,N_32900,N_32760);
xor U33273 (N_33273,N_32887,N_32923);
and U33274 (N_33274,N_32726,N_32994);
nor U33275 (N_33275,N_32605,N_32525);
xor U33276 (N_33276,N_32671,N_32916);
xnor U33277 (N_33277,N_32685,N_32693);
and U33278 (N_33278,N_32743,N_32611);
xor U33279 (N_33279,N_32620,N_32514);
xor U33280 (N_33280,N_32615,N_32514);
or U33281 (N_33281,N_32808,N_32614);
xor U33282 (N_33282,N_32635,N_32764);
and U33283 (N_33283,N_32929,N_32596);
nand U33284 (N_33284,N_32846,N_32551);
nand U33285 (N_33285,N_32688,N_32510);
nand U33286 (N_33286,N_32778,N_32883);
nor U33287 (N_33287,N_32739,N_32757);
xnor U33288 (N_33288,N_32906,N_32534);
xnor U33289 (N_33289,N_32734,N_32891);
and U33290 (N_33290,N_32923,N_32616);
xor U33291 (N_33291,N_32605,N_32514);
nand U33292 (N_33292,N_32829,N_32694);
and U33293 (N_33293,N_32770,N_32680);
xnor U33294 (N_33294,N_32953,N_32815);
nor U33295 (N_33295,N_32672,N_32696);
nand U33296 (N_33296,N_32629,N_32810);
or U33297 (N_33297,N_32706,N_32724);
or U33298 (N_33298,N_32723,N_32712);
nor U33299 (N_33299,N_32888,N_32989);
nand U33300 (N_33300,N_32735,N_32543);
nand U33301 (N_33301,N_32954,N_32929);
nor U33302 (N_33302,N_32665,N_32956);
nand U33303 (N_33303,N_32994,N_32959);
or U33304 (N_33304,N_32867,N_32524);
nand U33305 (N_33305,N_32868,N_32820);
nor U33306 (N_33306,N_32994,N_32534);
nor U33307 (N_33307,N_32976,N_32707);
and U33308 (N_33308,N_32984,N_32935);
or U33309 (N_33309,N_32738,N_32904);
xor U33310 (N_33310,N_32887,N_32991);
and U33311 (N_33311,N_32963,N_32589);
nand U33312 (N_33312,N_32728,N_32759);
nand U33313 (N_33313,N_32778,N_32751);
nor U33314 (N_33314,N_32601,N_32820);
and U33315 (N_33315,N_32624,N_32845);
nand U33316 (N_33316,N_32934,N_32945);
or U33317 (N_33317,N_32924,N_32665);
nand U33318 (N_33318,N_32822,N_32971);
and U33319 (N_33319,N_32693,N_32629);
and U33320 (N_33320,N_32567,N_32753);
nor U33321 (N_33321,N_32571,N_32874);
xnor U33322 (N_33322,N_32593,N_32528);
nor U33323 (N_33323,N_32568,N_32663);
or U33324 (N_33324,N_32717,N_32520);
nor U33325 (N_33325,N_32683,N_32719);
xnor U33326 (N_33326,N_32929,N_32712);
nand U33327 (N_33327,N_32727,N_32690);
nand U33328 (N_33328,N_32655,N_32892);
nand U33329 (N_33329,N_32533,N_32916);
and U33330 (N_33330,N_32637,N_32707);
or U33331 (N_33331,N_32528,N_32661);
nand U33332 (N_33332,N_32967,N_32963);
nand U33333 (N_33333,N_32922,N_32636);
or U33334 (N_33334,N_32855,N_32650);
nand U33335 (N_33335,N_32882,N_32806);
nor U33336 (N_33336,N_32823,N_32509);
and U33337 (N_33337,N_32992,N_32941);
or U33338 (N_33338,N_32968,N_32565);
and U33339 (N_33339,N_32819,N_32641);
nor U33340 (N_33340,N_32767,N_32876);
xnor U33341 (N_33341,N_32793,N_32906);
nor U33342 (N_33342,N_32711,N_32976);
nor U33343 (N_33343,N_32557,N_32927);
nand U33344 (N_33344,N_32901,N_32876);
and U33345 (N_33345,N_32537,N_32588);
nor U33346 (N_33346,N_32520,N_32952);
xnor U33347 (N_33347,N_32954,N_32937);
nor U33348 (N_33348,N_32725,N_32763);
nor U33349 (N_33349,N_32630,N_32759);
xor U33350 (N_33350,N_32783,N_32770);
and U33351 (N_33351,N_32740,N_32918);
and U33352 (N_33352,N_32885,N_32857);
or U33353 (N_33353,N_32507,N_32515);
xor U33354 (N_33354,N_32660,N_32900);
and U33355 (N_33355,N_32809,N_32824);
xnor U33356 (N_33356,N_32560,N_32536);
or U33357 (N_33357,N_32921,N_32594);
nand U33358 (N_33358,N_32530,N_32832);
nand U33359 (N_33359,N_32522,N_32898);
nor U33360 (N_33360,N_32690,N_32719);
and U33361 (N_33361,N_32501,N_32986);
nor U33362 (N_33362,N_32822,N_32697);
and U33363 (N_33363,N_32986,N_32879);
or U33364 (N_33364,N_32967,N_32853);
or U33365 (N_33365,N_32755,N_32848);
or U33366 (N_33366,N_32887,N_32535);
or U33367 (N_33367,N_32756,N_32980);
nand U33368 (N_33368,N_32814,N_32905);
nand U33369 (N_33369,N_32571,N_32534);
or U33370 (N_33370,N_32639,N_32935);
or U33371 (N_33371,N_32626,N_32827);
or U33372 (N_33372,N_32869,N_32719);
nor U33373 (N_33373,N_32801,N_32528);
xnor U33374 (N_33374,N_32812,N_32627);
nand U33375 (N_33375,N_32617,N_32803);
xnor U33376 (N_33376,N_32919,N_32666);
and U33377 (N_33377,N_32730,N_32874);
or U33378 (N_33378,N_32828,N_32850);
nand U33379 (N_33379,N_32572,N_32655);
or U33380 (N_33380,N_32684,N_32948);
or U33381 (N_33381,N_32672,N_32875);
and U33382 (N_33382,N_32566,N_32834);
and U33383 (N_33383,N_32638,N_32651);
nor U33384 (N_33384,N_32872,N_32726);
or U33385 (N_33385,N_32528,N_32527);
or U33386 (N_33386,N_32805,N_32999);
nand U33387 (N_33387,N_32517,N_32751);
nor U33388 (N_33388,N_32824,N_32669);
or U33389 (N_33389,N_32652,N_32542);
and U33390 (N_33390,N_32514,N_32937);
nor U33391 (N_33391,N_32559,N_32969);
xnor U33392 (N_33392,N_32865,N_32869);
and U33393 (N_33393,N_32674,N_32999);
nand U33394 (N_33394,N_32820,N_32918);
nor U33395 (N_33395,N_32789,N_32973);
and U33396 (N_33396,N_32573,N_32673);
xor U33397 (N_33397,N_32779,N_32717);
or U33398 (N_33398,N_32920,N_32907);
and U33399 (N_33399,N_32582,N_32796);
nand U33400 (N_33400,N_32561,N_32919);
or U33401 (N_33401,N_32910,N_32892);
nand U33402 (N_33402,N_32765,N_32744);
nand U33403 (N_33403,N_32852,N_32686);
and U33404 (N_33404,N_32999,N_32692);
and U33405 (N_33405,N_32621,N_32976);
and U33406 (N_33406,N_32640,N_32805);
xor U33407 (N_33407,N_32731,N_32521);
or U33408 (N_33408,N_32908,N_32922);
and U33409 (N_33409,N_32593,N_32999);
nor U33410 (N_33410,N_32668,N_32504);
xnor U33411 (N_33411,N_32604,N_32893);
and U33412 (N_33412,N_32905,N_32588);
and U33413 (N_33413,N_32532,N_32674);
and U33414 (N_33414,N_32919,N_32560);
nor U33415 (N_33415,N_32645,N_32586);
xor U33416 (N_33416,N_32882,N_32513);
nor U33417 (N_33417,N_32908,N_32507);
nand U33418 (N_33418,N_32760,N_32807);
xnor U33419 (N_33419,N_32838,N_32640);
or U33420 (N_33420,N_32830,N_32704);
and U33421 (N_33421,N_32850,N_32779);
nand U33422 (N_33422,N_32868,N_32809);
nand U33423 (N_33423,N_32528,N_32883);
nor U33424 (N_33424,N_32930,N_32526);
xnor U33425 (N_33425,N_32694,N_32624);
nand U33426 (N_33426,N_32813,N_32887);
xnor U33427 (N_33427,N_32961,N_32769);
or U33428 (N_33428,N_32908,N_32814);
and U33429 (N_33429,N_32574,N_32643);
or U33430 (N_33430,N_32940,N_32691);
xor U33431 (N_33431,N_32542,N_32718);
and U33432 (N_33432,N_32890,N_32674);
and U33433 (N_33433,N_32582,N_32631);
xnor U33434 (N_33434,N_32606,N_32967);
xor U33435 (N_33435,N_32973,N_32791);
nor U33436 (N_33436,N_32973,N_32880);
and U33437 (N_33437,N_32903,N_32817);
nand U33438 (N_33438,N_32654,N_32721);
xnor U33439 (N_33439,N_32744,N_32858);
or U33440 (N_33440,N_32647,N_32791);
nand U33441 (N_33441,N_32729,N_32700);
and U33442 (N_33442,N_32637,N_32700);
and U33443 (N_33443,N_32775,N_32770);
xor U33444 (N_33444,N_32972,N_32582);
xor U33445 (N_33445,N_32603,N_32626);
nor U33446 (N_33446,N_32925,N_32941);
xor U33447 (N_33447,N_32917,N_32596);
nand U33448 (N_33448,N_32584,N_32653);
xnor U33449 (N_33449,N_32701,N_32941);
xor U33450 (N_33450,N_32712,N_32576);
or U33451 (N_33451,N_32774,N_32944);
nand U33452 (N_33452,N_32630,N_32593);
nand U33453 (N_33453,N_32508,N_32664);
nor U33454 (N_33454,N_32519,N_32526);
and U33455 (N_33455,N_32639,N_32681);
nor U33456 (N_33456,N_32556,N_32941);
and U33457 (N_33457,N_32703,N_32925);
nand U33458 (N_33458,N_32700,N_32530);
nor U33459 (N_33459,N_32922,N_32750);
and U33460 (N_33460,N_32646,N_32986);
nand U33461 (N_33461,N_32631,N_32514);
or U33462 (N_33462,N_32995,N_32838);
or U33463 (N_33463,N_32671,N_32924);
nand U33464 (N_33464,N_32998,N_32656);
xor U33465 (N_33465,N_32563,N_32844);
or U33466 (N_33466,N_32882,N_32916);
nor U33467 (N_33467,N_32836,N_32959);
or U33468 (N_33468,N_32872,N_32771);
xnor U33469 (N_33469,N_32848,N_32771);
nand U33470 (N_33470,N_32983,N_32963);
nand U33471 (N_33471,N_32892,N_32845);
and U33472 (N_33472,N_32529,N_32806);
nand U33473 (N_33473,N_32905,N_32653);
or U33474 (N_33474,N_32563,N_32505);
nand U33475 (N_33475,N_32826,N_32628);
nor U33476 (N_33476,N_32630,N_32949);
or U33477 (N_33477,N_32674,N_32849);
or U33478 (N_33478,N_32515,N_32630);
and U33479 (N_33479,N_32681,N_32948);
or U33480 (N_33480,N_32976,N_32949);
nand U33481 (N_33481,N_32845,N_32781);
or U33482 (N_33482,N_32890,N_32887);
nor U33483 (N_33483,N_32796,N_32789);
or U33484 (N_33484,N_32882,N_32671);
or U33485 (N_33485,N_32567,N_32785);
nand U33486 (N_33486,N_32543,N_32608);
or U33487 (N_33487,N_32649,N_32750);
xnor U33488 (N_33488,N_32872,N_32983);
nor U33489 (N_33489,N_32699,N_32757);
and U33490 (N_33490,N_32556,N_32777);
or U33491 (N_33491,N_32952,N_32549);
xor U33492 (N_33492,N_32853,N_32706);
nand U33493 (N_33493,N_32849,N_32850);
xor U33494 (N_33494,N_32717,N_32749);
nor U33495 (N_33495,N_32971,N_32568);
or U33496 (N_33496,N_32865,N_32757);
nand U33497 (N_33497,N_32640,N_32962);
and U33498 (N_33498,N_32949,N_32607);
or U33499 (N_33499,N_32797,N_32659);
or U33500 (N_33500,N_33184,N_33159);
and U33501 (N_33501,N_33222,N_33356);
or U33502 (N_33502,N_33358,N_33274);
xor U33503 (N_33503,N_33178,N_33145);
and U33504 (N_33504,N_33200,N_33426);
xor U33505 (N_33505,N_33047,N_33316);
nand U33506 (N_33506,N_33215,N_33369);
or U33507 (N_33507,N_33080,N_33134);
or U33508 (N_33508,N_33071,N_33329);
nand U33509 (N_33509,N_33064,N_33227);
xor U33510 (N_33510,N_33138,N_33477);
or U33511 (N_33511,N_33401,N_33482);
and U33512 (N_33512,N_33385,N_33088);
nand U33513 (N_33513,N_33390,N_33366);
and U33514 (N_33514,N_33220,N_33190);
nand U33515 (N_33515,N_33201,N_33150);
xor U33516 (N_33516,N_33235,N_33449);
or U33517 (N_33517,N_33028,N_33219);
xor U33518 (N_33518,N_33381,N_33348);
or U33519 (N_33519,N_33133,N_33281);
nand U33520 (N_33520,N_33406,N_33428);
xnor U33521 (N_33521,N_33483,N_33130);
nand U33522 (N_33522,N_33164,N_33214);
nand U33523 (N_33523,N_33257,N_33173);
xor U33524 (N_33524,N_33113,N_33213);
nor U33525 (N_33525,N_33212,N_33490);
and U33526 (N_33526,N_33299,N_33306);
or U33527 (N_33527,N_33098,N_33497);
xnor U33528 (N_33528,N_33325,N_33059);
xor U33529 (N_33529,N_33140,N_33077);
and U33530 (N_33530,N_33045,N_33174);
xnor U33531 (N_33531,N_33270,N_33106);
nor U33532 (N_33532,N_33127,N_33421);
and U33533 (N_33533,N_33397,N_33155);
and U33534 (N_33534,N_33262,N_33414);
or U33535 (N_33535,N_33206,N_33353);
or U33536 (N_33536,N_33313,N_33240);
xor U33537 (N_33537,N_33117,N_33493);
or U33538 (N_33538,N_33055,N_33415);
nor U33539 (N_33539,N_33470,N_33333);
nor U33540 (N_33540,N_33437,N_33374);
or U33541 (N_33541,N_33139,N_33052);
nand U33542 (N_33542,N_33392,N_33443);
nand U33543 (N_33543,N_33442,N_33268);
or U33544 (N_33544,N_33244,N_33456);
xor U33545 (N_33545,N_33198,N_33065);
or U33546 (N_33546,N_33332,N_33312);
nor U33547 (N_33547,N_33157,N_33195);
and U33548 (N_33548,N_33249,N_33231);
and U33549 (N_33549,N_33375,N_33423);
nand U33550 (N_33550,N_33013,N_33296);
xor U33551 (N_33551,N_33376,N_33239);
nor U33552 (N_33552,N_33101,N_33492);
nor U33553 (N_33553,N_33438,N_33398);
and U33554 (N_33554,N_33409,N_33391);
or U33555 (N_33555,N_33417,N_33499);
and U33556 (N_33556,N_33057,N_33435);
xor U33557 (N_33557,N_33429,N_33453);
xnor U33558 (N_33558,N_33335,N_33310);
nor U33559 (N_33559,N_33458,N_33441);
and U33560 (N_33560,N_33091,N_33290);
and U33561 (N_33561,N_33051,N_33054);
nand U33562 (N_33562,N_33021,N_33166);
nand U33563 (N_33563,N_33293,N_33412);
and U33564 (N_33564,N_33181,N_33177);
nand U33565 (N_33565,N_33085,N_33189);
or U33566 (N_33566,N_33160,N_33108);
or U33567 (N_33567,N_33009,N_33183);
nor U33568 (N_33568,N_33046,N_33163);
xor U33569 (N_33569,N_33121,N_33258);
and U33570 (N_33570,N_33185,N_33143);
and U33571 (N_33571,N_33033,N_33191);
and U33572 (N_33572,N_33387,N_33093);
nor U33573 (N_33573,N_33169,N_33202);
xnor U33574 (N_33574,N_33430,N_33072);
nand U33575 (N_33575,N_33444,N_33000);
xnor U33576 (N_33576,N_33498,N_33095);
nand U33577 (N_33577,N_33084,N_33207);
xor U33578 (N_33578,N_33250,N_33115);
nand U33579 (N_33579,N_33125,N_33287);
or U33580 (N_33580,N_33131,N_33355);
xor U33581 (N_33581,N_33092,N_33342);
or U33582 (N_33582,N_33460,N_33188);
xnor U33583 (N_33583,N_33481,N_33246);
nor U33584 (N_33584,N_33330,N_33367);
nand U33585 (N_33585,N_33102,N_33336);
xor U33586 (N_33586,N_33010,N_33225);
nand U33587 (N_33587,N_33221,N_33344);
xor U33588 (N_33588,N_33408,N_33253);
xnor U33589 (N_33589,N_33479,N_33199);
xnor U33590 (N_33590,N_33286,N_33090);
xnor U33591 (N_33591,N_33022,N_33340);
nor U33592 (N_33592,N_33323,N_33269);
or U33593 (N_33593,N_33229,N_33067);
nand U33594 (N_33594,N_33129,N_33454);
xnor U33595 (N_33595,N_33056,N_33451);
nor U33596 (N_33596,N_33204,N_33350);
nor U33597 (N_33597,N_33315,N_33082);
and U33598 (N_33598,N_33378,N_33370);
and U33599 (N_33599,N_33211,N_33402);
nand U33600 (N_33600,N_33005,N_33165);
or U33601 (N_33601,N_33053,N_33389);
xor U33602 (N_33602,N_33124,N_33265);
nor U33603 (N_33603,N_33151,N_33100);
and U33604 (N_33604,N_33069,N_33485);
nand U33605 (N_33605,N_33447,N_33413);
xor U33606 (N_33606,N_33463,N_33388);
nand U33607 (N_33607,N_33464,N_33144);
xnor U33608 (N_33608,N_33345,N_33099);
nor U33609 (N_33609,N_33475,N_33436);
xnor U33610 (N_33610,N_33217,N_33301);
nor U33611 (N_33611,N_33284,N_33334);
nand U33612 (N_33612,N_33180,N_33007);
nor U33613 (N_33613,N_33360,N_33282);
nand U33614 (N_33614,N_33081,N_33132);
and U33615 (N_33615,N_33109,N_33309);
xnor U33616 (N_33616,N_33386,N_33276);
and U33617 (N_33617,N_33491,N_33318);
nor U33618 (N_33618,N_33289,N_33023);
or U33619 (N_33619,N_33128,N_33404);
or U33620 (N_33620,N_33186,N_33273);
nand U33621 (N_33621,N_33321,N_33450);
and U33622 (N_33622,N_33058,N_33017);
nand U33623 (N_33623,N_33030,N_33107);
xnor U33624 (N_33624,N_33152,N_33403);
nand U33625 (N_33625,N_33368,N_33148);
nand U33626 (N_33626,N_33048,N_33176);
xor U33627 (N_33627,N_33272,N_33226);
nor U33628 (N_33628,N_33288,N_33362);
nor U33629 (N_33629,N_33416,N_33419);
nor U33630 (N_33630,N_33234,N_33489);
and U33631 (N_33631,N_33086,N_33295);
or U33632 (N_33632,N_33083,N_33149);
xor U33633 (N_33633,N_33480,N_33486);
nand U33634 (N_33634,N_33062,N_33359);
xnor U33635 (N_33635,N_33252,N_33020);
nor U33636 (N_33636,N_33034,N_33372);
nand U33637 (N_33637,N_33110,N_33126);
and U33638 (N_33638,N_33431,N_33024);
nor U33639 (N_33639,N_33474,N_33352);
nor U33640 (N_33640,N_33147,N_33001);
nand U33641 (N_33641,N_33433,N_33019);
or U33642 (N_33642,N_33411,N_33255);
nand U33643 (N_33643,N_33462,N_33380);
nand U33644 (N_33644,N_33425,N_33236);
nand U33645 (N_33645,N_33223,N_33461);
xnor U33646 (N_33646,N_33043,N_33271);
xnor U33647 (N_33647,N_33011,N_33298);
and U33648 (N_33648,N_33297,N_33337);
nand U33649 (N_33649,N_33384,N_33264);
and U33650 (N_33650,N_33070,N_33142);
or U33651 (N_33651,N_33488,N_33029);
nor U33652 (N_33652,N_33209,N_33478);
or U33653 (N_33653,N_33407,N_33434);
xor U33654 (N_33654,N_33104,N_33156);
nand U33655 (N_33655,N_33187,N_33146);
nor U33656 (N_33656,N_33118,N_33153);
nand U33657 (N_33657,N_33373,N_33076);
or U33658 (N_33658,N_33006,N_33197);
xnor U33659 (N_33659,N_33158,N_33439);
and U33660 (N_33660,N_33120,N_33260);
nor U33661 (N_33661,N_33014,N_33161);
xnor U33662 (N_33662,N_33060,N_33050);
or U33663 (N_33663,N_33467,N_33291);
or U33664 (N_33664,N_33228,N_33324);
nor U33665 (N_33665,N_33018,N_33027);
nor U33666 (N_33666,N_33196,N_33237);
nor U33667 (N_33667,N_33472,N_33208);
nor U33668 (N_33668,N_33418,N_33171);
and U33669 (N_33669,N_33233,N_33025);
or U33670 (N_33670,N_33016,N_33194);
and U33671 (N_33671,N_33266,N_33357);
or U33672 (N_33672,N_33468,N_33382);
nor U33673 (N_33673,N_33445,N_33292);
xor U33674 (N_33674,N_33494,N_33136);
xor U33675 (N_33675,N_33305,N_33457);
and U33676 (N_33676,N_33326,N_33410);
xnor U33677 (N_33677,N_33210,N_33243);
and U33678 (N_33678,N_33218,N_33496);
and U33679 (N_33679,N_33031,N_33167);
nor U33680 (N_33680,N_33135,N_33327);
and U33681 (N_33681,N_33203,N_33394);
and U33682 (N_33682,N_33087,N_33331);
nor U33683 (N_33683,N_33094,N_33123);
xor U33684 (N_33684,N_33141,N_33427);
nand U33685 (N_33685,N_33383,N_33036);
nor U33686 (N_33686,N_33004,N_33300);
and U33687 (N_33687,N_33012,N_33363);
and U33688 (N_33688,N_33349,N_33371);
xnor U33689 (N_33689,N_33044,N_33103);
and U33690 (N_33690,N_33365,N_33277);
or U33691 (N_33691,N_33230,N_33170);
xnor U33692 (N_33692,N_33302,N_33259);
or U33693 (N_33693,N_33294,N_33396);
xnor U33694 (N_33694,N_33038,N_33002);
nand U33695 (N_33695,N_33039,N_33471);
nand U33696 (N_33696,N_33354,N_33049);
or U33697 (N_33697,N_33341,N_33484);
xor U33698 (N_33698,N_33193,N_33192);
xnor U33699 (N_33699,N_33320,N_33303);
nor U33700 (N_33700,N_33008,N_33168);
xnor U33701 (N_33701,N_33105,N_33377);
and U33702 (N_33702,N_33432,N_33304);
and U33703 (N_33703,N_33278,N_33420);
or U33704 (N_33704,N_33275,N_33232);
nor U33705 (N_33705,N_33179,N_33073);
nand U33706 (N_33706,N_33238,N_33311);
nand U33707 (N_33707,N_33122,N_33465);
and U33708 (N_33708,N_33096,N_33267);
nor U33709 (N_33709,N_33263,N_33162);
or U33710 (N_33710,N_33172,N_33400);
or U33711 (N_33711,N_33495,N_33308);
nand U33712 (N_33712,N_33361,N_33487);
or U33713 (N_33713,N_33319,N_33364);
or U33714 (N_33714,N_33254,N_33338);
and U33715 (N_33715,N_33446,N_33205);
and U33716 (N_33716,N_33041,N_33283);
or U33717 (N_33717,N_33015,N_33455);
nor U33718 (N_33718,N_33003,N_33347);
or U33719 (N_33719,N_33251,N_33343);
xnor U33720 (N_33720,N_33307,N_33035);
nand U33721 (N_33721,N_33111,N_33061);
nand U33722 (N_33722,N_33063,N_33248);
and U33723 (N_33723,N_33346,N_33241);
xnor U33724 (N_33724,N_33452,N_33245);
nor U33725 (N_33725,N_33317,N_33175);
or U33726 (N_33726,N_33075,N_33393);
xor U33727 (N_33727,N_33328,N_33112);
xnor U33728 (N_33728,N_33119,N_33440);
xor U33729 (N_33729,N_33339,N_33032);
xnor U33730 (N_33730,N_33097,N_33256);
nand U33731 (N_33731,N_33182,N_33247);
or U33732 (N_33732,N_33279,N_33079);
nor U33733 (N_33733,N_33216,N_33405);
and U33734 (N_33734,N_33114,N_33379);
nand U33735 (N_33735,N_33314,N_33285);
and U33736 (N_33736,N_33224,N_33422);
and U33737 (N_33737,N_33042,N_33322);
xnor U33738 (N_33738,N_33399,N_33395);
xnor U33739 (N_33739,N_33280,N_33066);
and U33740 (N_33740,N_33469,N_33078);
and U33741 (N_33741,N_33242,N_33068);
xnor U33742 (N_33742,N_33466,N_33137);
or U33743 (N_33743,N_33089,N_33154);
nand U33744 (N_33744,N_33351,N_33424);
nand U33745 (N_33745,N_33116,N_33476);
or U33746 (N_33746,N_33448,N_33037);
and U33747 (N_33747,N_33074,N_33261);
nor U33748 (N_33748,N_33459,N_33040);
nand U33749 (N_33749,N_33026,N_33473);
nor U33750 (N_33750,N_33238,N_33392);
and U33751 (N_33751,N_33195,N_33142);
nand U33752 (N_33752,N_33125,N_33075);
and U33753 (N_33753,N_33201,N_33450);
and U33754 (N_33754,N_33336,N_33134);
nand U33755 (N_33755,N_33374,N_33414);
nand U33756 (N_33756,N_33297,N_33209);
nand U33757 (N_33757,N_33340,N_33269);
xnor U33758 (N_33758,N_33010,N_33177);
or U33759 (N_33759,N_33389,N_33446);
and U33760 (N_33760,N_33128,N_33113);
nor U33761 (N_33761,N_33073,N_33208);
or U33762 (N_33762,N_33002,N_33048);
and U33763 (N_33763,N_33083,N_33261);
nand U33764 (N_33764,N_33140,N_33306);
xor U33765 (N_33765,N_33441,N_33220);
nor U33766 (N_33766,N_33002,N_33387);
nand U33767 (N_33767,N_33420,N_33457);
nand U33768 (N_33768,N_33293,N_33057);
nand U33769 (N_33769,N_33378,N_33424);
xor U33770 (N_33770,N_33285,N_33131);
and U33771 (N_33771,N_33405,N_33076);
and U33772 (N_33772,N_33048,N_33434);
xor U33773 (N_33773,N_33401,N_33402);
nor U33774 (N_33774,N_33216,N_33053);
nand U33775 (N_33775,N_33458,N_33327);
nor U33776 (N_33776,N_33206,N_33131);
xnor U33777 (N_33777,N_33187,N_33284);
or U33778 (N_33778,N_33131,N_33395);
xor U33779 (N_33779,N_33057,N_33266);
nand U33780 (N_33780,N_33000,N_33275);
nor U33781 (N_33781,N_33011,N_33472);
xor U33782 (N_33782,N_33323,N_33081);
nand U33783 (N_33783,N_33166,N_33223);
or U33784 (N_33784,N_33135,N_33339);
nand U33785 (N_33785,N_33159,N_33456);
nand U33786 (N_33786,N_33426,N_33459);
xor U33787 (N_33787,N_33290,N_33487);
nor U33788 (N_33788,N_33144,N_33217);
or U33789 (N_33789,N_33241,N_33442);
nand U33790 (N_33790,N_33400,N_33226);
xor U33791 (N_33791,N_33371,N_33352);
nor U33792 (N_33792,N_33276,N_33292);
and U33793 (N_33793,N_33420,N_33479);
xnor U33794 (N_33794,N_33136,N_33112);
or U33795 (N_33795,N_33115,N_33220);
xor U33796 (N_33796,N_33248,N_33262);
nand U33797 (N_33797,N_33089,N_33121);
xor U33798 (N_33798,N_33220,N_33439);
nand U33799 (N_33799,N_33271,N_33451);
and U33800 (N_33800,N_33453,N_33483);
nor U33801 (N_33801,N_33408,N_33203);
or U33802 (N_33802,N_33029,N_33188);
or U33803 (N_33803,N_33476,N_33403);
and U33804 (N_33804,N_33358,N_33114);
nor U33805 (N_33805,N_33175,N_33066);
xnor U33806 (N_33806,N_33246,N_33139);
nand U33807 (N_33807,N_33451,N_33419);
nand U33808 (N_33808,N_33442,N_33065);
and U33809 (N_33809,N_33195,N_33349);
and U33810 (N_33810,N_33258,N_33140);
and U33811 (N_33811,N_33323,N_33019);
nand U33812 (N_33812,N_33399,N_33264);
and U33813 (N_33813,N_33433,N_33194);
or U33814 (N_33814,N_33118,N_33239);
or U33815 (N_33815,N_33275,N_33359);
or U33816 (N_33816,N_33073,N_33352);
nor U33817 (N_33817,N_33006,N_33120);
or U33818 (N_33818,N_33483,N_33187);
nor U33819 (N_33819,N_33001,N_33454);
xnor U33820 (N_33820,N_33474,N_33388);
nand U33821 (N_33821,N_33097,N_33327);
nor U33822 (N_33822,N_33298,N_33176);
and U33823 (N_33823,N_33256,N_33029);
or U33824 (N_33824,N_33435,N_33280);
nand U33825 (N_33825,N_33396,N_33076);
nand U33826 (N_33826,N_33003,N_33182);
nor U33827 (N_33827,N_33087,N_33074);
nor U33828 (N_33828,N_33094,N_33469);
nand U33829 (N_33829,N_33211,N_33356);
and U33830 (N_33830,N_33485,N_33399);
nand U33831 (N_33831,N_33126,N_33331);
or U33832 (N_33832,N_33442,N_33056);
nand U33833 (N_33833,N_33415,N_33381);
and U33834 (N_33834,N_33478,N_33219);
nor U33835 (N_33835,N_33273,N_33476);
and U33836 (N_33836,N_33366,N_33228);
or U33837 (N_33837,N_33121,N_33331);
and U33838 (N_33838,N_33179,N_33204);
nand U33839 (N_33839,N_33372,N_33486);
and U33840 (N_33840,N_33019,N_33143);
nand U33841 (N_33841,N_33021,N_33465);
xnor U33842 (N_33842,N_33480,N_33490);
and U33843 (N_33843,N_33405,N_33416);
xnor U33844 (N_33844,N_33093,N_33497);
or U33845 (N_33845,N_33105,N_33080);
nand U33846 (N_33846,N_33260,N_33116);
and U33847 (N_33847,N_33306,N_33378);
and U33848 (N_33848,N_33427,N_33274);
nand U33849 (N_33849,N_33193,N_33362);
nor U33850 (N_33850,N_33074,N_33439);
and U33851 (N_33851,N_33158,N_33404);
nor U33852 (N_33852,N_33401,N_33478);
and U33853 (N_33853,N_33471,N_33332);
or U33854 (N_33854,N_33379,N_33421);
xnor U33855 (N_33855,N_33141,N_33065);
xor U33856 (N_33856,N_33215,N_33249);
and U33857 (N_33857,N_33160,N_33074);
nor U33858 (N_33858,N_33285,N_33250);
xnor U33859 (N_33859,N_33089,N_33228);
nand U33860 (N_33860,N_33497,N_33249);
nor U33861 (N_33861,N_33174,N_33466);
nor U33862 (N_33862,N_33082,N_33178);
or U33863 (N_33863,N_33495,N_33108);
and U33864 (N_33864,N_33113,N_33396);
nor U33865 (N_33865,N_33180,N_33093);
or U33866 (N_33866,N_33292,N_33016);
xor U33867 (N_33867,N_33144,N_33066);
xor U33868 (N_33868,N_33282,N_33301);
nand U33869 (N_33869,N_33403,N_33357);
nor U33870 (N_33870,N_33493,N_33348);
nand U33871 (N_33871,N_33090,N_33445);
xnor U33872 (N_33872,N_33392,N_33208);
and U33873 (N_33873,N_33474,N_33035);
nor U33874 (N_33874,N_33449,N_33026);
or U33875 (N_33875,N_33349,N_33050);
nand U33876 (N_33876,N_33427,N_33230);
xnor U33877 (N_33877,N_33112,N_33466);
and U33878 (N_33878,N_33352,N_33444);
xor U33879 (N_33879,N_33094,N_33287);
or U33880 (N_33880,N_33080,N_33262);
nand U33881 (N_33881,N_33243,N_33189);
and U33882 (N_33882,N_33292,N_33102);
or U33883 (N_33883,N_33495,N_33033);
nor U33884 (N_33884,N_33490,N_33149);
nor U33885 (N_33885,N_33137,N_33047);
or U33886 (N_33886,N_33125,N_33473);
xnor U33887 (N_33887,N_33343,N_33090);
or U33888 (N_33888,N_33304,N_33110);
nor U33889 (N_33889,N_33327,N_33280);
or U33890 (N_33890,N_33179,N_33414);
nor U33891 (N_33891,N_33067,N_33100);
nand U33892 (N_33892,N_33419,N_33059);
and U33893 (N_33893,N_33460,N_33308);
nand U33894 (N_33894,N_33388,N_33060);
or U33895 (N_33895,N_33478,N_33138);
nor U33896 (N_33896,N_33110,N_33137);
nand U33897 (N_33897,N_33454,N_33143);
nor U33898 (N_33898,N_33190,N_33406);
and U33899 (N_33899,N_33033,N_33486);
and U33900 (N_33900,N_33292,N_33206);
nand U33901 (N_33901,N_33336,N_33109);
and U33902 (N_33902,N_33300,N_33414);
nand U33903 (N_33903,N_33023,N_33455);
or U33904 (N_33904,N_33490,N_33378);
xor U33905 (N_33905,N_33134,N_33461);
nand U33906 (N_33906,N_33025,N_33198);
nand U33907 (N_33907,N_33492,N_33112);
nand U33908 (N_33908,N_33386,N_33237);
or U33909 (N_33909,N_33010,N_33132);
nor U33910 (N_33910,N_33484,N_33362);
xor U33911 (N_33911,N_33364,N_33359);
nor U33912 (N_33912,N_33484,N_33150);
or U33913 (N_33913,N_33281,N_33209);
xnor U33914 (N_33914,N_33349,N_33479);
and U33915 (N_33915,N_33181,N_33352);
xor U33916 (N_33916,N_33234,N_33491);
nand U33917 (N_33917,N_33158,N_33250);
and U33918 (N_33918,N_33156,N_33322);
nor U33919 (N_33919,N_33158,N_33337);
and U33920 (N_33920,N_33446,N_33405);
nand U33921 (N_33921,N_33162,N_33230);
and U33922 (N_33922,N_33382,N_33234);
nand U33923 (N_33923,N_33244,N_33211);
xnor U33924 (N_33924,N_33489,N_33352);
nand U33925 (N_33925,N_33058,N_33313);
and U33926 (N_33926,N_33126,N_33336);
nor U33927 (N_33927,N_33431,N_33359);
nand U33928 (N_33928,N_33101,N_33182);
xnor U33929 (N_33929,N_33037,N_33244);
xor U33930 (N_33930,N_33489,N_33142);
nor U33931 (N_33931,N_33071,N_33374);
nand U33932 (N_33932,N_33390,N_33036);
nand U33933 (N_33933,N_33272,N_33060);
and U33934 (N_33934,N_33033,N_33349);
and U33935 (N_33935,N_33228,N_33206);
nand U33936 (N_33936,N_33125,N_33314);
or U33937 (N_33937,N_33016,N_33043);
nand U33938 (N_33938,N_33126,N_33323);
nor U33939 (N_33939,N_33418,N_33289);
nand U33940 (N_33940,N_33073,N_33084);
xnor U33941 (N_33941,N_33107,N_33224);
and U33942 (N_33942,N_33322,N_33098);
nor U33943 (N_33943,N_33441,N_33186);
and U33944 (N_33944,N_33188,N_33498);
or U33945 (N_33945,N_33410,N_33021);
nor U33946 (N_33946,N_33409,N_33315);
xnor U33947 (N_33947,N_33219,N_33285);
nor U33948 (N_33948,N_33165,N_33207);
or U33949 (N_33949,N_33294,N_33407);
or U33950 (N_33950,N_33174,N_33192);
or U33951 (N_33951,N_33273,N_33034);
and U33952 (N_33952,N_33323,N_33086);
or U33953 (N_33953,N_33127,N_33130);
or U33954 (N_33954,N_33496,N_33324);
nand U33955 (N_33955,N_33020,N_33162);
nor U33956 (N_33956,N_33493,N_33005);
xnor U33957 (N_33957,N_33478,N_33389);
nor U33958 (N_33958,N_33385,N_33396);
or U33959 (N_33959,N_33162,N_33379);
nor U33960 (N_33960,N_33431,N_33034);
and U33961 (N_33961,N_33356,N_33306);
nand U33962 (N_33962,N_33198,N_33374);
nor U33963 (N_33963,N_33436,N_33158);
or U33964 (N_33964,N_33057,N_33233);
nand U33965 (N_33965,N_33112,N_33311);
nand U33966 (N_33966,N_33204,N_33030);
or U33967 (N_33967,N_33283,N_33389);
nor U33968 (N_33968,N_33083,N_33004);
xor U33969 (N_33969,N_33271,N_33239);
or U33970 (N_33970,N_33032,N_33335);
or U33971 (N_33971,N_33069,N_33424);
and U33972 (N_33972,N_33464,N_33416);
nand U33973 (N_33973,N_33252,N_33011);
nor U33974 (N_33974,N_33106,N_33450);
and U33975 (N_33975,N_33471,N_33192);
nor U33976 (N_33976,N_33239,N_33211);
or U33977 (N_33977,N_33239,N_33092);
and U33978 (N_33978,N_33043,N_33059);
nand U33979 (N_33979,N_33301,N_33008);
and U33980 (N_33980,N_33201,N_33193);
and U33981 (N_33981,N_33254,N_33191);
or U33982 (N_33982,N_33359,N_33356);
xor U33983 (N_33983,N_33423,N_33459);
or U33984 (N_33984,N_33371,N_33422);
xnor U33985 (N_33985,N_33213,N_33018);
nand U33986 (N_33986,N_33191,N_33490);
xor U33987 (N_33987,N_33460,N_33242);
xor U33988 (N_33988,N_33109,N_33119);
or U33989 (N_33989,N_33273,N_33324);
or U33990 (N_33990,N_33341,N_33207);
or U33991 (N_33991,N_33201,N_33323);
nand U33992 (N_33992,N_33105,N_33396);
or U33993 (N_33993,N_33183,N_33044);
and U33994 (N_33994,N_33444,N_33029);
or U33995 (N_33995,N_33006,N_33449);
nor U33996 (N_33996,N_33225,N_33419);
and U33997 (N_33997,N_33103,N_33480);
xor U33998 (N_33998,N_33321,N_33316);
nand U33999 (N_33999,N_33105,N_33266);
and U34000 (N_34000,N_33507,N_33609);
nand U34001 (N_34001,N_33619,N_33855);
and U34002 (N_34002,N_33898,N_33971);
or U34003 (N_34003,N_33529,N_33901);
or U34004 (N_34004,N_33754,N_33840);
nor U34005 (N_34005,N_33988,N_33767);
xnor U34006 (N_34006,N_33572,N_33586);
xor U34007 (N_34007,N_33624,N_33659);
nor U34008 (N_34008,N_33541,N_33642);
and U34009 (N_34009,N_33933,N_33625);
or U34010 (N_34010,N_33680,N_33641);
xor U34011 (N_34011,N_33501,N_33618);
or U34012 (N_34012,N_33819,N_33548);
xnor U34013 (N_34013,N_33599,N_33549);
nand U34014 (N_34014,N_33651,N_33929);
or U34015 (N_34015,N_33518,N_33513);
or U34016 (N_34016,N_33791,N_33993);
nor U34017 (N_34017,N_33965,N_33861);
nor U34018 (N_34018,N_33869,N_33639);
and U34019 (N_34019,N_33736,N_33908);
xor U34020 (N_34020,N_33950,N_33943);
or U34021 (N_34021,N_33662,N_33813);
or U34022 (N_34022,N_33916,N_33604);
and U34023 (N_34023,N_33796,N_33985);
xnor U34024 (N_34024,N_33877,N_33768);
nand U34025 (N_34025,N_33544,N_33788);
nor U34026 (N_34026,N_33991,N_33834);
or U34027 (N_34027,N_33782,N_33621);
or U34028 (N_34028,N_33966,N_33686);
or U34029 (N_34029,N_33706,N_33808);
nor U34030 (N_34030,N_33821,N_33620);
nor U34031 (N_34031,N_33930,N_33899);
or U34032 (N_34032,N_33725,N_33954);
xor U34033 (N_34033,N_33589,N_33709);
nor U34034 (N_34034,N_33849,N_33672);
or U34035 (N_34035,N_33661,N_33707);
and U34036 (N_34036,N_33718,N_33805);
nand U34037 (N_34037,N_33818,N_33814);
or U34038 (N_34038,N_33986,N_33728);
or U34039 (N_34039,N_33559,N_33558);
or U34040 (N_34040,N_33708,N_33912);
or U34041 (N_34041,N_33983,N_33597);
and U34042 (N_34042,N_33720,N_33932);
xor U34043 (N_34043,N_33536,N_33896);
xnor U34044 (N_34044,N_33775,N_33778);
and U34045 (N_34045,N_33947,N_33922);
and U34046 (N_34046,N_33666,N_33874);
nor U34047 (N_34047,N_33863,N_33810);
nand U34048 (N_34048,N_33967,N_33876);
nor U34049 (N_34049,N_33951,N_33670);
nand U34050 (N_34050,N_33928,N_33521);
and U34051 (N_34051,N_33553,N_33984);
nor U34052 (N_34052,N_33623,N_33601);
nor U34053 (N_34053,N_33615,N_33745);
and U34054 (N_34054,N_33524,N_33523);
nand U34055 (N_34055,N_33534,N_33598);
nor U34056 (N_34056,N_33585,N_33644);
nor U34057 (N_34057,N_33566,N_33531);
nand U34058 (N_34058,N_33793,N_33867);
or U34059 (N_34059,N_33817,N_33504);
or U34060 (N_34060,N_33887,N_33547);
nor U34061 (N_34061,N_33746,N_33786);
nand U34062 (N_34062,N_33935,N_33858);
nor U34063 (N_34063,N_33646,N_33860);
or U34064 (N_34064,N_33873,N_33979);
xnor U34065 (N_34065,N_33723,N_33561);
nor U34066 (N_34066,N_33636,N_33730);
nor U34067 (N_34067,N_33852,N_33937);
nor U34068 (N_34068,N_33578,N_33890);
xnor U34069 (N_34069,N_33797,N_33826);
nand U34070 (N_34070,N_33537,N_33582);
or U34071 (N_34071,N_33889,N_33520);
or U34072 (N_34072,N_33871,N_33833);
and U34073 (N_34073,N_33841,N_33946);
or U34074 (N_34074,N_33649,N_33587);
nand U34075 (N_34075,N_33738,N_33824);
and U34076 (N_34076,N_33570,N_33722);
xor U34077 (N_34077,N_33822,N_33744);
nand U34078 (N_34078,N_33968,N_33635);
xnor U34079 (N_34079,N_33792,N_33975);
or U34080 (N_34080,N_33776,N_33562);
nor U34081 (N_34081,N_33990,N_33881);
xor U34082 (N_34082,N_33920,N_33668);
and U34083 (N_34083,N_33903,N_33964);
nor U34084 (N_34084,N_33811,N_33883);
xnor U34085 (N_34085,N_33512,N_33569);
nor U34086 (N_34086,N_33804,N_33687);
nand U34087 (N_34087,N_33856,N_33839);
nor U34088 (N_34088,N_33679,N_33542);
and U34089 (N_34089,N_33969,N_33757);
nand U34090 (N_34090,N_33742,N_33685);
and U34091 (N_34091,N_33726,N_33576);
nand U34092 (N_34092,N_33823,N_33936);
or U34093 (N_34093,N_33934,N_33892);
nand U34094 (N_34094,N_33705,N_33753);
and U34095 (N_34095,N_33961,N_33550);
and U34096 (N_34096,N_33690,N_33764);
or U34097 (N_34097,N_33584,N_33794);
and U34098 (N_34098,N_33533,N_33882);
nor U34099 (N_34099,N_33581,N_33960);
nor U34100 (N_34100,N_33777,N_33627);
nor U34101 (N_34101,N_33508,N_33747);
and U34102 (N_34102,N_33552,N_33906);
or U34103 (N_34103,N_33634,N_33803);
nor U34104 (N_34104,N_33844,N_33854);
and U34105 (N_34105,N_33694,N_33565);
and U34106 (N_34106,N_33528,N_33829);
nand U34107 (N_34107,N_33614,N_33880);
nand U34108 (N_34108,N_33895,N_33998);
nand U34109 (N_34109,N_33606,N_33830);
nor U34110 (N_34110,N_33592,N_33682);
or U34111 (N_34111,N_33836,N_33645);
nand U34112 (N_34112,N_33905,N_33688);
nand U34113 (N_34113,N_33955,N_33693);
and U34114 (N_34114,N_33952,N_33653);
and U34115 (N_34115,N_33610,N_33941);
nand U34116 (N_34116,N_33981,N_33884);
xnor U34117 (N_34117,N_33827,N_33774);
and U34118 (N_34118,N_33719,N_33732);
xnor U34119 (N_34119,N_33756,N_33848);
nand U34120 (N_34120,N_33652,N_33923);
and U34121 (N_34121,N_33538,N_33626);
nand U34122 (N_34122,N_33807,N_33514);
and U34123 (N_34123,N_33783,N_33866);
and U34124 (N_34124,N_33658,N_33956);
and U34125 (N_34125,N_33798,N_33842);
xor U34126 (N_34126,N_33862,N_33751);
and U34127 (N_34127,N_33716,N_33697);
nor U34128 (N_34128,N_33760,N_33560);
nand U34129 (N_34129,N_33568,N_33510);
nor U34130 (N_34130,N_33580,N_33959);
xnor U34131 (N_34131,N_33973,N_33769);
or U34132 (N_34132,N_33663,N_33825);
and U34133 (N_34133,N_33838,N_33699);
nor U34134 (N_34134,N_33755,N_33766);
or U34135 (N_34135,N_33654,N_33571);
or U34136 (N_34136,N_33859,N_33885);
nand U34137 (N_34137,N_33735,N_33831);
nor U34138 (N_34138,N_33815,N_33588);
nand U34139 (N_34139,N_33927,N_33633);
nand U34140 (N_34140,N_33530,N_33556);
and U34141 (N_34141,N_33657,N_33799);
or U34142 (N_34142,N_33787,N_33888);
nor U34143 (N_34143,N_33689,N_33710);
nand U34144 (N_34144,N_33503,N_33784);
nand U34145 (N_34145,N_33669,N_33678);
and U34146 (N_34146,N_33749,N_33762);
xor U34147 (N_34147,N_33574,N_33847);
xnor U34148 (N_34148,N_33600,N_33593);
xor U34149 (N_34149,N_33795,N_33771);
nor U34150 (N_34150,N_33551,N_33712);
or U34151 (N_34151,N_33925,N_33674);
or U34152 (N_34152,N_33517,N_33527);
or U34153 (N_34153,N_33980,N_33579);
and U34154 (N_34154,N_33972,N_33870);
or U34155 (N_34155,N_33779,N_33978);
and U34156 (N_34156,N_33857,N_33772);
xor U34157 (N_34157,N_33676,N_33907);
or U34158 (N_34158,N_33976,N_33957);
nor U34159 (N_34159,N_33939,N_33773);
or U34160 (N_34160,N_33622,N_33655);
xor U34161 (N_34161,N_33945,N_33886);
xnor U34162 (N_34162,N_33546,N_33820);
xor U34163 (N_34163,N_33698,N_33879);
and U34164 (N_34164,N_33958,N_33702);
or U34165 (N_34165,N_33630,N_33743);
nor U34166 (N_34166,N_33739,N_33893);
xnor U34167 (N_34167,N_33944,N_33902);
nand U34168 (N_34168,N_33949,N_33974);
and U34169 (N_34169,N_33917,N_33809);
and U34170 (N_34170,N_33781,N_33897);
and U34171 (N_34171,N_33734,N_33721);
nor U34172 (N_34172,N_33872,N_33878);
and U34173 (N_34173,N_33785,N_33733);
and U34174 (N_34174,N_33577,N_33656);
nand U34175 (N_34175,N_33864,N_33910);
nor U34176 (N_34176,N_33713,N_33532);
nand U34177 (N_34177,N_33660,N_33590);
xor U34178 (N_34178,N_33843,N_33806);
nand U34179 (N_34179,N_33692,N_33703);
nor U34180 (N_34180,N_33963,N_33594);
nand U34181 (N_34181,N_33748,N_33545);
or U34182 (N_34182,N_33763,N_33802);
or U34183 (N_34183,N_33643,N_33640);
xor U34184 (N_34184,N_33846,N_33554);
nand U34185 (N_34185,N_33714,N_33540);
nor U34186 (N_34186,N_33677,N_33780);
xnor U34187 (N_34187,N_33607,N_33832);
or U34188 (N_34188,N_33696,N_33613);
and U34189 (N_34189,N_33612,N_33539);
and U34190 (N_34190,N_33611,N_33995);
and U34191 (N_34191,N_33801,N_33605);
xor U34192 (N_34192,N_33516,N_33837);
xnor U34193 (N_34193,N_33953,N_33853);
xor U34194 (N_34194,N_33564,N_33638);
nand U34195 (N_34195,N_33525,N_33759);
nor U34196 (N_34196,N_33535,N_33909);
nand U34197 (N_34197,N_33926,N_33790);
nor U34198 (N_34198,N_33695,N_33962);
xor U34199 (N_34199,N_33913,N_33608);
nand U34200 (N_34200,N_33989,N_33629);
or U34201 (N_34201,N_33828,N_33648);
xnor U34202 (N_34202,N_33915,N_33567);
nor U34203 (N_34203,N_33509,N_33812);
nor U34204 (N_34204,N_33602,N_33637);
nand U34205 (N_34205,N_33894,N_33506);
and U34206 (N_34206,N_33505,N_33868);
nor U34207 (N_34207,N_33931,N_33851);
nand U34208 (N_34208,N_33740,N_33684);
nor U34209 (N_34209,N_33816,N_33711);
nor U34210 (N_34210,N_33681,N_33800);
xor U34211 (N_34211,N_33583,N_33691);
xnor U34212 (N_34212,N_33717,N_33835);
or U34213 (N_34213,N_33675,N_33904);
and U34214 (N_34214,N_33500,N_33750);
xor U34215 (N_34215,N_33996,N_33526);
nor U34216 (N_34216,N_33573,N_33997);
nand U34217 (N_34217,N_33999,N_33575);
nor U34218 (N_34218,N_33727,N_33563);
nand U34219 (N_34219,N_33650,N_33671);
nand U34220 (N_34220,N_33770,N_33865);
nand U34221 (N_34221,N_33729,N_33522);
or U34222 (N_34222,N_33765,N_33511);
nand U34223 (N_34223,N_33940,N_33970);
nor U34224 (N_34224,N_33987,N_33631);
and U34225 (N_34225,N_33628,N_33502);
nand U34226 (N_34226,N_33914,N_33557);
nor U34227 (N_34227,N_33982,N_33737);
nand U34228 (N_34228,N_33977,N_33741);
and U34229 (N_34229,N_33596,N_33515);
nor U34230 (N_34230,N_33850,N_33616);
xor U34231 (N_34231,N_33900,N_33992);
xor U34232 (N_34232,N_33683,N_33700);
nand U34233 (N_34233,N_33595,N_33667);
nand U34234 (N_34234,N_33918,N_33724);
xor U34235 (N_34235,N_33603,N_33647);
nand U34236 (N_34236,N_33715,N_33942);
or U34237 (N_34237,N_33519,N_33591);
nor U34238 (N_34238,N_33617,N_33919);
and U34239 (N_34239,N_33891,N_33632);
nand U34240 (N_34240,N_33948,N_33924);
nor U34241 (N_34241,N_33673,N_33701);
and U34242 (N_34242,N_33921,N_33543);
nor U34243 (N_34243,N_33731,N_33875);
nor U34244 (N_34244,N_33664,N_33761);
and U34245 (N_34245,N_33789,N_33845);
nand U34246 (N_34246,N_33555,N_33758);
nor U34247 (N_34247,N_33938,N_33911);
and U34248 (N_34248,N_33704,N_33994);
nand U34249 (N_34249,N_33665,N_33752);
xnor U34250 (N_34250,N_33769,N_33822);
xor U34251 (N_34251,N_33882,N_33594);
and U34252 (N_34252,N_33891,N_33528);
and U34253 (N_34253,N_33785,N_33837);
or U34254 (N_34254,N_33705,N_33761);
or U34255 (N_34255,N_33861,N_33586);
or U34256 (N_34256,N_33880,N_33748);
or U34257 (N_34257,N_33617,N_33992);
and U34258 (N_34258,N_33705,N_33777);
nor U34259 (N_34259,N_33643,N_33842);
and U34260 (N_34260,N_33756,N_33604);
and U34261 (N_34261,N_33795,N_33938);
nand U34262 (N_34262,N_33633,N_33801);
or U34263 (N_34263,N_33539,N_33706);
nand U34264 (N_34264,N_33515,N_33957);
nor U34265 (N_34265,N_33766,N_33757);
or U34266 (N_34266,N_33587,N_33670);
xor U34267 (N_34267,N_33597,N_33889);
or U34268 (N_34268,N_33867,N_33980);
nor U34269 (N_34269,N_33605,N_33735);
and U34270 (N_34270,N_33632,N_33629);
xor U34271 (N_34271,N_33698,N_33614);
nand U34272 (N_34272,N_33663,N_33607);
nor U34273 (N_34273,N_33676,N_33797);
or U34274 (N_34274,N_33675,N_33968);
nor U34275 (N_34275,N_33841,N_33999);
xor U34276 (N_34276,N_33623,N_33924);
nor U34277 (N_34277,N_33936,N_33551);
nor U34278 (N_34278,N_33826,N_33725);
nor U34279 (N_34279,N_33831,N_33973);
or U34280 (N_34280,N_33755,N_33707);
nor U34281 (N_34281,N_33595,N_33503);
nand U34282 (N_34282,N_33676,N_33595);
nor U34283 (N_34283,N_33976,N_33872);
and U34284 (N_34284,N_33615,N_33754);
xor U34285 (N_34285,N_33612,N_33983);
nor U34286 (N_34286,N_33959,N_33558);
xnor U34287 (N_34287,N_33566,N_33744);
xnor U34288 (N_34288,N_33585,N_33538);
nand U34289 (N_34289,N_33704,N_33887);
or U34290 (N_34290,N_33528,N_33903);
or U34291 (N_34291,N_33503,N_33942);
and U34292 (N_34292,N_33574,N_33992);
or U34293 (N_34293,N_33780,N_33522);
or U34294 (N_34294,N_33806,N_33565);
and U34295 (N_34295,N_33852,N_33734);
xnor U34296 (N_34296,N_33974,N_33914);
or U34297 (N_34297,N_33697,N_33715);
or U34298 (N_34298,N_33741,N_33500);
and U34299 (N_34299,N_33941,N_33602);
or U34300 (N_34300,N_33560,N_33511);
and U34301 (N_34301,N_33963,N_33518);
nand U34302 (N_34302,N_33678,N_33620);
nand U34303 (N_34303,N_33859,N_33963);
or U34304 (N_34304,N_33877,N_33666);
or U34305 (N_34305,N_33614,N_33798);
or U34306 (N_34306,N_33945,N_33730);
xor U34307 (N_34307,N_33974,N_33524);
nand U34308 (N_34308,N_33734,N_33828);
and U34309 (N_34309,N_33763,N_33925);
and U34310 (N_34310,N_33507,N_33894);
and U34311 (N_34311,N_33920,N_33940);
and U34312 (N_34312,N_33589,N_33794);
nor U34313 (N_34313,N_33835,N_33834);
nor U34314 (N_34314,N_33689,N_33767);
nor U34315 (N_34315,N_33793,N_33775);
nor U34316 (N_34316,N_33727,N_33981);
nor U34317 (N_34317,N_33837,N_33746);
xor U34318 (N_34318,N_33526,N_33829);
nand U34319 (N_34319,N_33901,N_33810);
and U34320 (N_34320,N_33961,N_33558);
or U34321 (N_34321,N_33950,N_33648);
xnor U34322 (N_34322,N_33793,N_33937);
xnor U34323 (N_34323,N_33542,N_33540);
and U34324 (N_34324,N_33942,N_33704);
and U34325 (N_34325,N_33902,N_33567);
or U34326 (N_34326,N_33850,N_33943);
nand U34327 (N_34327,N_33888,N_33854);
nand U34328 (N_34328,N_33643,N_33610);
xnor U34329 (N_34329,N_33648,N_33971);
and U34330 (N_34330,N_33790,N_33596);
xor U34331 (N_34331,N_33851,N_33553);
nor U34332 (N_34332,N_33611,N_33811);
nor U34333 (N_34333,N_33615,N_33634);
nand U34334 (N_34334,N_33976,N_33666);
nand U34335 (N_34335,N_33943,N_33708);
and U34336 (N_34336,N_33648,N_33625);
nand U34337 (N_34337,N_33526,N_33555);
or U34338 (N_34338,N_33997,N_33788);
nand U34339 (N_34339,N_33619,N_33544);
nor U34340 (N_34340,N_33936,N_33629);
xnor U34341 (N_34341,N_33838,N_33764);
xnor U34342 (N_34342,N_33851,N_33657);
and U34343 (N_34343,N_33919,N_33632);
xnor U34344 (N_34344,N_33839,N_33851);
nand U34345 (N_34345,N_33553,N_33864);
nor U34346 (N_34346,N_33900,N_33907);
nor U34347 (N_34347,N_33624,N_33711);
xor U34348 (N_34348,N_33687,N_33779);
and U34349 (N_34349,N_33616,N_33979);
nor U34350 (N_34350,N_33781,N_33903);
nand U34351 (N_34351,N_33681,N_33679);
or U34352 (N_34352,N_33589,N_33586);
nand U34353 (N_34353,N_33759,N_33710);
nand U34354 (N_34354,N_33692,N_33748);
nor U34355 (N_34355,N_33691,N_33874);
xnor U34356 (N_34356,N_33718,N_33685);
or U34357 (N_34357,N_33642,N_33536);
nand U34358 (N_34358,N_33927,N_33556);
nand U34359 (N_34359,N_33628,N_33907);
and U34360 (N_34360,N_33924,N_33691);
nor U34361 (N_34361,N_33649,N_33848);
and U34362 (N_34362,N_33628,N_33936);
nand U34363 (N_34363,N_33656,N_33650);
nor U34364 (N_34364,N_33859,N_33957);
nand U34365 (N_34365,N_33965,N_33602);
nand U34366 (N_34366,N_33879,N_33748);
nand U34367 (N_34367,N_33789,N_33565);
nor U34368 (N_34368,N_33502,N_33853);
xor U34369 (N_34369,N_33878,N_33502);
nand U34370 (N_34370,N_33610,N_33601);
and U34371 (N_34371,N_33805,N_33709);
and U34372 (N_34372,N_33866,N_33861);
xnor U34373 (N_34373,N_33613,N_33655);
and U34374 (N_34374,N_33923,N_33832);
nand U34375 (N_34375,N_33830,N_33975);
and U34376 (N_34376,N_33578,N_33807);
xor U34377 (N_34377,N_33917,N_33853);
or U34378 (N_34378,N_33677,N_33787);
and U34379 (N_34379,N_33700,N_33744);
nor U34380 (N_34380,N_33534,N_33788);
and U34381 (N_34381,N_33507,N_33739);
or U34382 (N_34382,N_33921,N_33741);
nor U34383 (N_34383,N_33888,N_33957);
nand U34384 (N_34384,N_33832,N_33534);
xor U34385 (N_34385,N_33913,N_33548);
nor U34386 (N_34386,N_33909,N_33641);
nor U34387 (N_34387,N_33588,N_33758);
and U34388 (N_34388,N_33710,N_33667);
nor U34389 (N_34389,N_33763,N_33873);
or U34390 (N_34390,N_33809,N_33745);
nand U34391 (N_34391,N_33755,N_33745);
or U34392 (N_34392,N_33744,N_33657);
nand U34393 (N_34393,N_33584,N_33737);
and U34394 (N_34394,N_33737,N_33858);
xnor U34395 (N_34395,N_33747,N_33689);
xnor U34396 (N_34396,N_33666,N_33956);
nor U34397 (N_34397,N_33619,N_33684);
nand U34398 (N_34398,N_33635,N_33713);
nand U34399 (N_34399,N_33910,N_33513);
nor U34400 (N_34400,N_33946,N_33637);
or U34401 (N_34401,N_33837,N_33627);
xnor U34402 (N_34402,N_33921,N_33955);
nand U34403 (N_34403,N_33821,N_33518);
nand U34404 (N_34404,N_33983,N_33671);
nand U34405 (N_34405,N_33789,N_33611);
xor U34406 (N_34406,N_33827,N_33555);
or U34407 (N_34407,N_33901,N_33894);
xor U34408 (N_34408,N_33954,N_33702);
and U34409 (N_34409,N_33818,N_33637);
xnor U34410 (N_34410,N_33776,N_33642);
nor U34411 (N_34411,N_33606,N_33879);
or U34412 (N_34412,N_33724,N_33905);
and U34413 (N_34413,N_33726,N_33607);
or U34414 (N_34414,N_33660,N_33639);
and U34415 (N_34415,N_33716,N_33786);
and U34416 (N_34416,N_33897,N_33677);
or U34417 (N_34417,N_33693,N_33503);
xnor U34418 (N_34418,N_33752,N_33835);
and U34419 (N_34419,N_33613,N_33654);
and U34420 (N_34420,N_33791,N_33779);
or U34421 (N_34421,N_33518,N_33781);
xnor U34422 (N_34422,N_33555,N_33571);
xor U34423 (N_34423,N_33733,N_33954);
nor U34424 (N_34424,N_33535,N_33551);
nor U34425 (N_34425,N_33819,N_33980);
nor U34426 (N_34426,N_33874,N_33837);
nor U34427 (N_34427,N_33697,N_33990);
nor U34428 (N_34428,N_33999,N_33545);
nand U34429 (N_34429,N_33577,N_33560);
nor U34430 (N_34430,N_33957,N_33786);
nand U34431 (N_34431,N_33767,N_33771);
and U34432 (N_34432,N_33552,N_33818);
and U34433 (N_34433,N_33575,N_33553);
nor U34434 (N_34434,N_33552,N_33829);
or U34435 (N_34435,N_33669,N_33761);
or U34436 (N_34436,N_33855,N_33706);
and U34437 (N_34437,N_33924,N_33681);
nand U34438 (N_34438,N_33756,N_33875);
and U34439 (N_34439,N_33951,N_33817);
and U34440 (N_34440,N_33665,N_33786);
nor U34441 (N_34441,N_33961,N_33775);
xor U34442 (N_34442,N_33733,N_33585);
xor U34443 (N_34443,N_33743,N_33887);
or U34444 (N_34444,N_33908,N_33867);
or U34445 (N_34445,N_33665,N_33509);
nand U34446 (N_34446,N_33699,N_33965);
nand U34447 (N_34447,N_33571,N_33626);
xor U34448 (N_34448,N_33657,N_33515);
nand U34449 (N_34449,N_33721,N_33937);
or U34450 (N_34450,N_33723,N_33534);
and U34451 (N_34451,N_33903,N_33520);
nand U34452 (N_34452,N_33943,N_33908);
and U34453 (N_34453,N_33833,N_33976);
or U34454 (N_34454,N_33893,N_33603);
or U34455 (N_34455,N_33919,N_33669);
nand U34456 (N_34456,N_33706,N_33667);
nand U34457 (N_34457,N_33914,N_33620);
nor U34458 (N_34458,N_33852,N_33721);
and U34459 (N_34459,N_33562,N_33690);
or U34460 (N_34460,N_33644,N_33638);
nand U34461 (N_34461,N_33886,N_33534);
xnor U34462 (N_34462,N_33569,N_33871);
nand U34463 (N_34463,N_33981,N_33725);
xnor U34464 (N_34464,N_33815,N_33851);
or U34465 (N_34465,N_33667,N_33868);
nand U34466 (N_34466,N_33516,N_33726);
or U34467 (N_34467,N_33971,N_33576);
nand U34468 (N_34468,N_33768,N_33943);
and U34469 (N_34469,N_33648,N_33808);
or U34470 (N_34470,N_33853,N_33993);
or U34471 (N_34471,N_33837,N_33526);
or U34472 (N_34472,N_33959,N_33701);
or U34473 (N_34473,N_33974,N_33782);
nor U34474 (N_34474,N_33501,N_33630);
xnor U34475 (N_34475,N_33761,N_33960);
and U34476 (N_34476,N_33933,N_33635);
and U34477 (N_34477,N_33632,N_33971);
or U34478 (N_34478,N_33862,N_33826);
nand U34479 (N_34479,N_33728,N_33849);
nand U34480 (N_34480,N_33817,N_33587);
xnor U34481 (N_34481,N_33899,N_33977);
nor U34482 (N_34482,N_33544,N_33938);
nor U34483 (N_34483,N_33522,N_33898);
nand U34484 (N_34484,N_33873,N_33941);
and U34485 (N_34485,N_33755,N_33534);
xor U34486 (N_34486,N_33882,N_33859);
nor U34487 (N_34487,N_33665,N_33545);
or U34488 (N_34488,N_33585,N_33923);
or U34489 (N_34489,N_33568,N_33719);
and U34490 (N_34490,N_33706,N_33796);
and U34491 (N_34491,N_33542,N_33645);
and U34492 (N_34492,N_33558,N_33581);
or U34493 (N_34493,N_33792,N_33639);
xor U34494 (N_34494,N_33576,N_33686);
nor U34495 (N_34495,N_33879,N_33814);
nor U34496 (N_34496,N_33640,N_33833);
xor U34497 (N_34497,N_33661,N_33730);
or U34498 (N_34498,N_33762,N_33574);
xnor U34499 (N_34499,N_33935,N_33902);
xnor U34500 (N_34500,N_34005,N_34416);
and U34501 (N_34501,N_34004,N_34375);
xnor U34502 (N_34502,N_34303,N_34244);
or U34503 (N_34503,N_34079,N_34238);
nand U34504 (N_34504,N_34421,N_34318);
or U34505 (N_34505,N_34358,N_34446);
xnor U34506 (N_34506,N_34168,N_34135);
nand U34507 (N_34507,N_34192,N_34127);
and U34508 (N_34508,N_34143,N_34206);
xnor U34509 (N_34509,N_34454,N_34415);
nor U34510 (N_34510,N_34456,N_34360);
nand U34511 (N_34511,N_34184,N_34202);
nand U34512 (N_34512,N_34027,N_34103);
nor U34513 (N_34513,N_34367,N_34315);
xnor U34514 (N_34514,N_34099,N_34424);
or U34515 (N_34515,N_34074,N_34408);
or U34516 (N_34516,N_34341,N_34425);
and U34517 (N_34517,N_34444,N_34073);
nor U34518 (N_34518,N_34194,N_34000);
or U34519 (N_34519,N_34348,N_34092);
or U34520 (N_34520,N_34326,N_34115);
xor U34521 (N_34521,N_34188,N_34152);
and U34522 (N_34522,N_34384,N_34230);
or U34523 (N_34523,N_34376,N_34123);
and U34524 (N_34524,N_34086,N_34003);
nand U34525 (N_34525,N_34101,N_34149);
and U34526 (N_34526,N_34025,N_34329);
nand U34527 (N_34527,N_34273,N_34093);
nand U34528 (N_34528,N_34497,N_34331);
nand U34529 (N_34529,N_34110,N_34130);
and U34530 (N_34530,N_34288,N_34055);
nand U34531 (N_34531,N_34183,N_34429);
xnor U34532 (N_34532,N_34471,N_34451);
nand U34533 (N_34533,N_34419,N_34483);
nor U34534 (N_34534,N_34404,N_34452);
xnor U34535 (N_34535,N_34438,N_34434);
and U34536 (N_34536,N_34380,N_34498);
xnor U34537 (N_34537,N_34053,N_34282);
nand U34538 (N_34538,N_34138,N_34021);
xor U34539 (N_34539,N_34235,N_34010);
and U34540 (N_34540,N_34270,N_34211);
nor U34541 (N_34541,N_34255,N_34436);
nor U34542 (N_34542,N_34447,N_34204);
or U34543 (N_34543,N_34140,N_34124);
nand U34544 (N_34544,N_34155,N_34088);
nand U34545 (N_34545,N_34063,N_34495);
nand U34546 (N_34546,N_34491,N_34199);
nor U34547 (N_34547,N_34215,N_34233);
nor U34548 (N_34548,N_34281,N_34117);
nand U34549 (N_34549,N_34208,N_34223);
nand U34550 (N_34550,N_34040,N_34195);
and U34551 (N_34551,N_34359,N_34156);
and U34552 (N_34552,N_34467,N_34252);
xnor U34553 (N_34553,N_34344,N_34276);
nand U34554 (N_34554,N_34098,N_34104);
nand U34555 (N_34555,N_34033,N_34248);
xnor U34556 (N_34556,N_34200,N_34144);
xor U34557 (N_34557,N_34317,N_34263);
xor U34558 (N_34558,N_34141,N_34388);
nand U34559 (N_34559,N_34391,N_34442);
nor U34560 (N_34560,N_34189,N_34378);
and U34561 (N_34561,N_34251,N_34395);
nor U34562 (N_34562,N_34046,N_34089);
nor U34563 (N_34563,N_34488,N_34214);
nand U34564 (N_34564,N_34243,N_34136);
or U34565 (N_34565,N_34038,N_34173);
xor U34566 (N_34566,N_34197,N_34049);
and U34567 (N_34567,N_34325,N_34026);
and U34568 (N_34568,N_34170,N_34187);
xor U34569 (N_34569,N_34108,N_34056);
nor U34570 (N_34570,N_34213,N_34316);
xnor U34571 (N_34571,N_34019,N_34286);
xor U34572 (N_34572,N_34234,N_34043);
nor U34573 (N_34573,N_34091,N_34013);
nand U34574 (N_34574,N_34011,N_34285);
and U34575 (N_34575,N_34227,N_34403);
xnor U34576 (N_34576,N_34209,N_34128);
or U34577 (N_34577,N_34499,N_34496);
and U34578 (N_34578,N_34241,N_34486);
and U34579 (N_34579,N_34292,N_34356);
or U34580 (N_34580,N_34062,N_34295);
xor U34581 (N_34581,N_34362,N_34269);
nor U34582 (N_34582,N_34036,N_34245);
or U34583 (N_34583,N_34431,N_34453);
nor U34584 (N_34584,N_34057,N_34312);
nor U34585 (N_34585,N_34153,N_34232);
nand U34586 (N_34586,N_34253,N_34080);
nand U34587 (N_34587,N_34008,N_34015);
or U34588 (N_34588,N_34353,N_34284);
nand U34589 (N_34589,N_34361,N_34385);
or U34590 (N_34590,N_34205,N_34352);
xnor U34591 (N_34591,N_34068,N_34222);
nor U34592 (N_34592,N_34300,N_34085);
nor U34593 (N_34593,N_34133,N_34158);
nand U34594 (N_34594,N_34272,N_34116);
xnor U34595 (N_34595,N_34337,N_34476);
or U34596 (N_34596,N_34210,N_34106);
nand U34597 (N_34597,N_34406,N_34069);
xor U34598 (N_34598,N_34364,N_34335);
and U34599 (N_34599,N_34370,N_34417);
or U34600 (N_34600,N_34259,N_34455);
nand U34601 (N_34601,N_34287,N_34162);
xnor U34602 (N_34602,N_34163,N_34394);
xnor U34603 (N_34603,N_34299,N_34392);
nand U34604 (N_34604,N_34340,N_34226);
xor U34605 (N_34605,N_34097,N_34381);
nand U34606 (N_34606,N_34441,N_34107);
nor U34607 (N_34607,N_34409,N_34028);
xnor U34608 (N_34608,N_34389,N_34024);
nor U34609 (N_34609,N_34032,N_34161);
nand U34610 (N_34610,N_34065,N_34231);
or U34611 (N_34611,N_34469,N_34332);
or U34612 (N_34612,N_34308,N_34440);
nand U34613 (N_34613,N_34422,N_34041);
xnor U34614 (N_34614,N_34368,N_34363);
nor U34615 (N_34615,N_34338,N_34347);
and U34616 (N_34616,N_34035,N_34058);
nor U34617 (N_34617,N_34030,N_34077);
nand U34618 (N_34618,N_34430,N_34167);
and U34619 (N_34619,N_34023,N_34059);
nand U34620 (N_34620,N_34377,N_34250);
xor U34621 (N_34621,N_34054,N_34051);
nand U34622 (N_34622,N_34094,N_34387);
or U34623 (N_34623,N_34007,N_34012);
nand U34624 (N_34624,N_34307,N_34072);
or U34625 (N_34625,N_34264,N_34102);
or U34626 (N_34626,N_34443,N_34475);
and U34627 (N_34627,N_34428,N_34061);
xnor U34628 (N_34628,N_34279,N_34218);
or U34629 (N_34629,N_34267,N_34132);
nand U34630 (N_34630,N_34018,N_34224);
or U34631 (N_34631,N_34246,N_34111);
and U34632 (N_34632,N_34151,N_34240);
nand U34633 (N_34633,N_34171,N_34355);
nand U34634 (N_34634,N_34480,N_34304);
xnor U34635 (N_34635,N_34175,N_34229);
nand U34636 (N_34636,N_34181,N_34298);
and U34637 (N_34637,N_34017,N_34472);
and U34638 (N_34638,N_34477,N_34020);
nand U34639 (N_34639,N_34334,N_34071);
nand U34640 (N_34640,N_34142,N_34311);
nor U34641 (N_34641,N_34009,N_34228);
or U34642 (N_34642,N_34397,N_34082);
or U34643 (N_34643,N_34256,N_34042);
or U34644 (N_34644,N_34407,N_34494);
xnor U34645 (N_34645,N_34154,N_34216);
nor U34646 (N_34646,N_34122,N_34283);
xnor U34647 (N_34647,N_34309,N_34484);
or U34648 (N_34648,N_34321,N_34067);
nand U34649 (N_34649,N_34029,N_34176);
nor U34650 (N_34650,N_34435,N_34212);
and U34651 (N_34651,N_34217,N_34147);
nor U34652 (N_34652,N_34177,N_34450);
xor U34653 (N_34653,N_34157,N_34075);
or U34654 (N_34654,N_34474,N_34180);
nand U34655 (N_34655,N_34150,N_34119);
and U34656 (N_34656,N_34249,N_34393);
xor U34657 (N_34657,N_34191,N_34169);
or U34658 (N_34658,N_34277,N_34294);
and U34659 (N_34659,N_34260,N_34405);
nor U34660 (N_34660,N_34301,N_34120);
and U34661 (N_34661,N_34134,N_34289);
xor U34662 (N_34662,N_34349,N_34398);
nand U34663 (N_34663,N_34047,N_34070);
and U34664 (N_34664,N_34266,N_34468);
and U34665 (N_34665,N_34083,N_34293);
or U34666 (N_34666,N_34310,N_34478);
xor U34667 (N_34667,N_34060,N_34296);
and U34668 (N_34668,N_34372,N_34463);
or U34669 (N_34669,N_34411,N_34182);
nor U34670 (N_34670,N_34034,N_34165);
or U34671 (N_34671,N_34339,N_34433);
nor U34672 (N_34672,N_34445,N_34172);
or U34673 (N_34673,N_34137,N_34371);
xnor U34674 (N_34674,N_34268,N_34351);
nand U34675 (N_34675,N_34333,N_34114);
nand U34676 (N_34676,N_34420,N_34139);
xor U34677 (N_34677,N_34418,N_34002);
or U34678 (N_34678,N_34470,N_34305);
nand U34679 (N_34679,N_34159,N_34328);
and U34680 (N_34680,N_34373,N_34365);
xnor U34681 (N_34681,N_34146,N_34109);
nand U34682 (N_34682,N_34178,N_34126);
and U34683 (N_34683,N_34160,N_34048);
or U34684 (N_34684,N_34458,N_34105);
or U34685 (N_34685,N_34196,N_34280);
xnor U34686 (N_34686,N_34350,N_34278);
or U34687 (N_34687,N_34466,N_34369);
or U34688 (N_34688,N_34112,N_34464);
and U34689 (N_34689,N_34313,N_34490);
nor U34690 (N_34690,N_34258,N_34439);
or U34691 (N_34691,N_34437,N_34118);
xor U34692 (N_34692,N_34066,N_34399);
xor U34693 (N_34693,N_34050,N_34193);
and U34694 (N_34694,N_34297,N_34262);
nor U34695 (N_34695,N_34457,N_34247);
nor U34696 (N_34696,N_34131,N_34037);
or U34697 (N_34697,N_34039,N_34465);
xnor U34698 (N_34698,N_34096,N_34401);
xnor U34699 (N_34699,N_34129,N_34022);
nand U34700 (N_34700,N_34236,N_34459);
xor U34701 (N_34701,N_34125,N_34336);
and U34702 (N_34702,N_34045,N_34179);
and U34703 (N_34703,N_34271,N_34383);
nor U34704 (N_34704,N_34261,N_34319);
xnor U34705 (N_34705,N_34320,N_34427);
nor U34706 (N_34706,N_34221,N_34100);
or U34707 (N_34707,N_34482,N_34327);
nand U34708 (N_34708,N_34201,N_34410);
xnor U34709 (N_34709,N_34076,N_34064);
nor U34710 (N_34710,N_34095,N_34354);
and U34711 (N_34711,N_34052,N_34219);
xnor U34712 (N_34712,N_34044,N_34390);
nor U34713 (N_34713,N_34113,N_34449);
or U34714 (N_34714,N_34220,N_34084);
xor U34715 (N_34715,N_34487,N_34400);
or U34716 (N_34716,N_34090,N_34014);
xor U34717 (N_34717,N_34016,N_34031);
nor U34718 (N_34718,N_34225,N_34148);
nand U34719 (N_34719,N_34423,N_34081);
nand U34720 (N_34720,N_34121,N_34481);
nand U34721 (N_34721,N_34290,N_34461);
or U34722 (N_34722,N_34257,N_34473);
xnor U34723 (N_34723,N_34379,N_34342);
or U34724 (N_34724,N_34396,N_34448);
nand U34725 (N_34725,N_34001,N_34185);
nand U34726 (N_34726,N_34254,N_34186);
nand U34727 (N_34727,N_34302,N_34386);
and U34728 (N_34728,N_34237,N_34242);
xor U34729 (N_34729,N_34374,N_34203);
nor U34730 (N_34730,N_34412,N_34314);
nand U34731 (N_34731,N_34426,N_34460);
nor U34732 (N_34732,N_34492,N_34485);
xnor U34733 (N_34733,N_34198,N_34078);
nor U34734 (N_34734,N_34190,N_34322);
nor U34735 (N_34735,N_34366,N_34174);
nor U34736 (N_34736,N_34087,N_34306);
or U34737 (N_34737,N_34166,N_34291);
and U34738 (N_34738,N_34432,N_34274);
nor U34739 (N_34739,N_34343,N_34265);
or U34740 (N_34740,N_34413,N_34414);
xnor U34741 (N_34741,N_34345,N_34145);
xor U34742 (N_34742,N_34330,N_34346);
or U34743 (N_34743,N_34493,N_34275);
and U34744 (N_34744,N_34357,N_34164);
or U34745 (N_34745,N_34479,N_34402);
nor U34746 (N_34746,N_34324,N_34382);
xor U34747 (N_34747,N_34489,N_34239);
xnor U34748 (N_34748,N_34323,N_34462);
xor U34749 (N_34749,N_34006,N_34207);
nor U34750 (N_34750,N_34056,N_34208);
nand U34751 (N_34751,N_34376,N_34383);
nor U34752 (N_34752,N_34432,N_34312);
or U34753 (N_34753,N_34197,N_34499);
xnor U34754 (N_34754,N_34031,N_34495);
or U34755 (N_34755,N_34469,N_34408);
or U34756 (N_34756,N_34076,N_34215);
xnor U34757 (N_34757,N_34471,N_34292);
nor U34758 (N_34758,N_34445,N_34432);
and U34759 (N_34759,N_34279,N_34016);
nor U34760 (N_34760,N_34264,N_34459);
nor U34761 (N_34761,N_34461,N_34237);
or U34762 (N_34762,N_34008,N_34159);
nor U34763 (N_34763,N_34387,N_34304);
or U34764 (N_34764,N_34000,N_34170);
nand U34765 (N_34765,N_34457,N_34356);
xor U34766 (N_34766,N_34483,N_34459);
or U34767 (N_34767,N_34392,N_34239);
nor U34768 (N_34768,N_34363,N_34118);
xor U34769 (N_34769,N_34160,N_34214);
or U34770 (N_34770,N_34236,N_34335);
nand U34771 (N_34771,N_34481,N_34184);
xnor U34772 (N_34772,N_34267,N_34230);
and U34773 (N_34773,N_34240,N_34163);
and U34774 (N_34774,N_34427,N_34243);
nor U34775 (N_34775,N_34411,N_34142);
nor U34776 (N_34776,N_34061,N_34404);
and U34777 (N_34777,N_34025,N_34358);
nand U34778 (N_34778,N_34460,N_34292);
nor U34779 (N_34779,N_34431,N_34484);
xnor U34780 (N_34780,N_34483,N_34421);
or U34781 (N_34781,N_34089,N_34333);
nor U34782 (N_34782,N_34385,N_34454);
nand U34783 (N_34783,N_34417,N_34219);
or U34784 (N_34784,N_34037,N_34296);
nand U34785 (N_34785,N_34183,N_34082);
nand U34786 (N_34786,N_34178,N_34176);
nor U34787 (N_34787,N_34448,N_34360);
and U34788 (N_34788,N_34030,N_34443);
nor U34789 (N_34789,N_34309,N_34082);
or U34790 (N_34790,N_34256,N_34152);
nor U34791 (N_34791,N_34150,N_34478);
xnor U34792 (N_34792,N_34130,N_34245);
nand U34793 (N_34793,N_34196,N_34369);
or U34794 (N_34794,N_34005,N_34386);
or U34795 (N_34795,N_34339,N_34168);
and U34796 (N_34796,N_34360,N_34110);
or U34797 (N_34797,N_34296,N_34272);
xor U34798 (N_34798,N_34413,N_34321);
nand U34799 (N_34799,N_34394,N_34302);
xor U34800 (N_34800,N_34444,N_34452);
nand U34801 (N_34801,N_34434,N_34331);
nor U34802 (N_34802,N_34406,N_34134);
and U34803 (N_34803,N_34168,N_34219);
nand U34804 (N_34804,N_34073,N_34211);
xor U34805 (N_34805,N_34402,N_34358);
nand U34806 (N_34806,N_34423,N_34334);
nand U34807 (N_34807,N_34347,N_34178);
nor U34808 (N_34808,N_34070,N_34458);
nor U34809 (N_34809,N_34235,N_34368);
and U34810 (N_34810,N_34326,N_34178);
nor U34811 (N_34811,N_34248,N_34128);
or U34812 (N_34812,N_34443,N_34241);
nand U34813 (N_34813,N_34461,N_34008);
nor U34814 (N_34814,N_34164,N_34277);
and U34815 (N_34815,N_34498,N_34008);
xnor U34816 (N_34816,N_34021,N_34361);
nand U34817 (N_34817,N_34241,N_34348);
nor U34818 (N_34818,N_34037,N_34393);
or U34819 (N_34819,N_34192,N_34493);
and U34820 (N_34820,N_34257,N_34270);
xnor U34821 (N_34821,N_34445,N_34496);
nor U34822 (N_34822,N_34384,N_34456);
and U34823 (N_34823,N_34345,N_34174);
nand U34824 (N_34824,N_34324,N_34111);
nor U34825 (N_34825,N_34019,N_34386);
and U34826 (N_34826,N_34012,N_34355);
nor U34827 (N_34827,N_34310,N_34463);
or U34828 (N_34828,N_34332,N_34158);
nor U34829 (N_34829,N_34190,N_34112);
nor U34830 (N_34830,N_34046,N_34317);
nand U34831 (N_34831,N_34498,N_34130);
nor U34832 (N_34832,N_34153,N_34054);
xnor U34833 (N_34833,N_34260,N_34102);
xnor U34834 (N_34834,N_34128,N_34448);
and U34835 (N_34835,N_34044,N_34426);
nor U34836 (N_34836,N_34383,N_34269);
and U34837 (N_34837,N_34496,N_34242);
nor U34838 (N_34838,N_34272,N_34376);
nand U34839 (N_34839,N_34339,N_34125);
nand U34840 (N_34840,N_34065,N_34015);
nand U34841 (N_34841,N_34289,N_34484);
nand U34842 (N_34842,N_34444,N_34331);
and U34843 (N_34843,N_34080,N_34006);
or U34844 (N_34844,N_34069,N_34051);
nor U34845 (N_34845,N_34497,N_34011);
and U34846 (N_34846,N_34203,N_34339);
xor U34847 (N_34847,N_34481,N_34325);
and U34848 (N_34848,N_34188,N_34262);
nand U34849 (N_34849,N_34290,N_34471);
and U34850 (N_34850,N_34168,N_34058);
nor U34851 (N_34851,N_34372,N_34417);
and U34852 (N_34852,N_34318,N_34193);
xor U34853 (N_34853,N_34106,N_34014);
and U34854 (N_34854,N_34408,N_34392);
nand U34855 (N_34855,N_34021,N_34116);
and U34856 (N_34856,N_34018,N_34189);
xnor U34857 (N_34857,N_34372,N_34348);
nor U34858 (N_34858,N_34470,N_34313);
and U34859 (N_34859,N_34464,N_34431);
xor U34860 (N_34860,N_34336,N_34463);
or U34861 (N_34861,N_34197,N_34328);
or U34862 (N_34862,N_34235,N_34331);
and U34863 (N_34863,N_34498,N_34201);
xor U34864 (N_34864,N_34217,N_34134);
xor U34865 (N_34865,N_34452,N_34023);
or U34866 (N_34866,N_34332,N_34146);
and U34867 (N_34867,N_34465,N_34040);
nor U34868 (N_34868,N_34490,N_34044);
nand U34869 (N_34869,N_34236,N_34150);
nor U34870 (N_34870,N_34062,N_34036);
or U34871 (N_34871,N_34092,N_34158);
and U34872 (N_34872,N_34392,N_34050);
nor U34873 (N_34873,N_34237,N_34317);
or U34874 (N_34874,N_34424,N_34141);
and U34875 (N_34875,N_34318,N_34013);
xor U34876 (N_34876,N_34465,N_34412);
nor U34877 (N_34877,N_34135,N_34042);
nor U34878 (N_34878,N_34083,N_34264);
nor U34879 (N_34879,N_34345,N_34381);
nand U34880 (N_34880,N_34410,N_34166);
nor U34881 (N_34881,N_34305,N_34362);
nand U34882 (N_34882,N_34189,N_34215);
nand U34883 (N_34883,N_34042,N_34465);
and U34884 (N_34884,N_34444,N_34032);
xnor U34885 (N_34885,N_34091,N_34009);
or U34886 (N_34886,N_34443,N_34403);
nor U34887 (N_34887,N_34220,N_34368);
nor U34888 (N_34888,N_34425,N_34270);
or U34889 (N_34889,N_34345,N_34348);
nor U34890 (N_34890,N_34445,N_34231);
or U34891 (N_34891,N_34272,N_34361);
or U34892 (N_34892,N_34154,N_34231);
and U34893 (N_34893,N_34423,N_34466);
xor U34894 (N_34894,N_34032,N_34403);
xor U34895 (N_34895,N_34374,N_34071);
and U34896 (N_34896,N_34467,N_34309);
or U34897 (N_34897,N_34443,N_34089);
and U34898 (N_34898,N_34172,N_34429);
nand U34899 (N_34899,N_34201,N_34007);
nor U34900 (N_34900,N_34376,N_34340);
nor U34901 (N_34901,N_34350,N_34396);
nand U34902 (N_34902,N_34370,N_34447);
xor U34903 (N_34903,N_34140,N_34232);
nand U34904 (N_34904,N_34126,N_34140);
nand U34905 (N_34905,N_34312,N_34206);
and U34906 (N_34906,N_34063,N_34007);
nand U34907 (N_34907,N_34294,N_34256);
xnor U34908 (N_34908,N_34477,N_34441);
nand U34909 (N_34909,N_34100,N_34383);
and U34910 (N_34910,N_34233,N_34166);
xnor U34911 (N_34911,N_34144,N_34131);
xor U34912 (N_34912,N_34288,N_34068);
and U34913 (N_34913,N_34043,N_34039);
xor U34914 (N_34914,N_34499,N_34194);
and U34915 (N_34915,N_34464,N_34417);
and U34916 (N_34916,N_34069,N_34356);
or U34917 (N_34917,N_34494,N_34019);
or U34918 (N_34918,N_34392,N_34006);
nand U34919 (N_34919,N_34012,N_34063);
xor U34920 (N_34920,N_34064,N_34276);
nor U34921 (N_34921,N_34131,N_34429);
nand U34922 (N_34922,N_34133,N_34399);
or U34923 (N_34923,N_34397,N_34171);
nor U34924 (N_34924,N_34359,N_34485);
nand U34925 (N_34925,N_34065,N_34373);
nor U34926 (N_34926,N_34018,N_34230);
nand U34927 (N_34927,N_34249,N_34262);
nand U34928 (N_34928,N_34341,N_34141);
xnor U34929 (N_34929,N_34159,N_34331);
nand U34930 (N_34930,N_34155,N_34021);
nor U34931 (N_34931,N_34267,N_34192);
nor U34932 (N_34932,N_34481,N_34483);
or U34933 (N_34933,N_34248,N_34267);
and U34934 (N_34934,N_34418,N_34335);
and U34935 (N_34935,N_34177,N_34379);
and U34936 (N_34936,N_34238,N_34383);
or U34937 (N_34937,N_34100,N_34351);
or U34938 (N_34938,N_34073,N_34494);
nor U34939 (N_34939,N_34393,N_34112);
xnor U34940 (N_34940,N_34491,N_34459);
or U34941 (N_34941,N_34428,N_34395);
nor U34942 (N_34942,N_34493,N_34396);
xor U34943 (N_34943,N_34306,N_34067);
nand U34944 (N_34944,N_34252,N_34485);
xor U34945 (N_34945,N_34274,N_34472);
or U34946 (N_34946,N_34006,N_34290);
and U34947 (N_34947,N_34354,N_34138);
xor U34948 (N_34948,N_34355,N_34030);
and U34949 (N_34949,N_34331,N_34124);
xnor U34950 (N_34950,N_34015,N_34221);
and U34951 (N_34951,N_34311,N_34432);
or U34952 (N_34952,N_34087,N_34408);
xnor U34953 (N_34953,N_34381,N_34009);
or U34954 (N_34954,N_34074,N_34008);
nor U34955 (N_34955,N_34487,N_34354);
or U34956 (N_34956,N_34377,N_34395);
xor U34957 (N_34957,N_34245,N_34266);
nor U34958 (N_34958,N_34215,N_34379);
nor U34959 (N_34959,N_34316,N_34256);
xor U34960 (N_34960,N_34383,N_34413);
xnor U34961 (N_34961,N_34244,N_34071);
nand U34962 (N_34962,N_34178,N_34383);
xnor U34963 (N_34963,N_34313,N_34046);
nand U34964 (N_34964,N_34249,N_34177);
nor U34965 (N_34965,N_34212,N_34391);
or U34966 (N_34966,N_34039,N_34326);
nor U34967 (N_34967,N_34407,N_34395);
and U34968 (N_34968,N_34365,N_34281);
nor U34969 (N_34969,N_34407,N_34367);
and U34970 (N_34970,N_34368,N_34037);
and U34971 (N_34971,N_34242,N_34290);
xor U34972 (N_34972,N_34296,N_34428);
or U34973 (N_34973,N_34020,N_34044);
nand U34974 (N_34974,N_34141,N_34483);
and U34975 (N_34975,N_34070,N_34095);
xor U34976 (N_34976,N_34415,N_34188);
and U34977 (N_34977,N_34410,N_34356);
or U34978 (N_34978,N_34232,N_34276);
xor U34979 (N_34979,N_34130,N_34070);
and U34980 (N_34980,N_34330,N_34378);
and U34981 (N_34981,N_34421,N_34175);
or U34982 (N_34982,N_34346,N_34202);
nor U34983 (N_34983,N_34481,N_34170);
nor U34984 (N_34984,N_34403,N_34063);
and U34985 (N_34985,N_34344,N_34139);
nand U34986 (N_34986,N_34214,N_34059);
nor U34987 (N_34987,N_34033,N_34000);
xor U34988 (N_34988,N_34334,N_34157);
or U34989 (N_34989,N_34180,N_34449);
xnor U34990 (N_34990,N_34271,N_34281);
xnor U34991 (N_34991,N_34049,N_34471);
or U34992 (N_34992,N_34113,N_34300);
nand U34993 (N_34993,N_34061,N_34343);
and U34994 (N_34994,N_34403,N_34023);
and U34995 (N_34995,N_34143,N_34196);
nand U34996 (N_34996,N_34158,N_34387);
nand U34997 (N_34997,N_34329,N_34117);
xor U34998 (N_34998,N_34086,N_34103);
or U34999 (N_34999,N_34309,N_34357);
nand U35000 (N_35000,N_34723,N_34695);
or U35001 (N_35001,N_34854,N_34881);
nand U35002 (N_35002,N_34755,N_34795);
or U35003 (N_35003,N_34853,N_34749);
and U35004 (N_35004,N_34935,N_34816);
nand U35005 (N_35005,N_34883,N_34951);
nand U35006 (N_35006,N_34763,N_34778);
and U35007 (N_35007,N_34945,N_34963);
or U35008 (N_35008,N_34706,N_34910);
xnor U35009 (N_35009,N_34826,N_34739);
and U35010 (N_35010,N_34964,N_34995);
nand U35011 (N_35011,N_34685,N_34909);
xnor U35012 (N_35012,N_34893,N_34752);
xnor U35013 (N_35013,N_34738,N_34861);
and U35014 (N_35014,N_34998,N_34505);
xnor U35015 (N_35015,N_34650,N_34905);
and U35016 (N_35016,N_34788,N_34707);
xnor U35017 (N_35017,N_34570,N_34939);
and U35018 (N_35018,N_34686,N_34711);
nand U35019 (N_35019,N_34720,N_34625);
and U35020 (N_35020,N_34936,N_34990);
xnor U35021 (N_35021,N_34892,N_34700);
nand U35022 (N_35022,N_34934,N_34802);
nor U35023 (N_35023,N_34967,N_34803);
xor U35024 (N_35024,N_34585,N_34888);
or U35025 (N_35025,N_34798,N_34528);
xor U35026 (N_35026,N_34651,N_34593);
or U35027 (N_35027,N_34860,N_34732);
and U35028 (N_35028,N_34774,N_34846);
nand U35029 (N_35029,N_34506,N_34626);
or U35030 (N_35030,N_34722,N_34607);
and U35031 (N_35031,N_34710,N_34712);
xor U35032 (N_35032,N_34799,N_34938);
and U35033 (N_35033,N_34960,N_34823);
nor U35034 (N_35034,N_34927,N_34699);
xnor U35035 (N_35035,N_34573,N_34825);
nand U35036 (N_35036,N_34561,N_34996);
nor U35037 (N_35037,N_34745,N_34543);
and U35038 (N_35038,N_34628,N_34867);
and U35039 (N_35039,N_34737,N_34609);
xor U35040 (N_35040,N_34517,N_34701);
or U35041 (N_35041,N_34821,N_34828);
nor U35042 (N_35042,N_34809,N_34510);
and U35043 (N_35043,N_34591,N_34672);
nor U35044 (N_35044,N_34621,N_34636);
xor U35045 (N_35045,N_34662,N_34847);
xor U35046 (N_35046,N_34688,N_34834);
nand U35047 (N_35047,N_34843,N_34954);
and U35048 (N_35048,N_34742,N_34999);
or U35049 (N_35049,N_34741,N_34574);
xnor U35050 (N_35050,N_34839,N_34895);
nor U35051 (N_35051,N_34988,N_34582);
or U35052 (N_35052,N_34536,N_34751);
nand U35053 (N_35053,N_34776,N_34652);
nor U35054 (N_35054,N_34872,N_34703);
or U35055 (N_35055,N_34970,N_34586);
or U35056 (N_35056,N_34790,N_34684);
nand U35057 (N_35057,N_34793,N_34544);
or U35058 (N_35058,N_34777,N_34693);
and U35059 (N_35059,N_34978,N_34917);
xor U35060 (N_35060,N_34566,N_34962);
nand U35061 (N_35061,N_34618,N_34949);
or U35062 (N_35062,N_34982,N_34503);
nand U35063 (N_35063,N_34541,N_34523);
nor U35064 (N_35064,N_34810,N_34835);
or U35065 (N_35065,N_34911,N_34583);
xor U35066 (N_35066,N_34555,N_34740);
or U35067 (N_35067,N_34914,N_34950);
nor U35068 (N_35068,N_34972,N_34687);
xnor U35069 (N_35069,N_34973,N_34596);
nor U35070 (N_35070,N_34829,N_34635);
xnor U35071 (N_35071,N_34649,N_34511);
xnor U35072 (N_35072,N_34524,N_34946);
nor U35073 (N_35073,N_34731,N_34932);
and U35074 (N_35074,N_34780,N_34668);
and U35075 (N_35075,N_34841,N_34762);
or U35076 (N_35076,N_34806,N_34758);
xor U35077 (N_35077,N_34901,N_34539);
nor U35078 (N_35078,N_34754,N_34862);
or U35079 (N_35079,N_34500,N_34808);
or U35080 (N_35080,N_34886,N_34768);
nor U35081 (N_35081,N_34880,N_34772);
and U35082 (N_35082,N_34550,N_34871);
and U35083 (N_35083,N_34616,N_34985);
xor U35084 (N_35084,N_34726,N_34876);
nand U35085 (N_35085,N_34734,N_34540);
xnor U35086 (N_35086,N_34655,N_34767);
and U35087 (N_35087,N_34783,N_34851);
and U35088 (N_35088,N_34965,N_34606);
nor U35089 (N_35089,N_34771,N_34733);
and U35090 (N_35090,N_34522,N_34680);
nor U35091 (N_35091,N_34530,N_34631);
xnor U35092 (N_35092,N_34559,N_34844);
or U35093 (N_35093,N_34903,N_34981);
and U35094 (N_35094,N_34805,N_34761);
nor U35095 (N_35095,N_34997,N_34943);
or U35096 (N_35096,N_34610,N_34991);
xor U35097 (N_35097,N_34564,N_34989);
nand U35098 (N_35098,N_34614,N_34885);
and U35099 (N_35099,N_34894,N_34904);
or U35100 (N_35100,N_34671,N_34504);
nand U35101 (N_35101,N_34532,N_34842);
xnor U35102 (N_35102,N_34956,N_34715);
and U35103 (N_35103,N_34595,N_34908);
nor U35104 (N_35104,N_34928,N_34906);
or U35105 (N_35105,N_34801,N_34833);
xnor U35106 (N_35106,N_34526,N_34845);
or U35107 (N_35107,N_34660,N_34764);
xnor U35108 (N_35108,N_34830,N_34959);
or U35109 (N_35109,N_34879,N_34681);
xnor U35110 (N_35110,N_34576,N_34527);
xnor U35111 (N_35111,N_34900,N_34537);
nand U35112 (N_35112,N_34629,N_34804);
nor U35113 (N_35113,N_34800,N_34918);
nor U35114 (N_35114,N_34840,N_34584);
and U35115 (N_35115,N_34624,N_34924);
xnor U35116 (N_35116,N_34877,N_34902);
xor U35117 (N_35117,N_34704,N_34615);
xnor U35118 (N_35118,N_34766,N_34588);
or U35119 (N_35119,N_34980,N_34957);
or U35120 (N_35120,N_34728,N_34553);
and U35121 (N_35121,N_34944,N_34608);
or U35122 (N_35122,N_34630,N_34942);
or U35123 (N_35123,N_34887,N_34868);
and U35124 (N_35124,N_34508,N_34966);
nor U35125 (N_35125,N_34533,N_34640);
and U35126 (N_35126,N_34916,N_34592);
nor U35127 (N_35127,N_34765,N_34746);
nor U35128 (N_35128,N_34848,N_34647);
xnor U35129 (N_35129,N_34565,N_34604);
nand U35130 (N_35130,N_34569,N_34994);
xor U35131 (N_35131,N_34501,N_34557);
xor U35132 (N_35132,N_34797,N_34875);
and U35133 (N_35133,N_34874,N_34661);
xor U35134 (N_35134,N_34716,N_34969);
nor U35135 (N_35135,N_34787,N_34611);
or U35136 (N_35136,N_34992,N_34925);
and U35137 (N_35137,N_34775,N_34919);
or U35138 (N_35138,N_34976,N_34760);
nor U35139 (N_35139,N_34676,N_34708);
nand U35140 (N_35140,N_34789,N_34702);
and U35141 (N_35141,N_34941,N_34663);
nand U35142 (N_35142,N_34898,N_34856);
or U35143 (N_35143,N_34824,N_34929);
nand U35144 (N_35144,N_34792,N_34859);
and U35145 (N_35145,N_34646,N_34870);
and U35146 (N_35146,N_34884,N_34933);
xnor U35147 (N_35147,N_34547,N_34753);
nand U35148 (N_35148,N_34784,N_34679);
and U35149 (N_35149,N_34852,N_34642);
and U35150 (N_35150,N_34832,N_34556);
nand U35151 (N_35151,N_34613,N_34587);
nand U35152 (N_35152,N_34718,N_34838);
and U35153 (N_35153,N_34896,N_34743);
xnor U35154 (N_35154,N_34725,N_34858);
nand U35155 (N_35155,N_34975,N_34987);
or U35156 (N_35156,N_34721,N_34667);
nand U35157 (N_35157,N_34594,N_34907);
nor U35158 (N_35158,N_34882,N_34785);
nand U35159 (N_35159,N_34568,N_34915);
nor U35160 (N_35160,N_34648,N_34664);
nor U35161 (N_35161,N_34786,N_34534);
or U35162 (N_35162,N_34654,N_34682);
and U35163 (N_35163,N_34836,N_34571);
xor U35164 (N_35164,N_34698,N_34560);
and U35165 (N_35165,N_34580,N_34705);
or U35166 (N_35166,N_34669,N_34947);
and U35167 (N_35167,N_34552,N_34675);
nor U35168 (N_35168,N_34577,N_34612);
xnor U35169 (N_35169,N_34502,N_34831);
and U35170 (N_35170,N_34729,N_34756);
xnor U35171 (N_35171,N_34599,N_34549);
nor U35172 (N_35172,N_34757,N_34891);
nor U35173 (N_35173,N_34563,N_34779);
nor U35174 (N_35174,N_34986,N_34750);
nor U35175 (N_35175,N_34974,N_34813);
xor U35176 (N_35176,N_34713,N_34633);
nor U35177 (N_35177,N_34665,N_34694);
nand U35178 (N_35178,N_34794,N_34878);
and U35179 (N_35179,N_34730,N_34769);
nor U35180 (N_35180,N_34819,N_34634);
nand U35181 (N_35181,N_34638,N_34627);
or U35182 (N_35182,N_34677,N_34678);
and U35183 (N_35183,N_34656,N_34509);
nand U35184 (N_35184,N_34657,N_34578);
and U35185 (N_35185,N_34516,N_34822);
or U35186 (N_35186,N_34692,N_34619);
nand U35187 (N_35187,N_34659,N_34683);
or U35188 (N_35188,N_34558,N_34719);
and U35189 (N_35189,N_34773,N_34748);
xor U35190 (N_35190,N_34697,N_34968);
or U35191 (N_35191,N_34645,N_34952);
nand U35192 (N_35192,N_34953,N_34873);
nand U35193 (N_35193,N_34865,N_34670);
or U35194 (N_35194,N_34590,N_34581);
nand U35195 (N_35195,N_34744,N_34589);
nor U35196 (N_35196,N_34572,N_34827);
and U35197 (N_35197,N_34983,N_34600);
nand U35198 (N_35198,N_34617,N_34796);
and U35199 (N_35199,N_34538,N_34890);
nand U35200 (N_35200,N_34696,N_34545);
nor U35201 (N_35201,N_34770,N_34850);
nor U35202 (N_35202,N_34554,N_34811);
nor U35203 (N_35203,N_34747,N_34782);
nor U35204 (N_35204,N_34515,N_34512);
nor U35205 (N_35205,N_34689,N_34863);
or U35206 (N_35206,N_34622,N_34759);
or U35207 (N_35207,N_34736,N_34632);
nor U35208 (N_35208,N_34535,N_34507);
xor U35209 (N_35209,N_34542,N_34922);
nand U35210 (N_35210,N_34984,N_34546);
or U35211 (N_35211,N_34921,N_34727);
nor U35212 (N_35212,N_34817,N_34857);
or U35213 (N_35213,N_34815,N_34837);
xnor U35214 (N_35214,N_34913,N_34807);
nand U35215 (N_35215,N_34724,N_34518);
and U35216 (N_35216,N_34666,N_34519);
xor U35217 (N_35217,N_34714,N_34601);
or U35218 (N_35218,N_34781,N_34551);
and U35219 (N_35219,N_34931,N_34575);
nand U35220 (N_35220,N_34855,N_34889);
xnor U35221 (N_35221,N_34639,N_34948);
and U35222 (N_35222,N_34993,N_34525);
or U35223 (N_35223,N_34864,N_34602);
nand U35224 (N_35224,N_34644,N_34623);
and U35225 (N_35225,N_34812,N_34930);
xor U35226 (N_35226,N_34603,N_34620);
xnor U35227 (N_35227,N_34579,N_34691);
or U35228 (N_35228,N_34562,N_34597);
xor U35229 (N_35229,N_34717,N_34658);
and U35230 (N_35230,N_34977,N_34529);
nor U35231 (N_35231,N_34598,N_34567);
xor U35232 (N_35232,N_34940,N_34866);
nand U35233 (N_35233,N_34791,N_34814);
or U35234 (N_35234,N_34690,N_34514);
and U35235 (N_35235,N_34735,N_34641);
xnor U35236 (N_35236,N_34912,N_34849);
nand U35237 (N_35237,N_34674,N_34958);
and U35238 (N_35238,N_34979,N_34899);
or U35239 (N_35239,N_34673,N_34521);
nor U35240 (N_35240,N_34920,N_34923);
nand U35241 (N_35241,N_34513,N_34605);
nand U35242 (N_35242,N_34520,N_34820);
xor U35243 (N_35243,N_34653,N_34531);
nor U35244 (N_35244,N_34937,N_34897);
and U35245 (N_35245,N_34709,N_34869);
or U35246 (N_35246,N_34643,N_34818);
or U35247 (N_35247,N_34548,N_34961);
xor U35248 (N_35248,N_34637,N_34955);
nand U35249 (N_35249,N_34971,N_34926);
and U35250 (N_35250,N_34979,N_34501);
or U35251 (N_35251,N_34926,N_34500);
and U35252 (N_35252,N_34819,N_34602);
nand U35253 (N_35253,N_34649,N_34630);
nand U35254 (N_35254,N_34836,N_34932);
nor U35255 (N_35255,N_34703,N_34736);
and U35256 (N_35256,N_34779,N_34806);
nor U35257 (N_35257,N_34740,N_34530);
xor U35258 (N_35258,N_34719,N_34926);
or U35259 (N_35259,N_34601,N_34715);
and U35260 (N_35260,N_34899,N_34911);
or U35261 (N_35261,N_34836,N_34742);
or U35262 (N_35262,N_34960,N_34669);
nand U35263 (N_35263,N_34765,N_34799);
or U35264 (N_35264,N_34794,N_34637);
nand U35265 (N_35265,N_34585,N_34568);
nor U35266 (N_35266,N_34611,N_34688);
nor U35267 (N_35267,N_34777,N_34987);
xnor U35268 (N_35268,N_34512,N_34647);
nor U35269 (N_35269,N_34795,N_34907);
nor U35270 (N_35270,N_34976,N_34704);
and U35271 (N_35271,N_34730,N_34670);
nor U35272 (N_35272,N_34588,N_34836);
and U35273 (N_35273,N_34680,N_34997);
nor U35274 (N_35274,N_34816,N_34690);
and U35275 (N_35275,N_34778,N_34935);
or U35276 (N_35276,N_34679,N_34561);
or U35277 (N_35277,N_34543,N_34727);
nor U35278 (N_35278,N_34870,N_34975);
nand U35279 (N_35279,N_34530,N_34914);
nor U35280 (N_35280,N_34521,N_34645);
or U35281 (N_35281,N_34967,N_34812);
nand U35282 (N_35282,N_34572,N_34626);
xor U35283 (N_35283,N_34836,N_34838);
and U35284 (N_35284,N_34931,N_34851);
and U35285 (N_35285,N_34990,N_34841);
or U35286 (N_35286,N_34513,N_34896);
or U35287 (N_35287,N_34643,N_34860);
xor U35288 (N_35288,N_34566,N_34512);
nor U35289 (N_35289,N_34588,N_34648);
or U35290 (N_35290,N_34963,N_34975);
nand U35291 (N_35291,N_34564,N_34657);
xor U35292 (N_35292,N_34877,N_34591);
nand U35293 (N_35293,N_34742,N_34712);
and U35294 (N_35294,N_34664,N_34857);
or U35295 (N_35295,N_34870,N_34736);
nor U35296 (N_35296,N_34737,N_34976);
nor U35297 (N_35297,N_34503,N_34682);
nor U35298 (N_35298,N_34786,N_34591);
xor U35299 (N_35299,N_34580,N_34744);
or U35300 (N_35300,N_34950,N_34996);
nor U35301 (N_35301,N_34954,N_34905);
and U35302 (N_35302,N_34818,N_34652);
or U35303 (N_35303,N_34557,N_34931);
xnor U35304 (N_35304,N_34828,N_34506);
nor U35305 (N_35305,N_34793,N_34636);
nand U35306 (N_35306,N_34998,N_34654);
xnor U35307 (N_35307,N_34591,N_34630);
and U35308 (N_35308,N_34656,N_34615);
or U35309 (N_35309,N_34632,N_34611);
xor U35310 (N_35310,N_34945,N_34942);
xnor U35311 (N_35311,N_34517,N_34754);
and U35312 (N_35312,N_34564,N_34881);
xor U35313 (N_35313,N_34812,N_34823);
xnor U35314 (N_35314,N_34752,N_34563);
nand U35315 (N_35315,N_34585,N_34745);
or U35316 (N_35316,N_34864,N_34790);
nor U35317 (N_35317,N_34833,N_34518);
xnor U35318 (N_35318,N_34661,N_34985);
or U35319 (N_35319,N_34909,N_34554);
xnor U35320 (N_35320,N_34966,N_34545);
nand U35321 (N_35321,N_34763,N_34805);
nor U35322 (N_35322,N_34508,N_34874);
and U35323 (N_35323,N_34933,N_34522);
nor U35324 (N_35324,N_34557,N_34882);
or U35325 (N_35325,N_34666,N_34753);
and U35326 (N_35326,N_34548,N_34842);
nand U35327 (N_35327,N_34501,N_34735);
or U35328 (N_35328,N_34869,N_34829);
nor U35329 (N_35329,N_34881,N_34975);
xnor U35330 (N_35330,N_34634,N_34848);
nand U35331 (N_35331,N_34803,N_34735);
and U35332 (N_35332,N_34726,N_34695);
nand U35333 (N_35333,N_34625,N_34792);
nor U35334 (N_35334,N_34940,N_34578);
nand U35335 (N_35335,N_34509,N_34944);
xor U35336 (N_35336,N_34782,N_34591);
xor U35337 (N_35337,N_34798,N_34573);
and U35338 (N_35338,N_34663,N_34991);
xor U35339 (N_35339,N_34941,N_34682);
nor U35340 (N_35340,N_34644,N_34638);
nor U35341 (N_35341,N_34731,N_34963);
or U35342 (N_35342,N_34803,N_34734);
or U35343 (N_35343,N_34828,N_34665);
or U35344 (N_35344,N_34519,N_34676);
xor U35345 (N_35345,N_34870,N_34570);
nand U35346 (N_35346,N_34928,N_34857);
or U35347 (N_35347,N_34654,N_34745);
and U35348 (N_35348,N_34535,N_34632);
and U35349 (N_35349,N_34992,N_34527);
nand U35350 (N_35350,N_34904,N_34659);
or U35351 (N_35351,N_34661,N_34938);
and U35352 (N_35352,N_34532,N_34815);
nor U35353 (N_35353,N_34871,N_34758);
xor U35354 (N_35354,N_34892,N_34977);
nor U35355 (N_35355,N_34606,N_34744);
nand U35356 (N_35356,N_34531,N_34804);
xor U35357 (N_35357,N_34535,N_34791);
nand U35358 (N_35358,N_34699,N_34870);
or U35359 (N_35359,N_34826,N_34607);
xnor U35360 (N_35360,N_34755,N_34916);
nor U35361 (N_35361,N_34951,N_34895);
xnor U35362 (N_35362,N_34920,N_34793);
xnor U35363 (N_35363,N_34789,N_34984);
xnor U35364 (N_35364,N_34695,N_34810);
nand U35365 (N_35365,N_34570,N_34695);
and U35366 (N_35366,N_34523,N_34700);
or U35367 (N_35367,N_34882,N_34827);
xor U35368 (N_35368,N_34556,N_34616);
nor U35369 (N_35369,N_34817,N_34530);
xor U35370 (N_35370,N_34951,N_34594);
and U35371 (N_35371,N_34921,N_34597);
nand U35372 (N_35372,N_34541,N_34625);
or U35373 (N_35373,N_34921,N_34876);
or U35374 (N_35374,N_34803,N_34769);
and U35375 (N_35375,N_34969,N_34523);
nor U35376 (N_35376,N_34500,N_34932);
nand U35377 (N_35377,N_34520,N_34900);
nor U35378 (N_35378,N_34937,N_34886);
nor U35379 (N_35379,N_34758,N_34703);
nand U35380 (N_35380,N_34550,N_34545);
or U35381 (N_35381,N_34717,N_34512);
and U35382 (N_35382,N_34715,N_34859);
xor U35383 (N_35383,N_34515,N_34923);
and U35384 (N_35384,N_34822,N_34935);
or U35385 (N_35385,N_34665,N_34639);
nor U35386 (N_35386,N_34646,N_34836);
and U35387 (N_35387,N_34857,N_34846);
xnor U35388 (N_35388,N_34805,N_34874);
xor U35389 (N_35389,N_34549,N_34914);
and U35390 (N_35390,N_34712,N_34647);
xor U35391 (N_35391,N_34808,N_34622);
nor U35392 (N_35392,N_34644,N_34755);
or U35393 (N_35393,N_34811,N_34850);
or U35394 (N_35394,N_34975,N_34884);
or U35395 (N_35395,N_34807,N_34637);
nand U35396 (N_35396,N_34500,N_34776);
and U35397 (N_35397,N_34808,N_34530);
nand U35398 (N_35398,N_34557,N_34980);
nand U35399 (N_35399,N_34858,N_34736);
or U35400 (N_35400,N_34943,N_34578);
xor U35401 (N_35401,N_34749,N_34877);
nand U35402 (N_35402,N_34636,N_34873);
and U35403 (N_35403,N_34586,N_34874);
and U35404 (N_35404,N_34809,N_34668);
nor U35405 (N_35405,N_34502,N_34967);
nand U35406 (N_35406,N_34862,N_34592);
xnor U35407 (N_35407,N_34940,N_34864);
or U35408 (N_35408,N_34514,N_34774);
and U35409 (N_35409,N_34571,N_34548);
xor U35410 (N_35410,N_34928,N_34672);
or U35411 (N_35411,N_34564,N_34638);
and U35412 (N_35412,N_34670,N_34948);
xor U35413 (N_35413,N_34604,N_34954);
or U35414 (N_35414,N_34923,N_34794);
or U35415 (N_35415,N_34899,N_34898);
nor U35416 (N_35416,N_34726,N_34565);
nor U35417 (N_35417,N_34848,N_34799);
xor U35418 (N_35418,N_34546,N_34812);
and U35419 (N_35419,N_34873,N_34825);
xnor U35420 (N_35420,N_34865,N_34969);
or U35421 (N_35421,N_34899,N_34951);
xor U35422 (N_35422,N_34913,N_34593);
nand U35423 (N_35423,N_34561,N_34601);
xnor U35424 (N_35424,N_34794,N_34979);
nor U35425 (N_35425,N_34621,N_34805);
and U35426 (N_35426,N_34765,N_34713);
nor U35427 (N_35427,N_34685,N_34735);
and U35428 (N_35428,N_34663,N_34851);
nor U35429 (N_35429,N_34989,N_34848);
xnor U35430 (N_35430,N_34965,N_34540);
or U35431 (N_35431,N_34570,N_34508);
or U35432 (N_35432,N_34726,N_34581);
xor U35433 (N_35433,N_34946,N_34630);
nand U35434 (N_35434,N_34875,N_34680);
nand U35435 (N_35435,N_34637,N_34529);
nor U35436 (N_35436,N_34740,N_34805);
or U35437 (N_35437,N_34772,N_34743);
and U35438 (N_35438,N_34570,N_34892);
nand U35439 (N_35439,N_34594,N_34785);
xor U35440 (N_35440,N_34829,N_34940);
xor U35441 (N_35441,N_34556,N_34533);
or U35442 (N_35442,N_34976,N_34944);
and U35443 (N_35443,N_34899,N_34983);
nand U35444 (N_35444,N_34969,N_34957);
and U35445 (N_35445,N_34576,N_34656);
nand U35446 (N_35446,N_34603,N_34902);
xor U35447 (N_35447,N_34715,N_34845);
and U35448 (N_35448,N_34817,N_34815);
and U35449 (N_35449,N_34573,N_34873);
or U35450 (N_35450,N_34869,N_34842);
nor U35451 (N_35451,N_34947,N_34742);
or U35452 (N_35452,N_34905,N_34965);
xnor U35453 (N_35453,N_34977,N_34628);
and U35454 (N_35454,N_34702,N_34985);
and U35455 (N_35455,N_34890,N_34553);
or U35456 (N_35456,N_34575,N_34654);
or U35457 (N_35457,N_34782,N_34797);
nor U35458 (N_35458,N_34894,N_34635);
and U35459 (N_35459,N_34638,N_34517);
xor U35460 (N_35460,N_34982,N_34969);
xor U35461 (N_35461,N_34730,N_34750);
xnor U35462 (N_35462,N_34831,N_34901);
and U35463 (N_35463,N_34788,N_34671);
nand U35464 (N_35464,N_34959,N_34711);
and U35465 (N_35465,N_34746,N_34736);
or U35466 (N_35466,N_34810,N_34940);
nor U35467 (N_35467,N_34820,N_34574);
nand U35468 (N_35468,N_34626,N_34764);
xor U35469 (N_35469,N_34956,N_34719);
xor U35470 (N_35470,N_34921,N_34917);
nor U35471 (N_35471,N_34534,N_34887);
or U35472 (N_35472,N_34700,N_34894);
and U35473 (N_35473,N_34808,N_34675);
or U35474 (N_35474,N_34968,N_34715);
nand U35475 (N_35475,N_34645,N_34810);
xnor U35476 (N_35476,N_34559,N_34876);
or U35477 (N_35477,N_34884,N_34740);
or U35478 (N_35478,N_34587,N_34581);
xnor U35479 (N_35479,N_34978,N_34622);
xnor U35480 (N_35480,N_34753,N_34751);
xor U35481 (N_35481,N_34949,N_34568);
or U35482 (N_35482,N_34927,N_34698);
or U35483 (N_35483,N_34802,N_34898);
xnor U35484 (N_35484,N_34910,N_34954);
nand U35485 (N_35485,N_34519,N_34552);
nand U35486 (N_35486,N_34832,N_34983);
and U35487 (N_35487,N_34613,N_34891);
nand U35488 (N_35488,N_34901,N_34879);
and U35489 (N_35489,N_34838,N_34714);
nor U35490 (N_35490,N_34611,N_34931);
nor U35491 (N_35491,N_34752,N_34664);
or U35492 (N_35492,N_34835,N_34579);
and U35493 (N_35493,N_34819,N_34539);
or U35494 (N_35494,N_34836,N_34541);
and U35495 (N_35495,N_34574,N_34818);
or U35496 (N_35496,N_34624,N_34819);
xor U35497 (N_35497,N_34689,N_34502);
or U35498 (N_35498,N_34503,N_34523);
xor U35499 (N_35499,N_34867,N_34784);
nor U35500 (N_35500,N_35209,N_35210);
and U35501 (N_35501,N_35426,N_35479);
nor U35502 (N_35502,N_35365,N_35086);
nor U35503 (N_35503,N_35369,N_35101);
xor U35504 (N_35504,N_35115,N_35113);
nor U35505 (N_35505,N_35129,N_35457);
and U35506 (N_35506,N_35010,N_35316);
nand U35507 (N_35507,N_35036,N_35363);
xor U35508 (N_35508,N_35130,N_35243);
and U35509 (N_35509,N_35228,N_35362);
xnor U35510 (N_35510,N_35471,N_35372);
and U35511 (N_35511,N_35073,N_35399);
nand U35512 (N_35512,N_35070,N_35337);
nor U35513 (N_35513,N_35049,N_35205);
nor U35514 (N_35514,N_35047,N_35152);
and U35515 (N_35515,N_35343,N_35176);
nor U35516 (N_35516,N_35392,N_35389);
nor U35517 (N_35517,N_35112,N_35134);
xnor U35518 (N_35518,N_35037,N_35231);
or U35519 (N_35519,N_35242,N_35254);
nand U35520 (N_35520,N_35227,N_35040);
or U35521 (N_35521,N_35138,N_35436);
nor U35522 (N_35522,N_35361,N_35433);
or U35523 (N_35523,N_35018,N_35168);
nor U35524 (N_35524,N_35307,N_35038);
xnor U35525 (N_35525,N_35009,N_35470);
and U35526 (N_35526,N_35249,N_35345);
nand U35527 (N_35527,N_35095,N_35482);
nor U35528 (N_35528,N_35405,N_35376);
nand U35529 (N_35529,N_35067,N_35078);
and U35530 (N_35530,N_35258,N_35478);
and U35531 (N_35531,N_35270,N_35180);
or U35532 (N_35532,N_35380,N_35177);
or U35533 (N_35533,N_35481,N_35005);
and U35534 (N_35534,N_35306,N_35189);
and U35535 (N_35535,N_35207,N_35089);
nand U35536 (N_35536,N_35214,N_35483);
nor U35537 (N_35537,N_35052,N_35021);
nand U35538 (N_35538,N_35443,N_35072);
or U35539 (N_35539,N_35229,N_35348);
and U35540 (N_35540,N_35486,N_35050);
nand U35541 (N_35541,N_35248,N_35082);
xor U35542 (N_35542,N_35409,N_35293);
nand U35543 (N_35543,N_35442,N_35450);
xnor U35544 (N_35544,N_35401,N_35335);
and U35545 (N_35545,N_35211,N_35489);
and U35546 (N_35546,N_35480,N_35090);
and U35547 (N_35547,N_35104,N_35069);
nor U35548 (N_35548,N_35032,N_35358);
and U35549 (N_35549,N_35385,N_35497);
nand U35550 (N_35550,N_35011,N_35267);
and U35551 (N_35551,N_35271,N_35445);
or U35552 (N_35552,N_35240,N_35429);
xor U35553 (N_35553,N_35292,N_35212);
nand U35554 (N_35554,N_35336,N_35342);
nand U35555 (N_35555,N_35490,N_35034);
nor U35556 (N_35556,N_35331,N_35384);
nand U35557 (N_35557,N_35237,N_35048);
nand U35558 (N_35558,N_35432,N_35390);
or U35559 (N_35559,N_35057,N_35493);
nand U35560 (N_35560,N_35276,N_35300);
xnor U35561 (N_35561,N_35419,N_35066);
xnor U35562 (N_35562,N_35423,N_35430);
xor U35563 (N_35563,N_35294,N_35378);
nor U35564 (N_35564,N_35427,N_35455);
xor U35565 (N_35565,N_35288,N_35025);
nand U35566 (N_35566,N_35351,N_35280);
nand U35567 (N_35567,N_35076,N_35127);
and U35568 (N_35568,N_35060,N_35002);
xor U35569 (N_35569,N_35219,N_35435);
xnor U35570 (N_35570,N_35041,N_35422);
or U35571 (N_35571,N_35169,N_35183);
and U35572 (N_35572,N_35145,N_35408);
or U35573 (N_35573,N_35269,N_35261);
nor U35574 (N_35574,N_35016,N_35226);
and U35575 (N_35575,N_35403,N_35023);
or U35576 (N_35576,N_35260,N_35364);
nor U35577 (N_35577,N_35441,N_35461);
nor U35578 (N_35578,N_35417,N_35323);
nand U35579 (N_35579,N_35327,N_35264);
nand U35580 (N_35580,N_35383,N_35467);
xnor U35581 (N_35581,N_35175,N_35246);
and U35582 (N_35582,N_35239,N_35099);
xnor U35583 (N_35583,N_35084,N_35062);
xor U35584 (N_35584,N_35199,N_35125);
and U35585 (N_35585,N_35094,N_35424);
nor U35586 (N_35586,N_35301,N_35252);
xor U35587 (N_35587,N_35302,N_35371);
or U35588 (N_35588,N_35290,N_35488);
nor U35589 (N_35589,N_35349,N_35459);
xor U35590 (N_35590,N_35106,N_35298);
nor U35591 (N_35591,N_35204,N_35053);
and U35592 (N_35592,N_35100,N_35059);
nand U35593 (N_35593,N_35136,N_35310);
nand U35594 (N_35594,N_35291,N_35359);
and U35595 (N_35595,N_35157,N_35147);
nand U35596 (N_35596,N_35004,N_35303);
nor U35597 (N_35597,N_35140,N_35080);
or U35598 (N_35598,N_35453,N_35135);
xor U35599 (N_35599,N_35043,N_35071);
nor U35600 (N_35600,N_35161,N_35196);
or U35601 (N_35601,N_35028,N_35160);
nand U35602 (N_35602,N_35452,N_35200);
or U35603 (N_35603,N_35241,N_35313);
nand U35604 (N_35604,N_35232,N_35137);
or U35605 (N_35605,N_35054,N_35174);
and U35606 (N_35606,N_35332,N_35198);
nor U35607 (N_35607,N_35218,N_35353);
nand U35608 (N_35608,N_35495,N_35014);
or U35609 (N_35609,N_35223,N_35007);
nand U35610 (N_35610,N_35421,N_35042);
or U35611 (N_35611,N_35120,N_35274);
nand U35612 (N_35612,N_35491,N_35061);
xnor U35613 (N_35613,N_35289,N_35346);
nor U35614 (N_35614,N_35273,N_35186);
xor U35615 (N_35615,N_35284,N_35396);
and U35616 (N_35616,N_35206,N_35075);
nor U35617 (N_35617,N_35394,N_35247);
xnor U35618 (N_35618,N_35257,N_35485);
xor U35619 (N_35619,N_35121,N_35366);
or U35620 (N_35620,N_35251,N_35314);
nor U35621 (N_35621,N_35000,N_35416);
nor U35622 (N_35622,N_35097,N_35133);
and U35623 (N_35623,N_35311,N_35434);
xor U35624 (N_35624,N_35407,N_35081);
and U35625 (N_35625,N_35413,N_35119);
xor U35626 (N_35626,N_35146,N_35111);
nand U35627 (N_35627,N_35162,N_35150);
nand U35628 (N_35628,N_35245,N_35220);
or U35629 (N_35629,N_35304,N_35320);
and U35630 (N_35630,N_35318,N_35006);
nand U35631 (N_35631,N_35055,N_35039);
nor U35632 (N_35632,N_35494,N_35029);
or U35633 (N_35633,N_35144,N_35030);
and U35634 (N_35634,N_35464,N_35462);
xor U35635 (N_35635,N_35044,N_35265);
or U35636 (N_35636,N_35387,N_35122);
and U35637 (N_35637,N_35222,N_35330);
or U35638 (N_35638,N_35463,N_35020);
nand U35639 (N_35639,N_35397,N_35472);
nor U35640 (N_35640,N_35278,N_35456);
nor U35641 (N_35641,N_35440,N_35447);
and U35642 (N_35642,N_35143,N_35013);
xor U35643 (N_35643,N_35465,N_35286);
nor U35644 (N_35644,N_35236,N_35110);
nor U35645 (N_35645,N_35182,N_35213);
nand U35646 (N_35646,N_35128,N_35064);
or U35647 (N_35647,N_35297,N_35326);
nand U35648 (N_35648,N_35224,N_35215);
xor U35649 (N_35649,N_35329,N_35262);
and U35650 (N_35650,N_35194,N_35388);
nand U35651 (N_35651,N_35370,N_35355);
or U35652 (N_35652,N_35017,N_35468);
nand U35653 (N_35653,N_35312,N_35458);
nand U35654 (N_35654,N_35225,N_35352);
nor U35655 (N_35655,N_35309,N_35356);
nor U35656 (N_35656,N_35410,N_35360);
xnor U35657 (N_35657,N_35282,N_35446);
or U35658 (N_35658,N_35065,N_35420);
nor U35659 (N_35659,N_35322,N_35172);
nor U35660 (N_35660,N_35400,N_35338);
or U35661 (N_35661,N_35431,N_35003);
nor U35662 (N_35662,N_35170,N_35188);
xor U35663 (N_35663,N_35279,N_35124);
nand U35664 (N_35664,N_35492,N_35201);
xnor U35665 (N_35665,N_35367,N_35324);
nand U35666 (N_35666,N_35406,N_35448);
or U35667 (N_35667,N_35019,N_35103);
and U35668 (N_35668,N_35277,N_35068);
and U35669 (N_35669,N_35386,N_35414);
nand U35670 (N_35670,N_35454,N_35083);
nor U35671 (N_35671,N_35428,N_35117);
nor U35672 (N_35672,N_35192,N_35046);
nor U35673 (N_35673,N_35001,N_35233);
and U35674 (N_35674,N_35203,N_35317);
or U35675 (N_35675,N_35158,N_35375);
nor U35676 (N_35676,N_35382,N_35139);
xnor U35677 (N_35677,N_35012,N_35444);
nand U35678 (N_35678,N_35398,N_35368);
or U35679 (N_35679,N_35185,N_35171);
nand U35680 (N_35680,N_35022,N_35148);
nor U35681 (N_35681,N_35109,N_35116);
and U35682 (N_35682,N_35159,N_35108);
xnor U35683 (N_35683,N_35173,N_35027);
xnor U35684 (N_35684,N_35118,N_35141);
xor U35685 (N_35685,N_35305,N_35235);
or U35686 (N_35686,N_35285,N_35321);
and U35687 (N_35687,N_35466,N_35425);
nand U35688 (N_35688,N_35473,N_35469);
or U35689 (N_35689,N_35449,N_35451);
xnor U35690 (N_35690,N_35045,N_35238);
nor U35691 (N_35691,N_35096,N_35098);
xor U35692 (N_35692,N_35319,N_35031);
and U35693 (N_35693,N_35333,N_35340);
or U35694 (N_35694,N_35058,N_35296);
nor U35695 (N_35695,N_35193,N_35344);
or U35696 (N_35696,N_35149,N_35051);
nand U35697 (N_35697,N_35476,N_35381);
or U35698 (N_35698,N_35474,N_35256);
or U35699 (N_35699,N_35334,N_35377);
nand U35700 (N_35700,N_35087,N_35268);
nand U35701 (N_35701,N_35164,N_35093);
or U35702 (N_35702,N_35015,N_35484);
or U35703 (N_35703,N_35063,N_35114);
xor U35704 (N_35704,N_35165,N_35092);
or U35705 (N_35705,N_35259,N_35132);
nor U35706 (N_35706,N_35275,N_35153);
nand U35707 (N_35707,N_35328,N_35266);
nor U35708 (N_35708,N_35179,N_35167);
nand U35709 (N_35709,N_35035,N_35026);
nor U35710 (N_35710,N_35373,N_35077);
nand U35711 (N_35711,N_35074,N_35496);
and U35712 (N_35712,N_35178,N_35374);
or U35713 (N_35713,N_35339,N_35142);
or U35714 (N_35714,N_35230,N_35250);
or U35715 (N_35715,N_35056,N_35487);
nand U35716 (N_35716,N_35438,N_35079);
nand U35717 (N_35717,N_35315,N_35412);
xor U35718 (N_35718,N_35131,N_35299);
and U35719 (N_35719,N_35255,N_35308);
nor U35720 (N_35720,N_35091,N_35283);
nand U35721 (N_35721,N_35155,N_35379);
nand U35722 (N_35722,N_35460,N_35295);
xnor U35723 (N_35723,N_35393,N_35195);
nand U35724 (N_35724,N_35163,N_35085);
and U35725 (N_35725,N_35126,N_35499);
or U35726 (N_35726,N_35217,N_35402);
nor U35727 (N_35727,N_35350,N_35151);
nand U35728 (N_35728,N_35404,N_35439);
and U35729 (N_35729,N_35202,N_35008);
nor U35730 (N_35730,N_35088,N_35024);
nor U35731 (N_35731,N_35437,N_35197);
nand U35732 (N_35732,N_35411,N_35281);
nor U35733 (N_35733,N_35263,N_35156);
or U35734 (N_35734,N_35395,N_35244);
or U35735 (N_35735,N_35191,N_35102);
nor U35736 (N_35736,N_35184,N_35272);
nor U35737 (N_35737,N_35391,N_35154);
or U35738 (N_35738,N_35221,N_35166);
nand U35739 (N_35739,N_35181,N_35105);
and U35740 (N_35740,N_35234,N_35190);
nor U35741 (N_35741,N_35325,N_35418);
nand U35742 (N_35742,N_35354,N_35216);
nand U35743 (N_35743,N_35477,N_35498);
nor U35744 (N_35744,N_35187,N_35415);
xnor U35745 (N_35745,N_35033,N_35107);
nor U35746 (N_35746,N_35347,N_35287);
nand U35747 (N_35747,N_35341,N_35475);
or U35748 (N_35748,N_35253,N_35123);
xnor U35749 (N_35749,N_35357,N_35208);
nor U35750 (N_35750,N_35012,N_35424);
xnor U35751 (N_35751,N_35331,N_35111);
xor U35752 (N_35752,N_35171,N_35301);
xor U35753 (N_35753,N_35484,N_35440);
nor U35754 (N_35754,N_35009,N_35328);
nand U35755 (N_35755,N_35394,N_35480);
or U35756 (N_35756,N_35220,N_35490);
nand U35757 (N_35757,N_35313,N_35066);
or U35758 (N_35758,N_35241,N_35494);
or U35759 (N_35759,N_35097,N_35155);
nand U35760 (N_35760,N_35345,N_35370);
nor U35761 (N_35761,N_35151,N_35287);
and U35762 (N_35762,N_35076,N_35176);
xnor U35763 (N_35763,N_35114,N_35130);
nor U35764 (N_35764,N_35488,N_35423);
and U35765 (N_35765,N_35301,N_35119);
and U35766 (N_35766,N_35300,N_35100);
nor U35767 (N_35767,N_35117,N_35150);
and U35768 (N_35768,N_35260,N_35337);
nor U35769 (N_35769,N_35321,N_35231);
and U35770 (N_35770,N_35415,N_35114);
nand U35771 (N_35771,N_35011,N_35265);
or U35772 (N_35772,N_35288,N_35199);
or U35773 (N_35773,N_35006,N_35273);
nand U35774 (N_35774,N_35121,N_35436);
nor U35775 (N_35775,N_35213,N_35367);
xor U35776 (N_35776,N_35145,N_35082);
nor U35777 (N_35777,N_35340,N_35366);
or U35778 (N_35778,N_35014,N_35437);
or U35779 (N_35779,N_35417,N_35488);
and U35780 (N_35780,N_35064,N_35319);
nand U35781 (N_35781,N_35394,N_35272);
and U35782 (N_35782,N_35031,N_35266);
and U35783 (N_35783,N_35330,N_35487);
and U35784 (N_35784,N_35237,N_35352);
xnor U35785 (N_35785,N_35422,N_35432);
or U35786 (N_35786,N_35409,N_35172);
nand U35787 (N_35787,N_35161,N_35473);
nor U35788 (N_35788,N_35279,N_35058);
nand U35789 (N_35789,N_35088,N_35464);
nand U35790 (N_35790,N_35314,N_35482);
xnor U35791 (N_35791,N_35299,N_35192);
or U35792 (N_35792,N_35301,N_35278);
nor U35793 (N_35793,N_35157,N_35228);
or U35794 (N_35794,N_35400,N_35156);
nand U35795 (N_35795,N_35470,N_35242);
nand U35796 (N_35796,N_35114,N_35450);
nand U35797 (N_35797,N_35188,N_35404);
nor U35798 (N_35798,N_35203,N_35192);
and U35799 (N_35799,N_35462,N_35175);
nor U35800 (N_35800,N_35450,N_35428);
or U35801 (N_35801,N_35257,N_35004);
and U35802 (N_35802,N_35316,N_35365);
nand U35803 (N_35803,N_35302,N_35458);
nand U35804 (N_35804,N_35440,N_35433);
xnor U35805 (N_35805,N_35443,N_35418);
and U35806 (N_35806,N_35391,N_35376);
nor U35807 (N_35807,N_35229,N_35154);
xnor U35808 (N_35808,N_35020,N_35245);
nand U35809 (N_35809,N_35020,N_35226);
or U35810 (N_35810,N_35466,N_35133);
and U35811 (N_35811,N_35025,N_35101);
xnor U35812 (N_35812,N_35021,N_35056);
nand U35813 (N_35813,N_35388,N_35461);
nand U35814 (N_35814,N_35209,N_35052);
nand U35815 (N_35815,N_35237,N_35487);
xnor U35816 (N_35816,N_35299,N_35264);
and U35817 (N_35817,N_35400,N_35461);
nand U35818 (N_35818,N_35461,N_35042);
nor U35819 (N_35819,N_35202,N_35426);
or U35820 (N_35820,N_35332,N_35383);
and U35821 (N_35821,N_35237,N_35304);
nor U35822 (N_35822,N_35474,N_35499);
nor U35823 (N_35823,N_35042,N_35310);
nor U35824 (N_35824,N_35036,N_35430);
nand U35825 (N_35825,N_35095,N_35138);
nor U35826 (N_35826,N_35409,N_35396);
and U35827 (N_35827,N_35126,N_35111);
xnor U35828 (N_35828,N_35160,N_35296);
nor U35829 (N_35829,N_35471,N_35221);
nand U35830 (N_35830,N_35183,N_35344);
xnor U35831 (N_35831,N_35326,N_35414);
nand U35832 (N_35832,N_35387,N_35055);
xor U35833 (N_35833,N_35137,N_35023);
nand U35834 (N_35834,N_35009,N_35330);
xnor U35835 (N_35835,N_35435,N_35469);
and U35836 (N_35836,N_35309,N_35277);
nor U35837 (N_35837,N_35220,N_35385);
and U35838 (N_35838,N_35358,N_35084);
nor U35839 (N_35839,N_35335,N_35329);
xnor U35840 (N_35840,N_35113,N_35230);
and U35841 (N_35841,N_35376,N_35364);
nor U35842 (N_35842,N_35120,N_35412);
and U35843 (N_35843,N_35113,N_35186);
nand U35844 (N_35844,N_35480,N_35418);
and U35845 (N_35845,N_35454,N_35087);
xor U35846 (N_35846,N_35463,N_35129);
and U35847 (N_35847,N_35232,N_35399);
nor U35848 (N_35848,N_35143,N_35083);
nand U35849 (N_35849,N_35333,N_35327);
nand U35850 (N_35850,N_35455,N_35363);
nor U35851 (N_35851,N_35170,N_35016);
nor U35852 (N_35852,N_35426,N_35019);
or U35853 (N_35853,N_35092,N_35005);
xor U35854 (N_35854,N_35351,N_35220);
or U35855 (N_35855,N_35109,N_35073);
nor U35856 (N_35856,N_35277,N_35097);
nor U35857 (N_35857,N_35145,N_35476);
nor U35858 (N_35858,N_35377,N_35141);
and U35859 (N_35859,N_35173,N_35113);
nand U35860 (N_35860,N_35499,N_35264);
or U35861 (N_35861,N_35014,N_35223);
xnor U35862 (N_35862,N_35037,N_35080);
nor U35863 (N_35863,N_35170,N_35077);
or U35864 (N_35864,N_35023,N_35255);
xnor U35865 (N_35865,N_35435,N_35329);
or U35866 (N_35866,N_35231,N_35218);
or U35867 (N_35867,N_35417,N_35212);
or U35868 (N_35868,N_35279,N_35346);
nor U35869 (N_35869,N_35096,N_35318);
or U35870 (N_35870,N_35217,N_35188);
nor U35871 (N_35871,N_35148,N_35174);
and U35872 (N_35872,N_35197,N_35091);
nor U35873 (N_35873,N_35232,N_35489);
nand U35874 (N_35874,N_35135,N_35156);
or U35875 (N_35875,N_35061,N_35225);
xor U35876 (N_35876,N_35107,N_35318);
nand U35877 (N_35877,N_35052,N_35227);
xor U35878 (N_35878,N_35018,N_35355);
xor U35879 (N_35879,N_35187,N_35129);
or U35880 (N_35880,N_35136,N_35224);
or U35881 (N_35881,N_35007,N_35417);
nand U35882 (N_35882,N_35424,N_35283);
and U35883 (N_35883,N_35268,N_35219);
nor U35884 (N_35884,N_35487,N_35047);
and U35885 (N_35885,N_35060,N_35425);
xnor U35886 (N_35886,N_35429,N_35121);
or U35887 (N_35887,N_35343,N_35312);
and U35888 (N_35888,N_35021,N_35415);
nor U35889 (N_35889,N_35324,N_35027);
or U35890 (N_35890,N_35082,N_35201);
or U35891 (N_35891,N_35095,N_35129);
nor U35892 (N_35892,N_35053,N_35005);
xor U35893 (N_35893,N_35298,N_35415);
or U35894 (N_35894,N_35348,N_35470);
and U35895 (N_35895,N_35358,N_35367);
nand U35896 (N_35896,N_35495,N_35265);
or U35897 (N_35897,N_35137,N_35469);
xor U35898 (N_35898,N_35447,N_35226);
nand U35899 (N_35899,N_35438,N_35078);
and U35900 (N_35900,N_35275,N_35456);
nand U35901 (N_35901,N_35107,N_35100);
or U35902 (N_35902,N_35244,N_35128);
and U35903 (N_35903,N_35027,N_35002);
or U35904 (N_35904,N_35456,N_35008);
nand U35905 (N_35905,N_35398,N_35452);
or U35906 (N_35906,N_35468,N_35431);
nor U35907 (N_35907,N_35379,N_35182);
xor U35908 (N_35908,N_35201,N_35179);
xor U35909 (N_35909,N_35039,N_35111);
and U35910 (N_35910,N_35167,N_35481);
nor U35911 (N_35911,N_35284,N_35225);
nor U35912 (N_35912,N_35125,N_35117);
and U35913 (N_35913,N_35190,N_35498);
nor U35914 (N_35914,N_35010,N_35374);
xor U35915 (N_35915,N_35404,N_35402);
nor U35916 (N_35916,N_35376,N_35148);
nand U35917 (N_35917,N_35215,N_35273);
nand U35918 (N_35918,N_35274,N_35154);
and U35919 (N_35919,N_35309,N_35379);
or U35920 (N_35920,N_35086,N_35162);
or U35921 (N_35921,N_35168,N_35175);
nor U35922 (N_35922,N_35147,N_35356);
xnor U35923 (N_35923,N_35234,N_35130);
nand U35924 (N_35924,N_35251,N_35264);
or U35925 (N_35925,N_35414,N_35106);
nor U35926 (N_35926,N_35137,N_35178);
xor U35927 (N_35927,N_35186,N_35240);
xnor U35928 (N_35928,N_35147,N_35085);
nand U35929 (N_35929,N_35474,N_35007);
nor U35930 (N_35930,N_35087,N_35448);
and U35931 (N_35931,N_35429,N_35227);
nor U35932 (N_35932,N_35153,N_35026);
or U35933 (N_35933,N_35204,N_35405);
and U35934 (N_35934,N_35317,N_35232);
or U35935 (N_35935,N_35054,N_35322);
nand U35936 (N_35936,N_35038,N_35328);
or U35937 (N_35937,N_35207,N_35048);
nand U35938 (N_35938,N_35323,N_35496);
nand U35939 (N_35939,N_35096,N_35200);
and U35940 (N_35940,N_35172,N_35085);
xnor U35941 (N_35941,N_35449,N_35078);
nand U35942 (N_35942,N_35145,N_35053);
nor U35943 (N_35943,N_35132,N_35016);
or U35944 (N_35944,N_35234,N_35136);
or U35945 (N_35945,N_35273,N_35369);
or U35946 (N_35946,N_35162,N_35437);
nor U35947 (N_35947,N_35235,N_35411);
nand U35948 (N_35948,N_35363,N_35019);
and U35949 (N_35949,N_35295,N_35150);
xor U35950 (N_35950,N_35283,N_35019);
or U35951 (N_35951,N_35134,N_35252);
nand U35952 (N_35952,N_35126,N_35228);
and U35953 (N_35953,N_35449,N_35207);
and U35954 (N_35954,N_35207,N_35019);
xor U35955 (N_35955,N_35030,N_35133);
nand U35956 (N_35956,N_35229,N_35012);
xnor U35957 (N_35957,N_35114,N_35087);
and U35958 (N_35958,N_35362,N_35357);
and U35959 (N_35959,N_35249,N_35335);
xnor U35960 (N_35960,N_35235,N_35073);
or U35961 (N_35961,N_35206,N_35031);
or U35962 (N_35962,N_35158,N_35355);
and U35963 (N_35963,N_35125,N_35390);
and U35964 (N_35964,N_35436,N_35345);
nor U35965 (N_35965,N_35348,N_35144);
nand U35966 (N_35966,N_35234,N_35000);
and U35967 (N_35967,N_35457,N_35442);
nand U35968 (N_35968,N_35433,N_35297);
xor U35969 (N_35969,N_35001,N_35241);
xnor U35970 (N_35970,N_35328,N_35432);
or U35971 (N_35971,N_35053,N_35013);
xor U35972 (N_35972,N_35249,N_35483);
xor U35973 (N_35973,N_35065,N_35107);
nand U35974 (N_35974,N_35498,N_35081);
nor U35975 (N_35975,N_35051,N_35367);
xnor U35976 (N_35976,N_35135,N_35020);
or U35977 (N_35977,N_35276,N_35287);
and U35978 (N_35978,N_35409,N_35217);
xor U35979 (N_35979,N_35427,N_35200);
and U35980 (N_35980,N_35036,N_35319);
nand U35981 (N_35981,N_35238,N_35487);
xnor U35982 (N_35982,N_35149,N_35136);
nor U35983 (N_35983,N_35194,N_35201);
or U35984 (N_35984,N_35435,N_35246);
nand U35985 (N_35985,N_35129,N_35052);
nand U35986 (N_35986,N_35048,N_35173);
or U35987 (N_35987,N_35359,N_35212);
nand U35988 (N_35988,N_35007,N_35183);
nor U35989 (N_35989,N_35099,N_35198);
xor U35990 (N_35990,N_35363,N_35016);
nor U35991 (N_35991,N_35014,N_35228);
nand U35992 (N_35992,N_35363,N_35246);
or U35993 (N_35993,N_35089,N_35487);
nand U35994 (N_35994,N_35191,N_35138);
xnor U35995 (N_35995,N_35185,N_35206);
nand U35996 (N_35996,N_35355,N_35001);
and U35997 (N_35997,N_35304,N_35384);
nor U35998 (N_35998,N_35291,N_35169);
nor U35999 (N_35999,N_35248,N_35047);
nand U36000 (N_36000,N_35572,N_35802);
or U36001 (N_36001,N_35625,N_35939);
xnor U36002 (N_36002,N_35691,N_35795);
xor U36003 (N_36003,N_35711,N_35926);
and U36004 (N_36004,N_35845,N_35879);
nor U36005 (N_36005,N_35621,N_35657);
xor U36006 (N_36006,N_35922,N_35534);
nand U36007 (N_36007,N_35761,N_35908);
and U36008 (N_36008,N_35872,N_35983);
or U36009 (N_36009,N_35703,N_35723);
or U36010 (N_36010,N_35727,N_35624);
xnor U36011 (N_36011,N_35659,N_35950);
or U36012 (N_36012,N_35611,N_35655);
xnor U36013 (N_36013,N_35885,N_35897);
nor U36014 (N_36014,N_35675,N_35893);
and U36015 (N_36015,N_35620,N_35853);
or U36016 (N_36016,N_35769,N_35840);
xor U36017 (N_36017,N_35809,N_35902);
nor U36018 (N_36018,N_35751,N_35980);
and U36019 (N_36019,N_35821,N_35735);
xor U36020 (N_36020,N_35512,N_35518);
and U36021 (N_36021,N_35959,N_35822);
and U36022 (N_36022,N_35537,N_35634);
and U36023 (N_36023,N_35758,N_35837);
xor U36024 (N_36024,N_35511,N_35865);
xor U36025 (N_36025,N_35743,N_35500);
or U36026 (N_36026,N_35869,N_35789);
nor U36027 (N_36027,N_35694,N_35906);
nand U36028 (N_36028,N_35875,N_35506);
and U36029 (N_36029,N_35776,N_35683);
and U36030 (N_36030,N_35808,N_35843);
and U36031 (N_36031,N_35766,N_35686);
nor U36032 (N_36032,N_35828,N_35589);
nor U36033 (N_36033,N_35839,N_35651);
or U36034 (N_36034,N_35575,N_35842);
nor U36035 (N_36035,N_35979,N_35787);
and U36036 (N_36036,N_35904,N_35600);
nand U36037 (N_36037,N_35641,N_35924);
nand U36038 (N_36038,N_35891,N_35985);
xnor U36039 (N_36039,N_35756,N_35971);
nor U36040 (N_36040,N_35870,N_35955);
nand U36041 (N_36041,N_35501,N_35586);
xor U36042 (N_36042,N_35672,N_35811);
nor U36043 (N_36043,N_35567,N_35504);
or U36044 (N_36044,N_35740,N_35833);
nor U36045 (N_36045,N_35656,N_35606);
xor U36046 (N_36046,N_35949,N_35945);
and U36047 (N_36047,N_35946,N_35584);
xnor U36048 (N_36048,N_35529,N_35526);
and U36049 (N_36049,N_35903,N_35782);
and U36050 (N_36050,N_35911,N_35996);
nor U36051 (N_36051,N_35825,N_35707);
nand U36052 (N_36052,N_35610,N_35977);
nand U36053 (N_36053,N_35615,N_35684);
nor U36054 (N_36054,N_35889,N_35576);
xnor U36055 (N_36055,N_35588,N_35692);
nor U36056 (N_36056,N_35849,N_35535);
xnor U36057 (N_36057,N_35944,N_35559);
and U36058 (N_36058,N_35565,N_35665);
nand U36059 (N_36059,N_35682,N_35724);
nor U36060 (N_36060,N_35791,N_35508);
or U36061 (N_36061,N_35868,N_35856);
nand U36062 (N_36062,N_35716,N_35813);
nand U36063 (N_36063,N_35984,N_35585);
nand U36064 (N_36064,N_35550,N_35798);
nor U36065 (N_36065,N_35951,N_35750);
nor U36066 (N_36066,N_35744,N_35725);
nand U36067 (N_36067,N_35763,N_35919);
nor U36068 (N_36068,N_35706,N_35834);
xor U36069 (N_36069,N_35638,N_35661);
or U36070 (N_36070,N_35779,N_35505);
nor U36071 (N_36071,N_35730,N_35598);
or U36072 (N_36072,N_35548,N_35967);
or U36073 (N_36073,N_35732,N_35729);
xor U36074 (N_36074,N_35829,N_35742);
or U36075 (N_36075,N_35536,N_35639);
nor U36076 (N_36076,N_35649,N_35807);
xor U36077 (N_36077,N_35749,N_35583);
or U36078 (N_36078,N_35622,N_35545);
xor U36079 (N_36079,N_35876,N_35764);
nand U36080 (N_36080,N_35835,N_35823);
and U36081 (N_36081,N_35687,N_35998);
or U36082 (N_36082,N_35516,N_35737);
nand U36083 (N_36083,N_35883,N_35805);
nor U36084 (N_36084,N_35513,N_35633);
nand U36085 (N_36085,N_35968,N_35914);
nand U36086 (N_36086,N_35595,N_35558);
and U36087 (N_36087,N_35754,N_35982);
xor U36088 (N_36088,N_35676,N_35580);
and U36089 (N_36089,N_35770,N_35830);
or U36090 (N_36090,N_35817,N_35803);
and U36091 (N_36091,N_35969,N_35590);
and U36092 (N_36092,N_35881,N_35826);
nor U36093 (N_36093,N_35895,N_35582);
and U36094 (N_36094,N_35591,N_35918);
or U36095 (N_36095,N_35970,N_35768);
and U36096 (N_36096,N_35635,N_35820);
or U36097 (N_36097,N_35520,N_35522);
or U36098 (N_36098,N_35755,N_35936);
and U36099 (N_36099,N_35816,N_35882);
nor U36100 (N_36100,N_35748,N_35562);
xor U36101 (N_36101,N_35556,N_35757);
and U36102 (N_36102,N_35940,N_35960);
nand U36103 (N_36103,N_35767,N_35510);
and U36104 (N_36104,N_35759,N_35861);
and U36105 (N_36105,N_35608,N_35566);
nor U36106 (N_36106,N_35571,N_35896);
or U36107 (N_36107,N_35943,N_35956);
or U36108 (N_36108,N_35988,N_35653);
nand U36109 (N_36109,N_35827,N_35547);
nor U36110 (N_36110,N_35728,N_35643);
and U36111 (N_36111,N_35652,N_35991);
nor U36112 (N_36112,N_35752,N_35549);
xnor U36113 (N_36113,N_35577,N_35775);
or U36114 (N_36114,N_35890,N_35555);
nor U36115 (N_36115,N_35804,N_35831);
and U36116 (N_36116,N_35715,N_35542);
or U36117 (N_36117,N_35987,N_35973);
xor U36118 (N_36118,N_35954,N_35507);
nand U36119 (N_36119,N_35797,N_35910);
xnor U36120 (N_36120,N_35958,N_35877);
nand U36121 (N_36121,N_35931,N_35667);
nor U36122 (N_36122,N_35544,N_35688);
or U36123 (N_36123,N_35640,N_35601);
nand U36124 (N_36124,N_35623,N_35947);
xor U36125 (N_36125,N_35602,N_35539);
or U36126 (N_36126,N_35783,N_35609);
or U36127 (N_36127,N_35630,N_35898);
xor U36128 (N_36128,N_35697,N_35690);
or U36129 (N_36129,N_35866,N_35731);
and U36130 (N_36130,N_35760,N_35632);
and U36131 (N_36131,N_35670,N_35777);
nand U36132 (N_36132,N_35614,N_35972);
nor U36133 (N_36133,N_35934,N_35886);
nand U36134 (N_36134,N_35878,N_35525);
nand U36135 (N_36135,N_35978,N_35531);
xor U36136 (N_36136,N_35645,N_35784);
nand U36137 (N_36137,N_35712,N_35654);
or U36138 (N_36138,N_35709,N_35514);
or U36139 (N_36139,N_35663,N_35855);
or U36140 (N_36140,N_35933,N_35923);
nand U36141 (N_36141,N_35738,N_35894);
and U36142 (N_36142,N_35552,N_35810);
nor U36143 (N_36143,N_35648,N_35509);
and U36144 (N_36144,N_35819,N_35741);
xor U36145 (N_36145,N_35674,N_35786);
and U36146 (N_36146,N_35981,N_35921);
xor U36147 (N_36147,N_35992,N_35700);
xnor U36148 (N_36148,N_35907,N_35852);
and U36149 (N_36149,N_35905,N_35658);
xor U36150 (N_36150,N_35540,N_35935);
nor U36151 (N_36151,N_35938,N_35965);
xnor U36152 (N_36152,N_35989,N_35929);
and U36153 (N_36153,N_35720,N_35515);
nand U36154 (N_36154,N_35568,N_35806);
nand U36155 (N_36155,N_35796,N_35762);
and U36156 (N_36156,N_35530,N_35719);
or U36157 (N_36157,N_35662,N_35551);
or U36158 (N_36158,N_35746,N_35909);
and U36159 (N_36159,N_35773,N_35613);
nand U36160 (N_36160,N_35524,N_35689);
and U36161 (N_36161,N_35772,N_35618);
xor U36162 (N_36162,N_35859,N_35747);
or U36163 (N_36163,N_35696,N_35519);
xnor U36164 (N_36164,N_35592,N_35581);
nor U36165 (N_36165,N_35814,N_35527);
nor U36166 (N_36166,N_35650,N_35563);
nor U36167 (N_36167,N_35644,N_35607);
or U36168 (N_36168,N_35887,N_35781);
or U36169 (N_36169,N_35569,N_35948);
xnor U36170 (N_36170,N_35528,N_35593);
xnor U36171 (N_36171,N_35597,N_35701);
or U36172 (N_36172,N_35617,N_35966);
xor U36173 (N_36173,N_35850,N_35863);
and U36174 (N_36174,N_35847,N_35541);
or U36175 (N_36175,N_35708,N_35841);
or U36176 (N_36176,N_35864,N_35993);
xor U36177 (N_36177,N_35668,N_35680);
xor U36178 (N_36178,N_35642,N_35564);
xnor U36179 (N_36179,N_35932,N_35873);
xor U36180 (N_36180,N_35986,N_35521);
and U36181 (N_36181,N_35631,N_35874);
xor U36182 (N_36182,N_35599,N_35626);
or U36183 (N_36183,N_35884,N_35812);
nand U36184 (N_36184,N_35553,N_35937);
nor U36185 (N_36185,N_35554,N_35628);
nor U36186 (N_36186,N_35818,N_35961);
nor U36187 (N_36187,N_35900,N_35836);
xor U36188 (N_36188,N_35533,N_35679);
xnor U36189 (N_36189,N_35677,N_35920);
and U36190 (N_36190,N_35953,N_35603);
and U36191 (N_36191,N_35523,N_35627);
nor U36192 (N_36192,N_35976,N_35942);
xor U36193 (N_36193,N_35718,N_35578);
or U36194 (N_36194,N_35546,N_35774);
nand U36195 (N_36195,N_35792,N_35780);
nor U36196 (N_36196,N_35928,N_35517);
xor U36197 (N_36197,N_35801,N_35671);
nand U36198 (N_36198,N_35815,N_35605);
or U36199 (N_36199,N_35846,N_35994);
nor U36200 (N_36200,N_35794,N_35778);
nand U36201 (N_36201,N_35713,N_35594);
or U36202 (N_36202,N_35532,N_35733);
nand U36203 (N_36203,N_35666,N_35587);
nor U36204 (N_36204,N_35739,N_35579);
or U36205 (N_36205,N_35899,N_35570);
nor U36206 (N_36206,N_35800,N_35699);
or U36207 (N_36207,N_35880,N_35721);
and U36208 (N_36208,N_35636,N_35862);
xor U36209 (N_36209,N_35913,N_35619);
nor U36210 (N_36210,N_35765,N_35503);
nand U36211 (N_36211,N_35596,N_35616);
or U36212 (N_36212,N_35785,N_35705);
nand U36213 (N_36213,N_35664,N_35573);
or U36214 (N_36214,N_35927,N_35975);
nor U36215 (N_36215,N_35832,N_35952);
nor U36216 (N_36216,N_35858,N_35901);
xnor U36217 (N_36217,N_35854,N_35646);
and U36218 (N_36218,N_35963,N_35685);
and U36219 (N_36219,N_35717,N_35925);
and U36220 (N_36220,N_35647,N_35793);
nand U36221 (N_36221,N_35612,N_35714);
and U36222 (N_36222,N_35726,N_35790);
nor U36223 (N_36223,N_35710,N_35844);
nor U36224 (N_36224,N_35912,N_35736);
and U36225 (N_36225,N_35941,N_35990);
and U36226 (N_36226,N_35824,N_35848);
or U36227 (N_36227,N_35860,N_35574);
or U36228 (N_36228,N_35857,N_35930);
nor U36229 (N_36229,N_35867,N_35734);
or U36230 (N_36230,N_35915,N_35695);
nor U36231 (N_36231,N_35704,N_35788);
or U36232 (N_36232,N_35678,N_35722);
nor U36233 (N_36233,N_35502,N_35557);
and U36234 (N_36234,N_35693,N_35957);
and U36235 (N_36235,N_35838,N_35892);
nor U36236 (N_36236,N_35771,N_35962);
xor U36237 (N_36237,N_35995,N_35698);
xnor U36238 (N_36238,N_35745,N_35702);
nand U36239 (N_36239,N_35917,N_35629);
or U36240 (N_36240,N_35637,N_35974);
nand U36241 (N_36241,N_35561,N_35999);
xnor U36242 (N_36242,N_35753,N_35964);
and U36243 (N_36243,N_35538,N_35673);
or U36244 (N_36244,N_35604,N_35660);
nand U36245 (N_36245,N_35560,N_35871);
and U36246 (N_36246,N_35669,N_35681);
nand U36247 (N_36247,N_35543,N_35799);
xor U36248 (N_36248,N_35916,N_35888);
or U36249 (N_36249,N_35851,N_35997);
xnor U36250 (N_36250,N_35621,N_35774);
and U36251 (N_36251,N_35580,N_35825);
nand U36252 (N_36252,N_35678,N_35535);
and U36253 (N_36253,N_35954,N_35591);
and U36254 (N_36254,N_35618,N_35855);
xor U36255 (N_36255,N_35617,N_35510);
nor U36256 (N_36256,N_35735,N_35873);
xnor U36257 (N_36257,N_35745,N_35869);
xor U36258 (N_36258,N_35760,N_35527);
and U36259 (N_36259,N_35985,N_35719);
nand U36260 (N_36260,N_35596,N_35708);
nor U36261 (N_36261,N_35889,N_35935);
and U36262 (N_36262,N_35949,N_35533);
or U36263 (N_36263,N_35821,N_35922);
nand U36264 (N_36264,N_35686,N_35903);
or U36265 (N_36265,N_35646,N_35556);
xnor U36266 (N_36266,N_35708,N_35511);
or U36267 (N_36267,N_35871,N_35872);
nor U36268 (N_36268,N_35560,N_35504);
or U36269 (N_36269,N_35813,N_35671);
nand U36270 (N_36270,N_35592,N_35886);
or U36271 (N_36271,N_35888,N_35557);
xor U36272 (N_36272,N_35513,N_35934);
or U36273 (N_36273,N_35970,N_35910);
nand U36274 (N_36274,N_35827,N_35900);
and U36275 (N_36275,N_35997,N_35918);
and U36276 (N_36276,N_35909,N_35832);
or U36277 (N_36277,N_35577,N_35505);
xor U36278 (N_36278,N_35555,N_35614);
nor U36279 (N_36279,N_35574,N_35920);
xor U36280 (N_36280,N_35941,N_35621);
nor U36281 (N_36281,N_35957,N_35701);
nand U36282 (N_36282,N_35683,N_35729);
nand U36283 (N_36283,N_35893,N_35929);
xnor U36284 (N_36284,N_35680,N_35822);
nand U36285 (N_36285,N_35809,N_35634);
or U36286 (N_36286,N_35770,N_35926);
or U36287 (N_36287,N_35568,N_35655);
nand U36288 (N_36288,N_35564,N_35853);
nand U36289 (N_36289,N_35949,N_35767);
and U36290 (N_36290,N_35774,N_35754);
nand U36291 (N_36291,N_35738,N_35720);
or U36292 (N_36292,N_35726,N_35566);
nor U36293 (N_36293,N_35940,N_35985);
nor U36294 (N_36294,N_35818,N_35520);
xnor U36295 (N_36295,N_35970,N_35715);
nand U36296 (N_36296,N_35760,N_35973);
or U36297 (N_36297,N_35638,N_35957);
xnor U36298 (N_36298,N_35844,N_35824);
nand U36299 (N_36299,N_35945,N_35932);
nand U36300 (N_36300,N_35794,N_35677);
nand U36301 (N_36301,N_35914,N_35588);
nand U36302 (N_36302,N_35891,N_35524);
nor U36303 (N_36303,N_35594,N_35579);
or U36304 (N_36304,N_35830,N_35746);
xnor U36305 (N_36305,N_35747,N_35584);
nand U36306 (N_36306,N_35541,N_35543);
or U36307 (N_36307,N_35589,N_35669);
and U36308 (N_36308,N_35616,N_35831);
or U36309 (N_36309,N_35532,N_35584);
nor U36310 (N_36310,N_35581,N_35670);
nand U36311 (N_36311,N_35739,N_35998);
nor U36312 (N_36312,N_35892,N_35688);
nor U36313 (N_36313,N_35828,N_35658);
or U36314 (N_36314,N_35578,N_35930);
nand U36315 (N_36315,N_35865,N_35896);
nor U36316 (N_36316,N_35951,N_35788);
or U36317 (N_36317,N_35575,N_35945);
nor U36318 (N_36318,N_35790,N_35534);
or U36319 (N_36319,N_35976,N_35698);
and U36320 (N_36320,N_35587,N_35902);
or U36321 (N_36321,N_35513,N_35719);
xor U36322 (N_36322,N_35544,N_35805);
nand U36323 (N_36323,N_35644,N_35726);
nor U36324 (N_36324,N_35505,N_35582);
nand U36325 (N_36325,N_35596,N_35799);
nand U36326 (N_36326,N_35633,N_35514);
and U36327 (N_36327,N_35575,N_35775);
nor U36328 (N_36328,N_35591,N_35658);
xnor U36329 (N_36329,N_35835,N_35830);
and U36330 (N_36330,N_35890,N_35501);
nor U36331 (N_36331,N_35910,N_35730);
and U36332 (N_36332,N_35551,N_35931);
and U36333 (N_36333,N_35516,N_35537);
or U36334 (N_36334,N_35984,N_35587);
nor U36335 (N_36335,N_35510,N_35521);
and U36336 (N_36336,N_35682,N_35809);
nor U36337 (N_36337,N_35668,N_35621);
xnor U36338 (N_36338,N_35763,N_35564);
xnor U36339 (N_36339,N_35736,N_35962);
or U36340 (N_36340,N_35930,N_35746);
and U36341 (N_36341,N_35548,N_35793);
nand U36342 (N_36342,N_35803,N_35581);
and U36343 (N_36343,N_35594,N_35831);
nand U36344 (N_36344,N_35685,N_35634);
nor U36345 (N_36345,N_35502,N_35874);
nor U36346 (N_36346,N_35533,N_35662);
xor U36347 (N_36347,N_35786,N_35781);
xor U36348 (N_36348,N_35831,N_35588);
xor U36349 (N_36349,N_35675,N_35865);
nor U36350 (N_36350,N_35690,N_35819);
nor U36351 (N_36351,N_35901,N_35848);
nor U36352 (N_36352,N_35575,N_35814);
nor U36353 (N_36353,N_35880,N_35662);
nand U36354 (N_36354,N_35836,N_35671);
nor U36355 (N_36355,N_35902,N_35741);
and U36356 (N_36356,N_35649,N_35993);
nand U36357 (N_36357,N_35778,N_35721);
nand U36358 (N_36358,N_35687,N_35585);
nand U36359 (N_36359,N_35607,N_35892);
xor U36360 (N_36360,N_35629,N_35870);
and U36361 (N_36361,N_35995,N_35878);
nand U36362 (N_36362,N_35907,N_35991);
and U36363 (N_36363,N_35853,N_35872);
nor U36364 (N_36364,N_35559,N_35837);
nor U36365 (N_36365,N_35794,N_35841);
and U36366 (N_36366,N_35556,N_35625);
xnor U36367 (N_36367,N_35763,N_35591);
nand U36368 (N_36368,N_35653,N_35686);
xnor U36369 (N_36369,N_35635,N_35813);
and U36370 (N_36370,N_35848,N_35789);
xnor U36371 (N_36371,N_35954,N_35733);
or U36372 (N_36372,N_35739,N_35542);
nand U36373 (N_36373,N_35881,N_35934);
nor U36374 (N_36374,N_35657,N_35909);
or U36375 (N_36375,N_35817,N_35512);
nor U36376 (N_36376,N_35988,N_35896);
and U36377 (N_36377,N_35661,N_35789);
or U36378 (N_36378,N_35875,N_35518);
or U36379 (N_36379,N_35932,N_35652);
and U36380 (N_36380,N_35798,N_35942);
nor U36381 (N_36381,N_35714,N_35809);
xnor U36382 (N_36382,N_35835,N_35718);
or U36383 (N_36383,N_35671,N_35895);
nand U36384 (N_36384,N_35748,N_35842);
or U36385 (N_36385,N_35529,N_35621);
xor U36386 (N_36386,N_35811,N_35557);
xnor U36387 (N_36387,N_35866,N_35536);
nor U36388 (N_36388,N_35564,N_35765);
nor U36389 (N_36389,N_35548,N_35997);
or U36390 (N_36390,N_35592,N_35503);
nor U36391 (N_36391,N_35956,N_35994);
nor U36392 (N_36392,N_35593,N_35983);
or U36393 (N_36393,N_35838,N_35563);
and U36394 (N_36394,N_35535,N_35614);
xor U36395 (N_36395,N_35528,N_35679);
xnor U36396 (N_36396,N_35750,N_35577);
nand U36397 (N_36397,N_35786,N_35749);
and U36398 (N_36398,N_35576,N_35766);
xor U36399 (N_36399,N_35950,N_35965);
nor U36400 (N_36400,N_35549,N_35868);
nand U36401 (N_36401,N_35623,N_35789);
nand U36402 (N_36402,N_35743,N_35951);
xor U36403 (N_36403,N_35838,N_35861);
xor U36404 (N_36404,N_35729,N_35902);
or U36405 (N_36405,N_35937,N_35860);
or U36406 (N_36406,N_35535,N_35945);
nor U36407 (N_36407,N_35518,N_35511);
xnor U36408 (N_36408,N_35805,N_35602);
nor U36409 (N_36409,N_35785,N_35816);
nand U36410 (N_36410,N_35808,N_35738);
or U36411 (N_36411,N_35930,N_35795);
xor U36412 (N_36412,N_35584,N_35536);
or U36413 (N_36413,N_35750,N_35934);
nand U36414 (N_36414,N_35808,N_35693);
and U36415 (N_36415,N_35955,N_35927);
or U36416 (N_36416,N_35504,N_35653);
xnor U36417 (N_36417,N_35919,N_35706);
nor U36418 (N_36418,N_35510,N_35861);
nor U36419 (N_36419,N_35818,N_35617);
or U36420 (N_36420,N_35746,N_35675);
or U36421 (N_36421,N_35971,N_35833);
nor U36422 (N_36422,N_35840,N_35678);
nor U36423 (N_36423,N_35559,N_35957);
nand U36424 (N_36424,N_35766,N_35921);
nor U36425 (N_36425,N_35791,N_35641);
xor U36426 (N_36426,N_35661,N_35971);
or U36427 (N_36427,N_35720,N_35683);
or U36428 (N_36428,N_35801,N_35546);
nand U36429 (N_36429,N_35556,N_35585);
nor U36430 (N_36430,N_35807,N_35740);
xor U36431 (N_36431,N_35817,N_35881);
nand U36432 (N_36432,N_35835,N_35715);
nand U36433 (N_36433,N_35946,N_35987);
xnor U36434 (N_36434,N_35604,N_35608);
nor U36435 (N_36435,N_35692,N_35615);
and U36436 (N_36436,N_35645,N_35788);
nand U36437 (N_36437,N_35542,N_35886);
and U36438 (N_36438,N_35505,N_35554);
xnor U36439 (N_36439,N_35895,N_35958);
nand U36440 (N_36440,N_35788,N_35830);
nor U36441 (N_36441,N_35865,N_35539);
or U36442 (N_36442,N_35645,N_35527);
nand U36443 (N_36443,N_35723,N_35522);
nand U36444 (N_36444,N_35856,N_35989);
nor U36445 (N_36445,N_35899,N_35940);
nand U36446 (N_36446,N_35774,N_35853);
xnor U36447 (N_36447,N_35609,N_35545);
nor U36448 (N_36448,N_35551,N_35916);
nand U36449 (N_36449,N_35651,N_35632);
or U36450 (N_36450,N_35696,N_35927);
nand U36451 (N_36451,N_35875,N_35725);
xnor U36452 (N_36452,N_35728,N_35703);
nor U36453 (N_36453,N_35847,N_35808);
or U36454 (N_36454,N_35918,N_35786);
nand U36455 (N_36455,N_35567,N_35832);
nand U36456 (N_36456,N_35967,N_35853);
nand U36457 (N_36457,N_35564,N_35902);
or U36458 (N_36458,N_35763,N_35991);
or U36459 (N_36459,N_35746,N_35925);
xor U36460 (N_36460,N_35670,N_35977);
and U36461 (N_36461,N_35676,N_35842);
nor U36462 (N_36462,N_35797,N_35793);
and U36463 (N_36463,N_35817,N_35990);
xnor U36464 (N_36464,N_35810,N_35539);
nor U36465 (N_36465,N_35670,N_35953);
or U36466 (N_36466,N_35755,N_35745);
xor U36467 (N_36467,N_35706,N_35841);
and U36468 (N_36468,N_35991,N_35540);
xnor U36469 (N_36469,N_35792,N_35778);
or U36470 (N_36470,N_35691,N_35577);
nand U36471 (N_36471,N_35549,N_35935);
nor U36472 (N_36472,N_35932,N_35924);
and U36473 (N_36473,N_35680,N_35518);
nor U36474 (N_36474,N_35922,N_35880);
or U36475 (N_36475,N_35956,N_35675);
or U36476 (N_36476,N_35833,N_35546);
or U36477 (N_36477,N_35651,N_35603);
or U36478 (N_36478,N_35934,N_35656);
and U36479 (N_36479,N_35676,N_35763);
or U36480 (N_36480,N_35830,N_35530);
and U36481 (N_36481,N_35768,N_35950);
or U36482 (N_36482,N_35914,N_35731);
or U36483 (N_36483,N_35781,N_35952);
nand U36484 (N_36484,N_35834,N_35576);
or U36485 (N_36485,N_35742,N_35618);
or U36486 (N_36486,N_35644,N_35582);
xnor U36487 (N_36487,N_35596,N_35726);
xor U36488 (N_36488,N_35859,N_35806);
and U36489 (N_36489,N_35880,N_35590);
nand U36490 (N_36490,N_35800,N_35966);
nand U36491 (N_36491,N_35774,N_35955);
nor U36492 (N_36492,N_35795,N_35556);
nor U36493 (N_36493,N_35965,N_35995);
and U36494 (N_36494,N_35693,N_35603);
or U36495 (N_36495,N_35797,N_35723);
and U36496 (N_36496,N_35810,N_35986);
and U36497 (N_36497,N_35598,N_35873);
nand U36498 (N_36498,N_35683,N_35886);
nand U36499 (N_36499,N_35728,N_35961);
or U36500 (N_36500,N_36257,N_36294);
nand U36501 (N_36501,N_36400,N_36494);
and U36502 (N_36502,N_36442,N_36134);
and U36503 (N_36503,N_36077,N_36487);
and U36504 (N_36504,N_36206,N_36379);
nand U36505 (N_36505,N_36407,N_36090);
xor U36506 (N_36506,N_36410,N_36075);
nor U36507 (N_36507,N_36318,N_36251);
xnor U36508 (N_36508,N_36271,N_36327);
and U36509 (N_36509,N_36029,N_36338);
xor U36510 (N_36510,N_36373,N_36030);
nor U36511 (N_36511,N_36475,N_36466);
nand U36512 (N_36512,N_36478,N_36167);
xnor U36513 (N_36513,N_36147,N_36136);
or U36514 (N_36514,N_36279,N_36272);
or U36515 (N_36515,N_36158,N_36057);
nand U36516 (N_36516,N_36237,N_36320);
nor U36517 (N_36517,N_36114,N_36286);
nand U36518 (N_36518,N_36469,N_36086);
xnor U36519 (N_36519,N_36311,N_36062);
xor U36520 (N_36520,N_36094,N_36346);
and U36521 (N_36521,N_36002,N_36281);
nor U36522 (N_36522,N_36342,N_36103);
nor U36523 (N_36523,N_36026,N_36138);
nor U36524 (N_36524,N_36078,N_36444);
or U36525 (N_36525,N_36378,N_36447);
nor U36526 (N_36526,N_36126,N_36383);
xnor U36527 (N_36527,N_36421,N_36170);
or U36528 (N_36528,N_36081,N_36244);
or U36529 (N_36529,N_36211,N_36441);
xor U36530 (N_36530,N_36052,N_36248);
xnor U36531 (N_36531,N_36402,N_36071);
or U36532 (N_36532,N_36472,N_36437);
and U36533 (N_36533,N_36193,N_36282);
xor U36534 (N_36534,N_36467,N_36474);
xnor U36535 (N_36535,N_36095,N_36384);
nand U36536 (N_36536,N_36300,N_36098);
and U36537 (N_36537,N_36491,N_36331);
nand U36538 (N_36538,N_36395,N_36048);
xnor U36539 (N_36539,N_36208,N_36406);
nor U36540 (N_36540,N_36131,N_36285);
and U36541 (N_36541,N_36425,N_36390);
xnor U36542 (N_36542,N_36083,N_36305);
and U36543 (N_36543,N_36111,N_36133);
and U36544 (N_36544,N_36012,N_36435);
xor U36545 (N_36545,N_36238,N_36429);
nor U36546 (N_36546,N_36225,N_36124);
or U36547 (N_36547,N_36356,N_36184);
and U36548 (N_36548,N_36310,N_36038);
xor U36549 (N_36549,N_36313,N_36140);
nand U36550 (N_36550,N_36016,N_36341);
or U36551 (N_36551,N_36247,N_36139);
xnor U36552 (N_36552,N_36302,N_36157);
or U36553 (N_36553,N_36269,N_36200);
nor U36554 (N_36554,N_36382,N_36243);
nor U36555 (N_36555,N_36174,N_36363);
nand U36556 (N_36556,N_36426,N_36417);
nor U36557 (N_36557,N_36047,N_36003);
xnor U36558 (N_36558,N_36185,N_36462);
and U36559 (N_36559,N_36481,N_36091);
nor U36560 (N_36560,N_36359,N_36259);
nand U36561 (N_36561,N_36013,N_36207);
or U36562 (N_36562,N_36005,N_36160);
xor U36563 (N_36563,N_36042,N_36040);
xnor U36564 (N_36564,N_36190,N_36357);
and U36565 (N_36565,N_36468,N_36431);
or U36566 (N_36566,N_36000,N_36058);
nand U36567 (N_36567,N_36056,N_36393);
nor U36568 (N_36568,N_36290,N_36037);
or U36569 (N_36569,N_36448,N_36064);
nor U36570 (N_36570,N_36369,N_36416);
and U36571 (N_36571,N_36194,N_36499);
nand U36572 (N_36572,N_36112,N_36270);
and U36573 (N_36573,N_36180,N_36216);
nand U36574 (N_36574,N_36023,N_36358);
or U36575 (N_36575,N_36186,N_36368);
and U36576 (N_36576,N_36010,N_36014);
nor U36577 (N_36577,N_36486,N_36232);
or U36578 (N_36578,N_36340,N_36477);
or U36579 (N_36579,N_36428,N_36473);
and U36580 (N_36580,N_36353,N_36376);
or U36581 (N_36581,N_36059,N_36162);
xor U36582 (N_36582,N_36122,N_36088);
and U36583 (N_36583,N_36031,N_36001);
and U36584 (N_36584,N_36315,N_36165);
xor U36585 (N_36585,N_36253,N_36490);
and U36586 (N_36586,N_36060,N_36476);
or U36587 (N_36587,N_36072,N_36325);
and U36588 (N_36588,N_36479,N_36020);
nor U36589 (N_36589,N_36236,N_36354);
nand U36590 (N_36590,N_36427,N_36398);
xor U36591 (N_36591,N_36377,N_36192);
xor U36592 (N_36592,N_36113,N_36018);
and U36593 (N_36593,N_36488,N_36181);
nor U36594 (N_36594,N_36280,N_36260);
or U36595 (N_36595,N_36433,N_36006);
nor U36596 (N_36596,N_36166,N_36388);
nand U36597 (N_36597,N_36110,N_36349);
or U36598 (N_36598,N_36204,N_36362);
and U36599 (N_36599,N_36146,N_36326);
nand U36600 (N_36600,N_36198,N_36372);
or U36601 (N_36601,N_36385,N_36132);
nand U36602 (N_36602,N_36265,N_36409);
nand U36603 (N_36603,N_36221,N_36199);
nand U36604 (N_36604,N_36153,N_36201);
nand U36605 (N_36605,N_36189,N_36322);
or U36606 (N_36606,N_36480,N_36108);
nand U36607 (N_36607,N_36035,N_36336);
nand U36608 (N_36608,N_36004,N_36415);
or U36609 (N_36609,N_36191,N_36073);
or U36610 (N_36610,N_36044,N_36309);
xnor U36611 (N_36611,N_36347,N_36404);
or U36612 (N_36612,N_36420,N_36173);
nor U36613 (N_36613,N_36032,N_36156);
and U36614 (N_36614,N_36104,N_36460);
or U36615 (N_36615,N_36394,N_36306);
xnor U36616 (N_36616,N_36154,N_36125);
nand U36617 (N_36617,N_36403,N_36128);
xnor U36618 (N_36618,N_36364,N_36025);
nor U36619 (N_36619,N_36210,N_36120);
and U36620 (N_36620,N_36145,N_36386);
xor U36621 (N_36621,N_36109,N_36449);
xor U36622 (N_36622,N_36082,N_36219);
or U36623 (N_36623,N_36275,N_36312);
or U36624 (N_36624,N_36317,N_36401);
nor U36625 (N_36625,N_36345,N_36352);
or U36626 (N_36626,N_36118,N_36350);
nand U36627 (N_36627,N_36482,N_36424);
and U36628 (N_36628,N_36332,N_36414);
xor U36629 (N_36629,N_36278,N_36242);
and U36630 (N_36630,N_36164,N_36252);
xor U36631 (N_36631,N_36392,N_36365);
nor U36632 (N_36632,N_36419,N_36471);
xor U36633 (N_36633,N_36205,N_36493);
xor U36634 (N_36634,N_36096,N_36168);
xor U36635 (N_36635,N_36143,N_36067);
and U36636 (N_36636,N_36045,N_36066);
and U36637 (N_36637,N_36161,N_36223);
nand U36638 (N_36638,N_36187,N_36135);
xor U36639 (N_36639,N_36130,N_36413);
and U36640 (N_36640,N_36229,N_36183);
xnor U36641 (N_36641,N_36230,N_36245);
and U36642 (N_36642,N_36268,N_36446);
xor U36643 (N_36643,N_36291,N_36296);
and U36644 (N_36644,N_36105,N_36022);
xnor U36645 (N_36645,N_36049,N_36456);
and U36646 (N_36646,N_36051,N_36287);
nand U36647 (N_36647,N_36348,N_36498);
and U36648 (N_36648,N_36076,N_36224);
nor U36649 (N_36649,N_36228,N_36169);
xor U36650 (N_36650,N_36361,N_36202);
or U36651 (N_36651,N_36036,N_36314);
or U36652 (N_36652,N_36396,N_36121);
nand U36653 (N_36653,N_36182,N_36301);
nor U36654 (N_36654,N_36329,N_36065);
nand U36655 (N_36655,N_36262,N_36214);
and U36656 (N_36656,N_36289,N_36046);
or U36657 (N_36657,N_36496,N_36227);
xnor U36658 (N_36658,N_36092,N_36116);
xor U36659 (N_36659,N_36041,N_36335);
nor U36660 (N_36660,N_36222,N_36127);
xor U36661 (N_36661,N_36328,N_36397);
and U36662 (N_36662,N_36439,N_36445);
xor U36663 (N_36663,N_36436,N_36355);
or U36664 (N_36664,N_36144,N_36233);
and U36665 (N_36665,N_36106,N_36215);
and U36666 (N_36666,N_36293,N_36172);
nor U36667 (N_36667,N_36019,N_36339);
and U36668 (N_36668,N_36231,N_36264);
nor U36669 (N_36669,N_36277,N_36418);
and U36670 (N_36670,N_36387,N_36080);
nor U36671 (N_36671,N_36434,N_36151);
nand U36672 (N_36672,N_36034,N_36197);
or U36673 (N_36673,N_36027,N_36308);
nor U36674 (N_36674,N_36148,N_36389);
nor U36675 (N_36675,N_36323,N_36159);
and U36676 (N_36676,N_36371,N_36450);
and U36677 (N_36677,N_36171,N_36011);
nand U36678 (N_36678,N_36203,N_36033);
nor U36679 (N_36679,N_36028,N_36220);
and U36680 (N_36680,N_36440,N_36218);
or U36681 (N_36681,N_36274,N_36150);
and U36682 (N_36682,N_36337,N_36009);
or U36683 (N_36683,N_36254,N_36255);
nand U36684 (N_36684,N_36152,N_36470);
nor U36685 (N_36685,N_36188,N_36055);
xor U36686 (N_36686,N_36304,N_36485);
xor U36687 (N_36687,N_36217,N_36465);
or U36688 (N_36688,N_36155,N_36017);
xor U36689 (N_36689,N_36141,N_36008);
or U36690 (N_36690,N_36292,N_36079);
xnor U36691 (N_36691,N_36226,N_36464);
and U36692 (N_36692,N_36452,N_36024);
nand U36693 (N_36693,N_36249,N_36084);
nand U36694 (N_36694,N_36399,N_36370);
and U36695 (N_36695,N_36438,N_36344);
xor U36696 (N_36696,N_36176,N_36451);
and U36697 (N_36697,N_36177,N_36495);
xnor U36698 (N_36698,N_36039,N_36061);
xor U36699 (N_36699,N_36053,N_36246);
nand U36700 (N_36700,N_36484,N_36178);
nor U36701 (N_36701,N_36093,N_36234);
or U36702 (N_36702,N_36100,N_36209);
nor U36703 (N_36703,N_36241,N_36239);
nand U36704 (N_36704,N_36179,N_36250);
nand U36705 (N_36705,N_36266,N_36212);
or U36706 (N_36706,N_36119,N_36273);
xnor U36707 (N_36707,N_36054,N_36085);
and U36708 (N_36708,N_36063,N_36149);
or U36709 (N_36709,N_36069,N_36391);
xnor U36710 (N_36710,N_36021,N_36366);
nand U36711 (N_36711,N_36430,N_36196);
xor U36712 (N_36712,N_36213,N_36087);
or U36713 (N_36713,N_36163,N_36043);
nor U36714 (N_36714,N_36459,N_36375);
nand U36715 (N_36715,N_36333,N_36240);
and U36716 (N_36716,N_36089,N_36489);
xor U36717 (N_36717,N_36074,N_36195);
nand U36718 (N_36718,N_36068,N_36175);
xor U36719 (N_36719,N_36288,N_36276);
and U36720 (N_36720,N_36295,N_36261);
xor U36721 (N_36721,N_36412,N_36050);
nand U36722 (N_36722,N_36142,N_36123);
nand U36723 (N_36723,N_36483,N_36283);
nand U36724 (N_36724,N_36455,N_36303);
nand U36725 (N_36725,N_36324,N_36443);
nand U36726 (N_36726,N_36411,N_36297);
xnor U36727 (N_36727,N_36256,N_36099);
or U36728 (N_36728,N_36235,N_36007);
and U36729 (N_36729,N_36453,N_36015);
nand U36730 (N_36730,N_36137,N_36457);
xnor U36731 (N_36731,N_36097,N_36107);
nand U36732 (N_36732,N_36405,N_36422);
nand U36733 (N_36733,N_36343,N_36284);
nor U36734 (N_36734,N_36461,N_36367);
nor U36735 (N_36735,N_36432,N_36381);
or U36736 (N_36736,N_36298,N_36316);
nor U36737 (N_36737,N_36330,N_36497);
nor U36738 (N_36738,N_36334,N_36319);
xnor U36739 (N_36739,N_36263,N_36258);
nand U36740 (N_36740,N_36458,N_36423);
xnor U36741 (N_36741,N_36454,N_36115);
xnor U36742 (N_36742,N_36408,N_36492);
xor U36743 (N_36743,N_36463,N_36307);
or U36744 (N_36744,N_36351,N_36117);
nand U36745 (N_36745,N_36380,N_36374);
xor U36746 (N_36746,N_36267,N_36070);
or U36747 (N_36747,N_36101,N_36129);
or U36748 (N_36748,N_36299,N_36321);
nand U36749 (N_36749,N_36102,N_36360);
nor U36750 (N_36750,N_36081,N_36280);
and U36751 (N_36751,N_36292,N_36302);
nand U36752 (N_36752,N_36116,N_36213);
or U36753 (N_36753,N_36407,N_36354);
xnor U36754 (N_36754,N_36454,N_36450);
and U36755 (N_36755,N_36403,N_36275);
and U36756 (N_36756,N_36205,N_36065);
nor U36757 (N_36757,N_36036,N_36046);
and U36758 (N_36758,N_36121,N_36293);
nand U36759 (N_36759,N_36242,N_36128);
and U36760 (N_36760,N_36318,N_36032);
and U36761 (N_36761,N_36110,N_36097);
xnor U36762 (N_36762,N_36298,N_36465);
and U36763 (N_36763,N_36124,N_36040);
and U36764 (N_36764,N_36431,N_36439);
xor U36765 (N_36765,N_36280,N_36232);
xnor U36766 (N_36766,N_36296,N_36267);
nand U36767 (N_36767,N_36233,N_36288);
nand U36768 (N_36768,N_36333,N_36144);
nand U36769 (N_36769,N_36104,N_36439);
nor U36770 (N_36770,N_36256,N_36177);
nor U36771 (N_36771,N_36283,N_36209);
nand U36772 (N_36772,N_36091,N_36227);
nor U36773 (N_36773,N_36262,N_36127);
xor U36774 (N_36774,N_36182,N_36216);
or U36775 (N_36775,N_36124,N_36407);
or U36776 (N_36776,N_36306,N_36462);
or U36777 (N_36777,N_36174,N_36126);
and U36778 (N_36778,N_36056,N_36490);
nand U36779 (N_36779,N_36105,N_36423);
xor U36780 (N_36780,N_36172,N_36421);
or U36781 (N_36781,N_36483,N_36397);
nand U36782 (N_36782,N_36100,N_36048);
nand U36783 (N_36783,N_36064,N_36134);
nand U36784 (N_36784,N_36472,N_36045);
nand U36785 (N_36785,N_36012,N_36006);
or U36786 (N_36786,N_36170,N_36103);
or U36787 (N_36787,N_36221,N_36483);
xor U36788 (N_36788,N_36474,N_36326);
or U36789 (N_36789,N_36368,N_36078);
xor U36790 (N_36790,N_36319,N_36137);
nand U36791 (N_36791,N_36426,N_36342);
or U36792 (N_36792,N_36143,N_36230);
and U36793 (N_36793,N_36461,N_36303);
nor U36794 (N_36794,N_36226,N_36197);
nand U36795 (N_36795,N_36193,N_36353);
or U36796 (N_36796,N_36055,N_36390);
xnor U36797 (N_36797,N_36275,N_36016);
nand U36798 (N_36798,N_36162,N_36364);
nand U36799 (N_36799,N_36258,N_36198);
xor U36800 (N_36800,N_36157,N_36328);
or U36801 (N_36801,N_36421,N_36108);
or U36802 (N_36802,N_36390,N_36101);
and U36803 (N_36803,N_36244,N_36031);
nand U36804 (N_36804,N_36374,N_36486);
or U36805 (N_36805,N_36081,N_36295);
xor U36806 (N_36806,N_36294,N_36295);
nand U36807 (N_36807,N_36209,N_36008);
nand U36808 (N_36808,N_36250,N_36246);
or U36809 (N_36809,N_36076,N_36287);
nor U36810 (N_36810,N_36244,N_36060);
and U36811 (N_36811,N_36178,N_36437);
nor U36812 (N_36812,N_36294,N_36127);
or U36813 (N_36813,N_36253,N_36304);
xor U36814 (N_36814,N_36113,N_36367);
nand U36815 (N_36815,N_36013,N_36430);
nor U36816 (N_36816,N_36245,N_36104);
xnor U36817 (N_36817,N_36063,N_36303);
nand U36818 (N_36818,N_36201,N_36367);
or U36819 (N_36819,N_36374,N_36385);
nor U36820 (N_36820,N_36251,N_36062);
and U36821 (N_36821,N_36165,N_36022);
xnor U36822 (N_36822,N_36338,N_36101);
and U36823 (N_36823,N_36385,N_36138);
and U36824 (N_36824,N_36193,N_36383);
and U36825 (N_36825,N_36492,N_36227);
and U36826 (N_36826,N_36156,N_36081);
nor U36827 (N_36827,N_36293,N_36320);
nor U36828 (N_36828,N_36289,N_36434);
nor U36829 (N_36829,N_36408,N_36055);
or U36830 (N_36830,N_36343,N_36165);
xnor U36831 (N_36831,N_36320,N_36415);
nor U36832 (N_36832,N_36091,N_36389);
and U36833 (N_36833,N_36176,N_36212);
nor U36834 (N_36834,N_36269,N_36446);
nor U36835 (N_36835,N_36085,N_36358);
xnor U36836 (N_36836,N_36119,N_36405);
or U36837 (N_36837,N_36471,N_36389);
xor U36838 (N_36838,N_36084,N_36025);
nand U36839 (N_36839,N_36280,N_36188);
or U36840 (N_36840,N_36440,N_36414);
nand U36841 (N_36841,N_36239,N_36236);
and U36842 (N_36842,N_36015,N_36066);
xnor U36843 (N_36843,N_36238,N_36081);
or U36844 (N_36844,N_36310,N_36252);
nor U36845 (N_36845,N_36452,N_36087);
or U36846 (N_36846,N_36286,N_36464);
and U36847 (N_36847,N_36261,N_36097);
xnor U36848 (N_36848,N_36154,N_36307);
and U36849 (N_36849,N_36295,N_36397);
or U36850 (N_36850,N_36350,N_36083);
or U36851 (N_36851,N_36256,N_36326);
nor U36852 (N_36852,N_36494,N_36261);
nand U36853 (N_36853,N_36153,N_36180);
xnor U36854 (N_36854,N_36152,N_36255);
and U36855 (N_36855,N_36135,N_36029);
and U36856 (N_36856,N_36463,N_36066);
xor U36857 (N_36857,N_36449,N_36476);
and U36858 (N_36858,N_36153,N_36300);
nor U36859 (N_36859,N_36146,N_36387);
nand U36860 (N_36860,N_36435,N_36204);
nor U36861 (N_36861,N_36115,N_36147);
nor U36862 (N_36862,N_36453,N_36471);
nor U36863 (N_36863,N_36228,N_36482);
nor U36864 (N_36864,N_36037,N_36162);
and U36865 (N_36865,N_36091,N_36063);
nor U36866 (N_36866,N_36293,N_36130);
xor U36867 (N_36867,N_36196,N_36349);
nor U36868 (N_36868,N_36360,N_36190);
or U36869 (N_36869,N_36100,N_36375);
nor U36870 (N_36870,N_36214,N_36454);
or U36871 (N_36871,N_36366,N_36286);
nand U36872 (N_36872,N_36026,N_36466);
and U36873 (N_36873,N_36068,N_36035);
xnor U36874 (N_36874,N_36387,N_36027);
or U36875 (N_36875,N_36147,N_36247);
xor U36876 (N_36876,N_36263,N_36451);
and U36877 (N_36877,N_36023,N_36287);
or U36878 (N_36878,N_36416,N_36234);
xor U36879 (N_36879,N_36068,N_36078);
nand U36880 (N_36880,N_36496,N_36255);
nor U36881 (N_36881,N_36077,N_36197);
or U36882 (N_36882,N_36461,N_36447);
nor U36883 (N_36883,N_36454,N_36474);
xnor U36884 (N_36884,N_36172,N_36390);
nor U36885 (N_36885,N_36161,N_36031);
xnor U36886 (N_36886,N_36337,N_36497);
nand U36887 (N_36887,N_36062,N_36112);
nor U36888 (N_36888,N_36154,N_36238);
and U36889 (N_36889,N_36253,N_36278);
and U36890 (N_36890,N_36418,N_36221);
nor U36891 (N_36891,N_36194,N_36350);
and U36892 (N_36892,N_36054,N_36013);
and U36893 (N_36893,N_36400,N_36062);
or U36894 (N_36894,N_36193,N_36274);
and U36895 (N_36895,N_36259,N_36130);
or U36896 (N_36896,N_36228,N_36312);
nand U36897 (N_36897,N_36433,N_36400);
nor U36898 (N_36898,N_36433,N_36301);
xnor U36899 (N_36899,N_36221,N_36069);
xnor U36900 (N_36900,N_36342,N_36032);
and U36901 (N_36901,N_36376,N_36338);
nand U36902 (N_36902,N_36065,N_36475);
or U36903 (N_36903,N_36101,N_36393);
xnor U36904 (N_36904,N_36452,N_36051);
xor U36905 (N_36905,N_36069,N_36290);
nor U36906 (N_36906,N_36170,N_36003);
and U36907 (N_36907,N_36134,N_36148);
nor U36908 (N_36908,N_36042,N_36415);
xnor U36909 (N_36909,N_36172,N_36428);
or U36910 (N_36910,N_36164,N_36340);
or U36911 (N_36911,N_36080,N_36069);
and U36912 (N_36912,N_36327,N_36281);
xnor U36913 (N_36913,N_36482,N_36471);
nor U36914 (N_36914,N_36234,N_36390);
nand U36915 (N_36915,N_36479,N_36055);
or U36916 (N_36916,N_36387,N_36055);
xor U36917 (N_36917,N_36382,N_36151);
nor U36918 (N_36918,N_36093,N_36455);
nand U36919 (N_36919,N_36474,N_36343);
nand U36920 (N_36920,N_36414,N_36325);
nor U36921 (N_36921,N_36325,N_36053);
and U36922 (N_36922,N_36291,N_36490);
nor U36923 (N_36923,N_36404,N_36189);
nor U36924 (N_36924,N_36371,N_36317);
nor U36925 (N_36925,N_36417,N_36022);
nand U36926 (N_36926,N_36105,N_36029);
xnor U36927 (N_36927,N_36220,N_36465);
nand U36928 (N_36928,N_36355,N_36211);
and U36929 (N_36929,N_36400,N_36071);
xnor U36930 (N_36930,N_36157,N_36456);
or U36931 (N_36931,N_36409,N_36213);
and U36932 (N_36932,N_36459,N_36109);
and U36933 (N_36933,N_36410,N_36010);
nand U36934 (N_36934,N_36407,N_36494);
nor U36935 (N_36935,N_36413,N_36398);
or U36936 (N_36936,N_36034,N_36431);
or U36937 (N_36937,N_36415,N_36302);
nand U36938 (N_36938,N_36312,N_36024);
xnor U36939 (N_36939,N_36379,N_36404);
xnor U36940 (N_36940,N_36446,N_36497);
xor U36941 (N_36941,N_36249,N_36082);
or U36942 (N_36942,N_36035,N_36408);
and U36943 (N_36943,N_36286,N_36354);
xor U36944 (N_36944,N_36211,N_36417);
xnor U36945 (N_36945,N_36378,N_36343);
nor U36946 (N_36946,N_36224,N_36254);
and U36947 (N_36947,N_36482,N_36113);
nand U36948 (N_36948,N_36259,N_36085);
nand U36949 (N_36949,N_36438,N_36429);
and U36950 (N_36950,N_36118,N_36156);
or U36951 (N_36951,N_36402,N_36385);
nor U36952 (N_36952,N_36128,N_36419);
and U36953 (N_36953,N_36388,N_36184);
nor U36954 (N_36954,N_36484,N_36314);
and U36955 (N_36955,N_36488,N_36267);
xor U36956 (N_36956,N_36117,N_36182);
or U36957 (N_36957,N_36405,N_36444);
xnor U36958 (N_36958,N_36487,N_36381);
nand U36959 (N_36959,N_36458,N_36051);
nand U36960 (N_36960,N_36004,N_36308);
xnor U36961 (N_36961,N_36287,N_36428);
xnor U36962 (N_36962,N_36225,N_36181);
xnor U36963 (N_36963,N_36350,N_36405);
or U36964 (N_36964,N_36414,N_36395);
nand U36965 (N_36965,N_36153,N_36215);
and U36966 (N_36966,N_36211,N_36255);
nand U36967 (N_36967,N_36363,N_36142);
nor U36968 (N_36968,N_36145,N_36364);
and U36969 (N_36969,N_36300,N_36384);
nor U36970 (N_36970,N_36472,N_36101);
and U36971 (N_36971,N_36413,N_36203);
xor U36972 (N_36972,N_36005,N_36488);
xnor U36973 (N_36973,N_36433,N_36004);
and U36974 (N_36974,N_36345,N_36166);
and U36975 (N_36975,N_36212,N_36189);
nand U36976 (N_36976,N_36236,N_36244);
and U36977 (N_36977,N_36133,N_36372);
or U36978 (N_36978,N_36398,N_36166);
xnor U36979 (N_36979,N_36184,N_36333);
xor U36980 (N_36980,N_36358,N_36067);
xnor U36981 (N_36981,N_36082,N_36014);
and U36982 (N_36982,N_36388,N_36105);
xor U36983 (N_36983,N_36155,N_36101);
or U36984 (N_36984,N_36008,N_36202);
nand U36985 (N_36985,N_36294,N_36067);
nor U36986 (N_36986,N_36213,N_36055);
nand U36987 (N_36987,N_36178,N_36221);
xor U36988 (N_36988,N_36169,N_36266);
or U36989 (N_36989,N_36192,N_36493);
nand U36990 (N_36990,N_36143,N_36083);
and U36991 (N_36991,N_36183,N_36495);
nand U36992 (N_36992,N_36288,N_36109);
and U36993 (N_36993,N_36236,N_36165);
nand U36994 (N_36994,N_36049,N_36219);
or U36995 (N_36995,N_36482,N_36385);
nand U36996 (N_36996,N_36327,N_36252);
or U36997 (N_36997,N_36353,N_36499);
nor U36998 (N_36998,N_36309,N_36353);
xnor U36999 (N_36999,N_36023,N_36272);
or U37000 (N_37000,N_36547,N_36643);
or U37001 (N_37001,N_36544,N_36542);
nand U37002 (N_37002,N_36852,N_36677);
and U37003 (N_37003,N_36989,N_36641);
xnor U37004 (N_37004,N_36631,N_36799);
or U37005 (N_37005,N_36898,N_36530);
and U37006 (N_37006,N_36854,N_36500);
or U37007 (N_37007,N_36980,N_36859);
nand U37008 (N_37008,N_36976,N_36731);
xor U37009 (N_37009,N_36605,N_36981);
or U37010 (N_37010,N_36795,N_36746);
and U37011 (N_37011,N_36591,N_36907);
nand U37012 (N_37012,N_36900,N_36588);
nor U37013 (N_37013,N_36817,N_36932);
xor U37014 (N_37014,N_36628,N_36949);
xor U37015 (N_37015,N_36750,N_36866);
nor U37016 (N_37016,N_36915,N_36566);
nor U37017 (N_37017,N_36658,N_36992);
nand U37018 (N_37018,N_36742,N_36735);
or U37019 (N_37019,N_36702,N_36648);
or U37020 (N_37020,N_36765,N_36804);
nand U37021 (N_37021,N_36766,N_36574);
xor U37022 (N_37022,N_36726,N_36990);
or U37023 (N_37023,N_36539,N_36667);
nor U37024 (N_37024,N_36871,N_36853);
and U37025 (N_37025,N_36587,N_36708);
xor U37026 (N_37026,N_36729,N_36982);
xnor U37027 (N_37027,N_36665,N_36808);
or U37028 (N_37028,N_36576,N_36528);
xor U37029 (N_37029,N_36991,N_36621);
nor U37030 (N_37030,N_36843,N_36678);
or U37031 (N_37031,N_36759,N_36897);
and U37032 (N_37032,N_36724,N_36778);
nor U37033 (N_37033,N_36962,N_36944);
nor U37034 (N_37034,N_36770,N_36596);
nor U37035 (N_37035,N_36988,N_36793);
and U37036 (N_37036,N_36855,N_36771);
or U37037 (N_37037,N_36748,N_36821);
nor U37038 (N_37038,N_36856,N_36565);
and U37039 (N_37039,N_36790,N_36536);
nand U37040 (N_37040,N_36584,N_36783);
nor U37041 (N_37041,N_36986,N_36929);
or U37042 (N_37042,N_36590,N_36598);
xnor U37043 (N_37043,N_36619,N_36837);
and U37044 (N_37044,N_36922,N_36977);
nor U37045 (N_37045,N_36503,N_36510);
or U37046 (N_37046,N_36847,N_36664);
nor U37047 (N_37047,N_36796,N_36822);
and U37048 (N_37048,N_36521,N_36802);
xor U37049 (N_37049,N_36589,N_36662);
and U37050 (N_37050,N_36580,N_36827);
and U37051 (N_37051,N_36940,N_36921);
and U37052 (N_37052,N_36983,N_36654);
and U37053 (N_37053,N_36918,N_36970);
or U37054 (N_37054,N_36506,N_36823);
and U37055 (N_37055,N_36561,N_36908);
nor U37056 (N_37056,N_36762,N_36798);
xor U37057 (N_37057,N_36943,N_36519);
nand U37058 (N_37058,N_36692,N_36686);
xnor U37059 (N_37059,N_36541,N_36672);
xor U37060 (N_37060,N_36809,N_36937);
xor U37061 (N_37061,N_36518,N_36858);
xor U37062 (N_37062,N_36568,N_36999);
nor U37063 (N_37063,N_36893,N_36867);
nor U37064 (N_37064,N_36820,N_36706);
nand U37065 (N_37065,N_36913,N_36961);
and U37066 (N_37066,N_36743,N_36507);
or U37067 (N_37067,N_36603,N_36984);
xor U37068 (N_37068,N_36604,N_36681);
or U37069 (N_37069,N_36998,N_36563);
nand U37070 (N_37070,N_36673,N_36830);
nand U37071 (N_37071,N_36972,N_36780);
nor U37072 (N_37072,N_36951,N_36714);
xnor U37073 (N_37073,N_36652,N_36791);
and U37074 (N_37074,N_36693,N_36894);
or U37075 (N_37075,N_36878,N_36892);
nor U37076 (N_37076,N_36578,N_36734);
xnor U37077 (N_37077,N_36785,N_36501);
nor U37078 (N_37078,N_36575,N_36716);
nand U37079 (N_37079,N_36873,N_36535);
and U37080 (N_37080,N_36924,N_36527);
and U37081 (N_37081,N_36828,N_36602);
xnor U37082 (N_37082,N_36698,N_36857);
or U37083 (N_37083,N_36869,N_36711);
nand U37084 (N_37084,N_36845,N_36522);
nand U37085 (N_37085,N_36777,N_36829);
nor U37086 (N_37086,N_36747,N_36901);
and U37087 (N_37087,N_36646,N_36659);
nor U37088 (N_37088,N_36660,N_36933);
or U37089 (N_37089,N_36835,N_36567);
xnor U37090 (N_37090,N_36638,N_36649);
nand U37091 (N_37091,N_36966,N_36789);
xnor U37092 (N_37092,N_36755,N_36650);
xnor U37093 (N_37093,N_36640,N_36624);
or U37094 (N_37094,N_36959,N_36995);
xnor U37095 (N_37095,N_36850,N_36739);
nor U37096 (N_37096,N_36931,N_36722);
xnor U37097 (N_37097,N_36564,N_36801);
nor U37098 (N_37098,N_36571,N_36516);
and U37099 (N_37099,N_36926,N_36616);
xor U37100 (N_37100,N_36614,N_36668);
nor U37101 (N_37101,N_36888,N_36751);
and U37102 (N_37102,N_36537,N_36987);
or U37103 (N_37103,N_36582,N_36737);
or U37104 (N_37104,N_36644,N_36594);
xnor U37105 (N_37105,N_36890,N_36600);
nand U37106 (N_37106,N_36834,N_36816);
and U37107 (N_37107,N_36964,N_36680);
nand U37108 (N_37108,N_36841,N_36627);
nand U37109 (N_37109,N_36625,N_36675);
and U37110 (N_37110,N_36910,N_36942);
or U37111 (N_37111,N_36727,N_36691);
nor U37112 (N_37112,N_36552,N_36695);
nor U37113 (N_37113,N_36916,N_36904);
and U37114 (N_37114,N_36586,N_36776);
or U37115 (N_37115,N_36930,N_36917);
nand U37116 (N_37116,N_36811,N_36630);
nand U37117 (N_37117,N_36914,N_36657);
or U37118 (N_37118,N_36744,N_36532);
nand U37119 (N_37119,N_36872,N_36514);
xnor U37120 (N_37120,N_36774,N_36806);
or U37121 (N_37121,N_36760,N_36974);
nor U37122 (N_37122,N_36939,N_36736);
nand U37123 (N_37123,N_36938,N_36663);
nor U37124 (N_37124,N_36513,N_36697);
or U37125 (N_37125,N_36725,N_36612);
nor U37126 (N_37126,N_36676,N_36819);
nand U37127 (N_37127,N_36839,N_36842);
xnor U37128 (N_37128,N_36607,N_36875);
or U37129 (N_37129,N_36891,N_36953);
or U37130 (N_37130,N_36812,N_36669);
xor U37131 (N_37131,N_36963,N_36740);
or U37132 (N_37132,N_36548,N_36560);
xnor U37133 (N_37133,N_36965,N_36606);
and U37134 (N_37134,N_36905,N_36956);
or U37135 (N_37135,N_36865,N_36985);
xnor U37136 (N_37136,N_36868,N_36690);
or U37137 (N_37137,N_36769,N_36846);
or U37138 (N_37138,N_36849,N_36967);
or U37139 (N_37139,N_36557,N_36699);
or U37140 (N_37140,N_36874,N_36880);
nand U37141 (N_37141,N_36694,N_36703);
nand U37142 (N_37142,N_36832,N_36608);
or U37143 (N_37143,N_36794,N_36948);
and U37144 (N_37144,N_36733,N_36622);
or U37145 (N_37145,N_36800,N_36626);
xor U37146 (N_37146,N_36538,N_36623);
nand U37147 (N_37147,N_36807,N_36585);
and U37148 (N_37148,N_36840,N_36520);
nand U37149 (N_37149,N_36613,N_36844);
and U37150 (N_37150,N_36955,N_36745);
nor U37151 (N_37151,N_36969,N_36597);
xor U37152 (N_37152,N_36764,N_36524);
and U37153 (N_37153,N_36838,N_36958);
xnor U37154 (N_37154,N_36996,N_36579);
nand U37155 (N_37155,N_36687,N_36732);
and U37156 (N_37156,N_36583,N_36928);
nor U37157 (N_37157,N_36592,N_36884);
xor U37158 (N_37158,N_36719,N_36886);
xor U37159 (N_37159,N_36525,N_36670);
or U37160 (N_37160,N_36851,N_36912);
xnor U37161 (N_37161,N_36899,N_36863);
nor U37162 (N_37162,N_36814,N_36688);
nand U37163 (N_37163,N_36749,N_36753);
or U37164 (N_37164,N_36555,N_36666);
xor U37165 (N_37165,N_36876,N_36717);
nand U37166 (N_37166,N_36581,N_36730);
and U37167 (N_37167,N_36848,N_36639);
or U37168 (N_37168,N_36946,N_36954);
and U37169 (N_37169,N_36925,N_36610);
nand U37170 (N_37170,N_36718,N_36881);
nor U37171 (N_37171,N_36709,N_36710);
nand U37172 (N_37172,N_36927,N_36551);
nor U37173 (N_37173,N_36712,N_36685);
xor U37174 (N_37174,N_36601,N_36684);
nor U37175 (N_37175,N_36689,N_36636);
xnor U37176 (N_37176,N_36906,N_36818);
and U37177 (N_37177,N_36617,N_36788);
nand U37178 (N_37178,N_36833,N_36864);
xnor U37179 (N_37179,N_36994,N_36756);
xor U37180 (N_37180,N_36661,N_36651);
or U37181 (N_37181,N_36782,N_36887);
or U37182 (N_37182,N_36787,N_36637);
nor U37183 (N_37183,N_36653,N_36502);
xnor U37184 (N_37184,N_36883,N_36877);
and U37185 (N_37185,N_36505,N_36784);
xnor U37186 (N_37186,N_36618,N_36553);
nor U37187 (N_37187,N_36723,N_36549);
or U37188 (N_37188,N_36978,N_36655);
nor U37189 (N_37189,N_36550,N_36968);
and U37190 (N_37190,N_36936,N_36508);
xnor U37191 (N_37191,N_36920,N_36645);
nor U37192 (N_37192,N_36862,N_36570);
or U37193 (N_37193,N_36517,N_36803);
or U37194 (N_37194,N_36558,N_36772);
nor U37195 (N_37195,N_36629,N_36533);
and U37196 (N_37196,N_36810,N_36674);
xnor U37197 (N_37197,N_36879,N_36615);
xnor U37198 (N_37198,N_36781,N_36633);
nor U37199 (N_37199,N_36559,N_36611);
and U37200 (N_37200,N_36973,N_36775);
nand U37201 (N_37201,N_36504,N_36923);
nor U37202 (N_37202,N_36919,N_36902);
or U37203 (N_37203,N_36885,N_36761);
nand U37204 (N_37204,N_36721,N_36682);
xor U37205 (N_37205,N_36825,N_36993);
or U37206 (N_37206,N_36546,N_36741);
xor U37207 (N_37207,N_36554,N_36713);
nand U37208 (N_37208,N_36701,N_36700);
xnor U37209 (N_37209,N_36509,N_36909);
xnor U37210 (N_37210,N_36971,N_36599);
and U37211 (N_37211,N_36515,N_36813);
nand U37212 (N_37212,N_36556,N_36754);
xnor U37213 (N_37213,N_36805,N_36895);
or U37214 (N_37214,N_36534,N_36882);
and U37215 (N_37215,N_36935,N_36773);
or U37216 (N_37216,N_36786,N_36860);
nand U37217 (N_37217,N_36620,N_36950);
nor U37218 (N_37218,N_36836,N_36797);
nor U37219 (N_37219,N_36767,N_36632);
and U37220 (N_37220,N_36831,N_36934);
xnor U37221 (N_37221,N_36715,N_36941);
and U37222 (N_37222,N_36815,N_36523);
nor U37223 (N_37223,N_36569,N_36911);
xor U37224 (N_37224,N_36647,N_36683);
nand U37225 (N_37225,N_36572,N_36512);
or U37226 (N_37226,N_36824,N_36738);
nor U37227 (N_37227,N_36792,N_36511);
nor U37228 (N_37228,N_36526,N_36768);
or U37229 (N_37229,N_36896,N_36577);
nor U37230 (N_37230,N_36634,N_36529);
or U37231 (N_37231,N_36758,N_36543);
nor U37232 (N_37232,N_36679,N_36609);
and U37233 (N_37233,N_36696,N_36975);
or U37234 (N_37234,N_36562,N_36656);
nor U37235 (N_37235,N_36635,N_36671);
nand U37236 (N_37236,N_36903,N_36979);
or U37237 (N_37237,N_36763,N_36960);
xnor U37238 (N_37238,N_36704,N_36705);
nor U37239 (N_37239,N_36720,N_36573);
nand U37240 (N_37240,N_36752,N_36861);
or U37241 (N_37241,N_36870,N_36707);
nor U37242 (N_37242,N_36779,N_36826);
and U37243 (N_37243,N_36593,N_36531);
nand U37244 (N_37244,N_36642,N_36889);
and U37245 (N_37245,N_36952,N_36945);
nor U37246 (N_37246,N_36947,N_36957);
and U37247 (N_37247,N_36728,N_36545);
xor U37248 (N_37248,N_36595,N_36997);
and U37249 (N_37249,N_36540,N_36757);
xnor U37250 (N_37250,N_36633,N_36510);
nand U37251 (N_37251,N_36813,N_36985);
xor U37252 (N_37252,N_36864,N_36968);
nand U37253 (N_37253,N_36872,N_36982);
nand U37254 (N_37254,N_36910,N_36577);
or U37255 (N_37255,N_36953,N_36912);
nand U37256 (N_37256,N_36984,N_36675);
and U37257 (N_37257,N_36553,N_36877);
and U37258 (N_37258,N_36999,N_36960);
nand U37259 (N_37259,N_36886,N_36889);
and U37260 (N_37260,N_36599,N_36646);
xnor U37261 (N_37261,N_36729,N_36730);
xnor U37262 (N_37262,N_36528,N_36793);
nor U37263 (N_37263,N_36992,N_36536);
and U37264 (N_37264,N_36729,N_36826);
nand U37265 (N_37265,N_36687,N_36672);
nor U37266 (N_37266,N_36828,N_36841);
and U37267 (N_37267,N_36567,N_36532);
nor U37268 (N_37268,N_36712,N_36805);
xnor U37269 (N_37269,N_36720,N_36715);
or U37270 (N_37270,N_36972,N_36755);
and U37271 (N_37271,N_36710,N_36897);
xnor U37272 (N_37272,N_36920,N_36774);
and U37273 (N_37273,N_36940,N_36827);
or U37274 (N_37274,N_36540,N_36682);
xor U37275 (N_37275,N_36537,N_36648);
nand U37276 (N_37276,N_36760,N_36667);
xor U37277 (N_37277,N_36520,N_36599);
or U37278 (N_37278,N_36630,N_36767);
xnor U37279 (N_37279,N_36842,N_36787);
xor U37280 (N_37280,N_36509,N_36848);
and U37281 (N_37281,N_36711,N_36549);
and U37282 (N_37282,N_36899,N_36997);
and U37283 (N_37283,N_36973,N_36671);
nand U37284 (N_37284,N_36668,N_36520);
xor U37285 (N_37285,N_36683,N_36580);
nand U37286 (N_37286,N_36747,N_36537);
nand U37287 (N_37287,N_36529,N_36849);
or U37288 (N_37288,N_36844,N_36598);
and U37289 (N_37289,N_36771,N_36916);
nor U37290 (N_37290,N_36891,N_36722);
nor U37291 (N_37291,N_36876,N_36827);
nor U37292 (N_37292,N_36704,N_36926);
and U37293 (N_37293,N_36718,N_36626);
or U37294 (N_37294,N_36594,N_36753);
xnor U37295 (N_37295,N_36844,N_36892);
nor U37296 (N_37296,N_36637,N_36544);
nand U37297 (N_37297,N_36822,N_36644);
xnor U37298 (N_37298,N_36785,N_36600);
and U37299 (N_37299,N_36909,N_36856);
and U37300 (N_37300,N_36619,N_36635);
xor U37301 (N_37301,N_36998,N_36633);
nor U37302 (N_37302,N_36606,N_36788);
or U37303 (N_37303,N_36965,N_36810);
nor U37304 (N_37304,N_36582,N_36705);
nor U37305 (N_37305,N_36727,N_36980);
nor U37306 (N_37306,N_36684,N_36896);
xnor U37307 (N_37307,N_36821,N_36505);
nor U37308 (N_37308,N_36729,N_36529);
xor U37309 (N_37309,N_36649,N_36731);
nand U37310 (N_37310,N_36639,N_36859);
or U37311 (N_37311,N_36595,N_36736);
nand U37312 (N_37312,N_36531,N_36611);
and U37313 (N_37313,N_36702,N_36605);
nand U37314 (N_37314,N_36513,N_36970);
and U37315 (N_37315,N_36878,N_36578);
xnor U37316 (N_37316,N_36647,N_36712);
and U37317 (N_37317,N_36906,N_36902);
or U37318 (N_37318,N_36631,N_36812);
nor U37319 (N_37319,N_36537,N_36835);
and U37320 (N_37320,N_36774,N_36651);
xor U37321 (N_37321,N_36933,N_36590);
and U37322 (N_37322,N_36846,N_36553);
nor U37323 (N_37323,N_36820,N_36888);
nand U37324 (N_37324,N_36506,N_36584);
or U37325 (N_37325,N_36995,N_36795);
or U37326 (N_37326,N_36511,N_36986);
xnor U37327 (N_37327,N_36669,N_36633);
nand U37328 (N_37328,N_36634,N_36875);
nand U37329 (N_37329,N_36690,N_36569);
nand U37330 (N_37330,N_36662,N_36887);
and U37331 (N_37331,N_36513,N_36862);
xor U37332 (N_37332,N_36857,N_36639);
nor U37333 (N_37333,N_36957,N_36621);
nor U37334 (N_37334,N_36554,N_36956);
nor U37335 (N_37335,N_36916,N_36758);
xor U37336 (N_37336,N_36634,N_36561);
nand U37337 (N_37337,N_36995,N_36788);
or U37338 (N_37338,N_36777,N_36534);
xor U37339 (N_37339,N_36648,N_36766);
nor U37340 (N_37340,N_36866,N_36687);
xor U37341 (N_37341,N_36873,N_36596);
nor U37342 (N_37342,N_36954,N_36933);
nand U37343 (N_37343,N_36794,N_36509);
nor U37344 (N_37344,N_36581,N_36861);
nand U37345 (N_37345,N_36742,N_36921);
nand U37346 (N_37346,N_36557,N_36623);
nor U37347 (N_37347,N_36697,N_36724);
nor U37348 (N_37348,N_36580,N_36763);
nor U37349 (N_37349,N_36837,N_36688);
or U37350 (N_37350,N_36628,N_36551);
nand U37351 (N_37351,N_36946,N_36980);
or U37352 (N_37352,N_36733,N_36737);
and U37353 (N_37353,N_36538,N_36754);
or U37354 (N_37354,N_36812,N_36587);
xnor U37355 (N_37355,N_36596,N_36575);
nand U37356 (N_37356,N_36957,N_36775);
xor U37357 (N_37357,N_36738,N_36708);
nand U37358 (N_37358,N_36834,N_36662);
nand U37359 (N_37359,N_36804,N_36628);
nand U37360 (N_37360,N_36613,N_36897);
or U37361 (N_37361,N_36945,N_36562);
nor U37362 (N_37362,N_36901,N_36524);
nand U37363 (N_37363,N_36539,N_36560);
xor U37364 (N_37364,N_36632,N_36868);
nand U37365 (N_37365,N_36803,N_36775);
nand U37366 (N_37366,N_36620,N_36944);
nand U37367 (N_37367,N_36644,N_36872);
and U37368 (N_37368,N_36808,N_36789);
xnor U37369 (N_37369,N_36752,N_36943);
nand U37370 (N_37370,N_36798,N_36733);
or U37371 (N_37371,N_36618,N_36854);
nor U37372 (N_37372,N_36859,N_36529);
nor U37373 (N_37373,N_36531,N_36904);
and U37374 (N_37374,N_36727,N_36669);
xnor U37375 (N_37375,N_36587,N_36677);
or U37376 (N_37376,N_36802,N_36612);
or U37377 (N_37377,N_36619,N_36568);
nand U37378 (N_37378,N_36801,N_36887);
nand U37379 (N_37379,N_36672,N_36539);
and U37380 (N_37380,N_36731,N_36530);
xor U37381 (N_37381,N_36504,N_36513);
xnor U37382 (N_37382,N_36791,N_36843);
xnor U37383 (N_37383,N_36732,N_36887);
xor U37384 (N_37384,N_36754,N_36503);
nand U37385 (N_37385,N_36580,N_36690);
nand U37386 (N_37386,N_36601,N_36535);
nand U37387 (N_37387,N_36890,N_36584);
or U37388 (N_37388,N_36719,N_36607);
and U37389 (N_37389,N_36523,N_36538);
xnor U37390 (N_37390,N_36665,N_36636);
or U37391 (N_37391,N_36706,N_36933);
nor U37392 (N_37392,N_36530,N_36841);
nor U37393 (N_37393,N_36844,N_36810);
xor U37394 (N_37394,N_36808,N_36724);
nand U37395 (N_37395,N_36854,N_36661);
and U37396 (N_37396,N_36563,N_36937);
nor U37397 (N_37397,N_36934,N_36599);
xnor U37398 (N_37398,N_36766,N_36715);
nor U37399 (N_37399,N_36802,N_36614);
and U37400 (N_37400,N_36835,N_36633);
or U37401 (N_37401,N_36657,N_36571);
xnor U37402 (N_37402,N_36650,N_36866);
nor U37403 (N_37403,N_36976,N_36529);
xor U37404 (N_37404,N_36710,N_36926);
nor U37405 (N_37405,N_36557,N_36821);
nand U37406 (N_37406,N_36943,N_36690);
and U37407 (N_37407,N_36656,N_36762);
nand U37408 (N_37408,N_36683,N_36839);
nand U37409 (N_37409,N_36838,N_36632);
and U37410 (N_37410,N_36795,N_36714);
nand U37411 (N_37411,N_36609,N_36668);
nor U37412 (N_37412,N_36836,N_36904);
nand U37413 (N_37413,N_36786,N_36603);
nor U37414 (N_37414,N_36738,N_36672);
xnor U37415 (N_37415,N_36629,N_36613);
nand U37416 (N_37416,N_36733,N_36589);
and U37417 (N_37417,N_36583,N_36529);
xnor U37418 (N_37418,N_36608,N_36521);
or U37419 (N_37419,N_36867,N_36552);
and U37420 (N_37420,N_36560,N_36604);
or U37421 (N_37421,N_36879,N_36729);
xor U37422 (N_37422,N_36974,N_36611);
nor U37423 (N_37423,N_36858,N_36987);
or U37424 (N_37424,N_36635,N_36871);
nand U37425 (N_37425,N_36778,N_36718);
xnor U37426 (N_37426,N_36821,N_36972);
or U37427 (N_37427,N_36658,N_36631);
nand U37428 (N_37428,N_36657,N_36873);
nor U37429 (N_37429,N_36672,N_36511);
and U37430 (N_37430,N_36746,N_36879);
nand U37431 (N_37431,N_36720,N_36819);
and U37432 (N_37432,N_36968,N_36875);
nor U37433 (N_37433,N_36838,N_36514);
nand U37434 (N_37434,N_36701,N_36942);
nand U37435 (N_37435,N_36913,N_36887);
nor U37436 (N_37436,N_36904,N_36798);
or U37437 (N_37437,N_36919,N_36761);
xor U37438 (N_37438,N_36986,N_36979);
xnor U37439 (N_37439,N_36873,N_36646);
nand U37440 (N_37440,N_36692,N_36527);
nor U37441 (N_37441,N_36671,N_36527);
xor U37442 (N_37442,N_36591,N_36800);
nand U37443 (N_37443,N_36687,N_36821);
xnor U37444 (N_37444,N_36736,N_36585);
and U37445 (N_37445,N_36883,N_36978);
xor U37446 (N_37446,N_36565,N_36631);
or U37447 (N_37447,N_36511,N_36873);
nor U37448 (N_37448,N_36804,N_36974);
and U37449 (N_37449,N_36541,N_36604);
or U37450 (N_37450,N_36580,N_36555);
nor U37451 (N_37451,N_36896,N_36555);
xnor U37452 (N_37452,N_36827,N_36615);
nor U37453 (N_37453,N_36576,N_36562);
xnor U37454 (N_37454,N_36785,N_36759);
nor U37455 (N_37455,N_36758,N_36869);
nor U37456 (N_37456,N_36801,N_36647);
nand U37457 (N_37457,N_36881,N_36606);
xnor U37458 (N_37458,N_36536,N_36558);
or U37459 (N_37459,N_36699,N_36580);
nand U37460 (N_37460,N_36876,N_36544);
and U37461 (N_37461,N_36556,N_36648);
nand U37462 (N_37462,N_36725,N_36937);
or U37463 (N_37463,N_36897,N_36716);
or U37464 (N_37464,N_36768,N_36600);
nand U37465 (N_37465,N_36889,N_36501);
nor U37466 (N_37466,N_36558,N_36766);
nor U37467 (N_37467,N_36961,N_36916);
or U37468 (N_37468,N_36881,N_36529);
xor U37469 (N_37469,N_36885,N_36604);
xor U37470 (N_37470,N_36685,N_36714);
and U37471 (N_37471,N_36531,N_36834);
and U37472 (N_37472,N_36726,N_36850);
nor U37473 (N_37473,N_36502,N_36832);
nor U37474 (N_37474,N_36913,N_36935);
and U37475 (N_37475,N_36812,N_36975);
and U37476 (N_37476,N_36517,N_36505);
nand U37477 (N_37477,N_36810,N_36769);
and U37478 (N_37478,N_36983,N_36841);
nor U37479 (N_37479,N_36592,N_36700);
nand U37480 (N_37480,N_36587,N_36679);
nand U37481 (N_37481,N_36766,N_36810);
xnor U37482 (N_37482,N_36674,N_36742);
or U37483 (N_37483,N_36958,N_36601);
nand U37484 (N_37484,N_36815,N_36624);
nor U37485 (N_37485,N_36767,N_36919);
nand U37486 (N_37486,N_36821,N_36640);
nand U37487 (N_37487,N_36927,N_36670);
nor U37488 (N_37488,N_36929,N_36854);
xnor U37489 (N_37489,N_36760,N_36615);
nor U37490 (N_37490,N_36909,N_36858);
and U37491 (N_37491,N_36828,N_36985);
nand U37492 (N_37492,N_36865,N_36709);
or U37493 (N_37493,N_36629,N_36746);
or U37494 (N_37494,N_36677,N_36937);
and U37495 (N_37495,N_36952,N_36506);
or U37496 (N_37496,N_36772,N_36727);
nor U37497 (N_37497,N_36749,N_36715);
and U37498 (N_37498,N_36538,N_36710);
nor U37499 (N_37499,N_36639,N_36986);
or U37500 (N_37500,N_37173,N_37207);
xor U37501 (N_37501,N_37301,N_37454);
and U37502 (N_37502,N_37345,N_37441);
and U37503 (N_37503,N_37304,N_37372);
nand U37504 (N_37504,N_37434,N_37370);
and U37505 (N_37505,N_37340,N_37059);
nor U37506 (N_37506,N_37338,N_37130);
xnor U37507 (N_37507,N_37373,N_37410);
nor U37508 (N_37508,N_37228,N_37122);
nand U37509 (N_37509,N_37254,N_37295);
xor U37510 (N_37510,N_37077,N_37231);
nor U37511 (N_37511,N_37351,N_37405);
and U37512 (N_37512,N_37089,N_37492);
or U37513 (N_37513,N_37150,N_37296);
nor U37514 (N_37514,N_37385,N_37110);
or U37515 (N_37515,N_37083,N_37429);
nand U37516 (N_37516,N_37067,N_37220);
or U37517 (N_37517,N_37195,N_37055);
nor U37518 (N_37518,N_37136,N_37289);
xnor U37519 (N_37519,N_37018,N_37397);
nor U37520 (N_37520,N_37357,N_37411);
nand U37521 (N_37521,N_37256,N_37297);
nor U37522 (N_37522,N_37106,N_37316);
and U37523 (N_37523,N_37347,N_37158);
nor U37524 (N_37524,N_37471,N_37322);
nand U37525 (N_37525,N_37483,N_37148);
or U37526 (N_37526,N_37198,N_37174);
and U37527 (N_37527,N_37327,N_37024);
nor U37528 (N_37528,N_37144,N_37028);
nor U37529 (N_37529,N_37287,N_37336);
or U37530 (N_37530,N_37097,N_37216);
and U37531 (N_37531,N_37082,N_37423);
and U37532 (N_37532,N_37032,N_37152);
xnor U37533 (N_37533,N_37323,N_37470);
xor U37534 (N_37534,N_37466,N_37126);
nand U37535 (N_37535,N_37235,N_37249);
xnor U37536 (N_37536,N_37278,N_37350);
xnor U37537 (N_37537,N_37498,N_37314);
xor U37538 (N_37538,N_37282,N_37246);
and U37539 (N_37539,N_37149,N_37463);
or U37540 (N_37540,N_37214,N_37353);
or U37541 (N_37541,N_37062,N_37046);
or U37542 (N_37542,N_37145,N_37090);
or U37543 (N_37543,N_37000,N_37419);
or U37544 (N_37544,N_37300,N_37459);
and U37545 (N_37545,N_37293,N_37132);
and U37546 (N_37546,N_37180,N_37363);
and U37547 (N_37547,N_37001,N_37412);
nor U37548 (N_37548,N_37076,N_37307);
nor U37549 (N_37549,N_37375,N_37362);
or U37550 (N_37550,N_37212,N_37374);
nand U37551 (N_37551,N_37206,N_37113);
or U37552 (N_37552,N_37036,N_37320);
xnor U37553 (N_37553,N_37217,N_37017);
nand U37554 (N_37554,N_37448,N_37064);
nand U37555 (N_37555,N_37294,N_37175);
nand U37556 (N_37556,N_37050,N_37333);
xnor U37557 (N_37557,N_37467,N_37171);
xor U37558 (N_37558,N_37318,N_37033);
or U37559 (N_37559,N_37183,N_37436);
or U37560 (N_37560,N_37233,N_37119);
xnor U37561 (N_37561,N_37058,N_37066);
nand U37562 (N_37562,N_37496,N_37319);
nor U37563 (N_37563,N_37140,N_37329);
and U37564 (N_37564,N_37427,N_37384);
nand U37565 (N_37565,N_37291,N_37203);
nand U37566 (N_37566,N_37182,N_37081);
or U37567 (N_37567,N_37092,N_37424);
and U37568 (N_37568,N_37383,N_37257);
or U37569 (N_37569,N_37098,N_37103);
nand U37570 (N_37570,N_37049,N_37253);
nor U37571 (N_37571,N_37057,N_37061);
xor U37572 (N_37572,N_37117,N_37490);
nor U37573 (N_37573,N_37073,N_37305);
xnor U37574 (N_37574,N_37236,N_37269);
and U37575 (N_37575,N_37417,N_37400);
nor U37576 (N_37576,N_37187,N_37146);
nand U37577 (N_37577,N_37368,N_37205);
and U37578 (N_37578,N_37393,N_37308);
nor U37579 (N_37579,N_37242,N_37267);
or U37580 (N_37580,N_37121,N_37238);
xnor U37581 (N_37581,N_37151,N_37426);
and U37582 (N_37582,N_37263,N_37312);
nand U37583 (N_37583,N_37356,N_37260);
xnor U37584 (N_37584,N_37035,N_37484);
nand U37585 (N_37585,N_37003,N_37298);
nand U37586 (N_37586,N_37248,N_37041);
and U37587 (N_37587,N_37226,N_37112);
nand U37588 (N_37588,N_37455,N_37200);
nor U37589 (N_37589,N_37131,N_37219);
or U37590 (N_37590,N_37489,N_37355);
nor U37591 (N_37591,N_37288,N_37339);
nor U37592 (N_37592,N_37302,N_37209);
nand U37593 (N_37593,N_37264,N_37255);
or U37594 (N_37594,N_37334,N_37447);
and U37595 (N_37595,N_37086,N_37481);
nor U37596 (N_37596,N_37193,N_37366);
nor U37597 (N_37597,N_37396,N_37284);
and U37598 (N_37598,N_37190,N_37382);
or U37599 (N_37599,N_37252,N_37185);
or U37600 (N_37600,N_37428,N_37007);
xor U37601 (N_37601,N_37052,N_37309);
xor U37602 (N_37602,N_37321,N_37476);
xor U37603 (N_37603,N_37330,N_37364);
nor U37604 (N_37604,N_37387,N_37279);
and U37605 (N_37605,N_37044,N_37240);
nor U37606 (N_37606,N_37197,N_37211);
or U37607 (N_37607,N_37023,N_37078);
nand U37608 (N_37608,N_37127,N_37201);
or U37609 (N_37609,N_37290,N_37361);
and U37610 (N_37610,N_37051,N_37222);
xor U37611 (N_37611,N_37020,N_37072);
nand U37612 (N_37612,N_37486,N_37401);
xor U37613 (N_37613,N_37179,N_37433);
nand U37614 (N_37614,N_37225,N_37299);
nor U37615 (N_37615,N_37389,N_37421);
xnor U37616 (N_37616,N_37194,N_37425);
xor U37617 (N_37617,N_37399,N_37215);
and U37618 (N_37618,N_37039,N_37488);
or U37619 (N_37619,N_37475,N_37019);
xnor U37620 (N_37620,N_37430,N_37065);
and U37621 (N_37621,N_37354,N_37192);
and U37622 (N_37622,N_37349,N_37402);
nor U37623 (N_37623,N_37462,N_37111);
xnor U37624 (N_37624,N_37037,N_37005);
nand U37625 (N_37625,N_37071,N_37080);
nor U37626 (N_37626,N_37138,N_37141);
nor U37627 (N_37627,N_37325,N_37016);
nor U37628 (N_37628,N_37142,N_37162);
and U37629 (N_37629,N_37107,N_37188);
and U37630 (N_37630,N_37348,N_37063);
xnor U37631 (N_37631,N_37164,N_37196);
or U37632 (N_37632,N_37109,N_37497);
and U37633 (N_37633,N_37054,N_37128);
xnor U37634 (N_37634,N_37315,N_37168);
nand U37635 (N_37635,N_37189,N_37084);
nand U37636 (N_37636,N_37208,N_37004);
xor U37637 (N_37637,N_37344,N_37156);
nand U37638 (N_37638,N_37414,N_37123);
nor U37639 (N_37639,N_37465,N_37124);
nor U37640 (N_37640,N_37143,N_37341);
nand U37641 (N_37641,N_37234,N_37438);
xnor U37642 (N_37642,N_37102,N_37440);
nor U37643 (N_37643,N_37139,N_37491);
xnor U37644 (N_37644,N_37224,N_37258);
nor U37645 (N_37645,N_37241,N_37056);
xnor U37646 (N_37646,N_37159,N_37435);
and U37647 (N_37647,N_37025,N_37157);
or U37648 (N_37648,N_37409,N_37464);
or U37649 (N_37649,N_37391,N_37099);
and U37650 (N_37650,N_37457,N_37015);
and U37651 (N_37651,N_37251,N_37358);
and U37652 (N_37652,N_37352,N_37310);
or U37653 (N_37653,N_37229,N_37060);
xor U37654 (N_37654,N_37376,N_37116);
nand U37655 (N_37655,N_37105,N_37034);
nor U37656 (N_37656,N_37259,N_37456);
and U37657 (N_37657,N_37273,N_37413);
nor U37658 (N_37658,N_37276,N_37365);
and U37659 (N_37659,N_37237,N_37311);
and U37660 (N_37660,N_37115,N_37027);
nand U37661 (N_37661,N_37011,N_37094);
xor U37662 (N_37662,N_37335,N_37324);
nand U37663 (N_37663,N_37026,N_37331);
xnor U37664 (N_37664,N_37494,N_37468);
or U37665 (N_37665,N_37085,N_37495);
nand U37666 (N_37666,N_37169,N_37469);
nand U37667 (N_37667,N_37346,N_37479);
xor U37668 (N_37668,N_37445,N_37068);
and U37669 (N_37669,N_37499,N_37227);
nand U37670 (N_37670,N_37271,N_37091);
and U37671 (N_37671,N_37100,N_37461);
nor U37672 (N_37672,N_37332,N_37202);
nor U37673 (N_37673,N_37392,N_37167);
and U37674 (N_37674,N_37022,N_37038);
xnor U37675 (N_37675,N_37474,N_37277);
or U37676 (N_37676,N_37087,N_37006);
nand U37677 (N_37677,N_37047,N_37013);
nand U37678 (N_37678,N_37133,N_37451);
or U37679 (N_37679,N_37453,N_37154);
nand U37680 (N_37680,N_37493,N_37386);
nand U37681 (N_37681,N_37244,N_37303);
xnor U37682 (N_37682,N_37292,N_37118);
or U37683 (N_37683,N_37210,N_37170);
xor U37684 (N_37684,N_37030,N_37012);
nor U37685 (N_37685,N_37280,N_37281);
or U37686 (N_37686,N_37390,N_37270);
nor U37687 (N_37687,N_37101,N_37367);
nor U37688 (N_37688,N_37268,N_37381);
xnor U37689 (N_37689,N_37002,N_37328);
nor U37690 (N_37690,N_37218,N_37165);
xor U37691 (N_37691,N_37415,N_37010);
nand U37692 (N_37692,N_37108,N_37045);
nand U37693 (N_37693,N_37265,N_37250);
and U37694 (N_37694,N_37378,N_37388);
and U37695 (N_37695,N_37221,N_37176);
and U37696 (N_37696,N_37009,N_37342);
xor U37697 (N_37697,N_37135,N_37449);
and U37698 (N_37698,N_37266,N_37443);
nor U37699 (N_37699,N_37371,N_37079);
and U37700 (N_37700,N_37163,N_37137);
and U37701 (N_37701,N_37306,N_37199);
xnor U37702 (N_37702,N_37213,N_37431);
xnor U37703 (N_37703,N_37153,N_37369);
and U37704 (N_37704,N_37048,N_37398);
xor U37705 (N_37705,N_37186,N_37181);
or U37706 (N_37706,N_37272,N_37477);
nand U37707 (N_37707,N_37043,N_37223);
xnor U37708 (N_37708,N_37395,N_37286);
or U37709 (N_37709,N_37008,N_37031);
nor U37710 (N_37710,N_37129,N_37191);
or U37711 (N_37711,N_37093,N_37021);
xor U37712 (N_37712,N_37230,N_37403);
nor U37713 (N_37713,N_37074,N_37343);
and U37714 (N_37714,N_37285,N_37184);
and U37715 (N_37715,N_37095,N_37408);
nand U37716 (N_37716,N_37418,N_37487);
or U37717 (N_37717,N_37239,N_37377);
or U37718 (N_37718,N_37283,N_37014);
xor U37719 (N_37719,N_37446,N_37437);
and U37720 (N_37720,N_37360,N_37379);
xnor U37721 (N_37721,N_37416,N_37029);
or U37722 (N_37722,N_37450,N_37452);
and U37723 (N_37723,N_37439,N_37485);
and U37724 (N_37724,N_37125,N_37478);
or U37725 (N_37725,N_37444,N_37088);
and U37726 (N_37726,N_37359,N_37177);
nand U37727 (N_37727,N_37275,N_37069);
xnor U37728 (N_37728,N_37460,N_37313);
and U37729 (N_37729,N_37161,N_37096);
and U37730 (N_37730,N_37120,N_37245);
xor U37731 (N_37731,N_37204,N_37404);
xor U37732 (N_37732,N_37160,N_37040);
or U37733 (N_37733,N_37172,N_37232);
or U37734 (N_37734,N_37482,N_37247);
xor U37735 (N_37735,N_37104,N_37420);
and U37736 (N_37736,N_37053,N_37380);
and U37737 (N_37737,N_37326,N_37394);
xor U37738 (N_37738,N_37261,N_37042);
nand U37739 (N_37739,N_37114,N_37472);
and U37740 (N_37740,N_37406,N_37155);
nor U37741 (N_37741,N_37480,N_37442);
nand U37742 (N_37742,N_37075,N_37147);
and U37743 (N_37743,N_37274,N_37178);
and U37744 (N_37744,N_37422,N_37317);
or U37745 (N_37745,N_37432,N_37262);
nor U37746 (N_37746,N_37070,N_37407);
nor U37747 (N_37747,N_37458,N_37473);
or U37748 (N_37748,N_37243,N_37166);
nor U37749 (N_37749,N_37134,N_37337);
and U37750 (N_37750,N_37282,N_37078);
nor U37751 (N_37751,N_37193,N_37096);
or U37752 (N_37752,N_37011,N_37389);
xnor U37753 (N_37753,N_37143,N_37274);
nand U37754 (N_37754,N_37204,N_37033);
nor U37755 (N_37755,N_37161,N_37152);
xor U37756 (N_37756,N_37055,N_37177);
or U37757 (N_37757,N_37277,N_37397);
nor U37758 (N_37758,N_37202,N_37412);
xnor U37759 (N_37759,N_37022,N_37148);
xor U37760 (N_37760,N_37014,N_37186);
xor U37761 (N_37761,N_37377,N_37013);
nand U37762 (N_37762,N_37440,N_37354);
xor U37763 (N_37763,N_37335,N_37408);
nand U37764 (N_37764,N_37250,N_37297);
xor U37765 (N_37765,N_37185,N_37322);
or U37766 (N_37766,N_37323,N_37441);
nand U37767 (N_37767,N_37070,N_37414);
or U37768 (N_37768,N_37366,N_37351);
nand U37769 (N_37769,N_37061,N_37060);
and U37770 (N_37770,N_37197,N_37176);
or U37771 (N_37771,N_37436,N_37413);
or U37772 (N_37772,N_37056,N_37270);
nor U37773 (N_37773,N_37203,N_37047);
or U37774 (N_37774,N_37418,N_37286);
nor U37775 (N_37775,N_37084,N_37111);
xor U37776 (N_37776,N_37114,N_37117);
nand U37777 (N_37777,N_37474,N_37114);
and U37778 (N_37778,N_37462,N_37370);
nor U37779 (N_37779,N_37116,N_37396);
and U37780 (N_37780,N_37361,N_37109);
and U37781 (N_37781,N_37400,N_37365);
nand U37782 (N_37782,N_37051,N_37370);
nor U37783 (N_37783,N_37399,N_37385);
nor U37784 (N_37784,N_37499,N_37177);
and U37785 (N_37785,N_37270,N_37398);
xor U37786 (N_37786,N_37223,N_37161);
or U37787 (N_37787,N_37170,N_37035);
and U37788 (N_37788,N_37414,N_37445);
nor U37789 (N_37789,N_37477,N_37334);
or U37790 (N_37790,N_37098,N_37038);
or U37791 (N_37791,N_37445,N_37471);
and U37792 (N_37792,N_37015,N_37460);
xor U37793 (N_37793,N_37174,N_37183);
nor U37794 (N_37794,N_37204,N_37162);
xor U37795 (N_37795,N_37183,N_37384);
or U37796 (N_37796,N_37439,N_37066);
nand U37797 (N_37797,N_37264,N_37085);
xor U37798 (N_37798,N_37407,N_37477);
xor U37799 (N_37799,N_37264,N_37213);
or U37800 (N_37800,N_37376,N_37122);
nor U37801 (N_37801,N_37091,N_37318);
nor U37802 (N_37802,N_37355,N_37434);
nor U37803 (N_37803,N_37347,N_37165);
nor U37804 (N_37804,N_37192,N_37470);
nor U37805 (N_37805,N_37041,N_37105);
xnor U37806 (N_37806,N_37404,N_37330);
or U37807 (N_37807,N_37037,N_37327);
and U37808 (N_37808,N_37091,N_37387);
nand U37809 (N_37809,N_37169,N_37210);
or U37810 (N_37810,N_37346,N_37364);
xnor U37811 (N_37811,N_37369,N_37331);
nor U37812 (N_37812,N_37310,N_37376);
nand U37813 (N_37813,N_37159,N_37276);
or U37814 (N_37814,N_37340,N_37358);
xnor U37815 (N_37815,N_37215,N_37271);
xor U37816 (N_37816,N_37460,N_37205);
xnor U37817 (N_37817,N_37371,N_37281);
nor U37818 (N_37818,N_37042,N_37291);
and U37819 (N_37819,N_37238,N_37070);
nand U37820 (N_37820,N_37091,N_37323);
xnor U37821 (N_37821,N_37237,N_37252);
and U37822 (N_37822,N_37016,N_37033);
xor U37823 (N_37823,N_37210,N_37350);
xnor U37824 (N_37824,N_37140,N_37351);
nand U37825 (N_37825,N_37314,N_37347);
nand U37826 (N_37826,N_37427,N_37432);
xor U37827 (N_37827,N_37438,N_37081);
and U37828 (N_37828,N_37165,N_37328);
xor U37829 (N_37829,N_37451,N_37186);
nor U37830 (N_37830,N_37473,N_37043);
nand U37831 (N_37831,N_37367,N_37080);
nand U37832 (N_37832,N_37427,N_37403);
or U37833 (N_37833,N_37250,N_37275);
nor U37834 (N_37834,N_37254,N_37321);
nand U37835 (N_37835,N_37391,N_37080);
or U37836 (N_37836,N_37142,N_37101);
nand U37837 (N_37837,N_37254,N_37056);
or U37838 (N_37838,N_37468,N_37089);
or U37839 (N_37839,N_37087,N_37435);
or U37840 (N_37840,N_37238,N_37030);
nand U37841 (N_37841,N_37244,N_37294);
or U37842 (N_37842,N_37199,N_37309);
nand U37843 (N_37843,N_37039,N_37018);
and U37844 (N_37844,N_37361,N_37253);
and U37845 (N_37845,N_37308,N_37094);
or U37846 (N_37846,N_37039,N_37209);
and U37847 (N_37847,N_37223,N_37415);
nor U37848 (N_37848,N_37152,N_37020);
and U37849 (N_37849,N_37486,N_37246);
nor U37850 (N_37850,N_37255,N_37116);
and U37851 (N_37851,N_37358,N_37038);
and U37852 (N_37852,N_37348,N_37414);
nor U37853 (N_37853,N_37064,N_37493);
and U37854 (N_37854,N_37104,N_37042);
nand U37855 (N_37855,N_37409,N_37386);
nand U37856 (N_37856,N_37016,N_37232);
nor U37857 (N_37857,N_37089,N_37251);
and U37858 (N_37858,N_37358,N_37094);
nand U37859 (N_37859,N_37367,N_37104);
and U37860 (N_37860,N_37096,N_37055);
nand U37861 (N_37861,N_37456,N_37293);
or U37862 (N_37862,N_37397,N_37291);
and U37863 (N_37863,N_37344,N_37182);
nand U37864 (N_37864,N_37172,N_37252);
xor U37865 (N_37865,N_37192,N_37468);
and U37866 (N_37866,N_37407,N_37020);
or U37867 (N_37867,N_37191,N_37286);
and U37868 (N_37868,N_37148,N_37365);
or U37869 (N_37869,N_37110,N_37249);
xor U37870 (N_37870,N_37027,N_37194);
or U37871 (N_37871,N_37410,N_37159);
or U37872 (N_37872,N_37145,N_37259);
nand U37873 (N_37873,N_37270,N_37285);
nand U37874 (N_37874,N_37383,N_37094);
nor U37875 (N_37875,N_37202,N_37242);
and U37876 (N_37876,N_37456,N_37249);
xnor U37877 (N_37877,N_37225,N_37213);
nand U37878 (N_37878,N_37077,N_37104);
and U37879 (N_37879,N_37188,N_37242);
and U37880 (N_37880,N_37076,N_37441);
nor U37881 (N_37881,N_37492,N_37488);
nor U37882 (N_37882,N_37226,N_37111);
nor U37883 (N_37883,N_37296,N_37052);
nor U37884 (N_37884,N_37292,N_37286);
nor U37885 (N_37885,N_37208,N_37026);
or U37886 (N_37886,N_37412,N_37426);
and U37887 (N_37887,N_37357,N_37002);
and U37888 (N_37888,N_37350,N_37198);
or U37889 (N_37889,N_37209,N_37359);
xor U37890 (N_37890,N_37423,N_37007);
and U37891 (N_37891,N_37273,N_37194);
and U37892 (N_37892,N_37003,N_37380);
and U37893 (N_37893,N_37178,N_37057);
xor U37894 (N_37894,N_37288,N_37489);
nand U37895 (N_37895,N_37141,N_37254);
nand U37896 (N_37896,N_37066,N_37027);
xor U37897 (N_37897,N_37142,N_37391);
and U37898 (N_37898,N_37084,N_37184);
nor U37899 (N_37899,N_37467,N_37140);
or U37900 (N_37900,N_37134,N_37376);
xnor U37901 (N_37901,N_37026,N_37171);
and U37902 (N_37902,N_37444,N_37002);
and U37903 (N_37903,N_37196,N_37305);
nor U37904 (N_37904,N_37428,N_37350);
and U37905 (N_37905,N_37105,N_37147);
and U37906 (N_37906,N_37331,N_37437);
or U37907 (N_37907,N_37037,N_37186);
and U37908 (N_37908,N_37415,N_37452);
nand U37909 (N_37909,N_37487,N_37028);
or U37910 (N_37910,N_37328,N_37345);
and U37911 (N_37911,N_37393,N_37199);
and U37912 (N_37912,N_37292,N_37162);
and U37913 (N_37913,N_37147,N_37024);
nor U37914 (N_37914,N_37246,N_37455);
and U37915 (N_37915,N_37303,N_37258);
or U37916 (N_37916,N_37259,N_37479);
xor U37917 (N_37917,N_37299,N_37059);
nand U37918 (N_37918,N_37227,N_37088);
and U37919 (N_37919,N_37103,N_37418);
nand U37920 (N_37920,N_37032,N_37010);
xor U37921 (N_37921,N_37328,N_37489);
and U37922 (N_37922,N_37457,N_37484);
and U37923 (N_37923,N_37465,N_37449);
nor U37924 (N_37924,N_37382,N_37089);
nor U37925 (N_37925,N_37184,N_37261);
nand U37926 (N_37926,N_37208,N_37420);
xor U37927 (N_37927,N_37365,N_37466);
nor U37928 (N_37928,N_37221,N_37435);
and U37929 (N_37929,N_37244,N_37397);
or U37930 (N_37930,N_37241,N_37423);
nand U37931 (N_37931,N_37102,N_37065);
and U37932 (N_37932,N_37190,N_37449);
and U37933 (N_37933,N_37481,N_37057);
nand U37934 (N_37934,N_37266,N_37364);
and U37935 (N_37935,N_37283,N_37096);
nand U37936 (N_37936,N_37469,N_37161);
and U37937 (N_37937,N_37192,N_37355);
nand U37938 (N_37938,N_37199,N_37215);
xor U37939 (N_37939,N_37000,N_37243);
nand U37940 (N_37940,N_37242,N_37412);
and U37941 (N_37941,N_37432,N_37383);
xnor U37942 (N_37942,N_37062,N_37186);
and U37943 (N_37943,N_37475,N_37173);
nand U37944 (N_37944,N_37070,N_37297);
xnor U37945 (N_37945,N_37187,N_37283);
or U37946 (N_37946,N_37019,N_37303);
nand U37947 (N_37947,N_37373,N_37216);
and U37948 (N_37948,N_37331,N_37287);
xnor U37949 (N_37949,N_37308,N_37493);
or U37950 (N_37950,N_37303,N_37392);
nand U37951 (N_37951,N_37269,N_37412);
nor U37952 (N_37952,N_37336,N_37400);
nor U37953 (N_37953,N_37287,N_37286);
nor U37954 (N_37954,N_37282,N_37080);
and U37955 (N_37955,N_37340,N_37490);
and U37956 (N_37956,N_37288,N_37481);
xor U37957 (N_37957,N_37199,N_37197);
nand U37958 (N_37958,N_37476,N_37292);
nor U37959 (N_37959,N_37397,N_37469);
nor U37960 (N_37960,N_37127,N_37200);
nor U37961 (N_37961,N_37238,N_37211);
or U37962 (N_37962,N_37243,N_37290);
or U37963 (N_37963,N_37155,N_37144);
nor U37964 (N_37964,N_37018,N_37068);
or U37965 (N_37965,N_37402,N_37377);
xnor U37966 (N_37966,N_37417,N_37217);
and U37967 (N_37967,N_37192,N_37027);
and U37968 (N_37968,N_37457,N_37418);
xor U37969 (N_37969,N_37234,N_37317);
xnor U37970 (N_37970,N_37471,N_37047);
and U37971 (N_37971,N_37438,N_37498);
and U37972 (N_37972,N_37000,N_37344);
or U37973 (N_37973,N_37196,N_37263);
nor U37974 (N_37974,N_37076,N_37044);
and U37975 (N_37975,N_37003,N_37276);
or U37976 (N_37976,N_37041,N_37489);
nand U37977 (N_37977,N_37342,N_37432);
xnor U37978 (N_37978,N_37322,N_37189);
nor U37979 (N_37979,N_37436,N_37381);
xnor U37980 (N_37980,N_37153,N_37358);
and U37981 (N_37981,N_37035,N_37090);
nand U37982 (N_37982,N_37192,N_37106);
xor U37983 (N_37983,N_37317,N_37122);
nor U37984 (N_37984,N_37494,N_37436);
nand U37985 (N_37985,N_37067,N_37335);
and U37986 (N_37986,N_37467,N_37200);
nand U37987 (N_37987,N_37251,N_37354);
or U37988 (N_37988,N_37429,N_37492);
nand U37989 (N_37989,N_37436,N_37123);
and U37990 (N_37990,N_37367,N_37496);
nand U37991 (N_37991,N_37436,N_37082);
xor U37992 (N_37992,N_37331,N_37127);
nor U37993 (N_37993,N_37046,N_37435);
nor U37994 (N_37994,N_37162,N_37210);
nor U37995 (N_37995,N_37053,N_37196);
xnor U37996 (N_37996,N_37417,N_37357);
nand U37997 (N_37997,N_37018,N_37247);
nand U37998 (N_37998,N_37076,N_37203);
xor U37999 (N_37999,N_37479,N_37222);
or U38000 (N_38000,N_37908,N_37970);
nand U38001 (N_38001,N_37729,N_37631);
xor U38002 (N_38002,N_37515,N_37888);
and U38003 (N_38003,N_37846,N_37946);
xnor U38004 (N_38004,N_37579,N_37815);
xnor U38005 (N_38005,N_37980,N_37576);
or U38006 (N_38006,N_37606,N_37770);
nand U38007 (N_38007,N_37852,N_37581);
nand U38008 (N_38008,N_37660,N_37706);
and U38009 (N_38009,N_37819,N_37904);
xor U38010 (N_38010,N_37552,N_37509);
xor U38011 (N_38011,N_37664,N_37793);
nand U38012 (N_38012,N_37988,N_37855);
nand U38013 (N_38013,N_37713,N_37847);
xor U38014 (N_38014,N_37716,N_37944);
nor U38015 (N_38015,N_37835,N_37511);
nand U38016 (N_38016,N_37865,N_37635);
xor U38017 (N_38017,N_37799,N_37566);
nor U38018 (N_38018,N_37621,N_37694);
nand U38019 (N_38019,N_37754,N_37648);
or U38020 (N_38020,N_37913,N_37957);
nand U38021 (N_38021,N_37531,N_37707);
xor U38022 (N_38022,N_37671,N_37973);
xnor U38023 (N_38023,N_37705,N_37662);
nor U38024 (N_38024,N_37678,N_37998);
and U38025 (N_38025,N_37501,N_37889);
nor U38026 (N_38026,N_37887,N_37996);
nor U38027 (N_38027,N_37500,N_37876);
xnor U38028 (N_38028,N_37895,N_37561);
or U38029 (N_38029,N_37569,N_37696);
nand U38030 (N_38030,N_37986,N_37801);
nor U38031 (N_38031,N_37702,N_37931);
and U38032 (N_38032,N_37939,N_37935);
xor U38033 (N_38033,N_37984,N_37994);
or U38034 (N_38034,N_37872,N_37622);
or U38035 (N_38035,N_37937,N_37730);
or U38036 (N_38036,N_37650,N_37845);
xnor U38037 (N_38037,N_37590,N_37892);
xor U38038 (N_38038,N_37536,N_37616);
nand U38039 (N_38039,N_37744,N_37894);
nand U38040 (N_38040,N_37504,N_37543);
nor U38041 (N_38041,N_37684,N_37874);
nand U38042 (N_38042,N_37859,N_37585);
nand U38043 (N_38043,N_37764,N_37637);
and U38044 (N_38044,N_37964,N_37682);
nor U38045 (N_38045,N_37991,N_37580);
nor U38046 (N_38046,N_37703,N_37817);
nor U38047 (N_38047,N_37783,N_37936);
nor U38048 (N_38048,N_37724,N_37958);
and U38049 (N_38049,N_37735,N_37748);
and U38050 (N_38050,N_37655,N_37794);
nor U38051 (N_38051,N_37787,N_37586);
nor U38052 (N_38052,N_37797,N_37634);
and U38053 (N_38053,N_37761,N_37919);
nor U38054 (N_38054,N_37971,N_37915);
or U38055 (N_38055,N_37989,N_37731);
or U38056 (N_38056,N_37686,N_37699);
or U38057 (N_38057,N_37942,N_37689);
nor U38058 (N_38058,N_37860,N_37920);
or U38059 (N_38059,N_37567,N_37784);
nor U38060 (N_38060,N_37961,N_37921);
and U38061 (N_38061,N_37505,N_37548);
and U38062 (N_38062,N_37965,N_37547);
nor U38063 (N_38063,N_37844,N_37882);
xor U38064 (N_38064,N_37727,N_37644);
nand U38065 (N_38065,N_37698,N_37966);
nand U38066 (N_38066,N_37858,N_37862);
nor U38067 (N_38067,N_37987,N_37571);
and U38068 (N_38068,N_37837,N_37612);
or U38069 (N_38069,N_37832,N_37667);
xnor U38070 (N_38070,N_37791,N_37756);
nor U38071 (N_38071,N_37927,N_37789);
or U38072 (N_38072,N_37781,N_37593);
xor U38073 (N_38073,N_37544,N_37546);
nand U38074 (N_38074,N_37573,N_37578);
xor U38075 (N_38075,N_37800,N_37778);
nand U38076 (N_38076,N_37641,N_37757);
and U38077 (N_38077,N_37681,N_37992);
xor U38078 (N_38078,N_37891,N_37721);
nand U38079 (N_38079,N_37540,N_37897);
xnor U38080 (N_38080,N_37595,N_37691);
nor U38081 (N_38081,N_37912,N_37582);
xnor U38082 (N_38082,N_37527,N_37945);
and U38083 (N_38083,N_37602,N_37905);
nor U38084 (N_38084,N_37674,N_37866);
xor U38085 (N_38085,N_37629,N_37873);
nand U38086 (N_38086,N_37558,N_37893);
xnor U38087 (N_38087,N_37976,N_37584);
and U38088 (N_38088,N_37842,N_37722);
or U38089 (N_38089,N_37529,N_37753);
nor U38090 (N_38090,N_37823,N_37768);
nor U38091 (N_38091,N_37867,N_37652);
xnor U38092 (N_38092,N_37709,N_37983);
nor U38093 (N_38093,N_37712,N_37725);
and U38094 (N_38094,N_37693,N_37922);
xor U38095 (N_38095,N_37740,N_37816);
and U38096 (N_38096,N_37899,N_37656);
and U38097 (N_38097,N_37902,N_37843);
nand U38098 (N_38098,N_37881,N_37790);
nand U38099 (N_38099,N_37940,N_37508);
or U38100 (N_38100,N_37788,N_37930);
and U38101 (N_38101,N_37517,N_37972);
and U38102 (N_38102,N_37545,N_37520);
nor U38103 (N_38103,N_37525,N_37951);
xor U38104 (N_38104,N_37750,N_37538);
xor U38105 (N_38105,N_37625,N_37745);
or U38106 (N_38106,N_37550,N_37617);
nor U38107 (N_38107,N_37985,N_37642);
xnor U38108 (N_38108,N_37636,N_37568);
xnor U38109 (N_38109,N_37555,N_37795);
and U38110 (N_38110,N_37959,N_37836);
or U38111 (N_38111,N_37510,N_37723);
nand U38112 (N_38112,N_37798,N_37995);
xnor U38113 (N_38113,N_37771,N_37752);
nor U38114 (N_38114,N_37755,N_37743);
nor U38115 (N_38115,N_37763,N_37609);
xor U38116 (N_38116,N_37717,N_37896);
nor U38117 (N_38117,N_37982,N_37933);
or U38118 (N_38118,N_37647,N_37524);
or U38119 (N_38119,N_37890,N_37901);
nand U38120 (N_38120,N_37767,N_37979);
nor U38121 (N_38121,N_37878,N_37523);
nand U38122 (N_38122,N_37539,N_37619);
and U38123 (N_38123,N_37848,N_37687);
xnor U38124 (N_38124,N_37695,N_37954);
or U38125 (N_38125,N_37626,N_37557);
xnor U38126 (N_38126,N_37728,N_37572);
and U38127 (N_38127,N_37906,N_37804);
or U38128 (N_38128,N_37683,N_37513);
and U38129 (N_38129,N_37720,N_37685);
and U38130 (N_38130,N_37840,N_37828);
or U38131 (N_38131,N_37738,N_37575);
and U38132 (N_38132,N_37620,N_37911);
nand U38133 (N_38133,N_37741,N_37649);
nand U38134 (N_38134,N_37657,N_37646);
or U38135 (N_38135,N_37627,N_37903);
xnor U38136 (N_38136,N_37814,N_37885);
nand U38137 (N_38137,N_37688,N_37950);
and U38138 (N_38138,N_37948,N_37632);
or U38139 (N_38139,N_37680,N_37811);
or U38140 (N_38140,N_37556,N_37588);
and U38141 (N_38141,N_37537,N_37956);
and U38142 (N_38142,N_37551,N_37775);
and U38143 (N_38143,N_37653,N_37938);
nand U38144 (N_38144,N_37506,N_37810);
xnor U38145 (N_38145,N_37603,N_37955);
or U38146 (N_38146,N_37564,N_37661);
and U38147 (N_38147,N_37943,N_37864);
and U38148 (N_38148,N_37565,N_37673);
nor U38149 (N_38149,N_37628,N_37960);
nor U38150 (N_38150,N_37676,N_37630);
xor U38151 (N_38151,N_37883,N_37813);
and U38152 (N_38152,N_37596,N_37997);
xor U38153 (N_38153,N_37766,N_37762);
xor U38154 (N_38154,N_37774,N_37592);
or U38155 (N_38155,N_37553,N_37507);
nand U38156 (N_38156,N_37559,N_37926);
xor U38157 (N_38157,N_37697,N_37670);
or U38158 (N_38158,N_37675,N_37715);
and U38159 (N_38159,N_37963,N_37850);
xor U38160 (N_38160,N_37822,N_37786);
and U38161 (N_38161,N_37726,N_37877);
or U38162 (N_38162,N_37639,N_37577);
nand U38163 (N_38163,N_37829,N_37521);
nor U38164 (N_38164,N_37809,N_37884);
and U38165 (N_38165,N_37993,N_37962);
xnor U38166 (N_38166,N_37607,N_37777);
nor U38167 (N_38167,N_37776,N_37928);
xnor U38168 (N_38168,N_37785,N_37554);
nand U38169 (N_38169,N_37708,N_37796);
or U38170 (N_38170,N_37853,N_37880);
and U38171 (N_38171,N_37838,N_37665);
and U38172 (N_38172,N_37929,N_37854);
nor U38173 (N_38173,N_37604,N_37526);
nor U38174 (N_38174,N_37780,N_37967);
and U38175 (N_38175,N_37917,N_37714);
nand U38176 (N_38176,N_37643,N_37668);
nand U38177 (N_38177,N_37802,N_37666);
nor U38178 (N_38178,N_37583,N_37969);
nand U38179 (N_38179,N_37711,N_37734);
nand U38180 (N_38180,N_37907,N_37749);
or U38181 (N_38181,N_37949,N_37613);
nor U38182 (N_38182,N_37990,N_37841);
xnor U38183 (N_38183,N_37923,N_37690);
xor U38184 (N_38184,N_37947,N_37542);
and U38185 (N_38185,N_37773,N_37645);
or U38186 (N_38186,N_37746,N_37514);
or U38187 (N_38187,N_37700,N_37677);
and U38188 (N_38188,N_37719,N_37910);
xor U38189 (N_38189,N_37792,N_37615);
and U38190 (N_38190,N_37751,N_37679);
xnor U38191 (N_38191,N_37704,N_37618);
and U38192 (N_38192,N_37608,N_37808);
and U38193 (N_38193,N_37638,N_37654);
and U38194 (N_38194,N_37502,N_37601);
or U38195 (N_38195,N_37863,N_37570);
and U38196 (N_38196,N_37710,N_37516);
and U38197 (N_38197,N_37759,N_37701);
xnor U38198 (N_38198,N_37599,N_37534);
nor U38199 (N_38199,N_37782,N_37530);
and U38200 (N_38200,N_37772,N_37818);
or U38201 (N_38201,N_37924,N_37739);
nand U38202 (N_38202,N_37623,N_37941);
or U38203 (N_38203,N_37918,N_37736);
xnor U38204 (N_38204,N_37925,N_37598);
and U38205 (N_38205,N_37857,N_37820);
nand U38206 (N_38206,N_37591,N_37732);
xnor U38207 (N_38207,N_37589,N_37977);
and U38208 (N_38208,N_37600,N_37806);
xnor U38209 (N_38209,N_37742,N_37856);
nand U38210 (N_38210,N_37574,N_37834);
xor U38211 (N_38211,N_37562,N_37541);
nor U38212 (N_38212,N_37512,N_37851);
nor U38213 (N_38213,N_37968,N_37861);
xnor U38214 (N_38214,N_37805,N_37981);
nand U38215 (N_38215,N_37914,N_37886);
nor U38216 (N_38216,N_37605,N_37839);
and U38217 (N_38217,N_37898,N_37932);
nand U38218 (N_38218,N_37765,N_37952);
and U38219 (N_38219,N_37779,N_37831);
and U38220 (N_38220,N_37651,N_37663);
nor U38221 (N_38221,N_37830,N_37672);
and U38222 (N_38222,N_37934,N_37827);
and U38223 (N_38223,N_37760,N_37871);
nand U38224 (N_38224,N_37812,N_37519);
xnor U38225 (N_38225,N_37503,N_37587);
and U38226 (N_38226,N_37868,N_37879);
nor U38227 (N_38227,N_37825,N_37611);
xnor U38228 (N_38228,N_37833,N_37535);
xnor U38229 (N_38229,N_37718,N_37597);
or U38230 (N_38230,N_37849,N_37518);
xnor U38231 (N_38231,N_37563,N_37974);
and U38232 (N_38232,N_37533,N_37658);
or U38233 (N_38233,N_37769,N_37624);
nand U38234 (N_38234,N_37633,N_37747);
nand U38235 (N_38235,N_37532,N_37614);
xnor U38236 (N_38236,N_37826,N_37528);
nand U38237 (N_38237,N_37640,N_37999);
xnor U38238 (N_38238,N_37900,N_37870);
nor U38239 (N_38239,N_37560,N_37807);
nand U38240 (N_38240,N_37875,N_37978);
xor U38241 (N_38241,N_37916,N_37522);
nor U38242 (N_38242,N_37758,N_37610);
or U38243 (N_38243,N_37953,N_37659);
and U38244 (N_38244,N_37803,N_37737);
nand U38245 (N_38245,N_37869,N_37669);
or U38246 (N_38246,N_37733,N_37909);
nand U38247 (N_38247,N_37549,N_37824);
xor U38248 (N_38248,N_37975,N_37594);
or U38249 (N_38249,N_37821,N_37692);
xor U38250 (N_38250,N_37637,N_37529);
and U38251 (N_38251,N_37612,N_37698);
xnor U38252 (N_38252,N_37551,N_37874);
xor U38253 (N_38253,N_37976,N_37665);
and U38254 (N_38254,N_37788,N_37970);
nand U38255 (N_38255,N_37854,N_37733);
nand U38256 (N_38256,N_37506,N_37960);
and U38257 (N_38257,N_37732,N_37542);
xnor U38258 (N_38258,N_37659,N_37890);
nor U38259 (N_38259,N_37794,N_37780);
or U38260 (N_38260,N_37584,N_37729);
xnor U38261 (N_38261,N_37624,N_37972);
or U38262 (N_38262,N_37682,N_37752);
nand U38263 (N_38263,N_37990,N_37680);
nor U38264 (N_38264,N_37543,N_37540);
nand U38265 (N_38265,N_37706,N_37895);
xnor U38266 (N_38266,N_37577,N_37659);
xor U38267 (N_38267,N_37658,N_37984);
or U38268 (N_38268,N_37686,N_37614);
xor U38269 (N_38269,N_37887,N_37825);
or U38270 (N_38270,N_37937,N_37918);
xor U38271 (N_38271,N_37735,N_37591);
nand U38272 (N_38272,N_37765,N_37520);
nor U38273 (N_38273,N_37653,N_37591);
xnor U38274 (N_38274,N_37671,N_37947);
and U38275 (N_38275,N_37906,N_37695);
nand U38276 (N_38276,N_37674,N_37771);
xor U38277 (N_38277,N_37959,N_37987);
nor U38278 (N_38278,N_37951,N_37605);
and U38279 (N_38279,N_37769,N_37756);
or U38280 (N_38280,N_37983,N_37877);
or U38281 (N_38281,N_37910,N_37523);
or U38282 (N_38282,N_37606,N_37798);
and U38283 (N_38283,N_37767,N_37725);
xor U38284 (N_38284,N_37884,N_37553);
nand U38285 (N_38285,N_37936,N_37672);
and U38286 (N_38286,N_37818,N_37746);
and U38287 (N_38287,N_37924,N_37970);
and U38288 (N_38288,N_37884,N_37952);
and U38289 (N_38289,N_37948,N_37990);
nand U38290 (N_38290,N_37932,N_37952);
and U38291 (N_38291,N_37593,N_37632);
xnor U38292 (N_38292,N_37875,N_37867);
nand U38293 (N_38293,N_37976,N_37996);
nand U38294 (N_38294,N_37772,N_37820);
nor U38295 (N_38295,N_37778,N_37749);
and U38296 (N_38296,N_37831,N_37515);
nor U38297 (N_38297,N_37944,N_37936);
or U38298 (N_38298,N_37972,N_37606);
nand U38299 (N_38299,N_37841,N_37599);
nand U38300 (N_38300,N_37593,N_37908);
nand U38301 (N_38301,N_37991,N_37721);
nor U38302 (N_38302,N_37749,N_37859);
xnor U38303 (N_38303,N_37919,N_37741);
nand U38304 (N_38304,N_37550,N_37763);
nor U38305 (N_38305,N_37836,N_37957);
nand U38306 (N_38306,N_37616,N_37890);
nor U38307 (N_38307,N_37548,N_37859);
and U38308 (N_38308,N_37991,N_37501);
nand U38309 (N_38309,N_37872,N_37921);
xor U38310 (N_38310,N_37819,N_37696);
or U38311 (N_38311,N_37972,N_37623);
or U38312 (N_38312,N_37766,N_37730);
xnor U38313 (N_38313,N_37652,N_37750);
nand U38314 (N_38314,N_37772,N_37504);
nand U38315 (N_38315,N_37745,N_37959);
nor U38316 (N_38316,N_37883,N_37866);
or U38317 (N_38317,N_37998,N_37823);
nand U38318 (N_38318,N_37957,N_37737);
xnor U38319 (N_38319,N_37706,N_37848);
nor U38320 (N_38320,N_37720,N_37729);
or U38321 (N_38321,N_37973,N_37892);
and U38322 (N_38322,N_37504,N_37611);
nand U38323 (N_38323,N_37920,N_37503);
and U38324 (N_38324,N_37988,N_37602);
and U38325 (N_38325,N_37748,N_37526);
or U38326 (N_38326,N_37755,N_37849);
or U38327 (N_38327,N_37881,N_37621);
and U38328 (N_38328,N_37734,N_37586);
or U38329 (N_38329,N_37934,N_37828);
or U38330 (N_38330,N_37575,N_37846);
and U38331 (N_38331,N_37648,N_37625);
nand U38332 (N_38332,N_37627,N_37593);
xor U38333 (N_38333,N_37562,N_37675);
xnor U38334 (N_38334,N_37533,N_37792);
nand U38335 (N_38335,N_37914,N_37847);
xor U38336 (N_38336,N_37746,N_37990);
nand U38337 (N_38337,N_37609,N_37986);
nand U38338 (N_38338,N_37510,N_37816);
or U38339 (N_38339,N_37892,N_37792);
xor U38340 (N_38340,N_37753,N_37912);
or U38341 (N_38341,N_37802,N_37706);
xnor U38342 (N_38342,N_37782,N_37813);
and U38343 (N_38343,N_37651,N_37684);
or U38344 (N_38344,N_37959,N_37591);
xnor U38345 (N_38345,N_37983,N_37672);
nand U38346 (N_38346,N_37660,N_37635);
xor U38347 (N_38347,N_37638,N_37962);
nor U38348 (N_38348,N_37737,N_37671);
or U38349 (N_38349,N_37789,N_37817);
and U38350 (N_38350,N_37786,N_37964);
and U38351 (N_38351,N_37712,N_37651);
nand U38352 (N_38352,N_37643,N_37899);
and U38353 (N_38353,N_37525,N_37693);
xor U38354 (N_38354,N_37981,N_37626);
nor U38355 (N_38355,N_37578,N_37772);
xor U38356 (N_38356,N_37635,N_37891);
nand U38357 (N_38357,N_37671,N_37667);
and U38358 (N_38358,N_37691,N_37784);
nand U38359 (N_38359,N_37673,N_37823);
or U38360 (N_38360,N_37920,N_37717);
or U38361 (N_38361,N_37681,N_37903);
nand U38362 (N_38362,N_37686,N_37517);
xnor U38363 (N_38363,N_37989,N_37839);
or U38364 (N_38364,N_37845,N_37710);
xor U38365 (N_38365,N_37534,N_37823);
nand U38366 (N_38366,N_37986,N_37716);
or U38367 (N_38367,N_37794,N_37791);
or U38368 (N_38368,N_37859,N_37553);
nand U38369 (N_38369,N_37840,N_37816);
nand U38370 (N_38370,N_37759,N_37561);
nand U38371 (N_38371,N_37644,N_37912);
xor U38372 (N_38372,N_37880,N_37944);
nand U38373 (N_38373,N_37684,N_37588);
xnor U38374 (N_38374,N_37959,N_37518);
nor U38375 (N_38375,N_37551,N_37868);
and U38376 (N_38376,N_37901,N_37897);
or U38377 (N_38377,N_37819,N_37642);
or U38378 (N_38378,N_37599,N_37681);
nor U38379 (N_38379,N_37995,N_37672);
and U38380 (N_38380,N_37965,N_37737);
and U38381 (N_38381,N_37899,N_37834);
and U38382 (N_38382,N_37536,N_37622);
xnor U38383 (N_38383,N_37565,N_37678);
and U38384 (N_38384,N_37940,N_37960);
or U38385 (N_38385,N_37504,N_37560);
and U38386 (N_38386,N_37729,N_37593);
nand U38387 (N_38387,N_37991,N_37981);
nand U38388 (N_38388,N_37929,N_37887);
nor U38389 (N_38389,N_37772,N_37661);
or U38390 (N_38390,N_37829,N_37768);
xor U38391 (N_38391,N_37800,N_37537);
and U38392 (N_38392,N_37805,N_37894);
and U38393 (N_38393,N_37990,N_37799);
nor U38394 (N_38394,N_37866,N_37899);
xnor U38395 (N_38395,N_37793,N_37582);
nand U38396 (N_38396,N_37913,N_37625);
or U38397 (N_38397,N_37535,N_37546);
or U38398 (N_38398,N_37847,N_37768);
xnor U38399 (N_38399,N_37914,N_37747);
or U38400 (N_38400,N_37549,N_37837);
or U38401 (N_38401,N_37994,N_37616);
nor U38402 (N_38402,N_37694,N_37717);
nand U38403 (N_38403,N_37875,N_37903);
nor U38404 (N_38404,N_37585,N_37914);
nor U38405 (N_38405,N_37932,N_37742);
or U38406 (N_38406,N_37841,N_37529);
nor U38407 (N_38407,N_37931,N_37576);
or U38408 (N_38408,N_37505,N_37810);
and U38409 (N_38409,N_37819,N_37747);
and U38410 (N_38410,N_37561,N_37709);
xnor U38411 (N_38411,N_37789,N_37522);
and U38412 (N_38412,N_37668,N_37554);
nor U38413 (N_38413,N_37800,N_37713);
nor U38414 (N_38414,N_37911,N_37939);
nand U38415 (N_38415,N_37868,N_37765);
nor U38416 (N_38416,N_37560,N_37676);
or U38417 (N_38417,N_37807,N_37651);
nor U38418 (N_38418,N_37963,N_37526);
xnor U38419 (N_38419,N_37521,N_37512);
or U38420 (N_38420,N_37774,N_37739);
nor U38421 (N_38421,N_37807,N_37721);
or U38422 (N_38422,N_37897,N_37929);
nor U38423 (N_38423,N_37576,N_37815);
nor U38424 (N_38424,N_37611,N_37636);
xnor U38425 (N_38425,N_37720,N_37869);
and U38426 (N_38426,N_37754,N_37904);
xnor U38427 (N_38427,N_37862,N_37722);
and U38428 (N_38428,N_37761,N_37762);
nor U38429 (N_38429,N_37762,N_37959);
nand U38430 (N_38430,N_37793,N_37740);
nor U38431 (N_38431,N_37981,N_37875);
nor U38432 (N_38432,N_37590,N_37721);
xnor U38433 (N_38433,N_37639,N_37607);
nand U38434 (N_38434,N_37844,N_37644);
and U38435 (N_38435,N_37867,N_37813);
and U38436 (N_38436,N_37966,N_37999);
or U38437 (N_38437,N_37925,N_37531);
nand U38438 (N_38438,N_37896,N_37870);
nand U38439 (N_38439,N_37750,N_37764);
nor U38440 (N_38440,N_37620,N_37824);
or U38441 (N_38441,N_37857,N_37702);
and U38442 (N_38442,N_37800,N_37797);
nor U38443 (N_38443,N_37640,N_37507);
nand U38444 (N_38444,N_37983,N_37662);
and U38445 (N_38445,N_37998,N_37633);
nand U38446 (N_38446,N_37901,N_37535);
xor U38447 (N_38447,N_37528,N_37505);
or U38448 (N_38448,N_37897,N_37998);
or U38449 (N_38449,N_37522,N_37853);
and U38450 (N_38450,N_37804,N_37559);
or U38451 (N_38451,N_37922,N_37930);
nor U38452 (N_38452,N_37674,N_37544);
nand U38453 (N_38453,N_37718,N_37816);
nor U38454 (N_38454,N_37617,N_37689);
nand U38455 (N_38455,N_37915,N_37997);
nor U38456 (N_38456,N_37647,N_37907);
xor U38457 (N_38457,N_37859,N_37702);
and U38458 (N_38458,N_37916,N_37917);
and U38459 (N_38459,N_37833,N_37931);
or U38460 (N_38460,N_37813,N_37624);
nor U38461 (N_38461,N_37573,N_37980);
nor U38462 (N_38462,N_37917,N_37841);
nand U38463 (N_38463,N_37525,N_37995);
or U38464 (N_38464,N_37524,N_37917);
xor U38465 (N_38465,N_37752,N_37676);
xnor U38466 (N_38466,N_37534,N_37970);
nor U38467 (N_38467,N_37952,N_37526);
and U38468 (N_38468,N_37738,N_37742);
nor U38469 (N_38469,N_37574,N_37675);
and U38470 (N_38470,N_37612,N_37829);
or U38471 (N_38471,N_37831,N_37889);
xor U38472 (N_38472,N_37618,N_37713);
xor U38473 (N_38473,N_37981,N_37679);
nand U38474 (N_38474,N_37930,N_37844);
or U38475 (N_38475,N_37634,N_37661);
and U38476 (N_38476,N_37977,N_37684);
xnor U38477 (N_38477,N_37810,N_37697);
nor U38478 (N_38478,N_37500,N_37584);
xnor U38479 (N_38479,N_37579,N_37868);
xnor U38480 (N_38480,N_37929,N_37734);
and U38481 (N_38481,N_37871,N_37935);
xnor U38482 (N_38482,N_37647,N_37947);
xor U38483 (N_38483,N_37911,N_37958);
and U38484 (N_38484,N_37946,N_37601);
and U38485 (N_38485,N_37589,N_37633);
nor U38486 (N_38486,N_37606,N_37909);
or U38487 (N_38487,N_37645,N_37801);
xor U38488 (N_38488,N_37692,N_37847);
nor U38489 (N_38489,N_37989,N_37594);
nor U38490 (N_38490,N_37846,N_37954);
nor U38491 (N_38491,N_37965,N_37783);
nor U38492 (N_38492,N_37607,N_37537);
nand U38493 (N_38493,N_37556,N_37819);
nor U38494 (N_38494,N_37816,N_37588);
nand U38495 (N_38495,N_37615,N_37552);
nor U38496 (N_38496,N_37614,N_37631);
or U38497 (N_38497,N_37653,N_37991);
or U38498 (N_38498,N_37515,N_37844);
and U38499 (N_38499,N_37873,N_37551);
nand U38500 (N_38500,N_38002,N_38339);
nor U38501 (N_38501,N_38240,N_38237);
nand U38502 (N_38502,N_38455,N_38005);
and U38503 (N_38503,N_38236,N_38357);
or U38504 (N_38504,N_38088,N_38177);
xnor U38505 (N_38505,N_38018,N_38181);
or U38506 (N_38506,N_38221,N_38130);
nand U38507 (N_38507,N_38450,N_38457);
nor U38508 (N_38508,N_38045,N_38300);
xnor U38509 (N_38509,N_38163,N_38061);
xor U38510 (N_38510,N_38378,N_38128);
and U38511 (N_38511,N_38396,N_38449);
or U38512 (N_38512,N_38171,N_38447);
or U38513 (N_38513,N_38343,N_38229);
and U38514 (N_38514,N_38344,N_38085);
nor U38515 (N_38515,N_38133,N_38150);
nand U38516 (N_38516,N_38208,N_38287);
nand U38517 (N_38517,N_38093,N_38250);
and U38518 (N_38518,N_38188,N_38286);
xor U38519 (N_38519,N_38058,N_38126);
nor U38520 (N_38520,N_38411,N_38044);
xnor U38521 (N_38521,N_38161,N_38244);
or U38522 (N_38522,N_38474,N_38247);
xnor U38523 (N_38523,N_38272,N_38098);
nor U38524 (N_38524,N_38274,N_38360);
or U38525 (N_38525,N_38235,N_38309);
nand U38526 (N_38526,N_38362,N_38347);
xor U38527 (N_38527,N_38155,N_38151);
or U38528 (N_38528,N_38158,N_38209);
nor U38529 (N_38529,N_38011,N_38010);
nor U38530 (N_38530,N_38213,N_38263);
nor U38531 (N_38531,N_38113,N_38284);
and U38532 (N_38532,N_38094,N_38456);
nand U38533 (N_38533,N_38356,N_38030);
nor U38534 (N_38534,N_38086,N_38484);
nor U38535 (N_38535,N_38055,N_38428);
or U38536 (N_38536,N_38111,N_38325);
xnor U38537 (N_38537,N_38215,N_38108);
nand U38538 (N_38538,N_38160,N_38351);
or U38539 (N_38539,N_38063,N_38112);
and U38540 (N_38540,N_38348,N_38006);
and U38541 (N_38541,N_38310,N_38172);
nand U38542 (N_38542,N_38425,N_38073);
or U38543 (N_38543,N_38419,N_38424);
nand U38544 (N_38544,N_38008,N_38053);
and U38545 (N_38545,N_38448,N_38195);
xnor U38546 (N_38546,N_38267,N_38206);
or U38547 (N_38547,N_38222,N_38460);
xnor U38548 (N_38548,N_38436,N_38049);
and U38549 (N_38549,N_38226,N_38337);
or U38550 (N_38550,N_38273,N_38488);
xor U38551 (N_38551,N_38346,N_38101);
nand U38552 (N_38552,N_38083,N_38446);
xnor U38553 (N_38553,N_38296,N_38297);
xor U38554 (N_38554,N_38246,N_38464);
and U38555 (N_38555,N_38153,N_38214);
nand U38556 (N_38556,N_38000,N_38040);
nor U38557 (N_38557,N_38354,N_38389);
nor U38558 (N_38558,N_38034,N_38394);
xnor U38559 (N_38559,N_38127,N_38015);
and U38560 (N_38560,N_38279,N_38418);
xor U38561 (N_38561,N_38462,N_38147);
or U38562 (N_38562,N_38090,N_38285);
and U38563 (N_38563,N_38434,N_38435);
and U38564 (N_38564,N_38048,N_38290);
and U38565 (N_38565,N_38386,N_38335);
nor U38566 (N_38566,N_38084,N_38087);
or U38567 (N_38567,N_38349,N_38097);
or U38568 (N_38568,N_38311,N_38179);
or U38569 (N_38569,N_38019,N_38194);
or U38570 (N_38570,N_38451,N_38072);
nand U38571 (N_38571,N_38490,N_38404);
xor U38572 (N_38572,N_38412,N_38255);
nor U38573 (N_38573,N_38414,N_38099);
or U38574 (N_38574,N_38353,N_38369);
xor U38575 (N_38575,N_38374,N_38121);
nand U38576 (N_38576,N_38124,N_38067);
xor U38577 (N_38577,N_38403,N_38363);
nor U38578 (N_38578,N_38303,N_38117);
xnor U38579 (N_38579,N_38298,N_38134);
and U38580 (N_38580,N_38439,N_38430);
and U38581 (N_38581,N_38184,N_38245);
nor U38582 (N_38582,N_38307,N_38433);
and U38583 (N_38583,N_38050,N_38036);
nand U38584 (N_38584,N_38132,N_38463);
xor U38585 (N_38585,N_38288,N_38407);
nor U38586 (N_38586,N_38452,N_38390);
xnor U38587 (N_38587,N_38069,N_38257);
nand U38588 (N_38588,N_38224,N_38304);
or U38589 (N_38589,N_38413,N_38336);
nor U38590 (N_38590,N_38115,N_38202);
or U38591 (N_38591,N_38092,N_38345);
nor U38592 (N_38592,N_38355,N_38321);
and U38593 (N_38593,N_38327,N_38406);
or U38594 (N_38594,N_38294,N_38114);
nand U38595 (N_38595,N_38201,N_38375);
nand U38596 (N_38596,N_38495,N_38293);
nand U38597 (N_38597,N_38023,N_38021);
xor U38598 (N_38598,N_38468,N_38438);
or U38599 (N_38599,N_38278,N_38170);
or U38600 (N_38600,N_38301,N_38052);
nor U38601 (N_38601,N_38479,N_38079);
xnor U38602 (N_38602,N_38393,N_38059);
or U38603 (N_38603,N_38138,N_38173);
xor U38604 (N_38604,N_38329,N_38361);
or U38605 (N_38605,N_38070,N_38104);
nand U38606 (N_38606,N_38051,N_38024);
and U38607 (N_38607,N_38395,N_38186);
nor U38608 (N_38608,N_38004,N_38441);
or U38609 (N_38609,N_38371,N_38028);
and U38610 (N_38610,N_38308,N_38318);
or U38611 (N_38611,N_38306,N_38164);
xnor U38612 (N_38612,N_38204,N_38074);
and U38613 (N_38613,N_38198,N_38417);
xnor U38614 (N_38614,N_38239,N_38493);
or U38615 (N_38615,N_38109,N_38046);
nor U38616 (N_38616,N_38225,N_38039);
nand U38617 (N_38617,N_38068,N_38313);
nand U38618 (N_38618,N_38333,N_38075);
nand U38619 (N_38619,N_38323,N_38497);
or U38620 (N_38620,N_38217,N_38422);
nand U38621 (N_38621,N_38299,N_38332);
nor U38622 (N_38622,N_38248,N_38210);
or U38623 (N_38623,N_38013,N_38370);
nor U38624 (N_38624,N_38106,N_38107);
xor U38625 (N_38625,N_38496,N_38180);
and U38626 (N_38626,N_38320,N_38489);
and U38627 (N_38627,N_38373,N_38080);
nand U38628 (N_38628,N_38469,N_38189);
xor U38629 (N_38629,N_38388,N_38269);
xor U38630 (N_38630,N_38123,N_38096);
or U38631 (N_38631,N_38277,N_38027);
nand U38632 (N_38632,N_38176,N_38256);
or U38633 (N_38633,N_38182,N_38405);
or U38634 (N_38634,N_38427,N_38183);
or U38635 (N_38635,N_38401,N_38384);
nor U38636 (N_38636,N_38302,N_38228);
nand U38637 (N_38637,N_38319,N_38485);
xnor U38638 (N_38638,N_38031,N_38331);
and U38639 (N_38639,N_38007,N_38081);
nand U38640 (N_38640,N_38017,N_38400);
nand U38641 (N_38641,N_38232,N_38476);
nor U38642 (N_38642,N_38341,N_38342);
or U38643 (N_38643,N_38473,N_38152);
nand U38644 (N_38644,N_38139,N_38038);
xor U38645 (N_38645,N_38076,N_38271);
nor U38646 (N_38646,N_38459,N_38442);
nand U38647 (N_38647,N_38275,N_38233);
xnor U38648 (N_38648,N_38482,N_38242);
xor U38649 (N_38649,N_38416,N_38165);
and U38650 (N_38650,N_38477,N_38431);
and U38651 (N_38651,N_38258,N_38001);
nor U38652 (N_38652,N_38118,N_38056);
nand U38653 (N_38653,N_38366,N_38409);
or U38654 (N_38654,N_38191,N_38199);
nand U38655 (N_38655,N_38408,N_38491);
nor U38656 (N_38656,N_38203,N_38219);
xnor U38657 (N_38657,N_38281,N_38125);
or U38658 (N_38658,N_38499,N_38066);
nand U38659 (N_38659,N_38402,N_38003);
or U38660 (N_38660,N_38316,N_38260);
nand U38661 (N_38661,N_38383,N_38103);
xnor U38662 (N_38662,N_38014,N_38137);
nor U38663 (N_38663,N_38440,N_38078);
nor U38664 (N_38664,N_38033,N_38315);
or U38665 (N_38665,N_38205,N_38157);
or U38666 (N_38666,N_38145,N_38122);
and U38667 (N_38667,N_38196,N_38148);
nand U38668 (N_38668,N_38243,N_38207);
and U38669 (N_38669,N_38057,N_38326);
nand U38670 (N_38670,N_38054,N_38259);
xor U38671 (N_38671,N_38387,N_38314);
nor U38672 (N_38672,N_38095,N_38282);
nor U38673 (N_38673,N_38264,N_38483);
xnor U38674 (N_38674,N_38234,N_38144);
and U38675 (N_38675,N_38365,N_38350);
and U38676 (N_38676,N_38136,N_38494);
nand U38677 (N_38677,N_38283,N_38480);
nor U38678 (N_38678,N_38212,N_38420);
or U38679 (N_38679,N_38091,N_38110);
and U38680 (N_38680,N_38453,N_38487);
or U38681 (N_38681,N_38120,N_38359);
xnor U38682 (N_38682,N_38166,N_38142);
and U38683 (N_38683,N_38398,N_38169);
nand U38684 (N_38684,N_38060,N_38047);
and U38685 (N_38685,N_38478,N_38227);
nor U38686 (N_38686,N_38026,N_38218);
or U38687 (N_38687,N_38042,N_38012);
or U38688 (N_38688,N_38372,N_38379);
or U38689 (N_38689,N_38385,N_38156);
xor U38690 (N_38690,N_38466,N_38223);
nand U38691 (N_38691,N_38249,N_38043);
xnor U38692 (N_38692,N_38364,N_38143);
nor U38693 (N_38693,N_38025,N_38382);
xnor U38694 (N_38694,N_38280,N_38251);
and U38695 (N_38695,N_38035,N_38399);
nand U38696 (N_38696,N_38200,N_38220);
xnor U38697 (N_38697,N_38211,N_38082);
xor U38698 (N_38698,N_38238,N_38131);
nand U38699 (N_38699,N_38322,N_38185);
or U38700 (N_38700,N_38077,N_38432);
xor U38701 (N_38701,N_38089,N_38317);
nor U38702 (N_38702,N_38324,N_38175);
or U38703 (N_38703,N_38254,N_38071);
or U38704 (N_38704,N_38009,N_38437);
nand U38705 (N_38705,N_38178,N_38481);
and U38706 (N_38706,N_38141,N_38498);
xnor U38707 (N_38707,N_38029,N_38190);
and U38708 (N_38708,N_38140,N_38149);
and U38709 (N_38709,N_38197,N_38429);
and U38710 (N_38710,N_38100,N_38116);
nor U38711 (N_38711,N_38340,N_38266);
nand U38712 (N_38712,N_38475,N_38289);
xnor U38713 (N_38713,N_38305,N_38174);
or U38714 (N_38714,N_38065,N_38252);
nand U38715 (N_38715,N_38358,N_38458);
nand U38716 (N_38716,N_38241,N_38270);
or U38717 (N_38717,N_38486,N_38020);
xnor U38718 (N_38718,N_38334,N_38167);
nand U38719 (N_38719,N_38064,N_38470);
xnor U38720 (N_38720,N_38022,N_38410);
and U38721 (N_38721,N_38162,N_38041);
nand U38722 (N_38722,N_38062,N_38102);
nor U38723 (N_38723,N_38380,N_38465);
nor U38724 (N_38724,N_38268,N_38330);
and U38725 (N_38725,N_38216,N_38443);
nand U38726 (N_38726,N_38016,N_38231);
or U38727 (N_38727,N_38135,N_38421);
nor U38728 (N_38728,N_38105,N_38168);
nor U38729 (N_38729,N_38291,N_38261);
or U38730 (N_38730,N_38338,N_38292);
xnor U38731 (N_38731,N_38377,N_38312);
nand U38732 (N_38732,N_38037,N_38262);
nor U38733 (N_38733,N_38454,N_38193);
nand U38734 (N_38734,N_38192,N_38154);
xor U38735 (N_38735,N_38159,N_38423);
xor U38736 (N_38736,N_38328,N_38368);
and U38737 (N_38737,N_38129,N_38187);
xor U38738 (N_38738,N_38392,N_38230);
xnor U38739 (N_38739,N_38472,N_38295);
nand U38740 (N_38740,N_38492,N_38119);
nor U38741 (N_38741,N_38146,N_38376);
or U38742 (N_38742,N_38276,N_38253);
or U38743 (N_38743,N_38391,N_38367);
or U38744 (N_38744,N_38471,N_38352);
nand U38745 (N_38745,N_38444,N_38426);
or U38746 (N_38746,N_38265,N_38445);
and U38747 (N_38747,N_38415,N_38461);
nand U38748 (N_38748,N_38467,N_38397);
xnor U38749 (N_38749,N_38032,N_38381);
xor U38750 (N_38750,N_38469,N_38478);
nand U38751 (N_38751,N_38170,N_38386);
nand U38752 (N_38752,N_38055,N_38440);
or U38753 (N_38753,N_38320,N_38298);
or U38754 (N_38754,N_38067,N_38325);
nor U38755 (N_38755,N_38311,N_38424);
xor U38756 (N_38756,N_38449,N_38183);
nand U38757 (N_38757,N_38434,N_38477);
nand U38758 (N_38758,N_38301,N_38223);
xor U38759 (N_38759,N_38042,N_38347);
or U38760 (N_38760,N_38128,N_38497);
or U38761 (N_38761,N_38148,N_38041);
and U38762 (N_38762,N_38014,N_38226);
xor U38763 (N_38763,N_38197,N_38149);
and U38764 (N_38764,N_38489,N_38100);
nand U38765 (N_38765,N_38275,N_38321);
nor U38766 (N_38766,N_38177,N_38306);
nor U38767 (N_38767,N_38041,N_38199);
nor U38768 (N_38768,N_38013,N_38272);
xor U38769 (N_38769,N_38150,N_38337);
nor U38770 (N_38770,N_38464,N_38275);
and U38771 (N_38771,N_38159,N_38151);
nand U38772 (N_38772,N_38169,N_38023);
nand U38773 (N_38773,N_38296,N_38252);
and U38774 (N_38774,N_38224,N_38111);
nor U38775 (N_38775,N_38234,N_38255);
or U38776 (N_38776,N_38440,N_38135);
xor U38777 (N_38777,N_38368,N_38285);
and U38778 (N_38778,N_38337,N_38115);
xnor U38779 (N_38779,N_38170,N_38178);
and U38780 (N_38780,N_38249,N_38094);
xnor U38781 (N_38781,N_38202,N_38137);
or U38782 (N_38782,N_38261,N_38086);
nand U38783 (N_38783,N_38055,N_38013);
and U38784 (N_38784,N_38153,N_38163);
or U38785 (N_38785,N_38032,N_38418);
xor U38786 (N_38786,N_38256,N_38371);
nand U38787 (N_38787,N_38293,N_38348);
nor U38788 (N_38788,N_38407,N_38037);
xor U38789 (N_38789,N_38358,N_38248);
nor U38790 (N_38790,N_38390,N_38320);
nor U38791 (N_38791,N_38189,N_38288);
xnor U38792 (N_38792,N_38383,N_38388);
and U38793 (N_38793,N_38130,N_38287);
nand U38794 (N_38794,N_38104,N_38015);
nand U38795 (N_38795,N_38205,N_38434);
xor U38796 (N_38796,N_38430,N_38363);
nand U38797 (N_38797,N_38232,N_38339);
nand U38798 (N_38798,N_38144,N_38091);
and U38799 (N_38799,N_38111,N_38298);
nor U38800 (N_38800,N_38277,N_38411);
nor U38801 (N_38801,N_38350,N_38109);
and U38802 (N_38802,N_38293,N_38160);
xnor U38803 (N_38803,N_38474,N_38169);
or U38804 (N_38804,N_38385,N_38487);
or U38805 (N_38805,N_38279,N_38160);
xor U38806 (N_38806,N_38416,N_38024);
nor U38807 (N_38807,N_38450,N_38159);
or U38808 (N_38808,N_38042,N_38368);
nor U38809 (N_38809,N_38301,N_38305);
nor U38810 (N_38810,N_38376,N_38265);
and U38811 (N_38811,N_38487,N_38284);
nor U38812 (N_38812,N_38130,N_38044);
or U38813 (N_38813,N_38202,N_38227);
and U38814 (N_38814,N_38327,N_38050);
nor U38815 (N_38815,N_38103,N_38263);
xor U38816 (N_38816,N_38310,N_38369);
nor U38817 (N_38817,N_38481,N_38067);
nor U38818 (N_38818,N_38439,N_38291);
nand U38819 (N_38819,N_38232,N_38241);
or U38820 (N_38820,N_38408,N_38188);
xor U38821 (N_38821,N_38222,N_38122);
xor U38822 (N_38822,N_38278,N_38028);
and U38823 (N_38823,N_38121,N_38006);
nand U38824 (N_38824,N_38247,N_38256);
nor U38825 (N_38825,N_38368,N_38325);
nand U38826 (N_38826,N_38488,N_38169);
nor U38827 (N_38827,N_38106,N_38226);
and U38828 (N_38828,N_38436,N_38135);
nand U38829 (N_38829,N_38415,N_38200);
and U38830 (N_38830,N_38422,N_38190);
nor U38831 (N_38831,N_38376,N_38359);
or U38832 (N_38832,N_38034,N_38173);
nor U38833 (N_38833,N_38306,N_38206);
or U38834 (N_38834,N_38478,N_38470);
xnor U38835 (N_38835,N_38276,N_38103);
or U38836 (N_38836,N_38264,N_38046);
and U38837 (N_38837,N_38299,N_38340);
nand U38838 (N_38838,N_38019,N_38158);
nand U38839 (N_38839,N_38273,N_38425);
xor U38840 (N_38840,N_38241,N_38361);
and U38841 (N_38841,N_38334,N_38195);
nor U38842 (N_38842,N_38108,N_38084);
or U38843 (N_38843,N_38371,N_38219);
nand U38844 (N_38844,N_38380,N_38320);
nand U38845 (N_38845,N_38051,N_38008);
nor U38846 (N_38846,N_38031,N_38236);
xnor U38847 (N_38847,N_38031,N_38253);
xor U38848 (N_38848,N_38307,N_38440);
and U38849 (N_38849,N_38198,N_38382);
nand U38850 (N_38850,N_38369,N_38211);
and U38851 (N_38851,N_38398,N_38285);
nor U38852 (N_38852,N_38331,N_38468);
nor U38853 (N_38853,N_38043,N_38495);
xnor U38854 (N_38854,N_38224,N_38424);
and U38855 (N_38855,N_38196,N_38118);
or U38856 (N_38856,N_38251,N_38180);
nand U38857 (N_38857,N_38030,N_38488);
nor U38858 (N_38858,N_38355,N_38183);
nor U38859 (N_38859,N_38458,N_38255);
xnor U38860 (N_38860,N_38294,N_38426);
and U38861 (N_38861,N_38057,N_38153);
or U38862 (N_38862,N_38077,N_38429);
xnor U38863 (N_38863,N_38492,N_38424);
and U38864 (N_38864,N_38080,N_38459);
and U38865 (N_38865,N_38225,N_38157);
nor U38866 (N_38866,N_38278,N_38220);
and U38867 (N_38867,N_38010,N_38401);
or U38868 (N_38868,N_38424,N_38283);
nand U38869 (N_38869,N_38358,N_38446);
nor U38870 (N_38870,N_38176,N_38158);
or U38871 (N_38871,N_38234,N_38493);
or U38872 (N_38872,N_38091,N_38220);
nor U38873 (N_38873,N_38053,N_38343);
nor U38874 (N_38874,N_38497,N_38168);
or U38875 (N_38875,N_38047,N_38150);
nor U38876 (N_38876,N_38172,N_38072);
nor U38877 (N_38877,N_38304,N_38235);
and U38878 (N_38878,N_38342,N_38249);
nand U38879 (N_38879,N_38221,N_38264);
nor U38880 (N_38880,N_38404,N_38305);
and U38881 (N_38881,N_38493,N_38411);
nand U38882 (N_38882,N_38451,N_38120);
xor U38883 (N_38883,N_38463,N_38186);
or U38884 (N_38884,N_38340,N_38429);
nor U38885 (N_38885,N_38385,N_38421);
xor U38886 (N_38886,N_38223,N_38096);
nor U38887 (N_38887,N_38390,N_38035);
nor U38888 (N_38888,N_38358,N_38211);
or U38889 (N_38889,N_38018,N_38395);
xnor U38890 (N_38890,N_38455,N_38446);
nand U38891 (N_38891,N_38093,N_38264);
xor U38892 (N_38892,N_38009,N_38499);
or U38893 (N_38893,N_38343,N_38463);
xnor U38894 (N_38894,N_38273,N_38087);
and U38895 (N_38895,N_38291,N_38016);
nand U38896 (N_38896,N_38092,N_38385);
or U38897 (N_38897,N_38060,N_38203);
and U38898 (N_38898,N_38407,N_38045);
nand U38899 (N_38899,N_38094,N_38279);
nand U38900 (N_38900,N_38337,N_38038);
nand U38901 (N_38901,N_38355,N_38328);
or U38902 (N_38902,N_38066,N_38433);
nand U38903 (N_38903,N_38347,N_38471);
xnor U38904 (N_38904,N_38057,N_38140);
nor U38905 (N_38905,N_38249,N_38027);
xnor U38906 (N_38906,N_38124,N_38041);
nand U38907 (N_38907,N_38254,N_38123);
xnor U38908 (N_38908,N_38371,N_38283);
and U38909 (N_38909,N_38044,N_38479);
nand U38910 (N_38910,N_38061,N_38296);
nand U38911 (N_38911,N_38441,N_38226);
or U38912 (N_38912,N_38067,N_38240);
nor U38913 (N_38913,N_38309,N_38269);
xor U38914 (N_38914,N_38337,N_38415);
and U38915 (N_38915,N_38106,N_38463);
nand U38916 (N_38916,N_38173,N_38328);
nand U38917 (N_38917,N_38138,N_38191);
xnor U38918 (N_38918,N_38117,N_38020);
nor U38919 (N_38919,N_38427,N_38353);
nor U38920 (N_38920,N_38459,N_38331);
xor U38921 (N_38921,N_38038,N_38309);
xor U38922 (N_38922,N_38175,N_38095);
or U38923 (N_38923,N_38253,N_38366);
nand U38924 (N_38924,N_38488,N_38021);
nand U38925 (N_38925,N_38013,N_38444);
or U38926 (N_38926,N_38136,N_38251);
or U38927 (N_38927,N_38231,N_38239);
xor U38928 (N_38928,N_38236,N_38104);
xor U38929 (N_38929,N_38438,N_38152);
or U38930 (N_38930,N_38495,N_38408);
nor U38931 (N_38931,N_38067,N_38225);
and U38932 (N_38932,N_38294,N_38234);
xor U38933 (N_38933,N_38169,N_38196);
nor U38934 (N_38934,N_38414,N_38229);
nor U38935 (N_38935,N_38266,N_38311);
or U38936 (N_38936,N_38073,N_38374);
xor U38937 (N_38937,N_38300,N_38018);
nand U38938 (N_38938,N_38152,N_38198);
or U38939 (N_38939,N_38439,N_38141);
or U38940 (N_38940,N_38140,N_38005);
or U38941 (N_38941,N_38409,N_38117);
and U38942 (N_38942,N_38237,N_38496);
nor U38943 (N_38943,N_38251,N_38325);
nand U38944 (N_38944,N_38086,N_38453);
xnor U38945 (N_38945,N_38049,N_38450);
xor U38946 (N_38946,N_38075,N_38458);
or U38947 (N_38947,N_38308,N_38168);
xnor U38948 (N_38948,N_38374,N_38232);
xor U38949 (N_38949,N_38095,N_38461);
nand U38950 (N_38950,N_38191,N_38296);
xnor U38951 (N_38951,N_38406,N_38465);
xor U38952 (N_38952,N_38167,N_38046);
nor U38953 (N_38953,N_38341,N_38172);
or U38954 (N_38954,N_38310,N_38035);
nor U38955 (N_38955,N_38068,N_38021);
and U38956 (N_38956,N_38486,N_38356);
nand U38957 (N_38957,N_38104,N_38067);
xnor U38958 (N_38958,N_38098,N_38152);
xor U38959 (N_38959,N_38498,N_38286);
nand U38960 (N_38960,N_38303,N_38048);
or U38961 (N_38961,N_38040,N_38154);
or U38962 (N_38962,N_38383,N_38286);
nand U38963 (N_38963,N_38097,N_38241);
nand U38964 (N_38964,N_38486,N_38108);
or U38965 (N_38965,N_38295,N_38208);
and U38966 (N_38966,N_38483,N_38381);
xor U38967 (N_38967,N_38105,N_38340);
nand U38968 (N_38968,N_38241,N_38428);
or U38969 (N_38969,N_38348,N_38048);
nor U38970 (N_38970,N_38255,N_38387);
nor U38971 (N_38971,N_38339,N_38469);
nor U38972 (N_38972,N_38153,N_38002);
or U38973 (N_38973,N_38085,N_38413);
and U38974 (N_38974,N_38141,N_38300);
or U38975 (N_38975,N_38424,N_38418);
and U38976 (N_38976,N_38101,N_38096);
and U38977 (N_38977,N_38157,N_38007);
xor U38978 (N_38978,N_38234,N_38247);
nand U38979 (N_38979,N_38490,N_38016);
nor U38980 (N_38980,N_38189,N_38027);
xor U38981 (N_38981,N_38352,N_38388);
nand U38982 (N_38982,N_38131,N_38184);
or U38983 (N_38983,N_38184,N_38141);
and U38984 (N_38984,N_38004,N_38311);
xor U38985 (N_38985,N_38309,N_38462);
or U38986 (N_38986,N_38483,N_38286);
nor U38987 (N_38987,N_38495,N_38429);
nand U38988 (N_38988,N_38424,N_38342);
nand U38989 (N_38989,N_38193,N_38251);
xnor U38990 (N_38990,N_38371,N_38131);
nor U38991 (N_38991,N_38175,N_38079);
nand U38992 (N_38992,N_38378,N_38095);
and U38993 (N_38993,N_38259,N_38442);
and U38994 (N_38994,N_38499,N_38415);
or U38995 (N_38995,N_38344,N_38379);
nor U38996 (N_38996,N_38364,N_38301);
xor U38997 (N_38997,N_38400,N_38499);
nand U38998 (N_38998,N_38331,N_38145);
nand U38999 (N_38999,N_38247,N_38369);
nand U39000 (N_39000,N_38905,N_38744);
xnor U39001 (N_39001,N_38773,N_38544);
nand U39002 (N_39002,N_38872,N_38848);
nand U39003 (N_39003,N_38831,N_38596);
xnor U39004 (N_39004,N_38777,N_38524);
and U39005 (N_39005,N_38623,N_38951);
and U39006 (N_39006,N_38862,N_38709);
nand U39007 (N_39007,N_38741,N_38946);
nor U39008 (N_39008,N_38788,N_38801);
and U39009 (N_39009,N_38804,N_38520);
and U39010 (N_39010,N_38803,N_38707);
nand U39011 (N_39011,N_38641,N_38569);
nand U39012 (N_39012,N_38993,N_38971);
nand U39013 (N_39013,N_38716,N_38949);
and U39014 (N_39014,N_38594,N_38557);
xnor U39015 (N_39015,N_38834,N_38686);
or U39016 (N_39016,N_38600,N_38650);
xnor U39017 (N_39017,N_38964,N_38561);
and U39018 (N_39018,N_38554,N_38677);
nor U39019 (N_39019,N_38536,N_38797);
and U39020 (N_39020,N_38879,N_38620);
nand U39021 (N_39021,N_38713,N_38527);
xor U39022 (N_39022,N_38920,N_38984);
and U39023 (N_39023,N_38525,N_38692);
nand U39024 (N_39024,N_38723,N_38918);
or U39025 (N_39025,N_38756,N_38895);
and U39026 (N_39026,N_38994,N_38990);
xor U39027 (N_39027,N_38719,N_38654);
xor U39028 (N_39028,N_38830,N_38805);
or U39029 (N_39029,N_38588,N_38778);
and U39030 (N_39030,N_38669,N_38806);
nand U39031 (N_39031,N_38921,N_38986);
or U39032 (N_39032,N_38926,N_38816);
or U39033 (N_39033,N_38859,N_38606);
or U39034 (N_39034,N_38568,N_38865);
nor U39035 (N_39035,N_38590,N_38539);
xor U39036 (N_39036,N_38980,N_38891);
nand U39037 (N_39037,N_38663,N_38625);
nand U39038 (N_39038,N_38508,N_38708);
or U39039 (N_39039,N_38972,N_38607);
nand U39040 (N_39040,N_38583,N_38844);
and U39041 (N_39041,N_38978,N_38789);
and U39042 (N_39042,N_38821,N_38861);
or U39043 (N_39043,N_38573,N_38718);
nand U39044 (N_39044,N_38738,N_38792);
nor U39045 (N_39045,N_38802,N_38758);
xor U39046 (N_39046,N_38952,N_38846);
nor U39047 (N_39047,N_38842,N_38944);
and U39048 (N_39048,N_38706,N_38608);
or U39049 (N_39049,N_38874,N_38546);
and U39050 (N_39050,N_38882,N_38725);
nand U39051 (N_39051,N_38769,N_38500);
xnor U39052 (N_39052,N_38940,N_38985);
nand U39053 (N_39053,N_38526,N_38850);
nor U39054 (N_39054,N_38614,N_38515);
xor U39055 (N_39055,N_38914,N_38899);
nor U39056 (N_39056,N_38660,N_38693);
nor U39057 (N_39057,N_38814,N_38701);
xor U39058 (N_39058,N_38688,N_38672);
or U39059 (N_39059,N_38772,N_38668);
xnor U39060 (N_39060,N_38519,N_38950);
and U39061 (N_39061,N_38624,N_38791);
and U39062 (N_39062,N_38687,N_38819);
and U39063 (N_39063,N_38700,N_38784);
nor U39064 (N_39064,N_38617,N_38886);
nand U39065 (N_39065,N_38929,N_38699);
xor U39066 (N_39066,N_38676,N_38566);
or U39067 (N_39067,N_38545,N_38933);
nand U39068 (N_39068,N_38531,N_38832);
nand U39069 (N_39069,N_38960,N_38727);
xor U39070 (N_39070,N_38885,N_38647);
or U39071 (N_39071,N_38549,N_38763);
or U39072 (N_39072,N_38502,N_38551);
and U39073 (N_39073,N_38613,N_38888);
xnor U39074 (N_39074,N_38838,N_38742);
xor U39075 (N_39075,N_38637,N_38749);
nand U39076 (N_39076,N_38825,N_38904);
nand U39077 (N_39077,N_38992,N_38898);
or U39078 (N_39078,N_38796,N_38889);
and U39079 (N_39079,N_38948,N_38565);
and U39080 (N_39080,N_38643,N_38767);
nand U39081 (N_39081,N_38930,N_38998);
and U39082 (N_39082,N_38681,N_38538);
xor U39083 (N_39083,N_38934,N_38667);
and U39084 (N_39084,N_38932,N_38768);
nand U39085 (N_39085,N_38977,N_38562);
and U39086 (N_39086,N_38555,N_38649);
xnor U39087 (N_39087,N_38619,N_38683);
nand U39088 (N_39088,N_38967,N_38774);
and U39089 (N_39089,N_38956,N_38822);
or U39090 (N_39090,N_38799,N_38578);
nand U39091 (N_39091,N_38747,N_38824);
xnor U39092 (N_39092,N_38523,N_38746);
xor U39093 (N_39093,N_38868,N_38794);
xnor U39094 (N_39094,N_38757,N_38981);
or U39095 (N_39095,N_38983,N_38655);
nand U39096 (N_39096,N_38829,N_38552);
or U39097 (N_39097,N_38653,N_38745);
nor U39098 (N_39098,N_38712,N_38532);
and U39099 (N_39099,N_38969,N_38957);
or U39100 (N_39100,N_38908,N_38720);
xor U39101 (N_39101,N_38730,N_38941);
or U39102 (N_39102,N_38919,N_38997);
xor U39103 (N_39103,N_38581,N_38575);
and U39104 (N_39104,N_38864,N_38923);
nand U39105 (N_39105,N_38835,N_38633);
nand U39106 (N_39106,N_38776,N_38710);
nor U39107 (N_39107,N_38953,N_38671);
nor U39108 (N_39108,N_38759,N_38751);
or U39109 (N_39109,N_38942,N_38853);
nand U39110 (N_39110,N_38847,N_38626);
or U39111 (N_39111,N_38656,N_38631);
nand U39112 (N_39112,N_38636,N_38943);
and U39113 (N_39113,N_38947,N_38781);
nand U39114 (N_39114,N_38570,N_38572);
nand U39115 (N_39115,N_38505,N_38585);
or U39116 (N_39116,N_38558,N_38635);
nor U39117 (N_39117,N_38658,N_38764);
nor U39118 (N_39118,N_38839,N_38616);
nand U39119 (N_39119,N_38893,N_38646);
xnor U39120 (N_39120,N_38740,N_38775);
xor U39121 (N_39121,N_38987,N_38996);
and U39122 (N_39122,N_38761,N_38979);
nand U39123 (N_39123,N_38694,N_38779);
or U39124 (N_39124,N_38863,N_38766);
xnor U39125 (N_39125,N_38542,N_38813);
nor U39126 (N_39126,N_38743,N_38582);
nand U39127 (N_39127,N_38610,N_38915);
or U39128 (N_39128,N_38897,N_38703);
or U39129 (N_39129,N_38512,N_38627);
xnor U39130 (N_39130,N_38629,N_38896);
nor U39131 (N_39131,N_38630,N_38628);
or U39132 (N_39132,N_38609,N_38878);
nand U39133 (N_39133,N_38535,N_38715);
nor U39134 (N_39134,N_38876,N_38795);
xor U39135 (N_39135,N_38533,N_38529);
nor U39136 (N_39136,N_38851,N_38711);
or U39137 (N_39137,N_38912,N_38748);
and U39138 (N_39138,N_38737,N_38553);
or U39139 (N_39139,N_38673,N_38679);
nor U39140 (N_39140,N_38843,N_38513);
nand U39141 (N_39141,N_38845,N_38612);
and U39142 (N_39142,N_38511,N_38579);
nor U39143 (N_39143,N_38597,N_38662);
and U39144 (N_39144,N_38503,N_38962);
xor U39145 (N_39145,N_38540,N_38798);
nand U39146 (N_39146,N_38564,N_38659);
xnor U39147 (N_39147,N_38731,N_38982);
xor U39148 (N_39148,N_38753,N_38836);
xnor U39149 (N_39149,N_38808,N_38733);
nand U39150 (N_39150,N_38860,N_38858);
xor U39151 (N_39151,N_38690,N_38890);
xnor U39152 (N_39152,N_38622,N_38705);
or U39153 (N_39153,N_38675,N_38563);
xnor U39154 (N_39154,N_38697,N_38543);
nand U39155 (N_39155,N_38598,N_38724);
xor U39156 (N_39156,N_38674,N_38680);
and U39157 (N_39157,N_38604,N_38632);
and U39158 (N_39158,N_38556,N_38909);
nand U39159 (N_39159,N_38516,N_38867);
xnor U39160 (N_39160,N_38823,N_38849);
nand U39161 (N_39161,N_38547,N_38782);
or U39162 (N_39162,N_38639,N_38841);
xnor U39163 (N_39163,N_38871,N_38939);
xor U39164 (N_39164,N_38593,N_38935);
and U39165 (N_39165,N_38786,N_38765);
nand U39166 (N_39166,N_38780,N_38811);
nand U39167 (N_39167,N_38910,N_38584);
xor U39168 (N_39168,N_38726,N_38913);
or U39169 (N_39169,N_38602,N_38887);
nand U39170 (N_39170,N_38621,N_38991);
and U39171 (N_39171,N_38855,N_38501);
xnor U39172 (N_39172,N_38518,N_38818);
and U39173 (N_39173,N_38875,N_38685);
or U39174 (N_39174,N_38966,N_38522);
nor U39175 (N_39175,N_38704,N_38592);
xor U39176 (N_39176,N_38638,N_38884);
or U39177 (N_39177,N_38837,N_38587);
nand U39178 (N_39178,N_38927,N_38634);
or U39179 (N_39179,N_38856,N_38810);
nor U39180 (N_39180,N_38812,N_38900);
or U39181 (N_39181,N_38696,N_38541);
nor U39182 (N_39182,N_38534,N_38854);
and U39183 (N_39183,N_38580,N_38877);
nand U39184 (N_39184,N_38517,N_38973);
nor U39185 (N_39185,N_38873,N_38665);
and U39186 (N_39186,N_38754,N_38907);
and U39187 (N_39187,N_38640,N_38787);
xnor U39188 (N_39188,N_38928,N_38734);
nand U39189 (N_39189,N_38974,N_38828);
nand U39190 (N_39190,N_38793,N_38601);
xor U39191 (N_39191,N_38722,N_38682);
and U39192 (N_39192,N_38651,N_38894);
nand U39193 (N_39193,N_38881,N_38783);
nor U39194 (N_39194,N_38611,N_38755);
nand U39195 (N_39195,N_38510,N_38857);
xnor U39196 (N_39196,N_38975,N_38702);
nor U39197 (N_39197,N_38728,N_38615);
nor U39198 (N_39198,N_38550,N_38917);
nand U39199 (N_39199,N_38903,N_38937);
xor U39200 (N_39200,N_38714,N_38931);
and U39201 (N_39201,N_38559,N_38506);
nand U39202 (N_39202,N_38807,N_38901);
or U39203 (N_39203,N_38732,N_38827);
and U39204 (N_39204,N_38833,N_38880);
or U39205 (N_39205,N_38976,N_38883);
xor U39206 (N_39206,N_38902,N_38968);
xnor U39207 (N_39207,N_38691,N_38852);
and U39208 (N_39208,N_38869,N_38695);
xor U39209 (N_39209,N_38739,N_38605);
xnor U39210 (N_39210,N_38970,N_38925);
xor U39211 (N_39211,N_38574,N_38790);
or U39212 (N_39212,N_38999,N_38892);
nor U39213 (N_39213,N_38938,N_38995);
nand U39214 (N_39214,N_38586,N_38771);
nor U39215 (N_39215,N_38595,N_38664);
nor U39216 (N_39216,N_38954,N_38760);
nand U39217 (N_39217,N_38817,N_38911);
nor U39218 (N_39218,N_38752,N_38652);
or U39219 (N_39219,N_38698,N_38840);
nand U39220 (N_39220,N_38618,N_38815);
nor U39221 (N_39221,N_38762,N_38521);
nand U39222 (N_39222,N_38567,N_38729);
and U39223 (N_39223,N_38800,N_38571);
or U39224 (N_39224,N_38989,N_38963);
nand U39225 (N_39225,N_38750,N_38644);
and U39226 (N_39226,N_38530,N_38870);
xor U39227 (N_39227,N_38645,N_38678);
nor U39228 (N_39228,N_38603,N_38589);
nor U39229 (N_39229,N_38689,N_38577);
nor U39230 (N_39230,N_38826,N_38560);
nor U39231 (N_39231,N_38936,N_38736);
xnor U39232 (N_39232,N_38965,N_38528);
nand U39233 (N_39233,N_38770,N_38721);
nor U39234 (N_39234,N_38958,N_38670);
and U39235 (N_39235,N_38537,N_38955);
nand U39236 (N_39236,N_38988,N_38548);
nand U39237 (N_39237,N_38666,N_38924);
xnor U39238 (N_39238,N_38906,N_38507);
nand U39239 (N_39239,N_38504,N_38648);
nand U39240 (N_39240,N_38642,N_38591);
or U39241 (N_39241,N_38785,N_38509);
nor U39242 (N_39242,N_38661,N_38916);
or U39243 (N_39243,N_38809,N_38735);
nand U39244 (N_39244,N_38820,N_38945);
xor U39245 (N_39245,N_38959,N_38866);
or U39246 (N_39246,N_38717,N_38599);
and U39247 (N_39247,N_38961,N_38922);
nor U39248 (N_39248,N_38576,N_38684);
nand U39249 (N_39249,N_38657,N_38514);
nand U39250 (N_39250,N_38610,N_38864);
or U39251 (N_39251,N_38702,N_38562);
xor U39252 (N_39252,N_38916,N_38726);
or U39253 (N_39253,N_38783,N_38704);
nor U39254 (N_39254,N_38586,N_38974);
nor U39255 (N_39255,N_38588,N_38890);
and U39256 (N_39256,N_38688,N_38870);
xor U39257 (N_39257,N_38559,N_38713);
and U39258 (N_39258,N_38960,N_38807);
nor U39259 (N_39259,N_38809,N_38625);
nor U39260 (N_39260,N_38669,N_38919);
or U39261 (N_39261,N_38707,N_38751);
xor U39262 (N_39262,N_38844,N_38601);
nor U39263 (N_39263,N_38958,N_38649);
or U39264 (N_39264,N_38976,N_38570);
xnor U39265 (N_39265,N_38779,N_38708);
and U39266 (N_39266,N_38516,N_38514);
or U39267 (N_39267,N_38594,N_38874);
nand U39268 (N_39268,N_38630,N_38762);
xnor U39269 (N_39269,N_38704,N_38910);
nand U39270 (N_39270,N_38600,N_38752);
nand U39271 (N_39271,N_38996,N_38894);
nand U39272 (N_39272,N_38545,N_38881);
and U39273 (N_39273,N_38881,N_38999);
nor U39274 (N_39274,N_38657,N_38539);
nor U39275 (N_39275,N_38650,N_38965);
and U39276 (N_39276,N_38575,N_38969);
nand U39277 (N_39277,N_38714,N_38789);
xnor U39278 (N_39278,N_38968,N_38761);
and U39279 (N_39279,N_38852,N_38932);
nand U39280 (N_39280,N_38544,N_38702);
and U39281 (N_39281,N_38522,N_38686);
nor U39282 (N_39282,N_38588,N_38977);
nand U39283 (N_39283,N_38536,N_38750);
nand U39284 (N_39284,N_38563,N_38526);
or U39285 (N_39285,N_38685,N_38861);
nand U39286 (N_39286,N_38676,N_38835);
xor U39287 (N_39287,N_38623,N_38823);
nand U39288 (N_39288,N_38963,N_38958);
nand U39289 (N_39289,N_38948,N_38663);
nor U39290 (N_39290,N_38722,N_38860);
nand U39291 (N_39291,N_38925,N_38587);
nor U39292 (N_39292,N_38576,N_38991);
and U39293 (N_39293,N_38884,N_38608);
or U39294 (N_39294,N_38737,N_38895);
xnor U39295 (N_39295,N_38924,N_38652);
xor U39296 (N_39296,N_38532,N_38544);
nand U39297 (N_39297,N_38675,N_38731);
or U39298 (N_39298,N_38900,N_38532);
nand U39299 (N_39299,N_38755,N_38662);
or U39300 (N_39300,N_38732,N_38545);
nor U39301 (N_39301,N_38930,N_38661);
or U39302 (N_39302,N_38632,N_38868);
nand U39303 (N_39303,N_38569,N_38514);
and U39304 (N_39304,N_38909,N_38563);
or U39305 (N_39305,N_38670,N_38910);
or U39306 (N_39306,N_38610,N_38978);
or U39307 (N_39307,N_38642,N_38665);
or U39308 (N_39308,N_38600,N_38587);
and U39309 (N_39309,N_38905,N_38750);
nor U39310 (N_39310,N_38854,N_38543);
xnor U39311 (N_39311,N_38861,N_38736);
or U39312 (N_39312,N_38890,N_38844);
nor U39313 (N_39313,N_38877,N_38537);
xor U39314 (N_39314,N_38868,N_38752);
xor U39315 (N_39315,N_38779,N_38731);
or U39316 (N_39316,N_38549,N_38510);
nand U39317 (N_39317,N_38655,N_38678);
nand U39318 (N_39318,N_38977,N_38598);
and U39319 (N_39319,N_38868,N_38905);
and U39320 (N_39320,N_38592,N_38769);
nand U39321 (N_39321,N_38540,N_38796);
xor U39322 (N_39322,N_38971,N_38744);
nand U39323 (N_39323,N_38826,N_38999);
and U39324 (N_39324,N_38672,N_38696);
nand U39325 (N_39325,N_38596,N_38728);
nor U39326 (N_39326,N_38991,N_38716);
or U39327 (N_39327,N_38898,N_38883);
nand U39328 (N_39328,N_38538,N_38631);
nor U39329 (N_39329,N_38981,N_38662);
and U39330 (N_39330,N_38513,N_38981);
nor U39331 (N_39331,N_38528,N_38507);
or U39332 (N_39332,N_38540,N_38760);
nor U39333 (N_39333,N_38719,N_38558);
xor U39334 (N_39334,N_38930,N_38785);
xor U39335 (N_39335,N_38804,N_38741);
nor U39336 (N_39336,N_38544,N_38930);
nor U39337 (N_39337,N_38618,N_38819);
nand U39338 (N_39338,N_38725,N_38973);
nor U39339 (N_39339,N_38825,N_38613);
nand U39340 (N_39340,N_38800,N_38589);
nor U39341 (N_39341,N_38831,N_38709);
xnor U39342 (N_39342,N_38539,N_38661);
xnor U39343 (N_39343,N_38804,N_38589);
or U39344 (N_39344,N_38933,N_38517);
or U39345 (N_39345,N_38618,N_38636);
xor U39346 (N_39346,N_38616,N_38568);
or U39347 (N_39347,N_38909,N_38641);
and U39348 (N_39348,N_38729,N_38781);
or U39349 (N_39349,N_38896,N_38947);
or U39350 (N_39350,N_38534,N_38541);
xor U39351 (N_39351,N_38708,N_38755);
nor U39352 (N_39352,N_38714,N_38593);
and U39353 (N_39353,N_38756,N_38533);
nand U39354 (N_39354,N_38588,N_38801);
xnor U39355 (N_39355,N_38729,N_38790);
nand U39356 (N_39356,N_38951,N_38743);
nand U39357 (N_39357,N_38516,N_38689);
nor U39358 (N_39358,N_38783,N_38607);
nand U39359 (N_39359,N_38855,N_38557);
nand U39360 (N_39360,N_38719,N_38694);
nor U39361 (N_39361,N_38624,N_38658);
nand U39362 (N_39362,N_38554,N_38577);
nand U39363 (N_39363,N_38795,N_38792);
nor U39364 (N_39364,N_38826,N_38677);
and U39365 (N_39365,N_38908,N_38858);
nor U39366 (N_39366,N_38709,N_38879);
xnor U39367 (N_39367,N_38917,N_38541);
nor U39368 (N_39368,N_38515,N_38960);
nand U39369 (N_39369,N_38872,N_38975);
nand U39370 (N_39370,N_38676,N_38631);
and U39371 (N_39371,N_38769,N_38565);
xnor U39372 (N_39372,N_38627,N_38637);
xnor U39373 (N_39373,N_38691,N_38998);
nand U39374 (N_39374,N_38929,N_38997);
or U39375 (N_39375,N_38784,N_38886);
or U39376 (N_39376,N_38543,N_38835);
and U39377 (N_39377,N_38642,N_38879);
nand U39378 (N_39378,N_38778,N_38605);
xnor U39379 (N_39379,N_38511,N_38970);
and U39380 (N_39380,N_38761,N_38584);
nand U39381 (N_39381,N_38800,N_38717);
nand U39382 (N_39382,N_38668,N_38876);
xor U39383 (N_39383,N_38887,N_38996);
nand U39384 (N_39384,N_38584,N_38886);
and U39385 (N_39385,N_38979,N_38854);
xnor U39386 (N_39386,N_38769,N_38826);
xor U39387 (N_39387,N_38854,N_38858);
xnor U39388 (N_39388,N_38547,N_38584);
nand U39389 (N_39389,N_38800,N_38924);
nor U39390 (N_39390,N_38745,N_38518);
nor U39391 (N_39391,N_38662,N_38885);
or U39392 (N_39392,N_38773,N_38665);
xor U39393 (N_39393,N_38691,N_38593);
nand U39394 (N_39394,N_38810,N_38866);
nor U39395 (N_39395,N_38679,N_38544);
and U39396 (N_39396,N_38576,N_38939);
xnor U39397 (N_39397,N_38500,N_38626);
nand U39398 (N_39398,N_38675,N_38918);
xnor U39399 (N_39399,N_38775,N_38895);
nor U39400 (N_39400,N_38736,N_38916);
nand U39401 (N_39401,N_38820,N_38675);
nor U39402 (N_39402,N_38723,N_38939);
and U39403 (N_39403,N_38831,N_38783);
or U39404 (N_39404,N_38558,N_38729);
or U39405 (N_39405,N_38508,N_38651);
or U39406 (N_39406,N_38837,N_38552);
xor U39407 (N_39407,N_38630,N_38886);
nand U39408 (N_39408,N_38546,N_38926);
nand U39409 (N_39409,N_38837,N_38878);
nand U39410 (N_39410,N_38767,N_38783);
nand U39411 (N_39411,N_38984,N_38873);
and U39412 (N_39412,N_38836,N_38981);
and U39413 (N_39413,N_38934,N_38872);
nand U39414 (N_39414,N_38966,N_38973);
or U39415 (N_39415,N_38665,N_38604);
and U39416 (N_39416,N_38689,N_38948);
and U39417 (N_39417,N_38844,N_38805);
xor U39418 (N_39418,N_38661,N_38978);
and U39419 (N_39419,N_38857,N_38552);
xor U39420 (N_39420,N_38787,N_38907);
xor U39421 (N_39421,N_38679,N_38511);
xnor U39422 (N_39422,N_38979,N_38648);
and U39423 (N_39423,N_38734,N_38709);
nor U39424 (N_39424,N_38732,N_38549);
and U39425 (N_39425,N_38899,N_38520);
nor U39426 (N_39426,N_38902,N_38868);
or U39427 (N_39427,N_38525,N_38914);
nor U39428 (N_39428,N_38538,N_38518);
or U39429 (N_39429,N_38963,N_38518);
xor U39430 (N_39430,N_38890,N_38974);
nand U39431 (N_39431,N_38911,N_38819);
or U39432 (N_39432,N_38899,N_38844);
nor U39433 (N_39433,N_38915,N_38829);
xnor U39434 (N_39434,N_38617,N_38558);
or U39435 (N_39435,N_38624,N_38737);
nor U39436 (N_39436,N_38910,N_38920);
nand U39437 (N_39437,N_38738,N_38955);
and U39438 (N_39438,N_38992,N_38513);
and U39439 (N_39439,N_38972,N_38676);
nand U39440 (N_39440,N_38795,N_38581);
and U39441 (N_39441,N_38842,N_38956);
and U39442 (N_39442,N_38991,N_38948);
or U39443 (N_39443,N_38881,N_38915);
nor U39444 (N_39444,N_38615,N_38828);
and U39445 (N_39445,N_38566,N_38654);
and U39446 (N_39446,N_38725,N_38893);
or U39447 (N_39447,N_38796,N_38978);
nor U39448 (N_39448,N_38898,N_38751);
or U39449 (N_39449,N_38533,N_38692);
or U39450 (N_39450,N_38749,N_38705);
nor U39451 (N_39451,N_38898,N_38621);
nor U39452 (N_39452,N_38710,N_38940);
and U39453 (N_39453,N_38523,N_38689);
or U39454 (N_39454,N_38685,N_38891);
nand U39455 (N_39455,N_38728,N_38507);
xnor U39456 (N_39456,N_38506,N_38885);
nand U39457 (N_39457,N_38879,N_38633);
or U39458 (N_39458,N_38945,N_38822);
and U39459 (N_39459,N_38549,N_38595);
and U39460 (N_39460,N_38781,N_38822);
nor U39461 (N_39461,N_38527,N_38654);
xor U39462 (N_39462,N_38531,N_38790);
or U39463 (N_39463,N_38951,N_38702);
or U39464 (N_39464,N_38872,N_38675);
nand U39465 (N_39465,N_38838,N_38788);
nor U39466 (N_39466,N_38816,N_38863);
and U39467 (N_39467,N_38988,N_38819);
and U39468 (N_39468,N_38883,N_38625);
and U39469 (N_39469,N_38611,N_38505);
nor U39470 (N_39470,N_38582,N_38783);
nand U39471 (N_39471,N_38954,N_38600);
nor U39472 (N_39472,N_38504,N_38740);
nor U39473 (N_39473,N_38829,N_38777);
or U39474 (N_39474,N_38918,N_38554);
or U39475 (N_39475,N_38985,N_38616);
and U39476 (N_39476,N_38521,N_38677);
and U39477 (N_39477,N_38928,N_38614);
nand U39478 (N_39478,N_38959,N_38977);
or U39479 (N_39479,N_38764,N_38987);
and U39480 (N_39480,N_38851,N_38681);
nand U39481 (N_39481,N_38997,N_38523);
or U39482 (N_39482,N_38871,N_38932);
nand U39483 (N_39483,N_38770,N_38803);
xnor U39484 (N_39484,N_38834,N_38622);
nand U39485 (N_39485,N_38834,N_38657);
or U39486 (N_39486,N_38772,N_38878);
nor U39487 (N_39487,N_38808,N_38522);
and U39488 (N_39488,N_38679,N_38633);
nand U39489 (N_39489,N_38602,N_38695);
nor U39490 (N_39490,N_38753,N_38959);
and U39491 (N_39491,N_38600,N_38887);
or U39492 (N_39492,N_38707,N_38900);
or U39493 (N_39493,N_38660,N_38998);
or U39494 (N_39494,N_38621,N_38553);
or U39495 (N_39495,N_38928,N_38517);
or U39496 (N_39496,N_38762,N_38786);
or U39497 (N_39497,N_38996,N_38701);
nor U39498 (N_39498,N_38508,N_38747);
and U39499 (N_39499,N_38723,N_38863);
and U39500 (N_39500,N_39177,N_39487);
nand U39501 (N_39501,N_39160,N_39133);
xor U39502 (N_39502,N_39148,N_39123);
and U39503 (N_39503,N_39204,N_39316);
and U39504 (N_39504,N_39292,N_39052);
nand U39505 (N_39505,N_39215,N_39179);
xor U39506 (N_39506,N_39205,N_39285);
and U39507 (N_39507,N_39121,N_39159);
or U39508 (N_39508,N_39327,N_39294);
nand U39509 (N_39509,N_39282,N_39065);
nor U39510 (N_39510,N_39030,N_39266);
or U39511 (N_39511,N_39257,N_39134);
and U39512 (N_39512,N_39132,N_39088);
xor U39513 (N_39513,N_39197,N_39236);
nor U39514 (N_39514,N_39122,N_39259);
nor U39515 (N_39515,N_39361,N_39370);
or U39516 (N_39516,N_39054,N_39142);
and U39517 (N_39517,N_39139,N_39172);
or U39518 (N_39518,N_39375,N_39016);
xor U39519 (N_39519,N_39096,N_39492);
or U39520 (N_39520,N_39004,N_39305);
or U39521 (N_39521,N_39422,N_39064);
nor U39522 (N_39522,N_39042,N_39155);
or U39523 (N_39523,N_39483,N_39077);
xnor U39524 (N_39524,N_39240,N_39312);
or U39525 (N_39525,N_39095,N_39163);
nand U39526 (N_39526,N_39195,N_39250);
xnor U39527 (N_39527,N_39093,N_39329);
and U39528 (N_39528,N_39334,N_39319);
and U39529 (N_39529,N_39317,N_39263);
nor U39530 (N_39530,N_39390,N_39038);
and U39531 (N_39531,N_39265,N_39365);
and U39532 (N_39532,N_39458,N_39276);
and U39533 (N_39533,N_39391,N_39118);
and U39534 (N_39534,N_39033,N_39044);
xnor U39535 (N_39535,N_39482,N_39326);
and U39536 (N_39536,N_39393,N_39268);
or U39537 (N_39537,N_39384,N_39344);
and U39538 (N_39538,N_39014,N_39416);
and U39539 (N_39539,N_39057,N_39046);
and U39540 (N_39540,N_39438,N_39371);
or U39541 (N_39541,N_39070,N_39255);
or U39542 (N_39542,N_39015,N_39075);
xnor U39543 (N_39543,N_39140,N_39481);
and U39544 (N_39544,N_39144,N_39131);
xor U39545 (N_39545,N_39104,N_39418);
and U39546 (N_39546,N_39444,N_39165);
xnor U39547 (N_39547,N_39040,N_39185);
nand U39548 (N_39548,N_39499,N_39314);
nor U39549 (N_39549,N_39380,N_39174);
and U39550 (N_39550,N_39402,N_39494);
and U39551 (N_39551,N_39242,N_39192);
or U39552 (N_39552,N_39382,N_39388);
xor U39553 (N_39553,N_39228,N_39010);
xor U39554 (N_39554,N_39424,N_39290);
xnor U39555 (N_39555,N_39281,N_39022);
or U39556 (N_39556,N_39206,N_39394);
or U39557 (N_39557,N_39201,N_39403);
nor U39558 (N_39558,N_39034,N_39013);
nand U39559 (N_39559,N_39414,N_39287);
or U39560 (N_39560,N_39083,N_39275);
or U39561 (N_39561,N_39099,N_39237);
nor U39562 (N_39562,N_39158,N_39475);
xor U39563 (N_39563,N_39176,N_39182);
xnor U39564 (N_39564,N_39471,N_39293);
and U39565 (N_39565,N_39352,N_39078);
nand U39566 (N_39566,N_39169,N_39145);
nor U39567 (N_39567,N_39254,N_39049);
or U39568 (N_39568,N_39493,N_39067);
or U39569 (N_39569,N_39166,N_39440);
or U39570 (N_39570,N_39028,N_39063);
or U39571 (N_39571,N_39081,N_39048);
nand U39572 (N_39572,N_39366,N_39008);
xor U39573 (N_39573,N_39284,N_39423);
xor U39574 (N_39574,N_39343,N_39200);
nand U39575 (N_39575,N_39468,N_39011);
and U39576 (N_39576,N_39079,N_39459);
xnor U39577 (N_39577,N_39234,N_39225);
or U39578 (N_39578,N_39264,N_39198);
or U39579 (N_39579,N_39066,N_39400);
or U39580 (N_39580,N_39256,N_39445);
nand U39581 (N_39581,N_39338,N_39248);
nand U39582 (N_39582,N_39497,N_39466);
or U39583 (N_39583,N_39358,N_39351);
xnor U39584 (N_39584,N_39452,N_39398);
xor U39585 (N_39585,N_39120,N_39496);
nor U39586 (N_39586,N_39386,N_39367);
nor U39587 (N_39587,N_39359,N_39363);
nand U39588 (N_39588,N_39410,N_39180);
nand U39589 (N_39589,N_39340,N_39495);
and U39590 (N_39590,N_39019,N_39243);
and U39591 (N_39591,N_39100,N_39113);
or U39592 (N_39592,N_39446,N_39269);
or U39593 (N_39593,N_39005,N_39235);
and U39594 (N_39594,N_39267,N_39220);
or U39595 (N_39595,N_39227,N_39062);
or U39596 (N_39596,N_39374,N_39126);
or U39597 (N_39597,N_39056,N_39053);
xnor U39598 (N_39598,N_39125,N_39465);
and U39599 (N_39599,N_39320,N_39238);
and U39600 (N_39600,N_39333,N_39101);
or U39601 (N_39601,N_39190,N_39469);
or U39602 (N_39602,N_39491,N_39301);
and U39603 (N_39603,N_39449,N_39246);
xnor U39604 (N_39604,N_39472,N_39086);
or U39605 (N_39605,N_39325,N_39335);
nand U39606 (N_39606,N_39098,N_39392);
xnor U39607 (N_39607,N_39435,N_39464);
and U39608 (N_39608,N_39110,N_39442);
xnor U39609 (N_39609,N_39141,N_39478);
xnor U39610 (N_39610,N_39232,N_39059);
and U39611 (N_39611,N_39331,N_39203);
xor U39612 (N_39612,N_39194,N_39273);
or U39613 (N_39613,N_39296,N_39262);
and U39614 (N_39614,N_39309,N_39311);
nor U39615 (N_39615,N_39239,N_39337);
xor U39616 (N_39616,N_39007,N_39074);
or U39617 (N_39617,N_39069,N_39420);
and U39618 (N_39618,N_39153,N_39186);
nor U39619 (N_39619,N_39387,N_39330);
or U39620 (N_39620,N_39288,N_39379);
and U39621 (N_39621,N_39318,N_39406);
nand U39622 (N_39622,N_39479,N_39152);
or U39623 (N_39623,N_39085,N_39490);
and U39624 (N_39624,N_39233,N_39486);
xor U39625 (N_39625,N_39043,N_39026);
or U39626 (N_39626,N_39409,N_39241);
nand U39627 (N_39627,N_39024,N_39170);
and U39628 (N_39628,N_39323,N_39023);
nor U39629 (N_39629,N_39084,N_39278);
and U39630 (N_39630,N_39324,N_39451);
xor U39631 (N_39631,N_39137,N_39039);
nand U39632 (N_39632,N_39350,N_39304);
xnor U39633 (N_39633,N_39463,N_39389);
and U39634 (N_39634,N_39209,N_39112);
or U39635 (N_39635,N_39055,N_39457);
xnor U39636 (N_39636,N_39128,N_39157);
or U39637 (N_39637,N_39216,N_39454);
or U39638 (N_39638,N_39230,N_39455);
nand U39639 (N_39639,N_39441,N_39364);
nor U39640 (N_39640,N_39307,N_39087);
nor U39641 (N_39641,N_39031,N_39035);
xor U39642 (N_39642,N_39138,N_39261);
nand U39643 (N_39643,N_39355,N_39461);
nor U39644 (N_39644,N_39002,N_39408);
xor U39645 (N_39645,N_39421,N_39061);
xnor U39646 (N_39646,N_39226,N_39187);
xnor U39647 (N_39647,N_39476,N_39076);
xnor U39648 (N_39648,N_39353,N_39289);
xnor U39649 (N_39649,N_39072,N_39383);
or U39650 (N_39650,N_39328,N_39223);
nor U39651 (N_39651,N_39345,N_39447);
nor U39652 (N_39652,N_39115,N_39467);
and U39653 (N_39653,N_39362,N_39027);
or U39654 (N_39654,N_39191,N_39251);
and U39655 (N_39655,N_39149,N_39025);
and U39656 (N_39656,N_39000,N_39109);
and U39657 (N_39657,N_39274,N_39020);
xnor U39658 (N_39658,N_39017,N_39419);
or U39659 (N_39659,N_39183,N_39181);
xnor U39660 (N_39660,N_39489,N_39147);
and U39661 (N_39661,N_39407,N_39395);
nand U39662 (N_39662,N_39143,N_39193);
and U39663 (N_39663,N_39258,N_39298);
or U39664 (N_39664,N_39051,N_39199);
nand U39665 (N_39665,N_39184,N_39091);
and U39666 (N_39666,N_39006,N_39488);
nor U39667 (N_39667,N_39295,N_39453);
and U39668 (N_39668,N_39302,N_39127);
xor U39669 (N_39669,N_39354,N_39222);
xor U39670 (N_39670,N_39090,N_39041);
or U39671 (N_39671,N_39173,N_39308);
xor U39672 (N_39672,N_39092,N_39474);
or U39673 (N_39673,N_39356,N_39189);
and U39674 (N_39674,N_39080,N_39045);
or U39675 (N_39675,N_39432,N_39217);
nand U39676 (N_39676,N_39150,N_39089);
and U39677 (N_39677,N_39404,N_39135);
or U39678 (N_39678,N_39310,N_39108);
nand U39679 (N_39679,N_39372,N_39322);
nand U39680 (N_39680,N_39029,N_39213);
nand U39681 (N_39681,N_39313,N_39117);
or U39682 (N_39682,N_39094,N_39369);
nand U39683 (N_39683,N_39202,N_39146);
nand U39684 (N_39684,N_39376,N_39058);
nand U39685 (N_39685,N_39433,N_39437);
and U39686 (N_39686,N_39349,N_39470);
or U39687 (N_39687,N_39399,N_39477);
nand U39688 (N_39688,N_39396,N_39167);
or U39689 (N_39689,N_39448,N_39357);
nor U39690 (N_39690,N_39291,N_39373);
or U39691 (N_39691,N_39434,N_39124);
xnor U39692 (N_39692,N_39037,N_39210);
or U39693 (N_39693,N_39171,N_39286);
and U39694 (N_39694,N_39212,N_39018);
or U39695 (N_39695,N_39272,N_39428);
nand U39696 (N_39696,N_39411,N_39339);
and U39697 (N_39697,N_39103,N_39154);
nand U39698 (N_39698,N_39280,N_39111);
or U39699 (N_39699,N_39332,N_39136);
and U39700 (N_39700,N_39450,N_39211);
nand U39701 (N_39701,N_39431,N_39162);
nor U39702 (N_39702,N_39426,N_39341);
or U39703 (N_39703,N_39405,N_39168);
nand U39704 (N_39704,N_39119,N_39129);
and U39705 (N_39705,N_39208,N_39427);
or U39706 (N_39706,N_39050,N_39456);
or U39707 (N_39707,N_39214,N_39188);
xor U39708 (N_39708,N_39460,N_39277);
or U39709 (N_39709,N_39107,N_39068);
and U39710 (N_39710,N_39425,N_39009);
xor U39711 (N_39711,N_39175,N_39346);
nand U39712 (N_39712,N_39415,N_39377);
nor U39713 (N_39713,N_39196,N_39336);
or U39714 (N_39714,N_39413,N_39071);
and U39715 (N_39715,N_39164,N_39348);
or U39716 (N_39716,N_39036,N_39342);
or U39717 (N_39717,N_39231,N_39462);
xnor U39718 (N_39718,N_39260,N_39271);
or U39719 (N_39719,N_39300,N_39252);
xor U39720 (N_39720,N_39247,N_39161);
nand U39721 (N_39721,N_39401,N_39207);
and U39722 (N_39722,N_39012,N_39218);
nor U39723 (N_39723,N_39368,N_39412);
nor U39724 (N_39724,N_39315,N_39114);
nor U39725 (N_39725,N_39021,N_39224);
and U39726 (N_39726,N_39430,N_39060);
xnor U39727 (N_39727,N_39249,N_39047);
nand U39728 (N_39728,N_39253,N_39082);
and U39729 (N_39729,N_39001,N_39156);
or U39730 (N_39730,N_39244,N_39480);
or U39731 (N_39731,N_39130,N_39219);
nor U39732 (N_39732,N_39397,N_39436);
or U39733 (N_39733,N_39178,N_39299);
nand U39734 (N_39734,N_39297,N_39106);
or U39735 (N_39735,N_39245,N_39003);
nor U39736 (N_39736,N_39484,N_39347);
nor U39737 (N_39737,N_39229,N_39498);
xnor U39738 (N_39738,N_39279,N_39032);
nand U39739 (N_39739,N_39097,N_39303);
nor U39740 (N_39740,N_39105,N_39221);
or U39741 (N_39741,N_39321,N_39283);
and U39742 (N_39742,N_39417,N_39473);
and U39743 (N_39743,N_39102,N_39270);
nor U39744 (N_39744,N_39385,N_39439);
xor U39745 (N_39745,N_39378,N_39151);
nor U39746 (N_39746,N_39306,N_39443);
nor U39747 (N_39747,N_39381,N_39116);
xor U39748 (N_39748,N_39073,N_39429);
or U39749 (N_39749,N_39485,N_39360);
xor U39750 (N_39750,N_39031,N_39025);
or U39751 (N_39751,N_39419,N_39018);
or U39752 (N_39752,N_39206,N_39411);
nand U39753 (N_39753,N_39089,N_39036);
nand U39754 (N_39754,N_39465,N_39191);
or U39755 (N_39755,N_39405,N_39129);
or U39756 (N_39756,N_39079,N_39382);
and U39757 (N_39757,N_39332,N_39172);
or U39758 (N_39758,N_39359,N_39444);
and U39759 (N_39759,N_39398,N_39273);
nand U39760 (N_39760,N_39157,N_39102);
xnor U39761 (N_39761,N_39065,N_39287);
xor U39762 (N_39762,N_39185,N_39420);
nand U39763 (N_39763,N_39465,N_39369);
xnor U39764 (N_39764,N_39199,N_39461);
and U39765 (N_39765,N_39449,N_39333);
xnor U39766 (N_39766,N_39001,N_39406);
nor U39767 (N_39767,N_39473,N_39201);
and U39768 (N_39768,N_39166,N_39485);
xor U39769 (N_39769,N_39083,N_39210);
and U39770 (N_39770,N_39394,N_39221);
nand U39771 (N_39771,N_39307,N_39426);
and U39772 (N_39772,N_39259,N_39068);
xnor U39773 (N_39773,N_39135,N_39451);
nor U39774 (N_39774,N_39269,N_39041);
or U39775 (N_39775,N_39095,N_39253);
nor U39776 (N_39776,N_39123,N_39189);
or U39777 (N_39777,N_39032,N_39439);
and U39778 (N_39778,N_39457,N_39227);
and U39779 (N_39779,N_39287,N_39356);
or U39780 (N_39780,N_39312,N_39327);
nor U39781 (N_39781,N_39198,N_39282);
xnor U39782 (N_39782,N_39031,N_39239);
or U39783 (N_39783,N_39055,N_39463);
and U39784 (N_39784,N_39254,N_39004);
and U39785 (N_39785,N_39155,N_39419);
or U39786 (N_39786,N_39407,N_39042);
nor U39787 (N_39787,N_39359,N_39304);
nand U39788 (N_39788,N_39178,N_39134);
nand U39789 (N_39789,N_39457,N_39128);
nand U39790 (N_39790,N_39062,N_39456);
nand U39791 (N_39791,N_39188,N_39221);
nor U39792 (N_39792,N_39332,N_39231);
nor U39793 (N_39793,N_39326,N_39195);
and U39794 (N_39794,N_39144,N_39050);
nand U39795 (N_39795,N_39145,N_39336);
or U39796 (N_39796,N_39421,N_39390);
nor U39797 (N_39797,N_39072,N_39316);
or U39798 (N_39798,N_39006,N_39313);
or U39799 (N_39799,N_39133,N_39484);
xor U39800 (N_39800,N_39116,N_39457);
or U39801 (N_39801,N_39285,N_39206);
and U39802 (N_39802,N_39310,N_39071);
nor U39803 (N_39803,N_39463,N_39033);
or U39804 (N_39804,N_39384,N_39156);
and U39805 (N_39805,N_39412,N_39092);
xnor U39806 (N_39806,N_39491,N_39219);
nand U39807 (N_39807,N_39067,N_39350);
nand U39808 (N_39808,N_39341,N_39488);
nor U39809 (N_39809,N_39344,N_39432);
nand U39810 (N_39810,N_39095,N_39083);
or U39811 (N_39811,N_39249,N_39383);
or U39812 (N_39812,N_39103,N_39221);
nor U39813 (N_39813,N_39266,N_39014);
or U39814 (N_39814,N_39179,N_39376);
nor U39815 (N_39815,N_39328,N_39284);
or U39816 (N_39816,N_39222,N_39402);
xnor U39817 (N_39817,N_39490,N_39288);
xor U39818 (N_39818,N_39255,N_39137);
xor U39819 (N_39819,N_39139,N_39085);
xnor U39820 (N_39820,N_39307,N_39001);
or U39821 (N_39821,N_39279,N_39459);
nand U39822 (N_39822,N_39382,N_39263);
xor U39823 (N_39823,N_39287,N_39003);
and U39824 (N_39824,N_39240,N_39372);
xor U39825 (N_39825,N_39391,N_39363);
and U39826 (N_39826,N_39066,N_39175);
or U39827 (N_39827,N_39209,N_39179);
or U39828 (N_39828,N_39148,N_39266);
nor U39829 (N_39829,N_39224,N_39049);
nor U39830 (N_39830,N_39429,N_39126);
and U39831 (N_39831,N_39197,N_39186);
nor U39832 (N_39832,N_39084,N_39473);
nor U39833 (N_39833,N_39096,N_39021);
nor U39834 (N_39834,N_39014,N_39150);
and U39835 (N_39835,N_39423,N_39142);
nand U39836 (N_39836,N_39263,N_39249);
or U39837 (N_39837,N_39004,N_39133);
and U39838 (N_39838,N_39298,N_39488);
and U39839 (N_39839,N_39340,N_39411);
nor U39840 (N_39840,N_39016,N_39417);
and U39841 (N_39841,N_39413,N_39230);
nor U39842 (N_39842,N_39406,N_39098);
and U39843 (N_39843,N_39134,N_39300);
and U39844 (N_39844,N_39396,N_39404);
and U39845 (N_39845,N_39363,N_39188);
nand U39846 (N_39846,N_39421,N_39009);
nor U39847 (N_39847,N_39146,N_39219);
nand U39848 (N_39848,N_39011,N_39404);
xnor U39849 (N_39849,N_39402,N_39312);
and U39850 (N_39850,N_39264,N_39316);
nor U39851 (N_39851,N_39005,N_39309);
nand U39852 (N_39852,N_39309,N_39265);
and U39853 (N_39853,N_39242,N_39058);
xor U39854 (N_39854,N_39241,N_39102);
or U39855 (N_39855,N_39228,N_39453);
nand U39856 (N_39856,N_39386,N_39026);
nand U39857 (N_39857,N_39296,N_39129);
and U39858 (N_39858,N_39468,N_39162);
xnor U39859 (N_39859,N_39337,N_39376);
xor U39860 (N_39860,N_39499,N_39213);
xor U39861 (N_39861,N_39493,N_39291);
xor U39862 (N_39862,N_39266,N_39400);
nor U39863 (N_39863,N_39427,N_39280);
nand U39864 (N_39864,N_39417,N_39157);
xor U39865 (N_39865,N_39242,N_39191);
nand U39866 (N_39866,N_39357,N_39148);
nor U39867 (N_39867,N_39377,N_39299);
or U39868 (N_39868,N_39353,N_39382);
and U39869 (N_39869,N_39084,N_39461);
nor U39870 (N_39870,N_39133,N_39362);
and U39871 (N_39871,N_39071,N_39131);
xor U39872 (N_39872,N_39086,N_39368);
or U39873 (N_39873,N_39283,N_39223);
nor U39874 (N_39874,N_39188,N_39169);
xnor U39875 (N_39875,N_39189,N_39306);
and U39876 (N_39876,N_39490,N_39183);
xor U39877 (N_39877,N_39415,N_39359);
xor U39878 (N_39878,N_39485,N_39105);
or U39879 (N_39879,N_39300,N_39113);
or U39880 (N_39880,N_39432,N_39308);
xor U39881 (N_39881,N_39342,N_39022);
or U39882 (N_39882,N_39205,N_39493);
and U39883 (N_39883,N_39240,N_39475);
and U39884 (N_39884,N_39083,N_39006);
or U39885 (N_39885,N_39270,N_39236);
nand U39886 (N_39886,N_39294,N_39365);
and U39887 (N_39887,N_39493,N_39373);
nor U39888 (N_39888,N_39102,N_39275);
or U39889 (N_39889,N_39383,N_39128);
and U39890 (N_39890,N_39323,N_39226);
nand U39891 (N_39891,N_39180,N_39043);
nor U39892 (N_39892,N_39340,N_39488);
nor U39893 (N_39893,N_39146,N_39234);
xnor U39894 (N_39894,N_39134,N_39319);
xnor U39895 (N_39895,N_39440,N_39365);
nand U39896 (N_39896,N_39442,N_39349);
nor U39897 (N_39897,N_39201,N_39354);
xor U39898 (N_39898,N_39043,N_39383);
nand U39899 (N_39899,N_39197,N_39126);
and U39900 (N_39900,N_39236,N_39254);
nand U39901 (N_39901,N_39238,N_39031);
or U39902 (N_39902,N_39047,N_39453);
nand U39903 (N_39903,N_39442,N_39401);
xor U39904 (N_39904,N_39059,N_39223);
or U39905 (N_39905,N_39194,N_39470);
xor U39906 (N_39906,N_39194,N_39466);
and U39907 (N_39907,N_39299,N_39103);
nor U39908 (N_39908,N_39086,N_39280);
and U39909 (N_39909,N_39405,N_39225);
and U39910 (N_39910,N_39100,N_39394);
nor U39911 (N_39911,N_39312,N_39403);
nand U39912 (N_39912,N_39190,N_39066);
nand U39913 (N_39913,N_39411,N_39101);
nor U39914 (N_39914,N_39320,N_39121);
nand U39915 (N_39915,N_39180,N_39476);
or U39916 (N_39916,N_39298,N_39439);
nor U39917 (N_39917,N_39395,N_39314);
and U39918 (N_39918,N_39117,N_39255);
and U39919 (N_39919,N_39178,N_39166);
and U39920 (N_39920,N_39248,N_39126);
nor U39921 (N_39921,N_39424,N_39024);
xnor U39922 (N_39922,N_39075,N_39386);
nor U39923 (N_39923,N_39161,N_39206);
nand U39924 (N_39924,N_39149,N_39338);
nor U39925 (N_39925,N_39413,N_39214);
and U39926 (N_39926,N_39221,N_39151);
or U39927 (N_39927,N_39135,N_39018);
nand U39928 (N_39928,N_39491,N_39053);
nor U39929 (N_39929,N_39377,N_39140);
nor U39930 (N_39930,N_39186,N_39114);
nand U39931 (N_39931,N_39441,N_39445);
and U39932 (N_39932,N_39285,N_39015);
nor U39933 (N_39933,N_39290,N_39404);
nand U39934 (N_39934,N_39224,N_39354);
or U39935 (N_39935,N_39324,N_39023);
or U39936 (N_39936,N_39076,N_39119);
nor U39937 (N_39937,N_39252,N_39136);
xor U39938 (N_39938,N_39381,N_39327);
nand U39939 (N_39939,N_39180,N_39443);
xnor U39940 (N_39940,N_39348,N_39134);
and U39941 (N_39941,N_39347,N_39330);
nand U39942 (N_39942,N_39490,N_39458);
xnor U39943 (N_39943,N_39381,N_39129);
nand U39944 (N_39944,N_39483,N_39401);
nand U39945 (N_39945,N_39014,N_39130);
and U39946 (N_39946,N_39352,N_39459);
xor U39947 (N_39947,N_39275,N_39286);
or U39948 (N_39948,N_39036,N_39451);
or U39949 (N_39949,N_39356,N_39024);
nor U39950 (N_39950,N_39069,N_39193);
and U39951 (N_39951,N_39094,N_39020);
or U39952 (N_39952,N_39336,N_39338);
xor U39953 (N_39953,N_39240,N_39261);
nor U39954 (N_39954,N_39258,N_39168);
nor U39955 (N_39955,N_39422,N_39486);
or U39956 (N_39956,N_39265,N_39466);
nor U39957 (N_39957,N_39432,N_39286);
xor U39958 (N_39958,N_39011,N_39038);
nor U39959 (N_39959,N_39050,N_39066);
nor U39960 (N_39960,N_39010,N_39442);
or U39961 (N_39961,N_39440,N_39371);
or U39962 (N_39962,N_39389,N_39016);
nand U39963 (N_39963,N_39479,N_39194);
and U39964 (N_39964,N_39132,N_39337);
xnor U39965 (N_39965,N_39111,N_39394);
or U39966 (N_39966,N_39092,N_39051);
and U39967 (N_39967,N_39186,N_39091);
or U39968 (N_39968,N_39358,N_39100);
xnor U39969 (N_39969,N_39415,N_39181);
and U39970 (N_39970,N_39422,N_39103);
and U39971 (N_39971,N_39496,N_39436);
nand U39972 (N_39972,N_39269,N_39044);
nand U39973 (N_39973,N_39224,N_39475);
or U39974 (N_39974,N_39048,N_39239);
nor U39975 (N_39975,N_39101,N_39487);
nand U39976 (N_39976,N_39423,N_39367);
nand U39977 (N_39977,N_39332,N_39498);
xnor U39978 (N_39978,N_39358,N_39476);
nand U39979 (N_39979,N_39439,N_39003);
and U39980 (N_39980,N_39089,N_39448);
nand U39981 (N_39981,N_39110,N_39341);
xor U39982 (N_39982,N_39457,N_39234);
xor U39983 (N_39983,N_39375,N_39109);
xnor U39984 (N_39984,N_39375,N_39324);
nand U39985 (N_39985,N_39398,N_39428);
xnor U39986 (N_39986,N_39456,N_39144);
or U39987 (N_39987,N_39253,N_39370);
or U39988 (N_39988,N_39382,N_39342);
or U39989 (N_39989,N_39464,N_39187);
or U39990 (N_39990,N_39367,N_39183);
nand U39991 (N_39991,N_39004,N_39289);
nand U39992 (N_39992,N_39008,N_39153);
and U39993 (N_39993,N_39238,N_39107);
or U39994 (N_39994,N_39358,N_39481);
and U39995 (N_39995,N_39131,N_39074);
and U39996 (N_39996,N_39418,N_39043);
nor U39997 (N_39997,N_39111,N_39178);
xor U39998 (N_39998,N_39286,N_39246);
nor U39999 (N_39999,N_39184,N_39443);
nand U40000 (N_40000,N_39899,N_39559);
nand U40001 (N_40001,N_39594,N_39706);
xnor U40002 (N_40002,N_39863,N_39518);
nor U40003 (N_40003,N_39709,N_39891);
xnor U40004 (N_40004,N_39539,N_39750);
nand U40005 (N_40005,N_39575,N_39897);
nor U40006 (N_40006,N_39942,N_39693);
nand U40007 (N_40007,N_39603,N_39620);
nand U40008 (N_40008,N_39619,N_39935);
or U40009 (N_40009,N_39585,N_39826);
xor U40010 (N_40010,N_39756,N_39547);
and U40011 (N_40011,N_39574,N_39682);
nor U40012 (N_40012,N_39877,N_39802);
and U40013 (N_40013,N_39552,N_39917);
or U40014 (N_40014,N_39950,N_39663);
nand U40015 (N_40015,N_39849,N_39900);
xnor U40016 (N_40016,N_39673,N_39595);
nand U40017 (N_40017,N_39541,N_39854);
xor U40018 (N_40018,N_39681,N_39737);
and U40019 (N_40019,N_39570,N_39761);
and U40020 (N_40020,N_39872,N_39949);
and U40021 (N_40021,N_39748,N_39726);
xnor U40022 (N_40022,N_39718,N_39712);
nand U40023 (N_40023,N_39556,N_39501);
and U40024 (N_40024,N_39542,N_39876);
and U40025 (N_40025,N_39962,N_39698);
nand U40026 (N_40026,N_39655,N_39778);
nor U40027 (N_40027,N_39623,N_39880);
and U40028 (N_40028,N_39704,N_39845);
and U40029 (N_40029,N_39782,N_39636);
nand U40030 (N_40030,N_39557,N_39631);
and U40031 (N_40031,N_39892,N_39569);
nand U40032 (N_40032,N_39861,N_39525);
and U40033 (N_40033,N_39963,N_39801);
or U40034 (N_40034,N_39973,N_39974);
xnor U40035 (N_40035,N_39776,N_39651);
nand U40036 (N_40036,N_39784,N_39551);
nand U40037 (N_40037,N_39817,N_39831);
nor U40038 (N_40038,N_39987,N_39903);
nor U40039 (N_40039,N_39568,N_39610);
and U40040 (N_40040,N_39509,N_39689);
nand U40041 (N_40041,N_39504,N_39656);
nor U40042 (N_40042,N_39716,N_39928);
or U40043 (N_40043,N_39933,N_39508);
and U40044 (N_40044,N_39964,N_39835);
or U40045 (N_40045,N_39922,N_39611);
nand U40046 (N_40046,N_39824,N_39680);
nand U40047 (N_40047,N_39617,N_39540);
or U40048 (N_40048,N_39510,N_39792);
or U40049 (N_40049,N_39740,N_39760);
xnor U40050 (N_40050,N_39905,N_39844);
nand U40051 (N_40051,N_39885,N_39652);
and U40052 (N_40052,N_39781,N_39536);
xor U40053 (N_40053,N_39645,N_39630);
or U40054 (N_40054,N_39972,N_39660);
xor U40055 (N_40055,N_39520,N_39654);
xnor U40056 (N_40056,N_39507,N_39516);
nand U40057 (N_40057,N_39637,N_39976);
and U40058 (N_40058,N_39548,N_39772);
nand U40059 (N_40059,N_39530,N_39662);
nand U40060 (N_40060,N_39531,N_39930);
or U40061 (N_40061,N_39668,N_39956);
or U40062 (N_40062,N_39633,N_39780);
and U40063 (N_40063,N_39647,N_39785);
or U40064 (N_40064,N_39995,N_39939);
xor U40065 (N_40065,N_39884,N_39565);
and U40066 (N_40066,N_39538,N_39841);
or U40067 (N_40067,N_39572,N_39730);
nand U40068 (N_40068,N_39522,N_39747);
nand U40069 (N_40069,N_39519,N_39819);
xnor U40070 (N_40070,N_39832,N_39901);
or U40071 (N_40071,N_39998,N_39794);
and U40072 (N_40072,N_39825,N_39895);
nor U40073 (N_40073,N_39996,N_39758);
nor U40074 (N_40074,N_39582,N_39929);
nor U40075 (N_40075,N_39641,N_39699);
and U40076 (N_40076,N_39855,N_39627);
nand U40077 (N_40077,N_39634,N_39511);
nand U40078 (N_40078,N_39560,N_39715);
and U40079 (N_40079,N_39852,N_39601);
xor U40080 (N_40080,N_39881,N_39791);
and U40081 (N_40081,N_39561,N_39853);
and U40082 (N_40082,N_39944,N_39691);
and U40083 (N_40083,N_39717,N_39809);
or U40084 (N_40084,N_39606,N_39960);
xnor U40085 (N_40085,N_39829,N_39678);
nand U40086 (N_40086,N_39579,N_39923);
and U40087 (N_40087,N_39787,N_39789);
and U40088 (N_40088,N_39577,N_39598);
and U40089 (N_40089,N_39613,N_39586);
nor U40090 (N_40090,N_39688,N_39524);
and U40091 (N_40091,N_39834,N_39867);
and U40092 (N_40092,N_39755,N_39578);
or U40093 (N_40093,N_39564,N_39978);
and U40094 (N_40094,N_39943,N_39759);
nor U40095 (N_40095,N_39725,N_39988);
nor U40096 (N_40096,N_39544,N_39743);
or U40097 (N_40097,N_39692,N_39571);
and U40098 (N_40098,N_39909,N_39773);
xor U40099 (N_40099,N_39865,N_39906);
xnor U40100 (N_40100,N_39584,N_39590);
and U40101 (N_40101,N_39675,N_39968);
and U40102 (N_40102,N_39665,N_39573);
or U40103 (N_40103,N_39959,N_39528);
nand U40104 (N_40104,N_39851,N_39650);
or U40105 (N_40105,N_39607,N_39806);
or U40106 (N_40106,N_39874,N_39830);
or U40107 (N_40107,N_39934,N_39947);
nand U40108 (N_40108,N_39907,N_39741);
and U40109 (N_40109,N_39599,N_39646);
and U40110 (N_40110,N_39587,N_39866);
nand U40111 (N_40111,N_39875,N_39946);
nor U40112 (N_40112,N_39757,N_39970);
nand U40113 (N_40113,N_39957,N_39596);
nand U40114 (N_40114,N_39546,N_39527);
xnor U40115 (N_40115,N_39639,N_39969);
nor U40116 (N_40116,N_39925,N_39612);
xnor U40117 (N_40117,N_39958,N_39793);
xnor U40118 (N_40118,N_39979,N_39549);
and U40119 (N_40119,N_39764,N_39864);
xnor U40120 (N_40120,N_39770,N_39615);
xnor U40121 (N_40121,N_39768,N_39847);
and U40122 (N_40122,N_39670,N_39896);
xnor U40123 (N_40123,N_39767,N_39990);
and U40124 (N_40124,N_39703,N_39625);
nand U40125 (N_40125,N_39882,N_39889);
xor U40126 (N_40126,N_39608,N_39769);
or U40127 (N_40127,N_39989,N_39635);
nor U40128 (N_40128,N_39697,N_39797);
nand U40129 (N_40129,N_39734,N_39505);
or U40130 (N_40130,N_39961,N_39775);
xnor U40131 (N_40131,N_39529,N_39604);
and U40132 (N_40132,N_39813,N_39883);
xor U40133 (N_40133,N_39658,N_39719);
nor U40134 (N_40134,N_39711,N_39555);
nor U40135 (N_40135,N_39992,N_39839);
or U40136 (N_40136,N_39890,N_39811);
nor U40137 (N_40137,N_39954,N_39659);
xnor U40138 (N_40138,N_39567,N_39533);
or U40139 (N_40139,N_39975,N_39723);
nor U40140 (N_40140,N_39563,N_39669);
nor U40141 (N_40141,N_39931,N_39967);
xnor U40142 (N_40142,N_39948,N_39763);
xnor U40143 (N_40143,N_39671,N_39628);
or U40144 (N_40144,N_39937,N_39593);
nor U40145 (N_40145,N_39986,N_39643);
nor U40146 (N_40146,N_39815,N_39583);
nand U40147 (N_40147,N_39600,N_39677);
xnor U40148 (N_40148,N_39710,N_39821);
or U40149 (N_40149,N_39733,N_39997);
and U40150 (N_40150,N_39629,N_39796);
and U40151 (N_40151,N_39915,N_39614);
or U40152 (N_40152,N_39887,N_39859);
or U40153 (N_40153,N_39696,N_39843);
xor U40154 (N_40154,N_39744,N_39800);
and U40155 (N_40155,N_39640,N_39838);
xnor U40156 (N_40156,N_39690,N_39816);
nor U40157 (N_40157,N_39952,N_39945);
nand U40158 (N_40158,N_39532,N_39827);
xor U40159 (N_40159,N_39918,N_39914);
nand U40160 (N_40160,N_39856,N_39846);
and U40161 (N_40161,N_39705,N_39912);
and U40162 (N_40162,N_39514,N_39731);
or U40163 (N_40163,N_39862,N_39878);
or U40164 (N_40164,N_39842,N_39919);
xnor U40165 (N_40165,N_39624,N_39999);
or U40166 (N_40166,N_39666,N_39777);
nor U40167 (N_40167,N_39921,N_39732);
xor U40168 (N_40168,N_39728,N_39940);
and U40169 (N_40169,N_39537,N_39562);
nor U40170 (N_40170,N_39951,N_39700);
nand U40171 (N_40171,N_39902,N_39953);
xor U40172 (N_40172,N_39664,N_39984);
or U40173 (N_40173,N_39724,N_39526);
nor U40174 (N_40174,N_39870,N_39779);
nor U40175 (N_40175,N_39685,N_39893);
and U40176 (N_40176,N_39814,N_39736);
nor U40177 (N_40177,N_39983,N_39661);
nor U40178 (N_40178,N_39833,N_39910);
nor U40179 (N_40179,N_39674,N_39828);
or U40180 (N_40180,N_39840,N_39879);
and U40181 (N_40181,N_39808,N_39722);
xnor U40182 (N_40182,N_39762,N_39807);
xor U40183 (N_40183,N_39672,N_39980);
xnor U40184 (N_40184,N_39591,N_39994);
and U40185 (N_40185,N_39812,N_39676);
and U40186 (N_40186,N_39523,N_39913);
nor U40187 (N_40187,N_39965,N_39786);
and U40188 (N_40188,N_39517,N_39746);
nand U40189 (N_40189,N_39868,N_39871);
xor U40190 (N_40190,N_39727,N_39721);
nand U40191 (N_40191,N_39754,N_39920);
and U40192 (N_40192,N_39869,N_39550);
and U40193 (N_40193,N_39774,N_39941);
nand U40194 (N_40194,N_39687,N_39589);
and U40195 (N_40195,N_39771,N_39745);
and U40196 (N_40196,N_39581,N_39667);
nor U40197 (N_40197,N_39632,N_39795);
nor U40198 (N_40198,N_39805,N_39616);
or U40199 (N_40199,N_39597,N_39848);
and U40200 (N_40200,N_39626,N_39790);
xor U40201 (N_40201,N_39648,N_39837);
nand U40202 (N_40202,N_39908,N_39503);
nand U40203 (N_40203,N_39911,N_39738);
xnor U40204 (N_40204,N_39588,N_39515);
nor U40205 (N_40205,N_39729,N_39753);
nor U40206 (N_40206,N_39823,N_39810);
and U40207 (N_40207,N_39576,N_39642);
xnor U40208 (N_40208,N_39720,N_39554);
or U40209 (N_40209,N_39506,N_39708);
nand U40210 (N_40210,N_39512,N_39924);
nand U40211 (N_40211,N_39873,N_39713);
or U40212 (N_40212,N_39558,N_39886);
nand U40213 (N_40213,N_39981,N_39955);
nand U40214 (N_40214,N_39938,N_39534);
and U40215 (N_40215,N_39799,N_39857);
nand U40216 (N_40216,N_39888,N_39580);
nor U40217 (N_40217,N_39766,N_39638);
nand U40218 (N_40218,N_39535,N_39971);
nor U40219 (N_40219,N_39836,N_39977);
nand U40220 (N_40220,N_39818,N_39735);
and U40221 (N_40221,N_39860,N_39798);
and U40222 (N_40222,N_39543,N_39500);
or U40223 (N_40223,N_39742,N_39752);
xnor U40224 (N_40224,N_39751,N_39592);
nor U40225 (N_40225,N_39695,N_39649);
and U40226 (N_40226,N_39618,N_39602);
and U40227 (N_40227,N_39985,N_39904);
nand U40228 (N_40228,N_39694,N_39714);
and U40229 (N_40229,N_39783,N_39609);
or U40230 (N_40230,N_39858,N_39804);
nand U40231 (N_40231,N_39803,N_39657);
and U40232 (N_40232,N_39644,N_39916);
xnor U40233 (N_40233,N_39993,N_39684);
or U40234 (N_40234,N_39686,N_39621);
nor U40235 (N_40235,N_39822,N_39513);
and U40236 (N_40236,N_39702,N_39932);
xor U40237 (N_40237,N_39788,N_39545);
nor U40238 (N_40238,N_39765,N_39966);
or U40239 (N_40239,N_39926,N_39927);
nor U40240 (N_40240,N_39749,N_39502);
nand U40241 (N_40241,N_39605,N_39898);
xor U40242 (N_40242,N_39679,N_39936);
nor U40243 (N_40243,N_39739,N_39701);
nand U40244 (N_40244,N_39894,N_39991);
nor U40245 (N_40245,N_39683,N_39566);
and U40246 (N_40246,N_39820,N_39982);
nor U40247 (N_40247,N_39521,N_39850);
nor U40248 (N_40248,N_39553,N_39707);
nor U40249 (N_40249,N_39622,N_39653);
xor U40250 (N_40250,N_39943,N_39836);
xor U40251 (N_40251,N_39793,N_39715);
nor U40252 (N_40252,N_39536,N_39939);
nand U40253 (N_40253,N_39684,N_39518);
nand U40254 (N_40254,N_39822,N_39557);
nor U40255 (N_40255,N_39687,N_39559);
nor U40256 (N_40256,N_39570,N_39683);
and U40257 (N_40257,N_39608,N_39759);
and U40258 (N_40258,N_39978,N_39598);
and U40259 (N_40259,N_39939,N_39624);
nand U40260 (N_40260,N_39807,N_39687);
or U40261 (N_40261,N_39960,N_39686);
nor U40262 (N_40262,N_39995,N_39845);
and U40263 (N_40263,N_39629,N_39766);
nand U40264 (N_40264,N_39595,N_39706);
or U40265 (N_40265,N_39945,N_39532);
or U40266 (N_40266,N_39770,N_39838);
xor U40267 (N_40267,N_39564,N_39625);
xnor U40268 (N_40268,N_39502,N_39500);
or U40269 (N_40269,N_39693,N_39612);
or U40270 (N_40270,N_39976,N_39842);
nor U40271 (N_40271,N_39518,N_39833);
or U40272 (N_40272,N_39960,N_39539);
nand U40273 (N_40273,N_39928,N_39706);
nand U40274 (N_40274,N_39561,N_39573);
nor U40275 (N_40275,N_39810,N_39716);
or U40276 (N_40276,N_39510,N_39638);
nor U40277 (N_40277,N_39888,N_39958);
and U40278 (N_40278,N_39505,N_39915);
xnor U40279 (N_40279,N_39663,N_39995);
nor U40280 (N_40280,N_39935,N_39956);
nor U40281 (N_40281,N_39845,N_39705);
and U40282 (N_40282,N_39671,N_39557);
nand U40283 (N_40283,N_39982,N_39901);
nand U40284 (N_40284,N_39657,N_39729);
or U40285 (N_40285,N_39934,N_39538);
nand U40286 (N_40286,N_39633,N_39704);
or U40287 (N_40287,N_39793,N_39870);
nor U40288 (N_40288,N_39843,N_39793);
or U40289 (N_40289,N_39828,N_39866);
nor U40290 (N_40290,N_39898,N_39648);
or U40291 (N_40291,N_39987,N_39862);
nand U40292 (N_40292,N_39546,N_39979);
and U40293 (N_40293,N_39933,N_39795);
xnor U40294 (N_40294,N_39929,N_39647);
xnor U40295 (N_40295,N_39927,N_39512);
nor U40296 (N_40296,N_39807,N_39640);
and U40297 (N_40297,N_39918,N_39906);
xor U40298 (N_40298,N_39695,N_39948);
nor U40299 (N_40299,N_39624,N_39918);
nand U40300 (N_40300,N_39644,N_39565);
nor U40301 (N_40301,N_39525,N_39673);
or U40302 (N_40302,N_39829,N_39763);
nand U40303 (N_40303,N_39708,N_39810);
or U40304 (N_40304,N_39817,N_39551);
or U40305 (N_40305,N_39672,N_39609);
xnor U40306 (N_40306,N_39931,N_39933);
nand U40307 (N_40307,N_39951,N_39618);
xor U40308 (N_40308,N_39645,N_39682);
nor U40309 (N_40309,N_39954,N_39861);
nand U40310 (N_40310,N_39998,N_39903);
and U40311 (N_40311,N_39947,N_39959);
nor U40312 (N_40312,N_39975,N_39646);
xor U40313 (N_40313,N_39731,N_39748);
and U40314 (N_40314,N_39914,N_39676);
nand U40315 (N_40315,N_39536,N_39575);
xor U40316 (N_40316,N_39873,N_39952);
xnor U40317 (N_40317,N_39818,N_39514);
or U40318 (N_40318,N_39685,N_39568);
and U40319 (N_40319,N_39524,N_39666);
or U40320 (N_40320,N_39950,N_39557);
nand U40321 (N_40321,N_39739,N_39616);
and U40322 (N_40322,N_39995,N_39636);
nand U40323 (N_40323,N_39798,N_39695);
xor U40324 (N_40324,N_39998,N_39881);
nor U40325 (N_40325,N_39559,N_39996);
and U40326 (N_40326,N_39931,N_39786);
xnor U40327 (N_40327,N_39931,N_39560);
and U40328 (N_40328,N_39555,N_39861);
or U40329 (N_40329,N_39896,N_39917);
and U40330 (N_40330,N_39630,N_39959);
or U40331 (N_40331,N_39811,N_39574);
and U40332 (N_40332,N_39537,N_39999);
nand U40333 (N_40333,N_39679,N_39603);
and U40334 (N_40334,N_39705,N_39852);
nand U40335 (N_40335,N_39888,N_39893);
nor U40336 (N_40336,N_39776,N_39920);
and U40337 (N_40337,N_39807,N_39981);
nor U40338 (N_40338,N_39783,N_39874);
nor U40339 (N_40339,N_39724,N_39575);
nor U40340 (N_40340,N_39942,N_39806);
or U40341 (N_40341,N_39947,N_39515);
nor U40342 (N_40342,N_39974,N_39635);
or U40343 (N_40343,N_39775,N_39654);
nor U40344 (N_40344,N_39857,N_39587);
nor U40345 (N_40345,N_39726,N_39510);
and U40346 (N_40346,N_39928,N_39661);
or U40347 (N_40347,N_39842,N_39546);
nor U40348 (N_40348,N_39602,N_39859);
nand U40349 (N_40349,N_39626,N_39750);
and U40350 (N_40350,N_39856,N_39526);
nor U40351 (N_40351,N_39802,N_39522);
xor U40352 (N_40352,N_39621,N_39995);
or U40353 (N_40353,N_39742,N_39882);
nor U40354 (N_40354,N_39607,N_39515);
xor U40355 (N_40355,N_39881,N_39969);
nand U40356 (N_40356,N_39775,N_39616);
nor U40357 (N_40357,N_39696,N_39704);
and U40358 (N_40358,N_39817,N_39786);
nor U40359 (N_40359,N_39574,N_39591);
xor U40360 (N_40360,N_39903,N_39678);
or U40361 (N_40361,N_39625,N_39753);
or U40362 (N_40362,N_39794,N_39706);
or U40363 (N_40363,N_39500,N_39538);
or U40364 (N_40364,N_39599,N_39839);
nand U40365 (N_40365,N_39936,N_39515);
nand U40366 (N_40366,N_39579,N_39680);
or U40367 (N_40367,N_39562,N_39879);
nor U40368 (N_40368,N_39592,N_39908);
or U40369 (N_40369,N_39595,N_39511);
nor U40370 (N_40370,N_39844,N_39504);
and U40371 (N_40371,N_39928,N_39859);
and U40372 (N_40372,N_39607,N_39683);
and U40373 (N_40373,N_39500,N_39546);
xor U40374 (N_40374,N_39572,N_39737);
or U40375 (N_40375,N_39570,N_39529);
nor U40376 (N_40376,N_39611,N_39847);
nand U40377 (N_40377,N_39914,N_39660);
nand U40378 (N_40378,N_39694,N_39884);
and U40379 (N_40379,N_39660,N_39834);
or U40380 (N_40380,N_39595,N_39876);
nor U40381 (N_40381,N_39968,N_39500);
and U40382 (N_40382,N_39732,N_39692);
xor U40383 (N_40383,N_39503,N_39631);
and U40384 (N_40384,N_39917,N_39689);
xor U40385 (N_40385,N_39728,N_39864);
and U40386 (N_40386,N_39697,N_39886);
or U40387 (N_40387,N_39982,N_39864);
nand U40388 (N_40388,N_39993,N_39882);
or U40389 (N_40389,N_39860,N_39785);
xor U40390 (N_40390,N_39691,N_39592);
and U40391 (N_40391,N_39518,N_39819);
nor U40392 (N_40392,N_39943,N_39855);
nor U40393 (N_40393,N_39506,N_39875);
nand U40394 (N_40394,N_39800,N_39552);
nand U40395 (N_40395,N_39994,N_39995);
nor U40396 (N_40396,N_39831,N_39722);
nor U40397 (N_40397,N_39675,N_39783);
or U40398 (N_40398,N_39580,N_39763);
nand U40399 (N_40399,N_39586,N_39533);
nor U40400 (N_40400,N_39814,N_39891);
nor U40401 (N_40401,N_39678,N_39613);
and U40402 (N_40402,N_39796,N_39751);
and U40403 (N_40403,N_39513,N_39974);
nand U40404 (N_40404,N_39585,N_39763);
nand U40405 (N_40405,N_39511,N_39579);
or U40406 (N_40406,N_39615,N_39905);
nor U40407 (N_40407,N_39639,N_39773);
xnor U40408 (N_40408,N_39761,N_39565);
or U40409 (N_40409,N_39643,N_39960);
nand U40410 (N_40410,N_39996,N_39522);
or U40411 (N_40411,N_39708,N_39974);
and U40412 (N_40412,N_39770,N_39780);
nand U40413 (N_40413,N_39836,N_39548);
nand U40414 (N_40414,N_39686,N_39797);
or U40415 (N_40415,N_39823,N_39875);
and U40416 (N_40416,N_39636,N_39933);
nand U40417 (N_40417,N_39559,N_39732);
nor U40418 (N_40418,N_39984,N_39744);
nor U40419 (N_40419,N_39582,N_39788);
xor U40420 (N_40420,N_39634,N_39920);
and U40421 (N_40421,N_39911,N_39731);
xor U40422 (N_40422,N_39998,N_39702);
or U40423 (N_40423,N_39567,N_39677);
or U40424 (N_40424,N_39758,N_39670);
or U40425 (N_40425,N_39737,N_39999);
nand U40426 (N_40426,N_39685,N_39556);
or U40427 (N_40427,N_39618,N_39645);
and U40428 (N_40428,N_39903,N_39944);
or U40429 (N_40429,N_39519,N_39841);
nand U40430 (N_40430,N_39739,N_39835);
nor U40431 (N_40431,N_39750,N_39709);
or U40432 (N_40432,N_39755,N_39699);
nand U40433 (N_40433,N_39863,N_39614);
or U40434 (N_40434,N_39937,N_39707);
or U40435 (N_40435,N_39571,N_39586);
nor U40436 (N_40436,N_39732,N_39820);
nand U40437 (N_40437,N_39533,N_39768);
or U40438 (N_40438,N_39521,N_39556);
or U40439 (N_40439,N_39980,N_39855);
xnor U40440 (N_40440,N_39734,N_39763);
and U40441 (N_40441,N_39738,N_39736);
xnor U40442 (N_40442,N_39938,N_39874);
xor U40443 (N_40443,N_39953,N_39728);
xor U40444 (N_40444,N_39804,N_39857);
nand U40445 (N_40445,N_39703,N_39611);
nor U40446 (N_40446,N_39968,N_39962);
or U40447 (N_40447,N_39705,N_39782);
xor U40448 (N_40448,N_39876,N_39582);
xor U40449 (N_40449,N_39644,N_39796);
nor U40450 (N_40450,N_39780,N_39582);
xnor U40451 (N_40451,N_39563,N_39986);
nor U40452 (N_40452,N_39766,N_39798);
nor U40453 (N_40453,N_39585,N_39807);
nor U40454 (N_40454,N_39945,N_39660);
xor U40455 (N_40455,N_39769,N_39650);
and U40456 (N_40456,N_39500,N_39541);
nand U40457 (N_40457,N_39587,N_39578);
xnor U40458 (N_40458,N_39668,N_39617);
and U40459 (N_40459,N_39846,N_39715);
nand U40460 (N_40460,N_39656,N_39843);
and U40461 (N_40461,N_39646,N_39936);
xor U40462 (N_40462,N_39966,N_39950);
xnor U40463 (N_40463,N_39811,N_39992);
or U40464 (N_40464,N_39956,N_39548);
nor U40465 (N_40465,N_39582,N_39743);
or U40466 (N_40466,N_39826,N_39770);
or U40467 (N_40467,N_39869,N_39811);
nand U40468 (N_40468,N_39706,N_39901);
nor U40469 (N_40469,N_39515,N_39942);
and U40470 (N_40470,N_39508,N_39924);
nor U40471 (N_40471,N_39533,N_39605);
nand U40472 (N_40472,N_39771,N_39920);
nand U40473 (N_40473,N_39522,N_39902);
nor U40474 (N_40474,N_39985,N_39656);
nor U40475 (N_40475,N_39990,N_39950);
and U40476 (N_40476,N_39718,N_39779);
nand U40477 (N_40477,N_39545,N_39985);
nor U40478 (N_40478,N_39515,N_39586);
nor U40479 (N_40479,N_39596,N_39763);
nand U40480 (N_40480,N_39840,N_39586);
nand U40481 (N_40481,N_39680,N_39926);
nor U40482 (N_40482,N_39617,N_39829);
nand U40483 (N_40483,N_39815,N_39630);
and U40484 (N_40484,N_39869,N_39507);
xor U40485 (N_40485,N_39565,N_39971);
nand U40486 (N_40486,N_39527,N_39967);
nor U40487 (N_40487,N_39964,N_39518);
and U40488 (N_40488,N_39769,N_39850);
nand U40489 (N_40489,N_39505,N_39701);
or U40490 (N_40490,N_39861,N_39687);
or U40491 (N_40491,N_39874,N_39962);
xor U40492 (N_40492,N_39820,N_39933);
or U40493 (N_40493,N_39882,N_39603);
xor U40494 (N_40494,N_39595,N_39526);
or U40495 (N_40495,N_39859,N_39691);
xnor U40496 (N_40496,N_39988,N_39799);
xor U40497 (N_40497,N_39682,N_39909);
or U40498 (N_40498,N_39511,N_39856);
or U40499 (N_40499,N_39625,N_39771);
nor U40500 (N_40500,N_40360,N_40174);
or U40501 (N_40501,N_40445,N_40259);
and U40502 (N_40502,N_40364,N_40087);
and U40503 (N_40503,N_40398,N_40363);
nand U40504 (N_40504,N_40415,N_40099);
nand U40505 (N_40505,N_40182,N_40462);
nor U40506 (N_40506,N_40103,N_40160);
nand U40507 (N_40507,N_40092,N_40104);
and U40508 (N_40508,N_40412,N_40070);
and U40509 (N_40509,N_40424,N_40169);
nor U40510 (N_40510,N_40051,N_40325);
xnor U40511 (N_40511,N_40209,N_40002);
and U40512 (N_40512,N_40402,N_40061);
and U40513 (N_40513,N_40111,N_40423);
or U40514 (N_40514,N_40150,N_40467);
xnor U40515 (N_40515,N_40416,N_40188);
xor U40516 (N_40516,N_40373,N_40189);
or U40517 (N_40517,N_40277,N_40281);
nand U40518 (N_40518,N_40028,N_40449);
or U40519 (N_40519,N_40147,N_40330);
and U40520 (N_40520,N_40441,N_40022);
or U40521 (N_40521,N_40434,N_40359);
nor U40522 (N_40522,N_40027,N_40332);
nand U40523 (N_40523,N_40274,N_40153);
or U40524 (N_40524,N_40172,N_40013);
nor U40525 (N_40525,N_40256,N_40219);
nand U40526 (N_40526,N_40304,N_40431);
and U40527 (N_40527,N_40008,N_40474);
or U40528 (N_40528,N_40064,N_40119);
nor U40529 (N_40529,N_40260,N_40270);
nor U40530 (N_40530,N_40263,N_40163);
nand U40531 (N_40531,N_40378,N_40034);
nor U40532 (N_40532,N_40248,N_40131);
nand U40533 (N_40533,N_40037,N_40232);
xor U40534 (N_40534,N_40030,N_40183);
or U40535 (N_40535,N_40063,N_40149);
nand U40536 (N_40536,N_40354,N_40464);
nand U40537 (N_40537,N_40193,N_40102);
xor U40538 (N_40538,N_40021,N_40168);
xor U40539 (N_40539,N_40380,N_40144);
xnor U40540 (N_40540,N_40078,N_40164);
nor U40541 (N_40541,N_40116,N_40083);
nand U40542 (N_40542,N_40125,N_40101);
xor U40543 (N_40543,N_40447,N_40315);
xnor U40544 (N_40544,N_40276,N_40442);
or U40545 (N_40545,N_40026,N_40094);
nor U40546 (N_40546,N_40048,N_40459);
nand U40547 (N_40547,N_40298,N_40386);
and U40548 (N_40548,N_40140,N_40014);
or U40549 (N_40549,N_40450,N_40176);
and U40550 (N_40550,N_40479,N_40288);
and U40551 (N_40551,N_40370,N_40420);
or U40552 (N_40552,N_40042,N_40074);
nor U40553 (N_40553,N_40397,N_40293);
and U40554 (N_40554,N_40327,N_40371);
and U40555 (N_40555,N_40186,N_40292);
or U40556 (N_40556,N_40156,N_40179);
nand U40557 (N_40557,N_40046,N_40312);
or U40558 (N_40558,N_40165,N_40301);
nor U40559 (N_40559,N_40054,N_40426);
xnor U40560 (N_40560,N_40446,N_40495);
and U40561 (N_40561,N_40075,N_40494);
xor U40562 (N_40562,N_40199,N_40117);
and U40563 (N_40563,N_40480,N_40482);
xor U40564 (N_40564,N_40382,N_40353);
and U40565 (N_40565,N_40376,N_40085);
xor U40566 (N_40566,N_40234,N_40207);
or U40567 (N_40567,N_40129,N_40035);
or U40568 (N_40568,N_40145,N_40394);
nor U40569 (N_40569,N_40436,N_40461);
or U40570 (N_40570,N_40230,N_40218);
nor U40571 (N_40571,N_40250,N_40216);
nor U40572 (N_40572,N_40128,N_40499);
xnor U40573 (N_40573,N_40016,N_40226);
xor U40574 (N_40574,N_40201,N_40466);
nand U40575 (N_40575,N_40287,N_40247);
nor U40576 (N_40576,N_40133,N_40417);
nor U40577 (N_40577,N_40235,N_40289);
nand U40578 (N_40578,N_40214,N_40432);
nand U40579 (N_40579,N_40017,N_40478);
nand U40580 (N_40580,N_40228,N_40167);
and U40581 (N_40581,N_40107,N_40314);
nand U40582 (N_40582,N_40439,N_40178);
nor U40583 (N_40583,N_40379,N_40282);
or U40584 (N_40584,N_40491,N_40225);
xnor U40585 (N_40585,N_40001,N_40317);
or U40586 (N_40586,N_40497,N_40345);
and U40587 (N_40587,N_40134,N_40428);
nand U40588 (N_40588,N_40184,N_40444);
and U40589 (N_40589,N_40366,N_40024);
nor U40590 (N_40590,N_40224,N_40170);
and U40591 (N_40591,N_40192,N_40372);
xnor U40592 (N_40592,N_40357,N_40490);
or U40593 (N_40593,N_40076,N_40043);
nor U40594 (N_40594,N_40120,N_40262);
or U40595 (N_40595,N_40425,N_40137);
nand U40596 (N_40596,N_40056,N_40384);
and U40597 (N_40597,N_40005,N_40275);
and U40598 (N_40598,N_40419,N_40215);
xnor U40599 (N_40599,N_40197,N_40408);
xor U40600 (N_40600,N_40290,N_40211);
nor U40601 (N_40601,N_40391,N_40333);
and U40602 (N_40602,N_40095,N_40080);
or U40603 (N_40603,N_40081,N_40181);
or U40604 (N_40604,N_40227,N_40040);
xnor U40605 (N_40605,N_40036,N_40148);
and U40606 (N_40606,N_40460,N_40469);
and U40607 (N_40607,N_40033,N_40091);
nor U40608 (N_40608,N_40369,N_40246);
xnor U40609 (N_40609,N_40267,N_40110);
or U40610 (N_40610,N_40198,N_40212);
nand U40611 (N_40611,N_40321,N_40194);
or U40612 (N_40612,N_40489,N_40498);
and U40613 (N_40613,N_40217,N_40443);
nor U40614 (N_40614,N_40383,N_40114);
nor U40615 (N_40615,N_40452,N_40338);
or U40616 (N_40616,N_40121,N_40157);
xor U40617 (N_40617,N_40143,N_40427);
nand U40618 (N_40618,N_40066,N_40175);
xor U40619 (N_40619,N_40113,N_40341);
xnor U40620 (N_40620,N_40237,N_40297);
or U40621 (N_40621,N_40108,N_40328);
nor U40622 (N_40622,N_40238,N_40309);
or U40623 (N_40623,N_40481,N_40191);
and U40624 (N_40624,N_40352,N_40385);
xnor U40625 (N_40625,N_40316,N_40023);
nor U40626 (N_40626,N_40404,N_40390);
nor U40627 (N_40627,N_40003,N_40483);
nor U40628 (N_40628,N_40241,N_40039);
nor U40629 (N_40629,N_40331,N_40470);
nor U40630 (N_40630,N_40118,N_40493);
xor U40631 (N_40631,N_40272,N_40326);
nand U40632 (N_40632,N_40047,N_40465);
and U40633 (N_40633,N_40055,N_40433);
or U40634 (N_40634,N_40334,N_40392);
or U40635 (N_40635,N_40195,N_40278);
and U40636 (N_40636,N_40088,N_40180);
and U40637 (N_40637,N_40342,N_40285);
nand U40638 (N_40638,N_40100,N_40136);
or U40639 (N_40639,N_40071,N_40223);
nor U40640 (N_40640,N_40266,N_40388);
nor U40641 (N_40641,N_40032,N_40422);
nor U40642 (N_40642,N_40343,N_40429);
or U40643 (N_40643,N_40205,N_40041);
or U40644 (N_40644,N_40487,N_40213);
or U40645 (N_40645,N_40303,N_40322);
and U40646 (N_40646,N_40015,N_40239);
and U40647 (N_40647,N_40154,N_40093);
nand U40648 (N_40648,N_40323,N_40029);
nand U40649 (N_40649,N_40381,N_40155);
or U40650 (N_40650,N_40401,N_40038);
nor U40651 (N_40651,N_40090,N_40222);
xnor U40652 (N_40652,N_40318,N_40455);
and U40653 (N_40653,N_40031,N_40068);
nand U40654 (N_40654,N_40221,N_40486);
and U40655 (N_40655,N_40052,N_40413);
and U40656 (N_40656,N_40159,N_40067);
xor U40657 (N_40657,N_40210,N_40264);
xor U40658 (N_40658,N_40368,N_40112);
and U40659 (N_40659,N_40411,N_40437);
or U40660 (N_40660,N_40456,N_40045);
xnor U40661 (N_40661,N_40097,N_40069);
nor U40662 (N_40662,N_40018,N_40012);
or U40663 (N_40663,N_40361,N_40079);
nand U40664 (N_40664,N_40409,N_40135);
nand U40665 (N_40665,N_40105,N_40253);
and U40666 (N_40666,N_40362,N_40348);
nand U40667 (N_40667,N_40492,N_40115);
or U40668 (N_40668,N_40395,N_40336);
nand U40669 (N_40669,N_40283,N_40025);
xor U40670 (N_40670,N_40440,N_40187);
or U40671 (N_40671,N_40132,N_40242);
or U40672 (N_40672,N_40475,N_40280);
nor U40673 (N_40673,N_40463,N_40096);
and U40674 (N_40674,N_40240,N_40286);
or U40675 (N_40675,N_40202,N_40453);
xnor U40676 (N_40676,N_40393,N_40365);
xor U40677 (N_40677,N_40203,N_40123);
nand U40678 (N_40678,N_40377,N_40468);
and U40679 (N_40679,N_40268,N_40271);
xnor U40680 (N_40680,N_40471,N_40306);
or U40681 (N_40681,N_40457,N_40127);
and U40682 (N_40682,N_40396,N_40158);
or U40683 (N_40683,N_40488,N_40261);
nand U40684 (N_40684,N_40082,N_40233);
xor U40685 (N_40685,N_40231,N_40249);
nand U40686 (N_40686,N_40421,N_40019);
nor U40687 (N_40687,N_40448,N_40389);
nor U40688 (N_40688,N_40146,N_40245);
and U40689 (N_40689,N_40335,N_40313);
or U40690 (N_40690,N_40307,N_40185);
xor U40691 (N_40691,N_40273,N_40340);
nor U40692 (N_40692,N_40347,N_40124);
xor U40693 (N_40693,N_40251,N_40403);
and U40694 (N_40694,N_40295,N_40086);
and U40695 (N_40695,N_40407,N_40329);
or U40696 (N_40696,N_40355,N_40057);
nand U40697 (N_40697,N_40009,N_40059);
nor U40698 (N_40698,N_40060,N_40258);
or U40699 (N_40699,N_40294,N_40410);
nand U40700 (N_40700,N_40130,N_40451);
xnor U40701 (N_40701,N_40089,N_40349);
or U40702 (N_40702,N_40072,N_40265);
xor U40703 (N_40703,N_40337,N_40062);
or U40704 (N_40704,N_40200,N_40050);
or U40705 (N_40705,N_40496,N_40405);
nand U40706 (N_40706,N_40472,N_40344);
xnor U40707 (N_40707,N_40004,N_40077);
xnor U40708 (N_40708,N_40484,N_40296);
nand U40709 (N_40709,N_40399,N_40177);
or U40710 (N_40710,N_40350,N_40109);
and U40711 (N_40711,N_40367,N_40269);
or U40712 (N_40712,N_40319,N_40196);
or U40713 (N_40713,N_40430,N_40254);
and U40714 (N_40714,N_40311,N_40171);
or U40715 (N_40715,N_40300,N_40220);
or U40716 (N_40716,N_40320,N_40308);
or U40717 (N_40717,N_40058,N_40243);
or U40718 (N_40718,N_40414,N_40204);
and U40719 (N_40719,N_40356,N_40011);
or U40720 (N_40720,N_40142,N_40053);
nand U40721 (N_40721,N_40418,N_40208);
nand U40722 (N_40722,N_40152,N_40161);
nand U40723 (N_40723,N_40476,N_40324);
nand U40724 (N_40724,N_40073,N_40151);
and U40725 (N_40725,N_40106,N_40310);
xor U40726 (N_40726,N_40139,N_40122);
and U40727 (N_40727,N_40166,N_40084);
nand U40728 (N_40728,N_40190,N_40229);
or U40729 (N_40729,N_40284,N_40435);
xnor U40730 (N_40730,N_40252,N_40044);
xnor U40731 (N_40731,N_40006,N_40173);
xnor U40732 (N_40732,N_40454,N_40141);
nor U40733 (N_40733,N_40374,N_40126);
nor U40734 (N_40734,N_40049,N_40244);
nor U40735 (N_40735,N_40257,N_40065);
or U40736 (N_40736,N_40010,N_40485);
and U40737 (N_40737,N_40007,N_40458);
xor U40738 (N_40738,N_40236,N_40406);
xor U40739 (N_40739,N_40098,N_40000);
or U40740 (N_40740,N_40162,N_40279);
xor U40741 (N_40741,N_40400,N_40255);
or U40742 (N_40742,N_40346,N_40387);
nand U40743 (N_40743,N_40206,N_40020);
nand U40744 (N_40744,N_40138,N_40358);
nand U40745 (N_40745,N_40302,N_40291);
nand U40746 (N_40746,N_40305,N_40339);
nand U40747 (N_40747,N_40299,N_40351);
and U40748 (N_40748,N_40477,N_40438);
and U40749 (N_40749,N_40375,N_40473);
nand U40750 (N_40750,N_40372,N_40399);
and U40751 (N_40751,N_40492,N_40372);
nor U40752 (N_40752,N_40376,N_40229);
nor U40753 (N_40753,N_40305,N_40177);
and U40754 (N_40754,N_40465,N_40365);
nor U40755 (N_40755,N_40154,N_40378);
or U40756 (N_40756,N_40010,N_40251);
nand U40757 (N_40757,N_40273,N_40271);
xnor U40758 (N_40758,N_40190,N_40203);
nor U40759 (N_40759,N_40076,N_40265);
xor U40760 (N_40760,N_40472,N_40266);
and U40761 (N_40761,N_40476,N_40448);
xor U40762 (N_40762,N_40080,N_40406);
nand U40763 (N_40763,N_40344,N_40426);
or U40764 (N_40764,N_40418,N_40211);
nand U40765 (N_40765,N_40297,N_40411);
or U40766 (N_40766,N_40209,N_40273);
or U40767 (N_40767,N_40220,N_40007);
nand U40768 (N_40768,N_40240,N_40018);
xor U40769 (N_40769,N_40353,N_40087);
and U40770 (N_40770,N_40163,N_40097);
nand U40771 (N_40771,N_40304,N_40093);
nor U40772 (N_40772,N_40280,N_40304);
and U40773 (N_40773,N_40206,N_40183);
nor U40774 (N_40774,N_40231,N_40247);
nand U40775 (N_40775,N_40435,N_40188);
xnor U40776 (N_40776,N_40066,N_40228);
nor U40777 (N_40777,N_40125,N_40187);
and U40778 (N_40778,N_40165,N_40382);
or U40779 (N_40779,N_40451,N_40345);
nor U40780 (N_40780,N_40499,N_40152);
nor U40781 (N_40781,N_40330,N_40143);
nand U40782 (N_40782,N_40178,N_40113);
or U40783 (N_40783,N_40062,N_40069);
and U40784 (N_40784,N_40374,N_40245);
nand U40785 (N_40785,N_40019,N_40418);
or U40786 (N_40786,N_40369,N_40466);
and U40787 (N_40787,N_40405,N_40358);
and U40788 (N_40788,N_40449,N_40019);
nand U40789 (N_40789,N_40365,N_40410);
and U40790 (N_40790,N_40096,N_40115);
or U40791 (N_40791,N_40205,N_40135);
nand U40792 (N_40792,N_40155,N_40334);
nand U40793 (N_40793,N_40302,N_40416);
nor U40794 (N_40794,N_40208,N_40269);
xor U40795 (N_40795,N_40438,N_40376);
nor U40796 (N_40796,N_40033,N_40019);
or U40797 (N_40797,N_40075,N_40300);
or U40798 (N_40798,N_40155,N_40416);
xnor U40799 (N_40799,N_40153,N_40033);
and U40800 (N_40800,N_40358,N_40274);
or U40801 (N_40801,N_40194,N_40254);
xor U40802 (N_40802,N_40112,N_40213);
nand U40803 (N_40803,N_40337,N_40272);
nor U40804 (N_40804,N_40180,N_40395);
nand U40805 (N_40805,N_40426,N_40463);
nand U40806 (N_40806,N_40295,N_40395);
or U40807 (N_40807,N_40003,N_40245);
xnor U40808 (N_40808,N_40433,N_40095);
nand U40809 (N_40809,N_40299,N_40489);
nor U40810 (N_40810,N_40360,N_40100);
nand U40811 (N_40811,N_40087,N_40213);
xor U40812 (N_40812,N_40204,N_40273);
nor U40813 (N_40813,N_40338,N_40004);
nor U40814 (N_40814,N_40163,N_40141);
or U40815 (N_40815,N_40266,N_40341);
or U40816 (N_40816,N_40287,N_40161);
xnor U40817 (N_40817,N_40275,N_40136);
nand U40818 (N_40818,N_40258,N_40346);
and U40819 (N_40819,N_40112,N_40162);
nor U40820 (N_40820,N_40024,N_40325);
nor U40821 (N_40821,N_40330,N_40418);
and U40822 (N_40822,N_40416,N_40405);
xor U40823 (N_40823,N_40386,N_40002);
nand U40824 (N_40824,N_40239,N_40236);
and U40825 (N_40825,N_40316,N_40320);
nand U40826 (N_40826,N_40019,N_40445);
nand U40827 (N_40827,N_40032,N_40039);
nand U40828 (N_40828,N_40201,N_40322);
or U40829 (N_40829,N_40462,N_40378);
nand U40830 (N_40830,N_40191,N_40306);
xnor U40831 (N_40831,N_40198,N_40281);
nor U40832 (N_40832,N_40184,N_40372);
nand U40833 (N_40833,N_40446,N_40404);
xnor U40834 (N_40834,N_40327,N_40007);
nor U40835 (N_40835,N_40058,N_40263);
nor U40836 (N_40836,N_40267,N_40323);
nor U40837 (N_40837,N_40108,N_40415);
nand U40838 (N_40838,N_40056,N_40028);
nor U40839 (N_40839,N_40423,N_40145);
xnor U40840 (N_40840,N_40040,N_40342);
nor U40841 (N_40841,N_40186,N_40356);
xor U40842 (N_40842,N_40210,N_40421);
nand U40843 (N_40843,N_40173,N_40201);
nor U40844 (N_40844,N_40001,N_40153);
nor U40845 (N_40845,N_40316,N_40024);
xor U40846 (N_40846,N_40273,N_40059);
xnor U40847 (N_40847,N_40009,N_40198);
and U40848 (N_40848,N_40246,N_40113);
and U40849 (N_40849,N_40196,N_40091);
nor U40850 (N_40850,N_40483,N_40313);
xor U40851 (N_40851,N_40481,N_40071);
xnor U40852 (N_40852,N_40308,N_40073);
nor U40853 (N_40853,N_40230,N_40475);
and U40854 (N_40854,N_40190,N_40155);
nor U40855 (N_40855,N_40026,N_40020);
and U40856 (N_40856,N_40496,N_40441);
nand U40857 (N_40857,N_40199,N_40187);
nor U40858 (N_40858,N_40351,N_40286);
nand U40859 (N_40859,N_40367,N_40118);
nand U40860 (N_40860,N_40380,N_40255);
or U40861 (N_40861,N_40163,N_40189);
nand U40862 (N_40862,N_40178,N_40210);
nand U40863 (N_40863,N_40143,N_40347);
nor U40864 (N_40864,N_40026,N_40308);
or U40865 (N_40865,N_40122,N_40312);
xor U40866 (N_40866,N_40467,N_40432);
nand U40867 (N_40867,N_40145,N_40403);
xor U40868 (N_40868,N_40194,N_40263);
and U40869 (N_40869,N_40196,N_40009);
xor U40870 (N_40870,N_40274,N_40200);
nor U40871 (N_40871,N_40148,N_40206);
or U40872 (N_40872,N_40285,N_40081);
nor U40873 (N_40873,N_40274,N_40323);
nand U40874 (N_40874,N_40309,N_40039);
and U40875 (N_40875,N_40305,N_40047);
and U40876 (N_40876,N_40007,N_40260);
nor U40877 (N_40877,N_40336,N_40344);
and U40878 (N_40878,N_40033,N_40050);
nor U40879 (N_40879,N_40017,N_40311);
or U40880 (N_40880,N_40015,N_40046);
nor U40881 (N_40881,N_40447,N_40192);
nor U40882 (N_40882,N_40447,N_40138);
xor U40883 (N_40883,N_40314,N_40089);
or U40884 (N_40884,N_40205,N_40026);
and U40885 (N_40885,N_40150,N_40224);
or U40886 (N_40886,N_40183,N_40093);
nor U40887 (N_40887,N_40001,N_40089);
nand U40888 (N_40888,N_40124,N_40324);
nor U40889 (N_40889,N_40068,N_40136);
nand U40890 (N_40890,N_40485,N_40255);
or U40891 (N_40891,N_40396,N_40406);
or U40892 (N_40892,N_40257,N_40279);
and U40893 (N_40893,N_40281,N_40026);
nand U40894 (N_40894,N_40348,N_40359);
nor U40895 (N_40895,N_40310,N_40402);
nand U40896 (N_40896,N_40386,N_40040);
nand U40897 (N_40897,N_40255,N_40137);
nor U40898 (N_40898,N_40162,N_40060);
nor U40899 (N_40899,N_40419,N_40382);
nand U40900 (N_40900,N_40074,N_40137);
or U40901 (N_40901,N_40202,N_40268);
nor U40902 (N_40902,N_40025,N_40201);
nor U40903 (N_40903,N_40456,N_40082);
and U40904 (N_40904,N_40172,N_40408);
nor U40905 (N_40905,N_40293,N_40155);
or U40906 (N_40906,N_40274,N_40350);
and U40907 (N_40907,N_40140,N_40267);
and U40908 (N_40908,N_40010,N_40427);
xnor U40909 (N_40909,N_40234,N_40116);
and U40910 (N_40910,N_40476,N_40488);
nor U40911 (N_40911,N_40192,N_40236);
nor U40912 (N_40912,N_40450,N_40110);
nand U40913 (N_40913,N_40084,N_40486);
or U40914 (N_40914,N_40432,N_40408);
nand U40915 (N_40915,N_40121,N_40498);
and U40916 (N_40916,N_40441,N_40338);
nand U40917 (N_40917,N_40491,N_40384);
nand U40918 (N_40918,N_40040,N_40014);
or U40919 (N_40919,N_40178,N_40067);
or U40920 (N_40920,N_40220,N_40028);
or U40921 (N_40921,N_40056,N_40100);
nor U40922 (N_40922,N_40191,N_40437);
xor U40923 (N_40923,N_40167,N_40208);
xnor U40924 (N_40924,N_40307,N_40176);
and U40925 (N_40925,N_40391,N_40354);
nor U40926 (N_40926,N_40200,N_40420);
and U40927 (N_40927,N_40040,N_40290);
nand U40928 (N_40928,N_40071,N_40486);
xor U40929 (N_40929,N_40322,N_40068);
xor U40930 (N_40930,N_40031,N_40104);
and U40931 (N_40931,N_40198,N_40064);
nand U40932 (N_40932,N_40018,N_40408);
nor U40933 (N_40933,N_40344,N_40486);
nand U40934 (N_40934,N_40204,N_40456);
nor U40935 (N_40935,N_40068,N_40212);
nor U40936 (N_40936,N_40332,N_40241);
or U40937 (N_40937,N_40476,N_40387);
or U40938 (N_40938,N_40447,N_40457);
nor U40939 (N_40939,N_40418,N_40180);
nand U40940 (N_40940,N_40026,N_40314);
nand U40941 (N_40941,N_40159,N_40215);
nor U40942 (N_40942,N_40328,N_40174);
nand U40943 (N_40943,N_40389,N_40341);
xor U40944 (N_40944,N_40349,N_40459);
and U40945 (N_40945,N_40373,N_40321);
or U40946 (N_40946,N_40255,N_40468);
or U40947 (N_40947,N_40016,N_40260);
nor U40948 (N_40948,N_40299,N_40368);
xnor U40949 (N_40949,N_40339,N_40284);
xnor U40950 (N_40950,N_40191,N_40384);
and U40951 (N_40951,N_40227,N_40110);
and U40952 (N_40952,N_40036,N_40460);
or U40953 (N_40953,N_40187,N_40365);
xor U40954 (N_40954,N_40277,N_40498);
xnor U40955 (N_40955,N_40323,N_40421);
nor U40956 (N_40956,N_40431,N_40481);
xnor U40957 (N_40957,N_40462,N_40402);
or U40958 (N_40958,N_40051,N_40243);
xnor U40959 (N_40959,N_40399,N_40206);
or U40960 (N_40960,N_40346,N_40324);
or U40961 (N_40961,N_40380,N_40306);
xor U40962 (N_40962,N_40332,N_40245);
nor U40963 (N_40963,N_40267,N_40498);
nand U40964 (N_40964,N_40233,N_40143);
xnor U40965 (N_40965,N_40290,N_40356);
xnor U40966 (N_40966,N_40015,N_40100);
or U40967 (N_40967,N_40296,N_40003);
or U40968 (N_40968,N_40075,N_40097);
and U40969 (N_40969,N_40389,N_40466);
nand U40970 (N_40970,N_40097,N_40249);
nand U40971 (N_40971,N_40450,N_40426);
and U40972 (N_40972,N_40026,N_40186);
nand U40973 (N_40973,N_40437,N_40054);
and U40974 (N_40974,N_40094,N_40256);
nand U40975 (N_40975,N_40115,N_40145);
nor U40976 (N_40976,N_40200,N_40042);
or U40977 (N_40977,N_40184,N_40110);
xor U40978 (N_40978,N_40313,N_40348);
nand U40979 (N_40979,N_40293,N_40410);
nor U40980 (N_40980,N_40276,N_40441);
and U40981 (N_40981,N_40292,N_40362);
xnor U40982 (N_40982,N_40004,N_40140);
and U40983 (N_40983,N_40285,N_40100);
nor U40984 (N_40984,N_40424,N_40117);
nand U40985 (N_40985,N_40207,N_40079);
nor U40986 (N_40986,N_40388,N_40310);
and U40987 (N_40987,N_40286,N_40263);
and U40988 (N_40988,N_40057,N_40372);
nor U40989 (N_40989,N_40098,N_40291);
nor U40990 (N_40990,N_40108,N_40376);
and U40991 (N_40991,N_40415,N_40396);
and U40992 (N_40992,N_40453,N_40264);
and U40993 (N_40993,N_40284,N_40206);
nor U40994 (N_40994,N_40252,N_40153);
and U40995 (N_40995,N_40349,N_40458);
nor U40996 (N_40996,N_40392,N_40467);
nand U40997 (N_40997,N_40155,N_40094);
or U40998 (N_40998,N_40073,N_40480);
xor U40999 (N_40999,N_40427,N_40106);
nand U41000 (N_41000,N_40699,N_40824);
nor U41001 (N_41001,N_40841,N_40500);
xor U41002 (N_41002,N_40663,N_40732);
xor U41003 (N_41003,N_40795,N_40875);
nor U41004 (N_41004,N_40952,N_40957);
or U41005 (N_41005,N_40705,N_40560);
nor U41006 (N_41006,N_40870,N_40501);
xnor U41007 (N_41007,N_40528,N_40899);
nor U41008 (N_41008,N_40770,N_40558);
nor U41009 (N_41009,N_40533,N_40755);
nor U41010 (N_41010,N_40918,N_40610);
nand U41011 (N_41011,N_40849,N_40802);
or U41012 (N_41012,N_40966,N_40903);
or U41013 (N_41013,N_40972,N_40617);
and U41014 (N_41014,N_40974,N_40778);
nor U41015 (N_41015,N_40695,N_40806);
and U41016 (N_41016,N_40808,N_40730);
or U41017 (N_41017,N_40604,N_40557);
nand U41018 (N_41018,N_40947,N_40584);
nand U41019 (N_41019,N_40503,N_40780);
xor U41020 (N_41020,N_40840,N_40550);
and U41021 (N_41021,N_40864,N_40999);
or U41022 (N_41022,N_40735,N_40692);
nor U41023 (N_41023,N_40553,N_40860);
and U41024 (N_41024,N_40843,N_40862);
xor U41025 (N_41025,N_40998,N_40794);
nand U41026 (N_41026,N_40810,N_40716);
nand U41027 (N_41027,N_40512,N_40920);
or U41028 (N_41028,N_40856,N_40772);
and U41029 (N_41029,N_40836,N_40675);
or U41030 (N_41030,N_40767,N_40725);
and U41031 (N_41031,N_40603,N_40753);
and U41032 (N_41032,N_40756,N_40906);
and U41033 (N_41033,N_40956,N_40654);
nor U41034 (N_41034,N_40554,N_40514);
and U41035 (N_41035,N_40791,N_40750);
xor U41036 (N_41036,N_40986,N_40835);
nand U41037 (N_41037,N_40764,N_40607);
and U41038 (N_41038,N_40917,N_40988);
nand U41039 (N_41039,N_40520,N_40948);
nand U41040 (N_41040,N_40524,N_40763);
xnor U41041 (N_41041,N_40624,N_40653);
or U41042 (N_41042,N_40890,N_40967);
nor U41043 (N_41043,N_40537,N_40789);
nor U41044 (N_41044,N_40646,N_40896);
and U41045 (N_41045,N_40535,N_40713);
nand U41046 (N_41046,N_40641,N_40911);
nor U41047 (N_41047,N_40546,N_40830);
nand U41048 (N_41048,N_40828,N_40680);
nor U41049 (N_41049,N_40964,N_40597);
nor U41050 (N_41050,N_40958,N_40666);
xor U41051 (N_41051,N_40605,N_40814);
or U41052 (N_41052,N_40709,N_40950);
or U41053 (N_41053,N_40823,N_40724);
nor U41054 (N_41054,N_40635,N_40609);
nand U41055 (N_41055,N_40518,N_40880);
and U41056 (N_41056,N_40575,N_40866);
xor U41057 (N_41057,N_40572,N_40698);
xnor U41058 (N_41058,N_40811,N_40768);
and U41059 (N_41059,N_40519,N_40869);
or U41060 (N_41060,N_40733,N_40844);
xnor U41061 (N_41061,N_40509,N_40594);
or U41062 (N_41062,N_40687,N_40639);
nand U41063 (N_41063,N_40914,N_40701);
nor U41064 (N_41064,N_40760,N_40598);
or U41065 (N_41065,N_40962,N_40702);
or U41066 (N_41066,N_40686,N_40515);
xor U41067 (N_41067,N_40505,N_40939);
nand U41068 (N_41068,N_40771,N_40523);
and U41069 (N_41069,N_40997,N_40983);
and U41070 (N_41070,N_40961,N_40513);
xnor U41071 (N_41071,N_40743,N_40921);
or U41072 (N_41072,N_40820,N_40637);
and U41073 (N_41073,N_40766,N_40803);
xor U41074 (N_41074,N_40993,N_40989);
or U41075 (N_41075,N_40992,N_40944);
xor U41076 (N_41076,N_40670,N_40718);
xnor U41077 (N_41077,N_40877,N_40671);
nor U41078 (N_41078,N_40714,N_40951);
nand U41079 (N_41079,N_40865,N_40850);
nor U41080 (N_41080,N_40704,N_40925);
xor U41081 (N_41081,N_40879,N_40946);
or U41082 (N_41082,N_40991,N_40728);
nand U41083 (N_41083,N_40867,N_40818);
nand U41084 (N_41084,N_40996,N_40583);
or U41085 (N_41085,N_40874,N_40812);
xor U41086 (N_41086,N_40719,N_40532);
xor U41087 (N_41087,N_40580,N_40590);
or U41088 (N_41088,N_40536,N_40600);
xnor U41089 (N_41089,N_40531,N_40589);
and U41090 (N_41090,N_40749,N_40542);
xnor U41091 (N_41091,N_40676,N_40855);
and U41092 (N_41092,N_40540,N_40545);
and U41093 (N_41093,N_40656,N_40696);
nand U41094 (N_41094,N_40504,N_40759);
xnor U41095 (N_41095,N_40734,N_40723);
nor U41096 (N_41096,N_40662,N_40990);
nand U41097 (N_41097,N_40745,N_40930);
or U41098 (N_41098,N_40995,N_40897);
xnor U41099 (N_41099,N_40678,N_40574);
nor U41100 (N_41100,N_40926,N_40758);
and U41101 (N_41101,N_40581,N_40717);
and U41102 (N_41102,N_40851,N_40522);
nand U41103 (N_41103,N_40510,N_40891);
nor U41104 (N_41104,N_40555,N_40621);
nand U41105 (N_41105,N_40538,N_40736);
or U41106 (N_41106,N_40738,N_40541);
and U41107 (N_41107,N_40977,N_40661);
and U41108 (N_41108,N_40819,N_40650);
nand U41109 (N_41109,N_40544,N_40534);
nor U41110 (N_41110,N_40813,N_40618);
nand U41111 (N_41111,N_40588,N_40871);
nand U41112 (N_41112,N_40683,N_40682);
and U41113 (N_41113,N_40585,N_40579);
or U41114 (N_41114,N_40747,N_40796);
nand U41115 (N_41115,N_40872,N_40616);
xor U41116 (N_41116,N_40591,N_40882);
nor U41117 (N_41117,N_40798,N_40779);
nand U41118 (N_41118,N_40797,N_40691);
nor U41119 (N_41119,N_40774,N_40614);
xor U41120 (N_41120,N_40935,N_40907);
or U41121 (N_41121,N_40729,N_40612);
nor U41122 (N_41122,N_40506,N_40900);
nand U41123 (N_41123,N_40634,N_40684);
and U41124 (N_41124,N_40804,N_40673);
xnor U41125 (N_41125,N_40943,N_40690);
nor U41126 (N_41126,N_40984,N_40809);
nor U41127 (N_41127,N_40994,N_40721);
xor U41128 (N_41128,N_40878,N_40905);
and U41129 (N_41129,N_40884,N_40625);
or U41130 (N_41130,N_40885,N_40936);
and U41131 (N_41131,N_40576,N_40668);
and U41132 (N_41132,N_40978,N_40655);
or U41133 (N_41133,N_40910,N_40652);
xor U41134 (N_41134,N_40693,N_40893);
and U41135 (N_41135,N_40552,N_40769);
or U41136 (N_41136,N_40599,N_40715);
nor U41137 (N_41137,N_40568,N_40570);
or U41138 (N_41138,N_40927,N_40848);
nand U41139 (N_41139,N_40697,N_40628);
or U41140 (N_41140,N_40799,N_40822);
nand U41141 (N_41141,N_40633,N_40915);
xor U41142 (N_41142,N_40765,N_40648);
xor U41143 (N_41143,N_40839,N_40832);
nor U41144 (N_41144,N_40657,N_40960);
or U41145 (N_41145,N_40741,N_40945);
or U41146 (N_41146,N_40596,N_40928);
or U41147 (N_41147,N_40629,N_40913);
and U41148 (N_41148,N_40527,N_40782);
xor U41149 (N_41149,N_40924,N_40601);
xnor U41150 (N_41150,N_40644,N_40543);
xor U41151 (N_41151,N_40786,N_40846);
nand U41152 (N_41152,N_40619,N_40852);
and U41153 (N_41153,N_40593,N_40602);
xor U41154 (N_41154,N_40788,N_40980);
or U41155 (N_41155,N_40923,N_40929);
xnor U41156 (N_41156,N_40615,N_40831);
nor U41157 (N_41157,N_40858,N_40508);
xnor U41158 (N_41158,N_40502,N_40816);
xor U41159 (N_41159,N_40722,N_40595);
or U41160 (N_41160,N_40742,N_40526);
nand U41161 (N_41161,N_40651,N_40941);
nor U41162 (N_41162,N_40821,N_40773);
nor U41163 (N_41163,N_40746,N_40672);
and U41164 (N_41164,N_40551,N_40815);
nor U41165 (N_41165,N_40620,N_40606);
xor U41166 (N_41166,N_40781,N_40775);
and U41167 (N_41167,N_40562,N_40712);
nand U41168 (N_41168,N_40710,N_40530);
xor U41169 (N_41169,N_40507,N_40965);
nor U41170 (N_41170,N_40868,N_40976);
nor U41171 (N_41171,N_40790,N_40638);
and U41172 (N_41172,N_40883,N_40969);
and U41173 (N_41173,N_40861,N_40622);
nand U41174 (N_41174,N_40665,N_40955);
and U41175 (N_41175,N_40688,N_40985);
xnor U41176 (N_41176,N_40825,N_40744);
xor U41177 (N_41177,N_40694,N_40981);
and U41178 (N_41178,N_40889,N_40739);
nand U41179 (N_41179,N_40511,N_40640);
xnor U41180 (N_41180,N_40959,N_40829);
or U41181 (N_41181,N_40833,N_40854);
xnor U41182 (N_41182,N_40982,N_40556);
and U41183 (N_41183,N_40548,N_40949);
xor U41184 (N_41184,N_40707,N_40569);
and U41185 (N_41185,N_40807,N_40863);
or U41186 (N_41186,N_40549,N_40817);
nor U41187 (N_41187,N_40892,N_40901);
nand U41188 (N_41188,N_40922,N_40578);
nand U41189 (N_41189,N_40565,N_40626);
nand U41190 (N_41190,N_40887,N_40751);
xnor U41191 (N_41191,N_40658,N_40636);
xor U41192 (N_41192,N_40592,N_40934);
nand U41193 (N_41193,N_40571,N_40559);
nor U41194 (N_41194,N_40630,N_40970);
xnor U41195 (N_41195,N_40529,N_40837);
xnor U41196 (N_41196,N_40853,N_40664);
or U41197 (N_41197,N_40577,N_40834);
xor U41198 (N_41198,N_40669,N_40968);
nor U41199 (N_41199,N_40752,N_40902);
or U41200 (N_41200,N_40586,N_40873);
xor U41201 (N_41201,N_40792,N_40800);
nand U41202 (N_41202,N_40979,N_40582);
nand U41203 (N_41203,N_40826,N_40881);
and U41204 (N_41204,N_40631,N_40916);
xnor U41205 (N_41205,N_40787,N_40783);
xnor U41206 (N_41206,N_40613,N_40933);
or U41207 (N_41207,N_40627,N_40908);
or U41208 (N_41208,N_40942,N_40706);
nor U41209 (N_41209,N_40754,N_40859);
or U41210 (N_41210,N_40937,N_40679);
or U41211 (N_41211,N_40805,N_40777);
nor U41212 (N_41212,N_40931,N_40573);
nand U41213 (N_41213,N_40793,N_40726);
nand U41214 (N_41214,N_40708,N_40784);
nand U41215 (N_41215,N_40703,N_40971);
or U41216 (N_41216,N_40660,N_40827);
or U41217 (N_41217,N_40857,N_40737);
nand U41218 (N_41218,N_40727,N_40894);
nand U41219 (N_41219,N_40685,N_40517);
nand U41220 (N_41220,N_40642,N_40731);
and U41221 (N_41221,N_40711,N_40674);
or U41222 (N_41222,N_40566,N_40845);
or U41223 (N_41223,N_40785,N_40521);
xor U41224 (N_41224,N_40938,N_40623);
nand U41225 (N_41225,N_40895,N_40876);
nor U41226 (N_41226,N_40643,N_40940);
and U41227 (N_41227,N_40898,N_40700);
nand U41228 (N_41228,N_40547,N_40720);
nor U41229 (N_41229,N_40953,N_40838);
xor U41230 (N_41230,N_40847,N_40912);
and U41231 (N_41231,N_40762,N_40516);
nor U41232 (N_41232,N_40904,N_40987);
nor U41233 (N_41233,N_40645,N_40539);
and U41234 (N_41234,N_40909,N_40757);
and U41235 (N_41235,N_40689,N_40667);
and U41236 (N_41236,N_40525,N_40677);
and U41237 (N_41237,N_40564,N_40632);
and U41238 (N_41238,N_40801,N_40567);
xor U41239 (N_41239,N_40748,N_40932);
xor U41240 (N_41240,N_40954,N_40649);
or U41241 (N_41241,N_40776,N_40681);
nand U41242 (N_41242,N_40740,N_40963);
xnor U41243 (N_41243,N_40842,N_40587);
xnor U41244 (N_41244,N_40888,N_40561);
or U41245 (N_41245,N_40611,N_40973);
or U41246 (N_41246,N_40761,N_40659);
and U41247 (N_41247,N_40647,N_40919);
nor U41248 (N_41248,N_40886,N_40608);
xnor U41249 (N_41249,N_40563,N_40975);
nand U41250 (N_41250,N_40705,N_40651);
and U41251 (N_41251,N_40621,N_40848);
nor U41252 (N_41252,N_40554,N_40690);
nor U41253 (N_41253,N_40943,N_40728);
xor U41254 (N_41254,N_40722,N_40525);
xnor U41255 (N_41255,N_40949,N_40709);
xnor U41256 (N_41256,N_40790,N_40700);
and U41257 (N_41257,N_40826,N_40744);
xnor U41258 (N_41258,N_40546,N_40612);
and U41259 (N_41259,N_40845,N_40644);
xor U41260 (N_41260,N_40741,N_40610);
xnor U41261 (N_41261,N_40533,N_40995);
nor U41262 (N_41262,N_40746,N_40941);
and U41263 (N_41263,N_40773,N_40592);
nor U41264 (N_41264,N_40646,N_40966);
or U41265 (N_41265,N_40748,N_40982);
or U41266 (N_41266,N_40964,N_40586);
xor U41267 (N_41267,N_40911,N_40502);
nand U41268 (N_41268,N_40540,N_40701);
nand U41269 (N_41269,N_40877,N_40592);
nor U41270 (N_41270,N_40962,N_40895);
and U41271 (N_41271,N_40907,N_40742);
nor U41272 (N_41272,N_40659,N_40671);
or U41273 (N_41273,N_40718,N_40647);
xor U41274 (N_41274,N_40766,N_40866);
nand U41275 (N_41275,N_40657,N_40766);
nand U41276 (N_41276,N_40821,N_40920);
nor U41277 (N_41277,N_40813,N_40580);
nand U41278 (N_41278,N_40596,N_40772);
nand U41279 (N_41279,N_40568,N_40864);
nand U41280 (N_41280,N_40880,N_40602);
xnor U41281 (N_41281,N_40640,N_40813);
nand U41282 (N_41282,N_40874,N_40987);
or U41283 (N_41283,N_40785,N_40912);
or U41284 (N_41284,N_40662,N_40658);
and U41285 (N_41285,N_40847,N_40824);
nand U41286 (N_41286,N_40646,N_40699);
nand U41287 (N_41287,N_40770,N_40919);
nor U41288 (N_41288,N_40776,N_40782);
and U41289 (N_41289,N_40729,N_40731);
nand U41290 (N_41290,N_40967,N_40900);
xor U41291 (N_41291,N_40902,N_40574);
or U41292 (N_41292,N_40903,N_40825);
and U41293 (N_41293,N_40925,N_40736);
or U41294 (N_41294,N_40711,N_40688);
and U41295 (N_41295,N_40953,N_40770);
xnor U41296 (N_41296,N_40686,N_40881);
xor U41297 (N_41297,N_40812,N_40659);
and U41298 (N_41298,N_40960,N_40965);
xnor U41299 (N_41299,N_40718,N_40907);
nand U41300 (N_41300,N_40818,N_40670);
xnor U41301 (N_41301,N_40567,N_40889);
and U41302 (N_41302,N_40716,N_40925);
nand U41303 (N_41303,N_40708,N_40905);
and U41304 (N_41304,N_40504,N_40565);
nor U41305 (N_41305,N_40541,N_40944);
or U41306 (N_41306,N_40527,N_40726);
nand U41307 (N_41307,N_40998,N_40762);
and U41308 (N_41308,N_40728,N_40889);
nand U41309 (N_41309,N_40974,N_40561);
xor U41310 (N_41310,N_40821,N_40669);
nand U41311 (N_41311,N_40796,N_40986);
and U41312 (N_41312,N_40971,N_40759);
or U41313 (N_41313,N_40981,N_40766);
or U41314 (N_41314,N_40629,N_40748);
or U41315 (N_41315,N_40898,N_40661);
and U41316 (N_41316,N_40712,N_40983);
or U41317 (N_41317,N_40823,N_40622);
nor U41318 (N_41318,N_40842,N_40863);
nand U41319 (N_41319,N_40762,N_40802);
or U41320 (N_41320,N_40796,N_40726);
and U41321 (N_41321,N_40814,N_40925);
xnor U41322 (N_41322,N_40552,N_40748);
xor U41323 (N_41323,N_40902,N_40799);
or U41324 (N_41324,N_40903,N_40852);
or U41325 (N_41325,N_40680,N_40619);
nand U41326 (N_41326,N_40600,N_40974);
nand U41327 (N_41327,N_40889,N_40753);
or U41328 (N_41328,N_40882,N_40914);
nor U41329 (N_41329,N_40865,N_40826);
or U41330 (N_41330,N_40902,N_40660);
or U41331 (N_41331,N_40596,N_40717);
nand U41332 (N_41332,N_40582,N_40897);
xnor U41333 (N_41333,N_40684,N_40582);
nor U41334 (N_41334,N_40830,N_40760);
nand U41335 (N_41335,N_40655,N_40797);
nor U41336 (N_41336,N_40735,N_40769);
and U41337 (N_41337,N_40709,N_40502);
or U41338 (N_41338,N_40615,N_40519);
or U41339 (N_41339,N_40556,N_40677);
and U41340 (N_41340,N_40929,N_40946);
nor U41341 (N_41341,N_40594,N_40597);
or U41342 (N_41342,N_40650,N_40704);
or U41343 (N_41343,N_40822,N_40627);
or U41344 (N_41344,N_40505,N_40546);
and U41345 (N_41345,N_40699,N_40955);
and U41346 (N_41346,N_40874,N_40809);
nand U41347 (N_41347,N_40700,N_40891);
or U41348 (N_41348,N_40631,N_40669);
or U41349 (N_41349,N_40917,N_40700);
nand U41350 (N_41350,N_40589,N_40955);
nand U41351 (N_41351,N_40756,N_40723);
and U41352 (N_41352,N_40755,N_40961);
nor U41353 (N_41353,N_40996,N_40920);
xor U41354 (N_41354,N_40648,N_40661);
nand U41355 (N_41355,N_40628,N_40927);
or U41356 (N_41356,N_40582,N_40612);
or U41357 (N_41357,N_40850,N_40796);
xor U41358 (N_41358,N_40846,N_40744);
or U41359 (N_41359,N_40647,N_40960);
and U41360 (N_41360,N_40518,N_40971);
nor U41361 (N_41361,N_40792,N_40863);
nor U41362 (N_41362,N_40868,N_40644);
nand U41363 (N_41363,N_40788,N_40888);
or U41364 (N_41364,N_40916,N_40925);
xnor U41365 (N_41365,N_40992,N_40720);
or U41366 (N_41366,N_40636,N_40985);
xor U41367 (N_41367,N_40833,N_40928);
or U41368 (N_41368,N_40801,N_40910);
nor U41369 (N_41369,N_40711,N_40574);
and U41370 (N_41370,N_40557,N_40678);
nor U41371 (N_41371,N_40820,N_40752);
or U41372 (N_41372,N_40862,N_40704);
and U41373 (N_41373,N_40809,N_40750);
nand U41374 (N_41374,N_40532,N_40506);
xnor U41375 (N_41375,N_40702,N_40627);
and U41376 (N_41376,N_40581,N_40720);
and U41377 (N_41377,N_40844,N_40877);
xnor U41378 (N_41378,N_40704,N_40561);
nor U41379 (N_41379,N_40996,N_40718);
and U41380 (N_41380,N_40968,N_40940);
and U41381 (N_41381,N_40956,N_40624);
and U41382 (N_41382,N_40926,N_40825);
or U41383 (N_41383,N_40893,N_40904);
xor U41384 (N_41384,N_40628,N_40775);
nand U41385 (N_41385,N_40526,N_40571);
nor U41386 (N_41386,N_40871,N_40644);
xnor U41387 (N_41387,N_40749,N_40893);
and U41388 (N_41388,N_40759,N_40516);
or U41389 (N_41389,N_40720,N_40816);
nand U41390 (N_41390,N_40633,N_40716);
nand U41391 (N_41391,N_40979,N_40987);
nand U41392 (N_41392,N_40551,N_40749);
nor U41393 (N_41393,N_40750,N_40946);
or U41394 (N_41394,N_40729,N_40949);
and U41395 (N_41395,N_40873,N_40731);
nand U41396 (N_41396,N_40800,N_40697);
or U41397 (N_41397,N_40702,N_40878);
nand U41398 (N_41398,N_40856,N_40999);
or U41399 (N_41399,N_40594,N_40741);
nor U41400 (N_41400,N_40760,N_40679);
or U41401 (N_41401,N_40788,N_40993);
and U41402 (N_41402,N_40909,N_40715);
nand U41403 (N_41403,N_40677,N_40524);
nand U41404 (N_41404,N_40648,N_40613);
nor U41405 (N_41405,N_40886,N_40899);
or U41406 (N_41406,N_40953,N_40620);
or U41407 (N_41407,N_40593,N_40579);
xor U41408 (N_41408,N_40680,N_40690);
xor U41409 (N_41409,N_40611,N_40948);
or U41410 (N_41410,N_40606,N_40943);
nand U41411 (N_41411,N_40620,N_40638);
or U41412 (N_41412,N_40837,N_40685);
or U41413 (N_41413,N_40941,N_40840);
xnor U41414 (N_41414,N_40873,N_40647);
xnor U41415 (N_41415,N_40910,N_40790);
or U41416 (N_41416,N_40959,N_40841);
nor U41417 (N_41417,N_40779,N_40748);
and U41418 (N_41418,N_40723,N_40602);
or U41419 (N_41419,N_40772,N_40826);
xor U41420 (N_41420,N_40533,N_40796);
xnor U41421 (N_41421,N_40617,N_40613);
or U41422 (N_41422,N_40669,N_40598);
xor U41423 (N_41423,N_40733,N_40855);
xnor U41424 (N_41424,N_40745,N_40901);
or U41425 (N_41425,N_40797,N_40917);
or U41426 (N_41426,N_40635,N_40716);
nor U41427 (N_41427,N_40524,N_40511);
nand U41428 (N_41428,N_40685,N_40705);
xor U41429 (N_41429,N_40727,N_40792);
xor U41430 (N_41430,N_40749,N_40629);
xnor U41431 (N_41431,N_40813,N_40515);
or U41432 (N_41432,N_40846,N_40756);
nand U41433 (N_41433,N_40803,N_40703);
xor U41434 (N_41434,N_40928,N_40786);
xnor U41435 (N_41435,N_40941,N_40563);
or U41436 (N_41436,N_40884,N_40651);
and U41437 (N_41437,N_40572,N_40754);
and U41438 (N_41438,N_40610,N_40565);
nor U41439 (N_41439,N_40870,N_40679);
nor U41440 (N_41440,N_40777,N_40886);
and U41441 (N_41441,N_40546,N_40681);
xnor U41442 (N_41442,N_40749,N_40557);
and U41443 (N_41443,N_40958,N_40533);
xor U41444 (N_41444,N_40854,N_40796);
xnor U41445 (N_41445,N_40805,N_40545);
and U41446 (N_41446,N_40714,N_40608);
nor U41447 (N_41447,N_40671,N_40854);
nand U41448 (N_41448,N_40606,N_40924);
and U41449 (N_41449,N_40904,N_40719);
and U41450 (N_41450,N_40886,N_40587);
xor U41451 (N_41451,N_40566,N_40986);
or U41452 (N_41452,N_40709,N_40855);
and U41453 (N_41453,N_40777,N_40993);
and U41454 (N_41454,N_40839,N_40556);
and U41455 (N_41455,N_40794,N_40864);
or U41456 (N_41456,N_40789,N_40906);
nand U41457 (N_41457,N_40688,N_40971);
xor U41458 (N_41458,N_40968,N_40644);
and U41459 (N_41459,N_40602,N_40503);
and U41460 (N_41460,N_40528,N_40943);
nor U41461 (N_41461,N_40877,N_40838);
or U41462 (N_41462,N_40679,N_40591);
and U41463 (N_41463,N_40792,N_40760);
xor U41464 (N_41464,N_40525,N_40596);
and U41465 (N_41465,N_40780,N_40747);
xor U41466 (N_41466,N_40945,N_40933);
nand U41467 (N_41467,N_40678,N_40677);
nand U41468 (N_41468,N_40935,N_40559);
or U41469 (N_41469,N_40588,N_40984);
nor U41470 (N_41470,N_40652,N_40765);
nor U41471 (N_41471,N_40541,N_40865);
or U41472 (N_41472,N_40700,N_40963);
or U41473 (N_41473,N_40939,N_40842);
nand U41474 (N_41474,N_40636,N_40990);
or U41475 (N_41475,N_40795,N_40810);
nand U41476 (N_41476,N_40662,N_40727);
xor U41477 (N_41477,N_40821,N_40887);
or U41478 (N_41478,N_40606,N_40511);
nand U41479 (N_41479,N_40602,N_40820);
and U41480 (N_41480,N_40509,N_40666);
xor U41481 (N_41481,N_40553,N_40655);
and U41482 (N_41482,N_40910,N_40816);
nor U41483 (N_41483,N_40631,N_40650);
xor U41484 (N_41484,N_40510,N_40762);
and U41485 (N_41485,N_40732,N_40876);
or U41486 (N_41486,N_40580,N_40701);
or U41487 (N_41487,N_40597,N_40538);
nor U41488 (N_41488,N_40561,N_40574);
or U41489 (N_41489,N_40596,N_40671);
and U41490 (N_41490,N_40728,N_40644);
nor U41491 (N_41491,N_40610,N_40529);
or U41492 (N_41492,N_40796,N_40678);
nand U41493 (N_41493,N_40865,N_40871);
xnor U41494 (N_41494,N_40869,N_40997);
nor U41495 (N_41495,N_40501,N_40785);
nor U41496 (N_41496,N_40682,N_40946);
nand U41497 (N_41497,N_40600,N_40835);
nor U41498 (N_41498,N_40780,N_40641);
nand U41499 (N_41499,N_40521,N_40523);
nor U41500 (N_41500,N_41191,N_41067);
nor U41501 (N_41501,N_41342,N_41375);
nor U41502 (N_41502,N_41498,N_41247);
nor U41503 (N_41503,N_41369,N_41013);
xor U41504 (N_41504,N_41215,N_41448);
nand U41505 (N_41505,N_41006,N_41050);
and U41506 (N_41506,N_41317,N_41159);
and U41507 (N_41507,N_41051,N_41491);
xor U41508 (N_41508,N_41327,N_41167);
or U41509 (N_41509,N_41269,N_41205);
or U41510 (N_41510,N_41415,N_41461);
and U41511 (N_41511,N_41042,N_41071);
nor U41512 (N_41512,N_41363,N_41329);
and U41513 (N_41513,N_41260,N_41105);
xnor U41514 (N_41514,N_41427,N_41353);
xnor U41515 (N_41515,N_41240,N_41408);
nor U41516 (N_41516,N_41244,N_41397);
nand U41517 (N_41517,N_41401,N_41086);
xor U41518 (N_41518,N_41081,N_41282);
and U41519 (N_41519,N_41058,N_41366);
nor U41520 (N_41520,N_41188,N_41284);
nor U41521 (N_41521,N_41128,N_41177);
or U41522 (N_41522,N_41066,N_41136);
or U41523 (N_41523,N_41253,N_41328);
and U41524 (N_41524,N_41232,N_41277);
nor U41525 (N_41525,N_41256,N_41194);
xor U41526 (N_41526,N_41144,N_41307);
nand U41527 (N_41527,N_41083,N_41481);
nand U41528 (N_41528,N_41039,N_41122);
xnor U41529 (N_41529,N_41103,N_41404);
nand U41530 (N_41530,N_41254,N_41435);
nand U41531 (N_41531,N_41469,N_41044);
nand U41532 (N_41532,N_41093,N_41018);
xor U41533 (N_41533,N_41420,N_41199);
nor U41534 (N_41534,N_41484,N_41280);
and U41535 (N_41535,N_41399,N_41000);
nor U41536 (N_41536,N_41464,N_41162);
and U41537 (N_41537,N_41182,N_41489);
and U41538 (N_41538,N_41080,N_41168);
and U41539 (N_41539,N_41332,N_41387);
nand U41540 (N_41540,N_41364,N_41153);
xor U41541 (N_41541,N_41245,N_41338);
nor U41542 (N_41542,N_41056,N_41088);
nand U41543 (N_41543,N_41019,N_41017);
xnor U41544 (N_41544,N_41474,N_41176);
xnor U41545 (N_41545,N_41041,N_41340);
and U41546 (N_41546,N_41220,N_41362);
and U41547 (N_41547,N_41243,N_41189);
xnor U41548 (N_41548,N_41053,N_41212);
xnor U41549 (N_41549,N_41173,N_41446);
nor U41550 (N_41550,N_41034,N_41003);
and U41551 (N_41551,N_41116,N_41283);
or U41552 (N_41552,N_41270,N_41405);
or U41553 (N_41553,N_41365,N_41371);
nor U41554 (N_41554,N_41023,N_41298);
and U41555 (N_41555,N_41190,N_41110);
xnor U41556 (N_41556,N_41026,N_41303);
xor U41557 (N_41557,N_41265,N_41025);
nand U41558 (N_41558,N_41391,N_41228);
or U41559 (N_41559,N_41268,N_41460);
and U41560 (N_41560,N_41309,N_41216);
nor U41561 (N_41561,N_41314,N_41409);
and U41562 (N_41562,N_41038,N_41402);
nand U41563 (N_41563,N_41074,N_41312);
nand U41564 (N_41564,N_41281,N_41305);
or U41565 (N_41565,N_41131,N_41434);
nand U41566 (N_41566,N_41477,N_41002);
or U41567 (N_41567,N_41331,N_41180);
xnor U41568 (N_41568,N_41288,N_41049);
and U41569 (N_41569,N_41226,N_41478);
xnor U41570 (N_41570,N_41033,N_41463);
or U41571 (N_41571,N_41142,N_41459);
nand U41572 (N_41572,N_41467,N_41293);
nor U41573 (N_41573,N_41152,N_41490);
or U41574 (N_41574,N_41325,N_41135);
xnor U41575 (N_41575,N_41319,N_41470);
nor U41576 (N_41576,N_41137,N_41235);
or U41577 (N_41577,N_41263,N_41246);
nor U41578 (N_41578,N_41424,N_41027);
nand U41579 (N_41579,N_41486,N_41151);
xor U41580 (N_41580,N_41272,N_41451);
nor U41581 (N_41581,N_41238,N_41020);
and U41582 (N_41582,N_41179,N_41472);
or U41583 (N_41583,N_41198,N_41108);
or U41584 (N_41584,N_41248,N_41209);
nor U41585 (N_41585,N_41117,N_41429);
or U41586 (N_41586,N_41386,N_41061);
xnor U41587 (N_41587,N_41413,N_41012);
nand U41588 (N_41588,N_41107,N_41225);
and U41589 (N_41589,N_41473,N_41138);
nor U41590 (N_41590,N_41214,N_41040);
nor U41591 (N_41591,N_41274,N_41316);
or U41592 (N_41592,N_41271,N_41339);
xnor U41593 (N_41593,N_41048,N_41445);
nor U41594 (N_41594,N_41221,N_41453);
and U41595 (N_41595,N_41130,N_41416);
and U41596 (N_41596,N_41059,N_41388);
nand U41597 (N_41597,N_41032,N_41295);
or U41598 (N_41598,N_41279,N_41203);
and U41599 (N_41599,N_41351,N_41224);
or U41600 (N_41600,N_41326,N_41257);
and U41601 (N_41601,N_41157,N_41097);
nand U41602 (N_41602,N_41410,N_41311);
and U41603 (N_41603,N_41437,N_41062);
xor U41604 (N_41604,N_41037,N_41273);
xor U41605 (N_41605,N_41120,N_41380);
or U41606 (N_41606,N_41202,N_41333);
or U41607 (N_41607,N_41423,N_41087);
nand U41608 (N_41608,N_41302,N_41229);
or U41609 (N_41609,N_41145,N_41174);
and U41610 (N_41610,N_41098,N_41475);
nor U41611 (N_41611,N_41487,N_41161);
nand U41612 (N_41612,N_41236,N_41047);
nor U41613 (N_41613,N_41239,N_41230);
nor U41614 (N_41614,N_41406,N_41099);
xnor U41615 (N_41615,N_41418,N_41456);
or U41616 (N_41616,N_41115,N_41485);
xnor U41617 (N_41617,N_41350,N_41315);
nand U41618 (N_41618,N_41476,N_41304);
nor U41619 (N_41619,N_41252,N_41359);
xor U41620 (N_41620,N_41139,N_41368);
and U41621 (N_41621,N_41414,N_41084);
xnor U41622 (N_41622,N_41355,N_41170);
nand U41623 (N_41623,N_41419,N_41289);
nor U41624 (N_41624,N_41089,N_41140);
and U41625 (N_41625,N_41197,N_41372);
or U41626 (N_41626,N_41440,N_41267);
or U41627 (N_41627,N_41454,N_41150);
and U41628 (N_41628,N_41085,N_41109);
xor U41629 (N_41629,N_41296,N_41266);
nand U41630 (N_41630,N_41322,N_41035);
nor U41631 (N_41631,N_41301,N_41024);
nand U41632 (N_41632,N_41395,N_41373);
or U41633 (N_41633,N_41480,N_41165);
and U41634 (N_41634,N_41126,N_41421);
nor U41635 (N_41635,N_41146,N_41114);
nor U41636 (N_41636,N_41030,N_41045);
xnor U41637 (N_41637,N_41183,N_41292);
nor U41638 (N_41638,N_41113,N_41181);
xnor U41639 (N_41639,N_41433,N_41129);
nor U41640 (N_41640,N_41193,N_41337);
nor U41641 (N_41641,N_41495,N_41381);
and U41642 (N_41642,N_41354,N_41390);
nand U41643 (N_41643,N_41320,N_41436);
xor U41644 (N_41644,N_41187,N_41028);
xor U41645 (N_41645,N_41200,N_41184);
nor U41646 (N_41646,N_41286,N_41389);
nand U41647 (N_41647,N_41094,N_41222);
and U41648 (N_41648,N_41442,N_41431);
and U41649 (N_41649,N_41291,N_41009);
xnor U41650 (N_41650,N_41379,N_41360);
or U41651 (N_41651,N_41343,N_41164);
xor U41652 (N_41652,N_41210,N_41082);
and U41653 (N_41653,N_41412,N_41443);
or U41654 (N_41654,N_41010,N_41444);
xnor U41655 (N_41655,N_41217,N_41223);
nor U41656 (N_41656,N_41134,N_41290);
xor U41657 (N_41657,N_41466,N_41357);
or U41658 (N_41658,N_41425,N_41090);
nand U41659 (N_41659,N_41306,N_41449);
xnor U41660 (N_41660,N_41323,N_41211);
nor U41661 (N_41661,N_41143,N_41349);
xor U41662 (N_41662,N_41072,N_41356);
nor U41663 (N_41663,N_41207,N_41385);
xnor U41664 (N_41664,N_41417,N_41031);
and U41665 (N_41665,N_41060,N_41483);
nand U41666 (N_41666,N_41213,N_41335);
xor U41667 (N_41667,N_41384,N_41428);
or U41668 (N_41668,N_41111,N_41321);
nor U41669 (N_41669,N_41195,N_41204);
xnor U41670 (N_41670,N_41231,N_41055);
or U41671 (N_41671,N_41155,N_41285);
or U41672 (N_41672,N_41064,N_41014);
or U41673 (N_41673,N_41439,N_41073);
or U41674 (N_41674,N_41358,N_41070);
and U41675 (N_41675,N_41079,N_41336);
xor U41676 (N_41676,N_41341,N_41141);
nor U41677 (N_41677,N_41121,N_41393);
nand U41678 (N_41678,N_41218,N_41068);
nor U41679 (N_41679,N_41237,N_41377);
or U41680 (N_41680,N_41234,N_41344);
nor U41681 (N_41681,N_41075,N_41261);
nor U41682 (N_41682,N_41127,N_41471);
xnor U41683 (N_41683,N_41411,N_41219);
nand U41684 (N_41684,N_41029,N_41101);
or U41685 (N_41685,N_41208,N_41352);
or U41686 (N_41686,N_41186,N_41233);
or U41687 (N_41687,N_41330,N_41201);
nor U41688 (N_41688,N_41076,N_41096);
nor U41689 (N_41689,N_41275,N_41367);
or U41690 (N_41690,N_41438,N_41118);
and U41691 (N_41691,N_41132,N_41294);
nor U41692 (N_41692,N_41370,N_41492);
or U41693 (N_41693,N_41249,N_41422);
nand U41694 (N_41694,N_41313,N_41100);
nand U41695 (N_41695,N_41494,N_41102);
nand U41696 (N_41696,N_41361,N_41398);
and U41697 (N_41697,N_41345,N_41278);
nor U41698 (N_41698,N_41149,N_41250);
nor U41699 (N_41699,N_41258,N_41022);
xor U41700 (N_41700,N_41242,N_41148);
xnor U41701 (N_41701,N_41092,N_41077);
nand U41702 (N_41702,N_41348,N_41287);
and U41703 (N_41703,N_41123,N_41432);
nand U41704 (N_41704,N_41133,N_41468);
nor U41705 (N_41705,N_41493,N_41426);
nand U41706 (N_41706,N_41057,N_41015);
xnor U41707 (N_41707,N_41297,N_41324);
nor U41708 (N_41708,N_41259,N_41106);
nand U41709 (N_41709,N_41374,N_41171);
xnor U41710 (N_41710,N_41499,N_41004);
nor U41711 (N_41711,N_41069,N_41452);
xor U41712 (N_41712,N_41112,N_41078);
and U41713 (N_41713,N_41154,N_41206);
xnor U41714 (N_41714,N_41011,N_41021);
nand U41715 (N_41715,N_41063,N_41043);
xnor U41716 (N_41716,N_41496,N_41104);
nand U41717 (N_41717,N_41163,N_41008);
nand U41718 (N_41718,N_41383,N_41441);
nand U41719 (N_41719,N_41407,N_41052);
nand U41720 (N_41720,N_41378,N_41054);
nor U41721 (N_41721,N_41392,N_41192);
nor U41722 (N_41722,N_41172,N_41016);
xor U41723 (N_41723,N_41185,N_41178);
and U41724 (N_41724,N_41310,N_41458);
xnor U41725 (N_41725,N_41482,N_41160);
nor U41726 (N_41726,N_41091,N_41488);
and U41727 (N_41727,N_41394,N_41158);
nand U41728 (N_41728,N_41175,N_41430);
and U41729 (N_41729,N_41334,N_41241);
nand U41730 (N_41730,N_41147,N_41255);
nor U41731 (N_41731,N_41065,N_41005);
nand U41732 (N_41732,N_41396,N_41169);
xor U41733 (N_41733,N_41196,N_41450);
and U41734 (N_41734,N_41465,N_41300);
or U41735 (N_41735,N_41447,N_41347);
or U41736 (N_41736,N_41376,N_41251);
and U41737 (N_41737,N_41124,N_41299);
and U41738 (N_41738,N_41125,N_41001);
xnor U41739 (N_41739,N_41227,N_41400);
nor U41740 (N_41740,N_41166,N_41346);
xor U41741 (N_41741,N_41479,N_41382);
or U41742 (N_41742,N_41036,N_41264);
nand U41743 (N_41743,N_41119,N_41455);
xor U41744 (N_41744,N_41403,N_41156);
nand U41745 (N_41745,N_41457,N_41007);
nor U41746 (N_41746,N_41095,N_41462);
xor U41747 (N_41747,N_41262,N_41497);
nand U41748 (N_41748,N_41276,N_41046);
and U41749 (N_41749,N_41318,N_41308);
nand U41750 (N_41750,N_41103,N_41196);
and U41751 (N_41751,N_41454,N_41011);
nor U41752 (N_41752,N_41189,N_41016);
nand U41753 (N_41753,N_41031,N_41270);
nand U41754 (N_41754,N_41014,N_41036);
nor U41755 (N_41755,N_41239,N_41402);
or U41756 (N_41756,N_41159,N_41296);
and U41757 (N_41757,N_41417,N_41218);
nor U41758 (N_41758,N_41333,N_41412);
and U41759 (N_41759,N_41033,N_41423);
nand U41760 (N_41760,N_41484,N_41193);
xor U41761 (N_41761,N_41290,N_41094);
xnor U41762 (N_41762,N_41232,N_41229);
or U41763 (N_41763,N_41168,N_41332);
or U41764 (N_41764,N_41227,N_41279);
nand U41765 (N_41765,N_41462,N_41111);
nor U41766 (N_41766,N_41498,N_41189);
xor U41767 (N_41767,N_41412,N_41330);
and U41768 (N_41768,N_41469,N_41025);
nand U41769 (N_41769,N_41011,N_41394);
nand U41770 (N_41770,N_41179,N_41104);
and U41771 (N_41771,N_41462,N_41156);
nor U41772 (N_41772,N_41142,N_41179);
nand U41773 (N_41773,N_41031,N_41402);
xnor U41774 (N_41774,N_41131,N_41055);
and U41775 (N_41775,N_41061,N_41400);
or U41776 (N_41776,N_41296,N_41280);
nand U41777 (N_41777,N_41482,N_41457);
and U41778 (N_41778,N_41307,N_41250);
or U41779 (N_41779,N_41480,N_41143);
nand U41780 (N_41780,N_41129,N_41011);
nor U41781 (N_41781,N_41281,N_41211);
and U41782 (N_41782,N_41382,N_41338);
or U41783 (N_41783,N_41095,N_41317);
or U41784 (N_41784,N_41092,N_41127);
or U41785 (N_41785,N_41092,N_41432);
nor U41786 (N_41786,N_41003,N_41173);
nor U41787 (N_41787,N_41017,N_41298);
and U41788 (N_41788,N_41057,N_41226);
and U41789 (N_41789,N_41064,N_41482);
xor U41790 (N_41790,N_41492,N_41423);
nor U41791 (N_41791,N_41090,N_41154);
nand U41792 (N_41792,N_41105,N_41244);
and U41793 (N_41793,N_41169,N_41103);
xor U41794 (N_41794,N_41241,N_41155);
and U41795 (N_41795,N_41450,N_41490);
or U41796 (N_41796,N_41392,N_41219);
or U41797 (N_41797,N_41311,N_41164);
xor U41798 (N_41798,N_41295,N_41072);
nand U41799 (N_41799,N_41018,N_41480);
or U41800 (N_41800,N_41100,N_41076);
nor U41801 (N_41801,N_41390,N_41243);
xor U41802 (N_41802,N_41105,N_41476);
xor U41803 (N_41803,N_41267,N_41364);
nand U41804 (N_41804,N_41223,N_41211);
xor U41805 (N_41805,N_41077,N_41367);
xor U41806 (N_41806,N_41142,N_41001);
nand U41807 (N_41807,N_41379,N_41000);
nand U41808 (N_41808,N_41416,N_41128);
xor U41809 (N_41809,N_41329,N_41418);
xor U41810 (N_41810,N_41458,N_41367);
or U41811 (N_41811,N_41487,N_41426);
or U41812 (N_41812,N_41132,N_41064);
or U41813 (N_41813,N_41454,N_41374);
xor U41814 (N_41814,N_41000,N_41019);
nor U41815 (N_41815,N_41065,N_41092);
or U41816 (N_41816,N_41408,N_41146);
or U41817 (N_41817,N_41464,N_41293);
nand U41818 (N_41818,N_41387,N_41131);
nor U41819 (N_41819,N_41421,N_41160);
and U41820 (N_41820,N_41048,N_41006);
xnor U41821 (N_41821,N_41471,N_41455);
nand U41822 (N_41822,N_41232,N_41106);
nand U41823 (N_41823,N_41282,N_41450);
nor U41824 (N_41824,N_41283,N_41058);
and U41825 (N_41825,N_41359,N_41001);
and U41826 (N_41826,N_41166,N_41018);
nor U41827 (N_41827,N_41107,N_41203);
and U41828 (N_41828,N_41220,N_41330);
xnor U41829 (N_41829,N_41358,N_41019);
nor U41830 (N_41830,N_41275,N_41004);
nor U41831 (N_41831,N_41395,N_41215);
nand U41832 (N_41832,N_41133,N_41476);
nor U41833 (N_41833,N_41113,N_41304);
xnor U41834 (N_41834,N_41295,N_41230);
nor U41835 (N_41835,N_41067,N_41086);
or U41836 (N_41836,N_41218,N_41376);
nand U41837 (N_41837,N_41183,N_41334);
and U41838 (N_41838,N_41045,N_41074);
nand U41839 (N_41839,N_41364,N_41142);
or U41840 (N_41840,N_41342,N_41022);
nand U41841 (N_41841,N_41016,N_41028);
xor U41842 (N_41842,N_41455,N_41002);
or U41843 (N_41843,N_41027,N_41145);
nor U41844 (N_41844,N_41036,N_41441);
xor U41845 (N_41845,N_41376,N_41014);
xor U41846 (N_41846,N_41287,N_41182);
nand U41847 (N_41847,N_41190,N_41228);
or U41848 (N_41848,N_41279,N_41239);
and U41849 (N_41849,N_41169,N_41010);
and U41850 (N_41850,N_41418,N_41446);
or U41851 (N_41851,N_41110,N_41317);
nand U41852 (N_41852,N_41236,N_41312);
and U41853 (N_41853,N_41445,N_41294);
xnor U41854 (N_41854,N_41491,N_41149);
nor U41855 (N_41855,N_41146,N_41086);
or U41856 (N_41856,N_41085,N_41051);
nor U41857 (N_41857,N_41155,N_41013);
nor U41858 (N_41858,N_41108,N_41171);
xor U41859 (N_41859,N_41315,N_41364);
or U41860 (N_41860,N_41348,N_41442);
nor U41861 (N_41861,N_41228,N_41249);
nor U41862 (N_41862,N_41111,N_41058);
or U41863 (N_41863,N_41131,N_41051);
xnor U41864 (N_41864,N_41246,N_41289);
nor U41865 (N_41865,N_41148,N_41109);
and U41866 (N_41866,N_41268,N_41309);
nor U41867 (N_41867,N_41297,N_41196);
xor U41868 (N_41868,N_41061,N_41299);
nand U41869 (N_41869,N_41396,N_41398);
or U41870 (N_41870,N_41260,N_41494);
nand U41871 (N_41871,N_41105,N_41047);
and U41872 (N_41872,N_41491,N_41255);
and U41873 (N_41873,N_41363,N_41027);
nand U41874 (N_41874,N_41477,N_41279);
and U41875 (N_41875,N_41395,N_41420);
or U41876 (N_41876,N_41109,N_41096);
or U41877 (N_41877,N_41173,N_41415);
nor U41878 (N_41878,N_41145,N_41436);
and U41879 (N_41879,N_41473,N_41319);
nand U41880 (N_41880,N_41427,N_41467);
xor U41881 (N_41881,N_41464,N_41062);
xnor U41882 (N_41882,N_41061,N_41290);
nand U41883 (N_41883,N_41323,N_41279);
nand U41884 (N_41884,N_41354,N_41025);
xor U41885 (N_41885,N_41101,N_41388);
nand U41886 (N_41886,N_41118,N_41237);
nand U41887 (N_41887,N_41187,N_41367);
and U41888 (N_41888,N_41398,N_41462);
or U41889 (N_41889,N_41073,N_41116);
nor U41890 (N_41890,N_41382,N_41150);
or U41891 (N_41891,N_41433,N_41078);
xnor U41892 (N_41892,N_41052,N_41473);
xor U41893 (N_41893,N_41469,N_41298);
and U41894 (N_41894,N_41320,N_41137);
nand U41895 (N_41895,N_41125,N_41452);
xor U41896 (N_41896,N_41124,N_41282);
nor U41897 (N_41897,N_41202,N_41301);
xnor U41898 (N_41898,N_41028,N_41463);
and U41899 (N_41899,N_41049,N_41331);
and U41900 (N_41900,N_41417,N_41439);
and U41901 (N_41901,N_41139,N_41042);
nor U41902 (N_41902,N_41178,N_41307);
nand U41903 (N_41903,N_41320,N_41118);
or U41904 (N_41904,N_41118,N_41075);
and U41905 (N_41905,N_41309,N_41033);
and U41906 (N_41906,N_41284,N_41037);
nor U41907 (N_41907,N_41221,N_41413);
nand U41908 (N_41908,N_41289,N_41151);
or U41909 (N_41909,N_41198,N_41351);
xnor U41910 (N_41910,N_41155,N_41438);
nor U41911 (N_41911,N_41186,N_41048);
xnor U41912 (N_41912,N_41477,N_41311);
xor U41913 (N_41913,N_41176,N_41358);
nand U41914 (N_41914,N_41439,N_41141);
nand U41915 (N_41915,N_41249,N_41499);
nand U41916 (N_41916,N_41328,N_41260);
and U41917 (N_41917,N_41272,N_41003);
nand U41918 (N_41918,N_41464,N_41262);
or U41919 (N_41919,N_41349,N_41043);
xor U41920 (N_41920,N_41091,N_41139);
nor U41921 (N_41921,N_41088,N_41320);
xor U41922 (N_41922,N_41218,N_41244);
nor U41923 (N_41923,N_41264,N_41260);
xnor U41924 (N_41924,N_41348,N_41450);
nand U41925 (N_41925,N_41472,N_41204);
nor U41926 (N_41926,N_41047,N_41475);
and U41927 (N_41927,N_41184,N_41185);
and U41928 (N_41928,N_41388,N_41335);
or U41929 (N_41929,N_41144,N_41103);
and U41930 (N_41930,N_41230,N_41479);
nand U41931 (N_41931,N_41204,N_41198);
xor U41932 (N_41932,N_41300,N_41095);
nor U41933 (N_41933,N_41147,N_41481);
or U41934 (N_41934,N_41474,N_41205);
xor U41935 (N_41935,N_41034,N_41116);
nor U41936 (N_41936,N_41433,N_41187);
nor U41937 (N_41937,N_41311,N_41067);
xnor U41938 (N_41938,N_41123,N_41190);
and U41939 (N_41939,N_41260,N_41279);
nand U41940 (N_41940,N_41000,N_41401);
and U41941 (N_41941,N_41427,N_41087);
and U41942 (N_41942,N_41215,N_41457);
or U41943 (N_41943,N_41349,N_41189);
nand U41944 (N_41944,N_41279,N_41137);
nor U41945 (N_41945,N_41001,N_41247);
xor U41946 (N_41946,N_41063,N_41371);
and U41947 (N_41947,N_41315,N_41125);
and U41948 (N_41948,N_41107,N_41492);
nor U41949 (N_41949,N_41491,N_41453);
nand U41950 (N_41950,N_41092,N_41316);
or U41951 (N_41951,N_41053,N_41143);
or U41952 (N_41952,N_41347,N_41124);
and U41953 (N_41953,N_41122,N_41031);
nand U41954 (N_41954,N_41436,N_41393);
nand U41955 (N_41955,N_41197,N_41402);
nand U41956 (N_41956,N_41173,N_41031);
nand U41957 (N_41957,N_41027,N_41477);
nor U41958 (N_41958,N_41259,N_41167);
nor U41959 (N_41959,N_41103,N_41391);
nor U41960 (N_41960,N_41252,N_41159);
nor U41961 (N_41961,N_41387,N_41487);
and U41962 (N_41962,N_41055,N_41470);
nand U41963 (N_41963,N_41074,N_41440);
and U41964 (N_41964,N_41366,N_41226);
and U41965 (N_41965,N_41147,N_41035);
nand U41966 (N_41966,N_41465,N_41469);
nand U41967 (N_41967,N_41101,N_41234);
and U41968 (N_41968,N_41246,N_41381);
and U41969 (N_41969,N_41131,N_41121);
nand U41970 (N_41970,N_41399,N_41214);
and U41971 (N_41971,N_41146,N_41369);
nand U41972 (N_41972,N_41318,N_41236);
nor U41973 (N_41973,N_41290,N_41040);
and U41974 (N_41974,N_41026,N_41259);
nand U41975 (N_41975,N_41129,N_41378);
nor U41976 (N_41976,N_41463,N_41063);
and U41977 (N_41977,N_41261,N_41010);
xnor U41978 (N_41978,N_41220,N_41192);
xnor U41979 (N_41979,N_41110,N_41434);
nand U41980 (N_41980,N_41057,N_41170);
xor U41981 (N_41981,N_41192,N_41421);
nor U41982 (N_41982,N_41232,N_41044);
nor U41983 (N_41983,N_41439,N_41393);
xor U41984 (N_41984,N_41073,N_41136);
and U41985 (N_41985,N_41497,N_41249);
or U41986 (N_41986,N_41132,N_41484);
and U41987 (N_41987,N_41397,N_41041);
or U41988 (N_41988,N_41225,N_41173);
and U41989 (N_41989,N_41132,N_41200);
nor U41990 (N_41990,N_41162,N_41331);
or U41991 (N_41991,N_41291,N_41228);
xnor U41992 (N_41992,N_41263,N_41380);
or U41993 (N_41993,N_41111,N_41241);
or U41994 (N_41994,N_41466,N_41413);
and U41995 (N_41995,N_41192,N_41497);
and U41996 (N_41996,N_41218,N_41389);
nor U41997 (N_41997,N_41411,N_41196);
or U41998 (N_41998,N_41319,N_41112);
nor U41999 (N_41999,N_41113,N_41231);
xnor U42000 (N_42000,N_41902,N_41667);
or U42001 (N_42001,N_41935,N_41837);
nand U42002 (N_42002,N_41887,N_41592);
or U42003 (N_42003,N_41764,N_41572);
xor U42004 (N_42004,N_41968,N_41873);
nand U42005 (N_42005,N_41882,N_41692);
nand U42006 (N_42006,N_41796,N_41773);
nand U42007 (N_42007,N_41980,N_41896);
nand U42008 (N_42008,N_41787,N_41869);
nand U42009 (N_42009,N_41766,N_41827);
xnor U42010 (N_42010,N_41566,N_41506);
xor U42011 (N_42011,N_41910,N_41969);
or U42012 (N_42012,N_41850,N_41853);
or U42013 (N_42013,N_41582,N_41772);
or U42014 (N_42014,N_41841,N_41816);
nor U42015 (N_42015,N_41697,N_41635);
and U42016 (N_42016,N_41878,N_41733);
nor U42017 (N_42017,N_41771,N_41618);
or U42018 (N_42018,N_41507,N_41580);
nand U42019 (N_42019,N_41683,N_41893);
or U42020 (N_42020,N_41921,N_41824);
nor U42021 (N_42021,N_41690,N_41938);
nor U42022 (N_42022,N_41604,N_41852);
or U42023 (N_42023,N_41602,N_41742);
and U42024 (N_42024,N_41728,N_41735);
nor U42025 (N_42025,N_41718,N_41805);
xor U42026 (N_42026,N_41704,N_41584);
nor U42027 (N_42027,N_41623,N_41989);
and U42028 (N_42028,N_41722,N_41577);
and U42029 (N_42029,N_41942,N_41847);
xnor U42030 (N_42030,N_41628,N_41711);
xnor U42031 (N_42031,N_41844,N_41621);
nor U42032 (N_42032,N_41633,N_41648);
xor U42033 (N_42033,N_41525,N_41851);
xor U42034 (N_42034,N_41906,N_41778);
nand U42035 (N_42035,N_41681,N_41738);
or U42036 (N_42036,N_41937,N_41620);
nor U42037 (N_42037,N_41732,N_41570);
xor U42038 (N_42038,N_41693,N_41658);
nand U42039 (N_42039,N_41710,N_41625);
xnor U42040 (N_42040,N_41515,N_41613);
nand U42041 (N_42041,N_41992,N_41561);
xnor U42042 (N_42042,N_41627,N_41855);
and U42043 (N_42043,N_41644,N_41894);
and U42044 (N_42044,N_41698,N_41668);
nand U42045 (N_42045,N_41811,N_41883);
and U42046 (N_42046,N_41736,N_41651);
or U42047 (N_42047,N_41678,N_41940);
xnor U42048 (N_42048,N_41836,N_41977);
or U42049 (N_42049,N_41931,N_41634);
xnor U42050 (N_42050,N_41933,N_41573);
and U42051 (N_42051,N_41813,N_41846);
and U42052 (N_42052,N_41567,N_41911);
or U42053 (N_42053,N_41675,N_41981);
nor U42054 (N_42054,N_41756,N_41591);
and U42055 (N_42055,N_41637,N_41821);
nand U42056 (N_42056,N_41661,N_41993);
and U42057 (N_42057,N_41952,N_41900);
nor U42058 (N_42058,N_41825,N_41598);
and U42059 (N_42059,N_41838,N_41550);
nand U42060 (N_42060,N_41551,N_41785);
nor U42061 (N_42061,N_41964,N_41588);
or U42062 (N_42062,N_41503,N_41652);
or U42063 (N_42063,N_41513,N_41715);
or U42064 (N_42064,N_41747,N_41723);
and U42065 (N_42065,N_41545,N_41810);
nor U42066 (N_42066,N_41769,N_41960);
or U42067 (N_42067,N_41533,N_41708);
nand U42068 (N_42068,N_41880,N_41903);
and U42069 (N_42069,N_41721,N_41786);
nand U42070 (N_42070,N_41996,N_41780);
or U42071 (N_42071,N_41973,N_41779);
and U42072 (N_42072,N_41749,N_41656);
or U42073 (N_42073,N_41532,N_41829);
nand U42074 (N_42074,N_41726,N_41700);
nor U42075 (N_42075,N_41674,N_41927);
nand U42076 (N_42076,N_41881,N_41544);
or U42077 (N_42077,N_41929,N_41632);
and U42078 (N_42078,N_41731,N_41783);
and U42079 (N_42079,N_41839,N_41765);
nor U42080 (N_42080,N_41502,N_41677);
or U42081 (N_42081,N_41543,N_41770);
xor U42082 (N_42082,N_41858,N_41801);
or U42083 (N_42083,N_41793,N_41535);
nor U42084 (N_42084,N_41870,N_41640);
or U42085 (N_42085,N_41707,N_41564);
or U42086 (N_42086,N_41919,N_41600);
nand U42087 (N_42087,N_41806,N_41777);
nand U42088 (N_42088,N_41516,N_41671);
nand U42089 (N_42089,N_41541,N_41596);
or U42090 (N_42090,N_41712,N_41754);
or U42091 (N_42091,N_41717,N_41967);
xnor U42092 (N_42092,N_41760,N_41868);
nand U42093 (N_42093,N_41581,N_41750);
xnor U42094 (N_42094,N_41945,N_41594);
and U42095 (N_42095,N_41616,N_41788);
nand U42096 (N_42096,N_41845,N_41916);
nand U42097 (N_42097,N_41886,N_41961);
and U42098 (N_42098,N_41554,N_41534);
nor U42099 (N_42099,N_41737,N_41687);
nor U42100 (N_42100,N_41505,N_41745);
nor U42101 (N_42101,N_41862,N_41832);
nand U42102 (N_42102,N_41646,N_41724);
xor U42103 (N_42103,N_41559,N_41939);
and U42104 (N_42104,N_41912,N_41642);
or U42105 (N_42105,N_41645,N_41579);
nor U42106 (N_42106,N_41528,N_41751);
nor U42107 (N_42107,N_41755,N_41905);
xor U42108 (N_42108,N_41848,N_41734);
and U42109 (N_42109,N_41930,N_41775);
or U42110 (N_42110,N_41975,N_41798);
and U42111 (N_42111,N_41574,N_41800);
and U42112 (N_42112,N_41514,N_41899);
nor U42113 (N_42113,N_41917,N_41521);
xor U42114 (N_42114,N_41762,N_41542);
or U42115 (N_42115,N_41818,N_41556);
and U42116 (N_42116,N_41639,N_41913);
nor U42117 (N_42117,N_41877,N_41888);
and U42118 (N_42118,N_41609,N_41955);
xor U42119 (N_42119,N_41739,N_41595);
nand U42120 (N_42120,N_41638,N_41915);
and U42121 (N_42121,N_41695,N_41617);
xnor U42122 (N_42122,N_41907,N_41624);
nor U42123 (N_42123,N_41918,N_41812);
nand U42124 (N_42124,N_41589,N_41746);
nor U42125 (N_42125,N_41974,N_41607);
and U42126 (N_42126,N_41953,N_41986);
xor U42127 (N_42127,N_41776,N_41970);
xnor U42128 (N_42128,N_41767,N_41630);
nor U42129 (N_42129,N_41565,N_41826);
nor U42130 (N_42130,N_41619,N_41696);
or U42131 (N_42131,N_41615,N_41703);
and U42132 (N_42132,N_41520,N_41730);
and U42133 (N_42133,N_41833,N_41797);
and U42134 (N_42134,N_41972,N_41979);
nor U42135 (N_42135,N_41804,N_41571);
or U42136 (N_42136,N_41553,N_41954);
and U42137 (N_42137,N_41744,N_41593);
or U42138 (N_42138,N_41748,N_41643);
nor U42139 (N_42139,N_41823,N_41814);
nor U42140 (N_42140,N_41784,N_41684);
or U42141 (N_42141,N_41947,N_41928);
nor U42142 (N_42142,N_41509,N_41702);
nand U42143 (N_42143,N_41665,N_41612);
and U42144 (N_42144,N_41508,N_41799);
or U42145 (N_42145,N_41990,N_41562);
nand U42146 (N_42146,N_41659,N_41966);
or U42147 (N_42147,N_41957,N_41861);
or U42148 (N_42148,N_41789,N_41555);
or U42149 (N_42149,N_41991,N_41922);
xnor U42150 (N_42150,N_41781,N_41995);
nor U42151 (N_42151,N_41547,N_41904);
and U42152 (N_42152,N_41672,N_41854);
nand U42153 (N_42153,N_41701,N_41971);
nor U42154 (N_42154,N_41699,N_41819);
nand U42155 (N_42155,N_41761,N_41891);
nand U42156 (N_42156,N_41629,N_41546);
xnor U42157 (N_42157,N_41705,N_41537);
xor U42158 (N_42158,N_41831,N_41792);
nand U42159 (N_42159,N_41669,N_41663);
nand U42160 (N_42160,N_41828,N_41808);
and U42161 (N_42161,N_41864,N_41994);
and U42162 (N_42162,N_41670,N_41531);
and U42163 (N_42163,N_41822,N_41501);
and U42164 (N_42164,N_41720,N_41817);
xor U42165 (N_42165,N_41587,N_41709);
nor U42166 (N_42166,N_41923,N_41976);
nand U42167 (N_42167,N_41653,N_41830);
xnor U42168 (N_42168,N_41840,N_41926);
xor U42169 (N_42169,N_41597,N_41714);
nand U42170 (N_42170,N_41518,N_41599);
or U42171 (N_42171,N_41522,N_41965);
xnor U42172 (N_42172,N_41803,N_41949);
and U42173 (N_42173,N_41606,N_41662);
and U42174 (N_42174,N_41897,N_41859);
nor U42175 (N_42175,N_41527,N_41835);
nor U42176 (N_42176,N_41890,N_41757);
nand U42177 (N_42177,N_41794,N_41641);
xnor U42178 (N_42178,N_41815,N_41622);
or U42179 (N_42179,N_41611,N_41568);
and U42180 (N_42180,N_41889,N_41583);
xor U42181 (N_42181,N_41863,N_41951);
and U42182 (N_42182,N_41743,N_41950);
xnor U42183 (N_42183,N_41530,N_41909);
nand U42184 (N_42184,N_41569,N_41809);
nand U42185 (N_42185,N_41948,N_41631);
nand U42186 (N_42186,N_41782,N_41586);
xor U42187 (N_42187,N_41872,N_41590);
nor U42188 (N_42188,N_41999,N_41932);
xor U42189 (N_42189,N_41680,N_41774);
xnor U42190 (N_42190,N_41657,N_41519);
xor U42191 (N_42191,N_41768,N_41512);
xor U42192 (N_42192,N_41614,N_41987);
nor U42193 (N_42193,N_41807,N_41925);
or U42194 (N_42194,N_41959,N_41795);
xor U42195 (N_42195,N_41759,N_41998);
and U42196 (N_42196,N_41849,N_41576);
nor U42197 (N_42197,N_41908,N_41552);
or U42198 (N_42198,N_41654,N_41956);
nand U42199 (N_42199,N_41536,N_41865);
or U42200 (N_42200,N_41884,N_41510);
nor U42201 (N_42201,N_41983,N_41962);
and U42202 (N_42202,N_41985,N_41941);
or U42203 (N_42203,N_41867,N_41603);
nor U42204 (N_42204,N_41540,N_41524);
xor U42205 (N_42205,N_41673,N_41946);
or U42206 (N_42206,N_41585,N_41791);
nand U42207 (N_42207,N_41688,N_41860);
nor U42208 (N_42208,N_41511,N_41558);
nand U42209 (N_42209,N_41504,N_41682);
nand U42210 (N_42210,N_41713,N_41575);
and U42211 (N_42211,N_41649,N_41626);
nand U42212 (N_42212,N_41605,N_41666);
and U42213 (N_42213,N_41834,N_41843);
or U42214 (N_42214,N_41752,N_41914);
and U42215 (N_42215,N_41790,N_41526);
and U42216 (N_42216,N_41538,N_41901);
nor U42217 (N_42217,N_41842,N_41539);
and U42218 (N_42218,N_41920,N_41601);
xnor U42219 (N_42219,N_41647,N_41885);
nor U42220 (N_42220,N_41660,N_41729);
xor U42221 (N_42221,N_41943,N_41958);
xor U42222 (N_42222,N_41753,N_41523);
nand U42223 (N_42223,N_41924,N_41997);
xnor U42224 (N_42224,N_41871,N_41716);
nor U42225 (N_42225,N_41875,N_41664);
or U42226 (N_42226,N_41934,N_41988);
nor U42227 (N_42227,N_41676,N_41500);
or U42228 (N_42228,N_41741,N_41610);
or U42229 (N_42229,N_41898,N_41719);
xor U42230 (N_42230,N_41820,N_41856);
nor U42231 (N_42231,N_41963,N_41879);
nand U42232 (N_42232,N_41944,N_41517);
or U42233 (N_42233,N_41694,N_41876);
or U42234 (N_42234,N_41655,N_41689);
nand U42235 (N_42235,N_41549,N_41548);
nand U42236 (N_42236,N_41557,N_41608);
or U42237 (N_42237,N_41802,N_41727);
nand U42238 (N_42238,N_41560,N_41740);
nor U42239 (N_42239,N_41763,N_41866);
nand U42240 (N_42240,N_41679,N_41895);
nand U42241 (N_42241,N_41691,N_41563);
nor U42242 (N_42242,N_41892,N_41706);
xnor U42243 (N_42243,N_41984,N_41758);
nor U42244 (N_42244,N_41529,N_41685);
and U42245 (N_42245,N_41578,N_41650);
and U42246 (N_42246,N_41686,N_41982);
or U42247 (N_42247,N_41874,N_41936);
or U42248 (N_42248,N_41725,N_41857);
and U42249 (N_42249,N_41978,N_41636);
nor U42250 (N_42250,N_41692,N_41601);
or U42251 (N_42251,N_41577,N_41895);
and U42252 (N_42252,N_41707,N_41757);
and U42253 (N_42253,N_41850,N_41667);
or U42254 (N_42254,N_41702,N_41811);
xnor U42255 (N_42255,N_41778,N_41869);
nand U42256 (N_42256,N_41667,N_41818);
nand U42257 (N_42257,N_41853,N_41710);
nand U42258 (N_42258,N_41632,N_41635);
xnor U42259 (N_42259,N_41674,N_41686);
nor U42260 (N_42260,N_41974,N_41588);
and U42261 (N_42261,N_41736,N_41592);
nand U42262 (N_42262,N_41786,N_41642);
nand U42263 (N_42263,N_41532,N_41867);
nor U42264 (N_42264,N_41649,N_41680);
or U42265 (N_42265,N_41721,N_41534);
nor U42266 (N_42266,N_41731,N_41979);
and U42267 (N_42267,N_41990,N_41952);
xor U42268 (N_42268,N_41527,N_41808);
and U42269 (N_42269,N_41565,N_41500);
or U42270 (N_42270,N_41918,N_41935);
xnor U42271 (N_42271,N_41939,N_41734);
xnor U42272 (N_42272,N_41641,N_41751);
xor U42273 (N_42273,N_41531,N_41722);
nand U42274 (N_42274,N_41780,N_41676);
nor U42275 (N_42275,N_41810,N_41893);
or U42276 (N_42276,N_41797,N_41673);
and U42277 (N_42277,N_41531,N_41816);
xnor U42278 (N_42278,N_41516,N_41843);
nor U42279 (N_42279,N_41894,N_41890);
or U42280 (N_42280,N_41835,N_41531);
nor U42281 (N_42281,N_41960,N_41651);
nand U42282 (N_42282,N_41660,N_41792);
and U42283 (N_42283,N_41545,N_41770);
and U42284 (N_42284,N_41918,N_41768);
nor U42285 (N_42285,N_41930,N_41789);
xor U42286 (N_42286,N_41859,N_41578);
nand U42287 (N_42287,N_41746,N_41678);
and U42288 (N_42288,N_41694,N_41680);
and U42289 (N_42289,N_41728,N_41795);
nand U42290 (N_42290,N_41513,N_41869);
nand U42291 (N_42291,N_41546,N_41668);
or U42292 (N_42292,N_41575,N_41895);
xor U42293 (N_42293,N_41676,N_41508);
xor U42294 (N_42294,N_41803,N_41712);
nand U42295 (N_42295,N_41540,N_41742);
or U42296 (N_42296,N_41683,N_41702);
nand U42297 (N_42297,N_41818,N_41679);
and U42298 (N_42298,N_41658,N_41769);
nor U42299 (N_42299,N_41703,N_41833);
and U42300 (N_42300,N_41810,N_41830);
nand U42301 (N_42301,N_41759,N_41975);
nor U42302 (N_42302,N_41893,N_41836);
or U42303 (N_42303,N_41616,N_41859);
nand U42304 (N_42304,N_41715,N_41635);
or U42305 (N_42305,N_41823,N_41794);
xor U42306 (N_42306,N_41726,N_41650);
nand U42307 (N_42307,N_41641,N_41894);
or U42308 (N_42308,N_41928,N_41962);
or U42309 (N_42309,N_41947,N_41751);
xnor U42310 (N_42310,N_41986,N_41888);
or U42311 (N_42311,N_41837,N_41687);
or U42312 (N_42312,N_41598,N_41823);
nand U42313 (N_42313,N_41616,N_41622);
nand U42314 (N_42314,N_41546,N_41567);
and U42315 (N_42315,N_41704,N_41777);
xor U42316 (N_42316,N_41819,N_41547);
xnor U42317 (N_42317,N_41918,N_41941);
xnor U42318 (N_42318,N_41854,N_41611);
and U42319 (N_42319,N_41592,N_41928);
nand U42320 (N_42320,N_41529,N_41999);
xnor U42321 (N_42321,N_41992,N_41774);
and U42322 (N_42322,N_41853,N_41892);
xnor U42323 (N_42323,N_41502,N_41897);
nor U42324 (N_42324,N_41598,N_41819);
nor U42325 (N_42325,N_41770,N_41785);
nor U42326 (N_42326,N_41598,N_41828);
or U42327 (N_42327,N_41779,N_41991);
or U42328 (N_42328,N_41965,N_41764);
and U42329 (N_42329,N_41702,N_41856);
and U42330 (N_42330,N_41590,N_41850);
xor U42331 (N_42331,N_41864,N_41819);
and U42332 (N_42332,N_41600,N_41955);
or U42333 (N_42333,N_41521,N_41620);
nand U42334 (N_42334,N_41668,N_41802);
or U42335 (N_42335,N_41878,N_41933);
nand U42336 (N_42336,N_41978,N_41564);
nor U42337 (N_42337,N_41652,N_41762);
or U42338 (N_42338,N_41861,N_41812);
nand U42339 (N_42339,N_41555,N_41502);
or U42340 (N_42340,N_41933,N_41554);
nor U42341 (N_42341,N_41959,N_41914);
nor U42342 (N_42342,N_41861,N_41984);
xor U42343 (N_42343,N_41952,N_41505);
and U42344 (N_42344,N_41969,N_41610);
xor U42345 (N_42345,N_41697,N_41699);
xor U42346 (N_42346,N_41598,N_41836);
nor U42347 (N_42347,N_41898,N_41763);
and U42348 (N_42348,N_41634,N_41637);
nor U42349 (N_42349,N_41805,N_41959);
or U42350 (N_42350,N_41513,N_41944);
and U42351 (N_42351,N_41742,N_41853);
nand U42352 (N_42352,N_41986,N_41581);
and U42353 (N_42353,N_41760,N_41535);
or U42354 (N_42354,N_41568,N_41896);
or U42355 (N_42355,N_41830,N_41896);
nor U42356 (N_42356,N_41501,N_41840);
or U42357 (N_42357,N_41775,N_41681);
nor U42358 (N_42358,N_41859,N_41839);
nor U42359 (N_42359,N_41637,N_41941);
or U42360 (N_42360,N_41889,N_41662);
nand U42361 (N_42361,N_41832,N_41835);
xnor U42362 (N_42362,N_41904,N_41530);
nor U42363 (N_42363,N_41568,N_41744);
and U42364 (N_42364,N_41666,N_41577);
or U42365 (N_42365,N_41922,N_41529);
nor U42366 (N_42366,N_41873,N_41900);
xor U42367 (N_42367,N_41885,N_41502);
or U42368 (N_42368,N_41961,N_41894);
xor U42369 (N_42369,N_41562,N_41768);
nand U42370 (N_42370,N_41903,N_41676);
nand U42371 (N_42371,N_41530,N_41660);
or U42372 (N_42372,N_41787,N_41747);
xor U42373 (N_42373,N_41614,N_41524);
nand U42374 (N_42374,N_41627,N_41764);
nand U42375 (N_42375,N_41905,N_41734);
xor U42376 (N_42376,N_41881,N_41909);
xor U42377 (N_42377,N_41821,N_41706);
nand U42378 (N_42378,N_41776,N_41608);
xor U42379 (N_42379,N_41885,N_41521);
nor U42380 (N_42380,N_41921,N_41761);
and U42381 (N_42381,N_41689,N_41676);
and U42382 (N_42382,N_41863,N_41938);
nand U42383 (N_42383,N_41587,N_41911);
xnor U42384 (N_42384,N_41640,N_41792);
and U42385 (N_42385,N_41895,N_41587);
nor U42386 (N_42386,N_41600,N_41751);
xnor U42387 (N_42387,N_41991,N_41517);
and U42388 (N_42388,N_41601,N_41607);
or U42389 (N_42389,N_41874,N_41778);
xor U42390 (N_42390,N_41814,N_41731);
nor U42391 (N_42391,N_41579,N_41699);
nor U42392 (N_42392,N_41683,N_41509);
xor U42393 (N_42393,N_41757,N_41581);
nand U42394 (N_42394,N_41633,N_41570);
or U42395 (N_42395,N_41797,N_41602);
and U42396 (N_42396,N_41928,N_41501);
or U42397 (N_42397,N_41937,N_41948);
or U42398 (N_42398,N_41524,N_41979);
and U42399 (N_42399,N_41868,N_41927);
nand U42400 (N_42400,N_41524,N_41520);
or U42401 (N_42401,N_41756,N_41822);
nand U42402 (N_42402,N_41960,N_41994);
nor U42403 (N_42403,N_41736,N_41683);
xnor U42404 (N_42404,N_41579,N_41756);
nand U42405 (N_42405,N_41814,N_41862);
and U42406 (N_42406,N_41854,N_41555);
xor U42407 (N_42407,N_41660,N_41970);
and U42408 (N_42408,N_41709,N_41704);
or U42409 (N_42409,N_41776,N_41543);
xor U42410 (N_42410,N_41917,N_41874);
xor U42411 (N_42411,N_41691,N_41931);
and U42412 (N_42412,N_41971,N_41696);
and U42413 (N_42413,N_41617,N_41961);
and U42414 (N_42414,N_41884,N_41899);
nor U42415 (N_42415,N_41696,N_41561);
or U42416 (N_42416,N_41897,N_41659);
or U42417 (N_42417,N_41853,N_41639);
nor U42418 (N_42418,N_41862,N_41555);
nor U42419 (N_42419,N_41891,N_41805);
and U42420 (N_42420,N_41920,N_41883);
or U42421 (N_42421,N_41821,N_41946);
nand U42422 (N_42422,N_41737,N_41896);
xnor U42423 (N_42423,N_41521,N_41817);
nand U42424 (N_42424,N_41935,N_41760);
and U42425 (N_42425,N_41610,N_41563);
or U42426 (N_42426,N_41831,N_41895);
and U42427 (N_42427,N_41896,N_41621);
nor U42428 (N_42428,N_41828,N_41933);
and U42429 (N_42429,N_41807,N_41575);
nand U42430 (N_42430,N_41925,N_41776);
xor U42431 (N_42431,N_41914,N_41861);
nor U42432 (N_42432,N_41832,N_41597);
xor U42433 (N_42433,N_41680,N_41505);
xnor U42434 (N_42434,N_41919,N_41669);
nand U42435 (N_42435,N_41999,N_41600);
and U42436 (N_42436,N_41618,N_41533);
and U42437 (N_42437,N_41892,N_41612);
or U42438 (N_42438,N_41861,N_41661);
xor U42439 (N_42439,N_41548,N_41755);
nand U42440 (N_42440,N_41503,N_41509);
or U42441 (N_42441,N_41889,N_41999);
xor U42442 (N_42442,N_41974,N_41844);
nor U42443 (N_42443,N_41903,N_41996);
xor U42444 (N_42444,N_41694,N_41890);
xnor U42445 (N_42445,N_41592,N_41560);
xor U42446 (N_42446,N_41594,N_41593);
nand U42447 (N_42447,N_41904,N_41572);
or U42448 (N_42448,N_41569,N_41672);
or U42449 (N_42449,N_41568,N_41713);
and U42450 (N_42450,N_41652,N_41845);
and U42451 (N_42451,N_41535,N_41927);
and U42452 (N_42452,N_41895,N_41746);
xnor U42453 (N_42453,N_41904,N_41593);
and U42454 (N_42454,N_41613,N_41606);
xnor U42455 (N_42455,N_41622,N_41741);
xor U42456 (N_42456,N_41686,N_41768);
nor U42457 (N_42457,N_41948,N_41879);
xor U42458 (N_42458,N_41601,N_41664);
and U42459 (N_42459,N_41710,N_41551);
nand U42460 (N_42460,N_41609,N_41536);
xnor U42461 (N_42461,N_41813,N_41777);
and U42462 (N_42462,N_41834,N_41777);
and U42463 (N_42463,N_41760,N_41871);
or U42464 (N_42464,N_41999,N_41505);
nor U42465 (N_42465,N_41747,N_41773);
nand U42466 (N_42466,N_41619,N_41585);
nand U42467 (N_42467,N_41846,N_41530);
or U42468 (N_42468,N_41790,N_41981);
nor U42469 (N_42469,N_41707,N_41761);
or U42470 (N_42470,N_41784,N_41661);
xor U42471 (N_42471,N_41749,N_41960);
or U42472 (N_42472,N_41840,N_41532);
nor U42473 (N_42473,N_41635,N_41831);
xor U42474 (N_42474,N_41769,N_41844);
nand U42475 (N_42475,N_41933,N_41612);
nand U42476 (N_42476,N_41528,N_41646);
nor U42477 (N_42477,N_41899,N_41905);
nand U42478 (N_42478,N_41759,N_41764);
or U42479 (N_42479,N_41951,N_41583);
nand U42480 (N_42480,N_41520,N_41630);
nand U42481 (N_42481,N_41934,N_41672);
or U42482 (N_42482,N_41812,N_41957);
nor U42483 (N_42483,N_41887,N_41663);
or U42484 (N_42484,N_41776,N_41524);
xor U42485 (N_42485,N_41517,N_41516);
or U42486 (N_42486,N_41618,N_41839);
nor U42487 (N_42487,N_41924,N_41777);
xor U42488 (N_42488,N_41908,N_41935);
xor U42489 (N_42489,N_41695,N_41984);
and U42490 (N_42490,N_41677,N_41596);
nor U42491 (N_42491,N_41532,N_41528);
or U42492 (N_42492,N_41634,N_41705);
nand U42493 (N_42493,N_41689,N_41808);
nor U42494 (N_42494,N_41813,N_41863);
and U42495 (N_42495,N_41818,N_41938);
nand U42496 (N_42496,N_41525,N_41766);
or U42497 (N_42497,N_41983,N_41688);
nand U42498 (N_42498,N_41800,N_41631);
nand U42499 (N_42499,N_41846,N_41601);
or U42500 (N_42500,N_42335,N_42273);
or U42501 (N_42501,N_42050,N_42474);
nand U42502 (N_42502,N_42207,N_42060);
xor U42503 (N_42503,N_42321,N_42336);
nor U42504 (N_42504,N_42268,N_42077);
or U42505 (N_42505,N_42159,N_42492);
or U42506 (N_42506,N_42397,N_42279);
nand U42507 (N_42507,N_42491,N_42055);
and U42508 (N_42508,N_42252,N_42197);
or U42509 (N_42509,N_42436,N_42066);
or U42510 (N_42510,N_42497,N_42091);
nor U42511 (N_42511,N_42437,N_42391);
and U42512 (N_42512,N_42194,N_42428);
or U42513 (N_42513,N_42212,N_42153);
and U42514 (N_42514,N_42134,N_42456);
nor U42515 (N_42515,N_42215,N_42367);
and U42516 (N_42516,N_42243,N_42364);
and U42517 (N_42517,N_42465,N_42124);
nand U42518 (N_42518,N_42267,N_42018);
nand U42519 (N_42519,N_42021,N_42407);
nor U42520 (N_42520,N_42216,N_42111);
nor U42521 (N_42521,N_42461,N_42410);
or U42522 (N_42522,N_42355,N_42334);
or U42523 (N_42523,N_42486,N_42366);
nand U42524 (N_42524,N_42001,N_42265);
or U42525 (N_42525,N_42317,N_42405);
xor U42526 (N_42526,N_42094,N_42020);
and U42527 (N_42527,N_42189,N_42012);
or U42528 (N_42528,N_42261,N_42024);
nor U42529 (N_42529,N_42343,N_42220);
or U42530 (N_42530,N_42179,N_42183);
or U42531 (N_42531,N_42193,N_42223);
nor U42532 (N_42532,N_42118,N_42123);
or U42533 (N_42533,N_42435,N_42235);
and U42534 (N_42534,N_42203,N_42376);
nand U42535 (N_42535,N_42283,N_42447);
xor U42536 (N_42536,N_42038,N_42108);
xnor U42537 (N_42537,N_42096,N_42196);
nand U42538 (N_42538,N_42146,N_42044);
nor U42539 (N_42539,N_42051,N_42419);
nor U42540 (N_42540,N_42314,N_42454);
and U42541 (N_42541,N_42385,N_42290);
xnor U42542 (N_42542,N_42382,N_42301);
or U42543 (N_42543,N_42357,N_42065);
and U42544 (N_42544,N_42082,N_42042);
or U42545 (N_42545,N_42286,N_42272);
xnor U42546 (N_42546,N_42092,N_42316);
or U42547 (N_42547,N_42054,N_42069);
nand U42548 (N_42548,N_42190,N_42387);
xnor U42549 (N_42549,N_42141,N_42485);
and U42550 (N_42550,N_42247,N_42169);
nor U42551 (N_42551,N_42182,N_42351);
nor U42552 (N_42552,N_42043,N_42450);
xnor U42553 (N_42553,N_42112,N_42140);
xnor U42554 (N_42554,N_42409,N_42186);
and U42555 (N_42555,N_42295,N_42093);
nor U42556 (N_42556,N_42389,N_42148);
nor U42557 (N_42557,N_42284,N_42289);
nand U42558 (N_42558,N_42151,N_42156);
nor U42559 (N_42559,N_42218,N_42211);
nand U42560 (N_42560,N_42347,N_42463);
nand U42561 (N_42561,N_42188,N_42328);
and U42562 (N_42562,N_42341,N_42256);
xnor U42563 (N_42563,N_42324,N_42332);
nand U42564 (N_42564,N_42368,N_42070);
xor U42565 (N_42565,N_42128,N_42327);
nand U42566 (N_42566,N_42274,N_42199);
and U42567 (N_42567,N_42184,N_42131);
nand U42568 (N_42568,N_42348,N_42445);
and U42569 (N_42569,N_42308,N_42342);
xnor U42570 (N_42570,N_42312,N_42344);
nor U42571 (N_42571,N_42126,N_42296);
nand U42572 (N_42572,N_42424,N_42072);
xor U42573 (N_42573,N_42291,N_42408);
xor U42574 (N_42574,N_42191,N_42358);
nor U42575 (N_42575,N_42361,N_42469);
and U42576 (N_42576,N_42144,N_42488);
nor U42577 (N_42577,N_42175,N_42318);
nand U42578 (N_42578,N_42278,N_42299);
and U42579 (N_42579,N_42076,N_42281);
xor U42580 (N_42580,N_42306,N_42227);
nand U42581 (N_42581,N_42418,N_42239);
and U42582 (N_42582,N_42395,N_42310);
nand U42583 (N_42583,N_42476,N_42384);
and U42584 (N_42584,N_42237,N_42198);
nand U42585 (N_42585,N_42172,N_42241);
xnor U42586 (N_42586,N_42149,N_42285);
nor U42587 (N_42587,N_42443,N_42046);
xnor U42588 (N_42588,N_42319,N_42019);
xnor U42589 (N_42589,N_42249,N_42116);
or U42590 (N_42590,N_42154,N_42269);
xor U42591 (N_42591,N_42225,N_42244);
nand U42592 (N_42592,N_42023,N_42416);
or U42593 (N_42593,N_42171,N_42362);
xor U42594 (N_42594,N_42214,N_42113);
xor U42595 (N_42595,N_42400,N_42333);
or U42596 (N_42596,N_42311,N_42037);
nor U42597 (N_42597,N_42471,N_42170);
xor U42598 (N_42598,N_42147,N_42005);
or U42599 (N_42599,N_42487,N_42457);
xnor U42600 (N_42600,N_42423,N_42490);
xor U42601 (N_42601,N_42266,N_42090);
xnor U42602 (N_42602,N_42117,N_42204);
or U42603 (N_42603,N_42130,N_42099);
or U42604 (N_42604,N_42138,N_42426);
and U42605 (N_42605,N_42380,N_42036);
nand U42606 (N_42606,N_42280,N_42132);
or U42607 (N_42607,N_42015,N_42152);
and U42608 (N_42608,N_42217,N_42142);
xor U42609 (N_42609,N_42122,N_42434);
xor U42610 (N_42610,N_42399,N_42462);
xor U42611 (N_42611,N_42392,N_42228);
xor U42612 (N_42612,N_42078,N_42467);
and U42613 (N_42613,N_42420,N_42262);
nor U42614 (N_42614,N_42004,N_42449);
nand U42615 (N_42615,N_42232,N_42006);
nor U42616 (N_42616,N_42475,N_42466);
xor U42617 (N_42617,N_42103,N_42010);
nor U42618 (N_42618,N_42071,N_42095);
xor U42619 (N_42619,N_42390,N_42430);
or U42620 (N_42620,N_42255,N_42346);
xor U42621 (N_42621,N_42181,N_42323);
and U42622 (N_42622,N_42429,N_42287);
and U42623 (N_42623,N_42480,N_42097);
nand U42624 (N_42624,N_42119,N_42174);
and U42625 (N_42625,N_42254,N_42164);
or U42626 (N_42626,N_42242,N_42002);
and U42627 (N_42627,N_42478,N_42378);
xor U42628 (N_42628,N_42340,N_42027);
and U42629 (N_42629,N_42468,N_42026);
or U42630 (N_42630,N_42477,N_42143);
xnor U42631 (N_42631,N_42448,N_42135);
xnor U42632 (N_42632,N_42370,N_42201);
or U42633 (N_42633,N_42068,N_42352);
and U42634 (N_42634,N_42114,N_42438);
xnor U42635 (N_42635,N_42115,N_42464);
or U42636 (N_42636,N_42326,N_42062);
or U42637 (N_42637,N_42451,N_42209);
or U42638 (N_42638,N_42303,N_42022);
and U42639 (N_42639,N_42157,N_42298);
xnor U42640 (N_42640,N_42246,N_42176);
nor U42641 (N_42641,N_42275,N_42109);
or U42642 (N_42642,N_42433,N_42297);
nand U42643 (N_42643,N_42016,N_42185);
nand U42644 (N_42644,N_42425,N_42411);
or U42645 (N_42645,N_42263,N_42374);
nand U42646 (N_42646,N_42360,N_42472);
nand U42647 (N_42647,N_42208,N_42479);
and U42648 (N_42648,N_42402,N_42059);
xor U42649 (N_42649,N_42330,N_42041);
xnor U42650 (N_42650,N_42003,N_42393);
xnor U42651 (N_42651,N_42377,N_42253);
and U42652 (N_42652,N_42105,N_42056);
and U42653 (N_42653,N_42270,N_42089);
nand U42654 (N_42654,N_42388,N_42431);
xnor U42655 (N_42655,N_42187,N_42257);
and U42656 (N_42656,N_42180,N_42013);
nand U42657 (N_42657,N_42213,N_42309);
nor U42658 (N_42658,N_42271,N_42064);
or U42659 (N_42659,N_42133,N_42313);
or U42660 (N_42660,N_42231,N_42383);
or U42661 (N_42661,N_42300,N_42083);
nor U42662 (N_42662,N_42224,N_42258);
nand U42663 (N_42663,N_42173,N_42205);
xnor U42664 (N_42664,N_42292,N_42085);
nand U42665 (N_42665,N_42259,N_42039);
nand U42666 (N_42666,N_42030,N_42444);
nand U42667 (N_42667,N_42277,N_42079);
or U42668 (N_42668,N_42222,N_42167);
nand U42669 (N_42669,N_42088,N_42127);
nor U42670 (N_42670,N_42011,N_42034);
or U42671 (N_42671,N_42017,N_42315);
and U42672 (N_42672,N_42081,N_42087);
or U42673 (N_42673,N_42009,N_42307);
xnor U42674 (N_42674,N_42061,N_42048);
or U42675 (N_42675,N_42162,N_42337);
nand U42676 (N_42676,N_42052,N_42210);
nor U42677 (N_42677,N_42233,N_42339);
and U42678 (N_42678,N_42221,N_42356);
and U42679 (N_42679,N_42359,N_42440);
xnor U42680 (N_42680,N_42226,N_42481);
and U42681 (N_42681,N_42106,N_42245);
nor U42682 (N_42682,N_42029,N_42107);
and U42683 (N_42683,N_42294,N_42129);
and U42684 (N_42684,N_42484,N_42058);
or U42685 (N_42685,N_42495,N_42000);
or U42686 (N_42686,N_42483,N_42282);
and U42687 (N_42687,N_42033,N_42040);
xor U42688 (N_42688,N_42100,N_42349);
xor U42689 (N_42689,N_42240,N_42086);
xor U42690 (N_42690,N_42442,N_42473);
nor U42691 (N_42691,N_42178,N_42379);
nand U42692 (N_42692,N_42372,N_42369);
nand U42693 (N_42693,N_42104,N_42206);
nor U42694 (N_42694,N_42136,N_42238);
xor U42695 (N_42695,N_42120,N_42414);
nand U42696 (N_42696,N_42489,N_42073);
nand U42697 (N_42697,N_42412,N_42394);
nand U42698 (N_42698,N_42439,N_42053);
or U42699 (N_42699,N_42350,N_42381);
nor U42700 (N_42700,N_42032,N_42145);
xor U42701 (N_42701,N_42168,N_42063);
and U42702 (N_42702,N_42406,N_42421);
or U42703 (N_42703,N_42080,N_42028);
nand U42704 (N_42704,N_42322,N_42453);
or U42705 (N_42705,N_42452,N_42125);
nor U42706 (N_42706,N_42417,N_42415);
nand U42707 (N_42707,N_42413,N_42177);
xnor U42708 (N_42708,N_42320,N_42101);
or U42709 (N_42709,N_42251,N_42499);
xnor U42710 (N_42710,N_42338,N_42371);
and U42711 (N_42711,N_42396,N_42007);
and U42712 (N_42712,N_42161,N_42098);
and U42713 (N_42713,N_42345,N_42398);
and U42714 (N_42714,N_42446,N_42493);
or U42715 (N_42715,N_42137,N_42498);
and U42716 (N_42716,N_42363,N_42219);
and U42717 (N_42717,N_42288,N_42200);
xnor U42718 (N_42718,N_42496,N_42160);
nand U42719 (N_42719,N_42084,N_42494);
nand U42720 (N_42720,N_42401,N_42195);
and U42721 (N_42721,N_42158,N_42404);
xnor U42722 (N_42722,N_42427,N_42234);
or U42723 (N_42723,N_42166,N_42365);
or U42724 (N_42724,N_42403,N_42260);
and U42725 (N_42725,N_42264,N_42459);
nand U42726 (N_42726,N_42470,N_42075);
and U42727 (N_42727,N_42458,N_42230);
xnor U42728 (N_42728,N_42250,N_42293);
nand U42729 (N_42729,N_42305,N_42304);
xor U42730 (N_42730,N_42014,N_42202);
or U42731 (N_42731,N_42067,N_42248);
nor U42732 (N_42732,N_42155,N_42008);
nand U42733 (N_42733,N_42165,N_42025);
or U42734 (N_42734,N_42331,N_42139);
and U42735 (N_42735,N_42110,N_42031);
nor U42736 (N_42736,N_42432,N_42163);
nand U42737 (N_42737,N_42192,N_42121);
and U42738 (N_42738,N_42386,N_42236);
or U42739 (N_42739,N_42325,N_42102);
xnor U42740 (N_42740,N_42302,N_42229);
or U42741 (N_42741,N_42049,N_42057);
and U42742 (N_42742,N_42460,N_42329);
nor U42743 (N_42743,N_42353,N_42354);
nand U42744 (N_42744,N_42045,N_42276);
xnor U42745 (N_42745,N_42455,N_42035);
xnor U42746 (N_42746,N_42482,N_42074);
nand U42747 (N_42747,N_42441,N_42422);
xor U42748 (N_42748,N_42375,N_42047);
nor U42749 (N_42749,N_42373,N_42150);
xor U42750 (N_42750,N_42169,N_42287);
and U42751 (N_42751,N_42422,N_42015);
or U42752 (N_42752,N_42071,N_42160);
and U42753 (N_42753,N_42465,N_42299);
or U42754 (N_42754,N_42079,N_42037);
and U42755 (N_42755,N_42367,N_42214);
nand U42756 (N_42756,N_42090,N_42057);
and U42757 (N_42757,N_42456,N_42434);
xor U42758 (N_42758,N_42023,N_42336);
or U42759 (N_42759,N_42028,N_42434);
nor U42760 (N_42760,N_42063,N_42396);
and U42761 (N_42761,N_42445,N_42049);
xnor U42762 (N_42762,N_42223,N_42179);
xnor U42763 (N_42763,N_42269,N_42202);
nor U42764 (N_42764,N_42088,N_42315);
xor U42765 (N_42765,N_42396,N_42142);
xor U42766 (N_42766,N_42143,N_42214);
xor U42767 (N_42767,N_42210,N_42108);
xnor U42768 (N_42768,N_42484,N_42016);
and U42769 (N_42769,N_42058,N_42409);
and U42770 (N_42770,N_42455,N_42114);
nand U42771 (N_42771,N_42449,N_42304);
nor U42772 (N_42772,N_42088,N_42312);
xnor U42773 (N_42773,N_42330,N_42281);
or U42774 (N_42774,N_42383,N_42395);
and U42775 (N_42775,N_42355,N_42262);
or U42776 (N_42776,N_42107,N_42405);
xnor U42777 (N_42777,N_42175,N_42237);
nand U42778 (N_42778,N_42177,N_42143);
nor U42779 (N_42779,N_42179,N_42082);
nor U42780 (N_42780,N_42416,N_42205);
xor U42781 (N_42781,N_42479,N_42321);
nor U42782 (N_42782,N_42403,N_42405);
nor U42783 (N_42783,N_42019,N_42477);
nand U42784 (N_42784,N_42263,N_42470);
or U42785 (N_42785,N_42342,N_42347);
xor U42786 (N_42786,N_42110,N_42080);
or U42787 (N_42787,N_42315,N_42394);
or U42788 (N_42788,N_42302,N_42403);
and U42789 (N_42789,N_42215,N_42278);
and U42790 (N_42790,N_42271,N_42241);
nand U42791 (N_42791,N_42031,N_42122);
nand U42792 (N_42792,N_42284,N_42247);
or U42793 (N_42793,N_42475,N_42457);
or U42794 (N_42794,N_42124,N_42393);
xnor U42795 (N_42795,N_42055,N_42444);
xnor U42796 (N_42796,N_42322,N_42056);
and U42797 (N_42797,N_42240,N_42426);
xnor U42798 (N_42798,N_42470,N_42419);
or U42799 (N_42799,N_42305,N_42417);
xor U42800 (N_42800,N_42497,N_42376);
or U42801 (N_42801,N_42100,N_42483);
nor U42802 (N_42802,N_42409,N_42092);
xnor U42803 (N_42803,N_42113,N_42016);
and U42804 (N_42804,N_42340,N_42143);
xor U42805 (N_42805,N_42165,N_42098);
xor U42806 (N_42806,N_42069,N_42056);
xnor U42807 (N_42807,N_42074,N_42386);
or U42808 (N_42808,N_42451,N_42164);
and U42809 (N_42809,N_42229,N_42128);
nor U42810 (N_42810,N_42204,N_42072);
or U42811 (N_42811,N_42003,N_42464);
or U42812 (N_42812,N_42110,N_42273);
or U42813 (N_42813,N_42443,N_42442);
nand U42814 (N_42814,N_42029,N_42068);
or U42815 (N_42815,N_42064,N_42220);
and U42816 (N_42816,N_42405,N_42369);
or U42817 (N_42817,N_42052,N_42265);
and U42818 (N_42818,N_42214,N_42431);
and U42819 (N_42819,N_42377,N_42272);
and U42820 (N_42820,N_42231,N_42485);
nand U42821 (N_42821,N_42370,N_42498);
and U42822 (N_42822,N_42280,N_42165);
or U42823 (N_42823,N_42488,N_42395);
and U42824 (N_42824,N_42166,N_42470);
nand U42825 (N_42825,N_42404,N_42213);
and U42826 (N_42826,N_42495,N_42319);
nand U42827 (N_42827,N_42449,N_42392);
nor U42828 (N_42828,N_42170,N_42122);
and U42829 (N_42829,N_42106,N_42194);
nor U42830 (N_42830,N_42023,N_42225);
nor U42831 (N_42831,N_42135,N_42477);
or U42832 (N_42832,N_42156,N_42274);
or U42833 (N_42833,N_42367,N_42306);
nand U42834 (N_42834,N_42181,N_42207);
nand U42835 (N_42835,N_42001,N_42100);
nor U42836 (N_42836,N_42213,N_42091);
xor U42837 (N_42837,N_42238,N_42291);
or U42838 (N_42838,N_42162,N_42132);
xor U42839 (N_42839,N_42290,N_42412);
and U42840 (N_42840,N_42336,N_42366);
nand U42841 (N_42841,N_42470,N_42151);
nand U42842 (N_42842,N_42302,N_42072);
nand U42843 (N_42843,N_42123,N_42248);
nor U42844 (N_42844,N_42411,N_42112);
nand U42845 (N_42845,N_42259,N_42136);
and U42846 (N_42846,N_42135,N_42155);
xnor U42847 (N_42847,N_42416,N_42095);
and U42848 (N_42848,N_42104,N_42196);
nor U42849 (N_42849,N_42001,N_42344);
nor U42850 (N_42850,N_42236,N_42382);
nand U42851 (N_42851,N_42180,N_42070);
nor U42852 (N_42852,N_42051,N_42191);
nor U42853 (N_42853,N_42286,N_42328);
nand U42854 (N_42854,N_42286,N_42176);
and U42855 (N_42855,N_42359,N_42018);
nor U42856 (N_42856,N_42453,N_42244);
xor U42857 (N_42857,N_42098,N_42010);
nor U42858 (N_42858,N_42178,N_42043);
or U42859 (N_42859,N_42094,N_42310);
and U42860 (N_42860,N_42142,N_42352);
or U42861 (N_42861,N_42351,N_42384);
nor U42862 (N_42862,N_42246,N_42433);
nor U42863 (N_42863,N_42426,N_42324);
and U42864 (N_42864,N_42229,N_42210);
or U42865 (N_42865,N_42491,N_42028);
or U42866 (N_42866,N_42137,N_42067);
and U42867 (N_42867,N_42236,N_42033);
and U42868 (N_42868,N_42082,N_42364);
and U42869 (N_42869,N_42237,N_42358);
nand U42870 (N_42870,N_42471,N_42075);
or U42871 (N_42871,N_42356,N_42403);
xor U42872 (N_42872,N_42306,N_42475);
nand U42873 (N_42873,N_42400,N_42184);
xor U42874 (N_42874,N_42010,N_42160);
and U42875 (N_42875,N_42495,N_42316);
or U42876 (N_42876,N_42077,N_42207);
and U42877 (N_42877,N_42422,N_42198);
nand U42878 (N_42878,N_42258,N_42018);
nor U42879 (N_42879,N_42228,N_42329);
or U42880 (N_42880,N_42426,N_42232);
and U42881 (N_42881,N_42214,N_42362);
and U42882 (N_42882,N_42018,N_42466);
nand U42883 (N_42883,N_42257,N_42380);
and U42884 (N_42884,N_42393,N_42466);
nand U42885 (N_42885,N_42226,N_42066);
or U42886 (N_42886,N_42265,N_42475);
or U42887 (N_42887,N_42148,N_42488);
xnor U42888 (N_42888,N_42197,N_42402);
nand U42889 (N_42889,N_42265,N_42425);
xnor U42890 (N_42890,N_42471,N_42439);
or U42891 (N_42891,N_42166,N_42443);
nand U42892 (N_42892,N_42174,N_42279);
nand U42893 (N_42893,N_42384,N_42083);
xor U42894 (N_42894,N_42246,N_42069);
or U42895 (N_42895,N_42273,N_42417);
and U42896 (N_42896,N_42351,N_42342);
or U42897 (N_42897,N_42016,N_42099);
xor U42898 (N_42898,N_42365,N_42218);
or U42899 (N_42899,N_42059,N_42223);
nor U42900 (N_42900,N_42272,N_42175);
nand U42901 (N_42901,N_42001,N_42162);
nand U42902 (N_42902,N_42286,N_42081);
nand U42903 (N_42903,N_42482,N_42456);
xnor U42904 (N_42904,N_42234,N_42111);
nand U42905 (N_42905,N_42079,N_42386);
or U42906 (N_42906,N_42123,N_42247);
and U42907 (N_42907,N_42335,N_42400);
and U42908 (N_42908,N_42339,N_42426);
or U42909 (N_42909,N_42437,N_42027);
nor U42910 (N_42910,N_42119,N_42264);
nor U42911 (N_42911,N_42335,N_42448);
nand U42912 (N_42912,N_42053,N_42006);
or U42913 (N_42913,N_42306,N_42485);
xor U42914 (N_42914,N_42040,N_42260);
nor U42915 (N_42915,N_42394,N_42265);
or U42916 (N_42916,N_42357,N_42426);
and U42917 (N_42917,N_42278,N_42018);
nor U42918 (N_42918,N_42134,N_42124);
and U42919 (N_42919,N_42426,N_42137);
and U42920 (N_42920,N_42388,N_42232);
or U42921 (N_42921,N_42274,N_42000);
or U42922 (N_42922,N_42425,N_42476);
nand U42923 (N_42923,N_42066,N_42408);
and U42924 (N_42924,N_42318,N_42262);
xor U42925 (N_42925,N_42062,N_42179);
nand U42926 (N_42926,N_42309,N_42402);
or U42927 (N_42927,N_42052,N_42322);
or U42928 (N_42928,N_42155,N_42124);
nand U42929 (N_42929,N_42044,N_42412);
nor U42930 (N_42930,N_42114,N_42150);
and U42931 (N_42931,N_42263,N_42208);
nor U42932 (N_42932,N_42215,N_42042);
nor U42933 (N_42933,N_42221,N_42247);
nand U42934 (N_42934,N_42120,N_42278);
and U42935 (N_42935,N_42291,N_42329);
xor U42936 (N_42936,N_42300,N_42350);
and U42937 (N_42937,N_42305,N_42166);
or U42938 (N_42938,N_42283,N_42478);
xnor U42939 (N_42939,N_42041,N_42316);
and U42940 (N_42940,N_42316,N_42044);
and U42941 (N_42941,N_42023,N_42205);
nand U42942 (N_42942,N_42369,N_42222);
and U42943 (N_42943,N_42358,N_42440);
and U42944 (N_42944,N_42328,N_42092);
nor U42945 (N_42945,N_42494,N_42160);
nand U42946 (N_42946,N_42000,N_42117);
nand U42947 (N_42947,N_42427,N_42315);
xnor U42948 (N_42948,N_42366,N_42191);
xor U42949 (N_42949,N_42134,N_42172);
xnor U42950 (N_42950,N_42397,N_42093);
nor U42951 (N_42951,N_42050,N_42489);
nand U42952 (N_42952,N_42475,N_42209);
nand U42953 (N_42953,N_42159,N_42316);
and U42954 (N_42954,N_42423,N_42106);
nand U42955 (N_42955,N_42053,N_42339);
nand U42956 (N_42956,N_42118,N_42357);
nand U42957 (N_42957,N_42029,N_42306);
nand U42958 (N_42958,N_42090,N_42038);
nor U42959 (N_42959,N_42061,N_42492);
nor U42960 (N_42960,N_42427,N_42486);
xnor U42961 (N_42961,N_42166,N_42364);
nor U42962 (N_42962,N_42434,N_42222);
nand U42963 (N_42963,N_42121,N_42342);
or U42964 (N_42964,N_42150,N_42031);
or U42965 (N_42965,N_42081,N_42417);
and U42966 (N_42966,N_42001,N_42364);
nand U42967 (N_42967,N_42416,N_42237);
and U42968 (N_42968,N_42148,N_42462);
xor U42969 (N_42969,N_42081,N_42319);
nand U42970 (N_42970,N_42099,N_42163);
nand U42971 (N_42971,N_42106,N_42103);
or U42972 (N_42972,N_42118,N_42362);
xnor U42973 (N_42973,N_42179,N_42319);
xnor U42974 (N_42974,N_42420,N_42055);
nor U42975 (N_42975,N_42393,N_42024);
nor U42976 (N_42976,N_42164,N_42084);
nor U42977 (N_42977,N_42356,N_42169);
nor U42978 (N_42978,N_42363,N_42020);
and U42979 (N_42979,N_42318,N_42422);
or U42980 (N_42980,N_42057,N_42202);
and U42981 (N_42981,N_42047,N_42225);
xnor U42982 (N_42982,N_42050,N_42378);
and U42983 (N_42983,N_42063,N_42441);
nor U42984 (N_42984,N_42240,N_42092);
nor U42985 (N_42985,N_42031,N_42254);
or U42986 (N_42986,N_42276,N_42180);
nand U42987 (N_42987,N_42429,N_42469);
or U42988 (N_42988,N_42357,N_42441);
or U42989 (N_42989,N_42338,N_42410);
xnor U42990 (N_42990,N_42289,N_42007);
and U42991 (N_42991,N_42230,N_42393);
or U42992 (N_42992,N_42038,N_42242);
or U42993 (N_42993,N_42402,N_42055);
or U42994 (N_42994,N_42069,N_42401);
nor U42995 (N_42995,N_42386,N_42093);
and U42996 (N_42996,N_42218,N_42165);
or U42997 (N_42997,N_42149,N_42441);
or U42998 (N_42998,N_42379,N_42459);
xnor U42999 (N_42999,N_42238,N_42282);
and U43000 (N_43000,N_42861,N_42761);
nand U43001 (N_43001,N_42991,N_42688);
xnor U43002 (N_43002,N_42700,N_42945);
xnor U43003 (N_43003,N_42651,N_42915);
nor U43004 (N_43004,N_42649,N_42818);
nor U43005 (N_43005,N_42977,N_42607);
xor U43006 (N_43006,N_42880,N_42726);
and U43007 (N_43007,N_42696,N_42771);
nand U43008 (N_43008,N_42893,N_42703);
and U43009 (N_43009,N_42982,N_42691);
xor U43010 (N_43010,N_42512,N_42623);
and U43011 (N_43011,N_42645,N_42902);
nand U43012 (N_43012,N_42800,N_42657);
and U43013 (N_43013,N_42860,N_42821);
xor U43014 (N_43014,N_42981,N_42681);
or U43015 (N_43015,N_42823,N_42849);
or U43016 (N_43016,N_42674,N_42692);
nand U43017 (N_43017,N_42794,N_42807);
xor U43018 (N_43018,N_42805,N_42583);
and U43019 (N_43019,N_42628,N_42634);
nand U43020 (N_43020,N_42953,N_42752);
or U43021 (N_43021,N_42894,N_42716);
nand U43022 (N_43022,N_42775,N_42971);
or U43023 (N_43023,N_42882,N_42519);
nand U43024 (N_43024,N_42578,N_42906);
and U43025 (N_43025,N_42763,N_42970);
and U43026 (N_43026,N_42648,N_42784);
nor U43027 (N_43027,N_42773,N_42834);
xnor U43028 (N_43028,N_42878,N_42920);
or U43029 (N_43029,N_42898,N_42619);
xnor U43030 (N_43030,N_42711,N_42676);
and U43031 (N_43031,N_42741,N_42610);
nor U43032 (N_43032,N_42738,N_42613);
nor U43033 (N_43033,N_42647,N_42544);
nand U43034 (N_43034,N_42718,N_42901);
xnor U43035 (N_43035,N_42806,N_42632);
xnor U43036 (N_43036,N_42735,N_42660);
xnor U43037 (N_43037,N_42986,N_42956);
nor U43038 (N_43038,N_42922,N_42717);
nand U43039 (N_43039,N_42531,N_42702);
and U43040 (N_43040,N_42659,N_42847);
nor U43041 (N_43041,N_42586,N_42548);
nand U43042 (N_43042,N_42564,N_42995);
or U43043 (N_43043,N_42750,N_42863);
nor U43044 (N_43044,N_42809,N_42785);
or U43045 (N_43045,N_42677,N_42772);
or U43046 (N_43046,N_42862,N_42655);
xnor U43047 (N_43047,N_42639,N_42665);
nand U43048 (N_43048,N_42715,N_42984);
xor U43049 (N_43049,N_42932,N_42973);
or U43050 (N_43050,N_42875,N_42712);
or U43051 (N_43051,N_42916,N_42770);
nand U43052 (N_43052,N_42713,N_42527);
or U43053 (N_43053,N_42679,N_42796);
and U43054 (N_43054,N_42904,N_42903);
xor U43055 (N_43055,N_42781,N_42833);
nor U43056 (N_43056,N_42760,N_42988);
and U43057 (N_43057,N_42641,N_42517);
and U43058 (N_43058,N_42508,N_42615);
or U43059 (N_43059,N_42944,N_42708);
nand U43060 (N_43060,N_42671,N_42501);
xor U43061 (N_43061,N_42740,N_42857);
nor U43062 (N_43062,N_42686,N_42539);
nand U43063 (N_43063,N_42646,N_42502);
nor U43064 (N_43064,N_42558,N_42557);
nor U43065 (N_43065,N_42656,N_42574);
nand U43066 (N_43066,N_42598,N_42881);
nand U43067 (N_43067,N_42993,N_42859);
and U43068 (N_43068,N_42776,N_42758);
or U43069 (N_43069,N_42581,N_42840);
xor U43070 (N_43070,N_42798,N_42721);
nand U43071 (N_43071,N_42965,N_42745);
or U43072 (N_43072,N_42888,N_42816);
nor U43073 (N_43073,N_42998,N_42950);
or U43074 (N_43074,N_42852,N_42848);
nand U43075 (N_43075,N_42590,N_42941);
or U43076 (N_43076,N_42751,N_42670);
xor U43077 (N_43077,N_42789,N_42939);
nor U43078 (N_43078,N_42856,N_42839);
nand U43079 (N_43079,N_42997,N_42968);
and U43080 (N_43080,N_42573,N_42510);
or U43081 (N_43081,N_42966,N_42912);
nor U43082 (N_43082,N_42804,N_42780);
nand U43083 (N_43083,N_42680,N_42990);
or U43084 (N_43084,N_42961,N_42625);
xnor U43085 (N_43085,N_42536,N_42989);
nor U43086 (N_43086,N_42969,N_42710);
nor U43087 (N_43087,N_42528,N_42762);
xnor U43088 (N_43088,N_42795,N_42658);
nand U43089 (N_43089,N_42521,N_42801);
nor U43090 (N_43090,N_42778,N_42620);
nand U43091 (N_43091,N_42675,N_42533);
nor U43092 (N_43092,N_42911,N_42865);
and U43093 (N_43093,N_42522,N_42664);
nand U43094 (N_43094,N_42958,N_42940);
xor U43095 (N_43095,N_42782,N_42917);
or U43096 (N_43096,N_42790,N_42722);
or U43097 (N_43097,N_42684,N_42624);
xnor U43098 (N_43098,N_42803,N_42748);
nor U43099 (N_43099,N_42817,N_42814);
xnor U43100 (N_43100,N_42774,N_42899);
nor U43101 (N_43101,N_42541,N_42732);
nand U43102 (N_43102,N_42837,N_42720);
or U43103 (N_43103,N_42832,N_42886);
and U43104 (N_43104,N_42827,N_42829);
xnor U43105 (N_43105,N_42617,N_42864);
nand U43106 (N_43106,N_42608,N_42709);
nand U43107 (N_43107,N_42571,N_42652);
and U43108 (N_43108,N_42602,N_42727);
or U43109 (N_43109,N_42747,N_42810);
and U43110 (N_43110,N_42505,N_42570);
and U43111 (N_43111,N_42957,N_42719);
or U43112 (N_43112,N_42535,N_42767);
nor U43113 (N_43113,N_42537,N_42921);
and U43114 (N_43114,N_42813,N_42503);
or U43115 (N_43115,N_42918,N_42525);
xnor U43116 (N_43116,N_42695,N_42811);
and U43117 (N_43117,N_42855,N_42946);
nand U43118 (N_43118,N_42553,N_42947);
and U43119 (N_43119,N_42788,N_42975);
nand U43120 (N_43120,N_42900,N_42792);
or U43121 (N_43121,N_42520,N_42560);
and U43122 (N_43122,N_42577,N_42642);
xnor U43123 (N_43123,N_42985,N_42824);
xnor U43124 (N_43124,N_42601,N_42755);
and U43125 (N_43125,N_42669,N_42783);
or U43126 (N_43126,N_42731,N_42812);
nand U43127 (N_43127,N_42913,N_42643);
or U43128 (N_43128,N_42885,N_42593);
and U43129 (N_43129,N_42663,N_42928);
nand U43130 (N_43130,N_42538,N_42926);
xor U43131 (N_43131,N_42819,N_42935);
or U43132 (N_43132,N_42851,N_42756);
nand U43133 (N_43133,N_42938,N_42526);
xnor U43134 (N_43134,N_42631,N_42769);
and U43135 (N_43135,N_42908,N_42699);
nand U43136 (N_43136,N_42627,N_42714);
and U43137 (N_43137,N_42626,N_42568);
nor U43138 (N_43138,N_42737,N_42960);
nand U43139 (N_43139,N_42636,N_42511);
nand U43140 (N_43140,N_42614,N_42606);
and U43141 (N_43141,N_42838,N_42887);
nand U43142 (N_43142,N_42524,N_42513);
xor U43143 (N_43143,N_42869,N_42983);
and U43144 (N_43144,N_42556,N_42638);
or U43145 (N_43145,N_42575,N_42543);
xnor U43146 (N_43146,N_42846,N_42580);
nor U43147 (N_43147,N_42929,N_42516);
or U43148 (N_43148,N_42962,N_42959);
and U43149 (N_43149,N_42867,N_42698);
nor U43150 (N_43150,N_42919,N_42786);
nor U43151 (N_43151,N_42868,N_42640);
xnor U43152 (N_43152,N_42914,N_42948);
nor U43153 (N_43153,N_42896,N_42964);
nand U43154 (N_43154,N_42637,N_42994);
and U43155 (N_43155,N_42910,N_42793);
nand U43156 (N_43156,N_42844,N_42561);
and U43157 (N_43157,N_42843,N_42559);
and U43158 (N_43158,N_42723,N_42529);
nor U43159 (N_43159,N_42858,N_42841);
nand U43160 (N_43160,N_42579,N_42540);
xnor U43161 (N_43161,N_42611,N_42992);
or U43162 (N_43162,N_42890,N_42826);
nor U43163 (N_43163,N_42555,N_42584);
nand U43164 (N_43164,N_42588,N_42891);
or U43165 (N_43165,N_42980,N_42653);
and U43166 (N_43166,N_42753,N_42949);
xnor U43167 (N_43167,N_42542,N_42777);
xor U43168 (N_43168,N_42728,N_42854);
xor U43169 (N_43169,N_42759,N_42514);
nor U43170 (N_43170,N_42550,N_42853);
nor U43171 (N_43171,N_42974,N_42592);
nor U43172 (N_43172,N_42599,N_42565);
and U43173 (N_43173,N_42999,N_42546);
and U43174 (N_43174,N_42689,N_42621);
xnor U43175 (N_43175,N_42976,N_42884);
nand U43176 (N_43176,N_42654,N_42591);
nor U43177 (N_43177,N_42764,N_42567);
nor U43178 (N_43178,N_42706,N_42518);
nor U43179 (N_43179,N_42530,N_42551);
nor U43180 (N_43180,N_42683,N_42828);
xor U43181 (N_43181,N_42515,N_42967);
nor U43182 (N_43182,N_42630,N_42943);
nand U43183 (N_43183,N_42547,N_42933);
and U43184 (N_43184,N_42879,N_42927);
nor U43185 (N_43185,N_42729,N_42743);
nor U43186 (N_43186,N_42666,N_42820);
nand U43187 (N_43187,N_42797,N_42870);
nor U43188 (N_43188,N_42585,N_42616);
nand U43189 (N_43189,N_42566,N_42600);
nand U43190 (N_43190,N_42707,N_42787);
xnor U43191 (N_43191,N_42754,N_42835);
nor U43192 (N_43192,N_42701,N_42905);
nand U43193 (N_43193,N_42549,N_42594);
and U43194 (N_43194,N_42889,N_42799);
and U43195 (N_43195,N_42506,N_42609);
nand U43196 (N_43196,N_42831,N_42597);
xnor U43197 (N_43197,N_42576,N_42572);
nand U43198 (N_43198,N_42739,N_42768);
nor U43199 (N_43199,N_42589,N_42734);
nand U43200 (N_43200,N_42582,N_42872);
nand U43201 (N_43201,N_42825,N_42978);
nand U43202 (N_43202,N_42996,N_42936);
xor U43203 (N_43203,N_42629,N_42622);
nor U43204 (N_43204,N_42618,N_42633);
nor U43205 (N_43205,N_42987,N_42909);
or U43206 (N_43206,N_42907,N_42554);
and U43207 (N_43207,N_42563,N_42668);
xor U43208 (N_43208,N_42955,N_42523);
xor U43209 (N_43209,N_42963,N_42952);
or U43210 (N_43210,N_42500,N_42596);
xnor U43211 (N_43211,N_42562,N_42871);
or U43212 (N_43212,N_42667,N_42736);
and U43213 (N_43213,N_42746,N_42877);
or U43214 (N_43214,N_42866,N_42937);
and U43215 (N_43215,N_42690,N_42876);
and U43216 (N_43216,N_42534,N_42873);
nor U43217 (N_43217,N_42507,N_42842);
and U43218 (N_43218,N_42724,N_42730);
xor U43219 (N_43219,N_42874,N_42951);
nor U43220 (N_43220,N_42604,N_42704);
xor U43221 (N_43221,N_42509,N_42954);
nand U43222 (N_43222,N_42923,N_42694);
and U43223 (N_43223,N_42644,N_42979);
or U43224 (N_43224,N_42685,N_42765);
nand U43225 (N_43225,N_42836,N_42897);
nor U43226 (N_43226,N_42697,N_42749);
or U43227 (N_43227,N_42850,N_42552);
and U43228 (N_43228,N_42672,N_42612);
or U43229 (N_43229,N_42678,N_42742);
nand U43230 (N_43230,N_42766,N_42815);
and U43231 (N_43231,N_42605,N_42687);
and U43232 (N_43232,N_42504,N_42845);
nor U43233 (N_43233,N_42635,N_42883);
xnor U43234 (N_43234,N_42662,N_42587);
xor U43235 (N_43235,N_42830,N_42595);
nand U43236 (N_43236,N_42779,N_42791);
nor U43237 (N_43237,N_42808,N_42682);
nand U43238 (N_43238,N_42693,N_42930);
and U43239 (N_43239,N_42744,N_42650);
xnor U43240 (N_43240,N_42892,N_42822);
and U43241 (N_43241,N_42972,N_42931);
and U43242 (N_43242,N_42705,N_42733);
nand U43243 (N_43243,N_42569,N_42545);
xor U43244 (N_43244,N_42532,N_42924);
and U43245 (N_43245,N_42802,N_42934);
and U43246 (N_43246,N_42895,N_42725);
and U43247 (N_43247,N_42603,N_42661);
nand U43248 (N_43248,N_42925,N_42673);
and U43249 (N_43249,N_42942,N_42757);
xor U43250 (N_43250,N_42529,N_42941);
nor U43251 (N_43251,N_42954,N_42924);
nor U43252 (N_43252,N_42650,N_42536);
or U43253 (N_43253,N_42637,N_42883);
and U43254 (N_43254,N_42914,N_42974);
nor U43255 (N_43255,N_42781,N_42628);
and U43256 (N_43256,N_42793,N_42585);
or U43257 (N_43257,N_42891,N_42676);
and U43258 (N_43258,N_42511,N_42942);
nand U43259 (N_43259,N_42687,N_42844);
and U43260 (N_43260,N_42922,N_42991);
nand U43261 (N_43261,N_42510,N_42590);
and U43262 (N_43262,N_42837,N_42518);
nand U43263 (N_43263,N_42547,N_42571);
and U43264 (N_43264,N_42855,N_42629);
or U43265 (N_43265,N_42837,N_42582);
and U43266 (N_43266,N_42645,N_42719);
nor U43267 (N_43267,N_42896,N_42933);
nand U43268 (N_43268,N_42906,N_42781);
or U43269 (N_43269,N_42947,N_42780);
or U43270 (N_43270,N_42660,N_42975);
or U43271 (N_43271,N_42876,N_42829);
nand U43272 (N_43272,N_42687,N_42883);
and U43273 (N_43273,N_42556,N_42648);
nor U43274 (N_43274,N_42526,N_42891);
nand U43275 (N_43275,N_42572,N_42745);
nor U43276 (N_43276,N_42900,N_42931);
nand U43277 (N_43277,N_42977,N_42611);
and U43278 (N_43278,N_42570,N_42906);
and U43279 (N_43279,N_42971,N_42906);
or U43280 (N_43280,N_42919,N_42518);
or U43281 (N_43281,N_42538,N_42814);
nand U43282 (N_43282,N_42745,N_42855);
nor U43283 (N_43283,N_42700,N_42634);
nor U43284 (N_43284,N_42709,N_42813);
and U43285 (N_43285,N_42612,N_42718);
or U43286 (N_43286,N_42703,N_42936);
xnor U43287 (N_43287,N_42827,N_42593);
and U43288 (N_43288,N_42943,N_42993);
nor U43289 (N_43289,N_42501,N_42722);
and U43290 (N_43290,N_42988,N_42718);
nand U43291 (N_43291,N_42851,N_42814);
and U43292 (N_43292,N_42925,N_42891);
or U43293 (N_43293,N_42518,N_42736);
xor U43294 (N_43294,N_42889,N_42601);
nor U43295 (N_43295,N_42810,N_42619);
nand U43296 (N_43296,N_42743,N_42757);
nand U43297 (N_43297,N_42747,N_42966);
or U43298 (N_43298,N_42640,N_42512);
xnor U43299 (N_43299,N_42953,N_42725);
xor U43300 (N_43300,N_42664,N_42797);
and U43301 (N_43301,N_42504,N_42555);
nor U43302 (N_43302,N_42586,N_42620);
and U43303 (N_43303,N_42794,N_42574);
or U43304 (N_43304,N_42644,N_42838);
nand U43305 (N_43305,N_42885,N_42503);
xor U43306 (N_43306,N_42692,N_42689);
or U43307 (N_43307,N_42545,N_42802);
xor U43308 (N_43308,N_42961,N_42794);
and U43309 (N_43309,N_42731,N_42884);
or U43310 (N_43310,N_42549,N_42922);
nor U43311 (N_43311,N_42694,N_42603);
nor U43312 (N_43312,N_42977,N_42773);
and U43313 (N_43313,N_42835,N_42781);
or U43314 (N_43314,N_42501,N_42519);
xor U43315 (N_43315,N_42898,N_42734);
or U43316 (N_43316,N_42618,N_42622);
nor U43317 (N_43317,N_42503,N_42799);
xnor U43318 (N_43318,N_42760,N_42542);
nand U43319 (N_43319,N_42582,N_42784);
xor U43320 (N_43320,N_42976,N_42824);
or U43321 (N_43321,N_42907,N_42697);
and U43322 (N_43322,N_42908,N_42547);
or U43323 (N_43323,N_42621,N_42508);
xnor U43324 (N_43324,N_42863,N_42603);
nand U43325 (N_43325,N_42897,N_42743);
or U43326 (N_43326,N_42673,N_42803);
and U43327 (N_43327,N_42669,N_42722);
xor U43328 (N_43328,N_42897,N_42525);
nand U43329 (N_43329,N_42669,N_42589);
or U43330 (N_43330,N_42979,N_42686);
nand U43331 (N_43331,N_42786,N_42756);
xnor U43332 (N_43332,N_42645,N_42614);
or U43333 (N_43333,N_42786,N_42799);
nand U43334 (N_43334,N_42574,N_42501);
or U43335 (N_43335,N_42961,N_42686);
xor U43336 (N_43336,N_42522,N_42548);
or U43337 (N_43337,N_42993,N_42990);
xor U43338 (N_43338,N_42985,N_42603);
and U43339 (N_43339,N_42920,N_42986);
nor U43340 (N_43340,N_42878,N_42552);
and U43341 (N_43341,N_42511,N_42507);
or U43342 (N_43342,N_42963,N_42647);
nand U43343 (N_43343,N_42547,N_42647);
or U43344 (N_43344,N_42848,N_42854);
and U43345 (N_43345,N_42563,N_42819);
nand U43346 (N_43346,N_42575,N_42973);
nand U43347 (N_43347,N_42649,N_42908);
nor U43348 (N_43348,N_42616,N_42763);
nor U43349 (N_43349,N_42892,N_42867);
xnor U43350 (N_43350,N_42955,N_42755);
xor U43351 (N_43351,N_42702,N_42786);
or U43352 (N_43352,N_42703,N_42808);
nand U43353 (N_43353,N_42546,N_42920);
or U43354 (N_43354,N_42517,N_42950);
and U43355 (N_43355,N_42684,N_42660);
xor U43356 (N_43356,N_42583,N_42785);
xor U43357 (N_43357,N_42630,N_42876);
xor U43358 (N_43358,N_42933,N_42569);
xnor U43359 (N_43359,N_42965,N_42707);
nor U43360 (N_43360,N_42520,N_42854);
xor U43361 (N_43361,N_42948,N_42545);
and U43362 (N_43362,N_42802,N_42854);
or U43363 (N_43363,N_42961,N_42752);
nand U43364 (N_43364,N_42624,N_42880);
xnor U43365 (N_43365,N_42898,N_42763);
nand U43366 (N_43366,N_42982,N_42743);
and U43367 (N_43367,N_42605,N_42619);
or U43368 (N_43368,N_42846,N_42528);
or U43369 (N_43369,N_42812,N_42694);
or U43370 (N_43370,N_42952,N_42773);
nand U43371 (N_43371,N_42941,N_42636);
or U43372 (N_43372,N_42994,N_42715);
or U43373 (N_43373,N_42662,N_42506);
or U43374 (N_43374,N_42723,N_42876);
and U43375 (N_43375,N_42969,N_42813);
and U43376 (N_43376,N_42914,N_42846);
and U43377 (N_43377,N_42816,N_42708);
and U43378 (N_43378,N_42643,N_42697);
and U43379 (N_43379,N_42806,N_42634);
nand U43380 (N_43380,N_42675,N_42526);
nor U43381 (N_43381,N_42895,N_42612);
or U43382 (N_43382,N_42920,N_42929);
nand U43383 (N_43383,N_42746,N_42955);
or U43384 (N_43384,N_42542,N_42802);
or U43385 (N_43385,N_42576,N_42814);
xnor U43386 (N_43386,N_42727,N_42555);
nand U43387 (N_43387,N_42824,N_42826);
nand U43388 (N_43388,N_42998,N_42660);
nor U43389 (N_43389,N_42589,N_42608);
nand U43390 (N_43390,N_42696,N_42839);
nor U43391 (N_43391,N_42722,N_42519);
xor U43392 (N_43392,N_42776,N_42680);
or U43393 (N_43393,N_42692,N_42873);
and U43394 (N_43394,N_42515,N_42542);
xnor U43395 (N_43395,N_42927,N_42880);
and U43396 (N_43396,N_42922,N_42893);
xor U43397 (N_43397,N_42887,N_42659);
or U43398 (N_43398,N_42823,N_42736);
nor U43399 (N_43399,N_42941,N_42611);
and U43400 (N_43400,N_42800,N_42802);
nand U43401 (N_43401,N_42592,N_42505);
and U43402 (N_43402,N_42990,N_42894);
nand U43403 (N_43403,N_42562,N_42628);
nand U43404 (N_43404,N_42988,N_42727);
xnor U43405 (N_43405,N_42979,N_42786);
nor U43406 (N_43406,N_42891,N_42974);
or U43407 (N_43407,N_42997,N_42514);
and U43408 (N_43408,N_42903,N_42576);
nor U43409 (N_43409,N_42943,N_42519);
xor U43410 (N_43410,N_42513,N_42787);
nand U43411 (N_43411,N_42705,N_42559);
nor U43412 (N_43412,N_42945,N_42659);
or U43413 (N_43413,N_42608,N_42859);
nand U43414 (N_43414,N_42514,N_42727);
and U43415 (N_43415,N_42599,N_42931);
nor U43416 (N_43416,N_42581,N_42523);
and U43417 (N_43417,N_42791,N_42626);
nor U43418 (N_43418,N_42805,N_42593);
nand U43419 (N_43419,N_42555,N_42963);
nor U43420 (N_43420,N_42933,N_42644);
or U43421 (N_43421,N_42951,N_42725);
xnor U43422 (N_43422,N_42835,N_42977);
or U43423 (N_43423,N_42746,N_42870);
nand U43424 (N_43424,N_42998,N_42511);
xnor U43425 (N_43425,N_42744,N_42894);
xor U43426 (N_43426,N_42560,N_42912);
and U43427 (N_43427,N_42705,N_42997);
and U43428 (N_43428,N_42589,N_42983);
nor U43429 (N_43429,N_42566,N_42551);
or U43430 (N_43430,N_42987,N_42947);
nand U43431 (N_43431,N_42753,N_42964);
and U43432 (N_43432,N_42997,N_42885);
nand U43433 (N_43433,N_42852,N_42509);
xor U43434 (N_43434,N_42769,N_42781);
nand U43435 (N_43435,N_42581,N_42770);
or U43436 (N_43436,N_42567,N_42753);
nand U43437 (N_43437,N_42821,N_42522);
nor U43438 (N_43438,N_42844,N_42830);
or U43439 (N_43439,N_42611,N_42775);
xor U43440 (N_43440,N_42955,N_42597);
nand U43441 (N_43441,N_42714,N_42533);
nand U43442 (N_43442,N_42998,N_42548);
nand U43443 (N_43443,N_42618,N_42773);
and U43444 (N_43444,N_42685,N_42569);
and U43445 (N_43445,N_42673,N_42793);
and U43446 (N_43446,N_42828,N_42819);
or U43447 (N_43447,N_42800,N_42949);
and U43448 (N_43448,N_42510,N_42629);
and U43449 (N_43449,N_42813,N_42670);
xor U43450 (N_43450,N_42999,N_42525);
nand U43451 (N_43451,N_42515,N_42868);
nand U43452 (N_43452,N_42839,N_42644);
nand U43453 (N_43453,N_42551,N_42700);
or U43454 (N_43454,N_42649,N_42645);
xor U43455 (N_43455,N_42573,N_42995);
or U43456 (N_43456,N_42942,N_42876);
xnor U43457 (N_43457,N_42935,N_42759);
nor U43458 (N_43458,N_42675,N_42792);
or U43459 (N_43459,N_42794,N_42575);
and U43460 (N_43460,N_42787,N_42851);
nor U43461 (N_43461,N_42567,N_42826);
and U43462 (N_43462,N_42918,N_42709);
or U43463 (N_43463,N_42533,N_42541);
nand U43464 (N_43464,N_42683,N_42907);
xnor U43465 (N_43465,N_42672,N_42500);
nand U43466 (N_43466,N_42856,N_42622);
nor U43467 (N_43467,N_42730,N_42800);
or U43468 (N_43468,N_42875,N_42562);
or U43469 (N_43469,N_42532,N_42944);
nand U43470 (N_43470,N_42597,N_42825);
nand U43471 (N_43471,N_42656,N_42844);
and U43472 (N_43472,N_42829,N_42601);
and U43473 (N_43473,N_42771,N_42755);
nand U43474 (N_43474,N_42591,N_42831);
nor U43475 (N_43475,N_42852,N_42591);
xnor U43476 (N_43476,N_42602,N_42550);
or U43477 (N_43477,N_42626,N_42866);
xnor U43478 (N_43478,N_42756,N_42930);
and U43479 (N_43479,N_42817,N_42611);
nand U43480 (N_43480,N_42736,N_42604);
xor U43481 (N_43481,N_42530,N_42879);
nor U43482 (N_43482,N_42746,N_42928);
and U43483 (N_43483,N_42727,N_42733);
nand U43484 (N_43484,N_42898,N_42833);
nand U43485 (N_43485,N_42913,N_42965);
xnor U43486 (N_43486,N_42885,N_42716);
and U43487 (N_43487,N_42929,N_42978);
xnor U43488 (N_43488,N_42947,N_42817);
and U43489 (N_43489,N_42602,N_42553);
or U43490 (N_43490,N_42754,N_42893);
xor U43491 (N_43491,N_42735,N_42727);
nor U43492 (N_43492,N_42886,N_42806);
and U43493 (N_43493,N_42900,N_42781);
and U43494 (N_43494,N_42580,N_42990);
nor U43495 (N_43495,N_42606,N_42882);
and U43496 (N_43496,N_42937,N_42842);
and U43497 (N_43497,N_42816,N_42528);
nor U43498 (N_43498,N_42663,N_42522);
xor U43499 (N_43499,N_42641,N_42608);
nor U43500 (N_43500,N_43163,N_43084);
and U43501 (N_43501,N_43379,N_43407);
nor U43502 (N_43502,N_43293,N_43273);
and U43503 (N_43503,N_43030,N_43111);
nand U43504 (N_43504,N_43313,N_43005);
and U43505 (N_43505,N_43485,N_43083);
xor U43506 (N_43506,N_43035,N_43464);
nor U43507 (N_43507,N_43460,N_43275);
xor U43508 (N_43508,N_43126,N_43215);
or U43509 (N_43509,N_43272,N_43259);
xor U43510 (N_43510,N_43318,N_43423);
nand U43511 (N_43511,N_43238,N_43302);
or U43512 (N_43512,N_43101,N_43227);
or U43513 (N_43513,N_43297,N_43144);
xnor U43514 (N_43514,N_43374,N_43304);
nor U43515 (N_43515,N_43172,N_43298);
nor U43516 (N_43516,N_43489,N_43086);
nor U43517 (N_43517,N_43129,N_43003);
or U43518 (N_43518,N_43271,N_43384);
nor U43519 (N_43519,N_43036,N_43396);
xnor U43520 (N_43520,N_43029,N_43143);
xnor U43521 (N_43521,N_43109,N_43233);
nor U43522 (N_43522,N_43236,N_43353);
nand U43523 (N_43523,N_43355,N_43179);
nand U43524 (N_43524,N_43477,N_43327);
or U43525 (N_43525,N_43409,N_43173);
and U43526 (N_43526,N_43204,N_43322);
or U43527 (N_43527,N_43441,N_43157);
nand U43528 (N_43528,N_43066,N_43253);
and U43529 (N_43529,N_43419,N_43262);
or U43530 (N_43530,N_43132,N_43082);
or U43531 (N_43531,N_43010,N_43232);
nor U43532 (N_43532,N_43019,N_43367);
xor U43533 (N_43533,N_43100,N_43254);
nor U43534 (N_43534,N_43321,N_43376);
nand U43535 (N_43535,N_43094,N_43147);
nand U43536 (N_43536,N_43332,N_43424);
or U43537 (N_43537,N_43291,N_43231);
nor U43538 (N_43538,N_43133,N_43241);
nand U43539 (N_43539,N_43404,N_43440);
nor U43540 (N_43540,N_43124,N_43224);
and U43541 (N_43541,N_43288,N_43207);
nand U43542 (N_43542,N_43405,N_43043);
nand U43543 (N_43543,N_43027,N_43442);
xnor U43544 (N_43544,N_43471,N_43076);
nand U43545 (N_43545,N_43252,N_43198);
nor U43546 (N_43546,N_43316,N_43184);
nor U43547 (N_43547,N_43075,N_43209);
nor U43548 (N_43548,N_43142,N_43369);
nand U43549 (N_43549,N_43130,N_43039);
and U43550 (N_43550,N_43497,N_43145);
or U43551 (N_43551,N_43325,N_43337);
xor U43552 (N_43552,N_43072,N_43432);
nor U43553 (N_43553,N_43278,N_43422);
or U43554 (N_43554,N_43377,N_43438);
and U43555 (N_43555,N_43333,N_43170);
xnor U43556 (N_43556,N_43092,N_43156);
xor U43557 (N_43557,N_43223,N_43020);
nand U43558 (N_43558,N_43491,N_43340);
xor U43559 (N_43559,N_43052,N_43183);
nor U43560 (N_43560,N_43115,N_43444);
or U43561 (N_43561,N_43411,N_43475);
nor U43562 (N_43562,N_43166,N_43093);
nor U43563 (N_43563,N_43174,N_43118);
or U43564 (N_43564,N_43199,N_43201);
and U43565 (N_43565,N_43447,N_43339);
or U43566 (N_43566,N_43108,N_43021);
and U43567 (N_43567,N_43059,N_43090);
xnor U43568 (N_43568,N_43269,N_43373);
nand U43569 (N_43569,N_43364,N_43413);
or U43570 (N_43570,N_43014,N_43192);
xnor U43571 (N_43571,N_43081,N_43312);
xnor U43572 (N_43572,N_43496,N_43387);
xor U43573 (N_43573,N_43343,N_43177);
nor U43574 (N_43574,N_43200,N_43013);
xnor U43575 (N_43575,N_43079,N_43397);
or U43576 (N_43576,N_43127,N_43285);
or U43577 (N_43577,N_43452,N_43385);
or U43578 (N_43578,N_43239,N_43334);
nor U43579 (N_43579,N_43294,N_43160);
nand U43580 (N_43580,N_43435,N_43243);
or U43581 (N_43581,N_43328,N_43141);
nor U43582 (N_43582,N_43153,N_43481);
nand U43583 (N_43583,N_43168,N_43033);
nand U43584 (N_43584,N_43214,N_43457);
or U43585 (N_43585,N_43242,N_43360);
nor U43586 (N_43586,N_43336,N_43088);
nor U43587 (N_43587,N_43067,N_43063);
or U43588 (N_43588,N_43220,N_43182);
nand U43589 (N_43589,N_43000,N_43098);
and U43590 (N_43590,N_43228,N_43210);
xnor U43591 (N_43591,N_43078,N_43258);
xor U43592 (N_43592,N_43372,N_43046);
or U43593 (N_43593,N_43351,N_43483);
and U43594 (N_43594,N_43274,N_43261);
xnor U43595 (N_43595,N_43050,N_43037);
nor U43596 (N_43596,N_43468,N_43264);
and U43597 (N_43597,N_43329,N_43338);
nor U43598 (N_43598,N_43474,N_43265);
and U43599 (N_43599,N_43450,N_43426);
nor U43600 (N_43600,N_43017,N_43176);
or U43601 (N_43601,N_43068,N_43159);
xor U43602 (N_43602,N_43001,N_43097);
or U43603 (N_43603,N_43152,N_43248);
xor U43604 (N_43604,N_43197,N_43024);
or U43605 (N_43605,N_43064,N_43125);
nand U43606 (N_43606,N_43492,N_43401);
nand U43607 (N_43607,N_43493,N_43455);
and U43608 (N_43608,N_43465,N_43439);
or U43609 (N_43609,N_43410,N_43323);
nand U43610 (N_43610,N_43417,N_43317);
nand U43611 (N_43611,N_43008,N_43105);
and U43612 (N_43612,N_43453,N_43368);
or U43613 (N_43613,N_43263,N_43418);
or U43614 (N_43614,N_43416,N_43139);
or U43615 (N_43615,N_43018,N_43476);
nor U43616 (N_43616,N_43283,N_43301);
nor U43617 (N_43617,N_43307,N_43473);
xor U43618 (N_43618,N_43221,N_43131);
or U43619 (N_43619,N_43255,N_43038);
nand U43620 (N_43620,N_43470,N_43406);
nand U43621 (N_43621,N_43311,N_43023);
nand U43622 (N_43622,N_43106,N_43303);
and U43623 (N_43623,N_43393,N_43467);
nand U43624 (N_43624,N_43281,N_43110);
nor U43625 (N_43625,N_43390,N_43004);
and U43626 (N_43626,N_43137,N_43498);
or U43627 (N_43627,N_43292,N_43099);
nand U43628 (N_43628,N_43022,N_43349);
xor U43629 (N_43629,N_43234,N_43446);
and U43630 (N_43630,N_43026,N_43378);
and U43631 (N_43631,N_43382,N_43472);
nor U43632 (N_43632,N_43392,N_43122);
or U43633 (N_43633,N_43305,N_43226);
nand U43634 (N_43634,N_43451,N_43188);
nand U43635 (N_43635,N_43280,N_43459);
xnor U43636 (N_43636,N_43403,N_43314);
nor U43637 (N_43637,N_43429,N_43202);
or U43638 (N_43638,N_43400,N_43245);
and U43639 (N_43639,N_43454,N_43237);
xor U43640 (N_43640,N_43229,N_43268);
or U43641 (N_43641,N_43103,N_43345);
xor U43642 (N_43642,N_43140,N_43462);
and U43643 (N_43643,N_43434,N_43398);
and U43644 (N_43644,N_43060,N_43388);
or U43645 (N_43645,N_43062,N_43123);
nand U43646 (N_43646,N_43348,N_43162);
xnor U43647 (N_43647,N_43276,N_43296);
nand U43648 (N_43648,N_43138,N_43445);
or U43649 (N_43649,N_43203,N_43165);
nand U43650 (N_43650,N_43175,N_43433);
nand U43651 (N_43651,N_43495,N_43102);
nor U43652 (N_43652,N_43191,N_43117);
or U43653 (N_43653,N_43354,N_43344);
nand U43654 (N_43654,N_43194,N_43096);
or U43655 (N_43655,N_43015,N_43282);
xor U43656 (N_43656,N_43463,N_43150);
and U43657 (N_43657,N_43352,N_43213);
or U43658 (N_43658,N_43069,N_43412);
nor U43659 (N_43659,N_43222,N_43381);
or U43660 (N_43660,N_43295,N_43335);
and U43661 (N_43661,N_43246,N_43041);
or U43662 (N_43662,N_43119,N_43225);
nand U43663 (N_43663,N_43428,N_43324);
xor U43664 (N_43664,N_43486,N_43080);
and U43665 (N_43665,N_43217,N_43430);
nand U43666 (N_43666,N_43386,N_43134);
nor U43667 (N_43667,N_43040,N_43112);
and U43668 (N_43668,N_43308,N_43420);
and U43669 (N_43669,N_43421,N_43290);
nor U43670 (N_43670,N_43006,N_43186);
and U43671 (N_43671,N_43074,N_43104);
xor U43672 (N_43672,N_43009,N_43257);
and U43673 (N_43673,N_43116,N_43371);
and U43674 (N_43674,N_43151,N_43055);
nor U43675 (N_43675,N_43399,N_43331);
nand U43676 (N_43676,N_43011,N_43149);
and U43677 (N_43677,N_43230,N_43240);
or U43678 (N_43678,N_43048,N_43185);
nand U43679 (N_43679,N_43270,N_43427);
or U43680 (N_43680,N_43181,N_43095);
and U43681 (N_43681,N_43077,N_43089);
nand U43682 (N_43682,N_43414,N_43395);
xor U43683 (N_43683,N_43205,N_43437);
nand U43684 (N_43684,N_43330,N_43458);
xor U43685 (N_43685,N_43091,N_43286);
xnor U43686 (N_43686,N_43180,N_43206);
xnor U43687 (N_43687,N_43061,N_43361);
nand U43688 (N_43688,N_43365,N_43148);
and U43689 (N_43689,N_43244,N_43466);
xnor U43690 (N_43690,N_43190,N_43164);
and U43691 (N_43691,N_43025,N_43488);
and U43692 (N_43692,N_43034,N_43235);
or U43693 (N_43693,N_43251,N_43212);
nand U43694 (N_43694,N_43211,N_43267);
xnor U43695 (N_43695,N_43266,N_43249);
nor U43696 (N_43696,N_43047,N_43482);
xnor U43697 (N_43697,N_43044,N_43425);
nand U43698 (N_43698,N_43058,N_43320);
nand U43699 (N_43699,N_43260,N_43187);
nor U43700 (N_43700,N_43208,N_43449);
or U43701 (N_43701,N_43490,N_43049);
nand U43702 (N_43702,N_43277,N_43279);
or U43703 (N_43703,N_43402,N_43347);
nand U43704 (N_43704,N_43120,N_43341);
and U43705 (N_43705,N_43007,N_43287);
and U43706 (N_43706,N_43219,N_43107);
xnor U43707 (N_43707,N_43350,N_43216);
nand U43708 (N_43708,N_43073,N_43196);
and U43709 (N_43709,N_43358,N_43045);
nor U43710 (N_43710,N_43002,N_43370);
nand U43711 (N_43711,N_43146,N_43487);
nand U43712 (N_43712,N_43306,N_43250);
nand U43713 (N_43713,N_43389,N_43167);
nor U43714 (N_43714,N_43247,N_43016);
nand U43715 (N_43715,N_43478,N_43289);
nand U43716 (N_43716,N_43469,N_43443);
nand U43717 (N_43717,N_43342,N_43070);
and U43718 (N_43718,N_43408,N_43113);
or U43719 (N_43719,N_43031,N_43193);
nor U43720 (N_43720,N_43032,N_43284);
nand U43721 (N_43721,N_43456,N_43383);
and U43722 (N_43722,N_43054,N_43431);
nand U43723 (N_43723,N_43326,N_43494);
or U43724 (N_43724,N_43087,N_43499);
nand U43725 (N_43725,N_43359,N_43256);
nand U43726 (N_43726,N_43309,N_43218);
nor U43727 (N_43727,N_43394,N_43319);
nand U43728 (N_43728,N_43158,N_43357);
and U43729 (N_43729,N_43315,N_43356);
xor U43730 (N_43730,N_43178,N_43362);
nor U43731 (N_43731,N_43135,N_43380);
xor U43732 (N_43732,N_43480,N_43028);
or U43733 (N_43733,N_43366,N_43161);
nand U43734 (N_43734,N_43155,N_43057);
xor U43735 (N_43735,N_43299,N_43346);
and U43736 (N_43736,N_43310,N_43484);
nand U43737 (N_43737,N_43136,N_43051);
nand U43738 (N_43738,N_43189,N_43121);
or U43739 (N_43739,N_43461,N_43071);
xor U43740 (N_43740,N_43053,N_43195);
or U43741 (N_43741,N_43042,N_43065);
and U43742 (N_43742,N_43415,N_43479);
or U43743 (N_43743,N_43114,N_43300);
nand U43744 (N_43744,N_43169,N_43056);
xnor U43745 (N_43745,N_43012,N_43391);
or U43746 (N_43746,N_43128,N_43154);
xnor U43747 (N_43747,N_43363,N_43448);
nor U43748 (N_43748,N_43375,N_43436);
and U43749 (N_43749,N_43085,N_43171);
or U43750 (N_43750,N_43138,N_43297);
or U43751 (N_43751,N_43364,N_43087);
xor U43752 (N_43752,N_43455,N_43093);
nand U43753 (N_43753,N_43485,N_43374);
or U43754 (N_43754,N_43263,N_43028);
or U43755 (N_43755,N_43126,N_43106);
nor U43756 (N_43756,N_43253,N_43049);
and U43757 (N_43757,N_43405,N_43329);
nor U43758 (N_43758,N_43236,N_43270);
xnor U43759 (N_43759,N_43233,N_43342);
nor U43760 (N_43760,N_43279,N_43402);
xnor U43761 (N_43761,N_43039,N_43306);
or U43762 (N_43762,N_43111,N_43283);
or U43763 (N_43763,N_43212,N_43499);
nand U43764 (N_43764,N_43482,N_43245);
xnor U43765 (N_43765,N_43449,N_43407);
and U43766 (N_43766,N_43418,N_43182);
and U43767 (N_43767,N_43454,N_43372);
or U43768 (N_43768,N_43158,N_43134);
nand U43769 (N_43769,N_43492,N_43344);
nor U43770 (N_43770,N_43443,N_43008);
and U43771 (N_43771,N_43071,N_43107);
nor U43772 (N_43772,N_43382,N_43261);
nor U43773 (N_43773,N_43496,N_43104);
and U43774 (N_43774,N_43049,N_43154);
or U43775 (N_43775,N_43168,N_43389);
nor U43776 (N_43776,N_43232,N_43107);
xor U43777 (N_43777,N_43405,N_43412);
nor U43778 (N_43778,N_43259,N_43326);
xnor U43779 (N_43779,N_43439,N_43252);
and U43780 (N_43780,N_43472,N_43375);
and U43781 (N_43781,N_43405,N_43110);
nor U43782 (N_43782,N_43319,N_43385);
nand U43783 (N_43783,N_43366,N_43095);
nor U43784 (N_43784,N_43128,N_43015);
xnor U43785 (N_43785,N_43412,N_43388);
and U43786 (N_43786,N_43433,N_43251);
or U43787 (N_43787,N_43410,N_43491);
xor U43788 (N_43788,N_43155,N_43222);
or U43789 (N_43789,N_43175,N_43063);
and U43790 (N_43790,N_43288,N_43448);
or U43791 (N_43791,N_43038,N_43008);
or U43792 (N_43792,N_43468,N_43412);
and U43793 (N_43793,N_43004,N_43239);
nand U43794 (N_43794,N_43313,N_43421);
nand U43795 (N_43795,N_43448,N_43424);
or U43796 (N_43796,N_43411,N_43166);
nor U43797 (N_43797,N_43309,N_43065);
xnor U43798 (N_43798,N_43224,N_43150);
or U43799 (N_43799,N_43481,N_43308);
nand U43800 (N_43800,N_43111,N_43354);
or U43801 (N_43801,N_43068,N_43188);
nand U43802 (N_43802,N_43419,N_43318);
and U43803 (N_43803,N_43331,N_43397);
nand U43804 (N_43804,N_43468,N_43097);
xnor U43805 (N_43805,N_43152,N_43125);
nor U43806 (N_43806,N_43270,N_43452);
and U43807 (N_43807,N_43487,N_43194);
nand U43808 (N_43808,N_43379,N_43441);
and U43809 (N_43809,N_43141,N_43152);
xor U43810 (N_43810,N_43227,N_43165);
and U43811 (N_43811,N_43074,N_43492);
xor U43812 (N_43812,N_43408,N_43121);
or U43813 (N_43813,N_43262,N_43035);
nand U43814 (N_43814,N_43284,N_43087);
and U43815 (N_43815,N_43126,N_43206);
or U43816 (N_43816,N_43428,N_43206);
nand U43817 (N_43817,N_43005,N_43057);
nor U43818 (N_43818,N_43000,N_43077);
or U43819 (N_43819,N_43001,N_43187);
and U43820 (N_43820,N_43487,N_43449);
or U43821 (N_43821,N_43098,N_43241);
or U43822 (N_43822,N_43233,N_43331);
nor U43823 (N_43823,N_43065,N_43099);
xor U43824 (N_43824,N_43290,N_43001);
or U43825 (N_43825,N_43460,N_43465);
xnor U43826 (N_43826,N_43367,N_43084);
xnor U43827 (N_43827,N_43083,N_43215);
or U43828 (N_43828,N_43101,N_43186);
and U43829 (N_43829,N_43343,N_43262);
and U43830 (N_43830,N_43248,N_43238);
and U43831 (N_43831,N_43345,N_43251);
nor U43832 (N_43832,N_43292,N_43208);
nand U43833 (N_43833,N_43445,N_43394);
and U43834 (N_43834,N_43355,N_43470);
nand U43835 (N_43835,N_43141,N_43356);
and U43836 (N_43836,N_43120,N_43320);
or U43837 (N_43837,N_43358,N_43171);
nand U43838 (N_43838,N_43180,N_43186);
or U43839 (N_43839,N_43422,N_43361);
xor U43840 (N_43840,N_43486,N_43472);
nand U43841 (N_43841,N_43327,N_43219);
and U43842 (N_43842,N_43399,N_43297);
nor U43843 (N_43843,N_43302,N_43476);
nor U43844 (N_43844,N_43243,N_43413);
nand U43845 (N_43845,N_43376,N_43107);
or U43846 (N_43846,N_43007,N_43232);
or U43847 (N_43847,N_43339,N_43046);
or U43848 (N_43848,N_43229,N_43021);
or U43849 (N_43849,N_43138,N_43313);
xor U43850 (N_43850,N_43301,N_43460);
or U43851 (N_43851,N_43148,N_43461);
xor U43852 (N_43852,N_43146,N_43159);
nor U43853 (N_43853,N_43315,N_43305);
xor U43854 (N_43854,N_43189,N_43429);
nand U43855 (N_43855,N_43060,N_43069);
nor U43856 (N_43856,N_43213,N_43095);
nand U43857 (N_43857,N_43085,N_43084);
xnor U43858 (N_43858,N_43147,N_43353);
and U43859 (N_43859,N_43146,N_43206);
and U43860 (N_43860,N_43292,N_43004);
or U43861 (N_43861,N_43258,N_43396);
or U43862 (N_43862,N_43111,N_43369);
nand U43863 (N_43863,N_43259,N_43274);
nor U43864 (N_43864,N_43292,N_43253);
xnor U43865 (N_43865,N_43410,N_43168);
xnor U43866 (N_43866,N_43335,N_43366);
xnor U43867 (N_43867,N_43079,N_43194);
and U43868 (N_43868,N_43127,N_43216);
or U43869 (N_43869,N_43187,N_43013);
xor U43870 (N_43870,N_43405,N_43480);
xor U43871 (N_43871,N_43016,N_43017);
nor U43872 (N_43872,N_43451,N_43316);
or U43873 (N_43873,N_43482,N_43301);
and U43874 (N_43874,N_43197,N_43246);
nand U43875 (N_43875,N_43150,N_43130);
xnor U43876 (N_43876,N_43427,N_43220);
xor U43877 (N_43877,N_43175,N_43156);
xnor U43878 (N_43878,N_43234,N_43060);
nor U43879 (N_43879,N_43087,N_43311);
or U43880 (N_43880,N_43019,N_43036);
and U43881 (N_43881,N_43171,N_43148);
or U43882 (N_43882,N_43231,N_43410);
or U43883 (N_43883,N_43007,N_43238);
xnor U43884 (N_43884,N_43283,N_43464);
and U43885 (N_43885,N_43187,N_43241);
nand U43886 (N_43886,N_43274,N_43350);
xnor U43887 (N_43887,N_43276,N_43210);
xnor U43888 (N_43888,N_43341,N_43162);
and U43889 (N_43889,N_43178,N_43244);
or U43890 (N_43890,N_43343,N_43173);
or U43891 (N_43891,N_43365,N_43376);
and U43892 (N_43892,N_43223,N_43013);
or U43893 (N_43893,N_43461,N_43213);
and U43894 (N_43894,N_43341,N_43362);
nand U43895 (N_43895,N_43278,N_43344);
nand U43896 (N_43896,N_43365,N_43332);
nand U43897 (N_43897,N_43135,N_43229);
or U43898 (N_43898,N_43196,N_43027);
xor U43899 (N_43899,N_43165,N_43489);
and U43900 (N_43900,N_43429,N_43128);
or U43901 (N_43901,N_43093,N_43067);
nor U43902 (N_43902,N_43488,N_43463);
and U43903 (N_43903,N_43190,N_43159);
or U43904 (N_43904,N_43184,N_43325);
or U43905 (N_43905,N_43210,N_43159);
xnor U43906 (N_43906,N_43403,N_43059);
or U43907 (N_43907,N_43274,N_43051);
and U43908 (N_43908,N_43454,N_43140);
or U43909 (N_43909,N_43316,N_43383);
xor U43910 (N_43910,N_43466,N_43102);
or U43911 (N_43911,N_43418,N_43176);
nor U43912 (N_43912,N_43173,N_43076);
nor U43913 (N_43913,N_43283,N_43447);
or U43914 (N_43914,N_43498,N_43119);
and U43915 (N_43915,N_43452,N_43233);
nor U43916 (N_43916,N_43411,N_43442);
or U43917 (N_43917,N_43176,N_43214);
nor U43918 (N_43918,N_43403,N_43465);
and U43919 (N_43919,N_43117,N_43208);
xnor U43920 (N_43920,N_43299,N_43041);
and U43921 (N_43921,N_43276,N_43357);
nor U43922 (N_43922,N_43337,N_43029);
nor U43923 (N_43923,N_43487,N_43344);
nand U43924 (N_43924,N_43007,N_43052);
nand U43925 (N_43925,N_43037,N_43271);
nand U43926 (N_43926,N_43104,N_43174);
and U43927 (N_43927,N_43194,N_43033);
and U43928 (N_43928,N_43392,N_43246);
xnor U43929 (N_43929,N_43080,N_43365);
nand U43930 (N_43930,N_43113,N_43385);
xnor U43931 (N_43931,N_43319,N_43200);
and U43932 (N_43932,N_43167,N_43417);
or U43933 (N_43933,N_43452,N_43297);
or U43934 (N_43934,N_43167,N_43498);
or U43935 (N_43935,N_43250,N_43438);
or U43936 (N_43936,N_43162,N_43473);
nand U43937 (N_43937,N_43410,N_43285);
and U43938 (N_43938,N_43287,N_43031);
nor U43939 (N_43939,N_43211,N_43136);
and U43940 (N_43940,N_43490,N_43036);
xor U43941 (N_43941,N_43380,N_43298);
or U43942 (N_43942,N_43385,N_43107);
xor U43943 (N_43943,N_43383,N_43271);
xor U43944 (N_43944,N_43258,N_43019);
and U43945 (N_43945,N_43335,N_43494);
or U43946 (N_43946,N_43467,N_43160);
nand U43947 (N_43947,N_43131,N_43136);
and U43948 (N_43948,N_43267,N_43497);
xnor U43949 (N_43949,N_43242,N_43350);
xor U43950 (N_43950,N_43025,N_43250);
nand U43951 (N_43951,N_43297,N_43223);
nand U43952 (N_43952,N_43284,N_43081);
nor U43953 (N_43953,N_43151,N_43160);
or U43954 (N_43954,N_43235,N_43421);
and U43955 (N_43955,N_43202,N_43344);
and U43956 (N_43956,N_43192,N_43451);
or U43957 (N_43957,N_43471,N_43356);
or U43958 (N_43958,N_43005,N_43357);
nand U43959 (N_43959,N_43249,N_43448);
or U43960 (N_43960,N_43294,N_43384);
nand U43961 (N_43961,N_43182,N_43024);
nand U43962 (N_43962,N_43480,N_43042);
nor U43963 (N_43963,N_43460,N_43466);
nand U43964 (N_43964,N_43293,N_43434);
xnor U43965 (N_43965,N_43013,N_43052);
xnor U43966 (N_43966,N_43406,N_43325);
nand U43967 (N_43967,N_43385,N_43292);
nor U43968 (N_43968,N_43166,N_43420);
or U43969 (N_43969,N_43499,N_43149);
xnor U43970 (N_43970,N_43484,N_43046);
nand U43971 (N_43971,N_43340,N_43093);
xnor U43972 (N_43972,N_43287,N_43202);
nand U43973 (N_43973,N_43079,N_43388);
nand U43974 (N_43974,N_43157,N_43426);
and U43975 (N_43975,N_43094,N_43176);
or U43976 (N_43976,N_43350,N_43352);
nor U43977 (N_43977,N_43060,N_43119);
or U43978 (N_43978,N_43452,N_43381);
nand U43979 (N_43979,N_43488,N_43415);
and U43980 (N_43980,N_43481,N_43390);
xor U43981 (N_43981,N_43210,N_43344);
and U43982 (N_43982,N_43215,N_43053);
xor U43983 (N_43983,N_43327,N_43283);
or U43984 (N_43984,N_43050,N_43151);
xnor U43985 (N_43985,N_43294,N_43476);
or U43986 (N_43986,N_43438,N_43063);
or U43987 (N_43987,N_43095,N_43486);
or U43988 (N_43988,N_43329,N_43281);
nor U43989 (N_43989,N_43106,N_43318);
xnor U43990 (N_43990,N_43008,N_43136);
nor U43991 (N_43991,N_43339,N_43198);
nand U43992 (N_43992,N_43383,N_43192);
xnor U43993 (N_43993,N_43288,N_43412);
nor U43994 (N_43994,N_43018,N_43436);
and U43995 (N_43995,N_43161,N_43176);
or U43996 (N_43996,N_43422,N_43309);
nand U43997 (N_43997,N_43426,N_43259);
nand U43998 (N_43998,N_43188,N_43105);
or U43999 (N_43999,N_43111,N_43440);
or U44000 (N_44000,N_43543,N_43584);
xor U44001 (N_44001,N_43740,N_43980);
nor U44002 (N_44002,N_43718,N_43847);
and U44003 (N_44003,N_43904,N_43744);
xor U44004 (N_44004,N_43547,N_43967);
and U44005 (N_44005,N_43992,N_43998);
or U44006 (N_44006,N_43800,N_43766);
and U44007 (N_44007,N_43600,N_43641);
nand U44008 (N_44008,N_43646,N_43738);
xor U44009 (N_44009,N_43822,N_43725);
nand U44010 (N_44010,N_43510,N_43556);
nand U44011 (N_44011,N_43686,N_43970);
and U44012 (N_44012,N_43661,N_43680);
or U44013 (N_44013,N_43908,N_43669);
xor U44014 (N_44014,N_43785,N_43577);
or U44015 (N_44015,N_43912,N_43879);
or U44016 (N_44016,N_43805,N_43806);
nor U44017 (N_44017,N_43569,N_43799);
and U44018 (N_44018,N_43512,N_43628);
or U44019 (N_44019,N_43719,N_43524);
or U44020 (N_44020,N_43553,N_43561);
xor U44021 (N_44021,N_43837,N_43918);
and U44022 (N_44022,N_43645,N_43868);
nand U44023 (N_44023,N_43968,N_43890);
or U44024 (N_44024,N_43615,N_43591);
nor U44025 (N_44025,N_43691,N_43504);
and U44026 (N_44026,N_43827,N_43567);
nor U44027 (N_44027,N_43851,N_43951);
nand U44028 (N_44028,N_43902,N_43530);
nand U44029 (N_44029,N_43969,N_43937);
nand U44030 (N_44030,N_43947,N_43729);
nand U44031 (N_44031,N_43949,N_43915);
or U44032 (N_44032,N_43579,N_43790);
xnor U44033 (N_44033,N_43724,N_43728);
or U44034 (N_44034,N_43565,N_43555);
nand U44035 (N_44035,N_43849,N_43931);
and U44036 (N_44036,N_43546,N_43863);
nand U44037 (N_44037,N_43812,N_43501);
nand U44038 (N_44038,N_43830,N_43679);
nand U44039 (N_44039,N_43707,N_43558);
or U44040 (N_44040,N_43559,N_43757);
nand U44041 (N_44041,N_43739,N_43630);
or U44042 (N_44042,N_43989,N_43824);
or U44043 (N_44043,N_43694,N_43907);
or U44044 (N_44044,N_43919,N_43913);
and U44045 (N_44045,N_43995,N_43791);
or U44046 (N_44046,N_43942,N_43898);
nor U44047 (N_44047,N_43823,N_43576);
or U44048 (N_44048,N_43516,N_43783);
and U44049 (N_44049,N_43666,N_43672);
and U44050 (N_44050,N_43870,N_43659);
xnor U44051 (N_44051,N_43722,N_43786);
or U44052 (N_44052,N_43844,N_43977);
xor U44053 (N_44053,N_43713,N_43706);
nand U44054 (N_44054,N_43663,N_43716);
or U44055 (N_44055,N_43900,N_43835);
nand U44056 (N_44056,N_43508,N_43749);
nor U44057 (N_44057,N_43873,N_43855);
nor U44058 (N_44058,N_43751,N_43613);
nand U44059 (N_44059,N_43647,N_43982);
nor U44060 (N_44060,N_43509,N_43711);
and U44061 (N_44061,N_43668,N_43518);
and U44062 (N_44062,N_43606,N_43853);
or U44063 (N_44063,N_43637,N_43523);
and U44064 (N_44064,N_43604,N_43650);
nand U44065 (N_44065,N_43564,N_43976);
or U44066 (N_44066,N_43587,N_43633);
nand U44067 (N_44067,N_43727,N_43658);
nor U44068 (N_44068,N_43638,N_43816);
xnor U44069 (N_44069,N_43676,N_43994);
and U44070 (N_44070,N_43896,N_43581);
and U44071 (N_44071,N_43959,N_43956);
nand U44072 (N_44072,N_43924,N_43934);
nand U44073 (N_44073,N_43511,N_43624);
nand U44074 (N_44074,N_43943,N_43532);
or U44075 (N_44075,N_43828,N_43945);
xor U44076 (N_44076,N_43921,N_43617);
and U44077 (N_44077,N_43939,N_43726);
nand U44078 (N_44078,N_43608,N_43585);
or U44079 (N_44079,N_43793,N_43926);
nand U44080 (N_44080,N_43609,N_43983);
nand U44081 (N_44081,N_43897,N_43520);
or U44082 (N_44082,N_43657,N_43958);
nand U44083 (N_44083,N_43748,N_43528);
nand U44084 (N_44084,N_43648,N_43986);
or U44085 (N_44085,N_43610,N_43871);
nand U44086 (N_44086,N_43704,N_43715);
nor U44087 (N_44087,N_43614,N_43723);
and U44088 (N_44088,N_43521,N_43737);
or U44089 (N_44089,N_43687,N_43597);
nor U44090 (N_44090,N_43573,N_43954);
and U44091 (N_44091,N_43771,N_43880);
xnor U44092 (N_44092,N_43901,N_43549);
xnor U44093 (N_44093,N_43764,N_43963);
nor U44094 (N_44094,N_43531,N_43538);
xnor U44095 (N_44095,N_43563,N_43731);
nor U44096 (N_44096,N_43964,N_43888);
xor U44097 (N_44097,N_43845,N_43631);
nor U44098 (N_44098,N_43857,N_43838);
nor U44099 (N_44099,N_43861,N_43622);
nor U44100 (N_44100,N_43712,N_43583);
nor U44101 (N_44101,N_43789,N_43673);
or U44102 (N_44102,N_43971,N_43536);
and U44103 (N_44103,N_43818,N_43920);
xor U44104 (N_44104,N_43655,N_43575);
or U44105 (N_44105,N_43519,N_43632);
xnor U44106 (N_44106,N_43957,N_43697);
nor U44107 (N_44107,N_43693,N_43801);
nor U44108 (N_44108,N_43804,N_43906);
nand U44109 (N_44109,N_43758,N_43649);
or U44110 (N_44110,N_43689,N_43526);
nand U44111 (N_44111,N_43955,N_43582);
and U44112 (N_44112,N_43787,N_43752);
or U44113 (N_44113,N_43962,N_43574);
xnor U44114 (N_44114,N_43802,N_43634);
nand U44115 (N_44115,N_43933,N_43590);
or U44116 (N_44116,N_43517,N_43952);
xor U44117 (N_44117,N_43929,N_43708);
or U44118 (N_44118,N_43506,N_43938);
or U44119 (N_44119,N_43843,N_43621);
or U44120 (N_44120,N_43775,N_43544);
xor U44121 (N_44121,N_43965,N_43776);
and U44122 (N_44122,N_43570,N_43683);
and U44123 (N_44123,N_43747,N_43651);
or U44124 (N_44124,N_43571,N_43960);
nor U44125 (N_44125,N_43560,N_43782);
nor U44126 (N_44126,N_43923,N_43753);
nand U44127 (N_44127,N_43742,N_43765);
nor U44128 (N_44128,N_43500,N_43627);
and U44129 (N_44129,N_43601,N_43656);
xor U44130 (N_44130,N_43777,N_43911);
xnor U44131 (N_44131,N_43554,N_43914);
xnor U44132 (N_44132,N_43732,N_43850);
or U44133 (N_44133,N_43932,N_43692);
or U44134 (N_44134,N_43681,N_43714);
xnor U44135 (N_44135,N_43829,N_43755);
nor U44136 (N_44136,N_43548,N_43674);
nor U44137 (N_44137,N_43767,N_43662);
and U44138 (N_44138,N_43936,N_43852);
or U44139 (N_44139,N_43808,N_43593);
nand U44140 (N_44140,N_43730,N_43644);
or U44141 (N_44141,N_43759,N_43842);
xnor U44142 (N_44142,N_43865,N_43545);
xnor U44143 (N_44143,N_43788,N_43568);
nand U44144 (N_44144,N_43618,N_43522);
nor U44145 (N_44145,N_43984,N_43503);
and U44146 (N_44146,N_43887,N_43595);
xnor U44147 (N_44147,N_43605,N_43763);
and U44148 (N_44148,N_43607,N_43925);
nor U44149 (N_44149,N_43684,N_43993);
nand U44150 (N_44150,N_43514,N_43572);
xor U44151 (N_44151,N_43889,N_43750);
nor U44152 (N_44152,N_43741,N_43746);
or U44153 (N_44153,N_43940,N_43710);
nor U44154 (N_44154,N_43602,N_43670);
or U44155 (N_44155,N_43917,N_43978);
or U44156 (N_44156,N_43598,N_43792);
or U44157 (N_44157,N_43988,N_43720);
xnor U44158 (N_44158,N_43909,N_43660);
or U44159 (N_44159,N_43831,N_43507);
nand U44160 (N_44160,N_43916,N_43635);
or U44161 (N_44161,N_43781,N_43770);
and U44162 (N_44162,N_43525,N_43690);
or U44163 (N_44163,N_43966,N_43769);
nor U44164 (N_44164,N_43623,N_43540);
nor U44165 (N_44165,N_43810,N_43675);
or U44166 (N_44166,N_43884,N_43819);
or U44167 (N_44167,N_43754,N_43619);
or U44168 (N_44168,N_43682,N_43784);
nor U44169 (N_44169,N_43580,N_43768);
and U44170 (N_44170,N_43639,N_43513);
or U44171 (N_44171,N_43814,N_43695);
xnor U44172 (N_44172,N_43973,N_43505);
nand U44173 (N_44173,N_43612,N_43780);
xnor U44174 (N_44174,N_43566,N_43859);
xor U44175 (N_44175,N_43987,N_43699);
or U44176 (N_44176,N_43653,N_43832);
xnor U44177 (N_44177,N_43717,N_43864);
xor U44178 (N_44178,N_43745,N_43841);
nand U44179 (N_44179,N_43778,N_43834);
and U44180 (N_44180,N_43603,N_43975);
nor U44181 (N_44181,N_43874,N_43935);
nor U44182 (N_44182,N_43700,N_43654);
xnor U44183 (N_44183,N_43885,N_43826);
nor U44184 (N_44184,N_43990,N_43541);
nor U44185 (N_44185,N_43698,N_43772);
or U44186 (N_44186,N_43535,N_43948);
and U44187 (N_44187,N_43667,N_43893);
or U44188 (N_44188,N_43981,N_43905);
nand U44189 (N_44189,N_43833,N_43922);
and U44190 (N_44190,N_43709,N_43736);
nor U44191 (N_44191,N_43652,N_43903);
or U44192 (N_44192,N_43869,N_43756);
and U44193 (N_44193,N_43537,N_43552);
xor U44194 (N_44194,N_43941,N_43991);
xor U44195 (N_44195,N_43856,N_43592);
nand U44196 (N_44196,N_43562,N_43815);
xor U44197 (N_44197,N_43910,N_43846);
nor U44198 (N_44198,N_43578,N_43773);
xnor U44199 (N_44199,N_43997,N_43734);
and U44200 (N_44200,N_43616,N_43701);
and U44201 (N_44201,N_43643,N_43671);
or U44202 (N_44202,N_43735,N_43599);
nor U44203 (N_44203,N_43928,N_43533);
xor U44204 (N_44204,N_43813,N_43854);
or U44205 (N_44205,N_43596,N_43797);
nand U44206 (N_44206,N_43803,N_43611);
and U44207 (N_44207,N_43867,N_43877);
nand U44208 (N_44208,N_43534,N_43858);
xor U44209 (N_44209,N_43860,N_43999);
and U44210 (N_44210,N_43825,N_43985);
or U44211 (N_44211,N_43620,N_43950);
nand U44212 (N_44212,N_43539,N_43809);
xnor U44213 (N_44213,N_43625,N_43953);
xor U44214 (N_44214,N_43703,N_43820);
xor U44215 (N_44215,N_43862,N_43642);
nor U44216 (N_44216,N_43840,N_43586);
or U44217 (N_44217,N_43702,N_43946);
and U44218 (N_44218,N_43761,N_43894);
and U44219 (N_44219,N_43721,N_43502);
nand U44220 (N_44220,N_43961,N_43836);
and U44221 (N_44221,N_43839,N_43878);
nand U44222 (N_44222,N_43762,N_43795);
and U44223 (N_44223,N_43875,N_43588);
xnor U44224 (N_44224,N_43883,N_43866);
xor U44225 (N_44225,N_43796,N_43743);
and U44226 (N_44226,N_43542,N_43677);
and U44227 (N_44227,N_43821,N_43705);
nand U44228 (N_44228,N_43892,N_43881);
or U44229 (N_44229,N_43848,N_43972);
or U44230 (N_44230,N_43589,N_43817);
nor U44231 (N_44231,N_43529,N_43944);
xnor U44232 (N_44232,N_43678,N_43640);
and U44233 (N_44233,N_43974,N_43774);
xnor U44234 (N_44234,N_43626,N_43760);
or U44235 (N_44235,N_43876,N_43515);
nor U44236 (N_44236,N_43551,N_43996);
xor U44237 (N_44237,N_43550,N_43688);
or U44238 (N_44238,N_43891,N_43527);
xor U44239 (N_44239,N_43665,N_43807);
or U44240 (N_44240,N_43733,N_43664);
or U44241 (N_44241,N_43557,N_43779);
and U44242 (N_44242,N_43685,N_43979);
nand U44243 (N_44243,N_43899,N_43927);
nand U44244 (N_44244,N_43594,N_43930);
nand U44245 (N_44245,N_43798,N_43882);
xor U44246 (N_44246,N_43811,N_43629);
xor U44247 (N_44247,N_43696,N_43636);
nor U44248 (N_44248,N_43895,N_43886);
and U44249 (N_44249,N_43872,N_43794);
nand U44250 (N_44250,N_43593,N_43911);
nor U44251 (N_44251,N_43749,N_43804);
nand U44252 (N_44252,N_43823,N_43844);
and U44253 (N_44253,N_43628,N_43669);
nand U44254 (N_44254,N_43679,N_43783);
or U44255 (N_44255,N_43786,N_43642);
nor U44256 (N_44256,N_43593,N_43769);
nor U44257 (N_44257,N_43860,N_43993);
xor U44258 (N_44258,N_43525,N_43853);
nor U44259 (N_44259,N_43505,N_43659);
nand U44260 (N_44260,N_43532,N_43886);
nand U44261 (N_44261,N_43911,N_43561);
or U44262 (N_44262,N_43755,N_43516);
and U44263 (N_44263,N_43952,N_43966);
and U44264 (N_44264,N_43503,N_43513);
nor U44265 (N_44265,N_43983,N_43657);
nand U44266 (N_44266,N_43833,N_43860);
and U44267 (N_44267,N_43733,N_43695);
or U44268 (N_44268,N_43976,N_43981);
or U44269 (N_44269,N_43782,N_43935);
and U44270 (N_44270,N_43870,N_43725);
nor U44271 (N_44271,N_43651,N_43770);
nor U44272 (N_44272,N_43595,N_43568);
or U44273 (N_44273,N_43734,N_43848);
nor U44274 (N_44274,N_43571,N_43679);
xor U44275 (N_44275,N_43536,N_43794);
xnor U44276 (N_44276,N_43550,N_43994);
or U44277 (N_44277,N_43818,N_43639);
and U44278 (N_44278,N_43707,N_43637);
nor U44279 (N_44279,N_43773,N_43571);
or U44280 (N_44280,N_43934,N_43982);
nor U44281 (N_44281,N_43545,N_43569);
xor U44282 (N_44282,N_43931,N_43547);
xor U44283 (N_44283,N_43844,N_43943);
nor U44284 (N_44284,N_43968,N_43600);
and U44285 (N_44285,N_43512,N_43732);
or U44286 (N_44286,N_43923,N_43787);
or U44287 (N_44287,N_43531,N_43823);
xor U44288 (N_44288,N_43972,N_43841);
and U44289 (N_44289,N_43539,N_43891);
and U44290 (N_44290,N_43709,N_43757);
nand U44291 (N_44291,N_43794,N_43700);
or U44292 (N_44292,N_43785,N_43700);
nor U44293 (N_44293,N_43570,N_43510);
or U44294 (N_44294,N_43597,N_43840);
nor U44295 (N_44295,N_43724,N_43571);
xor U44296 (N_44296,N_43656,N_43579);
nor U44297 (N_44297,N_43720,N_43511);
nand U44298 (N_44298,N_43635,N_43888);
and U44299 (N_44299,N_43735,N_43915);
and U44300 (N_44300,N_43572,N_43654);
nand U44301 (N_44301,N_43633,N_43993);
nand U44302 (N_44302,N_43523,N_43645);
nor U44303 (N_44303,N_43656,N_43536);
nand U44304 (N_44304,N_43643,N_43597);
and U44305 (N_44305,N_43620,N_43644);
and U44306 (N_44306,N_43717,N_43614);
nand U44307 (N_44307,N_43758,N_43898);
or U44308 (N_44308,N_43771,N_43838);
xnor U44309 (N_44309,N_43534,N_43648);
and U44310 (N_44310,N_43937,N_43979);
nor U44311 (N_44311,N_43957,N_43670);
nor U44312 (N_44312,N_43596,N_43825);
and U44313 (N_44313,N_43571,N_43725);
xor U44314 (N_44314,N_43999,N_43521);
nand U44315 (N_44315,N_43527,N_43673);
xnor U44316 (N_44316,N_43592,N_43722);
nor U44317 (N_44317,N_43517,N_43566);
nand U44318 (N_44318,N_43522,N_43667);
and U44319 (N_44319,N_43854,N_43670);
nand U44320 (N_44320,N_43610,N_43819);
and U44321 (N_44321,N_43814,N_43662);
nor U44322 (N_44322,N_43790,N_43539);
xor U44323 (N_44323,N_43591,N_43803);
xor U44324 (N_44324,N_43661,N_43735);
xor U44325 (N_44325,N_43822,N_43529);
xnor U44326 (N_44326,N_43513,N_43875);
nor U44327 (N_44327,N_43540,N_43530);
xor U44328 (N_44328,N_43810,N_43717);
nor U44329 (N_44329,N_43761,N_43775);
and U44330 (N_44330,N_43909,N_43911);
and U44331 (N_44331,N_43601,N_43884);
nor U44332 (N_44332,N_43919,N_43731);
nand U44333 (N_44333,N_43793,N_43735);
and U44334 (N_44334,N_43585,N_43544);
nand U44335 (N_44335,N_43973,N_43672);
and U44336 (N_44336,N_43575,N_43914);
xnor U44337 (N_44337,N_43592,N_43738);
xor U44338 (N_44338,N_43918,N_43924);
nand U44339 (N_44339,N_43640,N_43833);
or U44340 (N_44340,N_43736,N_43808);
or U44341 (N_44341,N_43986,N_43806);
and U44342 (N_44342,N_43963,N_43702);
nand U44343 (N_44343,N_43981,N_43952);
xnor U44344 (N_44344,N_43635,N_43691);
nand U44345 (N_44345,N_43645,N_43549);
and U44346 (N_44346,N_43633,N_43845);
or U44347 (N_44347,N_43918,N_43693);
nor U44348 (N_44348,N_43626,N_43759);
xnor U44349 (N_44349,N_43691,N_43725);
xor U44350 (N_44350,N_43851,N_43749);
xor U44351 (N_44351,N_43810,N_43975);
or U44352 (N_44352,N_43616,N_43633);
nor U44353 (N_44353,N_43574,N_43759);
xor U44354 (N_44354,N_43752,N_43701);
xor U44355 (N_44355,N_43557,N_43897);
or U44356 (N_44356,N_43894,N_43731);
nand U44357 (N_44357,N_43970,N_43761);
and U44358 (N_44358,N_43618,N_43552);
or U44359 (N_44359,N_43994,N_43693);
and U44360 (N_44360,N_43601,N_43959);
and U44361 (N_44361,N_43635,N_43580);
and U44362 (N_44362,N_43634,N_43971);
xnor U44363 (N_44363,N_43556,N_43891);
and U44364 (N_44364,N_43603,N_43923);
nand U44365 (N_44365,N_43845,N_43793);
xnor U44366 (N_44366,N_43781,N_43971);
xor U44367 (N_44367,N_43746,N_43929);
and U44368 (N_44368,N_43855,N_43627);
nand U44369 (N_44369,N_43998,N_43879);
nor U44370 (N_44370,N_43961,N_43707);
or U44371 (N_44371,N_43946,N_43822);
or U44372 (N_44372,N_43894,N_43561);
nor U44373 (N_44373,N_43660,N_43525);
nand U44374 (N_44374,N_43820,N_43984);
and U44375 (N_44375,N_43524,N_43852);
nor U44376 (N_44376,N_43672,N_43560);
and U44377 (N_44377,N_43795,N_43600);
nor U44378 (N_44378,N_43689,N_43597);
xnor U44379 (N_44379,N_43900,N_43808);
or U44380 (N_44380,N_43729,N_43778);
nand U44381 (N_44381,N_43742,N_43670);
nor U44382 (N_44382,N_43504,N_43922);
and U44383 (N_44383,N_43877,N_43691);
or U44384 (N_44384,N_43943,N_43909);
nand U44385 (N_44385,N_43693,N_43666);
xnor U44386 (N_44386,N_43753,N_43959);
xnor U44387 (N_44387,N_43793,N_43537);
or U44388 (N_44388,N_43780,N_43847);
and U44389 (N_44389,N_43896,N_43946);
or U44390 (N_44390,N_43704,N_43573);
nor U44391 (N_44391,N_43516,N_43644);
nand U44392 (N_44392,N_43915,N_43580);
nand U44393 (N_44393,N_43700,N_43603);
nor U44394 (N_44394,N_43550,N_43788);
and U44395 (N_44395,N_43789,N_43526);
nor U44396 (N_44396,N_43893,N_43743);
nand U44397 (N_44397,N_43784,N_43576);
xor U44398 (N_44398,N_43652,N_43633);
xor U44399 (N_44399,N_43606,N_43797);
xor U44400 (N_44400,N_43552,N_43976);
nor U44401 (N_44401,N_43805,N_43775);
and U44402 (N_44402,N_43950,N_43703);
nor U44403 (N_44403,N_43551,N_43853);
and U44404 (N_44404,N_43685,N_43918);
or U44405 (N_44405,N_43803,N_43792);
nor U44406 (N_44406,N_43958,N_43515);
nor U44407 (N_44407,N_43821,N_43602);
xnor U44408 (N_44408,N_43833,N_43834);
and U44409 (N_44409,N_43831,N_43971);
or U44410 (N_44410,N_43771,N_43953);
or U44411 (N_44411,N_43558,N_43564);
nor U44412 (N_44412,N_43908,N_43555);
nand U44413 (N_44413,N_43803,N_43837);
and U44414 (N_44414,N_43920,N_43575);
nor U44415 (N_44415,N_43633,N_43775);
or U44416 (N_44416,N_43726,N_43870);
xor U44417 (N_44417,N_43655,N_43750);
and U44418 (N_44418,N_43932,N_43700);
or U44419 (N_44419,N_43775,N_43742);
nand U44420 (N_44420,N_43620,N_43566);
nor U44421 (N_44421,N_43878,N_43815);
nor U44422 (N_44422,N_43902,N_43698);
nor U44423 (N_44423,N_43926,N_43614);
and U44424 (N_44424,N_43906,N_43560);
and U44425 (N_44425,N_43563,N_43681);
nor U44426 (N_44426,N_43709,N_43669);
or U44427 (N_44427,N_43632,N_43777);
and U44428 (N_44428,N_43937,N_43551);
nor U44429 (N_44429,N_43947,N_43546);
nand U44430 (N_44430,N_43785,N_43999);
nand U44431 (N_44431,N_43576,N_43711);
and U44432 (N_44432,N_43896,N_43691);
nor U44433 (N_44433,N_43890,N_43616);
and U44434 (N_44434,N_43830,N_43547);
nor U44435 (N_44435,N_43503,N_43771);
or U44436 (N_44436,N_43948,N_43812);
nand U44437 (N_44437,N_43904,N_43501);
nor U44438 (N_44438,N_43830,N_43667);
nor U44439 (N_44439,N_43845,N_43682);
and U44440 (N_44440,N_43777,N_43631);
nand U44441 (N_44441,N_43541,N_43811);
nor U44442 (N_44442,N_43786,N_43948);
and U44443 (N_44443,N_43953,N_43658);
nand U44444 (N_44444,N_43517,N_43645);
or U44445 (N_44445,N_43591,N_43951);
or U44446 (N_44446,N_43946,N_43933);
or U44447 (N_44447,N_43873,N_43813);
nand U44448 (N_44448,N_43833,N_43575);
nor U44449 (N_44449,N_43917,N_43938);
xor U44450 (N_44450,N_43857,N_43581);
xor U44451 (N_44451,N_43875,N_43696);
and U44452 (N_44452,N_43946,N_43528);
and U44453 (N_44453,N_43673,N_43593);
and U44454 (N_44454,N_43688,N_43656);
nor U44455 (N_44455,N_43886,N_43848);
and U44456 (N_44456,N_43941,N_43547);
nor U44457 (N_44457,N_43889,N_43859);
and U44458 (N_44458,N_43626,N_43624);
nor U44459 (N_44459,N_43941,N_43661);
and U44460 (N_44460,N_43969,N_43611);
and U44461 (N_44461,N_43769,N_43561);
or U44462 (N_44462,N_43643,N_43961);
nor U44463 (N_44463,N_43680,N_43969);
nor U44464 (N_44464,N_43870,N_43583);
xor U44465 (N_44465,N_43566,N_43534);
or U44466 (N_44466,N_43781,N_43866);
or U44467 (N_44467,N_43788,N_43737);
and U44468 (N_44468,N_43875,N_43624);
xnor U44469 (N_44469,N_43548,N_43860);
or U44470 (N_44470,N_43669,N_43847);
or U44471 (N_44471,N_43940,N_43781);
or U44472 (N_44472,N_43632,N_43977);
and U44473 (N_44473,N_43724,N_43623);
or U44474 (N_44474,N_43691,N_43700);
or U44475 (N_44475,N_43941,N_43829);
nand U44476 (N_44476,N_43684,N_43581);
nor U44477 (N_44477,N_43618,N_43899);
or U44478 (N_44478,N_43632,N_43654);
and U44479 (N_44479,N_43799,N_43639);
and U44480 (N_44480,N_43548,N_43636);
xnor U44481 (N_44481,N_43791,N_43993);
nor U44482 (N_44482,N_43517,N_43902);
or U44483 (N_44483,N_43953,N_43687);
and U44484 (N_44484,N_43723,N_43573);
xor U44485 (N_44485,N_43640,N_43862);
or U44486 (N_44486,N_43841,N_43836);
and U44487 (N_44487,N_43547,N_43887);
and U44488 (N_44488,N_43823,N_43910);
nand U44489 (N_44489,N_43878,N_43523);
and U44490 (N_44490,N_43558,N_43511);
and U44491 (N_44491,N_43935,N_43736);
or U44492 (N_44492,N_43770,N_43850);
nand U44493 (N_44493,N_43836,N_43604);
nand U44494 (N_44494,N_43901,N_43590);
nor U44495 (N_44495,N_43675,N_43771);
nand U44496 (N_44496,N_43803,N_43698);
or U44497 (N_44497,N_43873,N_43749);
nor U44498 (N_44498,N_43969,N_43608);
and U44499 (N_44499,N_43706,N_43750);
xnor U44500 (N_44500,N_44218,N_44141);
xnor U44501 (N_44501,N_44213,N_44015);
nand U44502 (N_44502,N_44112,N_44028);
xor U44503 (N_44503,N_44014,N_44421);
or U44504 (N_44504,N_44365,N_44043);
xor U44505 (N_44505,N_44388,N_44228);
nor U44506 (N_44506,N_44072,N_44019);
nor U44507 (N_44507,N_44401,N_44198);
nor U44508 (N_44508,N_44430,N_44338);
and U44509 (N_44509,N_44428,N_44268);
xnor U44510 (N_44510,N_44064,N_44270);
xnor U44511 (N_44511,N_44358,N_44169);
nor U44512 (N_44512,N_44295,N_44332);
or U44513 (N_44513,N_44390,N_44315);
xor U44514 (N_44514,N_44306,N_44487);
xnor U44515 (N_44515,N_44140,N_44386);
nand U44516 (N_44516,N_44088,N_44345);
and U44517 (N_44517,N_44127,N_44216);
xnor U44518 (N_44518,N_44320,N_44102);
or U44519 (N_44519,N_44284,N_44298);
xnor U44520 (N_44520,N_44468,N_44057);
and U44521 (N_44521,N_44287,N_44172);
xor U44522 (N_44522,N_44147,N_44134);
or U44523 (N_44523,N_44469,N_44079);
nand U44524 (N_44524,N_44137,N_44318);
nor U44525 (N_44525,N_44477,N_44067);
nand U44526 (N_44526,N_44203,N_44050);
nor U44527 (N_44527,N_44403,N_44340);
and U44528 (N_44528,N_44397,N_44008);
and U44529 (N_44529,N_44209,N_44272);
nor U44530 (N_44530,N_44256,N_44275);
xor U44531 (N_44531,N_44223,N_44308);
nand U44532 (N_44532,N_44266,N_44289);
or U44533 (N_44533,N_44179,N_44461);
nand U44534 (N_44534,N_44262,N_44382);
nand U44535 (N_44535,N_44493,N_44370);
or U44536 (N_44536,N_44394,N_44431);
and U44537 (N_44537,N_44291,N_44490);
xnor U44538 (N_44538,N_44475,N_44448);
or U44539 (N_44539,N_44126,N_44138);
and U44540 (N_44540,N_44080,N_44085);
nor U44541 (N_44541,N_44035,N_44076);
nor U44542 (N_44542,N_44485,N_44410);
nand U44543 (N_44543,N_44491,N_44247);
and U44544 (N_44544,N_44447,N_44139);
xnor U44545 (N_44545,N_44457,N_44023);
nor U44546 (N_44546,N_44093,N_44440);
nand U44547 (N_44547,N_44154,N_44416);
xnor U44548 (N_44548,N_44177,N_44250);
nor U44549 (N_44549,N_44368,N_44413);
and U44550 (N_44550,N_44217,N_44344);
and U44551 (N_44551,N_44305,N_44105);
nor U44552 (N_44552,N_44162,N_44068);
or U44553 (N_44553,N_44279,N_44124);
xor U44554 (N_44554,N_44060,N_44337);
xor U44555 (N_44555,N_44010,N_44161);
nor U44556 (N_44556,N_44013,N_44155);
nor U44557 (N_44557,N_44463,N_44438);
nand U44558 (N_44558,N_44481,N_44464);
and U44559 (N_44559,N_44460,N_44148);
nor U44560 (N_44560,N_44012,N_44374);
and U44561 (N_44561,N_44201,N_44474);
nor U44562 (N_44562,N_44237,N_44196);
or U44563 (N_44563,N_44273,N_44423);
and U44564 (N_44564,N_44024,N_44492);
xor U44565 (N_44565,N_44480,N_44353);
or U44566 (N_44566,N_44054,N_44163);
and U44567 (N_44567,N_44205,N_44167);
nand U44568 (N_44568,N_44441,N_44281);
nor U44569 (N_44569,N_44354,N_44407);
and U44570 (N_44570,N_44009,N_44197);
xnor U44571 (N_44571,N_44233,N_44007);
and U44572 (N_44572,N_44135,N_44395);
and U44573 (N_44573,N_44181,N_44389);
nand U44574 (N_44574,N_44096,N_44283);
xnor U44575 (N_44575,N_44107,N_44255);
or U44576 (N_44576,N_44360,N_44212);
or U44577 (N_44577,N_44158,N_44065);
and U44578 (N_44578,N_44082,N_44331);
xor U44579 (N_44579,N_44323,N_44357);
and U44580 (N_44580,N_44059,N_44210);
and U44581 (N_44581,N_44325,N_44222);
or U44582 (N_44582,N_44031,N_44446);
or U44583 (N_44583,N_44378,N_44249);
xnor U44584 (N_44584,N_44176,N_44120);
and U44585 (N_44585,N_44104,N_44097);
and U44586 (N_44586,N_44478,N_44373);
xnor U44587 (N_44587,N_44499,N_44494);
nor U44588 (N_44588,N_44253,N_44336);
and U44589 (N_44589,N_44341,N_44351);
nor U44590 (N_44590,N_44225,N_44027);
nand U44591 (N_44591,N_44226,N_44412);
or U44592 (N_44592,N_44496,N_44380);
and U44593 (N_44593,N_44215,N_44355);
nor U44594 (N_44594,N_44221,N_44118);
nor U44595 (N_44595,N_44425,N_44280);
nand U44596 (N_44596,N_44405,N_44489);
and U44597 (N_44597,N_44311,N_44452);
nand U44598 (N_44598,N_44251,N_44192);
nand U44599 (N_44599,N_44239,N_44302);
xor U44600 (N_44600,N_44087,N_44070);
and U44601 (N_44601,N_44058,N_44396);
xnor U44602 (N_44602,N_44333,N_44170);
and U44603 (N_44603,N_44453,N_44185);
nor U44604 (N_44604,N_44399,N_44178);
nor U44605 (N_44605,N_44269,N_44300);
nor U44606 (N_44606,N_44330,N_44435);
nand U44607 (N_44607,N_44328,N_44375);
nand U44608 (N_44608,N_44352,N_44146);
and U44609 (N_44609,N_44114,N_44377);
nor U44610 (N_44610,N_44202,N_44117);
or U44611 (N_44611,N_44108,N_44470);
or U44612 (N_44612,N_44227,N_44404);
and U44613 (N_44613,N_44439,N_44149);
xnor U44614 (N_44614,N_44159,N_44191);
nand U44615 (N_44615,N_44437,N_44037);
nand U44616 (N_44616,N_44398,N_44483);
and U44617 (N_44617,N_44263,N_44303);
nor U44618 (N_44618,N_44495,N_44246);
or U44619 (N_44619,N_44030,N_44032);
nand U44620 (N_44620,N_44219,N_44041);
xnor U44621 (N_44621,N_44426,N_44466);
nand U44622 (N_44622,N_44186,N_44433);
nand U44623 (N_44623,N_44415,N_44095);
nand U44624 (N_44624,N_44376,N_44123);
nor U44625 (N_44625,N_44274,N_44366);
and U44626 (N_44626,N_44290,N_44075);
and U44627 (N_44627,N_44436,N_44317);
nor U44628 (N_44628,N_44304,N_44450);
nand U44629 (N_44629,N_44276,N_44301);
or U44630 (N_44630,N_44116,N_44271);
nand U44631 (N_44631,N_44265,N_44455);
nand U44632 (N_44632,N_44039,N_44346);
xnor U44633 (N_44633,N_44168,N_44156);
nand U44634 (N_44634,N_44409,N_44051);
xnor U44635 (N_44635,N_44004,N_44111);
and U44636 (N_44636,N_44190,N_44005);
nor U44637 (N_44637,N_44073,N_44106);
nand U44638 (N_44638,N_44100,N_44220);
nor U44639 (N_44639,N_44094,N_44310);
nor U44640 (N_44640,N_44362,N_44131);
xnor U44641 (N_44641,N_44391,N_44419);
xnor U44642 (N_44642,N_44422,N_44349);
xnor U44643 (N_44643,N_44165,N_44125);
nand U44644 (N_44644,N_44115,N_44018);
nor U44645 (N_44645,N_44078,N_44194);
nand U44646 (N_44646,N_44254,N_44160);
nand U44647 (N_44647,N_44136,N_44069);
nand U44648 (N_44648,N_44327,N_44016);
or U44649 (N_44649,N_44025,N_44129);
and U44650 (N_44650,N_44314,N_44350);
or U44651 (N_44651,N_44242,N_44456);
nor U44652 (N_44652,N_44400,N_44183);
or U44653 (N_44653,N_44372,N_44454);
xor U44654 (N_44654,N_44184,N_44252);
nor U44655 (N_44655,N_44406,N_44150);
nor U44656 (N_44656,N_44451,N_44240);
xnor U44657 (N_44657,N_44498,N_44049);
or U44658 (N_44658,N_44066,N_44449);
xor U44659 (N_44659,N_44040,N_44445);
nand U44660 (N_44660,N_44145,N_44195);
nand U44661 (N_44661,N_44429,N_44420);
and U44662 (N_44662,N_44359,N_44214);
xor U44663 (N_44663,N_44189,N_44047);
or U44664 (N_44664,N_44241,N_44443);
nand U44665 (N_44665,N_44393,N_44022);
xnor U44666 (N_44666,N_44482,N_44174);
nor U44667 (N_44667,N_44387,N_44379);
xnor U44668 (N_44668,N_44371,N_44099);
and U44669 (N_44669,N_44312,N_44038);
xor U44670 (N_44670,N_44121,N_44128);
and U44671 (N_44671,N_44224,N_44044);
and U44672 (N_44672,N_44036,N_44098);
and U44673 (N_44673,N_44232,N_44153);
or U44674 (N_44674,N_44144,N_44414);
and U44675 (N_44675,N_44091,N_44130);
and U44676 (N_44676,N_44236,N_44322);
nor U44677 (N_44677,N_44363,N_44321);
or U44678 (N_44678,N_44029,N_44048);
and U44679 (N_44679,N_44294,N_44385);
xor U44680 (N_44680,N_44292,N_44077);
nand U44681 (N_44681,N_44465,N_44101);
nor U44682 (N_44682,N_44171,N_44180);
or U44683 (N_44683,N_44459,N_44484);
xnor U44684 (N_44684,N_44342,N_44417);
and U44685 (N_44685,N_44293,N_44335);
nor U44686 (N_44686,N_44248,N_44257);
xor U44687 (N_44687,N_44316,N_44231);
nor U44688 (N_44688,N_44367,N_44151);
or U44689 (N_44689,N_44261,N_44084);
xor U44690 (N_44690,N_44000,N_44187);
or U44691 (N_44691,N_44488,N_44486);
or U44692 (N_44692,N_44017,N_44244);
or U44693 (N_44693,N_44444,N_44199);
or U44694 (N_44694,N_44381,N_44297);
and U44695 (N_44695,N_44133,N_44383);
nand U44696 (N_44696,N_44074,N_44055);
nor U44697 (N_44697,N_44083,N_44235);
nor U44698 (N_44698,N_44001,N_44157);
and U44699 (N_44699,N_44056,N_44434);
nand U44700 (N_44700,N_44245,N_44045);
xor U44701 (N_44701,N_44206,N_44286);
or U44702 (N_44702,N_44424,N_44277);
xnor U44703 (N_44703,N_44173,N_44230);
nor U44704 (N_44704,N_44238,N_44208);
nand U44705 (N_44705,N_44063,N_44473);
and U44706 (N_44706,N_44334,N_44418);
or U44707 (N_44707,N_44207,N_44109);
and U44708 (N_44708,N_44119,N_44392);
nand U44709 (N_44709,N_44061,N_44260);
xor U44710 (N_44710,N_44166,N_44442);
or U44711 (N_44711,N_44113,N_44329);
or U44712 (N_44712,N_44188,N_44313);
xor U44713 (N_44713,N_44200,N_44021);
nand U44714 (N_44714,N_44006,N_44081);
and U44715 (N_44715,N_44467,N_44347);
nor U44716 (N_44716,N_44364,N_44071);
nand U44717 (N_44717,N_44259,N_44296);
and U44718 (N_44718,N_44476,N_44062);
xnor U44719 (N_44719,N_44267,N_44324);
nor U44720 (N_44720,N_44132,N_44011);
or U44721 (N_44721,N_44033,N_44110);
or U44722 (N_44722,N_44408,N_44307);
and U44723 (N_44723,N_44046,N_44026);
nor U44724 (N_44724,N_44402,N_44278);
and U44725 (N_44725,N_44182,N_44002);
nand U44726 (N_44726,N_44384,N_44427);
nor U44727 (N_44727,N_44348,N_44299);
or U44728 (N_44728,N_44472,N_44339);
xor U44729 (N_44729,N_44258,N_44411);
or U44730 (N_44730,N_44211,N_44471);
xnor U44731 (N_44731,N_44264,N_44243);
nand U44732 (N_44732,N_44122,N_44175);
nand U44733 (N_44733,N_44479,N_44052);
xnor U44734 (N_44734,N_44020,N_44432);
nand U44735 (N_44735,N_44143,N_44086);
or U44736 (N_44736,N_44042,N_44053);
nor U44737 (N_44737,N_44089,N_44369);
or U44738 (N_44738,N_44356,N_44034);
xnor U44739 (N_44739,N_44497,N_44458);
nor U44740 (N_44740,N_44164,N_44103);
nor U44741 (N_44741,N_44092,N_44319);
and U44742 (N_44742,N_44285,N_44142);
nor U44743 (N_44743,N_44361,N_44234);
xor U44744 (N_44744,N_44090,N_44288);
and U44745 (N_44745,N_44152,N_44309);
and U44746 (N_44746,N_44326,N_44343);
xnor U44747 (N_44747,N_44462,N_44003);
or U44748 (N_44748,N_44282,N_44204);
nor U44749 (N_44749,N_44193,N_44229);
xor U44750 (N_44750,N_44079,N_44453);
xor U44751 (N_44751,N_44452,N_44494);
xor U44752 (N_44752,N_44239,N_44042);
nand U44753 (N_44753,N_44254,N_44300);
and U44754 (N_44754,N_44319,N_44239);
or U44755 (N_44755,N_44339,N_44191);
or U44756 (N_44756,N_44136,N_44375);
or U44757 (N_44757,N_44193,N_44358);
nor U44758 (N_44758,N_44382,N_44446);
nor U44759 (N_44759,N_44128,N_44161);
nor U44760 (N_44760,N_44364,N_44094);
nand U44761 (N_44761,N_44351,N_44066);
and U44762 (N_44762,N_44138,N_44179);
xnor U44763 (N_44763,N_44439,N_44233);
and U44764 (N_44764,N_44004,N_44441);
nor U44765 (N_44765,N_44347,N_44005);
and U44766 (N_44766,N_44317,N_44053);
xnor U44767 (N_44767,N_44286,N_44137);
xnor U44768 (N_44768,N_44409,N_44344);
and U44769 (N_44769,N_44294,N_44108);
nand U44770 (N_44770,N_44101,N_44373);
and U44771 (N_44771,N_44472,N_44004);
nor U44772 (N_44772,N_44423,N_44432);
xnor U44773 (N_44773,N_44276,N_44141);
nand U44774 (N_44774,N_44460,N_44007);
and U44775 (N_44775,N_44311,N_44137);
nand U44776 (N_44776,N_44122,N_44005);
and U44777 (N_44777,N_44250,N_44350);
nand U44778 (N_44778,N_44106,N_44441);
and U44779 (N_44779,N_44403,N_44006);
or U44780 (N_44780,N_44479,N_44210);
nor U44781 (N_44781,N_44295,N_44216);
and U44782 (N_44782,N_44248,N_44343);
xor U44783 (N_44783,N_44071,N_44007);
or U44784 (N_44784,N_44023,N_44318);
xor U44785 (N_44785,N_44434,N_44090);
nand U44786 (N_44786,N_44369,N_44251);
or U44787 (N_44787,N_44372,N_44102);
nand U44788 (N_44788,N_44242,N_44019);
nor U44789 (N_44789,N_44118,N_44044);
or U44790 (N_44790,N_44367,N_44093);
xor U44791 (N_44791,N_44072,N_44148);
nor U44792 (N_44792,N_44234,N_44099);
or U44793 (N_44793,N_44161,N_44364);
nand U44794 (N_44794,N_44082,N_44371);
nor U44795 (N_44795,N_44400,N_44202);
nand U44796 (N_44796,N_44399,N_44219);
or U44797 (N_44797,N_44070,N_44264);
xnor U44798 (N_44798,N_44494,N_44090);
nor U44799 (N_44799,N_44319,N_44457);
nand U44800 (N_44800,N_44301,N_44458);
nor U44801 (N_44801,N_44267,N_44223);
nor U44802 (N_44802,N_44441,N_44467);
nor U44803 (N_44803,N_44330,N_44390);
and U44804 (N_44804,N_44432,N_44244);
nor U44805 (N_44805,N_44484,N_44491);
or U44806 (N_44806,N_44474,N_44252);
xor U44807 (N_44807,N_44272,N_44268);
and U44808 (N_44808,N_44478,N_44227);
nor U44809 (N_44809,N_44380,N_44136);
nor U44810 (N_44810,N_44143,N_44127);
nand U44811 (N_44811,N_44338,N_44154);
and U44812 (N_44812,N_44336,N_44095);
and U44813 (N_44813,N_44372,N_44032);
and U44814 (N_44814,N_44453,N_44050);
xor U44815 (N_44815,N_44368,N_44141);
nor U44816 (N_44816,N_44217,N_44225);
xnor U44817 (N_44817,N_44025,N_44078);
nand U44818 (N_44818,N_44064,N_44326);
or U44819 (N_44819,N_44299,N_44489);
nor U44820 (N_44820,N_44250,N_44006);
nor U44821 (N_44821,N_44180,N_44177);
xor U44822 (N_44822,N_44095,N_44412);
nor U44823 (N_44823,N_44432,N_44088);
or U44824 (N_44824,N_44262,N_44210);
nand U44825 (N_44825,N_44427,N_44166);
xor U44826 (N_44826,N_44267,N_44212);
or U44827 (N_44827,N_44069,N_44164);
and U44828 (N_44828,N_44203,N_44005);
nor U44829 (N_44829,N_44264,N_44411);
nand U44830 (N_44830,N_44447,N_44210);
and U44831 (N_44831,N_44478,N_44347);
nor U44832 (N_44832,N_44037,N_44094);
xor U44833 (N_44833,N_44461,N_44404);
and U44834 (N_44834,N_44082,N_44165);
or U44835 (N_44835,N_44161,N_44463);
xor U44836 (N_44836,N_44478,N_44447);
or U44837 (N_44837,N_44153,N_44070);
and U44838 (N_44838,N_44113,N_44466);
nand U44839 (N_44839,N_44053,N_44293);
nor U44840 (N_44840,N_44438,N_44394);
or U44841 (N_44841,N_44122,N_44462);
or U44842 (N_44842,N_44048,N_44145);
xor U44843 (N_44843,N_44241,N_44340);
and U44844 (N_44844,N_44099,N_44463);
nor U44845 (N_44845,N_44275,N_44013);
and U44846 (N_44846,N_44132,N_44160);
xnor U44847 (N_44847,N_44337,N_44260);
nand U44848 (N_44848,N_44489,N_44414);
or U44849 (N_44849,N_44300,N_44166);
xor U44850 (N_44850,N_44048,N_44259);
nor U44851 (N_44851,N_44401,N_44365);
nand U44852 (N_44852,N_44423,N_44177);
or U44853 (N_44853,N_44222,N_44149);
nand U44854 (N_44854,N_44417,N_44105);
or U44855 (N_44855,N_44133,N_44304);
and U44856 (N_44856,N_44138,N_44248);
and U44857 (N_44857,N_44440,N_44049);
and U44858 (N_44858,N_44339,N_44141);
or U44859 (N_44859,N_44431,N_44206);
nor U44860 (N_44860,N_44109,N_44316);
and U44861 (N_44861,N_44051,N_44435);
nor U44862 (N_44862,N_44458,N_44352);
nor U44863 (N_44863,N_44109,N_44383);
nand U44864 (N_44864,N_44330,N_44008);
nand U44865 (N_44865,N_44427,N_44080);
or U44866 (N_44866,N_44203,N_44166);
xnor U44867 (N_44867,N_44349,N_44182);
and U44868 (N_44868,N_44141,N_44033);
and U44869 (N_44869,N_44261,N_44445);
or U44870 (N_44870,N_44439,N_44454);
xnor U44871 (N_44871,N_44386,N_44121);
nand U44872 (N_44872,N_44249,N_44294);
nand U44873 (N_44873,N_44105,N_44390);
xor U44874 (N_44874,N_44008,N_44425);
and U44875 (N_44875,N_44287,N_44389);
or U44876 (N_44876,N_44329,N_44193);
and U44877 (N_44877,N_44342,N_44459);
xnor U44878 (N_44878,N_44169,N_44401);
nor U44879 (N_44879,N_44297,N_44333);
and U44880 (N_44880,N_44464,N_44340);
and U44881 (N_44881,N_44178,N_44494);
xnor U44882 (N_44882,N_44158,N_44450);
xor U44883 (N_44883,N_44075,N_44169);
and U44884 (N_44884,N_44312,N_44146);
nand U44885 (N_44885,N_44377,N_44166);
or U44886 (N_44886,N_44496,N_44063);
or U44887 (N_44887,N_44003,N_44057);
xor U44888 (N_44888,N_44389,N_44113);
nor U44889 (N_44889,N_44353,N_44205);
nand U44890 (N_44890,N_44279,N_44016);
and U44891 (N_44891,N_44112,N_44189);
or U44892 (N_44892,N_44236,N_44073);
nor U44893 (N_44893,N_44460,N_44311);
xnor U44894 (N_44894,N_44185,N_44233);
and U44895 (N_44895,N_44213,N_44365);
xnor U44896 (N_44896,N_44479,N_44089);
nand U44897 (N_44897,N_44157,N_44151);
and U44898 (N_44898,N_44259,N_44004);
nand U44899 (N_44899,N_44469,N_44321);
nor U44900 (N_44900,N_44435,N_44013);
xnor U44901 (N_44901,N_44030,N_44361);
and U44902 (N_44902,N_44050,N_44499);
nor U44903 (N_44903,N_44475,N_44152);
nor U44904 (N_44904,N_44063,N_44374);
xor U44905 (N_44905,N_44368,N_44279);
nor U44906 (N_44906,N_44295,N_44006);
nor U44907 (N_44907,N_44230,N_44239);
nor U44908 (N_44908,N_44188,N_44281);
and U44909 (N_44909,N_44046,N_44280);
xor U44910 (N_44910,N_44153,N_44401);
nand U44911 (N_44911,N_44034,N_44471);
nand U44912 (N_44912,N_44399,N_44377);
nor U44913 (N_44913,N_44136,N_44097);
nand U44914 (N_44914,N_44026,N_44258);
nand U44915 (N_44915,N_44092,N_44229);
xnor U44916 (N_44916,N_44328,N_44446);
or U44917 (N_44917,N_44283,N_44393);
or U44918 (N_44918,N_44230,N_44127);
nand U44919 (N_44919,N_44051,N_44335);
nor U44920 (N_44920,N_44260,N_44080);
nor U44921 (N_44921,N_44296,N_44117);
and U44922 (N_44922,N_44003,N_44291);
nand U44923 (N_44923,N_44485,N_44248);
nand U44924 (N_44924,N_44274,N_44320);
or U44925 (N_44925,N_44023,N_44491);
and U44926 (N_44926,N_44496,N_44003);
xnor U44927 (N_44927,N_44088,N_44119);
nand U44928 (N_44928,N_44160,N_44289);
and U44929 (N_44929,N_44015,N_44236);
xnor U44930 (N_44930,N_44341,N_44148);
xor U44931 (N_44931,N_44324,N_44109);
nand U44932 (N_44932,N_44216,N_44039);
nor U44933 (N_44933,N_44473,N_44071);
and U44934 (N_44934,N_44224,N_44230);
xnor U44935 (N_44935,N_44369,N_44423);
nor U44936 (N_44936,N_44423,N_44165);
or U44937 (N_44937,N_44057,N_44404);
nand U44938 (N_44938,N_44373,N_44076);
or U44939 (N_44939,N_44192,N_44033);
nor U44940 (N_44940,N_44416,N_44480);
and U44941 (N_44941,N_44358,N_44399);
nor U44942 (N_44942,N_44474,N_44321);
or U44943 (N_44943,N_44420,N_44196);
nand U44944 (N_44944,N_44258,N_44260);
and U44945 (N_44945,N_44242,N_44099);
nand U44946 (N_44946,N_44412,N_44172);
xnor U44947 (N_44947,N_44313,N_44193);
xnor U44948 (N_44948,N_44329,N_44357);
and U44949 (N_44949,N_44457,N_44020);
nand U44950 (N_44950,N_44388,N_44301);
nand U44951 (N_44951,N_44435,N_44212);
xnor U44952 (N_44952,N_44112,N_44313);
nor U44953 (N_44953,N_44112,N_44294);
or U44954 (N_44954,N_44485,N_44107);
nand U44955 (N_44955,N_44425,N_44015);
xor U44956 (N_44956,N_44011,N_44351);
nand U44957 (N_44957,N_44412,N_44169);
and U44958 (N_44958,N_44427,N_44390);
nor U44959 (N_44959,N_44121,N_44145);
and U44960 (N_44960,N_44321,N_44344);
nor U44961 (N_44961,N_44249,N_44248);
nand U44962 (N_44962,N_44061,N_44186);
nor U44963 (N_44963,N_44437,N_44143);
or U44964 (N_44964,N_44014,N_44220);
and U44965 (N_44965,N_44469,N_44043);
nand U44966 (N_44966,N_44307,N_44058);
or U44967 (N_44967,N_44056,N_44493);
nor U44968 (N_44968,N_44396,N_44171);
nor U44969 (N_44969,N_44346,N_44049);
nand U44970 (N_44970,N_44377,N_44458);
and U44971 (N_44971,N_44332,N_44229);
or U44972 (N_44972,N_44241,N_44360);
nand U44973 (N_44973,N_44254,N_44241);
nand U44974 (N_44974,N_44173,N_44433);
nand U44975 (N_44975,N_44436,N_44351);
xnor U44976 (N_44976,N_44360,N_44041);
and U44977 (N_44977,N_44444,N_44260);
or U44978 (N_44978,N_44250,N_44356);
xor U44979 (N_44979,N_44315,N_44349);
or U44980 (N_44980,N_44411,N_44465);
or U44981 (N_44981,N_44150,N_44230);
nand U44982 (N_44982,N_44096,N_44336);
nand U44983 (N_44983,N_44054,N_44086);
or U44984 (N_44984,N_44179,N_44354);
or U44985 (N_44985,N_44256,N_44222);
xor U44986 (N_44986,N_44020,N_44081);
nor U44987 (N_44987,N_44240,N_44219);
nor U44988 (N_44988,N_44463,N_44247);
xor U44989 (N_44989,N_44472,N_44306);
nand U44990 (N_44990,N_44169,N_44327);
nand U44991 (N_44991,N_44208,N_44361);
nor U44992 (N_44992,N_44412,N_44332);
xor U44993 (N_44993,N_44078,N_44408);
xnor U44994 (N_44994,N_44253,N_44332);
xor U44995 (N_44995,N_44157,N_44131);
xnor U44996 (N_44996,N_44267,N_44244);
xnor U44997 (N_44997,N_44169,N_44457);
and U44998 (N_44998,N_44256,N_44267);
and U44999 (N_44999,N_44276,N_44143);
or U45000 (N_45000,N_44893,N_44956);
or U45001 (N_45001,N_44900,N_44527);
nand U45002 (N_45002,N_44688,N_44886);
nor U45003 (N_45003,N_44866,N_44834);
xor U45004 (N_45004,N_44521,N_44560);
nor U45005 (N_45005,N_44986,N_44518);
and U45006 (N_45006,N_44717,N_44915);
nor U45007 (N_45007,N_44975,N_44620);
xor U45008 (N_45008,N_44860,N_44971);
nand U45009 (N_45009,N_44730,N_44988);
and U45010 (N_45010,N_44757,N_44574);
and U45011 (N_45011,N_44762,N_44695);
xnor U45012 (N_45012,N_44919,N_44796);
nand U45013 (N_45013,N_44949,N_44644);
nor U45014 (N_45014,N_44947,N_44830);
nor U45015 (N_45015,N_44957,N_44610);
nor U45016 (N_45016,N_44711,N_44908);
xnor U45017 (N_45017,N_44787,N_44655);
nor U45018 (N_45018,N_44780,N_44768);
nand U45019 (N_45019,N_44827,N_44510);
and U45020 (N_45020,N_44870,N_44748);
nand U45021 (N_45021,N_44671,N_44928);
nor U45022 (N_45022,N_44775,N_44739);
xnor U45023 (N_45023,N_44989,N_44679);
nor U45024 (N_45024,N_44643,N_44592);
xnor U45025 (N_45025,N_44641,N_44579);
or U45026 (N_45026,N_44666,N_44639);
xor U45027 (N_45027,N_44516,N_44501);
and U45028 (N_45028,N_44794,N_44985);
xnor U45029 (N_45029,N_44788,N_44702);
nor U45030 (N_45030,N_44898,N_44998);
xor U45031 (N_45031,N_44615,N_44699);
nand U45032 (N_45032,N_44868,N_44664);
or U45033 (N_45033,N_44909,N_44759);
or U45034 (N_45034,N_44647,N_44704);
nand U45035 (N_45035,N_44724,N_44809);
or U45036 (N_45036,N_44933,N_44853);
or U45037 (N_45037,N_44546,N_44571);
and U45038 (N_45038,N_44715,N_44941);
or U45039 (N_45039,N_44551,N_44686);
or U45040 (N_45040,N_44554,N_44541);
and U45041 (N_45041,N_44912,N_44667);
and U45042 (N_45042,N_44525,N_44875);
or U45043 (N_45043,N_44774,N_44595);
nand U45044 (N_45044,N_44879,N_44509);
xnor U45045 (N_45045,N_44980,N_44994);
nor U45046 (N_45046,N_44614,N_44533);
nor U45047 (N_45047,N_44669,N_44732);
nor U45048 (N_45048,N_44718,N_44802);
and U45049 (N_45049,N_44857,N_44531);
and U45050 (N_45050,N_44995,N_44631);
xor U45051 (N_45051,N_44935,N_44781);
nand U45052 (N_45052,N_44992,N_44741);
xnor U45053 (N_45053,N_44656,N_44712);
nand U45054 (N_45054,N_44619,N_44654);
and U45055 (N_45055,N_44921,N_44874);
nand U45056 (N_45056,N_44856,N_44734);
nand U45057 (N_45057,N_44709,N_44826);
or U45058 (N_45058,N_44676,N_44943);
and U45059 (N_45059,N_44895,N_44858);
nand U45060 (N_45060,N_44700,N_44897);
nand U45061 (N_45061,N_44969,N_44645);
or U45062 (N_45062,N_44884,N_44630);
xor U45063 (N_45063,N_44637,N_44653);
nand U45064 (N_45064,N_44539,N_44810);
nor U45065 (N_45065,N_44596,N_44511);
and U45066 (N_45066,N_44790,N_44569);
and U45067 (N_45067,N_44763,N_44814);
and U45068 (N_45068,N_44825,N_44607);
nand U45069 (N_45069,N_44609,N_44508);
xor U45070 (N_45070,N_44881,N_44566);
nand U45071 (N_45071,N_44681,N_44634);
and U45072 (N_45072,N_44758,N_44638);
nor U45073 (N_45073,N_44589,N_44737);
nor U45074 (N_45074,N_44795,N_44515);
nor U45075 (N_45075,N_44804,N_44512);
nand U45076 (N_45076,N_44976,N_44618);
nand U45077 (N_45077,N_44694,N_44911);
xnor U45078 (N_45078,N_44564,N_44864);
or U45079 (N_45079,N_44824,N_44940);
xnor U45080 (N_45080,N_44880,N_44602);
or U45081 (N_45081,N_44851,N_44685);
nor U45082 (N_45082,N_44613,N_44678);
and U45083 (N_45083,N_44764,N_44954);
nand U45084 (N_45084,N_44575,N_44913);
and U45085 (N_45085,N_44823,N_44828);
and U45086 (N_45086,N_44628,N_44966);
nand U45087 (N_45087,N_44777,N_44651);
or U45088 (N_45088,N_44728,N_44996);
and U45089 (N_45089,N_44968,N_44953);
nor U45090 (N_45090,N_44783,N_44663);
and U45091 (N_45091,N_44740,N_44529);
or U45092 (N_45092,N_44659,N_44594);
or U45093 (N_45093,N_44835,N_44997);
nor U45094 (N_45094,N_44677,N_44576);
nor U45095 (N_45095,N_44934,N_44812);
or U45096 (N_45096,N_44500,N_44627);
nand U45097 (N_45097,N_44789,N_44929);
and U45098 (N_45098,N_44549,N_44692);
or U45099 (N_45099,N_44832,N_44682);
nand U45100 (N_45100,N_44885,N_44977);
nand U45101 (N_45101,N_44670,N_44859);
xor U45102 (N_45102,N_44738,N_44605);
nand U45103 (N_45103,N_44865,N_44993);
or U45104 (N_45104,N_44693,N_44749);
xnor U45105 (N_45105,N_44601,N_44747);
nor U45106 (N_45106,N_44842,N_44567);
or U45107 (N_45107,N_44733,N_44506);
or U45108 (N_45108,N_44782,N_44930);
xnor U45109 (N_45109,N_44640,N_44914);
and U45110 (N_45110,N_44582,N_44650);
nand U45111 (N_45111,N_44672,N_44815);
or U45112 (N_45112,N_44552,N_44766);
and U45113 (N_45113,N_44562,N_44565);
nor U45114 (N_45114,N_44652,N_44863);
and U45115 (N_45115,N_44608,N_44550);
and U45116 (N_45116,N_44598,N_44513);
or U45117 (N_45117,N_44517,N_44773);
nor U45118 (N_45118,N_44904,N_44593);
nand U45119 (N_45119,N_44855,N_44603);
nand U45120 (N_45120,N_44792,N_44999);
or U45121 (N_45121,N_44807,N_44636);
nand U45122 (N_45122,N_44642,N_44751);
or U45123 (N_45123,N_44535,N_44877);
nand U45124 (N_45124,N_44945,N_44987);
nand U45125 (N_45125,N_44534,N_44816);
and U45126 (N_45126,N_44833,N_44697);
xnor U45127 (N_45127,N_44726,N_44746);
or U45128 (N_45128,N_44557,N_44960);
and U45129 (N_45129,N_44952,N_44545);
xnor U45130 (N_45130,N_44570,N_44955);
xnor U45131 (N_45131,N_44854,N_44963);
nor U45132 (N_45132,N_44590,N_44979);
nand U45133 (N_45133,N_44982,N_44710);
nand U45134 (N_45134,N_44990,N_44573);
xor U45135 (N_45135,N_44745,N_44821);
nor U45136 (N_45136,N_44536,N_44936);
nor U45137 (N_45137,N_44519,N_44735);
xor U45138 (N_45138,N_44705,N_44800);
and U45139 (N_45139,N_44837,N_44767);
nand U45140 (N_45140,N_44831,N_44840);
or U45141 (N_45141,N_44714,N_44938);
nor U45142 (N_45142,N_44632,N_44958);
nand U45143 (N_45143,N_44896,N_44923);
or U45144 (N_45144,N_44970,N_44984);
xnor U45145 (N_45145,N_44731,N_44578);
or U45146 (N_45146,N_44927,N_44950);
nor U45147 (N_45147,N_44588,N_44648);
and U45148 (N_45148,N_44756,N_44625);
nand U45149 (N_45149,N_44532,N_44665);
and U45150 (N_45150,N_44743,N_44873);
xor U45151 (N_45151,N_44503,N_44587);
xnor U45152 (N_45152,N_44722,N_44701);
or U45153 (N_45153,N_44887,N_44811);
nand U45154 (N_45154,N_44577,N_44600);
xnor U45155 (N_45155,N_44937,N_44661);
nand U45156 (N_45156,N_44612,N_44523);
or U45157 (N_45157,N_44611,N_44597);
and U45158 (N_45158,N_44752,N_44528);
nor U45159 (N_45159,N_44843,N_44755);
and U45160 (N_45160,N_44524,N_44680);
nand U45161 (N_45161,N_44961,N_44635);
or U45162 (N_45162,N_44925,N_44948);
and U45163 (N_45163,N_44836,N_44683);
and U45164 (N_45164,N_44778,N_44848);
nor U45165 (N_45165,N_44606,N_44706);
nand U45166 (N_45166,N_44698,N_44585);
nand U45167 (N_45167,N_44959,N_44708);
nor U45168 (N_45168,N_44725,N_44829);
and U45169 (N_45169,N_44617,N_44844);
nor U45170 (N_45170,N_44805,N_44526);
and U45171 (N_45171,N_44537,N_44504);
or U45172 (N_45172,N_44727,N_44553);
or U45173 (N_45173,N_44901,N_44750);
or U45174 (N_45174,N_44852,N_44522);
nor U45175 (N_45175,N_44916,N_44703);
nand U45176 (N_45176,N_44798,N_44931);
nor U45177 (N_45177,N_44662,N_44902);
nand U45178 (N_45178,N_44818,N_44894);
and U45179 (N_45179,N_44801,N_44910);
nand U45180 (N_45180,N_44660,N_44540);
or U45181 (N_45181,N_44820,N_44753);
nand U45182 (N_45182,N_44696,N_44806);
nor U45183 (N_45183,N_44784,N_44719);
xnor U45184 (N_45184,N_44538,N_44861);
nor U45185 (N_45185,N_44922,N_44555);
nand U45186 (N_45186,N_44530,N_44920);
nor U45187 (N_45187,N_44689,N_44964);
xor U45188 (N_45188,N_44721,N_44559);
or U45189 (N_45189,N_44769,N_44657);
or U45190 (N_45190,N_44974,N_44972);
nor U45191 (N_45191,N_44978,N_44899);
or U45192 (N_45192,N_44568,N_44808);
xor U45193 (N_45193,N_44736,N_44547);
xnor U45194 (N_45194,N_44505,N_44983);
xnor U45195 (N_45195,N_44819,N_44707);
nor U45196 (N_45196,N_44556,N_44723);
nor U45197 (N_45197,N_44907,N_44799);
and U45198 (N_45198,N_44867,N_44507);
nor U45199 (N_45199,N_44583,N_44646);
nor U45200 (N_45200,N_44889,N_44621);
nor U45201 (N_45201,N_44862,N_44542);
xnor U45202 (N_45202,N_44845,N_44770);
nand U45203 (N_45203,N_44572,N_44888);
and U45204 (N_45204,N_44761,N_44744);
nor U45205 (N_45205,N_44797,N_44754);
and U45206 (N_45206,N_44918,N_44876);
nand U45207 (N_45207,N_44684,N_44586);
nor U45208 (N_45208,N_44942,N_44839);
or U45209 (N_45209,N_44944,N_44793);
or U45210 (N_45210,N_44924,N_44558);
nor U45211 (N_45211,N_44991,N_44878);
or U45212 (N_45212,N_44838,N_44520);
nor U45213 (N_45213,N_44981,N_44917);
nor U45214 (N_45214,N_44591,N_44813);
or U45215 (N_45215,N_44563,N_44720);
nand U45216 (N_45216,N_44883,N_44502);
or U45217 (N_45217,N_44687,N_44849);
xnor U45218 (N_45218,N_44713,N_44890);
nor U45219 (N_45219,N_44729,N_44846);
nand U45220 (N_45220,N_44742,N_44906);
and U45221 (N_45221,N_44882,N_44599);
or U45222 (N_45222,N_44892,N_44548);
or U45223 (N_45223,N_44649,N_44847);
nor U45224 (N_45224,N_44765,N_44624);
or U45225 (N_45225,N_44771,N_44674);
or U45226 (N_45226,N_44932,N_44622);
and U45227 (N_45227,N_44658,N_44872);
and U45228 (N_45228,N_44965,N_44772);
nor U45229 (N_45229,N_44785,N_44668);
xnor U45230 (N_45230,N_44544,N_44779);
or U45231 (N_45231,N_44891,N_44791);
or U45232 (N_45232,N_44629,N_44850);
xnor U45233 (N_45233,N_44973,N_44716);
nand U45234 (N_45234,N_44673,N_44903);
or U45235 (N_45235,N_44946,N_44817);
and U45236 (N_45236,N_44633,N_44951);
nor U45237 (N_45237,N_44561,N_44776);
nor U45238 (N_45238,N_44760,N_44967);
nand U45239 (N_45239,N_44926,N_44786);
and U45240 (N_45240,N_44803,N_44869);
xor U45241 (N_45241,N_44514,N_44675);
or U45242 (N_45242,N_44626,N_44841);
and U45243 (N_45243,N_44871,N_44691);
nand U45244 (N_45244,N_44616,N_44905);
nand U45245 (N_45245,N_44822,N_44584);
xor U45246 (N_45246,N_44543,N_44604);
xnor U45247 (N_45247,N_44580,N_44939);
nand U45248 (N_45248,N_44581,N_44690);
nor U45249 (N_45249,N_44962,N_44623);
and U45250 (N_45250,N_44789,N_44792);
or U45251 (N_45251,N_44805,N_44860);
nand U45252 (N_45252,N_44696,N_44867);
nand U45253 (N_45253,N_44993,N_44661);
and U45254 (N_45254,N_44901,N_44951);
nand U45255 (N_45255,N_44604,N_44788);
xnor U45256 (N_45256,N_44973,N_44783);
nor U45257 (N_45257,N_44984,N_44977);
or U45258 (N_45258,N_44693,N_44828);
or U45259 (N_45259,N_44722,N_44925);
and U45260 (N_45260,N_44605,N_44973);
nor U45261 (N_45261,N_44519,N_44650);
and U45262 (N_45262,N_44982,N_44751);
nor U45263 (N_45263,N_44873,N_44889);
or U45264 (N_45264,N_44788,N_44934);
xor U45265 (N_45265,N_44830,N_44523);
nor U45266 (N_45266,N_44749,N_44598);
xor U45267 (N_45267,N_44747,N_44941);
or U45268 (N_45268,N_44924,N_44787);
and U45269 (N_45269,N_44959,N_44733);
or U45270 (N_45270,N_44798,N_44812);
nand U45271 (N_45271,N_44867,N_44998);
nor U45272 (N_45272,N_44861,N_44571);
nor U45273 (N_45273,N_44952,N_44883);
xnor U45274 (N_45274,N_44501,N_44849);
xor U45275 (N_45275,N_44957,N_44766);
nand U45276 (N_45276,N_44846,N_44898);
xnor U45277 (N_45277,N_44660,N_44587);
or U45278 (N_45278,N_44761,N_44525);
or U45279 (N_45279,N_44791,N_44763);
nor U45280 (N_45280,N_44704,N_44927);
or U45281 (N_45281,N_44898,N_44723);
xor U45282 (N_45282,N_44543,N_44821);
nor U45283 (N_45283,N_44883,N_44949);
or U45284 (N_45284,N_44753,N_44576);
nor U45285 (N_45285,N_44831,N_44635);
nand U45286 (N_45286,N_44705,N_44684);
and U45287 (N_45287,N_44645,N_44802);
or U45288 (N_45288,N_44937,N_44725);
and U45289 (N_45289,N_44662,N_44713);
and U45290 (N_45290,N_44663,N_44996);
and U45291 (N_45291,N_44648,N_44886);
or U45292 (N_45292,N_44965,N_44741);
and U45293 (N_45293,N_44955,N_44782);
nor U45294 (N_45294,N_44684,N_44776);
xnor U45295 (N_45295,N_44758,N_44516);
nand U45296 (N_45296,N_44937,N_44573);
or U45297 (N_45297,N_44780,N_44711);
xor U45298 (N_45298,N_44508,N_44977);
nand U45299 (N_45299,N_44558,N_44989);
nand U45300 (N_45300,N_44981,N_44677);
nand U45301 (N_45301,N_44931,N_44989);
nand U45302 (N_45302,N_44603,N_44549);
and U45303 (N_45303,N_44550,N_44680);
xor U45304 (N_45304,N_44867,N_44685);
nand U45305 (N_45305,N_44566,N_44545);
or U45306 (N_45306,N_44606,N_44689);
or U45307 (N_45307,N_44911,N_44804);
nor U45308 (N_45308,N_44883,N_44648);
xor U45309 (N_45309,N_44804,N_44992);
and U45310 (N_45310,N_44702,N_44564);
xor U45311 (N_45311,N_44798,N_44851);
xor U45312 (N_45312,N_44793,N_44542);
xor U45313 (N_45313,N_44840,N_44924);
nor U45314 (N_45314,N_44936,N_44960);
xnor U45315 (N_45315,N_44781,N_44807);
nand U45316 (N_45316,N_44566,N_44964);
or U45317 (N_45317,N_44508,N_44944);
nor U45318 (N_45318,N_44815,N_44547);
nand U45319 (N_45319,N_44764,N_44702);
nand U45320 (N_45320,N_44733,N_44935);
or U45321 (N_45321,N_44990,N_44641);
nor U45322 (N_45322,N_44702,N_44913);
nor U45323 (N_45323,N_44880,N_44663);
and U45324 (N_45324,N_44595,N_44650);
nor U45325 (N_45325,N_44643,N_44903);
nor U45326 (N_45326,N_44997,N_44858);
or U45327 (N_45327,N_44792,N_44827);
xnor U45328 (N_45328,N_44938,N_44890);
xnor U45329 (N_45329,N_44669,N_44529);
and U45330 (N_45330,N_44706,N_44829);
and U45331 (N_45331,N_44811,N_44842);
nand U45332 (N_45332,N_44525,N_44962);
nand U45333 (N_45333,N_44918,N_44732);
xor U45334 (N_45334,N_44568,N_44873);
and U45335 (N_45335,N_44593,N_44791);
or U45336 (N_45336,N_44768,N_44586);
nor U45337 (N_45337,N_44760,N_44657);
xnor U45338 (N_45338,N_44539,N_44875);
nand U45339 (N_45339,N_44712,N_44676);
or U45340 (N_45340,N_44585,N_44633);
nand U45341 (N_45341,N_44521,N_44976);
xnor U45342 (N_45342,N_44844,N_44894);
and U45343 (N_45343,N_44913,N_44708);
xnor U45344 (N_45344,N_44783,N_44986);
and U45345 (N_45345,N_44667,N_44553);
nor U45346 (N_45346,N_44787,N_44898);
and U45347 (N_45347,N_44654,N_44589);
xnor U45348 (N_45348,N_44776,N_44537);
or U45349 (N_45349,N_44666,N_44952);
and U45350 (N_45350,N_44515,N_44566);
nand U45351 (N_45351,N_44611,N_44956);
nor U45352 (N_45352,N_44886,N_44635);
and U45353 (N_45353,N_44549,N_44919);
or U45354 (N_45354,N_44532,N_44564);
nor U45355 (N_45355,N_44501,N_44883);
xor U45356 (N_45356,N_44515,N_44695);
or U45357 (N_45357,N_44605,N_44502);
or U45358 (N_45358,N_44826,N_44811);
nor U45359 (N_45359,N_44895,N_44850);
nand U45360 (N_45360,N_44531,N_44509);
nor U45361 (N_45361,N_44650,N_44843);
nand U45362 (N_45362,N_44736,N_44577);
xnor U45363 (N_45363,N_44845,N_44674);
and U45364 (N_45364,N_44708,N_44836);
xor U45365 (N_45365,N_44549,N_44749);
or U45366 (N_45366,N_44764,N_44815);
nor U45367 (N_45367,N_44912,N_44687);
nand U45368 (N_45368,N_44948,N_44520);
and U45369 (N_45369,N_44953,N_44680);
nor U45370 (N_45370,N_44522,N_44849);
and U45371 (N_45371,N_44910,N_44664);
xor U45372 (N_45372,N_44990,N_44968);
xor U45373 (N_45373,N_44677,N_44911);
xor U45374 (N_45374,N_44732,N_44653);
or U45375 (N_45375,N_44589,N_44977);
or U45376 (N_45376,N_44593,N_44866);
xnor U45377 (N_45377,N_44782,N_44594);
or U45378 (N_45378,N_44656,N_44658);
nand U45379 (N_45379,N_44794,N_44543);
or U45380 (N_45380,N_44855,N_44770);
or U45381 (N_45381,N_44983,N_44742);
or U45382 (N_45382,N_44692,N_44884);
nor U45383 (N_45383,N_44943,N_44995);
nand U45384 (N_45384,N_44828,N_44537);
nor U45385 (N_45385,N_44861,N_44791);
nand U45386 (N_45386,N_44698,N_44539);
nand U45387 (N_45387,N_44694,N_44840);
or U45388 (N_45388,N_44852,N_44815);
or U45389 (N_45389,N_44884,N_44880);
and U45390 (N_45390,N_44636,N_44672);
and U45391 (N_45391,N_44787,N_44789);
xnor U45392 (N_45392,N_44707,N_44751);
and U45393 (N_45393,N_44688,N_44818);
or U45394 (N_45394,N_44842,N_44776);
xor U45395 (N_45395,N_44510,N_44511);
or U45396 (N_45396,N_44954,N_44861);
nor U45397 (N_45397,N_44966,N_44598);
and U45398 (N_45398,N_44742,N_44818);
or U45399 (N_45399,N_44872,N_44827);
or U45400 (N_45400,N_44674,N_44659);
nand U45401 (N_45401,N_44833,N_44901);
or U45402 (N_45402,N_44504,N_44930);
xnor U45403 (N_45403,N_44848,N_44791);
or U45404 (N_45404,N_44613,N_44764);
nand U45405 (N_45405,N_44767,N_44567);
nor U45406 (N_45406,N_44546,N_44577);
and U45407 (N_45407,N_44723,N_44637);
and U45408 (N_45408,N_44992,N_44625);
or U45409 (N_45409,N_44774,N_44633);
and U45410 (N_45410,N_44611,N_44607);
nand U45411 (N_45411,N_44593,N_44967);
and U45412 (N_45412,N_44649,N_44980);
nor U45413 (N_45413,N_44999,N_44778);
or U45414 (N_45414,N_44832,N_44601);
xnor U45415 (N_45415,N_44854,N_44856);
nor U45416 (N_45416,N_44996,N_44924);
or U45417 (N_45417,N_44904,N_44573);
and U45418 (N_45418,N_44688,N_44992);
xnor U45419 (N_45419,N_44530,N_44899);
or U45420 (N_45420,N_44867,N_44900);
nor U45421 (N_45421,N_44781,N_44682);
and U45422 (N_45422,N_44801,N_44670);
and U45423 (N_45423,N_44979,N_44839);
xnor U45424 (N_45424,N_44580,N_44752);
xor U45425 (N_45425,N_44984,N_44825);
nand U45426 (N_45426,N_44527,N_44747);
nand U45427 (N_45427,N_44965,N_44617);
and U45428 (N_45428,N_44833,N_44505);
nand U45429 (N_45429,N_44943,N_44812);
and U45430 (N_45430,N_44669,N_44931);
xnor U45431 (N_45431,N_44870,N_44624);
or U45432 (N_45432,N_44625,N_44708);
xor U45433 (N_45433,N_44793,N_44538);
or U45434 (N_45434,N_44839,N_44728);
or U45435 (N_45435,N_44682,N_44744);
and U45436 (N_45436,N_44756,N_44982);
nand U45437 (N_45437,N_44600,N_44722);
or U45438 (N_45438,N_44933,N_44953);
and U45439 (N_45439,N_44789,N_44960);
and U45440 (N_45440,N_44693,N_44926);
nand U45441 (N_45441,N_44894,N_44644);
and U45442 (N_45442,N_44762,N_44881);
or U45443 (N_45443,N_44914,N_44523);
and U45444 (N_45444,N_44841,N_44501);
xor U45445 (N_45445,N_44825,N_44723);
xor U45446 (N_45446,N_44913,N_44994);
and U45447 (N_45447,N_44576,N_44956);
xor U45448 (N_45448,N_44741,N_44979);
nor U45449 (N_45449,N_44547,N_44708);
nand U45450 (N_45450,N_44688,N_44752);
xor U45451 (N_45451,N_44759,N_44620);
or U45452 (N_45452,N_44583,N_44642);
nor U45453 (N_45453,N_44972,N_44955);
xnor U45454 (N_45454,N_44538,N_44852);
nor U45455 (N_45455,N_44939,N_44534);
nor U45456 (N_45456,N_44937,N_44985);
nor U45457 (N_45457,N_44689,N_44935);
nand U45458 (N_45458,N_44595,N_44574);
and U45459 (N_45459,N_44723,N_44783);
nand U45460 (N_45460,N_44987,N_44697);
or U45461 (N_45461,N_44987,N_44760);
nand U45462 (N_45462,N_44939,N_44984);
or U45463 (N_45463,N_44756,N_44520);
or U45464 (N_45464,N_44702,N_44910);
xor U45465 (N_45465,N_44617,N_44652);
or U45466 (N_45466,N_44851,N_44546);
or U45467 (N_45467,N_44760,N_44897);
or U45468 (N_45468,N_44789,N_44645);
or U45469 (N_45469,N_44615,N_44835);
nor U45470 (N_45470,N_44554,N_44794);
nand U45471 (N_45471,N_44577,N_44879);
nor U45472 (N_45472,N_44859,N_44939);
nand U45473 (N_45473,N_44554,N_44622);
and U45474 (N_45474,N_44623,N_44580);
nand U45475 (N_45475,N_44508,N_44638);
or U45476 (N_45476,N_44986,N_44929);
nand U45477 (N_45477,N_44843,N_44740);
nand U45478 (N_45478,N_44533,N_44793);
nand U45479 (N_45479,N_44525,N_44717);
nand U45480 (N_45480,N_44597,N_44971);
nand U45481 (N_45481,N_44848,N_44929);
or U45482 (N_45482,N_44535,N_44946);
or U45483 (N_45483,N_44703,N_44968);
nand U45484 (N_45484,N_44871,N_44558);
nor U45485 (N_45485,N_44764,N_44709);
xor U45486 (N_45486,N_44623,N_44537);
xnor U45487 (N_45487,N_44631,N_44507);
and U45488 (N_45488,N_44588,N_44995);
or U45489 (N_45489,N_44983,N_44916);
or U45490 (N_45490,N_44574,N_44840);
or U45491 (N_45491,N_44941,N_44899);
xor U45492 (N_45492,N_44964,N_44584);
xor U45493 (N_45493,N_44785,N_44724);
xor U45494 (N_45494,N_44933,N_44751);
nor U45495 (N_45495,N_44543,N_44882);
nor U45496 (N_45496,N_44776,N_44615);
nand U45497 (N_45497,N_44795,N_44630);
nand U45498 (N_45498,N_44619,N_44973);
nand U45499 (N_45499,N_44831,N_44998);
xnor U45500 (N_45500,N_45458,N_45329);
nor U45501 (N_45501,N_45229,N_45260);
and U45502 (N_45502,N_45222,N_45184);
or U45503 (N_45503,N_45336,N_45287);
or U45504 (N_45504,N_45461,N_45266);
xor U45505 (N_45505,N_45049,N_45367);
nor U45506 (N_45506,N_45245,N_45435);
or U45507 (N_45507,N_45206,N_45077);
and U45508 (N_45508,N_45160,N_45491);
or U45509 (N_45509,N_45182,N_45442);
and U45510 (N_45510,N_45110,N_45129);
nand U45511 (N_45511,N_45490,N_45489);
nor U45512 (N_45512,N_45333,N_45072);
nand U45513 (N_45513,N_45263,N_45045);
or U45514 (N_45514,N_45488,N_45412);
nor U45515 (N_45515,N_45004,N_45403);
and U45516 (N_45516,N_45348,N_45462);
and U45517 (N_45517,N_45324,N_45423);
and U45518 (N_45518,N_45478,N_45471);
xnor U45519 (N_45519,N_45092,N_45413);
nor U45520 (N_45520,N_45362,N_45002);
nand U45521 (N_45521,N_45031,N_45425);
nor U45522 (N_45522,N_45296,N_45047);
nand U45523 (N_45523,N_45464,N_45411);
and U45524 (N_45524,N_45181,N_45390);
nand U45525 (N_45525,N_45215,N_45019);
nand U45526 (N_45526,N_45056,N_45289);
or U45527 (N_45527,N_45032,N_45434);
or U45528 (N_45528,N_45060,N_45451);
xor U45529 (N_45529,N_45247,N_45108);
and U45530 (N_45530,N_45431,N_45179);
nor U45531 (N_45531,N_45386,N_45028);
nor U45532 (N_45532,N_45109,N_45205);
nor U45533 (N_45533,N_45354,N_45283);
nand U45534 (N_45534,N_45365,N_45428);
and U45535 (N_45535,N_45363,N_45375);
nand U45536 (N_45536,N_45382,N_45204);
xor U45537 (N_45537,N_45409,N_45497);
nand U45538 (N_45538,N_45143,N_45420);
nand U45539 (N_45539,N_45317,N_45339);
or U45540 (N_45540,N_45437,N_45255);
and U45541 (N_45541,N_45378,N_45054);
xor U45542 (N_45542,N_45356,N_45188);
xor U45543 (N_45543,N_45278,N_45327);
xnor U45544 (N_45544,N_45029,N_45249);
nor U45545 (N_45545,N_45114,N_45292);
or U45546 (N_45546,N_45262,N_45430);
or U45547 (N_45547,N_45122,N_45210);
nand U45548 (N_45548,N_45083,N_45025);
xnor U45549 (N_45549,N_45001,N_45162);
xnor U45550 (N_45550,N_45294,N_45233);
and U45551 (N_45551,N_45472,N_45086);
nand U45552 (N_45552,N_45419,N_45172);
or U45553 (N_45553,N_45057,N_45117);
xnor U45554 (N_45554,N_45357,N_45220);
or U45555 (N_45555,N_45351,N_45223);
nor U45556 (N_45556,N_45246,N_45218);
or U45557 (N_45557,N_45325,N_45044);
or U45558 (N_45558,N_45498,N_45052);
or U45559 (N_45559,N_45318,N_45141);
and U45560 (N_45560,N_45163,N_45147);
nor U45561 (N_45561,N_45370,N_45020);
and U45562 (N_45562,N_45364,N_45446);
xor U45563 (N_45563,N_45165,N_45041);
and U45564 (N_45564,N_45368,N_45250);
and U45565 (N_45565,N_45225,N_45048);
xnor U45566 (N_45566,N_45046,N_45008);
or U45567 (N_45567,N_45011,N_45353);
nor U45568 (N_45568,N_45265,N_45142);
xnor U45569 (N_45569,N_45416,N_45268);
and U45570 (N_45570,N_45064,N_45207);
nor U45571 (N_45571,N_45078,N_45105);
and U45572 (N_45572,N_45331,N_45447);
xnor U45573 (N_45573,N_45426,N_45274);
and U45574 (N_45574,N_45422,N_45256);
nor U45575 (N_45575,N_45201,N_45404);
nor U45576 (N_45576,N_45460,N_45280);
xor U45577 (N_45577,N_45071,N_45017);
nand U45578 (N_45578,N_45113,N_45007);
or U45579 (N_45579,N_45192,N_45187);
nand U45580 (N_45580,N_45455,N_45272);
or U45581 (N_45581,N_45065,N_45376);
nand U45582 (N_45582,N_45337,N_45394);
and U45583 (N_45583,N_45059,N_45074);
nand U45584 (N_45584,N_45308,N_45061);
nor U45585 (N_45585,N_45066,N_45009);
xnor U45586 (N_45586,N_45022,N_45290);
nand U45587 (N_45587,N_45427,N_45196);
nand U45588 (N_45588,N_45212,N_45194);
xor U45589 (N_45589,N_45469,N_45213);
nand U45590 (N_45590,N_45091,N_45115);
or U45591 (N_45591,N_45235,N_45227);
and U45592 (N_45592,N_45393,N_45116);
nor U45593 (N_45593,N_45082,N_45178);
or U45594 (N_45594,N_45173,N_45444);
or U45595 (N_45595,N_45107,N_45015);
and U45596 (N_45596,N_45417,N_45093);
xor U45597 (N_45597,N_45369,N_45334);
nand U45598 (N_45598,N_45299,N_45097);
nand U45599 (N_45599,N_45088,N_45102);
and U45600 (N_45600,N_45135,N_45146);
xnor U45601 (N_45601,N_45456,N_45033);
or U45602 (N_45602,N_45421,N_45106);
nand U45603 (N_45603,N_45343,N_45133);
xnor U45604 (N_45604,N_45342,N_45193);
and U45605 (N_45605,N_45476,N_45312);
xnor U45606 (N_45606,N_45448,N_45480);
and U45607 (N_45607,N_45099,N_45180);
and U45608 (N_45608,N_45286,N_45344);
nand U45609 (N_45609,N_45140,N_45171);
nand U45610 (N_45610,N_45381,N_45440);
xnor U45611 (N_45611,N_45258,N_45118);
and U45612 (N_45612,N_45144,N_45494);
nand U45613 (N_45613,N_45094,N_45176);
nor U45614 (N_45614,N_45479,N_45030);
nor U45615 (N_45615,N_45096,N_45429);
nand U45616 (N_45616,N_45377,N_45081);
xor U45617 (N_45617,N_45282,N_45226);
or U45618 (N_45618,N_45112,N_45481);
and U45619 (N_45619,N_45499,N_45003);
nand U45620 (N_45620,N_45137,N_45387);
xnor U45621 (N_45621,N_45358,N_45175);
and U45622 (N_45622,N_45230,N_45131);
or U45623 (N_45623,N_45384,N_45068);
or U45624 (N_45624,N_45306,N_45027);
and U45625 (N_45625,N_45269,N_45298);
and U45626 (N_45626,N_45359,N_45053);
nor U45627 (N_45627,N_45148,N_45195);
xnor U45628 (N_45628,N_45104,N_45257);
nand U45629 (N_45629,N_45153,N_45475);
xor U45630 (N_45630,N_45161,N_45211);
and U45631 (N_45631,N_45132,N_45401);
xor U45632 (N_45632,N_45254,N_45005);
nand U45633 (N_45633,N_45070,N_45408);
and U45634 (N_45634,N_45076,N_45311);
and U45635 (N_45635,N_45277,N_45310);
nor U45636 (N_45636,N_45452,N_45085);
nor U45637 (N_45637,N_45295,N_45373);
or U45638 (N_45638,N_45349,N_45040);
nand U45639 (N_45639,N_45214,N_45016);
and U45640 (N_45640,N_45418,N_45034);
nand U45641 (N_45641,N_45039,N_45051);
or U45642 (N_45642,N_45410,N_45360);
nor U45643 (N_45643,N_45439,N_45264);
and U45644 (N_45644,N_45232,N_45457);
or U45645 (N_45645,N_45170,N_45186);
and U45646 (N_45646,N_45155,N_45159);
xnor U45647 (N_45647,N_45062,N_45284);
and U45648 (N_45648,N_45197,N_45013);
or U45649 (N_45649,N_45219,N_45397);
xnor U45650 (N_45650,N_45152,N_45379);
nand U45651 (N_45651,N_45242,N_45090);
xor U45652 (N_45652,N_45101,N_45396);
nor U45653 (N_45653,N_45319,N_45482);
nor U45654 (N_45654,N_45128,N_45372);
or U45655 (N_45655,N_45326,N_45493);
nand U45656 (N_45656,N_45035,N_45466);
or U45657 (N_45657,N_45496,N_45454);
xnor U45658 (N_45658,N_45139,N_45198);
nand U45659 (N_45659,N_45300,N_45276);
and U45660 (N_45660,N_45345,N_45243);
nand U45661 (N_45661,N_45388,N_45126);
xnor U45662 (N_45662,N_45248,N_45405);
nand U45663 (N_45663,N_45314,N_45224);
nand U45664 (N_45664,N_45151,N_45089);
nand U45665 (N_45665,N_45177,N_45252);
nor U45666 (N_45666,N_45485,N_45487);
nor U45667 (N_45667,N_45402,N_45293);
nor U45668 (N_45668,N_45267,N_45473);
and U45669 (N_45669,N_45483,N_45352);
and U45670 (N_45670,N_45273,N_45239);
nand U45671 (N_45671,N_45145,N_45157);
nor U45672 (N_45672,N_45234,N_45084);
xor U45673 (N_45673,N_45332,N_45361);
xor U45674 (N_45674,N_45075,N_45398);
nand U45675 (N_45675,N_45315,N_45183);
nor U45676 (N_45676,N_45166,N_45018);
xnor U45677 (N_45677,N_45050,N_45125);
xor U45678 (N_45678,N_45209,N_45036);
nand U45679 (N_45679,N_45309,N_45474);
or U45680 (N_45680,N_45468,N_45236);
xnor U45681 (N_45681,N_45169,N_45199);
nand U45682 (N_45682,N_45459,N_45433);
xnor U45683 (N_45683,N_45316,N_45055);
xnor U45684 (N_45684,N_45441,N_45484);
nor U45685 (N_45685,N_45149,N_45203);
or U45686 (N_45686,N_45014,N_45453);
nand U45687 (N_45687,N_45414,N_45385);
xor U45688 (N_45688,N_45399,N_45167);
nand U45689 (N_45689,N_45406,N_45335);
nor U45690 (N_45690,N_45231,N_45087);
nand U45691 (N_45691,N_45150,N_45288);
nor U45692 (N_45692,N_45067,N_45470);
xnor U45693 (N_45693,N_45058,N_45240);
nor U45694 (N_45694,N_45038,N_45012);
or U45695 (N_45695,N_45037,N_45043);
nor U45696 (N_45696,N_45244,N_45024);
nor U45697 (N_45697,N_45338,N_45275);
and U45698 (N_45698,N_45119,N_45297);
and U45699 (N_45699,N_45080,N_45303);
and U45700 (N_45700,N_45400,N_45320);
and U45701 (N_45701,N_45424,N_45328);
and U45702 (N_45702,N_45120,N_45449);
or U45703 (N_45703,N_45392,N_45371);
nor U45704 (N_45704,N_45190,N_45130);
or U45705 (N_45705,N_45330,N_45208);
nand U45706 (N_45706,N_45279,N_45168);
xnor U45707 (N_45707,N_45138,N_45191);
nor U45708 (N_45708,N_45042,N_45495);
nor U45709 (N_45709,N_45301,N_45216);
xor U45710 (N_45710,N_45253,N_45238);
nand U45711 (N_45711,N_45021,N_45010);
nor U45712 (N_45712,N_45217,N_45228);
nor U45713 (N_45713,N_45302,N_45237);
or U45714 (N_45714,N_45445,N_45006);
xnor U45715 (N_45715,N_45281,N_45069);
and U45716 (N_45716,N_45486,N_45438);
xor U45717 (N_45717,N_45305,N_45136);
xnor U45718 (N_45718,N_45221,N_45291);
and U45719 (N_45719,N_45436,N_45241);
nand U45720 (N_45720,N_45383,N_45340);
nor U45721 (N_45721,N_45123,N_45251);
nor U45722 (N_45722,N_45355,N_45366);
nand U45723 (N_45723,N_45415,N_45380);
or U45724 (N_45724,N_45346,N_45095);
nor U45725 (N_45725,N_45443,N_45259);
or U45726 (N_45726,N_45477,N_45200);
or U45727 (N_45727,N_45391,N_45347);
or U45728 (N_45728,N_45313,N_45465);
nand U45729 (N_45729,N_45285,N_45395);
xor U45730 (N_45730,N_45467,N_45127);
or U45731 (N_45731,N_45389,N_45121);
or U45732 (N_45732,N_45321,N_45063);
nand U45733 (N_45733,N_45154,N_45323);
nand U45734 (N_45734,N_45341,N_45103);
nand U45735 (N_45735,N_45270,N_45073);
xnor U45736 (N_45736,N_45164,N_45026);
nand U45737 (N_45737,N_45124,N_45000);
and U45738 (N_45738,N_45432,N_45261);
nor U45739 (N_45739,N_45156,N_45463);
and U45740 (N_45740,N_45100,N_45271);
nand U45741 (N_45741,N_45450,N_45174);
and U45742 (N_45742,N_45374,N_45307);
xnor U45743 (N_45743,N_45407,N_45492);
xor U45744 (N_45744,N_45111,N_45322);
or U45745 (N_45745,N_45189,N_45185);
or U45746 (N_45746,N_45158,N_45202);
nor U45747 (N_45747,N_45350,N_45134);
or U45748 (N_45748,N_45304,N_45079);
and U45749 (N_45749,N_45098,N_45023);
or U45750 (N_45750,N_45067,N_45035);
and U45751 (N_45751,N_45253,N_45490);
and U45752 (N_45752,N_45419,N_45112);
or U45753 (N_45753,N_45243,N_45164);
xor U45754 (N_45754,N_45143,N_45033);
nor U45755 (N_45755,N_45391,N_45237);
or U45756 (N_45756,N_45224,N_45270);
nor U45757 (N_45757,N_45051,N_45363);
nand U45758 (N_45758,N_45304,N_45260);
xor U45759 (N_45759,N_45473,N_45146);
or U45760 (N_45760,N_45472,N_45349);
and U45761 (N_45761,N_45241,N_45015);
nor U45762 (N_45762,N_45289,N_45177);
and U45763 (N_45763,N_45461,N_45325);
nand U45764 (N_45764,N_45113,N_45285);
or U45765 (N_45765,N_45218,N_45287);
or U45766 (N_45766,N_45440,N_45380);
and U45767 (N_45767,N_45023,N_45471);
nor U45768 (N_45768,N_45255,N_45347);
nand U45769 (N_45769,N_45161,N_45104);
or U45770 (N_45770,N_45257,N_45154);
nand U45771 (N_45771,N_45482,N_45430);
or U45772 (N_45772,N_45451,N_45433);
xor U45773 (N_45773,N_45000,N_45225);
nand U45774 (N_45774,N_45286,N_45316);
nor U45775 (N_45775,N_45051,N_45452);
or U45776 (N_45776,N_45220,N_45457);
nand U45777 (N_45777,N_45342,N_45435);
or U45778 (N_45778,N_45034,N_45051);
nand U45779 (N_45779,N_45384,N_45262);
nor U45780 (N_45780,N_45115,N_45318);
or U45781 (N_45781,N_45154,N_45277);
nor U45782 (N_45782,N_45442,N_45224);
xor U45783 (N_45783,N_45133,N_45041);
or U45784 (N_45784,N_45240,N_45272);
xor U45785 (N_45785,N_45405,N_45360);
or U45786 (N_45786,N_45344,N_45007);
nor U45787 (N_45787,N_45032,N_45386);
and U45788 (N_45788,N_45019,N_45306);
nand U45789 (N_45789,N_45117,N_45208);
and U45790 (N_45790,N_45484,N_45037);
or U45791 (N_45791,N_45330,N_45011);
nor U45792 (N_45792,N_45427,N_45030);
or U45793 (N_45793,N_45346,N_45312);
nor U45794 (N_45794,N_45042,N_45332);
and U45795 (N_45795,N_45276,N_45158);
nor U45796 (N_45796,N_45031,N_45411);
nor U45797 (N_45797,N_45265,N_45386);
nand U45798 (N_45798,N_45089,N_45126);
and U45799 (N_45799,N_45044,N_45057);
or U45800 (N_45800,N_45271,N_45229);
nand U45801 (N_45801,N_45113,N_45103);
nor U45802 (N_45802,N_45280,N_45049);
nand U45803 (N_45803,N_45310,N_45283);
xor U45804 (N_45804,N_45004,N_45467);
and U45805 (N_45805,N_45073,N_45051);
xor U45806 (N_45806,N_45078,N_45398);
nand U45807 (N_45807,N_45071,N_45484);
and U45808 (N_45808,N_45332,N_45224);
xor U45809 (N_45809,N_45153,N_45006);
nor U45810 (N_45810,N_45365,N_45417);
and U45811 (N_45811,N_45241,N_45258);
xnor U45812 (N_45812,N_45337,N_45222);
nand U45813 (N_45813,N_45082,N_45219);
nor U45814 (N_45814,N_45258,N_45242);
nand U45815 (N_45815,N_45058,N_45182);
and U45816 (N_45816,N_45385,N_45477);
xnor U45817 (N_45817,N_45138,N_45118);
or U45818 (N_45818,N_45251,N_45249);
xor U45819 (N_45819,N_45331,N_45156);
nor U45820 (N_45820,N_45085,N_45217);
nand U45821 (N_45821,N_45111,N_45064);
and U45822 (N_45822,N_45406,N_45124);
or U45823 (N_45823,N_45009,N_45319);
or U45824 (N_45824,N_45078,N_45300);
nand U45825 (N_45825,N_45341,N_45274);
and U45826 (N_45826,N_45460,N_45428);
nor U45827 (N_45827,N_45270,N_45007);
or U45828 (N_45828,N_45019,N_45313);
nand U45829 (N_45829,N_45122,N_45388);
and U45830 (N_45830,N_45185,N_45263);
xnor U45831 (N_45831,N_45339,N_45368);
nand U45832 (N_45832,N_45390,N_45005);
xor U45833 (N_45833,N_45270,N_45416);
xnor U45834 (N_45834,N_45069,N_45402);
and U45835 (N_45835,N_45198,N_45264);
or U45836 (N_45836,N_45007,N_45129);
or U45837 (N_45837,N_45003,N_45458);
nor U45838 (N_45838,N_45014,N_45072);
nor U45839 (N_45839,N_45364,N_45375);
nor U45840 (N_45840,N_45051,N_45208);
nor U45841 (N_45841,N_45252,N_45082);
or U45842 (N_45842,N_45194,N_45367);
nand U45843 (N_45843,N_45228,N_45385);
and U45844 (N_45844,N_45237,N_45183);
xor U45845 (N_45845,N_45222,N_45229);
xnor U45846 (N_45846,N_45356,N_45494);
nor U45847 (N_45847,N_45088,N_45179);
nand U45848 (N_45848,N_45471,N_45181);
nand U45849 (N_45849,N_45300,N_45047);
nor U45850 (N_45850,N_45186,N_45344);
xor U45851 (N_45851,N_45146,N_45177);
xor U45852 (N_45852,N_45236,N_45083);
nor U45853 (N_45853,N_45346,N_45048);
nand U45854 (N_45854,N_45142,N_45250);
xnor U45855 (N_45855,N_45378,N_45212);
and U45856 (N_45856,N_45333,N_45160);
xnor U45857 (N_45857,N_45203,N_45328);
or U45858 (N_45858,N_45080,N_45452);
nand U45859 (N_45859,N_45212,N_45136);
xor U45860 (N_45860,N_45080,N_45358);
nand U45861 (N_45861,N_45046,N_45469);
nand U45862 (N_45862,N_45127,N_45162);
nor U45863 (N_45863,N_45015,N_45445);
nor U45864 (N_45864,N_45301,N_45209);
nand U45865 (N_45865,N_45191,N_45047);
nor U45866 (N_45866,N_45247,N_45005);
and U45867 (N_45867,N_45317,N_45186);
and U45868 (N_45868,N_45481,N_45200);
nor U45869 (N_45869,N_45237,N_45468);
nor U45870 (N_45870,N_45282,N_45215);
and U45871 (N_45871,N_45047,N_45343);
nor U45872 (N_45872,N_45406,N_45056);
and U45873 (N_45873,N_45340,N_45027);
nor U45874 (N_45874,N_45441,N_45260);
or U45875 (N_45875,N_45371,N_45329);
and U45876 (N_45876,N_45022,N_45393);
xor U45877 (N_45877,N_45095,N_45225);
nor U45878 (N_45878,N_45141,N_45146);
nand U45879 (N_45879,N_45223,N_45146);
nand U45880 (N_45880,N_45031,N_45150);
or U45881 (N_45881,N_45428,N_45130);
nand U45882 (N_45882,N_45142,N_45382);
or U45883 (N_45883,N_45153,N_45086);
or U45884 (N_45884,N_45252,N_45217);
and U45885 (N_45885,N_45368,N_45136);
xor U45886 (N_45886,N_45125,N_45196);
nor U45887 (N_45887,N_45015,N_45064);
nor U45888 (N_45888,N_45133,N_45312);
or U45889 (N_45889,N_45255,N_45382);
nor U45890 (N_45890,N_45069,N_45108);
nand U45891 (N_45891,N_45192,N_45277);
and U45892 (N_45892,N_45144,N_45095);
nor U45893 (N_45893,N_45219,N_45292);
nor U45894 (N_45894,N_45041,N_45009);
nor U45895 (N_45895,N_45049,N_45227);
nor U45896 (N_45896,N_45193,N_45031);
and U45897 (N_45897,N_45155,N_45324);
or U45898 (N_45898,N_45220,N_45249);
or U45899 (N_45899,N_45435,N_45242);
and U45900 (N_45900,N_45156,N_45171);
or U45901 (N_45901,N_45230,N_45449);
nor U45902 (N_45902,N_45480,N_45192);
nand U45903 (N_45903,N_45221,N_45083);
nor U45904 (N_45904,N_45114,N_45451);
nor U45905 (N_45905,N_45185,N_45098);
and U45906 (N_45906,N_45429,N_45478);
nand U45907 (N_45907,N_45166,N_45351);
xnor U45908 (N_45908,N_45426,N_45171);
xnor U45909 (N_45909,N_45235,N_45043);
and U45910 (N_45910,N_45237,N_45247);
or U45911 (N_45911,N_45097,N_45452);
and U45912 (N_45912,N_45263,N_45461);
nand U45913 (N_45913,N_45404,N_45251);
nor U45914 (N_45914,N_45460,N_45099);
xnor U45915 (N_45915,N_45296,N_45194);
nor U45916 (N_45916,N_45314,N_45254);
or U45917 (N_45917,N_45034,N_45181);
or U45918 (N_45918,N_45121,N_45233);
or U45919 (N_45919,N_45444,N_45238);
xnor U45920 (N_45920,N_45279,N_45098);
nor U45921 (N_45921,N_45111,N_45063);
and U45922 (N_45922,N_45379,N_45039);
nand U45923 (N_45923,N_45429,N_45222);
and U45924 (N_45924,N_45294,N_45104);
nand U45925 (N_45925,N_45003,N_45095);
and U45926 (N_45926,N_45433,N_45315);
nand U45927 (N_45927,N_45374,N_45253);
and U45928 (N_45928,N_45066,N_45287);
nand U45929 (N_45929,N_45328,N_45438);
nand U45930 (N_45930,N_45096,N_45157);
or U45931 (N_45931,N_45230,N_45041);
nor U45932 (N_45932,N_45309,N_45416);
xor U45933 (N_45933,N_45181,N_45193);
or U45934 (N_45934,N_45341,N_45328);
or U45935 (N_45935,N_45100,N_45204);
nor U45936 (N_45936,N_45421,N_45329);
xor U45937 (N_45937,N_45332,N_45205);
or U45938 (N_45938,N_45170,N_45485);
xor U45939 (N_45939,N_45393,N_45062);
nand U45940 (N_45940,N_45082,N_45355);
nand U45941 (N_45941,N_45103,N_45274);
nor U45942 (N_45942,N_45119,N_45400);
nand U45943 (N_45943,N_45343,N_45221);
or U45944 (N_45944,N_45092,N_45486);
xnor U45945 (N_45945,N_45283,N_45014);
or U45946 (N_45946,N_45211,N_45059);
or U45947 (N_45947,N_45048,N_45016);
nor U45948 (N_45948,N_45465,N_45214);
nor U45949 (N_45949,N_45438,N_45444);
nand U45950 (N_45950,N_45060,N_45377);
and U45951 (N_45951,N_45419,N_45440);
xnor U45952 (N_45952,N_45267,N_45313);
and U45953 (N_45953,N_45012,N_45034);
nand U45954 (N_45954,N_45013,N_45126);
nor U45955 (N_45955,N_45337,N_45150);
and U45956 (N_45956,N_45071,N_45081);
or U45957 (N_45957,N_45000,N_45169);
xnor U45958 (N_45958,N_45229,N_45402);
xor U45959 (N_45959,N_45344,N_45340);
nand U45960 (N_45960,N_45057,N_45143);
nor U45961 (N_45961,N_45240,N_45135);
xor U45962 (N_45962,N_45002,N_45224);
and U45963 (N_45963,N_45353,N_45155);
and U45964 (N_45964,N_45382,N_45093);
xor U45965 (N_45965,N_45003,N_45070);
or U45966 (N_45966,N_45453,N_45316);
nor U45967 (N_45967,N_45070,N_45116);
xor U45968 (N_45968,N_45127,N_45174);
and U45969 (N_45969,N_45266,N_45103);
xnor U45970 (N_45970,N_45092,N_45097);
nand U45971 (N_45971,N_45166,N_45435);
nand U45972 (N_45972,N_45293,N_45099);
xnor U45973 (N_45973,N_45323,N_45015);
and U45974 (N_45974,N_45177,N_45212);
and U45975 (N_45975,N_45092,N_45063);
nor U45976 (N_45976,N_45494,N_45294);
or U45977 (N_45977,N_45317,N_45057);
or U45978 (N_45978,N_45368,N_45018);
xor U45979 (N_45979,N_45410,N_45477);
or U45980 (N_45980,N_45104,N_45404);
nor U45981 (N_45981,N_45232,N_45219);
xor U45982 (N_45982,N_45144,N_45343);
or U45983 (N_45983,N_45134,N_45490);
nor U45984 (N_45984,N_45245,N_45027);
and U45985 (N_45985,N_45154,N_45380);
or U45986 (N_45986,N_45128,N_45177);
or U45987 (N_45987,N_45337,N_45169);
nor U45988 (N_45988,N_45314,N_45313);
or U45989 (N_45989,N_45469,N_45192);
nand U45990 (N_45990,N_45086,N_45393);
xnor U45991 (N_45991,N_45484,N_45172);
and U45992 (N_45992,N_45260,N_45077);
nand U45993 (N_45993,N_45445,N_45104);
xnor U45994 (N_45994,N_45402,N_45196);
nor U45995 (N_45995,N_45091,N_45378);
or U45996 (N_45996,N_45291,N_45082);
nor U45997 (N_45997,N_45255,N_45433);
xnor U45998 (N_45998,N_45393,N_45339);
or U45999 (N_45999,N_45184,N_45352);
xnor U46000 (N_46000,N_45590,N_45565);
xor U46001 (N_46001,N_45848,N_45600);
nand U46002 (N_46002,N_45850,N_45718);
xor U46003 (N_46003,N_45883,N_45659);
and U46004 (N_46004,N_45938,N_45835);
and U46005 (N_46005,N_45501,N_45559);
nand U46006 (N_46006,N_45530,N_45866);
or U46007 (N_46007,N_45789,N_45690);
and U46008 (N_46008,N_45933,N_45822);
and U46009 (N_46009,N_45792,N_45527);
xnor U46010 (N_46010,N_45512,N_45628);
nand U46011 (N_46011,N_45855,N_45920);
and U46012 (N_46012,N_45516,N_45844);
nand U46013 (N_46013,N_45763,N_45661);
nor U46014 (N_46014,N_45924,N_45767);
nand U46015 (N_46015,N_45837,N_45646);
and U46016 (N_46016,N_45941,N_45931);
or U46017 (N_46017,N_45687,N_45821);
nand U46018 (N_46018,N_45871,N_45964);
nor U46019 (N_46019,N_45984,N_45673);
nand U46020 (N_46020,N_45776,N_45680);
and U46021 (N_46021,N_45874,N_45803);
or U46022 (N_46022,N_45846,N_45774);
xnor U46023 (N_46023,N_45531,N_45532);
or U46024 (N_46024,N_45670,N_45961);
or U46025 (N_46025,N_45733,N_45651);
nand U46026 (N_46026,N_45574,N_45609);
nor U46027 (N_46027,N_45591,N_45905);
nand U46028 (N_46028,N_45840,N_45765);
nand U46029 (N_46029,N_45607,N_45704);
xnor U46030 (N_46030,N_45580,N_45599);
nand U46031 (N_46031,N_45809,N_45503);
nand U46032 (N_46032,N_45640,N_45819);
xnor U46033 (N_46033,N_45621,N_45948);
nand U46034 (N_46034,N_45854,N_45947);
xor U46035 (N_46035,N_45943,N_45973);
nand U46036 (N_46036,N_45608,N_45692);
and U46037 (N_46037,N_45875,N_45633);
and U46038 (N_46038,N_45613,N_45894);
xor U46039 (N_46039,N_45726,N_45965);
nand U46040 (N_46040,N_45707,N_45836);
nand U46041 (N_46041,N_45790,N_45696);
and U46042 (N_46042,N_45968,N_45829);
nor U46043 (N_46043,N_45877,N_45798);
and U46044 (N_46044,N_45695,N_45643);
nand U46045 (N_46045,N_45597,N_45614);
and U46046 (N_46046,N_45625,N_45885);
xnor U46047 (N_46047,N_45721,N_45969);
or U46048 (N_46048,N_45669,N_45998);
nand U46049 (N_46049,N_45999,N_45691);
xnor U46050 (N_46050,N_45754,N_45978);
or U46051 (N_46051,N_45760,N_45594);
or U46052 (N_46052,N_45912,N_45557);
nand U46053 (N_46053,N_45826,N_45517);
nand U46054 (N_46054,N_45824,N_45800);
xor U46055 (N_46055,N_45783,N_45593);
nand U46056 (N_46056,N_45980,N_45538);
or U46057 (N_46057,N_45811,N_45572);
or U46058 (N_46058,N_45768,N_45917);
and U46059 (N_46059,N_45554,N_45505);
xor U46060 (N_46060,N_45683,N_45890);
xor U46061 (N_46061,N_45723,N_45934);
nand U46062 (N_46062,N_45719,N_45701);
or U46063 (N_46063,N_45658,N_45955);
nand U46064 (N_46064,N_45750,N_45863);
and U46065 (N_46065,N_45911,N_45975);
nand U46066 (N_46066,N_45903,N_45518);
and U46067 (N_46067,N_45868,N_45963);
xnor U46068 (N_46068,N_45734,N_45992);
and U46069 (N_46069,N_45578,N_45898);
nand U46070 (N_46070,N_45960,N_45888);
or U46071 (N_46071,N_45676,N_45828);
or U46072 (N_46072,N_45663,N_45981);
or U46073 (N_46073,N_45936,N_45810);
nand U46074 (N_46074,N_45511,N_45852);
and U46075 (N_46075,N_45534,N_45678);
or U46076 (N_46076,N_45504,N_45839);
xnor U46077 (N_46077,N_45629,N_45714);
xnor U46078 (N_46078,N_45588,N_45649);
xnor U46079 (N_46079,N_45583,N_45862);
and U46080 (N_46080,N_45652,N_45910);
nand U46081 (N_46081,N_45575,N_45513);
or U46082 (N_46082,N_45856,N_45675);
nand U46083 (N_46083,N_45508,N_45841);
nand U46084 (N_46084,N_45681,N_45568);
xor U46085 (N_46085,N_45756,N_45878);
or U46086 (N_46086,N_45864,N_45648);
nand U46087 (N_46087,N_45728,N_45758);
and U46088 (N_46088,N_45705,N_45547);
and U46089 (N_46089,N_45660,N_45786);
or U46090 (N_46090,N_45672,N_45994);
xor U46091 (N_46091,N_45944,N_45526);
or U46092 (N_46092,N_45779,N_45677);
nor U46093 (N_46093,N_45967,N_45736);
xnor U46094 (N_46094,N_45951,N_45713);
xnor U46095 (N_46095,N_45823,N_45805);
xnor U46096 (N_46096,N_45569,N_45684);
nand U46097 (N_46097,N_45742,N_45971);
or U46098 (N_46098,N_45586,N_45612);
or U46099 (N_46099,N_45759,N_45579);
or U46100 (N_46100,N_45989,N_45830);
xor U46101 (N_46101,N_45622,N_45639);
or U46102 (N_46102,N_45617,N_45623);
and U46103 (N_46103,N_45956,N_45757);
and U46104 (N_46104,N_45869,N_45694);
xnor U46105 (N_46105,N_45642,N_45630);
xor U46106 (N_46106,N_45781,N_45551);
xor U46107 (N_46107,N_45710,N_45686);
or U46108 (N_46108,N_45730,N_45748);
xnor U46109 (N_46109,N_45747,N_45553);
and U46110 (N_46110,N_45679,N_45515);
nand U46111 (N_46111,N_45884,N_45901);
xnor U46112 (N_46112,N_45537,N_45950);
xor U46113 (N_46113,N_45667,N_45794);
nor U46114 (N_46114,N_45814,N_45571);
and U46115 (N_46115,N_45528,N_45555);
and U46116 (N_46116,N_45619,N_45550);
nand U46117 (N_46117,N_45922,N_45627);
nand U46118 (N_46118,N_45560,N_45778);
nor U46119 (N_46119,N_45573,N_45804);
nor U46120 (N_46120,N_45769,N_45521);
nor U46121 (N_46121,N_45787,N_45953);
nor U46122 (N_46122,N_45653,N_45815);
xnor U46123 (N_46123,N_45698,N_45732);
xnor U46124 (N_46124,N_45596,N_45558);
nand U46125 (N_46125,N_45566,N_45520);
nand U46126 (N_46126,N_45775,N_45927);
nand U46127 (N_46127,N_45749,N_45570);
and U46128 (N_46128,N_45782,N_45847);
xor U46129 (N_46129,N_45785,N_45602);
nand U46130 (N_46130,N_45682,N_45780);
nor U46131 (N_46131,N_45977,N_45706);
or U46132 (N_46132,N_45509,N_45812);
xnor U46133 (N_46133,N_45935,N_45631);
or U46134 (N_46134,N_45949,N_45740);
nand U46135 (N_46135,N_45548,N_45584);
nor U46136 (N_46136,N_45895,N_45729);
and U46137 (N_46137,N_45891,N_45539);
nor U46138 (N_46138,N_45793,N_45595);
and U46139 (N_46139,N_45549,N_45751);
xor U46140 (N_46140,N_45788,N_45900);
nand U46141 (N_46141,N_45795,N_45715);
or U46142 (N_46142,N_45746,N_45816);
nor U46143 (N_46143,N_45909,N_45561);
or U46144 (N_46144,N_45522,N_45519);
xnor U46145 (N_46145,N_45817,N_45688);
xnor U46146 (N_46146,N_45618,N_45657);
nor U46147 (N_46147,N_45611,N_45562);
xor U46148 (N_46148,N_45946,N_45604);
nor U46149 (N_46149,N_45666,N_45834);
nor U46150 (N_46150,N_45791,N_45589);
and U46151 (N_46151,N_45882,N_45879);
or U46152 (N_46152,N_45893,N_45529);
nor U46153 (N_46153,N_45697,N_45873);
or U46154 (N_46154,N_45725,N_45603);
nor U46155 (N_46155,N_45876,N_45716);
xnor U46156 (N_46156,N_45818,N_45708);
or U46157 (N_46157,N_45752,N_45693);
or U46158 (N_46158,N_45867,N_45958);
or U46159 (N_46159,N_45797,N_45932);
or U46160 (N_46160,N_45654,N_45655);
xnor U46161 (N_46161,N_45907,N_45929);
xor U46162 (N_46162,N_45906,N_45544);
and U46163 (N_46163,N_45926,N_45510);
nor U46164 (N_46164,N_45974,N_45506);
nor U46165 (N_46165,N_45889,N_45870);
and U46166 (N_46166,N_45923,N_45671);
and U46167 (N_46167,N_45857,N_45770);
and U46168 (N_46168,N_45880,N_45576);
xnor U46169 (N_46169,N_45914,N_45616);
and U46170 (N_46170,N_45982,N_45674);
or U46171 (N_46171,N_45919,N_45916);
or U46172 (N_46172,N_45536,N_45668);
and U46173 (N_46173,N_45500,N_45928);
or U46174 (N_46174,N_45892,N_45921);
and U46175 (N_46175,N_45582,N_45925);
nand U46176 (N_46176,N_45820,N_45753);
or U46177 (N_46177,N_45664,N_45886);
or U46178 (N_46178,N_45845,N_45606);
xnor U46179 (N_46179,N_45831,N_45983);
xnor U46180 (N_46180,N_45996,N_45842);
nand U46181 (N_46181,N_45802,N_45620);
nor U46182 (N_46182,N_45897,N_45641);
nand U46183 (N_46183,N_45644,N_45535);
nand U46184 (N_46184,N_45540,N_45542);
or U46185 (N_46185,N_45796,N_45700);
xnor U46186 (N_46186,N_45722,N_45615);
or U46187 (N_46187,N_45985,N_45737);
or U46188 (N_46188,N_45662,N_45899);
or U46189 (N_46189,N_45711,N_45533);
xnor U46190 (N_46190,N_45717,N_45624);
nor U46191 (N_46191,N_45703,N_45861);
xnor U46192 (N_46192,N_45634,N_45720);
or U46193 (N_46193,N_45918,N_45952);
nor U46194 (N_46194,N_45638,N_45959);
or U46195 (N_46195,N_45970,N_45702);
nand U46196 (N_46196,N_45843,N_45712);
nor U46197 (N_46197,N_45945,N_45645);
or U46198 (N_46198,N_45865,N_45913);
and U46199 (N_46199,N_45849,N_45896);
nor U46200 (N_46200,N_45853,N_45808);
xor U46201 (N_46201,N_45632,N_45784);
and U46202 (N_46202,N_45979,N_45656);
xnor U46203 (N_46203,N_45564,N_45825);
or U46204 (N_46204,N_45727,N_45772);
xor U46205 (N_46205,N_45902,N_45685);
or U46206 (N_46206,N_45581,N_45709);
or U46207 (N_46207,N_45807,N_45601);
or U46208 (N_46208,N_45689,N_45915);
or U46209 (N_46209,N_45990,N_45777);
nor U46210 (N_46210,N_45567,N_45563);
xnor U46211 (N_46211,N_45773,N_45523);
nor U46212 (N_46212,N_45626,N_45764);
nand U46213 (N_46213,N_45592,N_45993);
and U46214 (N_46214,N_45525,N_45988);
and U46215 (N_46215,N_45587,N_45724);
and U46216 (N_46216,N_45524,N_45939);
nor U46217 (N_46217,N_45543,N_45745);
and U46218 (N_46218,N_45881,N_45851);
and U46219 (N_46219,N_45908,N_45514);
and U46220 (N_46220,N_45577,N_45799);
nand U46221 (N_46221,N_45546,N_45940);
nand U46222 (N_46222,N_45647,N_45762);
xor U46223 (N_46223,N_45771,N_45827);
and U46224 (N_46224,N_45997,N_45872);
nand U46225 (N_46225,N_45904,N_45552);
nor U46226 (N_46226,N_45743,N_45887);
nand U46227 (N_46227,N_45838,N_45650);
and U46228 (N_46228,N_45585,N_45635);
or U46229 (N_46229,N_45858,N_45942);
and U46230 (N_46230,N_45545,N_45860);
and U46231 (N_46231,N_45637,N_45976);
xnor U46232 (N_46232,N_45744,N_45598);
xor U46233 (N_46233,N_45987,N_45541);
xor U46234 (N_46234,N_45738,N_45801);
xor U46235 (N_46235,N_45502,N_45832);
xnor U46236 (N_46236,N_45986,N_45556);
nand U46237 (N_46237,N_45962,N_45937);
or U46238 (N_46238,N_45954,N_45930);
and U46239 (N_46239,N_45699,N_45766);
and U46240 (N_46240,N_45833,N_45813);
and U46241 (N_46241,N_45806,N_45966);
nor U46242 (N_46242,N_45739,N_45735);
xor U46243 (N_46243,N_45731,N_45859);
and U46244 (N_46244,N_45957,N_45755);
nand U46245 (N_46245,N_45605,N_45761);
and U46246 (N_46246,N_45610,N_45995);
and U46247 (N_46247,N_45972,N_45507);
and U46248 (N_46248,N_45741,N_45665);
and U46249 (N_46249,N_45636,N_45991);
xnor U46250 (N_46250,N_45929,N_45995);
and U46251 (N_46251,N_45693,N_45616);
nand U46252 (N_46252,N_45776,N_45915);
xor U46253 (N_46253,N_45654,N_45822);
or U46254 (N_46254,N_45748,N_45677);
xor U46255 (N_46255,N_45872,N_45676);
nand U46256 (N_46256,N_45987,N_45941);
nand U46257 (N_46257,N_45718,N_45591);
or U46258 (N_46258,N_45818,N_45673);
nand U46259 (N_46259,N_45631,N_45566);
nor U46260 (N_46260,N_45719,N_45831);
nand U46261 (N_46261,N_45726,N_45527);
nand U46262 (N_46262,N_45645,N_45541);
nor U46263 (N_46263,N_45926,N_45603);
nor U46264 (N_46264,N_45793,N_45632);
nor U46265 (N_46265,N_45538,N_45894);
xnor U46266 (N_46266,N_45551,N_45933);
nor U46267 (N_46267,N_45932,N_45965);
and U46268 (N_46268,N_45597,N_45723);
nor U46269 (N_46269,N_45629,N_45535);
nor U46270 (N_46270,N_45601,N_45823);
and U46271 (N_46271,N_45513,N_45589);
and U46272 (N_46272,N_45519,N_45711);
or U46273 (N_46273,N_45846,N_45527);
nor U46274 (N_46274,N_45820,N_45674);
nand U46275 (N_46275,N_45583,N_45828);
and U46276 (N_46276,N_45721,N_45609);
and U46277 (N_46277,N_45971,N_45574);
or U46278 (N_46278,N_45662,N_45572);
nand U46279 (N_46279,N_45697,N_45645);
xnor U46280 (N_46280,N_45972,N_45511);
or U46281 (N_46281,N_45509,N_45842);
nor U46282 (N_46282,N_45986,N_45929);
xor U46283 (N_46283,N_45885,N_45998);
or U46284 (N_46284,N_45886,N_45771);
and U46285 (N_46285,N_45583,N_45704);
and U46286 (N_46286,N_45812,N_45831);
nand U46287 (N_46287,N_45593,N_45525);
and U46288 (N_46288,N_45900,N_45895);
and U46289 (N_46289,N_45672,N_45778);
or U46290 (N_46290,N_45506,N_45793);
nand U46291 (N_46291,N_45795,N_45930);
nor U46292 (N_46292,N_45818,N_45850);
nor U46293 (N_46293,N_45771,N_45901);
xor U46294 (N_46294,N_45662,N_45717);
or U46295 (N_46295,N_45856,N_45691);
and U46296 (N_46296,N_45909,N_45588);
nor U46297 (N_46297,N_45519,N_45981);
and U46298 (N_46298,N_45813,N_45949);
xor U46299 (N_46299,N_45707,N_45500);
or U46300 (N_46300,N_45962,N_45607);
nor U46301 (N_46301,N_45820,N_45885);
or U46302 (N_46302,N_45849,N_45835);
or U46303 (N_46303,N_45958,N_45944);
xnor U46304 (N_46304,N_45630,N_45960);
nor U46305 (N_46305,N_45980,N_45802);
nand U46306 (N_46306,N_45877,N_45915);
nor U46307 (N_46307,N_45510,N_45538);
nand U46308 (N_46308,N_45703,N_45859);
and U46309 (N_46309,N_45916,N_45961);
nor U46310 (N_46310,N_45729,N_45821);
nand U46311 (N_46311,N_45550,N_45746);
or U46312 (N_46312,N_45703,N_45982);
or U46313 (N_46313,N_45821,N_45999);
nor U46314 (N_46314,N_45522,N_45745);
or U46315 (N_46315,N_45619,N_45582);
nand U46316 (N_46316,N_45725,N_45775);
nand U46317 (N_46317,N_45941,N_45858);
nand U46318 (N_46318,N_45886,N_45576);
and U46319 (N_46319,N_45749,N_45957);
nor U46320 (N_46320,N_45510,N_45541);
or U46321 (N_46321,N_45695,N_45962);
xor U46322 (N_46322,N_45869,N_45692);
nand U46323 (N_46323,N_45793,N_45916);
nand U46324 (N_46324,N_45990,N_45594);
nor U46325 (N_46325,N_45629,N_45778);
nor U46326 (N_46326,N_45514,N_45983);
nand U46327 (N_46327,N_45727,N_45640);
xnor U46328 (N_46328,N_45653,N_45811);
nand U46329 (N_46329,N_45902,N_45507);
nor U46330 (N_46330,N_45880,N_45848);
or U46331 (N_46331,N_45536,N_45750);
or U46332 (N_46332,N_45949,N_45688);
nand U46333 (N_46333,N_45578,N_45676);
or U46334 (N_46334,N_45524,N_45683);
xnor U46335 (N_46335,N_45729,N_45932);
nand U46336 (N_46336,N_45506,N_45664);
nand U46337 (N_46337,N_45885,N_45726);
nor U46338 (N_46338,N_45818,N_45634);
nor U46339 (N_46339,N_45774,N_45725);
xnor U46340 (N_46340,N_45951,N_45599);
nor U46341 (N_46341,N_45764,N_45782);
nand U46342 (N_46342,N_45898,N_45607);
or U46343 (N_46343,N_45672,N_45774);
nor U46344 (N_46344,N_45966,N_45815);
or U46345 (N_46345,N_45513,N_45509);
nor U46346 (N_46346,N_45598,N_45914);
and U46347 (N_46347,N_45563,N_45652);
xor U46348 (N_46348,N_45769,N_45646);
and U46349 (N_46349,N_45943,N_45902);
xor U46350 (N_46350,N_45671,N_45847);
or U46351 (N_46351,N_45541,N_45767);
nand U46352 (N_46352,N_45640,N_45698);
xnor U46353 (N_46353,N_45857,N_45949);
and U46354 (N_46354,N_45525,N_45648);
nor U46355 (N_46355,N_45744,N_45795);
or U46356 (N_46356,N_45608,N_45525);
nor U46357 (N_46357,N_45564,N_45972);
or U46358 (N_46358,N_45998,N_45822);
and U46359 (N_46359,N_45813,N_45638);
and U46360 (N_46360,N_45722,N_45563);
and U46361 (N_46361,N_45873,N_45552);
or U46362 (N_46362,N_45798,N_45507);
xor U46363 (N_46363,N_45639,N_45959);
xor U46364 (N_46364,N_45739,N_45882);
nor U46365 (N_46365,N_45986,N_45578);
nand U46366 (N_46366,N_45962,N_45859);
xor U46367 (N_46367,N_45816,N_45883);
or U46368 (N_46368,N_45831,N_45525);
xor U46369 (N_46369,N_45555,N_45665);
nor U46370 (N_46370,N_45989,N_45654);
nor U46371 (N_46371,N_45517,N_45819);
nor U46372 (N_46372,N_45730,N_45911);
xor U46373 (N_46373,N_45655,N_45716);
nand U46374 (N_46374,N_45862,N_45792);
and U46375 (N_46375,N_45653,N_45969);
nand U46376 (N_46376,N_45932,N_45945);
nor U46377 (N_46377,N_45897,N_45656);
nand U46378 (N_46378,N_45662,N_45847);
nor U46379 (N_46379,N_45800,N_45890);
nor U46380 (N_46380,N_45661,N_45966);
xor U46381 (N_46381,N_45949,N_45840);
xnor U46382 (N_46382,N_45558,N_45872);
nand U46383 (N_46383,N_45718,N_45797);
nand U46384 (N_46384,N_45840,N_45694);
nand U46385 (N_46385,N_45764,N_45826);
nand U46386 (N_46386,N_45511,N_45910);
and U46387 (N_46387,N_45575,N_45950);
nor U46388 (N_46388,N_45678,N_45736);
xnor U46389 (N_46389,N_45733,N_45566);
or U46390 (N_46390,N_45911,N_45589);
nand U46391 (N_46391,N_45635,N_45666);
nor U46392 (N_46392,N_45659,N_45729);
and U46393 (N_46393,N_45546,N_45910);
or U46394 (N_46394,N_45886,N_45747);
nor U46395 (N_46395,N_45979,N_45739);
and U46396 (N_46396,N_45837,N_45621);
xnor U46397 (N_46397,N_45652,N_45502);
and U46398 (N_46398,N_45829,N_45955);
and U46399 (N_46399,N_45863,N_45825);
and U46400 (N_46400,N_45890,N_45777);
or U46401 (N_46401,N_45546,N_45831);
or U46402 (N_46402,N_45966,N_45848);
xnor U46403 (N_46403,N_45946,N_45699);
xor U46404 (N_46404,N_45756,N_45823);
xnor U46405 (N_46405,N_45931,N_45605);
nor U46406 (N_46406,N_45908,N_45799);
xnor U46407 (N_46407,N_45514,N_45611);
or U46408 (N_46408,N_45859,N_45721);
nor U46409 (N_46409,N_45743,N_45560);
and U46410 (N_46410,N_45945,N_45912);
or U46411 (N_46411,N_45528,N_45593);
nand U46412 (N_46412,N_45875,N_45975);
xnor U46413 (N_46413,N_45830,N_45554);
nor U46414 (N_46414,N_45521,N_45679);
nor U46415 (N_46415,N_45629,N_45857);
and U46416 (N_46416,N_45888,N_45680);
or U46417 (N_46417,N_45996,N_45559);
nor U46418 (N_46418,N_45981,N_45891);
or U46419 (N_46419,N_45656,N_45858);
nand U46420 (N_46420,N_45883,N_45529);
and U46421 (N_46421,N_45905,N_45990);
and U46422 (N_46422,N_45581,N_45567);
nor U46423 (N_46423,N_45658,N_45518);
xnor U46424 (N_46424,N_45699,N_45955);
nor U46425 (N_46425,N_45761,N_45712);
nand U46426 (N_46426,N_45951,N_45838);
nand U46427 (N_46427,N_45548,N_45844);
or U46428 (N_46428,N_45660,N_45663);
and U46429 (N_46429,N_45954,N_45772);
nand U46430 (N_46430,N_45562,N_45888);
nand U46431 (N_46431,N_45970,N_45985);
xor U46432 (N_46432,N_45734,N_45980);
nor U46433 (N_46433,N_45653,N_45709);
or U46434 (N_46434,N_45534,N_45554);
xnor U46435 (N_46435,N_45988,N_45775);
nor U46436 (N_46436,N_45830,N_45781);
and U46437 (N_46437,N_45987,N_45961);
nor U46438 (N_46438,N_45987,N_45974);
and U46439 (N_46439,N_45995,N_45897);
or U46440 (N_46440,N_45708,N_45830);
or U46441 (N_46441,N_45736,N_45751);
xor U46442 (N_46442,N_45763,N_45768);
or U46443 (N_46443,N_45704,N_45509);
and U46444 (N_46444,N_45986,N_45585);
or U46445 (N_46445,N_45949,N_45503);
nor U46446 (N_46446,N_45855,N_45746);
or U46447 (N_46447,N_45930,N_45793);
or U46448 (N_46448,N_45669,N_45665);
xor U46449 (N_46449,N_45950,N_45998);
and U46450 (N_46450,N_45536,N_45699);
and U46451 (N_46451,N_45711,N_45764);
and U46452 (N_46452,N_45767,N_45595);
and U46453 (N_46453,N_45579,N_45571);
or U46454 (N_46454,N_45511,N_45893);
and U46455 (N_46455,N_45530,N_45995);
and U46456 (N_46456,N_45673,N_45829);
nor U46457 (N_46457,N_45937,N_45735);
nand U46458 (N_46458,N_45676,N_45548);
nor U46459 (N_46459,N_45628,N_45539);
xor U46460 (N_46460,N_45520,N_45892);
nand U46461 (N_46461,N_45780,N_45746);
xnor U46462 (N_46462,N_45677,N_45861);
nand U46463 (N_46463,N_45711,N_45563);
xnor U46464 (N_46464,N_45607,N_45624);
nor U46465 (N_46465,N_45632,N_45763);
and U46466 (N_46466,N_45829,N_45549);
and U46467 (N_46467,N_45834,N_45905);
or U46468 (N_46468,N_45704,N_45908);
nand U46469 (N_46469,N_45607,N_45531);
or U46470 (N_46470,N_45909,N_45750);
nor U46471 (N_46471,N_45759,N_45999);
xnor U46472 (N_46472,N_45814,N_45952);
or U46473 (N_46473,N_45636,N_45533);
and U46474 (N_46474,N_45854,N_45696);
nor U46475 (N_46475,N_45589,N_45977);
nor U46476 (N_46476,N_45838,N_45611);
or U46477 (N_46477,N_45646,N_45893);
or U46478 (N_46478,N_45672,N_45642);
nand U46479 (N_46479,N_45576,N_45574);
nand U46480 (N_46480,N_45583,N_45951);
nor U46481 (N_46481,N_45532,N_45681);
or U46482 (N_46482,N_45940,N_45840);
xor U46483 (N_46483,N_45544,N_45662);
and U46484 (N_46484,N_45650,N_45804);
or U46485 (N_46485,N_45843,N_45868);
or U46486 (N_46486,N_45550,N_45970);
and U46487 (N_46487,N_45755,N_45898);
and U46488 (N_46488,N_45892,N_45633);
or U46489 (N_46489,N_45644,N_45931);
and U46490 (N_46490,N_45540,N_45613);
nand U46491 (N_46491,N_45598,N_45665);
nor U46492 (N_46492,N_45936,N_45512);
xnor U46493 (N_46493,N_45717,N_45617);
or U46494 (N_46494,N_45554,N_45891);
nand U46495 (N_46495,N_45700,N_45976);
nand U46496 (N_46496,N_45846,N_45556);
or U46497 (N_46497,N_45968,N_45593);
or U46498 (N_46498,N_45948,N_45594);
xnor U46499 (N_46499,N_45765,N_45556);
nand U46500 (N_46500,N_46245,N_46464);
nand U46501 (N_46501,N_46278,N_46408);
xor U46502 (N_46502,N_46164,N_46400);
or U46503 (N_46503,N_46198,N_46039);
and U46504 (N_46504,N_46131,N_46075);
nand U46505 (N_46505,N_46376,N_46055);
nand U46506 (N_46506,N_46048,N_46280);
nor U46507 (N_46507,N_46314,N_46490);
xor U46508 (N_46508,N_46178,N_46140);
and U46509 (N_46509,N_46410,N_46390);
xnor U46510 (N_46510,N_46033,N_46392);
and U46511 (N_46511,N_46115,N_46316);
xnor U46512 (N_46512,N_46356,N_46391);
and U46513 (N_46513,N_46241,N_46344);
or U46514 (N_46514,N_46208,N_46035);
and U46515 (N_46515,N_46082,N_46433);
nand U46516 (N_46516,N_46149,N_46155);
nor U46517 (N_46517,N_46239,N_46006);
nand U46518 (N_46518,N_46494,N_46444);
and U46519 (N_46519,N_46188,N_46419);
and U46520 (N_46520,N_46050,N_46201);
nand U46521 (N_46521,N_46374,N_46475);
nand U46522 (N_46522,N_46125,N_46018);
nand U46523 (N_46523,N_46121,N_46322);
or U46524 (N_46524,N_46414,N_46284);
xnor U46525 (N_46525,N_46441,N_46065);
or U46526 (N_46526,N_46047,N_46158);
xor U46527 (N_46527,N_46171,N_46247);
xnor U46528 (N_46528,N_46199,N_46308);
xnor U46529 (N_46529,N_46383,N_46249);
xor U46530 (N_46530,N_46409,N_46486);
nand U46531 (N_46531,N_46498,N_46398);
xnor U46532 (N_46532,N_46237,N_46371);
and U46533 (N_46533,N_46029,N_46088);
and U46534 (N_46534,N_46362,N_46429);
nor U46535 (N_46535,N_46445,N_46386);
xor U46536 (N_46536,N_46217,N_46091);
or U46537 (N_46537,N_46016,N_46000);
nand U46538 (N_46538,N_46258,N_46477);
xnor U46539 (N_46539,N_46273,N_46160);
nor U46540 (N_46540,N_46313,N_46437);
or U46541 (N_46541,N_46312,N_46244);
nor U46542 (N_46542,N_46220,N_46305);
nand U46543 (N_46543,N_46087,N_46238);
xnor U46544 (N_46544,N_46421,N_46030);
nor U46545 (N_46545,N_46084,N_46484);
xnor U46546 (N_46546,N_46274,N_46123);
nor U46547 (N_46547,N_46195,N_46223);
and U46548 (N_46548,N_46031,N_46072);
and U46549 (N_46549,N_46222,N_46270);
nand U46550 (N_46550,N_46372,N_46009);
or U46551 (N_46551,N_46355,N_46460);
and U46552 (N_46552,N_46487,N_46397);
and U46553 (N_46553,N_46328,N_46012);
and U46554 (N_46554,N_46251,N_46483);
xor U46555 (N_46555,N_46299,N_46379);
and U46556 (N_46556,N_46387,N_46364);
xnor U46557 (N_46557,N_46458,N_46282);
nor U46558 (N_46558,N_46167,N_46022);
and U46559 (N_46559,N_46059,N_46097);
and U46560 (N_46560,N_46044,N_46004);
xnor U46561 (N_46561,N_46393,N_46028);
xnor U46562 (N_46562,N_46169,N_46331);
nor U46563 (N_46563,N_46315,N_46434);
xnor U46564 (N_46564,N_46061,N_46230);
xor U46565 (N_46565,N_46026,N_46343);
or U46566 (N_46566,N_46024,N_46262);
and U46567 (N_46567,N_46259,N_46263);
xnor U46568 (N_46568,N_46384,N_46177);
or U46569 (N_46569,N_46389,N_46333);
or U46570 (N_46570,N_46302,N_46066);
nand U46571 (N_46571,N_46481,N_46395);
or U46572 (N_46572,N_46112,N_46010);
xor U46573 (N_46573,N_46404,N_46277);
nand U46574 (N_46574,N_46037,N_46204);
and U46575 (N_46575,N_46211,N_46272);
nor U46576 (N_46576,N_46341,N_46459);
nand U46577 (N_46577,N_46126,N_46041);
or U46578 (N_46578,N_46034,N_46021);
and U46579 (N_46579,N_46426,N_46093);
xor U46580 (N_46580,N_46168,N_46170);
or U46581 (N_46581,N_46268,N_46349);
or U46582 (N_46582,N_46424,N_46099);
nor U46583 (N_46583,N_46428,N_46334);
xor U46584 (N_46584,N_46493,N_46467);
xnor U46585 (N_46585,N_46005,N_46447);
nor U46586 (N_46586,N_46076,N_46233);
xor U46587 (N_46587,N_46180,N_46157);
or U46588 (N_46588,N_46068,N_46250);
nand U46589 (N_46589,N_46219,N_46103);
nor U46590 (N_46590,N_46154,N_46163);
and U46591 (N_46591,N_46473,N_46200);
or U46592 (N_46592,N_46064,N_46435);
nand U46593 (N_46593,N_46260,N_46406);
nor U46594 (N_46594,N_46214,N_46221);
or U46595 (N_46595,N_46472,N_46422);
and U46596 (N_46596,N_46193,N_46118);
or U46597 (N_46597,N_46056,N_46046);
nand U46598 (N_46598,N_46095,N_46127);
nand U46599 (N_46599,N_46488,N_46363);
or U46600 (N_46600,N_46116,N_46216);
nor U46601 (N_46601,N_46176,N_46373);
or U46602 (N_46602,N_46412,N_46360);
and U46603 (N_46603,N_46296,N_46063);
xor U46604 (N_46604,N_46416,N_46367);
and U46605 (N_46605,N_46209,N_46069);
or U46606 (N_46606,N_46017,N_46456);
nor U46607 (N_46607,N_46318,N_46287);
or U46608 (N_46608,N_46080,N_46179);
and U46609 (N_46609,N_46020,N_46073);
xor U46610 (N_46610,N_46276,N_46196);
xnor U46611 (N_46611,N_46348,N_46206);
xnor U46612 (N_46612,N_46388,N_46492);
nand U46613 (N_46613,N_46338,N_46189);
or U46614 (N_46614,N_46045,N_46011);
or U46615 (N_46615,N_46114,N_46086);
and U46616 (N_46616,N_46161,N_46329);
nor U46617 (N_46617,N_46070,N_46215);
nand U46618 (N_46618,N_46254,N_46210);
nor U46619 (N_46619,N_46440,N_46134);
nand U46620 (N_46620,N_46330,N_46148);
nand U46621 (N_46621,N_46346,N_46181);
xnor U46622 (N_46622,N_46446,N_46147);
xor U46623 (N_46623,N_46124,N_46358);
xnor U46624 (N_46624,N_46347,N_46365);
nand U46625 (N_46625,N_46120,N_46232);
and U46626 (N_46626,N_46049,N_46234);
nor U46627 (N_46627,N_46345,N_46415);
xnor U46628 (N_46628,N_46236,N_46117);
and U46629 (N_46629,N_46256,N_46079);
xor U46630 (N_46630,N_46101,N_46336);
nor U46631 (N_46631,N_46288,N_46153);
xor U46632 (N_46632,N_46165,N_46067);
xnor U46633 (N_46633,N_46420,N_46340);
xnor U46634 (N_46634,N_46166,N_46190);
xnor U46635 (N_46635,N_46471,N_46156);
xnor U46636 (N_46636,N_46089,N_46227);
and U46637 (N_46637,N_46466,N_46369);
nand U46638 (N_46638,N_46394,N_46071);
nand U46639 (N_46639,N_46401,N_46417);
nor U46640 (N_46640,N_46378,N_46192);
xnor U46641 (N_46641,N_46354,N_46423);
nor U46642 (N_46642,N_46051,N_46310);
nand U46643 (N_46643,N_46111,N_46174);
and U46644 (N_46644,N_46271,N_46242);
xor U46645 (N_46645,N_46332,N_46275);
nor U46646 (N_46646,N_46130,N_46159);
or U46647 (N_46647,N_46311,N_46455);
nand U46648 (N_46648,N_46141,N_46324);
or U46649 (N_46649,N_46146,N_46054);
xnor U46650 (N_46650,N_46451,N_46339);
and U46651 (N_46651,N_46100,N_46499);
xor U46652 (N_46652,N_46052,N_46013);
nand U46653 (N_46653,N_46443,N_46301);
xor U46654 (N_46654,N_46300,N_46057);
nand U46655 (N_46655,N_46307,N_46032);
and U46656 (N_46656,N_46261,N_46269);
xnor U46657 (N_46657,N_46468,N_46139);
xnor U46658 (N_46658,N_46438,N_46497);
nand U46659 (N_46659,N_46402,N_46025);
and U46660 (N_46660,N_46042,N_46002);
nand U46661 (N_46661,N_46295,N_46491);
and U46662 (N_46662,N_46294,N_46145);
and U46663 (N_46663,N_46496,N_46135);
or U46664 (N_46664,N_46293,N_46436);
or U46665 (N_46665,N_46023,N_46027);
nor U46666 (N_46666,N_46399,N_46357);
or U46667 (N_46667,N_46474,N_46203);
and U46668 (N_46668,N_46137,N_46430);
nor U46669 (N_46669,N_46224,N_46187);
and U46670 (N_46670,N_46425,N_46062);
xor U46671 (N_46671,N_46335,N_46407);
or U46672 (N_46672,N_46418,N_46370);
nor U46673 (N_46673,N_46136,N_46366);
nand U46674 (N_46674,N_46291,N_46462);
nand U46675 (N_46675,N_46382,N_46479);
or U46676 (N_46676,N_46279,N_46337);
xor U46677 (N_46677,N_46183,N_46359);
nor U46678 (N_46678,N_46143,N_46102);
nand U46679 (N_46679,N_46194,N_46454);
nor U46680 (N_46680,N_46185,N_46197);
or U46681 (N_46681,N_46319,N_46213);
or U46682 (N_46682,N_46083,N_46298);
xor U46683 (N_46683,N_46150,N_46240);
xor U46684 (N_46684,N_46323,N_46375);
nand U46685 (N_46685,N_46105,N_46128);
or U46686 (N_46686,N_46252,N_46122);
nor U46687 (N_46687,N_46353,N_46439);
or U46688 (N_46688,N_46266,N_46038);
and U46689 (N_46689,N_46476,N_46077);
nand U46690 (N_46690,N_46133,N_46281);
nand U46691 (N_46691,N_46306,N_46463);
nand U46692 (N_46692,N_46442,N_46094);
nor U46693 (N_46693,N_46457,N_46304);
xnor U46694 (N_46694,N_46368,N_46350);
nand U46695 (N_46695,N_46053,N_46283);
or U46696 (N_46696,N_46001,N_46152);
nand U46697 (N_46697,N_46007,N_46081);
nand U46698 (N_46698,N_46186,N_46231);
and U46699 (N_46699,N_46182,N_46292);
nor U46700 (N_46700,N_46207,N_46119);
or U46701 (N_46701,N_46290,N_46377);
nor U46702 (N_46702,N_46380,N_46202);
nor U46703 (N_46703,N_46184,N_46453);
and U46704 (N_46704,N_46449,N_46036);
or U46705 (N_46705,N_46225,N_46151);
or U46706 (N_46706,N_46320,N_46008);
xor U46707 (N_46707,N_46162,N_46060);
and U46708 (N_46708,N_46205,N_46058);
nor U46709 (N_46709,N_46172,N_46092);
and U46710 (N_46710,N_46450,N_46495);
nand U46711 (N_46711,N_46489,N_46264);
xnor U46712 (N_46712,N_46352,N_46403);
or U46713 (N_46713,N_46043,N_46074);
nor U46714 (N_46714,N_46226,N_46265);
xnor U46715 (N_46715,N_46015,N_46108);
nor U46716 (N_46716,N_46248,N_46431);
or U46717 (N_46717,N_46144,N_46303);
and U46718 (N_46718,N_46142,N_46411);
or U46719 (N_46719,N_46325,N_46246);
or U46720 (N_46720,N_46173,N_46327);
nand U46721 (N_46721,N_46342,N_46289);
or U46722 (N_46722,N_46452,N_46286);
nor U46723 (N_46723,N_46175,N_46106);
or U46724 (N_46724,N_46229,N_46482);
nor U46725 (N_46725,N_46480,N_46109);
xnor U46726 (N_46726,N_46090,N_46427);
or U46727 (N_46727,N_46113,N_46218);
xnor U46728 (N_46728,N_46321,N_46212);
nor U46729 (N_46729,N_46019,N_46465);
nor U46730 (N_46730,N_46078,N_46096);
and U46731 (N_46731,N_46413,N_46461);
and U46732 (N_46732,N_46235,N_46309);
nor U46733 (N_46733,N_46485,N_46243);
xnor U46734 (N_46734,N_46385,N_46129);
or U46735 (N_46735,N_46253,N_46326);
or U46736 (N_46736,N_46448,N_46470);
xnor U46737 (N_46737,N_46432,N_46040);
xor U46738 (N_46738,N_46255,N_46085);
or U46739 (N_46739,N_46469,N_46285);
or U46740 (N_46740,N_46003,N_46191);
xor U46741 (N_46741,N_46104,N_46267);
nor U46742 (N_46742,N_46014,N_46110);
and U46743 (N_46743,N_46361,N_46351);
nor U46744 (N_46744,N_46107,N_46132);
xnor U46745 (N_46745,N_46478,N_46381);
or U46746 (N_46746,N_46297,N_46257);
nor U46747 (N_46747,N_46405,N_46098);
xnor U46748 (N_46748,N_46317,N_46396);
and U46749 (N_46749,N_46138,N_46228);
xnor U46750 (N_46750,N_46343,N_46230);
xnor U46751 (N_46751,N_46124,N_46325);
xnor U46752 (N_46752,N_46349,N_46456);
and U46753 (N_46753,N_46295,N_46054);
and U46754 (N_46754,N_46416,N_46144);
nand U46755 (N_46755,N_46196,N_46069);
xor U46756 (N_46756,N_46498,N_46281);
xnor U46757 (N_46757,N_46439,N_46025);
nand U46758 (N_46758,N_46473,N_46070);
and U46759 (N_46759,N_46432,N_46025);
nor U46760 (N_46760,N_46411,N_46178);
nor U46761 (N_46761,N_46207,N_46126);
and U46762 (N_46762,N_46471,N_46313);
and U46763 (N_46763,N_46475,N_46357);
nor U46764 (N_46764,N_46236,N_46203);
nor U46765 (N_46765,N_46404,N_46288);
or U46766 (N_46766,N_46394,N_46283);
nor U46767 (N_46767,N_46370,N_46306);
and U46768 (N_46768,N_46193,N_46079);
xnor U46769 (N_46769,N_46323,N_46075);
xor U46770 (N_46770,N_46162,N_46433);
nand U46771 (N_46771,N_46266,N_46422);
nand U46772 (N_46772,N_46013,N_46102);
nand U46773 (N_46773,N_46059,N_46068);
and U46774 (N_46774,N_46035,N_46098);
nor U46775 (N_46775,N_46155,N_46076);
nor U46776 (N_46776,N_46171,N_46350);
xnor U46777 (N_46777,N_46334,N_46349);
nor U46778 (N_46778,N_46229,N_46416);
nor U46779 (N_46779,N_46206,N_46405);
or U46780 (N_46780,N_46053,N_46018);
nor U46781 (N_46781,N_46114,N_46446);
xnor U46782 (N_46782,N_46295,N_46083);
nand U46783 (N_46783,N_46062,N_46216);
or U46784 (N_46784,N_46308,N_46161);
or U46785 (N_46785,N_46411,N_46215);
or U46786 (N_46786,N_46341,N_46400);
xnor U46787 (N_46787,N_46041,N_46424);
nand U46788 (N_46788,N_46494,N_46073);
and U46789 (N_46789,N_46166,N_46217);
nor U46790 (N_46790,N_46448,N_46406);
and U46791 (N_46791,N_46023,N_46358);
and U46792 (N_46792,N_46025,N_46488);
xor U46793 (N_46793,N_46229,N_46248);
xnor U46794 (N_46794,N_46488,N_46001);
or U46795 (N_46795,N_46298,N_46137);
or U46796 (N_46796,N_46456,N_46072);
and U46797 (N_46797,N_46096,N_46265);
or U46798 (N_46798,N_46439,N_46255);
and U46799 (N_46799,N_46257,N_46045);
or U46800 (N_46800,N_46491,N_46147);
or U46801 (N_46801,N_46065,N_46413);
nor U46802 (N_46802,N_46403,N_46007);
xnor U46803 (N_46803,N_46485,N_46126);
xnor U46804 (N_46804,N_46227,N_46351);
or U46805 (N_46805,N_46065,N_46416);
nand U46806 (N_46806,N_46225,N_46211);
nand U46807 (N_46807,N_46327,N_46199);
xnor U46808 (N_46808,N_46039,N_46496);
and U46809 (N_46809,N_46007,N_46005);
nand U46810 (N_46810,N_46049,N_46354);
or U46811 (N_46811,N_46262,N_46260);
nand U46812 (N_46812,N_46435,N_46207);
xnor U46813 (N_46813,N_46395,N_46405);
or U46814 (N_46814,N_46143,N_46082);
nand U46815 (N_46815,N_46495,N_46406);
nor U46816 (N_46816,N_46372,N_46459);
and U46817 (N_46817,N_46334,N_46093);
and U46818 (N_46818,N_46321,N_46485);
xnor U46819 (N_46819,N_46096,N_46076);
nand U46820 (N_46820,N_46242,N_46215);
nand U46821 (N_46821,N_46111,N_46185);
xnor U46822 (N_46822,N_46216,N_46160);
or U46823 (N_46823,N_46159,N_46305);
nand U46824 (N_46824,N_46181,N_46231);
nand U46825 (N_46825,N_46223,N_46293);
or U46826 (N_46826,N_46261,N_46268);
or U46827 (N_46827,N_46125,N_46032);
or U46828 (N_46828,N_46205,N_46200);
xor U46829 (N_46829,N_46171,N_46088);
or U46830 (N_46830,N_46091,N_46175);
xor U46831 (N_46831,N_46317,N_46131);
xor U46832 (N_46832,N_46125,N_46223);
and U46833 (N_46833,N_46187,N_46241);
or U46834 (N_46834,N_46457,N_46255);
nand U46835 (N_46835,N_46249,N_46222);
and U46836 (N_46836,N_46280,N_46255);
nor U46837 (N_46837,N_46150,N_46235);
nand U46838 (N_46838,N_46386,N_46166);
or U46839 (N_46839,N_46497,N_46012);
nor U46840 (N_46840,N_46324,N_46401);
nand U46841 (N_46841,N_46114,N_46045);
nor U46842 (N_46842,N_46138,N_46151);
or U46843 (N_46843,N_46487,N_46291);
or U46844 (N_46844,N_46428,N_46249);
and U46845 (N_46845,N_46369,N_46417);
or U46846 (N_46846,N_46122,N_46190);
or U46847 (N_46847,N_46386,N_46438);
xnor U46848 (N_46848,N_46123,N_46489);
nand U46849 (N_46849,N_46142,N_46066);
xnor U46850 (N_46850,N_46426,N_46239);
xor U46851 (N_46851,N_46263,N_46021);
nor U46852 (N_46852,N_46070,N_46170);
nand U46853 (N_46853,N_46489,N_46259);
nand U46854 (N_46854,N_46179,N_46371);
xnor U46855 (N_46855,N_46368,N_46192);
xor U46856 (N_46856,N_46144,N_46097);
nor U46857 (N_46857,N_46295,N_46064);
and U46858 (N_46858,N_46079,N_46304);
xor U46859 (N_46859,N_46483,N_46255);
nor U46860 (N_46860,N_46380,N_46431);
xor U46861 (N_46861,N_46418,N_46351);
xnor U46862 (N_46862,N_46054,N_46495);
nand U46863 (N_46863,N_46129,N_46315);
nand U46864 (N_46864,N_46164,N_46031);
and U46865 (N_46865,N_46451,N_46326);
nand U46866 (N_46866,N_46192,N_46455);
or U46867 (N_46867,N_46329,N_46498);
and U46868 (N_46868,N_46471,N_46319);
xnor U46869 (N_46869,N_46002,N_46125);
nor U46870 (N_46870,N_46455,N_46322);
xor U46871 (N_46871,N_46256,N_46184);
nor U46872 (N_46872,N_46328,N_46017);
nand U46873 (N_46873,N_46085,N_46050);
xnor U46874 (N_46874,N_46473,N_46213);
nand U46875 (N_46875,N_46427,N_46121);
or U46876 (N_46876,N_46375,N_46004);
nor U46877 (N_46877,N_46104,N_46360);
or U46878 (N_46878,N_46472,N_46291);
xnor U46879 (N_46879,N_46162,N_46211);
nand U46880 (N_46880,N_46439,N_46094);
nor U46881 (N_46881,N_46487,N_46349);
and U46882 (N_46882,N_46436,N_46287);
nor U46883 (N_46883,N_46389,N_46011);
or U46884 (N_46884,N_46133,N_46323);
or U46885 (N_46885,N_46006,N_46336);
or U46886 (N_46886,N_46226,N_46188);
xor U46887 (N_46887,N_46158,N_46232);
nor U46888 (N_46888,N_46443,N_46053);
or U46889 (N_46889,N_46434,N_46186);
nand U46890 (N_46890,N_46208,N_46291);
and U46891 (N_46891,N_46253,N_46318);
xnor U46892 (N_46892,N_46183,N_46106);
nand U46893 (N_46893,N_46188,N_46497);
and U46894 (N_46894,N_46065,N_46415);
or U46895 (N_46895,N_46296,N_46431);
and U46896 (N_46896,N_46434,N_46311);
and U46897 (N_46897,N_46046,N_46192);
nand U46898 (N_46898,N_46037,N_46483);
nand U46899 (N_46899,N_46057,N_46481);
or U46900 (N_46900,N_46194,N_46432);
or U46901 (N_46901,N_46362,N_46258);
and U46902 (N_46902,N_46032,N_46256);
or U46903 (N_46903,N_46456,N_46298);
nor U46904 (N_46904,N_46160,N_46258);
xnor U46905 (N_46905,N_46012,N_46212);
or U46906 (N_46906,N_46274,N_46288);
or U46907 (N_46907,N_46494,N_46397);
or U46908 (N_46908,N_46470,N_46351);
nor U46909 (N_46909,N_46054,N_46444);
xnor U46910 (N_46910,N_46256,N_46348);
nor U46911 (N_46911,N_46390,N_46059);
or U46912 (N_46912,N_46149,N_46478);
or U46913 (N_46913,N_46031,N_46152);
xor U46914 (N_46914,N_46183,N_46005);
or U46915 (N_46915,N_46065,N_46004);
xnor U46916 (N_46916,N_46117,N_46229);
or U46917 (N_46917,N_46389,N_46321);
or U46918 (N_46918,N_46494,N_46027);
or U46919 (N_46919,N_46272,N_46128);
or U46920 (N_46920,N_46205,N_46170);
and U46921 (N_46921,N_46290,N_46329);
and U46922 (N_46922,N_46352,N_46160);
nor U46923 (N_46923,N_46201,N_46329);
nor U46924 (N_46924,N_46316,N_46093);
and U46925 (N_46925,N_46055,N_46489);
and U46926 (N_46926,N_46374,N_46356);
or U46927 (N_46927,N_46368,N_46206);
and U46928 (N_46928,N_46253,N_46255);
or U46929 (N_46929,N_46256,N_46037);
nand U46930 (N_46930,N_46367,N_46222);
xnor U46931 (N_46931,N_46390,N_46350);
nor U46932 (N_46932,N_46049,N_46484);
and U46933 (N_46933,N_46393,N_46449);
and U46934 (N_46934,N_46149,N_46013);
and U46935 (N_46935,N_46481,N_46340);
xnor U46936 (N_46936,N_46150,N_46084);
and U46937 (N_46937,N_46397,N_46091);
xor U46938 (N_46938,N_46482,N_46364);
nand U46939 (N_46939,N_46179,N_46135);
xnor U46940 (N_46940,N_46251,N_46088);
xor U46941 (N_46941,N_46176,N_46060);
and U46942 (N_46942,N_46266,N_46020);
xor U46943 (N_46943,N_46408,N_46008);
nand U46944 (N_46944,N_46341,N_46145);
and U46945 (N_46945,N_46344,N_46133);
nand U46946 (N_46946,N_46188,N_46117);
and U46947 (N_46947,N_46342,N_46274);
or U46948 (N_46948,N_46471,N_46381);
and U46949 (N_46949,N_46084,N_46033);
nand U46950 (N_46950,N_46302,N_46124);
or U46951 (N_46951,N_46257,N_46067);
xor U46952 (N_46952,N_46477,N_46409);
or U46953 (N_46953,N_46336,N_46024);
nor U46954 (N_46954,N_46240,N_46191);
nor U46955 (N_46955,N_46429,N_46191);
xor U46956 (N_46956,N_46038,N_46483);
xor U46957 (N_46957,N_46032,N_46079);
xnor U46958 (N_46958,N_46404,N_46287);
and U46959 (N_46959,N_46029,N_46032);
and U46960 (N_46960,N_46267,N_46439);
xor U46961 (N_46961,N_46361,N_46344);
xor U46962 (N_46962,N_46015,N_46463);
or U46963 (N_46963,N_46416,N_46186);
nor U46964 (N_46964,N_46070,N_46106);
and U46965 (N_46965,N_46018,N_46352);
or U46966 (N_46966,N_46364,N_46314);
nor U46967 (N_46967,N_46353,N_46417);
nor U46968 (N_46968,N_46075,N_46363);
xnor U46969 (N_46969,N_46396,N_46207);
and U46970 (N_46970,N_46487,N_46402);
nor U46971 (N_46971,N_46342,N_46238);
or U46972 (N_46972,N_46244,N_46044);
and U46973 (N_46973,N_46263,N_46430);
xnor U46974 (N_46974,N_46110,N_46007);
nand U46975 (N_46975,N_46028,N_46243);
nand U46976 (N_46976,N_46214,N_46289);
xnor U46977 (N_46977,N_46205,N_46469);
nor U46978 (N_46978,N_46146,N_46072);
and U46979 (N_46979,N_46015,N_46062);
or U46980 (N_46980,N_46167,N_46214);
nand U46981 (N_46981,N_46454,N_46305);
or U46982 (N_46982,N_46054,N_46451);
nor U46983 (N_46983,N_46251,N_46245);
and U46984 (N_46984,N_46469,N_46408);
nand U46985 (N_46985,N_46134,N_46362);
or U46986 (N_46986,N_46113,N_46099);
nor U46987 (N_46987,N_46380,N_46460);
and U46988 (N_46988,N_46100,N_46470);
or U46989 (N_46989,N_46303,N_46048);
and U46990 (N_46990,N_46182,N_46252);
and U46991 (N_46991,N_46230,N_46237);
or U46992 (N_46992,N_46261,N_46169);
nand U46993 (N_46993,N_46042,N_46462);
xnor U46994 (N_46994,N_46127,N_46051);
xor U46995 (N_46995,N_46039,N_46366);
or U46996 (N_46996,N_46416,N_46434);
xor U46997 (N_46997,N_46323,N_46301);
or U46998 (N_46998,N_46021,N_46055);
and U46999 (N_46999,N_46068,N_46269);
nand U47000 (N_47000,N_46755,N_46741);
nand U47001 (N_47001,N_46659,N_46635);
and U47002 (N_47002,N_46670,N_46545);
nor U47003 (N_47003,N_46607,N_46542);
and U47004 (N_47004,N_46900,N_46901);
nor U47005 (N_47005,N_46722,N_46743);
and U47006 (N_47006,N_46618,N_46819);
xnor U47007 (N_47007,N_46947,N_46798);
and U47008 (N_47008,N_46753,N_46522);
xnor U47009 (N_47009,N_46658,N_46966);
and U47010 (N_47010,N_46802,N_46525);
or U47011 (N_47011,N_46827,N_46527);
or U47012 (N_47012,N_46533,N_46984);
or U47013 (N_47013,N_46588,N_46976);
and U47014 (N_47014,N_46895,N_46694);
or U47015 (N_47015,N_46597,N_46509);
nor U47016 (N_47016,N_46760,N_46752);
nand U47017 (N_47017,N_46929,N_46845);
xnor U47018 (N_47018,N_46631,N_46651);
and U47019 (N_47019,N_46706,N_46595);
xnor U47020 (N_47020,N_46803,N_46555);
nand U47021 (N_47021,N_46603,N_46678);
xnor U47022 (N_47022,N_46933,N_46645);
xor U47023 (N_47023,N_46530,N_46677);
nand U47024 (N_47024,N_46875,N_46785);
or U47025 (N_47025,N_46911,N_46728);
and U47026 (N_47026,N_46746,N_46705);
xor U47027 (N_47027,N_46890,N_46758);
or U47028 (N_47028,N_46671,N_46896);
and U47029 (N_47029,N_46503,N_46647);
nor U47030 (N_47030,N_46872,N_46546);
nand U47031 (N_47031,N_46638,N_46903);
or U47032 (N_47032,N_46809,N_46849);
nor U47033 (N_47033,N_46780,N_46717);
nand U47034 (N_47034,N_46855,N_46958);
and U47035 (N_47035,N_46637,N_46702);
nor U47036 (N_47036,N_46990,N_46816);
nor U47037 (N_47037,N_46774,N_46939);
or U47038 (N_47038,N_46766,N_46515);
nand U47039 (N_47039,N_46615,N_46520);
and U47040 (N_47040,N_46943,N_46910);
or U47041 (N_47041,N_46871,N_46569);
nand U47042 (N_47042,N_46844,N_46514);
or U47043 (N_47043,N_46862,N_46822);
nor U47044 (N_47044,N_46719,N_46586);
xnor U47045 (N_47045,N_46781,N_46869);
nand U47046 (N_47046,N_46674,N_46796);
nor U47047 (N_47047,N_46624,N_46642);
or U47048 (N_47048,N_46567,N_46812);
and U47049 (N_47049,N_46544,N_46927);
or U47050 (N_47050,N_46581,N_46662);
xnor U47051 (N_47051,N_46925,N_46600);
nor U47052 (N_47052,N_46557,N_46536);
nand U47053 (N_47053,N_46561,N_46593);
or U47054 (N_47054,N_46696,N_46757);
nor U47055 (N_47055,N_46777,N_46936);
or U47056 (N_47056,N_46949,N_46516);
xnor U47057 (N_47057,N_46634,N_46535);
or U47058 (N_47058,N_46742,N_46873);
nor U47059 (N_47059,N_46981,N_46721);
xnor U47060 (N_47060,N_46937,N_46710);
xnor U47061 (N_47061,N_46504,N_46711);
xor U47062 (N_47062,N_46661,N_46842);
xnor U47063 (N_47063,N_46913,N_46926);
and U47064 (N_47064,N_46889,N_46799);
or U47065 (N_47065,N_46616,N_46897);
nand U47066 (N_47066,N_46578,N_46541);
nand U47067 (N_47067,N_46598,N_46914);
xor U47068 (N_47068,N_46679,N_46953);
and U47069 (N_47069,N_46640,N_46693);
or U47070 (N_47070,N_46614,N_46830);
nor U47071 (N_47071,N_46532,N_46859);
nor U47072 (N_47072,N_46992,N_46921);
xnor U47073 (N_47073,N_46691,N_46553);
or U47074 (N_47074,N_46979,N_46865);
xnor U47075 (N_47075,N_46843,N_46863);
or U47076 (N_47076,N_46905,N_46962);
nand U47077 (N_47077,N_46629,N_46681);
or U47078 (N_47078,N_46539,N_46575);
xnor U47079 (N_47079,N_46619,N_46594);
nor U47080 (N_47080,N_46874,N_46831);
nand U47081 (N_47081,N_46762,N_46963);
or U47082 (N_47082,N_46834,N_46519);
or U47083 (N_47083,N_46868,N_46652);
nand U47084 (N_47084,N_46673,N_46825);
and U47085 (N_47085,N_46808,N_46683);
xnor U47086 (N_47086,N_46988,N_46824);
nor U47087 (N_47087,N_46574,N_46997);
nand U47088 (N_47088,N_46771,N_46961);
nor U47089 (N_47089,N_46570,N_46521);
nor U47090 (N_47090,N_46685,N_46818);
or U47091 (N_47091,N_46828,N_46924);
and U47092 (N_47092,N_46931,N_46986);
nor U47093 (N_47093,N_46604,N_46759);
nand U47094 (N_47094,N_46836,N_46582);
xnor U47095 (N_47095,N_46583,N_46712);
nand U47096 (N_47096,N_46622,N_46954);
nand U47097 (N_47097,N_46704,N_46946);
and U47098 (N_47098,N_46589,N_46880);
and U47099 (N_47099,N_46980,N_46568);
or U47100 (N_47100,N_46891,N_46887);
xnor U47101 (N_47101,N_46650,N_46814);
or U47102 (N_47102,N_46633,N_46739);
nor U47103 (N_47103,N_46867,N_46554);
xor U47104 (N_47104,N_46695,N_46754);
or U47105 (N_47105,N_46571,N_46648);
and U47106 (N_47106,N_46860,N_46973);
or U47107 (N_47107,N_46585,N_46592);
nor U47108 (N_47108,N_46787,N_46708);
nor U47109 (N_47109,N_46950,N_46501);
nor U47110 (N_47110,N_46850,N_46686);
nand U47111 (N_47111,N_46821,N_46912);
xnor U47112 (N_47112,N_46538,N_46733);
nand U47113 (N_47113,N_46716,N_46657);
xor U47114 (N_47114,N_46829,N_46602);
nand U47115 (N_47115,N_46632,N_46715);
and U47116 (N_47116,N_46833,N_46587);
nor U47117 (N_47117,N_46566,N_46930);
nand U47118 (N_47118,N_46779,N_46738);
or U47119 (N_47119,N_46641,N_46878);
nor U47120 (N_47120,N_46955,N_46737);
nand U47121 (N_47121,N_46969,N_46885);
and U47122 (N_47122,N_46537,N_46940);
nor U47123 (N_47123,N_46770,N_46944);
xnor U47124 (N_47124,N_46580,N_46894);
and U47125 (N_47125,N_46888,N_46899);
and U47126 (N_47126,N_46551,N_46718);
or U47127 (N_47127,N_46573,N_46881);
nand U47128 (N_47128,N_46701,N_46500);
nand U47129 (N_47129,N_46810,N_46727);
and U47130 (N_47130,N_46982,N_46938);
nor U47131 (N_47131,N_46807,N_46606);
or U47132 (N_47132,N_46639,N_46884);
and U47133 (N_47133,N_46558,N_46666);
nand U47134 (N_47134,N_46791,N_46505);
nand U47135 (N_47135,N_46745,N_46556);
xor U47136 (N_47136,N_46951,N_46934);
and U47137 (N_47137,N_46877,N_46692);
or U47138 (N_47138,N_46960,N_46775);
nor U47139 (N_47139,N_46731,N_46552);
or U47140 (N_47140,N_46627,N_46730);
nor U47141 (N_47141,N_46994,N_46599);
or U47142 (N_47142,N_46841,N_46848);
nor U47143 (N_47143,N_46572,N_46513);
or U47144 (N_47144,N_46703,N_46768);
and U47145 (N_47145,N_46789,N_46999);
nand U47146 (N_47146,N_46655,N_46893);
nand U47147 (N_47147,N_46534,N_46918);
nand U47148 (N_47148,N_46861,N_46676);
xor U47149 (N_47149,N_46653,N_46792);
xnor U47150 (N_47150,N_46610,N_46660);
or U47151 (N_47151,N_46526,N_46735);
and U47152 (N_47152,N_46811,N_46654);
nand U47153 (N_47153,N_46790,N_46776);
xor U47154 (N_47154,N_46548,N_46761);
nand U47155 (N_47155,N_46883,N_46915);
or U47156 (N_47156,N_46511,N_46726);
xor U47157 (N_47157,N_46621,N_46563);
xor U47158 (N_47158,N_46932,N_46856);
nor U47159 (N_47159,N_46613,N_46690);
xor U47160 (N_47160,N_46646,N_46805);
or U47161 (N_47161,N_46916,N_46923);
nor U47162 (N_47162,N_46956,N_46684);
or U47163 (N_47163,N_46508,N_46817);
or U47164 (N_47164,N_46765,N_46784);
nand U47165 (N_47165,N_46920,N_46749);
xor U47166 (N_47166,N_46783,N_46643);
nand U47167 (N_47167,N_46851,N_46797);
xor U47168 (N_47168,N_46700,N_46987);
and U47169 (N_47169,N_46751,N_46769);
nand U47170 (N_47170,N_46750,N_46698);
xor U47171 (N_47171,N_46547,N_46617);
or U47172 (N_47172,N_46709,N_46748);
and U47173 (N_47173,N_46853,N_46531);
and U47174 (N_47174,N_46626,N_46794);
and U47175 (N_47175,N_46996,N_46815);
and U47176 (N_47176,N_46625,N_46879);
nor U47177 (N_47177,N_46724,N_46747);
and U47178 (N_47178,N_46675,N_46736);
or U47179 (N_47179,N_46993,N_46502);
or U47180 (N_47180,N_46506,N_46672);
nor U47181 (N_47181,N_46838,N_46864);
xnor U47182 (N_47182,N_46837,N_46804);
and U47183 (N_47183,N_46876,N_46591);
xor U47184 (N_47184,N_46907,N_46945);
xnor U47185 (N_47185,N_46906,N_46959);
xnor U47186 (N_47186,N_46596,N_46576);
or U47187 (N_47187,N_46935,N_46967);
nand U47188 (N_47188,N_46732,N_46978);
and U47189 (N_47189,N_46782,N_46518);
and U47190 (N_47190,N_46628,N_46763);
nor U47191 (N_47191,N_46565,N_46656);
nor U47192 (N_47192,N_46826,N_46813);
xnor U47193 (N_47193,N_46820,N_46847);
nor U47194 (N_47194,N_46854,N_46697);
or U47195 (N_47195,N_46795,N_46649);
nand U47196 (N_47196,N_46540,N_46975);
xor U47197 (N_47197,N_46744,N_46866);
or U47198 (N_47198,N_46590,N_46840);
nor U47199 (N_47199,N_46584,N_46560);
xor U47200 (N_47200,N_46523,N_46941);
and U47201 (N_47201,N_46852,N_46680);
or U47202 (N_47202,N_46892,N_46965);
and U47203 (N_47203,N_46983,N_46773);
and U47204 (N_47204,N_46507,N_46917);
nor U47205 (N_47205,N_46682,N_46517);
and U47206 (N_47206,N_46524,N_46699);
nor U47207 (N_47207,N_46948,N_46665);
xor U47208 (N_47208,N_46772,N_46786);
and U47209 (N_47209,N_46970,N_46688);
or U47210 (N_47210,N_46577,N_46714);
or U47211 (N_47211,N_46909,N_46922);
xor U47212 (N_47212,N_46964,N_46612);
nand U47213 (N_47213,N_46952,N_46870);
and U47214 (N_47214,N_46974,N_46977);
nand U47215 (N_47215,N_46904,N_46605);
nand U47216 (N_47216,N_46663,N_46971);
nand U47217 (N_47217,N_46902,N_46664);
nor U47218 (N_47218,N_46991,N_46886);
xnor U47219 (N_47219,N_46998,N_46667);
and U47220 (N_47220,N_46644,N_46839);
and U47221 (N_47221,N_46611,N_46549);
nor U47222 (N_47222,N_46767,N_46689);
and U47223 (N_47223,N_46756,N_46630);
nand U47224 (N_47224,N_46942,N_46793);
or U47225 (N_47225,N_46985,N_46668);
or U47226 (N_47226,N_46832,N_46740);
xor U47227 (N_47227,N_46550,N_46636);
and U47228 (N_47228,N_46669,N_46623);
and U47229 (N_47229,N_46919,N_46846);
and U47230 (N_47230,N_46801,N_46725);
nand U47231 (N_47231,N_46972,N_46529);
and U47232 (N_47232,N_46559,N_46609);
or U47233 (N_47233,N_46601,N_46989);
and U47234 (N_47234,N_46857,N_46928);
nand U47235 (N_47235,N_46608,N_46713);
nand U47236 (N_47236,N_46882,N_46564);
and U47237 (N_47237,N_46823,N_46729);
or U47238 (N_47238,N_46720,N_46723);
or U47239 (N_47239,N_46806,N_46579);
nand U47240 (N_47240,N_46898,N_46562);
xor U47241 (N_47241,N_46800,N_46778);
and U47242 (N_47242,N_46543,N_46995);
and U47243 (N_47243,N_46835,N_46687);
nor U47244 (N_47244,N_46512,N_46957);
nand U47245 (N_47245,N_46858,N_46707);
nor U47246 (N_47246,N_46510,N_46788);
or U47247 (N_47247,N_46528,N_46734);
nand U47248 (N_47248,N_46764,N_46620);
nand U47249 (N_47249,N_46968,N_46908);
nand U47250 (N_47250,N_46801,N_46720);
nor U47251 (N_47251,N_46838,N_46765);
and U47252 (N_47252,N_46808,N_46994);
nand U47253 (N_47253,N_46614,N_46682);
nor U47254 (N_47254,N_46772,N_46872);
nor U47255 (N_47255,N_46642,N_46539);
or U47256 (N_47256,N_46722,N_46703);
nand U47257 (N_47257,N_46820,N_46875);
nand U47258 (N_47258,N_46812,N_46528);
xor U47259 (N_47259,N_46874,N_46643);
and U47260 (N_47260,N_46657,N_46998);
xor U47261 (N_47261,N_46501,N_46855);
or U47262 (N_47262,N_46747,N_46901);
nand U47263 (N_47263,N_46883,N_46886);
nand U47264 (N_47264,N_46781,N_46718);
nor U47265 (N_47265,N_46796,N_46669);
and U47266 (N_47266,N_46694,N_46786);
and U47267 (N_47267,N_46606,N_46855);
nor U47268 (N_47268,N_46650,N_46565);
nand U47269 (N_47269,N_46828,N_46913);
or U47270 (N_47270,N_46765,N_46751);
nand U47271 (N_47271,N_46909,N_46669);
nor U47272 (N_47272,N_46635,N_46981);
xnor U47273 (N_47273,N_46732,N_46840);
xnor U47274 (N_47274,N_46674,N_46525);
nand U47275 (N_47275,N_46640,N_46619);
xor U47276 (N_47276,N_46657,N_46626);
nand U47277 (N_47277,N_46529,N_46559);
xor U47278 (N_47278,N_46811,N_46788);
and U47279 (N_47279,N_46729,N_46996);
and U47280 (N_47280,N_46967,N_46949);
or U47281 (N_47281,N_46663,N_46740);
nor U47282 (N_47282,N_46664,N_46665);
and U47283 (N_47283,N_46993,N_46872);
nor U47284 (N_47284,N_46708,N_46869);
nor U47285 (N_47285,N_46541,N_46593);
and U47286 (N_47286,N_46535,N_46982);
or U47287 (N_47287,N_46693,N_46916);
and U47288 (N_47288,N_46575,N_46639);
nor U47289 (N_47289,N_46901,N_46532);
or U47290 (N_47290,N_46692,N_46809);
and U47291 (N_47291,N_46683,N_46924);
and U47292 (N_47292,N_46760,N_46954);
nand U47293 (N_47293,N_46730,N_46561);
xnor U47294 (N_47294,N_46797,N_46641);
nand U47295 (N_47295,N_46674,N_46872);
xor U47296 (N_47296,N_46880,N_46969);
or U47297 (N_47297,N_46713,N_46750);
xnor U47298 (N_47298,N_46684,N_46921);
nor U47299 (N_47299,N_46708,N_46561);
and U47300 (N_47300,N_46664,N_46677);
nand U47301 (N_47301,N_46530,N_46880);
nor U47302 (N_47302,N_46997,N_46791);
nand U47303 (N_47303,N_46629,N_46505);
and U47304 (N_47304,N_46547,N_46957);
or U47305 (N_47305,N_46708,N_46602);
or U47306 (N_47306,N_46639,N_46529);
nand U47307 (N_47307,N_46685,N_46873);
xnor U47308 (N_47308,N_46760,N_46808);
xnor U47309 (N_47309,N_46711,N_46878);
or U47310 (N_47310,N_46953,N_46530);
nand U47311 (N_47311,N_46940,N_46818);
or U47312 (N_47312,N_46830,N_46929);
or U47313 (N_47313,N_46602,N_46685);
or U47314 (N_47314,N_46708,N_46791);
and U47315 (N_47315,N_46683,N_46875);
nand U47316 (N_47316,N_46557,N_46574);
and U47317 (N_47317,N_46756,N_46804);
nor U47318 (N_47318,N_46677,N_46963);
and U47319 (N_47319,N_46631,N_46643);
xor U47320 (N_47320,N_46900,N_46831);
nand U47321 (N_47321,N_46765,N_46831);
and U47322 (N_47322,N_46567,N_46952);
xor U47323 (N_47323,N_46550,N_46876);
xor U47324 (N_47324,N_46883,N_46582);
or U47325 (N_47325,N_46781,N_46505);
nor U47326 (N_47326,N_46748,N_46589);
nor U47327 (N_47327,N_46816,N_46682);
and U47328 (N_47328,N_46523,N_46771);
xnor U47329 (N_47329,N_46711,N_46665);
nor U47330 (N_47330,N_46589,N_46534);
xnor U47331 (N_47331,N_46805,N_46698);
xor U47332 (N_47332,N_46730,N_46855);
and U47333 (N_47333,N_46829,N_46955);
or U47334 (N_47334,N_46611,N_46724);
nor U47335 (N_47335,N_46732,N_46637);
and U47336 (N_47336,N_46560,N_46737);
xor U47337 (N_47337,N_46784,N_46627);
nand U47338 (N_47338,N_46903,N_46820);
or U47339 (N_47339,N_46800,N_46828);
nand U47340 (N_47340,N_46956,N_46742);
nand U47341 (N_47341,N_46933,N_46862);
nor U47342 (N_47342,N_46952,N_46881);
nor U47343 (N_47343,N_46716,N_46500);
nand U47344 (N_47344,N_46701,N_46536);
nand U47345 (N_47345,N_46712,N_46781);
and U47346 (N_47346,N_46718,N_46847);
nor U47347 (N_47347,N_46867,N_46973);
xor U47348 (N_47348,N_46563,N_46983);
or U47349 (N_47349,N_46938,N_46628);
xor U47350 (N_47350,N_46692,N_46638);
nand U47351 (N_47351,N_46626,N_46567);
nand U47352 (N_47352,N_46630,N_46915);
xor U47353 (N_47353,N_46584,N_46595);
nand U47354 (N_47354,N_46561,N_46843);
or U47355 (N_47355,N_46611,N_46754);
nor U47356 (N_47356,N_46734,N_46781);
or U47357 (N_47357,N_46819,N_46546);
nor U47358 (N_47358,N_46735,N_46853);
xor U47359 (N_47359,N_46537,N_46818);
nand U47360 (N_47360,N_46512,N_46660);
xnor U47361 (N_47361,N_46744,N_46758);
nand U47362 (N_47362,N_46975,N_46684);
nand U47363 (N_47363,N_46551,N_46527);
and U47364 (N_47364,N_46571,N_46599);
nand U47365 (N_47365,N_46769,N_46652);
nor U47366 (N_47366,N_46567,N_46902);
nor U47367 (N_47367,N_46999,N_46824);
xor U47368 (N_47368,N_46668,N_46725);
xor U47369 (N_47369,N_46691,N_46838);
and U47370 (N_47370,N_46845,N_46864);
or U47371 (N_47371,N_46988,N_46823);
xnor U47372 (N_47372,N_46571,N_46781);
or U47373 (N_47373,N_46887,N_46509);
nand U47374 (N_47374,N_46650,N_46780);
nor U47375 (N_47375,N_46942,N_46957);
or U47376 (N_47376,N_46959,N_46676);
nor U47377 (N_47377,N_46662,N_46872);
xnor U47378 (N_47378,N_46596,N_46621);
nor U47379 (N_47379,N_46625,N_46662);
xor U47380 (N_47380,N_46888,N_46532);
nand U47381 (N_47381,N_46795,N_46720);
or U47382 (N_47382,N_46579,N_46792);
or U47383 (N_47383,N_46749,N_46559);
nor U47384 (N_47384,N_46741,N_46619);
nand U47385 (N_47385,N_46950,N_46985);
and U47386 (N_47386,N_46628,N_46835);
xnor U47387 (N_47387,N_46704,N_46561);
nand U47388 (N_47388,N_46795,N_46809);
nand U47389 (N_47389,N_46685,N_46618);
nand U47390 (N_47390,N_46640,N_46560);
or U47391 (N_47391,N_46606,N_46614);
and U47392 (N_47392,N_46942,N_46752);
nand U47393 (N_47393,N_46888,N_46603);
xnor U47394 (N_47394,N_46674,N_46557);
nor U47395 (N_47395,N_46742,N_46648);
xnor U47396 (N_47396,N_46730,N_46898);
or U47397 (N_47397,N_46918,N_46780);
or U47398 (N_47398,N_46838,N_46644);
xor U47399 (N_47399,N_46900,N_46745);
nor U47400 (N_47400,N_46799,N_46783);
xnor U47401 (N_47401,N_46742,N_46617);
nand U47402 (N_47402,N_46942,N_46516);
xor U47403 (N_47403,N_46951,N_46745);
nor U47404 (N_47404,N_46973,N_46775);
nand U47405 (N_47405,N_46513,N_46815);
and U47406 (N_47406,N_46548,N_46641);
nand U47407 (N_47407,N_46689,N_46870);
nand U47408 (N_47408,N_46623,N_46676);
xor U47409 (N_47409,N_46774,N_46883);
or U47410 (N_47410,N_46560,N_46736);
or U47411 (N_47411,N_46589,N_46885);
nor U47412 (N_47412,N_46958,N_46687);
xnor U47413 (N_47413,N_46874,N_46912);
nand U47414 (N_47414,N_46812,N_46715);
or U47415 (N_47415,N_46666,N_46806);
and U47416 (N_47416,N_46849,N_46523);
or U47417 (N_47417,N_46750,N_46868);
or U47418 (N_47418,N_46635,N_46876);
xor U47419 (N_47419,N_46791,N_46684);
or U47420 (N_47420,N_46584,N_46664);
nor U47421 (N_47421,N_46831,N_46712);
or U47422 (N_47422,N_46575,N_46934);
xor U47423 (N_47423,N_46762,N_46551);
nor U47424 (N_47424,N_46831,N_46529);
xor U47425 (N_47425,N_46846,N_46586);
nand U47426 (N_47426,N_46514,N_46877);
or U47427 (N_47427,N_46542,N_46509);
or U47428 (N_47428,N_46824,N_46842);
and U47429 (N_47429,N_46664,N_46656);
nand U47430 (N_47430,N_46506,N_46811);
xnor U47431 (N_47431,N_46995,N_46826);
and U47432 (N_47432,N_46934,N_46869);
and U47433 (N_47433,N_46907,N_46880);
xor U47434 (N_47434,N_46971,N_46903);
or U47435 (N_47435,N_46830,N_46908);
nor U47436 (N_47436,N_46566,N_46848);
nor U47437 (N_47437,N_46969,N_46591);
nand U47438 (N_47438,N_46690,N_46906);
nand U47439 (N_47439,N_46928,N_46625);
nor U47440 (N_47440,N_46696,N_46522);
nand U47441 (N_47441,N_46841,N_46721);
and U47442 (N_47442,N_46889,N_46683);
or U47443 (N_47443,N_46634,N_46983);
xnor U47444 (N_47444,N_46657,N_46698);
nand U47445 (N_47445,N_46587,N_46571);
xor U47446 (N_47446,N_46561,N_46844);
nor U47447 (N_47447,N_46868,N_46816);
or U47448 (N_47448,N_46724,N_46798);
nand U47449 (N_47449,N_46661,N_46611);
xnor U47450 (N_47450,N_46887,N_46828);
nor U47451 (N_47451,N_46601,N_46636);
nand U47452 (N_47452,N_46985,N_46634);
or U47453 (N_47453,N_46728,N_46533);
or U47454 (N_47454,N_46623,N_46827);
or U47455 (N_47455,N_46755,N_46990);
nand U47456 (N_47456,N_46535,N_46836);
or U47457 (N_47457,N_46577,N_46725);
nand U47458 (N_47458,N_46870,N_46788);
or U47459 (N_47459,N_46679,N_46581);
or U47460 (N_47460,N_46565,N_46849);
or U47461 (N_47461,N_46620,N_46807);
or U47462 (N_47462,N_46571,N_46915);
nand U47463 (N_47463,N_46672,N_46859);
nand U47464 (N_47464,N_46896,N_46760);
and U47465 (N_47465,N_46690,N_46917);
or U47466 (N_47466,N_46529,N_46593);
or U47467 (N_47467,N_46659,N_46910);
and U47468 (N_47468,N_46557,N_46682);
and U47469 (N_47469,N_46616,N_46965);
nand U47470 (N_47470,N_46686,N_46500);
and U47471 (N_47471,N_46790,N_46838);
or U47472 (N_47472,N_46735,N_46767);
or U47473 (N_47473,N_46552,N_46970);
and U47474 (N_47474,N_46823,N_46597);
nor U47475 (N_47475,N_46978,N_46658);
nand U47476 (N_47476,N_46905,N_46623);
or U47477 (N_47477,N_46876,N_46601);
nor U47478 (N_47478,N_46849,N_46981);
nand U47479 (N_47479,N_46899,N_46584);
nor U47480 (N_47480,N_46919,N_46877);
nand U47481 (N_47481,N_46584,N_46833);
or U47482 (N_47482,N_46766,N_46830);
and U47483 (N_47483,N_46511,N_46596);
xnor U47484 (N_47484,N_46814,N_46794);
nor U47485 (N_47485,N_46795,N_46658);
and U47486 (N_47486,N_46735,N_46729);
nand U47487 (N_47487,N_46758,N_46774);
nand U47488 (N_47488,N_46863,N_46920);
xor U47489 (N_47489,N_46822,N_46972);
and U47490 (N_47490,N_46755,N_46964);
nand U47491 (N_47491,N_46995,N_46638);
and U47492 (N_47492,N_46956,N_46919);
xor U47493 (N_47493,N_46771,N_46904);
or U47494 (N_47494,N_46717,N_46988);
and U47495 (N_47495,N_46523,N_46518);
xor U47496 (N_47496,N_46704,N_46672);
nor U47497 (N_47497,N_46517,N_46886);
and U47498 (N_47498,N_46604,N_46786);
or U47499 (N_47499,N_46513,N_46505);
xnor U47500 (N_47500,N_47338,N_47239);
or U47501 (N_47501,N_47153,N_47390);
xnor U47502 (N_47502,N_47374,N_47137);
nor U47503 (N_47503,N_47087,N_47224);
or U47504 (N_47504,N_47114,N_47093);
or U47505 (N_47505,N_47301,N_47332);
xor U47506 (N_47506,N_47134,N_47179);
and U47507 (N_47507,N_47078,N_47198);
nor U47508 (N_47508,N_47321,N_47013);
nand U47509 (N_47509,N_47185,N_47328);
nor U47510 (N_47510,N_47211,N_47091);
nand U47511 (N_47511,N_47326,N_47496);
xor U47512 (N_47512,N_47381,N_47122);
nand U47513 (N_47513,N_47107,N_47204);
or U47514 (N_47514,N_47424,N_47306);
xor U47515 (N_47515,N_47109,N_47457);
or U47516 (N_47516,N_47043,N_47303);
and U47517 (N_47517,N_47064,N_47040);
nand U47518 (N_47518,N_47044,N_47261);
or U47519 (N_47519,N_47181,N_47408);
nor U47520 (N_47520,N_47150,N_47451);
or U47521 (N_47521,N_47092,N_47106);
and U47522 (N_47522,N_47099,N_47395);
or U47523 (N_47523,N_47489,N_47141);
nor U47524 (N_47524,N_47159,N_47162);
xnor U47525 (N_47525,N_47059,N_47305);
or U47526 (N_47526,N_47254,N_47209);
xnor U47527 (N_47527,N_47431,N_47052);
nor U47528 (N_47528,N_47411,N_47314);
and U47529 (N_47529,N_47005,N_47067);
nand U47530 (N_47530,N_47131,N_47265);
nand U47531 (N_47531,N_47195,N_47017);
nand U47532 (N_47532,N_47001,N_47475);
nand U47533 (N_47533,N_47333,N_47393);
or U47534 (N_47534,N_47278,N_47135);
or U47535 (N_47535,N_47373,N_47351);
nor U47536 (N_47536,N_47484,N_47330);
xor U47537 (N_47537,N_47037,N_47075);
nand U47538 (N_47538,N_47284,N_47046);
or U47539 (N_47539,N_47088,N_47450);
or U47540 (N_47540,N_47383,N_47486);
xor U47541 (N_47541,N_47102,N_47490);
nand U47542 (N_47542,N_47028,N_47363);
or U47543 (N_47543,N_47473,N_47319);
or U47544 (N_47544,N_47245,N_47119);
or U47545 (N_47545,N_47290,N_47167);
nor U47546 (N_47546,N_47325,N_47230);
or U47547 (N_47547,N_47336,N_47125);
nand U47548 (N_47548,N_47487,N_47029);
nand U47549 (N_47549,N_47104,N_47343);
nor U47550 (N_47550,N_47208,N_47292);
nand U47551 (N_47551,N_47060,N_47474);
and U47552 (N_47552,N_47349,N_47334);
and U47553 (N_47553,N_47483,N_47316);
nand U47554 (N_47554,N_47294,N_47112);
and U47555 (N_47555,N_47171,N_47251);
or U47556 (N_47556,N_47323,N_47397);
nand U47557 (N_47557,N_47427,N_47191);
nor U47558 (N_47558,N_47176,N_47024);
or U47559 (N_47559,N_47063,N_47404);
or U47560 (N_47560,N_47173,N_47414);
nand U47561 (N_47561,N_47158,N_47281);
nor U47562 (N_47562,N_47366,N_47000);
or U47563 (N_47563,N_47342,N_47241);
and U47564 (N_47564,N_47187,N_47156);
nor U47565 (N_47565,N_47236,N_47441);
and U47566 (N_47566,N_47468,N_47297);
xnor U47567 (N_47567,N_47493,N_47207);
or U47568 (N_47568,N_47465,N_47377);
nor U47569 (N_47569,N_47481,N_47340);
or U47570 (N_47570,N_47085,N_47276);
xnor U47571 (N_47571,N_47200,N_47497);
and U47572 (N_47572,N_47440,N_47205);
xor U47573 (N_47573,N_47409,N_47249);
xnor U47574 (N_47574,N_47177,N_47433);
xor U47575 (N_47575,N_47152,N_47042);
or U47576 (N_47576,N_47266,N_47247);
nand U47577 (N_47577,N_47006,N_47233);
nor U47578 (N_47578,N_47108,N_47070);
xor U47579 (N_47579,N_47226,N_47391);
or U47580 (N_47580,N_47412,N_47188);
xor U47581 (N_47581,N_47256,N_47053);
nor U47582 (N_47582,N_47380,N_47184);
nor U47583 (N_47583,N_47288,N_47379);
nand U47584 (N_47584,N_47454,N_47300);
nor U47585 (N_47585,N_47094,N_47232);
nor U47586 (N_47586,N_47180,N_47199);
nor U47587 (N_47587,N_47403,N_47304);
nor U47588 (N_47588,N_47136,N_47477);
nor U47589 (N_47589,N_47317,N_47382);
and U47590 (N_47590,N_47215,N_47074);
xor U47591 (N_47591,N_47008,N_47057);
or U47592 (N_47592,N_47169,N_47217);
nor U47593 (N_47593,N_47347,N_47252);
nor U47594 (N_47594,N_47129,N_47161);
or U47595 (N_47595,N_47143,N_47258);
nand U47596 (N_47596,N_47289,N_47105);
or U47597 (N_47597,N_47138,N_47189);
xor U47598 (N_47598,N_47183,N_47234);
nor U47599 (N_47599,N_47058,N_47032);
xor U47600 (N_47600,N_47166,N_47170);
nor U47601 (N_47601,N_47248,N_47011);
nor U47602 (N_47602,N_47010,N_47255);
and U47603 (N_47603,N_47387,N_47375);
nor U47604 (N_47604,N_47268,N_47140);
nand U47605 (N_47605,N_47172,N_47145);
or U47606 (N_47606,N_47160,N_47469);
or U47607 (N_47607,N_47362,N_47313);
nand U47608 (N_47608,N_47429,N_47275);
nand U47609 (N_47609,N_47420,N_47025);
or U47610 (N_47610,N_47163,N_47369);
and U47611 (N_47611,N_47445,N_47022);
nor U47612 (N_47612,N_47360,N_47378);
nand U47613 (N_47613,N_47318,N_47257);
nand U47614 (N_47614,N_47113,N_47376);
or U47615 (N_47615,N_47026,N_47214);
and U47616 (N_47616,N_47045,N_47157);
xor U47617 (N_47617,N_47364,N_47036);
nand U47618 (N_47618,N_47339,N_47421);
and U47619 (N_47619,N_47417,N_47090);
nor U47620 (N_47620,N_47423,N_47110);
nor U47621 (N_47621,N_47485,N_47081);
nor U47622 (N_47622,N_47231,N_47196);
and U47623 (N_47623,N_47186,N_47219);
and U47624 (N_47624,N_47220,N_47461);
xor U47625 (N_47625,N_47126,N_47460);
or U47626 (N_47626,N_47307,N_47470);
nor U47627 (N_47627,N_47324,N_47123);
or U47628 (N_47628,N_47407,N_47020);
nand U47629 (N_47629,N_47050,N_47240);
nor U47630 (N_47630,N_47178,N_47315);
nand U47631 (N_47631,N_47447,N_47353);
nand U47632 (N_47632,N_47021,N_47448);
and U47633 (N_47633,N_47359,N_47410);
or U47634 (N_47634,N_47228,N_47269);
and U47635 (N_47635,N_47435,N_47030);
or U47636 (N_47636,N_47016,N_47154);
xor U47637 (N_47637,N_47415,N_47229);
nand U47638 (N_47638,N_47201,N_47480);
xor U47639 (N_47639,N_47033,N_47210);
or U47640 (N_47640,N_47139,N_47174);
and U47641 (N_47641,N_47462,N_47133);
and U47642 (N_47642,N_47388,N_47100);
and U47643 (N_47643,N_47371,N_47293);
or U47644 (N_47644,N_47452,N_47331);
or U47645 (N_47645,N_47309,N_47055);
xnor U47646 (N_47646,N_47002,N_47368);
nor U47647 (N_47647,N_47443,N_47132);
nand U47648 (N_47648,N_47068,N_47413);
nor U47649 (N_47649,N_47216,N_47270);
nor U47650 (N_47650,N_47066,N_47308);
nor U47651 (N_47651,N_47422,N_47384);
nor U47652 (N_47652,N_47392,N_47295);
nor U47653 (N_47653,N_47048,N_47164);
and U47654 (N_47654,N_47147,N_47206);
nand U47655 (N_47655,N_47335,N_47399);
xor U47656 (N_47656,N_47494,N_47083);
or U47657 (N_47657,N_47287,N_47047);
nand U47658 (N_47658,N_47009,N_47111);
nor U47659 (N_47659,N_47004,N_47182);
and U47660 (N_47660,N_47076,N_47434);
nand U47661 (N_47661,N_47069,N_47051);
and U47662 (N_47662,N_47014,N_47348);
and U47663 (N_47663,N_47498,N_47244);
nand U47664 (N_47664,N_47262,N_47466);
nand U47665 (N_47665,N_47367,N_47175);
or U47666 (N_47666,N_47296,N_47401);
xnor U47667 (N_47667,N_47488,N_47130);
nor U47668 (N_47668,N_47283,N_47225);
or U47669 (N_47669,N_47322,N_47235);
nor U47670 (N_47670,N_47355,N_47432);
nand U47671 (N_47671,N_47003,N_47472);
or U47672 (N_47672,N_47405,N_47015);
or U47673 (N_47673,N_47459,N_47344);
xor U47674 (N_47674,N_47436,N_47142);
nor U47675 (N_47675,N_47389,N_47400);
nor U47676 (N_47676,N_47192,N_47084);
nand U47677 (N_47677,N_47082,N_47077);
xnor U47678 (N_47678,N_47065,N_47385);
nor U47679 (N_47679,N_47213,N_47190);
nor U47680 (N_47680,N_47264,N_47345);
nor U47681 (N_47681,N_47416,N_47073);
nor U47682 (N_47682,N_47212,N_47223);
nor U47683 (N_47683,N_47482,N_47193);
nand U47684 (N_47684,N_47118,N_47027);
or U47685 (N_47685,N_47280,N_47124);
nand U47686 (N_47686,N_47194,N_47372);
and U47687 (N_47687,N_47341,N_47128);
and U47688 (N_47688,N_47458,N_47467);
xnor U47689 (N_47689,N_47165,N_47430);
nor U47690 (N_47690,N_47272,N_47444);
nand U47691 (N_47691,N_47253,N_47035);
nor U47692 (N_47692,N_47311,N_47034);
nand U47693 (N_47693,N_47079,N_47428);
nor U47694 (N_47694,N_47398,N_47273);
and U47695 (N_47695,N_47054,N_47394);
or U47696 (N_47696,N_47365,N_47056);
and U47697 (N_47697,N_47396,N_47476);
nor U47698 (N_47698,N_47302,N_47438);
nor U47699 (N_47699,N_47495,N_47464);
nand U47700 (N_47700,N_47049,N_47298);
nor U47701 (N_47701,N_47116,N_47149);
xnor U47702 (N_47702,N_47097,N_47012);
or U47703 (N_47703,N_47120,N_47061);
nand U47704 (N_47704,N_47243,N_47146);
and U47705 (N_47705,N_47471,N_47267);
or U47706 (N_47706,N_47098,N_47115);
nor U47707 (N_47707,N_47019,N_47449);
nor U47708 (N_47708,N_47437,N_47031);
xnor U47709 (N_47709,N_47168,N_47299);
nor U47710 (N_47710,N_47221,N_47279);
nand U47711 (N_47711,N_47463,N_47023);
or U47712 (N_47712,N_47039,N_47453);
and U47713 (N_47713,N_47337,N_47260);
or U47714 (N_47714,N_47426,N_47442);
nand U47715 (N_47715,N_47358,N_47203);
and U47716 (N_47716,N_47096,N_47080);
nand U47717 (N_47717,N_47117,N_47346);
nor U47718 (N_47718,N_47499,N_47478);
nand U47719 (N_47719,N_47062,N_47386);
and U47720 (N_47720,N_47439,N_47222);
nor U47721 (N_47721,N_47148,N_47327);
or U47722 (N_47722,N_47312,N_47350);
xnor U47723 (N_47723,N_47356,N_47018);
or U47724 (N_47724,N_47286,N_47038);
xor U47725 (N_47725,N_47227,N_47041);
or U47726 (N_47726,N_47357,N_47250);
or U47727 (N_47727,N_47086,N_47151);
or U47728 (N_47728,N_47071,N_47202);
nand U47729 (N_47729,N_47418,N_47446);
nand U47730 (N_47730,N_47237,N_47456);
and U47731 (N_47731,N_47361,N_47007);
or U47732 (N_47732,N_47419,N_47277);
xor U47733 (N_47733,N_47491,N_47072);
nand U47734 (N_47734,N_47089,N_47274);
nand U47735 (N_47735,N_47354,N_47329);
and U47736 (N_47736,N_47320,N_47282);
or U47737 (N_47737,N_47259,N_47492);
xor U47738 (N_47738,N_47121,N_47197);
nor U47739 (N_47739,N_47238,N_47455);
xnor U47740 (N_47740,N_47144,N_47406);
or U47741 (N_47741,N_47479,N_47271);
nand U47742 (N_47742,N_47103,N_47352);
xnor U47743 (N_47743,N_47127,N_47095);
nand U47744 (N_47744,N_47402,N_47101);
and U47745 (N_47745,N_47155,N_47246);
nor U47746 (N_47746,N_47425,N_47242);
nand U47747 (N_47747,N_47263,N_47310);
xor U47748 (N_47748,N_47218,N_47285);
nor U47749 (N_47749,N_47370,N_47291);
and U47750 (N_47750,N_47058,N_47479);
nor U47751 (N_47751,N_47117,N_47358);
or U47752 (N_47752,N_47002,N_47167);
xor U47753 (N_47753,N_47264,N_47266);
and U47754 (N_47754,N_47483,N_47269);
nor U47755 (N_47755,N_47395,N_47063);
and U47756 (N_47756,N_47397,N_47377);
or U47757 (N_47757,N_47135,N_47246);
xor U47758 (N_47758,N_47281,N_47084);
nor U47759 (N_47759,N_47300,N_47436);
nor U47760 (N_47760,N_47193,N_47198);
nor U47761 (N_47761,N_47394,N_47091);
or U47762 (N_47762,N_47285,N_47324);
or U47763 (N_47763,N_47121,N_47357);
nand U47764 (N_47764,N_47405,N_47489);
nor U47765 (N_47765,N_47100,N_47138);
xor U47766 (N_47766,N_47343,N_47306);
nand U47767 (N_47767,N_47490,N_47387);
or U47768 (N_47768,N_47048,N_47170);
xor U47769 (N_47769,N_47200,N_47069);
nand U47770 (N_47770,N_47421,N_47431);
nor U47771 (N_47771,N_47237,N_47247);
xor U47772 (N_47772,N_47212,N_47424);
or U47773 (N_47773,N_47105,N_47135);
nor U47774 (N_47774,N_47432,N_47393);
and U47775 (N_47775,N_47070,N_47457);
and U47776 (N_47776,N_47467,N_47014);
and U47777 (N_47777,N_47112,N_47286);
xnor U47778 (N_47778,N_47327,N_47296);
nand U47779 (N_47779,N_47385,N_47014);
or U47780 (N_47780,N_47271,N_47319);
xor U47781 (N_47781,N_47476,N_47067);
nand U47782 (N_47782,N_47335,N_47073);
xnor U47783 (N_47783,N_47270,N_47224);
and U47784 (N_47784,N_47202,N_47209);
and U47785 (N_47785,N_47492,N_47413);
nand U47786 (N_47786,N_47302,N_47072);
or U47787 (N_47787,N_47299,N_47329);
nand U47788 (N_47788,N_47173,N_47345);
or U47789 (N_47789,N_47490,N_47298);
nand U47790 (N_47790,N_47449,N_47041);
nand U47791 (N_47791,N_47475,N_47497);
or U47792 (N_47792,N_47106,N_47147);
nor U47793 (N_47793,N_47081,N_47006);
nand U47794 (N_47794,N_47220,N_47103);
and U47795 (N_47795,N_47163,N_47064);
and U47796 (N_47796,N_47140,N_47163);
xor U47797 (N_47797,N_47292,N_47003);
and U47798 (N_47798,N_47319,N_47302);
and U47799 (N_47799,N_47373,N_47053);
or U47800 (N_47800,N_47081,N_47088);
nor U47801 (N_47801,N_47006,N_47091);
and U47802 (N_47802,N_47176,N_47396);
or U47803 (N_47803,N_47150,N_47278);
nor U47804 (N_47804,N_47112,N_47299);
and U47805 (N_47805,N_47057,N_47163);
and U47806 (N_47806,N_47437,N_47062);
xnor U47807 (N_47807,N_47491,N_47027);
xnor U47808 (N_47808,N_47437,N_47250);
nand U47809 (N_47809,N_47309,N_47225);
and U47810 (N_47810,N_47250,N_47201);
nand U47811 (N_47811,N_47126,N_47331);
and U47812 (N_47812,N_47417,N_47380);
xor U47813 (N_47813,N_47212,N_47018);
xor U47814 (N_47814,N_47011,N_47393);
nand U47815 (N_47815,N_47327,N_47008);
or U47816 (N_47816,N_47003,N_47340);
or U47817 (N_47817,N_47128,N_47079);
xor U47818 (N_47818,N_47137,N_47261);
nor U47819 (N_47819,N_47471,N_47465);
nand U47820 (N_47820,N_47466,N_47430);
nor U47821 (N_47821,N_47224,N_47001);
xor U47822 (N_47822,N_47226,N_47012);
and U47823 (N_47823,N_47471,N_47187);
nand U47824 (N_47824,N_47391,N_47408);
nor U47825 (N_47825,N_47132,N_47112);
or U47826 (N_47826,N_47240,N_47395);
nor U47827 (N_47827,N_47273,N_47356);
or U47828 (N_47828,N_47228,N_47222);
nand U47829 (N_47829,N_47014,N_47462);
or U47830 (N_47830,N_47421,N_47348);
or U47831 (N_47831,N_47106,N_47442);
nor U47832 (N_47832,N_47238,N_47045);
xor U47833 (N_47833,N_47298,N_47014);
xnor U47834 (N_47834,N_47416,N_47295);
and U47835 (N_47835,N_47472,N_47049);
nand U47836 (N_47836,N_47491,N_47033);
xnor U47837 (N_47837,N_47268,N_47296);
nand U47838 (N_47838,N_47350,N_47370);
xnor U47839 (N_47839,N_47180,N_47314);
nor U47840 (N_47840,N_47422,N_47458);
nor U47841 (N_47841,N_47223,N_47407);
or U47842 (N_47842,N_47291,N_47269);
nand U47843 (N_47843,N_47139,N_47285);
xnor U47844 (N_47844,N_47105,N_47309);
or U47845 (N_47845,N_47421,N_47315);
nand U47846 (N_47846,N_47307,N_47032);
and U47847 (N_47847,N_47263,N_47433);
xor U47848 (N_47848,N_47191,N_47167);
nand U47849 (N_47849,N_47263,N_47052);
nand U47850 (N_47850,N_47232,N_47322);
and U47851 (N_47851,N_47223,N_47051);
and U47852 (N_47852,N_47157,N_47076);
or U47853 (N_47853,N_47266,N_47440);
nor U47854 (N_47854,N_47055,N_47071);
or U47855 (N_47855,N_47134,N_47237);
nor U47856 (N_47856,N_47266,N_47432);
and U47857 (N_47857,N_47047,N_47061);
and U47858 (N_47858,N_47015,N_47071);
nor U47859 (N_47859,N_47127,N_47122);
nand U47860 (N_47860,N_47168,N_47096);
xnor U47861 (N_47861,N_47196,N_47193);
xor U47862 (N_47862,N_47451,N_47013);
and U47863 (N_47863,N_47047,N_47170);
nor U47864 (N_47864,N_47144,N_47346);
nand U47865 (N_47865,N_47129,N_47402);
or U47866 (N_47866,N_47301,N_47434);
and U47867 (N_47867,N_47096,N_47077);
and U47868 (N_47868,N_47415,N_47261);
nand U47869 (N_47869,N_47426,N_47109);
nand U47870 (N_47870,N_47105,N_47131);
nand U47871 (N_47871,N_47225,N_47032);
and U47872 (N_47872,N_47187,N_47415);
nor U47873 (N_47873,N_47458,N_47231);
nand U47874 (N_47874,N_47201,N_47228);
xnor U47875 (N_47875,N_47142,N_47317);
or U47876 (N_47876,N_47235,N_47383);
or U47877 (N_47877,N_47498,N_47211);
or U47878 (N_47878,N_47095,N_47497);
or U47879 (N_47879,N_47386,N_47136);
nor U47880 (N_47880,N_47191,N_47310);
nand U47881 (N_47881,N_47217,N_47133);
nand U47882 (N_47882,N_47390,N_47132);
or U47883 (N_47883,N_47091,N_47313);
nor U47884 (N_47884,N_47308,N_47100);
xor U47885 (N_47885,N_47107,N_47135);
or U47886 (N_47886,N_47447,N_47440);
nor U47887 (N_47887,N_47166,N_47182);
nor U47888 (N_47888,N_47164,N_47149);
or U47889 (N_47889,N_47319,N_47318);
xnor U47890 (N_47890,N_47002,N_47429);
xnor U47891 (N_47891,N_47395,N_47377);
or U47892 (N_47892,N_47230,N_47366);
or U47893 (N_47893,N_47420,N_47314);
and U47894 (N_47894,N_47109,N_47186);
nand U47895 (N_47895,N_47340,N_47243);
xor U47896 (N_47896,N_47335,N_47360);
nand U47897 (N_47897,N_47348,N_47225);
or U47898 (N_47898,N_47065,N_47277);
and U47899 (N_47899,N_47482,N_47343);
nand U47900 (N_47900,N_47463,N_47498);
or U47901 (N_47901,N_47063,N_47073);
and U47902 (N_47902,N_47249,N_47485);
or U47903 (N_47903,N_47024,N_47391);
xnor U47904 (N_47904,N_47151,N_47138);
nor U47905 (N_47905,N_47150,N_47447);
and U47906 (N_47906,N_47195,N_47112);
or U47907 (N_47907,N_47123,N_47396);
nor U47908 (N_47908,N_47465,N_47090);
or U47909 (N_47909,N_47403,N_47272);
nand U47910 (N_47910,N_47389,N_47468);
nand U47911 (N_47911,N_47358,N_47003);
and U47912 (N_47912,N_47037,N_47244);
or U47913 (N_47913,N_47290,N_47135);
nand U47914 (N_47914,N_47093,N_47477);
nand U47915 (N_47915,N_47447,N_47133);
or U47916 (N_47916,N_47397,N_47163);
and U47917 (N_47917,N_47042,N_47258);
and U47918 (N_47918,N_47175,N_47255);
or U47919 (N_47919,N_47347,N_47380);
nor U47920 (N_47920,N_47150,N_47489);
xor U47921 (N_47921,N_47310,N_47452);
or U47922 (N_47922,N_47250,N_47439);
or U47923 (N_47923,N_47139,N_47103);
and U47924 (N_47924,N_47401,N_47457);
or U47925 (N_47925,N_47170,N_47302);
and U47926 (N_47926,N_47076,N_47424);
nand U47927 (N_47927,N_47408,N_47001);
and U47928 (N_47928,N_47168,N_47070);
xnor U47929 (N_47929,N_47482,N_47332);
nand U47930 (N_47930,N_47048,N_47488);
xnor U47931 (N_47931,N_47160,N_47424);
nor U47932 (N_47932,N_47342,N_47066);
and U47933 (N_47933,N_47359,N_47026);
xnor U47934 (N_47934,N_47243,N_47058);
and U47935 (N_47935,N_47223,N_47184);
or U47936 (N_47936,N_47060,N_47082);
xor U47937 (N_47937,N_47323,N_47386);
and U47938 (N_47938,N_47127,N_47218);
xor U47939 (N_47939,N_47142,N_47190);
or U47940 (N_47940,N_47153,N_47069);
xnor U47941 (N_47941,N_47416,N_47137);
nand U47942 (N_47942,N_47404,N_47096);
nand U47943 (N_47943,N_47284,N_47450);
nand U47944 (N_47944,N_47318,N_47345);
xnor U47945 (N_47945,N_47474,N_47401);
nor U47946 (N_47946,N_47393,N_47375);
nand U47947 (N_47947,N_47234,N_47010);
and U47948 (N_47948,N_47176,N_47335);
or U47949 (N_47949,N_47321,N_47479);
or U47950 (N_47950,N_47216,N_47457);
or U47951 (N_47951,N_47423,N_47386);
xor U47952 (N_47952,N_47207,N_47078);
xnor U47953 (N_47953,N_47329,N_47360);
nand U47954 (N_47954,N_47298,N_47011);
xnor U47955 (N_47955,N_47082,N_47363);
or U47956 (N_47956,N_47279,N_47198);
and U47957 (N_47957,N_47009,N_47089);
xnor U47958 (N_47958,N_47036,N_47393);
nand U47959 (N_47959,N_47195,N_47438);
xnor U47960 (N_47960,N_47308,N_47328);
and U47961 (N_47961,N_47343,N_47296);
nor U47962 (N_47962,N_47096,N_47091);
nor U47963 (N_47963,N_47090,N_47383);
nand U47964 (N_47964,N_47341,N_47394);
nand U47965 (N_47965,N_47005,N_47064);
and U47966 (N_47966,N_47064,N_47192);
nand U47967 (N_47967,N_47352,N_47179);
nor U47968 (N_47968,N_47348,N_47281);
xnor U47969 (N_47969,N_47099,N_47325);
nor U47970 (N_47970,N_47345,N_47428);
or U47971 (N_47971,N_47140,N_47146);
nand U47972 (N_47972,N_47027,N_47188);
and U47973 (N_47973,N_47266,N_47456);
or U47974 (N_47974,N_47274,N_47068);
nor U47975 (N_47975,N_47080,N_47484);
and U47976 (N_47976,N_47462,N_47171);
nand U47977 (N_47977,N_47120,N_47370);
or U47978 (N_47978,N_47272,N_47261);
nand U47979 (N_47979,N_47281,N_47094);
and U47980 (N_47980,N_47036,N_47413);
nor U47981 (N_47981,N_47130,N_47216);
xnor U47982 (N_47982,N_47244,N_47179);
xor U47983 (N_47983,N_47413,N_47074);
xor U47984 (N_47984,N_47047,N_47214);
xor U47985 (N_47985,N_47135,N_47020);
and U47986 (N_47986,N_47123,N_47294);
and U47987 (N_47987,N_47385,N_47058);
nand U47988 (N_47988,N_47062,N_47432);
or U47989 (N_47989,N_47440,N_47438);
xnor U47990 (N_47990,N_47429,N_47174);
nor U47991 (N_47991,N_47088,N_47323);
or U47992 (N_47992,N_47233,N_47472);
and U47993 (N_47993,N_47362,N_47221);
nor U47994 (N_47994,N_47144,N_47449);
nor U47995 (N_47995,N_47400,N_47129);
or U47996 (N_47996,N_47445,N_47430);
nor U47997 (N_47997,N_47174,N_47074);
and U47998 (N_47998,N_47397,N_47133);
and U47999 (N_47999,N_47450,N_47417);
or U48000 (N_48000,N_47638,N_47918);
or U48001 (N_48001,N_47680,N_47672);
and U48002 (N_48002,N_47590,N_47930);
nand U48003 (N_48003,N_47934,N_47632);
nand U48004 (N_48004,N_47987,N_47780);
or U48005 (N_48005,N_47521,N_47889);
nand U48006 (N_48006,N_47654,N_47950);
xor U48007 (N_48007,N_47929,N_47796);
and U48008 (N_48008,N_47718,N_47967);
nor U48009 (N_48009,N_47728,N_47757);
nand U48010 (N_48010,N_47702,N_47914);
and U48011 (N_48011,N_47798,N_47819);
nor U48012 (N_48012,N_47651,N_47969);
xor U48013 (N_48013,N_47817,N_47971);
nor U48014 (N_48014,N_47942,N_47512);
xnor U48015 (N_48015,N_47980,N_47885);
and U48016 (N_48016,N_47856,N_47542);
nor U48017 (N_48017,N_47938,N_47847);
xnor U48018 (N_48018,N_47562,N_47848);
and U48019 (N_48019,N_47818,N_47553);
nor U48020 (N_48020,N_47804,N_47623);
nand U48021 (N_48021,N_47835,N_47519);
nand U48022 (N_48022,N_47840,N_47713);
nand U48023 (N_48023,N_47573,N_47705);
nor U48024 (N_48024,N_47721,N_47744);
xnor U48025 (N_48025,N_47671,N_47745);
nor U48026 (N_48026,N_47740,N_47838);
and U48027 (N_48027,N_47583,N_47944);
nand U48028 (N_48028,N_47800,N_47621);
nand U48029 (N_48029,N_47598,N_47961);
nor U48030 (N_48030,N_47755,N_47582);
xor U48031 (N_48031,N_47986,N_47701);
xor U48032 (N_48032,N_47907,N_47567);
nand U48033 (N_48033,N_47895,N_47826);
xnor U48034 (N_48034,N_47979,N_47712);
or U48035 (N_48035,N_47606,N_47915);
or U48036 (N_48036,N_47549,N_47832);
or U48037 (N_48037,N_47683,N_47710);
xor U48038 (N_48038,N_47875,N_47649);
nor U48039 (N_48039,N_47630,N_47593);
nand U48040 (N_48040,N_47834,N_47715);
xor U48041 (N_48041,N_47697,N_47788);
nor U48042 (N_48042,N_47836,N_47855);
nor U48043 (N_48043,N_47673,N_47896);
or U48044 (N_48044,N_47978,N_47596);
or U48045 (N_48045,N_47816,N_47505);
and U48046 (N_48046,N_47510,N_47877);
or U48047 (N_48047,N_47501,N_47793);
and U48048 (N_48048,N_47734,N_47642);
or U48049 (N_48049,N_47554,N_47663);
and U48050 (N_48050,N_47524,N_47741);
or U48051 (N_48051,N_47903,N_47974);
or U48052 (N_48052,N_47933,N_47503);
or U48053 (N_48053,N_47991,N_47584);
nand U48054 (N_48054,N_47650,N_47733);
xnor U48055 (N_48055,N_47940,N_47911);
or U48056 (N_48056,N_47926,N_47865);
nand U48057 (N_48057,N_47628,N_47694);
or U48058 (N_48058,N_47758,N_47749);
xor U48059 (N_48059,N_47677,N_47775);
or U48060 (N_48060,N_47791,N_47823);
and U48061 (N_48061,N_47666,N_47668);
nor U48062 (N_48062,N_47787,N_47679);
nor U48063 (N_48063,N_47686,N_47891);
or U48064 (N_48064,N_47575,N_47846);
nand U48065 (N_48065,N_47676,N_47892);
nor U48066 (N_48066,N_47808,N_47990);
and U48067 (N_48067,N_47965,N_47552);
nand U48068 (N_48068,N_47629,N_47858);
and U48069 (N_48069,N_47812,N_47597);
nor U48070 (N_48070,N_47664,N_47594);
and U48071 (N_48071,N_47727,N_47704);
nor U48072 (N_48072,N_47906,N_47556);
and U48073 (N_48073,N_47587,N_47941);
or U48074 (N_48074,N_47620,N_47852);
and U48075 (N_48075,N_47912,N_47658);
nor U48076 (N_48076,N_47964,N_47994);
xnor U48077 (N_48077,N_47960,N_47997);
and U48078 (N_48078,N_47528,N_47548);
nor U48079 (N_48079,N_47609,N_47878);
or U48080 (N_48080,N_47534,N_47772);
nor U48081 (N_48081,N_47563,N_47529);
xnor U48082 (N_48082,N_47936,N_47627);
xor U48083 (N_48083,N_47983,N_47670);
xnor U48084 (N_48084,N_47917,N_47899);
nand U48085 (N_48085,N_47866,N_47689);
or U48086 (N_48086,N_47633,N_47561);
or U48087 (N_48087,N_47514,N_47830);
nor U48088 (N_48088,N_47531,N_47693);
nor U48089 (N_48089,N_47982,N_47883);
and U48090 (N_48090,N_47853,N_47770);
nor U48091 (N_48091,N_47833,N_47854);
xnor U48092 (N_48092,N_47970,N_47643);
nor U48093 (N_48093,N_47760,N_47935);
nor U48094 (N_48094,N_47726,N_47972);
or U48095 (N_48095,N_47515,N_47943);
and U48096 (N_48096,N_47873,N_47523);
nor U48097 (N_48097,N_47558,N_47829);
and U48098 (N_48098,N_47973,N_47618);
nand U48099 (N_48099,N_47736,N_47952);
or U48100 (N_48100,N_47636,N_47611);
nand U48101 (N_48101,N_47814,N_47536);
nor U48102 (N_48102,N_47998,N_47882);
nor U48103 (N_48103,N_47706,N_47996);
nand U48104 (N_48104,N_47585,N_47541);
nor U48105 (N_48105,N_47748,N_47500);
nand U48106 (N_48106,N_47828,N_47779);
or U48107 (N_48107,N_47566,N_47859);
nor U48108 (N_48108,N_47752,N_47842);
nor U48109 (N_48109,N_47517,N_47526);
and U48110 (N_48110,N_47862,N_47844);
and U48111 (N_48111,N_47886,N_47731);
xor U48112 (N_48112,N_47735,N_47684);
nand U48113 (N_48113,N_47580,N_47999);
xnor U48114 (N_48114,N_47586,N_47525);
and U48115 (N_48115,N_47747,N_47550);
or U48116 (N_48116,N_47698,N_47708);
and U48117 (N_48117,N_47504,N_47872);
nor U48118 (N_48118,N_47923,N_47781);
and U48119 (N_48119,N_47902,N_47669);
nand U48120 (N_48120,N_47551,N_47884);
nand U48121 (N_48121,N_47954,N_47900);
xnor U48122 (N_48122,N_47719,N_47574);
nand U48123 (N_48123,N_47690,N_47894);
nand U48124 (N_48124,N_47678,N_47615);
nand U48125 (N_48125,N_47756,N_47932);
nand U48126 (N_48126,N_47540,N_47822);
and U48127 (N_48127,N_47841,N_47916);
xnor U48128 (N_48128,N_47951,N_47695);
nor U48129 (N_48129,N_47762,N_47730);
or U48130 (N_48130,N_47774,N_47839);
and U48131 (N_48131,N_47616,N_47685);
nor U48132 (N_48132,N_47813,N_47724);
nand U48133 (N_48133,N_47778,N_47769);
or U48134 (N_48134,N_47624,N_47837);
and U48135 (N_48135,N_47981,N_47592);
or U48136 (N_48136,N_47559,N_47539);
nand U48137 (N_48137,N_47555,N_47924);
or U48138 (N_48138,N_47975,N_47645);
xnor U48139 (N_48139,N_47958,N_47544);
nand U48140 (N_48140,N_47904,N_47963);
and U48141 (N_48141,N_47675,N_47945);
nand U48142 (N_48142,N_47513,N_47532);
nand U48143 (N_48143,N_47568,N_47985);
nand U48144 (N_48144,N_47545,N_47992);
nand U48145 (N_48145,N_47720,N_47723);
nor U48146 (N_48146,N_47700,N_47546);
or U48147 (N_48147,N_47761,N_47861);
and U48148 (N_48148,N_47605,N_47977);
nand U48149 (N_48149,N_47639,N_47782);
xor U48150 (N_48150,N_47516,N_47893);
and U48151 (N_48151,N_47810,N_47931);
nor U48152 (N_48152,N_47845,N_47647);
or U48153 (N_48153,N_47876,N_47599);
and U48154 (N_48154,N_47763,N_47984);
nor U48155 (N_48155,N_47610,N_47644);
or U48156 (N_48156,N_47809,N_47802);
and U48157 (N_48157,N_47785,N_47790);
nand U48158 (N_48158,N_47857,N_47820);
xor U48159 (N_48159,N_47682,N_47959);
nor U48160 (N_48160,N_47827,N_47789);
and U48161 (N_48161,N_47527,N_47688);
and U48162 (N_48162,N_47619,N_47622);
or U48163 (N_48163,N_47655,N_47759);
or U48164 (N_48164,N_47995,N_47625);
nand U48165 (N_48165,N_47920,N_47949);
xor U48166 (N_48166,N_47711,N_47732);
or U48167 (N_48167,N_47767,N_47581);
nand U48168 (N_48168,N_47898,N_47976);
or U48169 (N_48169,N_47947,N_47612);
or U48170 (N_48170,N_47577,N_47910);
nor U48171 (N_48171,N_47714,N_47707);
nor U48172 (N_48172,N_47824,N_47795);
and U48173 (N_48173,N_47777,N_47921);
nand U48174 (N_48174,N_47870,N_47955);
and U48175 (N_48175,N_47722,N_47530);
nor U48176 (N_48176,N_47806,N_47538);
xor U48177 (N_48177,N_47589,N_47508);
nor U48178 (N_48178,N_47662,N_47871);
and U48179 (N_48179,N_47968,N_47617);
xor U48180 (N_48180,N_47913,N_47956);
nand U48181 (N_48181,N_47815,N_47771);
and U48182 (N_48182,N_47863,N_47699);
nand U48183 (N_48183,N_47867,N_47881);
xnor U48184 (N_48184,N_47608,N_47709);
nand U48185 (N_48185,N_47989,N_47656);
or U48186 (N_48186,N_47604,N_47887);
and U48187 (N_48187,N_47773,N_47507);
xor U48188 (N_48188,N_47603,N_47860);
nand U48189 (N_48189,N_47879,N_47716);
nor U48190 (N_48190,N_47803,N_47890);
or U48191 (N_48191,N_47657,N_47753);
nand U48192 (N_48192,N_47533,N_47880);
and U48193 (N_48193,N_47601,N_47653);
xor U48194 (N_48194,N_47850,N_47908);
xnor U48195 (N_48195,N_47901,N_47725);
and U48196 (N_48196,N_47953,N_47737);
and U48197 (N_48197,N_47600,N_47799);
nor U48198 (N_48198,N_47743,N_47742);
nand U48199 (N_48199,N_47674,N_47626);
and U48200 (N_48200,N_47948,N_47572);
nor U48201 (N_48201,N_47768,N_47631);
xnor U48202 (N_48202,N_47843,N_47776);
and U48203 (N_48203,N_47831,N_47506);
nand U48204 (N_48204,N_47784,N_47560);
xnor U48205 (N_48205,N_47535,N_47905);
or U48206 (N_48206,N_47579,N_47874);
nand U48207 (N_48207,N_47634,N_47739);
xnor U48208 (N_48208,N_47557,N_47646);
xnor U48209 (N_48209,N_47825,N_47993);
and U48210 (N_48210,N_47957,N_47888);
nand U48211 (N_48211,N_47511,N_47864);
nor U48212 (N_48212,N_47637,N_47652);
or U48213 (N_48213,N_47751,N_47635);
nand U48214 (N_48214,N_47518,N_47919);
nand U48215 (N_48215,N_47570,N_47851);
nand U48216 (N_48216,N_47691,N_47746);
and U48217 (N_48217,N_47807,N_47805);
nor U48218 (N_48218,N_47661,N_47687);
nand U48219 (N_48219,N_47607,N_47922);
and U48220 (N_48220,N_47576,N_47738);
or U48221 (N_48221,N_47794,N_47641);
or U48222 (N_48222,N_47569,N_47648);
xnor U48223 (N_48223,N_47537,N_47717);
or U48224 (N_48224,N_47925,N_47946);
or U48225 (N_48225,N_47939,N_47588);
nand U48226 (N_48226,N_47750,N_47571);
and U48227 (N_48227,N_47729,N_47821);
nor U48228 (N_48228,N_47522,N_47909);
or U48229 (N_48229,N_47966,N_47591);
nand U48230 (N_48230,N_47543,N_47783);
nand U48231 (N_48231,N_47988,N_47502);
nand U48232 (N_48232,N_47764,N_47640);
xor U48233 (N_48233,N_47696,N_47937);
or U48234 (N_48234,N_47801,N_47927);
and U48235 (N_48235,N_47565,N_47520);
nand U48236 (N_48236,N_47602,N_47692);
nand U48237 (N_48237,N_47849,N_47754);
xor U48238 (N_48238,N_47928,N_47869);
or U48239 (N_48239,N_47962,N_47564);
xor U48240 (N_48240,N_47667,N_47614);
xor U48241 (N_48241,N_47578,N_47509);
or U48242 (N_48242,N_47868,N_47897);
and U48243 (N_48243,N_47703,N_47797);
xnor U48244 (N_48244,N_47665,N_47792);
and U48245 (N_48245,N_47659,N_47786);
nand U48246 (N_48246,N_47595,N_47660);
and U48247 (N_48247,N_47811,N_47613);
and U48248 (N_48248,N_47681,N_47547);
or U48249 (N_48249,N_47765,N_47766);
nand U48250 (N_48250,N_47553,N_47812);
xor U48251 (N_48251,N_47830,N_47698);
xnor U48252 (N_48252,N_47840,N_47703);
nand U48253 (N_48253,N_47969,N_47641);
xor U48254 (N_48254,N_47937,N_47506);
or U48255 (N_48255,N_47578,N_47870);
xor U48256 (N_48256,N_47780,N_47563);
nand U48257 (N_48257,N_47738,N_47638);
or U48258 (N_48258,N_47668,N_47905);
nand U48259 (N_48259,N_47520,N_47883);
xnor U48260 (N_48260,N_47761,N_47641);
nor U48261 (N_48261,N_47608,N_47749);
nand U48262 (N_48262,N_47986,N_47659);
nand U48263 (N_48263,N_47748,N_47995);
and U48264 (N_48264,N_47990,N_47660);
nand U48265 (N_48265,N_47978,N_47883);
xor U48266 (N_48266,N_47777,N_47604);
and U48267 (N_48267,N_47599,N_47996);
or U48268 (N_48268,N_47522,N_47792);
xnor U48269 (N_48269,N_47508,N_47814);
nand U48270 (N_48270,N_47508,N_47564);
or U48271 (N_48271,N_47786,N_47751);
nand U48272 (N_48272,N_47661,N_47766);
or U48273 (N_48273,N_47787,N_47756);
or U48274 (N_48274,N_47981,N_47705);
nor U48275 (N_48275,N_47664,N_47767);
nor U48276 (N_48276,N_47515,N_47911);
xnor U48277 (N_48277,N_47530,N_47623);
xor U48278 (N_48278,N_47840,N_47885);
and U48279 (N_48279,N_47738,N_47664);
xnor U48280 (N_48280,N_47779,N_47851);
xor U48281 (N_48281,N_47583,N_47916);
and U48282 (N_48282,N_47760,N_47693);
xor U48283 (N_48283,N_47705,N_47640);
nand U48284 (N_48284,N_47907,N_47666);
or U48285 (N_48285,N_47965,N_47503);
xnor U48286 (N_48286,N_47631,N_47777);
or U48287 (N_48287,N_47587,N_47911);
nor U48288 (N_48288,N_47955,N_47621);
nand U48289 (N_48289,N_47797,N_47694);
and U48290 (N_48290,N_47528,N_47836);
nand U48291 (N_48291,N_47932,N_47565);
or U48292 (N_48292,N_47643,N_47567);
or U48293 (N_48293,N_47732,N_47626);
nand U48294 (N_48294,N_47714,N_47917);
xnor U48295 (N_48295,N_47558,N_47825);
or U48296 (N_48296,N_47992,N_47993);
xor U48297 (N_48297,N_47981,N_47726);
nor U48298 (N_48298,N_47895,N_47574);
nor U48299 (N_48299,N_47933,N_47623);
or U48300 (N_48300,N_47887,N_47957);
nand U48301 (N_48301,N_47689,N_47604);
nand U48302 (N_48302,N_47682,N_47507);
xnor U48303 (N_48303,N_47620,N_47644);
and U48304 (N_48304,N_47960,N_47852);
or U48305 (N_48305,N_47879,N_47506);
xnor U48306 (N_48306,N_47730,N_47555);
xnor U48307 (N_48307,N_47574,N_47834);
xnor U48308 (N_48308,N_47599,N_47825);
and U48309 (N_48309,N_47852,N_47973);
nor U48310 (N_48310,N_47747,N_47563);
xnor U48311 (N_48311,N_47813,N_47965);
nand U48312 (N_48312,N_47647,N_47949);
nand U48313 (N_48313,N_47729,N_47819);
and U48314 (N_48314,N_47564,N_47989);
nand U48315 (N_48315,N_47770,N_47623);
nand U48316 (N_48316,N_47916,N_47668);
xor U48317 (N_48317,N_47753,N_47673);
and U48318 (N_48318,N_47843,N_47929);
nand U48319 (N_48319,N_47989,N_47683);
and U48320 (N_48320,N_47640,N_47841);
xor U48321 (N_48321,N_47973,N_47672);
and U48322 (N_48322,N_47985,N_47981);
and U48323 (N_48323,N_47907,N_47942);
xor U48324 (N_48324,N_47865,N_47691);
xor U48325 (N_48325,N_47779,N_47776);
or U48326 (N_48326,N_47904,N_47626);
or U48327 (N_48327,N_47673,N_47594);
nor U48328 (N_48328,N_47948,N_47711);
xor U48329 (N_48329,N_47533,N_47518);
nand U48330 (N_48330,N_47881,N_47882);
nor U48331 (N_48331,N_47998,N_47932);
xnor U48332 (N_48332,N_47541,N_47863);
xnor U48333 (N_48333,N_47733,N_47758);
nor U48334 (N_48334,N_47862,N_47950);
and U48335 (N_48335,N_47814,N_47739);
xor U48336 (N_48336,N_47968,N_47813);
nor U48337 (N_48337,N_47986,N_47508);
nor U48338 (N_48338,N_47543,N_47566);
xnor U48339 (N_48339,N_47986,N_47989);
nor U48340 (N_48340,N_47985,N_47718);
nand U48341 (N_48341,N_47597,N_47837);
xor U48342 (N_48342,N_47620,N_47904);
or U48343 (N_48343,N_47788,N_47540);
xor U48344 (N_48344,N_47572,N_47850);
nand U48345 (N_48345,N_47912,N_47730);
xnor U48346 (N_48346,N_47554,N_47913);
nor U48347 (N_48347,N_47736,N_47670);
xor U48348 (N_48348,N_47966,N_47930);
or U48349 (N_48349,N_47571,N_47867);
xor U48350 (N_48350,N_47895,N_47686);
or U48351 (N_48351,N_47635,N_47556);
nand U48352 (N_48352,N_47684,N_47951);
and U48353 (N_48353,N_47894,N_47934);
or U48354 (N_48354,N_47708,N_47712);
nor U48355 (N_48355,N_47979,N_47905);
and U48356 (N_48356,N_47873,N_47511);
and U48357 (N_48357,N_47605,N_47966);
nand U48358 (N_48358,N_47892,N_47961);
or U48359 (N_48359,N_47733,N_47658);
xor U48360 (N_48360,N_47518,N_47766);
and U48361 (N_48361,N_47682,N_47861);
nor U48362 (N_48362,N_47869,N_47942);
and U48363 (N_48363,N_47564,N_47548);
nand U48364 (N_48364,N_47727,N_47634);
nand U48365 (N_48365,N_47683,N_47644);
xor U48366 (N_48366,N_47534,N_47768);
nand U48367 (N_48367,N_47771,N_47966);
nand U48368 (N_48368,N_47627,N_47561);
xor U48369 (N_48369,N_47839,N_47587);
nand U48370 (N_48370,N_47784,N_47514);
or U48371 (N_48371,N_47912,N_47611);
nand U48372 (N_48372,N_47857,N_47950);
nor U48373 (N_48373,N_47915,N_47893);
and U48374 (N_48374,N_47667,N_47923);
nand U48375 (N_48375,N_47770,N_47634);
nand U48376 (N_48376,N_47970,N_47921);
or U48377 (N_48377,N_47815,N_47606);
nand U48378 (N_48378,N_47530,N_47590);
xnor U48379 (N_48379,N_47996,N_47715);
nand U48380 (N_48380,N_47867,N_47652);
nand U48381 (N_48381,N_47966,N_47737);
nor U48382 (N_48382,N_47868,N_47683);
and U48383 (N_48383,N_47657,N_47929);
nor U48384 (N_48384,N_47521,N_47756);
and U48385 (N_48385,N_47504,N_47664);
or U48386 (N_48386,N_47735,N_47504);
or U48387 (N_48387,N_47907,N_47891);
xnor U48388 (N_48388,N_47726,N_47514);
or U48389 (N_48389,N_47684,N_47800);
or U48390 (N_48390,N_47506,N_47756);
nor U48391 (N_48391,N_47933,N_47768);
or U48392 (N_48392,N_47891,N_47923);
and U48393 (N_48393,N_47549,N_47866);
nand U48394 (N_48394,N_47618,N_47817);
nor U48395 (N_48395,N_47754,N_47847);
or U48396 (N_48396,N_47983,N_47974);
nor U48397 (N_48397,N_47623,N_47561);
nand U48398 (N_48398,N_47914,N_47732);
nand U48399 (N_48399,N_47551,N_47698);
nand U48400 (N_48400,N_47982,N_47788);
xor U48401 (N_48401,N_47892,N_47574);
and U48402 (N_48402,N_47641,N_47702);
nand U48403 (N_48403,N_47944,N_47652);
and U48404 (N_48404,N_47729,N_47518);
or U48405 (N_48405,N_47977,N_47886);
nor U48406 (N_48406,N_47856,N_47809);
and U48407 (N_48407,N_47862,N_47650);
and U48408 (N_48408,N_47529,N_47786);
or U48409 (N_48409,N_47566,N_47559);
and U48410 (N_48410,N_47805,N_47798);
and U48411 (N_48411,N_47865,N_47846);
or U48412 (N_48412,N_47716,N_47749);
nor U48413 (N_48413,N_47555,N_47884);
or U48414 (N_48414,N_47775,N_47709);
nand U48415 (N_48415,N_47817,N_47838);
or U48416 (N_48416,N_47829,N_47807);
xor U48417 (N_48417,N_47915,N_47632);
or U48418 (N_48418,N_47519,N_47864);
xnor U48419 (N_48419,N_47739,N_47784);
nor U48420 (N_48420,N_47896,N_47532);
nor U48421 (N_48421,N_47849,N_47534);
or U48422 (N_48422,N_47675,N_47698);
nand U48423 (N_48423,N_47512,N_47852);
nand U48424 (N_48424,N_47702,N_47816);
or U48425 (N_48425,N_47764,N_47955);
nor U48426 (N_48426,N_47800,N_47711);
and U48427 (N_48427,N_47625,N_47694);
nor U48428 (N_48428,N_47848,N_47840);
nor U48429 (N_48429,N_47511,N_47978);
nand U48430 (N_48430,N_47516,N_47892);
and U48431 (N_48431,N_47808,N_47667);
or U48432 (N_48432,N_47847,N_47779);
xor U48433 (N_48433,N_47822,N_47939);
and U48434 (N_48434,N_47844,N_47673);
nand U48435 (N_48435,N_47874,N_47572);
and U48436 (N_48436,N_47674,N_47639);
or U48437 (N_48437,N_47774,N_47816);
nor U48438 (N_48438,N_47754,N_47604);
nand U48439 (N_48439,N_47954,N_47879);
xnor U48440 (N_48440,N_47698,N_47722);
or U48441 (N_48441,N_47881,N_47818);
nor U48442 (N_48442,N_47835,N_47898);
or U48443 (N_48443,N_47859,N_47694);
nor U48444 (N_48444,N_47992,N_47724);
and U48445 (N_48445,N_47694,N_47720);
nor U48446 (N_48446,N_47687,N_47849);
or U48447 (N_48447,N_47615,N_47562);
or U48448 (N_48448,N_47813,N_47811);
or U48449 (N_48449,N_47966,N_47530);
or U48450 (N_48450,N_47597,N_47802);
xnor U48451 (N_48451,N_47666,N_47508);
or U48452 (N_48452,N_47622,N_47916);
and U48453 (N_48453,N_47519,N_47643);
and U48454 (N_48454,N_47902,N_47883);
or U48455 (N_48455,N_47635,N_47620);
nor U48456 (N_48456,N_47648,N_47659);
nand U48457 (N_48457,N_47688,N_47640);
xnor U48458 (N_48458,N_47826,N_47796);
and U48459 (N_48459,N_47556,N_47768);
xor U48460 (N_48460,N_47971,N_47989);
and U48461 (N_48461,N_47883,N_47718);
or U48462 (N_48462,N_47920,N_47527);
xor U48463 (N_48463,N_47914,N_47910);
and U48464 (N_48464,N_47838,N_47815);
and U48465 (N_48465,N_47585,N_47536);
or U48466 (N_48466,N_47900,N_47987);
nand U48467 (N_48467,N_47994,N_47650);
nand U48468 (N_48468,N_47568,N_47892);
and U48469 (N_48469,N_47855,N_47653);
and U48470 (N_48470,N_47687,N_47510);
nor U48471 (N_48471,N_47675,N_47962);
nand U48472 (N_48472,N_47733,N_47664);
or U48473 (N_48473,N_47802,N_47721);
xnor U48474 (N_48474,N_47509,N_47783);
or U48475 (N_48475,N_47796,N_47682);
or U48476 (N_48476,N_47949,N_47767);
and U48477 (N_48477,N_47873,N_47704);
and U48478 (N_48478,N_47694,N_47806);
or U48479 (N_48479,N_47844,N_47550);
xor U48480 (N_48480,N_47698,N_47702);
nor U48481 (N_48481,N_47755,N_47971);
and U48482 (N_48482,N_47516,N_47708);
xor U48483 (N_48483,N_47931,N_47809);
nor U48484 (N_48484,N_47845,N_47713);
or U48485 (N_48485,N_47902,N_47897);
xor U48486 (N_48486,N_47908,N_47500);
xor U48487 (N_48487,N_47500,N_47618);
or U48488 (N_48488,N_47996,N_47975);
and U48489 (N_48489,N_47791,N_47564);
nor U48490 (N_48490,N_47870,N_47866);
and U48491 (N_48491,N_47754,N_47836);
and U48492 (N_48492,N_47539,N_47504);
xor U48493 (N_48493,N_47707,N_47777);
xnor U48494 (N_48494,N_47727,N_47895);
or U48495 (N_48495,N_47793,N_47696);
or U48496 (N_48496,N_47825,N_47932);
and U48497 (N_48497,N_47566,N_47658);
nor U48498 (N_48498,N_47750,N_47775);
and U48499 (N_48499,N_47986,N_47587);
xor U48500 (N_48500,N_48293,N_48351);
nor U48501 (N_48501,N_48040,N_48330);
nand U48502 (N_48502,N_48276,N_48005);
nor U48503 (N_48503,N_48016,N_48286);
or U48504 (N_48504,N_48116,N_48490);
nand U48505 (N_48505,N_48080,N_48349);
and U48506 (N_48506,N_48170,N_48001);
nand U48507 (N_48507,N_48290,N_48429);
or U48508 (N_48508,N_48288,N_48191);
or U48509 (N_48509,N_48274,N_48063);
or U48510 (N_48510,N_48099,N_48424);
nand U48511 (N_48511,N_48243,N_48294);
and U48512 (N_48512,N_48095,N_48051);
nand U48513 (N_48513,N_48245,N_48162);
and U48514 (N_48514,N_48093,N_48186);
nor U48515 (N_48515,N_48184,N_48432);
or U48516 (N_48516,N_48129,N_48239);
xor U48517 (N_48517,N_48345,N_48299);
nor U48518 (N_48518,N_48096,N_48034);
nor U48519 (N_48519,N_48339,N_48205);
xor U48520 (N_48520,N_48120,N_48378);
nand U48521 (N_48521,N_48206,N_48145);
nor U48522 (N_48522,N_48173,N_48121);
and U48523 (N_48523,N_48049,N_48444);
or U48524 (N_48524,N_48178,N_48317);
nor U48525 (N_48525,N_48418,N_48315);
or U48526 (N_48526,N_48371,N_48018);
or U48527 (N_48527,N_48227,N_48430);
nor U48528 (N_48528,N_48013,N_48219);
nand U48529 (N_48529,N_48411,N_48254);
and U48530 (N_48530,N_48118,N_48039);
xor U48531 (N_48531,N_48390,N_48014);
xnor U48532 (N_48532,N_48217,N_48468);
nor U48533 (N_48533,N_48123,N_48332);
nand U48534 (N_48534,N_48259,N_48450);
and U48535 (N_48535,N_48214,N_48305);
xnor U48536 (N_48536,N_48155,N_48037);
and U48537 (N_48537,N_48238,N_48374);
and U48538 (N_48538,N_48078,N_48140);
or U48539 (N_48539,N_48019,N_48327);
xor U48540 (N_48540,N_48314,N_48434);
xnor U48541 (N_48541,N_48175,N_48365);
nand U48542 (N_48542,N_48142,N_48149);
nor U48543 (N_48543,N_48225,N_48190);
xnor U48544 (N_48544,N_48253,N_48114);
xor U48545 (N_48545,N_48158,N_48043);
or U48546 (N_48546,N_48394,N_48348);
or U48547 (N_48547,N_48475,N_48012);
xnor U48548 (N_48548,N_48202,N_48221);
nor U48549 (N_48549,N_48073,N_48367);
xor U48550 (N_48550,N_48174,N_48067);
nand U48551 (N_48551,N_48493,N_48313);
and U48552 (N_48552,N_48210,N_48406);
nand U48553 (N_48553,N_48117,N_48104);
xnor U48554 (N_48554,N_48248,N_48060);
nand U48555 (N_48555,N_48062,N_48364);
xor U48556 (N_48556,N_48420,N_48204);
nor U48557 (N_48557,N_48124,N_48192);
or U48558 (N_48558,N_48464,N_48194);
xnor U48559 (N_48559,N_48074,N_48359);
nor U48560 (N_48560,N_48168,N_48494);
and U48561 (N_48561,N_48201,N_48488);
nand U48562 (N_48562,N_48296,N_48237);
and U48563 (N_48563,N_48391,N_48179);
nand U48564 (N_48564,N_48182,N_48209);
xor U48565 (N_48565,N_48047,N_48350);
and U48566 (N_48566,N_48025,N_48403);
xor U48567 (N_48567,N_48446,N_48386);
nand U48568 (N_48568,N_48109,N_48233);
xor U48569 (N_48569,N_48368,N_48112);
xnor U48570 (N_48570,N_48193,N_48366);
nor U48571 (N_48571,N_48222,N_48106);
or U48572 (N_48572,N_48007,N_48415);
nand U48573 (N_48573,N_48304,N_48275);
nand U48574 (N_48574,N_48277,N_48100);
and U48575 (N_48575,N_48393,N_48387);
and U48576 (N_48576,N_48224,N_48460);
xor U48577 (N_48577,N_48108,N_48144);
nor U48578 (N_48578,N_48402,N_48401);
nand U48579 (N_48579,N_48260,N_48269);
and U48580 (N_48580,N_48115,N_48427);
or U48581 (N_48581,N_48303,N_48309);
or U48582 (N_48582,N_48491,N_48256);
nor U48583 (N_48583,N_48297,N_48384);
nand U48584 (N_48584,N_48483,N_48130);
nand U48585 (N_48585,N_48101,N_48030);
xnor U48586 (N_48586,N_48215,N_48485);
nor U48587 (N_48587,N_48328,N_48375);
or U48588 (N_48588,N_48150,N_48456);
xor U48589 (N_48589,N_48031,N_48183);
xnor U48590 (N_48590,N_48344,N_48022);
nand U48591 (N_48591,N_48058,N_48477);
nand U48592 (N_48592,N_48203,N_48362);
nand U48593 (N_48593,N_48311,N_48467);
nor U48594 (N_48594,N_48153,N_48133);
and U48595 (N_48595,N_48492,N_48033);
and U48596 (N_48596,N_48268,N_48340);
nand U48597 (N_48597,N_48481,N_48449);
and U48598 (N_48598,N_48141,N_48353);
nor U48599 (N_48599,N_48105,N_48176);
or U48600 (N_48600,N_48015,N_48357);
nand U48601 (N_48601,N_48342,N_48271);
xor U48602 (N_48602,N_48041,N_48180);
nand U48603 (N_48603,N_48377,N_48052);
or U48604 (N_48604,N_48316,N_48321);
nand U48605 (N_48605,N_48090,N_48474);
and U48606 (N_48606,N_48138,N_48451);
or U48607 (N_48607,N_48066,N_48181);
nor U48608 (N_48608,N_48002,N_48208);
or U48609 (N_48609,N_48281,N_48472);
xnor U48610 (N_48610,N_48068,N_48382);
and U48611 (N_48611,N_48128,N_48482);
or U48612 (N_48612,N_48486,N_48171);
nand U48613 (N_48613,N_48071,N_48300);
or U48614 (N_48614,N_48172,N_48278);
nor U48615 (N_48615,N_48355,N_48098);
or U48616 (N_48616,N_48032,N_48319);
nand U48617 (N_48617,N_48438,N_48157);
xor U48618 (N_48618,N_48479,N_48360);
nand U48619 (N_48619,N_48495,N_48165);
or U48620 (N_48620,N_48498,N_48480);
and U48621 (N_48621,N_48189,N_48084);
nand U48622 (N_48622,N_48197,N_48087);
or U48623 (N_48623,N_48396,N_48307);
xor U48624 (N_48624,N_48050,N_48246);
nor U48625 (N_48625,N_48466,N_48159);
and U48626 (N_48626,N_48267,N_48126);
nand U48627 (N_48627,N_48426,N_48207);
nor U48628 (N_48628,N_48053,N_48465);
nor U48629 (N_48629,N_48452,N_48111);
nor U48630 (N_48630,N_48461,N_48335);
nor U48631 (N_48631,N_48326,N_48000);
or U48632 (N_48632,N_48419,N_48092);
and U48633 (N_48633,N_48017,N_48035);
xor U48634 (N_48634,N_48410,N_48265);
xor U48635 (N_48635,N_48038,N_48287);
xor U48636 (N_48636,N_48272,N_48441);
and U48637 (N_48637,N_48228,N_48242);
nor U48638 (N_48638,N_48318,N_48160);
and U48639 (N_48639,N_48082,N_48496);
nand U48640 (N_48640,N_48369,N_48487);
xnor U48641 (N_48641,N_48200,N_48395);
nand U48642 (N_48642,N_48440,N_48185);
xnor U48643 (N_48643,N_48136,N_48301);
nand U48644 (N_48644,N_48008,N_48151);
nor U48645 (N_48645,N_48196,N_48337);
nor U48646 (N_48646,N_48347,N_48076);
nor U48647 (N_48647,N_48388,N_48336);
nor U48648 (N_48648,N_48004,N_48251);
and U48649 (N_48649,N_48270,N_48003);
nand U48650 (N_48650,N_48028,N_48029);
xor U48651 (N_48651,N_48139,N_48223);
and U48652 (N_48652,N_48416,N_48134);
nor U48653 (N_48653,N_48292,N_48262);
nor U48654 (N_48654,N_48069,N_48011);
nor U48655 (N_48655,N_48244,N_48216);
or U48656 (N_48656,N_48166,N_48107);
and U48657 (N_48657,N_48372,N_48295);
nand U48658 (N_48658,N_48164,N_48373);
xor U48659 (N_48659,N_48021,N_48442);
xor U48660 (N_48660,N_48252,N_48195);
and U48661 (N_48661,N_48046,N_48322);
xor U48662 (N_48662,N_48356,N_48273);
xor U48663 (N_48663,N_48188,N_48381);
nor U48664 (N_48664,N_48370,N_48198);
xor U48665 (N_48665,N_48445,N_48024);
nand U48666 (N_48666,N_48255,N_48081);
and U48667 (N_48667,N_48497,N_48094);
xnor U48668 (N_48668,N_48457,N_48212);
and U48669 (N_48669,N_48261,N_48122);
nand U48670 (N_48670,N_48435,N_48263);
or U48671 (N_48671,N_48343,N_48392);
or U48672 (N_48672,N_48405,N_48334);
nor U48673 (N_48673,N_48454,N_48226);
nor U48674 (N_48674,N_48436,N_48110);
nor U48675 (N_48675,N_48177,N_48102);
xnor U48676 (N_48676,N_48379,N_48250);
nor U48677 (N_48677,N_48163,N_48064);
or U48678 (N_48678,N_48346,N_48079);
and U48679 (N_48679,N_48397,N_48146);
xnor U48680 (N_48680,N_48308,N_48042);
or U48681 (N_48681,N_48075,N_48103);
nor U48682 (N_48682,N_48065,N_48338);
or U48683 (N_48683,N_48232,N_48234);
xnor U48684 (N_48684,N_48421,N_48113);
xor U48685 (N_48685,N_48471,N_48072);
xor U48686 (N_48686,N_48266,N_48125);
nor U48687 (N_48687,N_48484,N_48409);
xnor U48688 (N_48688,N_48462,N_48413);
nor U48689 (N_48689,N_48341,N_48323);
nand U48690 (N_48690,N_48324,N_48306);
nor U48691 (N_48691,N_48229,N_48070);
xor U48692 (N_48692,N_48036,N_48329);
xnor U48693 (N_48693,N_48431,N_48478);
xnor U48694 (N_48694,N_48131,N_48055);
xor U48695 (N_48695,N_48358,N_48333);
nand U48696 (N_48696,N_48363,N_48325);
and U48697 (N_48697,N_48167,N_48161);
nor U48698 (N_48698,N_48135,N_48054);
xor U48699 (N_48699,N_48220,N_48056);
nand U48700 (N_48700,N_48414,N_48380);
or U48701 (N_48701,N_48407,N_48023);
nor U48702 (N_48702,N_48354,N_48399);
xnor U48703 (N_48703,N_48291,N_48152);
nor U48704 (N_48704,N_48009,N_48282);
or U48705 (N_48705,N_48447,N_48088);
and U48706 (N_48706,N_48218,N_48473);
and U48707 (N_48707,N_48458,N_48089);
or U48708 (N_48708,N_48026,N_48469);
xor U48709 (N_48709,N_48077,N_48091);
or U48710 (N_48710,N_48476,N_48437);
and U48711 (N_48711,N_48085,N_48119);
and U48712 (N_48712,N_48147,N_48086);
nand U48713 (N_48713,N_48048,N_48240);
and U48714 (N_48714,N_48169,N_48027);
nor U48715 (N_48715,N_48247,N_48331);
or U48716 (N_48716,N_48470,N_48284);
or U48717 (N_48717,N_48422,N_48310);
nand U48718 (N_48718,N_48057,N_48463);
and U48719 (N_48719,N_48398,N_48289);
and U48720 (N_48720,N_48137,N_48061);
xnor U48721 (N_48721,N_48285,N_48156);
or U48722 (N_48722,N_48404,N_48361);
and U48723 (N_48723,N_48298,N_48280);
or U48724 (N_48724,N_48376,N_48154);
xor U48725 (N_48725,N_48433,N_48312);
nor U48726 (N_48726,N_48408,N_48489);
nor U48727 (N_48727,N_48059,N_48127);
nand U48728 (N_48728,N_48283,N_48389);
or U48729 (N_48729,N_48412,N_48279);
nor U48730 (N_48730,N_48148,N_48235);
or U48731 (N_48731,N_48236,N_48083);
nand U48732 (N_48732,N_48020,N_48006);
and U48733 (N_48733,N_48499,N_48453);
and U48734 (N_48734,N_48352,N_48400);
nand U48735 (N_48735,N_48320,N_48443);
xnor U48736 (N_48736,N_48211,N_48383);
nand U48737 (N_48737,N_48010,N_48428);
and U48738 (N_48738,N_48249,N_48143);
xor U48739 (N_48739,N_48231,N_48045);
nand U48740 (N_48740,N_48417,N_48302);
nand U48741 (N_48741,N_48264,N_48241);
nand U48742 (N_48742,N_48258,N_48230);
nand U48743 (N_48743,N_48425,N_48423);
xnor U48744 (N_48744,N_48439,N_48455);
nor U48745 (N_48745,N_48257,N_48097);
nand U48746 (N_48746,N_48459,N_48213);
and U48747 (N_48747,N_48448,N_48385);
or U48748 (N_48748,N_48044,N_48132);
xnor U48749 (N_48749,N_48187,N_48199);
xor U48750 (N_48750,N_48414,N_48431);
or U48751 (N_48751,N_48137,N_48312);
nand U48752 (N_48752,N_48021,N_48284);
and U48753 (N_48753,N_48143,N_48308);
or U48754 (N_48754,N_48420,N_48080);
or U48755 (N_48755,N_48008,N_48292);
xor U48756 (N_48756,N_48220,N_48319);
nor U48757 (N_48757,N_48199,N_48056);
nor U48758 (N_48758,N_48284,N_48410);
xor U48759 (N_48759,N_48258,N_48265);
xnor U48760 (N_48760,N_48169,N_48003);
and U48761 (N_48761,N_48097,N_48338);
xnor U48762 (N_48762,N_48185,N_48372);
or U48763 (N_48763,N_48282,N_48296);
and U48764 (N_48764,N_48106,N_48375);
nand U48765 (N_48765,N_48434,N_48467);
nand U48766 (N_48766,N_48060,N_48414);
nor U48767 (N_48767,N_48491,N_48190);
or U48768 (N_48768,N_48490,N_48415);
nand U48769 (N_48769,N_48033,N_48484);
and U48770 (N_48770,N_48283,N_48474);
and U48771 (N_48771,N_48399,N_48452);
nand U48772 (N_48772,N_48269,N_48361);
and U48773 (N_48773,N_48044,N_48151);
and U48774 (N_48774,N_48002,N_48009);
and U48775 (N_48775,N_48316,N_48075);
nand U48776 (N_48776,N_48224,N_48466);
xor U48777 (N_48777,N_48155,N_48108);
or U48778 (N_48778,N_48195,N_48454);
nand U48779 (N_48779,N_48238,N_48127);
nor U48780 (N_48780,N_48239,N_48407);
nand U48781 (N_48781,N_48115,N_48429);
and U48782 (N_48782,N_48262,N_48350);
and U48783 (N_48783,N_48346,N_48152);
nor U48784 (N_48784,N_48119,N_48484);
xnor U48785 (N_48785,N_48425,N_48266);
xnor U48786 (N_48786,N_48341,N_48167);
xnor U48787 (N_48787,N_48199,N_48308);
or U48788 (N_48788,N_48097,N_48456);
nand U48789 (N_48789,N_48490,N_48079);
nor U48790 (N_48790,N_48384,N_48151);
nor U48791 (N_48791,N_48004,N_48270);
nand U48792 (N_48792,N_48071,N_48477);
and U48793 (N_48793,N_48339,N_48461);
xnor U48794 (N_48794,N_48061,N_48492);
and U48795 (N_48795,N_48212,N_48106);
and U48796 (N_48796,N_48252,N_48018);
nand U48797 (N_48797,N_48071,N_48221);
xnor U48798 (N_48798,N_48241,N_48065);
nor U48799 (N_48799,N_48363,N_48194);
and U48800 (N_48800,N_48356,N_48290);
xor U48801 (N_48801,N_48119,N_48102);
or U48802 (N_48802,N_48219,N_48395);
and U48803 (N_48803,N_48078,N_48404);
xnor U48804 (N_48804,N_48371,N_48348);
and U48805 (N_48805,N_48246,N_48183);
and U48806 (N_48806,N_48268,N_48247);
nand U48807 (N_48807,N_48039,N_48395);
and U48808 (N_48808,N_48216,N_48473);
or U48809 (N_48809,N_48332,N_48264);
nand U48810 (N_48810,N_48075,N_48423);
xor U48811 (N_48811,N_48485,N_48025);
and U48812 (N_48812,N_48073,N_48149);
xnor U48813 (N_48813,N_48061,N_48087);
nand U48814 (N_48814,N_48335,N_48003);
xnor U48815 (N_48815,N_48164,N_48407);
and U48816 (N_48816,N_48392,N_48175);
nor U48817 (N_48817,N_48281,N_48421);
nor U48818 (N_48818,N_48245,N_48264);
or U48819 (N_48819,N_48238,N_48298);
or U48820 (N_48820,N_48377,N_48200);
nor U48821 (N_48821,N_48073,N_48057);
nand U48822 (N_48822,N_48439,N_48085);
nand U48823 (N_48823,N_48151,N_48121);
xor U48824 (N_48824,N_48334,N_48053);
or U48825 (N_48825,N_48087,N_48027);
nor U48826 (N_48826,N_48332,N_48309);
xnor U48827 (N_48827,N_48271,N_48206);
or U48828 (N_48828,N_48301,N_48129);
or U48829 (N_48829,N_48142,N_48176);
nor U48830 (N_48830,N_48061,N_48408);
nor U48831 (N_48831,N_48442,N_48027);
nand U48832 (N_48832,N_48415,N_48005);
nand U48833 (N_48833,N_48302,N_48361);
xnor U48834 (N_48834,N_48394,N_48027);
nand U48835 (N_48835,N_48033,N_48113);
nand U48836 (N_48836,N_48225,N_48372);
xor U48837 (N_48837,N_48020,N_48029);
and U48838 (N_48838,N_48064,N_48140);
nand U48839 (N_48839,N_48358,N_48092);
nand U48840 (N_48840,N_48301,N_48082);
nor U48841 (N_48841,N_48470,N_48259);
nand U48842 (N_48842,N_48431,N_48215);
and U48843 (N_48843,N_48241,N_48214);
or U48844 (N_48844,N_48028,N_48405);
or U48845 (N_48845,N_48066,N_48095);
xnor U48846 (N_48846,N_48057,N_48024);
nor U48847 (N_48847,N_48256,N_48419);
xor U48848 (N_48848,N_48336,N_48118);
and U48849 (N_48849,N_48367,N_48256);
and U48850 (N_48850,N_48470,N_48409);
nor U48851 (N_48851,N_48327,N_48242);
or U48852 (N_48852,N_48337,N_48262);
nand U48853 (N_48853,N_48299,N_48298);
and U48854 (N_48854,N_48479,N_48332);
nand U48855 (N_48855,N_48098,N_48161);
nor U48856 (N_48856,N_48211,N_48222);
and U48857 (N_48857,N_48019,N_48409);
xnor U48858 (N_48858,N_48200,N_48182);
nand U48859 (N_48859,N_48201,N_48470);
and U48860 (N_48860,N_48383,N_48154);
nand U48861 (N_48861,N_48336,N_48275);
nor U48862 (N_48862,N_48100,N_48364);
nand U48863 (N_48863,N_48197,N_48359);
xnor U48864 (N_48864,N_48064,N_48473);
and U48865 (N_48865,N_48335,N_48341);
and U48866 (N_48866,N_48420,N_48206);
xnor U48867 (N_48867,N_48208,N_48464);
or U48868 (N_48868,N_48492,N_48260);
nor U48869 (N_48869,N_48246,N_48415);
xnor U48870 (N_48870,N_48064,N_48337);
nor U48871 (N_48871,N_48180,N_48381);
nand U48872 (N_48872,N_48110,N_48132);
or U48873 (N_48873,N_48128,N_48377);
nand U48874 (N_48874,N_48343,N_48126);
or U48875 (N_48875,N_48221,N_48268);
nand U48876 (N_48876,N_48296,N_48380);
and U48877 (N_48877,N_48323,N_48089);
xnor U48878 (N_48878,N_48254,N_48468);
xnor U48879 (N_48879,N_48243,N_48134);
and U48880 (N_48880,N_48014,N_48420);
xor U48881 (N_48881,N_48337,N_48454);
and U48882 (N_48882,N_48129,N_48338);
nor U48883 (N_48883,N_48085,N_48448);
or U48884 (N_48884,N_48484,N_48182);
nand U48885 (N_48885,N_48383,N_48156);
nor U48886 (N_48886,N_48375,N_48105);
xor U48887 (N_48887,N_48439,N_48395);
and U48888 (N_48888,N_48473,N_48007);
nand U48889 (N_48889,N_48449,N_48314);
and U48890 (N_48890,N_48334,N_48082);
xor U48891 (N_48891,N_48188,N_48273);
nand U48892 (N_48892,N_48397,N_48147);
nand U48893 (N_48893,N_48488,N_48211);
xnor U48894 (N_48894,N_48381,N_48318);
nand U48895 (N_48895,N_48323,N_48475);
nand U48896 (N_48896,N_48481,N_48373);
xor U48897 (N_48897,N_48373,N_48209);
or U48898 (N_48898,N_48260,N_48271);
nand U48899 (N_48899,N_48281,N_48049);
nand U48900 (N_48900,N_48247,N_48160);
xor U48901 (N_48901,N_48285,N_48466);
xor U48902 (N_48902,N_48106,N_48481);
xor U48903 (N_48903,N_48220,N_48080);
and U48904 (N_48904,N_48164,N_48032);
or U48905 (N_48905,N_48482,N_48071);
nor U48906 (N_48906,N_48408,N_48097);
or U48907 (N_48907,N_48205,N_48380);
nor U48908 (N_48908,N_48243,N_48341);
and U48909 (N_48909,N_48255,N_48162);
nand U48910 (N_48910,N_48016,N_48444);
xnor U48911 (N_48911,N_48302,N_48188);
or U48912 (N_48912,N_48392,N_48312);
nor U48913 (N_48913,N_48138,N_48153);
nor U48914 (N_48914,N_48108,N_48306);
xor U48915 (N_48915,N_48235,N_48319);
nor U48916 (N_48916,N_48247,N_48479);
and U48917 (N_48917,N_48221,N_48289);
nand U48918 (N_48918,N_48231,N_48311);
nand U48919 (N_48919,N_48267,N_48289);
or U48920 (N_48920,N_48060,N_48079);
xor U48921 (N_48921,N_48479,N_48088);
and U48922 (N_48922,N_48484,N_48317);
or U48923 (N_48923,N_48255,N_48342);
xor U48924 (N_48924,N_48491,N_48083);
or U48925 (N_48925,N_48373,N_48039);
nor U48926 (N_48926,N_48460,N_48477);
nor U48927 (N_48927,N_48035,N_48475);
xor U48928 (N_48928,N_48318,N_48071);
or U48929 (N_48929,N_48312,N_48329);
xnor U48930 (N_48930,N_48210,N_48485);
xnor U48931 (N_48931,N_48395,N_48088);
xor U48932 (N_48932,N_48389,N_48273);
nand U48933 (N_48933,N_48030,N_48142);
and U48934 (N_48934,N_48218,N_48178);
xor U48935 (N_48935,N_48350,N_48420);
nor U48936 (N_48936,N_48424,N_48088);
and U48937 (N_48937,N_48244,N_48318);
xnor U48938 (N_48938,N_48031,N_48115);
or U48939 (N_48939,N_48047,N_48415);
and U48940 (N_48940,N_48094,N_48324);
nor U48941 (N_48941,N_48412,N_48393);
and U48942 (N_48942,N_48305,N_48497);
and U48943 (N_48943,N_48322,N_48088);
and U48944 (N_48944,N_48269,N_48247);
xor U48945 (N_48945,N_48033,N_48149);
and U48946 (N_48946,N_48426,N_48052);
nor U48947 (N_48947,N_48241,N_48396);
xor U48948 (N_48948,N_48239,N_48456);
and U48949 (N_48949,N_48033,N_48402);
xnor U48950 (N_48950,N_48421,N_48422);
and U48951 (N_48951,N_48354,N_48412);
nand U48952 (N_48952,N_48354,N_48230);
or U48953 (N_48953,N_48353,N_48140);
and U48954 (N_48954,N_48413,N_48436);
or U48955 (N_48955,N_48192,N_48077);
and U48956 (N_48956,N_48483,N_48175);
and U48957 (N_48957,N_48350,N_48359);
and U48958 (N_48958,N_48375,N_48020);
or U48959 (N_48959,N_48383,N_48339);
or U48960 (N_48960,N_48056,N_48454);
nor U48961 (N_48961,N_48437,N_48001);
nor U48962 (N_48962,N_48245,N_48105);
nor U48963 (N_48963,N_48148,N_48454);
nand U48964 (N_48964,N_48448,N_48360);
nor U48965 (N_48965,N_48222,N_48300);
xor U48966 (N_48966,N_48167,N_48452);
and U48967 (N_48967,N_48415,N_48019);
xnor U48968 (N_48968,N_48461,N_48490);
or U48969 (N_48969,N_48204,N_48237);
or U48970 (N_48970,N_48328,N_48098);
and U48971 (N_48971,N_48092,N_48171);
nand U48972 (N_48972,N_48290,N_48143);
or U48973 (N_48973,N_48079,N_48319);
xnor U48974 (N_48974,N_48398,N_48401);
nor U48975 (N_48975,N_48110,N_48273);
xnor U48976 (N_48976,N_48221,N_48449);
xnor U48977 (N_48977,N_48300,N_48354);
or U48978 (N_48978,N_48379,N_48071);
xnor U48979 (N_48979,N_48405,N_48383);
or U48980 (N_48980,N_48472,N_48391);
and U48981 (N_48981,N_48310,N_48347);
or U48982 (N_48982,N_48380,N_48482);
xor U48983 (N_48983,N_48356,N_48157);
and U48984 (N_48984,N_48364,N_48144);
or U48985 (N_48985,N_48175,N_48387);
xnor U48986 (N_48986,N_48435,N_48172);
nor U48987 (N_48987,N_48131,N_48398);
and U48988 (N_48988,N_48361,N_48235);
nand U48989 (N_48989,N_48470,N_48134);
and U48990 (N_48990,N_48242,N_48184);
nor U48991 (N_48991,N_48488,N_48013);
or U48992 (N_48992,N_48072,N_48012);
and U48993 (N_48993,N_48459,N_48054);
or U48994 (N_48994,N_48325,N_48071);
xor U48995 (N_48995,N_48386,N_48073);
nand U48996 (N_48996,N_48381,N_48197);
nor U48997 (N_48997,N_48048,N_48129);
and U48998 (N_48998,N_48139,N_48010);
xor U48999 (N_48999,N_48157,N_48181);
and U49000 (N_49000,N_48503,N_48551);
nand U49001 (N_49001,N_48658,N_48747);
nand U49002 (N_49002,N_48715,N_48543);
or U49003 (N_49003,N_48893,N_48524);
and U49004 (N_49004,N_48765,N_48668);
xor U49005 (N_49005,N_48937,N_48995);
nor U49006 (N_49006,N_48904,N_48771);
nand U49007 (N_49007,N_48990,N_48667);
and U49008 (N_49008,N_48812,N_48623);
and U49009 (N_49009,N_48870,N_48615);
nand U49010 (N_49010,N_48819,N_48565);
xor U49011 (N_49011,N_48519,N_48829);
xnor U49012 (N_49012,N_48982,N_48891);
xnor U49013 (N_49013,N_48730,N_48506);
or U49014 (N_49014,N_48802,N_48756);
nor U49015 (N_49015,N_48627,N_48619);
and U49016 (N_49016,N_48865,N_48897);
and U49017 (N_49017,N_48626,N_48996);
or U49018 (N_49018,N_48635,N_48523);
or U49019 (N_49019,N_48844,N_48846);
or U49020 (N_49020,N_48835,N_48535);
nand U49021 (N_49021,N_48559,N_48942);
nor U49022 (N_49022,N_48707,N_48872);
and U49023 (N_49023,N_48815,N_48590);
xnor U49024 (N_49024,N_48818,N_48640);
and U49025 (N_49025,N_48936,N_48515);
nor U49026 (N_49026,N_48855,N_48783);
nand U49027 (N_49027,N_48949,N_48605);
and U49028 (N_49028,N_48613,N_48510);
and U49029 (N_49029,N_48621,N_48595);
and U49030 (N_49030,N_48769,N_48951);
xnor U49031 (N_49031,N_48702,N_48881);
and U49032 (N_49032,N_48629,N_48743);
nor U49033 (N_49033,N_48918,N_48649);
nor U49034 (N_49034,N_48789,N_48761);
or U49035 (N_49035,N_48900,N_48563);
and U49036 (N_49036,N_48796,N_48955);
and U49037 (N_49037,N_48727,N_48974);
and U49038 (N_49038,N_48999,N_48839);
xor U49039 (N_49039,N_48977,N_48801);
or U49040 (N_49040,N_48957,N_48689);
or U49041 (N_49041,N_48913,N_48699);
nand U49042 (N_49042,N_48708,N_48901);
and U49043 (N_49043,N_48916,N_48539);
or U49044 (N_49044,N_48726,N_48827);
nor U49045 (N_49045,N_48764,N_48928);
nand U49046 (N_49046,N_48687,N_48873);
xor U49047 (N_49047,N_48571,N_48500);
nor U49048 (N_49048,N_48542,N_48863);
nand U49049 (N_49049,N_48509,N_48940);
or U49050 (N_49050,N_48603,N_48958);
nand U49051 (N_49051,N_48867,N_48666);
and U49052 (N_49052,N_48596,N_48722);
nor U49053 (N_49053,N_48665,N_48947);
nor U49054 (N_49054,N_48734,N_48856);
or U49055 (N_49055,N_48610,N_48880);
or U49056 (N_49056,N_48507,N_48832);
nand U49057 (N_49057,N_48575,N_48987);
or U49058 (N_49058,N_48800,N_48549);
and U49059 (N_49059,N_48755,N_48532);
nor U49060 (N_49060,N_48816,N_48840);
nor U49061 (N_49061,N_48676,N_48577);
nor U49062 (N_49062,N_48860,N_48866);
or U49063 (N_49063,N_48879,N_48930);
xnor U49064 (N_49064,N_48671,N_48922);
nor U49065 (N_49065,N_48620,N_48959);
nor U49066 (N_49066,N_48625,N_48975);
xor U49067 (N_49067,N_48562,N_48622);
nand U49068 (N_49068,N_48710,N_48868);
nand U49069 (N_49069,N_48717,N_48541);
nand U49070 (N_49070,N_48908,N_48883);
xor U49071 (N_49071,N_48616,N_48588);
and U49072 (N_49072,N_48754,N_48617);
xor U49073 (N_49073,N_48723,N_48932);
or U49074 (N_49074,N_48703,N_48910);
and U49075 (N_49075,N_48886,N_48560);
nor U49076 (N_49076,N_48534,N_48614);
nor U49077 (N_49077,N_48552,N_48749);
or U49078 (N_49078,N_48953,N_48646);
nor U49079 (N_49079,N_48971,N_48825);
or U49080 (N_49080,N_48858,N_48774);
or U49081 (N_49081,N_48998,N_48721);
or U49082 (N_49082,N_48760,N_48701);
and U49083 (N_49083,N_48594,N_48972);
xnor U49084 (N_49084,N_48821,N_48954);
xnor U49085 (N_49085,N_48598,N_48655);
and U49086 (N_49086,N_48669,N_48573);
xor U49087 (N_49087,N_48536,N_48763);
and U49088 (N_49088,N_48989,N_48714);
nand U49089 (N_49089,N_48944,N_48554);
nand U49090 (N_49090,N_48602,N_48528);
or U49091 (N_49091,N_48583,N_48700);
and U49092 (N_49092,N_48798,N_48962);
xor U49093 (N_49093,N_48823,N_48768);
and U49094 (N_49094,N_48529,N_48806);
and U49095 (N_49095,N_48512,N_48567);
nor U49096 (N_49096,N_48853,N_48965);
nand U49097 (N_49097,N_48729,N_48793);
xnor U49098 (N_49098,N_48612,N_48585);
nand U49099 (N_49099,N_48837,N_48683);
and U49100 (N_49100,N_48943,N_48511);
and U49101 (N_49101,N_48690,N_48555);
nand U49102 (N_49102,N_48847,N_48653);
nand U49103 (N_49103,N_48546,N_48976);
xor U49104 (N_49104,N_48637,N_48917);
xnor U49105 (N_49105,N_48762,N_48923);
and U49106 (N_49106,N_48663,N_48788);
nand U49107 (N_49107,N_48890,N_48804);
xnor U49108 (N_49108,N_48744,N_48630);
or U49109 (N_49109,N_48750,N_48961);
xor U49110 (N_49110,N_48877,N_48556);
xor U49111 (N_49111,N_48533,N_48952);
xor U49112 (N_49112,N_48724,N_48903);
xnor U49113 (N_49113,N_48862,N_48960);
and U49114 (N_49114,N_48914,N_48824);
nor U49115 (N_49115,N_48887,N_48579);
nand U49116 (N_49116,N_48894,N_48647);
or U49117 (N_49117,N_48878,N_48526);
nor U49118 (N_49118,N_48624,N_48841);
nand U49119 (N_49119,N_48662,N_48697);
nor U49120 (N_49120,N_48516,N_48664);
nor U49121 (N_49121,N_48651,N_48912);
nand U49122 (N_49122,N_48979,N_48831);
xor U49123 (N_49123,N_48681,N_48520);
or U49124 (N_49124,N_48656,N_48591);
nand U49125 (N_49125,N_48686,N_48898);
and U49126 (N_49126,N_48692,N_48738);
xnor U49127 (N_49127,N_48736,N_48808);
and U49128 (N_49128,N_48902,N_48570);
nor U49129 (N_49129,N_48696,N_48836);
nand U49130 (N_49130,N_48964,N_48733);
nor U49131 (N_49131,N_48935,N_48527);
and U49132 (N_49132,N_48748,N_48680);
nand U49133 (N_49133,N_48892,N_48777);
or U49134 (N_49134,N_48850,N_48864);
nand U49135 (N_49135,N_48633,N_48857);
and U49136 (N_49136,N_48973,N_48817);
nand U49137 (N_49137,N_48911,N_48589);
xnor U49138 (N_49138,N_48779,N_48548);
nor U49139 (N_49139,N_48948,N_48618);
xor U49140 (N_49140,N_48550,N_48843);
and U49141 (N_49141,N_48746,N_48606);
or U49142 (N_49142,N_48628,N_48776);
nand U49143 (N_49143,N_48608,N_48632);
or U49144 (N_49144,N_48650,N_48826);
and U49145 (N_49145,N_48909,N_48518);
nor U49146 (N_49146,N_48593,N_48713);
and U49147 (N_49147,N_48688,N_48674);
and U49148 (N_49148,N_48716,N_48791);
and U49149 (N_49149,N_48992,N_48660);
or U49150 (N_49150,N_48934,N_48884);
xnor U49151 (N_49151,N_48871,N_48905);
nor U49152 (N_49152,N_48672,N_48581);
nand U49153 (N_49153,N_48530,N_48631);
nor U49154 (N_49154,N_48963,N_48787);
and U49155 (N_49155,N_48654,N_48986);
nor U49156 (N_49156,N_48670,N_48557);
or U49157 (N_49157,N_48600,N_48792);
or U49158 (N_49158,N_48673,N_48525);
xor U49159 (N_49159,N_48807,N_48978);
nand U49160 (N_49160,N_48876,N_48742);
xnor U49161 (N_49161,N_48704,N_48694);
nand U49162 (N_49162,N_48712,N_48641);
or U49163 (N_49163,N_48770,N_48741);
or U49164 (N_49164,N_48517,N_48767);
and U49165 (N_49165,N_48725,N_48657);
xnor U49166 (N_49166,N_48502,N_48849);
and U49167 (N_49167,N_48514,N_48969);
nor U49168 (N_49168,N_48785,N_48985);
and U49169 (N_49169,N_48820,N_48582);
and U49170 (N_49170,N_48643,N_48587);
xnor U49171 (N_49171,N_48848,N_48574);
or U49172 (N_49172,N_48899,N_48970);
xor U49173 (N_49173,N_48569,N_48693);
nor U49174 (N_49174,N_48597,N_48981);
and U49175 (N_49175,N_48652,N_48709);
or U49176 (N_49176,N_48967,N_48926);
nand U49177 (N_49177,N_48984,N_48685);
or U49178 (N_49178,N_48920,N_48566);
nand U49179 (N_49179,N_48636,N_48698);
nand U49180 (N_49180,N_48732,N_48759);
nor U49181 (N_49181,N_48945,N_48997);
nor U49182 (N_49182,N_48838,N_48691);
xnor U49183 (N_49183,N_48859,N_48719);
and U49184 (N_49184,N_48834,N_48572);
and U49185 (N_49185,N_48811,N_48980);
and U49186 (N_49186,N_48682,N_48993);
xor U49187 (N_49187,N_48941,N_48956);
nor U49188 (N_49188,N_48983,N_48513);
nor U49189 (N_49189,N_48584,N_48896);
nand U49190 (N_49190,N_48861,N_48521);
xor U49191 (N_49191,N_48828,N_48639);
nand U49192 (N_49192,N_48659,N_48813);
xnor U49193 (N_49193,N_48677,N_48580);
or U49194 (N_49194,N_48609,N_48786);
or U49195 (N_49195,N_48924,N_48805);
and U49196 (N_49196,N_48578,N_48780);
or U49197 (N_49197,N_48875,N_48505);
or U49198 (N_49198,N_48814,N_48946);
or U49199 (N_49199,N_48753,N_48933);
xor U49200 (N_49200,N_48939,N_48558);
or U49201 (N_49201,N_48869,N_48803);
nor U49202 (N_49202,N_48695,N_48751);
nand U49203 (N_49203,N_48739,N_48851);
nand U49204 (N_49204,N_48784,N_48508);
and U49205 (N_49205,N_48718,N_48852);
nand U49206 (N_49206,N_48799,N_48994);
or U49207 (N_49207,N_48797,N_48711);
nand U49208 (N_49208,N_48830,N_48906);
or U49209 (N_49209,N_48545,N_48772);
or U49210 (N_49210,N_48919,N_48678);
xor U49211 (N_49211,N_48586,N_48684);
nor U49212 (N_49212,N_48925,N_48611);
and U49213 (N_49213,N_48795,N_48988);
or U49214 (N_49214,N_48790,N_48929);
nor U49215 (N_49215,N_48645,N_48822);
nor U49216 (N_49216,N_48842,N_48504);
nor U49217 (N_49217,N_48931,N_48745);
or U49218 (N_49218,N_48531,N_48921);
nor U49219 (N_49219,N_48889,N_48644);
nor U49220 (N_49220,N_48915,N_48576);
nor U49221 (N_49221,N_48547,N_48679);
and U49222 (N_49222,N_48833,N_48540);
or U49223 (N_49223,N_48794,N_48553);
xnor U49224 (N_49224,N_48778,N_48599);
and U49225 (N_49225,N_48882,N_48501);
nand U49226 (N_49226,N_48991,N_48938);
or U49227 (N_49227,N_48706,N_48564);
xor U49228 (N_49228,N_48874,N_48601);
nand U49229 (N_49229,N_48766,N_48607);
nor U49230 (N_49230,N_48642,N_48810);
or U49231 (N_49231,N_48638,N_48752);
or U49232 (N_49232,N_48773,N_48661);
nand U49233 (N_49233,N_48592,N_48728);
nand U49234 (N_49234,N_48544,N_48538);
xor U49235 (N_49235,N_48757,N_48781);
nand U49236 (N_49236,N_48950,N_48809);
xor U49237 (N_49237,N_48522,N_48731);
or U49238 (N_49238,N_48740,N_48720);
and U49239 (N_49239,N_48907,N_48561);
xor U49240 (N_49240,N_48735,N_48888);
nor U49241 (N_49241,N_48845,N_48966);
and U49242 (N_49242,N_48537,N_48758);
xor U49243 (N_49243,N_48604,N_48775);
xnor U49244 (N_49244,N_48927,N_48634);
and U49245 (N_49245,N_48648,N_48737);
and U49246 (N_49246,N_48675,N_48885);
and U49247 (N_49247,N_48895,N_48854);
and U49248 (N_49248,N_48968,N_48568);
nand U49249 (N_49249,N_48782,N_48705);
or U49250 (N_49250,N_48742,N_48601);
and U49251 (N_49251,N_48871,N_48627);
nor U49252 (N_49252,N_48873,N_48786);
and U49253 (N_49253,N_48679,N_48623);
xnor U49254 (N_49254,N_48542,N_48605);
or U49255 (N_49255,N_48774,N_48510);
or U49256 (N_49256,N_48664,N_48645);
or U49257 (N_49257,N_48627,N_48725);
xnor U49258 (N_49258,N_48861,N_48806);
xor U49259 (N_49259,N_48913,N_48644);
nor U49260 (N_49260,N_48616,N_48734);
xnor U49261 (N_49261,N_48803,N_48881);
nand U49262 (N_49262,N_48728,N_48813);
xor U49263 (N_49263,N_48649,N_48621);
nor U49264 (N_49264,N_48722,N_48885);
nor U49265 (N_49265,N_48721,N_48994);
nand U49266 (N_49266,N_48737,N_48582);
nand U49267 (N_49267,N_48727,N_48918);
nand U49268 (N_49268,N_48790,N_48566);
nand U49269 (N_49269,N_48593,N_48794);
nor U49270 (N_49270,N_48718,N_48961);
nor U49271 (N_49271,N_48750,N_48558);
nor U49272 (N_49272,N_48702,N_48792);
and U49273 (N_49273,N_48882,N_48982);
or U49274 (N_49274,N_48796,N_48798);
nand U49275 (N_49275,N_48817,N_48897);
or U49276 (N_49276,N_48537,N_48635);
xor U49277 (N_49277,N_48782,N_48553);
nor U49278 (N_49278,N_48539,N_48780);
xnor U49279 (N_49279,N_48743,N_48995);
and U49280 (N_49280,N_48557,N_48820);
or U49281 (N_49281,N_48892,N_48625);
and U49282 (N_49282,N_48688,N_48758);
nor U49283 (N_49283,N_48625,N_48771);
and U49284 (N_49284,N_48684,N_48963);
and U49285 (N_49285,N_48791,N_48851);
xnor U49286 (N_49286,N_48676,N_48721);
nor U49287 (N_49287,N_48718,N_48641);
or U49288 (N_49288,N_48542,N_48820);
xor U49289 (N_49289,N_48827,N_48858);
and U49290 (N_49290,N_48886,N_48768);
or U49291 (N_49291,N_48579,N_48543);
and U49292 (N_49292,N_48867,N_48825);
xnor U49293 (N_49293,N_48682,N_48612);
xor U49294 (N_49294,N_48866,N_48831);
nand U49295 (N_49295,N_48524,N_48982);
nand U49296 (N_49296,N_48852,N_48538);
nand U49297 (N_49297,N_48878,N_48987);
and U49298 (N_49298,N_48522,N_48990);
nor U49299 (N_49299,N_48754,N_48905);
and U49300 (N_49300,N_48991,N_48613);
or U49301 (N_49301,N_48851,N_48583);
and U49302 (N_49302,N_48898,N_48670);
nor U49303 (N_49303,N_48877,N_48733);
nor U49304 (N_49304,N_48586,N_48978);
xor U49305 (N_49305,N_48527,N_48900);
xnor U49306 (N_49306,N_48589,N_48978);
or U49307 (N_49307,N_48524,N_48512);
xor U49308 (N_49308,N_48526,N_48784);
nor U49309 (N_49309,N_48518,N_48694);
or U49310 (N_49310,N_48885,N_48529);
nor U49311 (N_49311,N_48614,N_48908);
and U49312 (N_49312,N_48928,N_48989);
nand U49313 (N_49313,N_48812,N_48952);
xor U49314 (N_49314,N_48991,N_48842);
nand U49315 (N_49315,N_48873,N_48905);
nand U49316 (N_49316,N_48547,N_48616);
nand U49317 (N_49317,N_48945,N_48683);
nor U49318 (N_49318,N_48632,N_48595);
xnor U49319 (N_49319,N_48526,N_48533);
or U49320 (N_49320,N_48644,N_48741);
and U49321 (N_49321,N_48891,N_48859);
nand U49322 (N_49322,N_48979,N_48668);
nor U49323 (N_49323,N_48532,N_48942);
or U49324 (N_49324,N_48965,N_48557);
or U49325 (N_49325,N_48897,N_48598);
nor U49326 (N_49326,N_48514,N_48906);
nor U49327 (N_49327,N_48941,N_48811);
nand U49328 (N_49328,N_48692,N_48857);
nor U49329 (N_49329,N_48585,N_48863);
nand U49330 (N_49330,N_48539,N_48706);
nor U49331 (N_49331,N_48686,N_48757);
and U49332 (N_49332,N_48904,N_48814);
or U49333 (N_49333,N_48998,N_48584);
xor U49334 (N_49334,N_48931,N_48669);
nor U49335 (N_49335,N_48896,N_48856);
nand U49336 (N_49336,N_48773,N_48651);
nor U49337 (N_49337,N_48529,N_48808);
nand U49338 (N_49338,N_48987,N_48533);
nand U49339 (N_49339,N_48825,N_48972);
nand U49340 (N_49340,N_48535,N_48795);
nand U49341 (N_49341,N_48631,N_48730);
xor U49342 (N_49342,N_48779,N_48520);
xor U49343 (N_49343,N_48799,N_48800);
or U49344 (N_49344,N_48924,N_48960);
nor U49345 (N_49345,N_48723,N_48846);
and U49346 (N_49346,N_48707,N_48534);
and U49347 (N_49347,N_48791,N_48526);
or U49348 (N_49348,N_48925,N_48809);
or U49349 (N_49349,N_48983,N_48832);
xnor U49350 (N_49350,N_48789,N_48667);
nand U49351 (N_49351,N_48883,N_48939);
nand U49352 (N_49352,N_48555,N_48926);
or U49353 (N_49353,N_48732,N_48701);
xnor U49354 (N_49354,N_48527,N_48746);
xnor U49355 (N_49355,N_48716,N_48645);
nor U49356 (N_49356,N_48639,N_48802);
xor U49357 (N_49357,N_48538,N_48740);
nor U49358 (N_49358,N_48686,N_48730);
xnor U49359 (N_49359,N_48738,N_48640);
xor U49360 (N_49360,N_48702,N_48889);
or U49361 (N_49361,N_48658,N_48573);
or U49362 (N_49362,N_48524,N_48872);
and U49363 (N_49363,N_48705,N_48565);
and U49364 (N_49364,N_48886,N_48791);
xor U49365 (N_49365,N_48588,N_48866);
xnor U49366 (N_49366,N_48652,N_48939);
nand U49367 (N_49367,N_48822,N_48983);
xor U49368 (N_49368,N_48519,N_48848);
or U49369 (N_49369,N_48970,N_48983);
or U49370 (N_49370,N_48562,N_48865);
and U49371 (N_49371,N_48643,N_48652);
xor U49372 (N_49372,N_48926,N_48560);
and U49373 (N_49373,N_48521,N_48669);
and U49374 (N_49374,N_48828,N_48966);
nand U49375 (N_49375,N_48825,N_48589);
nand U49376 (N_49376,N_48954,N_48697);
nand U49377 (N_49377,N_48710,N_48899);
or U49378 (N_49378,N_48575,N_48776);
nand U49379 (N_49379,N_48636,N_48907);
nor U49380 (N_49380,N_48735,N_48628);
xor U49381 (N_49381,N_48650,N_48789);
xnor U49382 (N_49382,N_48671,N_48815);
or U49383 (N_49383,N_48793,N_48592);
nand U49384 (N_49384,N_48758,N_48892);
nor U49385 (N_49385,N_48749,N_48687);
nand U49386 (N_49386,N_48986,N_48818);
and U49387 (N_49387,N_48677,N_48524);
and U49388 (N_49388,N_48556,N_48885);
nor U49389 (N_49389,N_48706,N_48953);
or U49390 (N_49390,N_48654,N_48502);
nor U49391 (N_49391,N_48678,N_48567);
or U49392 (N_49392,N_48680,N_48912);
nand U49393 (N_49393,N_48501,N_48757);
and U49394 (N_49394,N_48575,N_48839);
nand U49395 (N_49395,N_48653,N_48728);
and U49396 (N_49396,N_48549,N_48973);
and U49397 (N_49397,N_48594,N_48748);
nand U49398 (N_49398,N_48618,N_48615);
nor U49399 (N_49399,N_48927,N_48940);
nand U49400 (N_49400,N_48503,N_48692);
or U49401 (N_49401,N_48966,N_48817);
nand U49402 (N_49402,N_48993,N_48692);
or U49403 (N_49403,N_48769,N_48893);
nand U49404 (N_49404,N_48960,N_48792);
and U49405 (N_49405,N_48909,N_48831);
xor U49406 (N_49406,N_48760,N_48583);
nand U49407 (N_49407,N_48545,N_48751);
and U49408 (N_49408,N_48826,N_48673);
or U49409 (N_49409,N_48979,N_48542);
and U49410 (N_49410,N_48765,N_48844);
nand U49411 (N_49411,N_48582,N_48705);
xor U49412 (N_49412,N_48671,N_48684);
nor U49413 (N_49413,N_48796,N_48764);
xnor U49414 (N_49414,N_48641,N_48614);
and U49415 (N_49415,N_48641,N_48600);
or U49416 (N_49416,N_48656,N_48755);
nand U49417 (N_49417,N_48981,N_48967);
nor U49418 (N_49418,N_48951,N_48758);
nand U49419 (N_49419,N_48619,N_48800);
nor U49420 (N_49420,N_48833,N_48998);
xor U49421 (N_49421,N_48550,N_48928);
and U49422 (N_49422,N_48581,N_48509);
nor U49423 (N_49423,N_48874,N_48708);
or U49424 (N_49424,N_48953,N_48815);
or U49425 (N_49425,N_48627,N_48772);
nor U49426 (N_49426,N_48732,N_48727);
or U49427 (N_49427,N_48954,N_48798);
xor U49428 (N_49428,N_48675,N_48849);
nand U49429 (N_49429,N_48545,N_48620);
xor U49430 (N_49430,N_48712,N_48640);
or U49431 (N_49431,N_48799,N_48884);
nor U49432 (N_49432,N_48690,N_48907);
xnor U49433 (N_49433,N_48640,N_48617);
xnor U49434 (N_49434,N_48728,N_48557);
nand U49435 (N_49435,N_48514,N_48599);
xor U49436 (N_49436,N_48708,N_48945);
xor U49437 (N_49437,N_48911,N_48938);
or U49438 (N_49438,N_48558,N_48777);
xnor U49439 (N_49439,N_48616,N_48674);
nor U49440 (N_49440,N_48715,N_48869);
nor U49441 (N_49441,N_48980,N_48503);
nor U49442 (N_49442,N_48707,N_48547);
or U49443 (N_49443,N_48853,N_48606);
and U49444 (N_49444,N_48783,N_48658);
xor U49445 (N_49445,N_48516,N_48546);
or U49446 (N_49446,N_48863,N_48934);
nand U49447 (N_49447,N_48907,N_48770);
nor U49448 (N_49448,N_48675,N_48554);
nor U49449 (N_49449,N_48825,N_48849);
or U49450 (N_49450,N_48680,N_48954);
nand U49451 (N_49451,N_48736,N_48514);
xnor U49452 (N_49452,N_48753,N_48776);
xnor U49453 (N_49453,N_48751,N_48626);
nand U49454 (N_49454,N_48699,N_48624);
or U49455 (N_49455,N_48672,N_48945);
nand U49456 (N_49456,N_48915,N_48858);
and U49457 (N_49457,N_48701,N_48537);
nor U49458 (N_49458,N_48576,N_48752);
or U49459 (N_49459,N_48843,N_48661);
nand U49460 (N_49460,N_48902,N_48817);
or U49461 (N_49461,N_48888,N_48931);
and U49462 (N_49462,N_48512,N_48900);
or U49463 (N_49463,N_48614,N_48769);
nand U49464 (N_49464,N_48883,N_48877);
and U49465 (N_49465,N_48828,N_48613);
nand U49466 (N_49466,N_48792,N_48998);
nand U49467 (N_49467,N_48871,N_48863);
xor U49468 (N_49468,N_48684,N_48929);
or U49469 (N_49469,N_48741,N_48943);
xnor U49470 (N_49470,N_48781,N_48588);
nand U49471 (N_49471,N_48904,N_48614);
nor U49472 (N_49472,N_48822,N_48502);
nand U49473 (N_49473,N_48614,N_48559);
or U49474 (N_49474,N_48749,N_48763);
and U49475 (N_49475,N_48809,N_48634);
or U49476 (N_49476,N_48976,N_48690);
and U49477 (N_49477,N_48582,N_48599);
or U49478 (N_49478,N_48883,N_48552);
nand U49479 (N_49479,N_48941,N_48617);
or U49480 (N_49480,N_48892,N_48960);
xor U49481 (N_49481,N_48747,N_48609);
and U49482 (N_49482,N_48838,N_48558);
xnor U49483 (N_49483,N_48730,N_48867);
or U49484 (N_49484,N_48843,N_48621);
or U49485 (N_49485,N_48711,N_48988);
nand U49486 (N_49486,N_48675,N_48708);
nand U49487 (N_49487,N_48972,N_48859);
and U49488 (N_49488,N_48994,N_48658);
and U49489 (N_49489,N_48939,N_48552);
nor U49490 (N_49490,N_48794,N_48813);
or U49491 (N_49491,N_48715,N_48638);
xor U49492 (N_49492,N_48908,N_48514);
nand U49493 (N_49493,N_48691,N_48730);
nand U49494 (N_49494,N_48570,N_48986);
xnor U49495 (N_49495,N_48808,N_48734);
or U49496 (N_49496,N_48890,N_48717);
or U49497 (N_49497,N_48612,N_48712);
xor U49498 (N_49498,N_48751,N_48697);
nand U49499 (N_49499,N_48975,N_48919);
or U49500 (N_49500,N_49481,N_49315);
nor U49501 (N_49501,N_49178,N_49430);
nand U49502 (N_49502,N_49112,N_49389);
nand U49503 (N_49503,N_49130,N_49199);
nand U49504 (N_49504,N_49233,N_49158);
or U49505 (N_49505,N_49181,N_49168);
and U49506 (N_49506,N_49426,N_49323);
and U49507 (N_49507,N_49296,N_49206);
nand U49508 (N_49508,N_49232,N_49342);
nor U49509 (N_49509,N_49444,N_49380);
xnor U49510 (N_49510,N_49121,N_49048);
xnor U49511 (N_49511,N_49093,N_49462);
nor U49512 (N_49512,N_49212,N_49194);
nand U49513 (N_49513,N_49150,N_49231);
nor U49514 (N_49514,N_49155,N_49031);
and U49515 (N_49515,N_49077,N_49053);
xor U49516 (N_49516,N_49289,N_49018);
and U49517 (N_49517,N_49271,N_49468);
and U49518 (N_49518,N_49407,N_49151);
nand U49519 (N_49519,N_49333,N_49131);
nand U49520 (N_49520,N_49344,N_49080);
nor U49521 (N_49521,N_49331,N_49105);
or U49522 (N_49522,N_49184,N_49498);
nand U49523 (N_49523,N_49237,N_49379);
and U49524 (N_49524,N_49182,N_49371);
xor U49525 (N_49525,N_49055,N_49147);
nor U49526 (N_49526,N_49397,N_49076);
xnor U49527 (N_49527,N_49453,N_49224);
nor U49528 (N_49528,N_49293,N_49338);
nor U49529 (N_49529,N_49424,N_49364);
nor U49530 (N_49530,N_49256,N_49134);
xor U49531 (N_49531,N_49169,N_49035);
nor U49532 (N_49532,N_49038,N_49026);
xor U49533 (N_49533,N_49287,N_49272);
or U49534 (N_49534,N_49395,N_49264);
and U49535 (N_49535,N_49402,N_49316);
nor U49536 (N_49536,N_49477,N_49399);
nand U49537 (N_49537,N_49259,N_49409);
xnor U49538 (N_49538,N_49085,N_49154);
and U49539 (N_49539,N_49336,N_49177);
and U49540 (N_49540,N_49023,N_49161);
xnor U49541 (N_49541,N_49291,N_49490);
and U49542 (N_49542,N_49072,N_49068);
nor U49543 (N_49543,N_49001,N_49408);
nand U49544 (N_49544,N_49183,N_49386);
nor U49545 (N_49545,N_49006,N_49273);
nor U49546 (N_49546,N_49017,N_49449);
and U49547 (N_49547,N_49180,N_49227);
and U49548 (N_49548,N_49210,N_49170);
nand U49549 (N_49549,N_49050,N_49304);
xor U49550 (N_49550,N_49089,N_49146);
xor U49551 (N_49551,N_49175,N_49135);
or U49552 (N_49552,N_49419,N_49470);
xor U49553 (N_49553,N_49120,N_49042);
nand U49554 (N_49554,N_49142,N_49197);
and U49555 (N_49555,N_49110,N_49459);
and U49556 (N_49556,N_49025,N_49241);
or U49557 (N_49557,N_49473,N_49354);
nand U49558 (N_49558,N_49179,N_49450);
nand U49559 (N_49559,N_49024,N_49270);
xor U49560 (N_49560,N_49357,N_49176);
nand U49561 (N_49561,N_49061,N_49242);
or U49562 (N_49562,N_49356,N_49465);
nor U49563 (N_49563,N_49172,N_49153);
xnor U49564 (N_49564,N_49167,N_49229);
nor U49565 (N_49565,N_49369,N_49084);
nor U49566 (N_49566,N_49013,N_49116);
nor U49567 (N_49567,N_49464,N_49491);
xor U49568 (N_49568,N_49349,N_49051);
and U49569 (N_49569,N_49215,N_49137);
or U49570 (N_49570,N_49128,N_49448);
or U49571 (N_49571,N_49149,N_49162);
xor U49572 (N_49572,N_49095,N_49418);
and U49573 (N_49573,N_49253,N_49127);
or U49574 (N_49574,N_49226,N_49066);
xor U49575 (N_49575,N_49204,N_49405);
nand U49576 (N_49576,N_49415,N_49340);
nor U49577 (N_49577,N_49099,N_49251);
nor U49578 (N_49578,N_49351,N_49214);
and U49579 (N_49579,N_49455,N_49325);
and U49580 (N_49580,N_49207,N_49329);
and U49581 (N_49581,N_49058,N_49339);
or U49582 (N_49582,N_49070,N_49432);
and U49583 (N_49583,N_49148,N_49119);
or U49584 (N_49584,N_49159,N_49312);
nand U49585 (N_49585,N_49484,N_49348);
and U49586 (N_49586,N_49046,N_49276);
nand U49587 (N_49587,N_49486,N_49103);
or U49588 (N_49588,N_49274,N_49497);
xnor U49589 (N_49589,N_49187,N_49311);
or U49590 (N_49590,N_49203,N_49301);
nand U49591 (N_49591,N_49236,N_49009);
and U49592 (N_49592,N_49345,N_49300);
xor U49593 (N_49593,N_49361,N_49234);
nand U49594 (N_49594,N_49143,N_49447);
nand U49595 (N_49595,N_49263,N_49420);
xor U49596 (N_49596,N_49034,N_49219);
nand U49597 (N_49597,N_49257,N_49140);
nor U49598 (N_49598,N_49283,N_49044);
or U49599 (N_49599,N_49318,N_49422);
nand U49600 (N_49600,N_49189,N_49358);
nor U49601 (N_49601,N_49008,N_49047);
xor U49602 (N_49602,N_49094,N_49383);
nand U49603 (N_49603,N_49032,N_49370);
or U49604 (N_49604,N_49456,N_49429);
nand U49605 (N_49605,N_49075,N_49275);
or U49606 (N_49606,N_49320,N_49021);
nor U49607 (N_49607,N_49466,N_49057);
and U49608 (N_49608,N_49029,N_49284);
and U49609 (N_49609,N_49347,N_49185);
nor U49610 (N_49610,N_49373,N_49489);
nor U49611 (N_49611,N_49431,N_49117);
or U49612 (N_49612,N_49310,N_49160);
or U49613 (N_49613,N_49111,N_49254);
or U49614 (N_49614,N_49216,N_49043);
xnor U49615 (N_49615,N_49113,N_49406);
or U49616 (N_49616,N_49480,N_49244);
nor U49617 (N_49617,N_49308,N_49136);
xnor U49618 (N_49618,N_49368,N_49106);
xnor U49619 (N_49619,N_49049,N_49393);
nor U49620 (N_49620,N_49196,N_49045);
and U49621 (N_49621,N_49262,N_49209);
nor U49622 (N_49622,N_49328,N_49166);
nor U49623 (N_49623,N_49208,N_49438);
or U49624 (N_49624,N_49437,N_49114);
or U49625 (N_49625,N_49156,N_49446);
nand U49626 (N_49626,N_49381,N_49390);
xor U49627 (N_49627,N_49281,N_49285);
or U49628 (N_49628,N_49260,N_49016);
or U49629 (N_49629,N_49343,N_49404);
nor U49630 (N_49630,N_49277,N_49388);
nand U49631 (N_49631,N_49478,N_49163);
xnor U49632 (N_49632,N_49375,N_49295);
xor U49633 (N_49633,N_49282,N_49141);
or U49634 (N_49634,N_49247,N_49417);
and U49635 (N_49635,N_49040,N_49139);
nor U49636 (N_49636,N_49314,N_49485);
and U49637 (N_49637,N_49441,N_49221);
xnor U49638 (N_49638,N_49401,N_49267);
nand U49639 (N_49639,N_49416,N_49082);
or U49640 (N_49640,N_49353,N_49190);
nor U49641 (N_49641,N_49475,N_49442);
nand U49642 (N_49642,N_49374,N_49088);
nand U49643 (N_49643,N_49074,N_49012);
and U49644 (N_49644,N_49334,N_49337);
nor U49645 (N_49645,N_49469,N_49092);
nor U49646 (N_49646,N_49324,N_49280);
and U49647 (N_49647,N_49372,N_49268);
nand U49648 (N_49648,N_49487,N_49412);
nand U49649 (N_49649,N_49144,N_49265);
nand U49650 (N_49650,N_49133,N_49499);
or U49651 (N_49651,N_49100,N_49365);
and U49652 (N_49652,N_49243,N_49494);
or U49653 (N_49653,N_49129,N_49425);
xnor U49654 (N_49654,N_49191,N_49164);
nor U49655 (N_49655,N_49115,N_49467);
or U49656 (N_49656,N_49200,N_49352);
nor U49657 (N_49657,N_49322,N_49248);
xnor U49658 (N_49658,N_49228,N_49240);
or U49659 (N_49659,N_49245,N_49174);
or U49660 (N_49660,N_49073,N_49359);
and U49661 (N_49661,N_49157,N_49421);
or U49662 (N_49662,N_49015,N_49479);
or U49663 (N_49663,N_49064,N_49173);
nor U49664 (N_49664,N_49217,N_49460);
and U49665 (N_49665,N_49385,N_49414);
or U49666 (N_49666,N_49279,N_49266);
and U49667 (N_49667,N_49218,N_49327);
xnor U49668 (N_49668,N_49413,N_49246);
nand U49669 (N_49669,N_49458,N_49222);
nor U49670 (N_49670,N_49433,N_49319);
nand U49671 (N_49671,N_49202,N_49002);
xnor U49672 (N_49672,N_49086,N_49238);
nand U49673 (N_49673,N_49317,N_49124);
nand U49674 (N_49674,N_49299,N_49303);
or U49675 (N_49675,N_49495,N_49443);
nor U49676 (N_49676,N_49145,N_49198);
nor U49677 (N_49677,N_49483,N_49063);
and U49678 (N_49678,N_49250,N_49230);
nor U49679 (N_49679,N_49220,N_49036);
xor U49680 (N_49680,N_49278,N_49461);
nor U49681 (N_49681,N_49065,N_49067);
and U49682 (N_49682,N_49225,N_49188);
xor U49683 (N_49683,N_49297,N_49004);
and U49684 (N_49684,N_49445,N_49022);
nor U49685 (N_49685,N_49452,N_49019);
and U49686 (N_49686,N_49078,N_49427);
or U49687 (N_49687,N_49186,N_49081);
xnor U49688 (N_49688,N_49213,N_49109);
nor U49689 (N_49689,N_49041,N_49439);
xor U49690 (N_49690,N_49382,N_49062);
nor U49691 (N_49691,N_49108,N_49335);
or U49692 (N_49692,N_49104,N_49463);
and U49693 (N_49693,N_49118,N_49192);
or U49694 (N_49694,N_49005,N_49492);
nor U49695 (N_49695,N_49107,N_49014);
or U49696 (N_49696,N_49096,N_49239);
xnor U49697 (N_49697,N_49403,N_49052);
or U49698 (N_49698,N_49123,N_49252);
nand U49699 (N_49699,N_49010,N_49341);
xnor U49700 (N_49700,N_49428,N_49472);
and U49701 (N_49701,N_49195,N_49362);
nand U49702 (N_49702,N_49007,N_49258);
nor U49703 (N_49703,N_49235,N_49307);
or U49704 (N_49704,N_49377,N_49102);
or U49705 (N_49705,N_49326,N_49451);
and U49706 (N_49706,N_49306,N_49360);
xnor U49707 (N_49707,N_49054,N_49027);
nand U49708 (N_49708,N_49305,N_49488);
nand U49709 (N_49709,N_49400,N_49152);
or U49710 (N_49710,N_49211,N_49474);
nand U49711 (N_49711,N_49309,N_49423);
or U49712 (N_49712,N_49020,N_49033);
or U49713 (N_49713,N_49294,N_49436);
or U49714 (N_49714,N_49391,N_49288);
nor U49715 (N_49715,N_49396,N_49087);
nor U49716 (N_49716,N_49454,N_49097);
nand U49717 (N_49717,N_49090,N_49290);
xnor U49718 (N_49718,N_49060,N_49126);
nand U49719 (N_49719,N_49384,N_49079);
or U49720 (N_49720,N_49138,N_49091);
and U49721 (N_49721,N_49471,N_49171);
nand U49722 (N_49722,N_49378,N_49071);
nor U49723 (N_49723,N_49269,N_49132);
nor U49724 (N_49724,N_49298,N_49392);
xnor U49725 (N_49725,N_49125,N_49394);
and U49726 (N_49726,N_49411,N_49286);
xor U49727 (N_49727,N_49098,N_49201);
nand U49728 (N_49728,N_49346,N_49482);
xor U49729 (N_49729,N_49037,N_49000);
and U49730 (N_49730,N_49493,N_49330);
nor U49731 (N_49731,N_49355,N_49313);
nor U49732 (N_49732,N_49476,N_49056);
and U49733 (N_49733,N_49249,N_49030);
nor U49734 (N_49734,N_49011,N_49223);
and U49735 (N_49735,N_49083,N_49261);
and U49736 (N_49736,N_49028,N_49367);
nor U49737 (N_49737,N_49435,N_49302);
nand U49738 (N_49738,N_49292,N_49440);
nor U49739 (N_49739,N_49410,N_49101);
nor U49740 (N_49740,N_49434,N_49366);
or U49741 (N_49741,N_49398,N_49069);
or U49742 (N_49742,N_49122,N_49003);
xor U49743 (N_49743,N_49496,N_49165);
nand U49744 (N_49744,N_49332,N_49321);
or U49745 (N_49745,N_49039,N_49376);
and U49746 (N_49746,N_49205,N_49363);
and U49747 (N_49747,N_49387,N_49457);
or U49748 (N_49748,N_49350,N_49255);
and U49749 (N_49749,N_49193,N_49059);
nor U49750 (N_49750,N_49298,N_49039);
xor U49751 (N_49751,N_49294,N_49194);
and U49752 (N_49752,N_49182,N_49168);
or U49753 (N_49753,N_49399,N_49487);
xor U49754 (N_49754,N_49143,N_49037);
xor U49755 (N_49755,N_49373,N_49007);
xnor U49756 (N_49756,N_49286,N_49479);
or U49757 (N_49757,N_49034,N_49363);
nor U49758 (N_49758,N_49310,N_49120);
or U49759 (N_49759,N_49150,N_49479);
and U49760 (N_49760,N_49294,N_49316);
nand U49761 (N_49761,N_49393,N_49164);
nor U49762 (N_49762,N_49362,N_49160);
or U49763 (N_49763,N_49115,N_49419);
or U49764 (N_49764,N_49383,N_49043);
nor U49765 (N_49765,N_49383,N_49078);
nor U49766 (N_49766,N_49131,N_49265);
and U49767 (N_49767,N_49398,N_49050);
xnor U49768 (N_49768,N_49249,N_49492);
or U49769 (N_49769,N_49187,N_49412);
nor U49770 (N_49770,N_49302,N_49056);
nand U49771 (N_49771,N_49104,N_49346);
and U49772 (N_49772,N_49443,N_49157);
xor U49773 (N_49773,N_49366,N_49097);
and U49774 (N_49774,N_49053,N_49080);
or U49775 (N_49775,N_49278,N_49096);
and U49776 (N_49776,N_49391,N_49224);
nand U49777 (N_49777,N_49354,N_49179);
xnor U49778 (N_49778,N_49256,N_49174);
nand U49779 (N_49779,N_49083,N_49392);
nor U49780 (N_49780,N_49101,N_49224);
xor U49781 (N_49781,N_49181,N_49330);
or U49782 (N_49782,N_49164,N_49491);
nand U49783 (N_49783,N_49489,N_49302);
xor U49784 (N_49784,N_49074,N_49232);
xnor U49785 (N_49785,N_49182,N_49059);
and U49786 (N_49786,N_49365,N_49387);
or U49787 (N_49787,N_49341,N_49123);
or U49788 (N_49788,N_49462,N_49138);
nand U49789 (N_49789,N_49290,N_49313);
nand U49790 (N_49790,N_49337,N_49146);
nand U49791 (N_49791,N_49036,N_49289);
xor U49792 (N_49792,N_49263,N_49324);
xor U49793 (N_49793,N_49264,N_49316);
or U49794 (N_49794,N_49176,N_49051);
nand U49795 (N_49795,N_49429,N_49374);
nor U49796 (N_49796,N_49383,N_49023);
xnor U49797 (N_49797,N_49276,N_49034);
nor U49798 (N_49798,N_49089,N_49371);
xor U49799 (N_49799,N_49369,N_49044);
nand U49800 (N_49800,N_49325,N_49393);
or U49801 (N_49801,N_49056,N_49452);
and U49802 (N_49802,N_49332,N_49249);
xor U49803 (N_49803,N_49040,N_49049);
or U49804 (N_49804,N_49282,N_49127);
and U49805 (N_49805,N_49218,N_49448);
nand U49806 (N_49806,N_49264,N_49233);
nor U49807 (N_49807,N_49164,N_49416);
nand U49808 (N_49808,N_49356,N_49437);
and U49809 (N_49809,N_49449,N_49041);
or U49810 (N_49810,N_49363,N_49065);
nand U49811 (N_49811,N_49225,N_49428);
nand U49812 (N_49812,N_49108,N_49410);
and U49813 (N_49813,N_49485,N_49428);
and U49814 (N_49814,N_49166,N_49039);
nand U49815 (N_49815,N_49278,N_49397);
nor U49816 (N_49816,N_49177,N_49006);
nand U49817 (N_49817,N_49425,N_49022);
xnor U49818 (N_49818,N_49186,N_49267);
xnor U49819 (N_49819,N_49353,N_49010);
nor U49820 (N_49820,N_49227,N_49234);
and U49821 (N_49821,N_49222,N_49406);
nor U49822 (N_49822,N_49333,N_49467);
nor U49823 (N_49823,N_49415,N_49032);
nand U49824 (N_49824,N_49390,N_49188);
xnor U49825 (N_49825,N_49214,N_49026);
or U49826 (N_49826,N_49428,N_49245);
xnor U49827 (N_49827,N_49260,N_49436);
nor U49828 (N_49828,N_49126,N_49210);
nor U49829 (N_49829,N_49334,N_49353);
nor U49830 (N_49830,N_49234,N_49330);
xnor U49831 (N_49831,N_49090,N_49432);
nand U49832 (N_49832,N_49496,N_49199);
or U49833 (N_49833,N_49134,N_49062);
or U49834 (N_49834,N_49288,N_49471);
and U49835 (N_49835,N_49334,N_49242);
nor U49836 (N_49836,N_49267,N_49322);
xor U49837 (N_49837,N_49202,N_49020);
nand U49838 (N_49838,N_49175,N_49304);
or U49839 (N_49839,N_49452,N_49334);
nor U49840 (N_49840,N_49209,N_49486);
nand U49841 (N_49841,N_49491,N_49239);
xor U49842 (N_49842,N_49236,N_49182);
xnor U49843 (N_49843,N_49138,N_49269);
xor U49844 (N_49844,N_49059,N_49048);
nor U49845 (N_49845,N_49007,N_49093);
nor U49846 (N_49846,N_49270,N_49231);
and U49847 (N_49847,N_49081,N_49000);
nor U49848 (N_49848,N_49011,N_49383);
xor U49849 (N_49849,N_49100,N_49257);
nand U49850 (N_49850,N_49330,N_49148);
or U49851 (N_49851,N_49371,N_49174);
xor U49852 (N_49852,N_49166,N_49413);
nand U49853 (N_49853,N_49446,N_49116);
nand U49854 (N_49854,N_49285,N_49216);
xnor U49855 (N_49855,N_49280,N_49033);
nor U49856 (N_49856,N_49354,N_49095);
and U49857 (N_49857,N_49370,N_49179);
or U49858 (N_49858,N_49282,N_49289);
xnor U49859 (N_49859,N_49068,N_49264);
xnor U49860 (N_49860,N_49174,N_49184);
nor U49861 (N_49861,N_49402,N_49480);
xor U49862 (N_49862,N_49438,N_49369);
or U49863 (N_49863,N_49227,N_49435);
xor U49864 (N_49864,N_49471,N_49486);
nor U49865 (N_49865,N_49270,N_49010);
nor U49866 (N_49866,N_49063,N_49376);
or U49867 (N_49867,N_49460,N_49457);
and U49868 (N_49868,N_49168,N_49119);
xor U49869 (N_49869,N_49464,N_49414);
xnor U49870 (N_49870,N_49104,N_49254);
nand U49871 (N_49871,N_49260,N_49316);
and U49872 (N_49872,N_49410,N_49384);
or U49873 (N_49873,N_49197,N_49261);
nor U49874 (N_49874,N_49368,N_49427);
nand U49875 (N_49875,N_49469,N_49497);
or U49876 (N_49876,N_49184,N_49006);
and U49877 (N_49877,N_49488,N_49044);
or U49878 (N_49878,N_49396,N_49033);
nor U49879 (N_49879,N_49155,N_49359);
or U49880 (N_49880,N_49406,N_49340);
nand U49881 (N_49881,N_49401,N_49075);
xnor U49882 (N_49882,N_49139,N_49486);
nand U49883 (N_49883,N_49194,N_49099);
nor U49884 (N_49884,N_49194,N_49002);
and U49885 (N_49885,N_49457,N_49183);
or U49886 (N_49886,N_49431,N_49182);
or U49887 (N_49887,N_49276,N_49073);
nor U49888 (N_49888,N_49190,N_49286);
and U49889 (N_49889,N_49203,N_49188);
or U49890 (N_49890,N_49014,N_49099);
or U49891 (N_49891,N_49461,N_49186);
xor U49892 (N_49892,N_49150,N_49252);
nor U49893 (N_49893,N_49431,N_49447);
or U49894 (N_49894,N_49471,N_49106);
and U49895 (N_49895,N_49369,N_49082);
nand U49896 (N_49896,N_49004,N_49355);
and U49897 (N_49897,N_49364,N_49060);
and U49898 (N_49898,N_49395,N_49045);
nand U49899 (N_49899,N_49435,N_49487);
or U49900 (N_49900,N_49059,N_49105);
nor U49901 (N_49901,N_49359,N_49153);
nor U49902 (N_49902,N_49164,N_49215);
nand U49903 (N_49903,N_49144,N_49140);
nand U49904 (N_49904,N_49094,N_49103);
nor U49905 (N_49905,N_49430,N_49084);
nor U49906 (N_49906,N_49051,N_49120);
or U49907 (N_49907,N_49014,N_49197);
xnor U49908 (N_49908,N_49474,N_49468);
xnor U49909 (N_49909,N_49016,N_49226);
or U49910 (N_49910,N_49002,N_49464);
and U49911 (N_49911,N_49496,N_49344);
nand U49912 (N_49912,N_49484,N_49282);
nor U49913 (N_49913,N_49169,N_49395);
nand U49914 (N_49914,N_49107,N_49177);
xnor U49915 (N_49915,N_49135,N_49094);
or U49916 (N_49916,N_49047,N_49216);
or U49917 (N_49917,N_49304,N_49319);
and U49918 (N_49918,N_49179,N_49009);
or U49919 (N_49919,N_49435,N_49238);
or U49920 (N_49920,N_49494,N_49177);
nor U49921 (N_49921,N_49494,N_49472);
and U49922 (N_49922,N_49306,N_49168);
and U49923 (N_49923,N_49344,N_49414);
nor U49924 (N_49924,N_49199,N_49015);
nor U49925 (N_49925,N_49125,N_49477);
or U49926 (N_49926,N_49172,N_49170);
and U49927 (N_49927,N_49487,N_49427);
xnor U49928 (N_49928,N_49389,N_49107);
nand U49929 (N_49929,N_49411,N_49049);
and U49930 (N_49930,N_49497,N_49144);
nand U49931 (N_49931,N_49427,N_49061);
or U49932 (N_49932,N_49444,N_49481);
or U49933 (N_49933,N_49269,N_49413);
and U49934 (N_49934,N_49174,N_49140);
nor U49935 (N_49935,N_49109,N_49491);
xor U49936 (N_49936,N_49232,N_49221);
nor U49937 (N_49937,N_49191,N_49440);
or U49938 (N_49938,N_49128,N_49278);
and U49939 (N_49939,N_49448,N_49077);
xor U49940 (N_49940,N_49250,N_49001);
and U49941 (N_49941,N_49413,N_49455);
xor U49942 (N_49942,N_49493,N_49005);
and U49943 (N_49943,N_49106,N_49116);
and U49944 (N_49944,N_49175,N_49142);
or U49945 (N_49945,N_49470,N_49076);
nor U49946 (N_49946,N_49312,N_49427);
xnor U49947 (N_49947,N_49379,N_49091);
or U49948 (N_49948,N_49062,N_49141);
and U49949 (N_49949,N_49283,N_49085);
nand U49950 (N_49950,N_49430,N_49391);
nor U49951 (N_49951,N_49220,N_49471);
nand U49952 (N_49952,N_49013,N_49361);
xor U49953 (N_49953,N_49309,N_49398);
and U49954 (N_49954,N_49189,N_49424);
nor U49955 (N_49955,N_49093,N_49003);
nand U49956 (N_49956,N_49048,N_49239);
nor U49957 (N_49957,N_49256,N_49288);
nand U49958 (N_49958,N_49242,N_49233);
and U49959 (N_49959,N_49342,N_49347);
nor U49960 (N_49960,N_49482,N_49182);
nor U49961 (N_49961,N_49185,N_49392);
nor U49962 (N_49962,N_49250,N_49363);
xnor U49963 (N_49963,N_49219,N_49073);
or U49964 (N_49964,N_49070,N_49002);
and U49965 (N_49965,N_49292,N_49006);
nor U49966 (N_49966,N_49271,N_49098);
xor U49967 (N_49967,N_49135,N_49384);
nor U49968 (N_49968,N_49399,N_49045);
xnor U49969 (N_49969,N_49322,N_49438);
and U49970 (N_49970,N_49393,N_49117);
nor U49971 (N_49971,N_49344,N_49010);
nand U49972 (N_49972,N_49027,N_49424);
and U49973 (N_49973,N_49033,N_49476);
nor U49974 (N_49974,N_49106,N_49040);
and U49975 (N_49975,N_49018,N_49488);
nand U49976 (N_49976,N_49102,N_49042);
nand U49977 (N_49977,N_49254,N_49385);
nor U49978 (N_49978,N_49008,N_49095);
nand U49979 (N_49979,N_49230,N_49196);
nand U49980 (N_49980,N_49278,N_49160);
and U49981 (N_49981,N_49054,N_49334);
nor U49982 (N_49982,N_49123,N_49178);
nand U49983 (N_49983,N_49321,N_49367);
and U49984 (N_49984,N_49352,N_49366);
or U49985 (N_49985,N_49060,N_49189);
nand U49986 (N_49986,N_49497,N_49388);
xor U49987 (N_49987,N_49383,N_49385);
or U49988 (N_49988,N_49343,N_49437);
nand U49989 (N_49989,N_49222,N_49015);
or U49990 (N_49990,N_49434,N_49169);
nand U49991 (N_49991,N_49033,N_49032);
xnor U49992 (N_49992,N_49162,N_49404);
xnor U49993 (N_49993,N_49495,N_49146);
nand U49994 (N_49994,N_49493,N_49422);
xnor U49995 (N_49995,N_49279,N_49223);
or U49996 (N_49996,N_49058,N_49236);
or U49997 (N_49997,N_49194,N_49422);
nand U49998 (N_49998,N_49417,N_49270);
and U49999 (N_49999,N_49168,N_49010);
xor UO_0 (O_0,N_49812,N_49751);
xor UO_1 (O_1,N_49623,N_49570);
or UO_2 (O_2,N_49767,N_49647);
nor UO_3 (O_3,N_49771,N_49849);
nor UO_4 (O_4,N_49993,N_49973);
nor UO_5 (O_5,N_49723,N_49853);
nor UO_6 (O_6,N_49589,N_49824);
nand UO_7 (O_7,N_49947,N_49813);
nor UO_8 (O_8,N_49980,N_49713);
and UO_9 (O_9,N_49890,N_49537);
nor UO_10 (O_10,N_49925,N_49869);
nor UO_11 (O_11,N_49660,N_49881);
and UO_12 (O_12,N_49631,N_49913);
nor UO_13 (O_13,N_49833,N_49880);
xnor UO_14 (O_14,N_49856,N_49875);
xnor UO_15 (O_15,N_49750,N_49523);
xor UO_16 (O_16,N_49800,N_49991);
or UO_17 (O_17,N_49722,N_49807);
xor UO_18 (O_18,N_49546,N_49682);
nand UO_19 (O_19,N_49953,N_49950);
or UO_20 (O_20,N_49539,N_49970);
or UO_21 (O_21,N_49607,N_49939);
nor UO_22 (O_22,N_49815,N_49638);
nor UO_23 (O_23,N_49739,N_49936);
nand UO_24 (O_24,N_49691,N_49714);
nor UO_25 (O_25,N_49898,N_49787);
nand UO_26 (O_26,N_49779,N_49557);
xnor UO_27 (O_27,N_49586,N_49692);
nor UO_28 (O_28,N_49903,N_49593);
nor UO_29 (O_29,N_49923,N_49552);
and UO_30 (O_30,N_49958,N_49838);
nand UO_31 (O_31,N_49511,N_49761);
and UO_32 (O_32,N_49500,N_49572);
nor UO_33 (O_33,N_49885,N_49995);
and UO_34 (O_34,N_49636,N_49677);
and UO_35 (O_35,N_49749,N_49984);
nand UO_36 (O_36,N_49628,N_49707);
or UO_37 (O_37,N_49542,N_49769);
and UO_38 (O_38,N_49520,N_49826);
and UO_39 (O_39,N_49782,N_49582);
xor UO_40 (O_40,N_49770,N_49509);
nor UO_41 (O_41,N_49610,N_49775);
or UO_42 (O_42,N_49961,N_49621);
and UO_43 (O_43,N_49627,N_49652);
nor UO_44 (O_44,N_49503,N_49730);
and UO_45 (O_45,N_49906,N_49781);
xnor UO_46 (O_46,N_49559,N_49614);
xor UO_47 (O_47,N_49711,N_49697);
and UO_48 (O_48,N_49565,N_49907);
nand UO_49 (O_49,N_49835,N_49651);
nand UO_50 (O_50,N_49954,N_49522);
and UO_51 (O_51,N_49596,N_49884);
nor UO_52 (O_52,N_49555,N_49857);
nand UO_53 (O_53,N_49791,N_49603);
or UO_54 (O_54,N_49989,N_49892);
nor UO_55 (O_55,N_49780,N_49528);
or UO_56 (O_56,N_49602,N_49673);
and UO_57 (O_57,N_49599,N_49635);
xnor UO_58 (O_58,N_49764,N_49914);
and UO_59 (O_59,N_49549,N_49744);
xnor UO_60 (O_60,N_49731,N_49922);
or UO_61 (O_61,N_49540,N_49967);
nand UO_62 (O_62,N_49785,N_49883);
xnor UO_63 (O_63,N_49959,N_49616);
xnor UO_64 (O_64,N_49832,N_49578);
nor UO_65 (O_65,N_49855,N_49605);
xor UO_66 (O_66,N_49741,N_49579);
xnor UO_67 (O_67,N_49728,N_49551);
or UO_68 (O_68,N_49902,N_49861);
or UO_69 (O_69,N_49620,N_49844);
nand UO_70 (O_70,N_49850,N_49740);
nor UO_71 (O_71,N_49910,N_49569);
and UO_72 (O_72,N_49726,N_49684);
nand UO_73 (O_73,N_49932,N_49762);
and UO_74 (O_74,N_49505,N_49686);
nor UO_75 (O_75,N_49705,N_49930);
or UO_76 (O_76,N_49878,N_49734);
nor UO_77 (O_77,N_49580,N_49618);
nand UO_78 (O_78,N_49680,N_49533);
nand UO_79 (O_79,N_49574,N_49576);
xor UO_80 (O_80,N_49735,N_49654);
xor UO_81 (O_81,N_49633,N_49985);
xor UO_82 (O_82,N_49604,N_49920);
or UO_83 (O_83,N_49790,N_49649);
xor UO_84 (O_84,N_49653,N_49891);
and UO_85 (O_85,N_49667,N_49597);
or UO_86 (O_86,N_49753,N_49561);
xor UO_87 (O_87,N_49564,N_49554);
xnor UO_88 (O_88,N_49748,N_49567);
or UO_89 (O_89,N_49823,N_49577);
and UO_90 (O_90,N_49590,N_49957);
or UO_91 (O_91,N_49931,N_49994);
or UO_92 (O_92,N_49525,N_49810);
nor UO_93 (O_93,N_49909,N_49532);
nand UO_94 (O_94,N_49611,N_49942);
nor UO_95 (O_95,N_49512,N_49772);
or UO_96 (O_96,N_49831,N_49752);
nand UO_97 (O_97,N_49658,N_49632);
xor UO_98 (O_98,N_49986,N_49797);
and UO_99 (O_99,N_49513,N_49688);
xor UO_100 (O_100,N_49821,N_49687);
nor UO_101 (O_101,N_49699,N_49927);
and UO_102 (O_102,N_49661,N_49981);
xnor UO_103 (O_103,N_49516,N_49895);
xnor UO_104 (O_104,N_49746,N_49659);
nand UO_105 (O_105,N_49608,N_49613);
or UO_106 (O_106,N_49836,N_49738);
nand UO_107 (O_107,N_49745,N_49820);
or UO_108 (O_108,N_49556,N_49594);
and UO_109 (O_109,N_49971,N_49786);
and UO_110 (O_110,N_49837,N_49657);
and UO_111 (O_111,N_49872,N_49563);
xnor UO_112 (O_112,N_49601,N_49612);
xnor UO_113 (O_113,N_49547,N_49758);
xnor UO_114 (O_114,N_49882,N_49972);
and UO_115 (O_115,N_49889,N_49901);
or UO_116 (O_116,N_49646,N_49867);
or UO_117 (O_117,N_49982,N_49763);
nand UO_118 (O_118,N_49733,N_49587);
nor UO_119 (O_119,N_49575,N_49640);
nor UO_120 (O_120,N_49672,N_49679);
nand UO_121 (O_121,N_49917,N_49894);
nand UO_122 (O_122,N_49664,N_49962);
nor UO_123 (O_123,N_49940,N_49701);
nor UO_124 (O_124,N_49689,N_49999);
nor UO_125 (O_125,N_49765,N_49521);
nand UO_126 (O_126,N_49581,N_49648);
and UO_127 (O_127,N_49504,N_49788);
or UO_128 (O_128,N_49834,N_49553);
xnor UO_129 (O_129,N_49963,N_49754);
nor UO_130 (O_130,N_49719,N_49757);
xor UO_131 (O_131,N_49600,N_49543);
or UO_132 (O_132,N_49768,N_49825);
xnor UO_133 (O_133,N_49566,N_49798);
and UO_134 (O_134,N_49702,N_49774);
and UO_135 (O_135,N_49560,N_49721);
nand UO_136 (O_136,N_49703,N_49756);
and UO_137 (O_137,N_49839,N_49650);
nand UO_138 (O_138,N_49584,N_49960);
and UO_139 (O_139,N_49615,N_49924);
xor UO_140 (O_140,N_49865,N_49830);
nor UO_141 (O_141,N_49715,N_49915);
or UO_142 (O_142,N_49671,N_49926);
nand UO_143 (O_143,N_49736,N_49822);
and UO_144 (O_144,N_49755,N_49796);
or UO_145 (O_145,N_49643,N_49676);
xnor UO_146 (O_146,N_49956,N_49864);
and UO_147 (O_147,N_49515,N_49716);
or UO_148 (O_148,N_49571,N_49949);
or UO_149 (O_149,N_49585,N_49747);
nor UO_150 (O_150,N_49545,N_49617);
nor UO_151 (O_151,N_49933,N_49847);
nand UO_152 (O_152,N_49665,N_49783);
nand UO_153 (O_153,N_49929,N_49866);
xor UO_154 (O_154,N_49870,N_49535);
and UO_155 (O_155,N_49904,N_49841);
or UO_156 (O_156,N_49606,N_49698);
xor UO_157 (O_157,N_49987,N_49979);
xnor UO_158 (O_158,N_49655,N_49519);
xor UO_159 (O_159,N_49639,N_49899);
xor UO_160 (O_160,N_49696,N_49819);
xor UO_161 (O_161,N_49937,N_49911);
xnor UO_162 (O_162,N_49704,N_49921);
nand UO_163 (O_163,N_49801,N_49946);
xor UO_164 (O_164,N_49694,N_49886);
or UO_165 (O_165,N_49951,N_49879);
nor UO_166 (O_166,N_49792,N_49729);
nand UO_167 (O_167,N_49527,N_49966);
nand UO_168 (O_168,N_49529,N_49806);
or UO_169 (O_169,N_49641,N_49845);
xor UO_170 (O_170,N_49541,N_49952);
xnor UO_171 (O_171,N_49843,N_49789);
xnor UO_172 (O_172,N_49842,N_49663);
nand UO_173 (O_173,N_49544,N_49988);
xnor UO_174 (O_174,N_49724,N_49625);
nand UO_175 (O_175,N_49595,N_49955);
and UO_176 (O_176,N_49969,N_49700);
nand UO_177 (O_177,N_49619,N_49773);
nand UO_178 (O_178,N_49863,N_49662);
and UO_179 (O_179,N_49854,N_49592);
xor UO_180 (O_180,N_49510,N_49965);
nor UO_181 (O_181,N_49828,N_49524);
or UO_182 (O_182,N_49997,N_49905);
and UO_183 (O_183,N_49802,N_49766);
nor UO_184 (O_184,N_49637,N_49919);
nor UO_185 (O_185,N_49945,N_49888);
xor UO_186 (O_186,N_49710,N_49727);
and UO_187 (O_187,N_49868,N_49859);
xor UO_188 (O_188,N_49873,N_49976);
nor UO_189 (O_189,N_49678,N_49674);
nand UO_190 (O_190,N_49693,N_49778);
nor UO_191 (O_191,N_49514,N_49508);
or UO_192 (O_192,N_49871,N_49626);
nand UO_193 (O_193,N_49759,N_49794);
nand UO_194 (O_194,N_49670,N_49829);
xnor UO_195 (O_195,N_49977,N_49912);
nand UO_196 (O_196,N_49695,N_49558);
and UO_197 (O_197,N_49816,N_49928);
or UO_198 (O_198,N_49846,N_49675);
nand UO_199 (O_199,N_49811,N_49501);
or UO_200 (O_200,N_49803,N_49874);
and UO_201 (O_201,N_49732,N_49896);
or UO_202 (O_202,N_49996,N_49918);
and UO_203 (O_203,N_49645,N_49990);
nor UO_204 (O_204,N_49609,N_49848);
xnor UO_205 (O_205,N_49550,N_49548);
nor UO_206 (O_206,N_49760,N_49799);
or UO_207 (O_207,N_49506,N_49502);
or UO_208 (O_208,N_49983,N_49944);
and UO_209 (O_209,N_49517,N_49858);
or UO_210 (O_210,N_49562,N_49588);
xor UO_211 (O_211,N_49777,N_49809);
xor UO_212 (O_212,N_49573,N_49742);
or UO_213 (O_213,N_49784,N_49818);
nand UO_214 (O_214,N_49876,N_49743);
or UO_215 (O_215,N_49887,N_49893);
nor UO_216 (O_216,N_49793,N_49656);
and UO_217 (O_217,N_49943,N_49591);
nor UO_218 (O_218,N_49583,N_49974);
or UO_219 (O_219,N_49622,N_49776);
xnor UO_220 (O_220,N_49534,N_49598);
and UO_221 (O_221,N_49968,N_49814);
nor UO_222 (O_222,N_49934,N_49998);
and UO_223 (O_223,N_49978,N_49568);
or UO_224 (O_224,N_49805,N_49538);
nor UO_225 (O_225,N_49804,N_49935);
xnor UO_226 (O_226,N_49908,N_49536);
xnor UO_227 (O_227,N_49827,N_49852);
nor UO_228 (O_228,N_49795,N_49668);
or UO_229 (O_229,N_49948,N_49629);
or UO_230 (O_230,N_49530,N_49630);
or UO_231 (O_231,N_49685,N_49817);
and UO_232 (O_232,N_49642,N_49860);
nand UO_233 (O_233,N_49964,N_49531);
nand UO_234 (O_234,N_49900,N_49624);
and UO_235 (O_235,N_49526,N_49897);
nor UO_236 (O_236,N_49706,N_49709);
xor UO_237 (O_237,N_49941,N_49720);
and UO_238 (O_238,N_49808,N_49862);
or UO_239 (O_239,N_49683,N_49518);
nor UO_240 (O_240,N_49938,N_49690);
nor UO_241 (O_241,N_49737,N_49669);
xor UO_242 (O_242,N_49717,N_49725);
and UO_243 (O_243,N_49718,N_49851);
nand UO_244 (O_244,N_49708,N_49975);
or UO_245 (O_245,N_49681,N_49634);
and UO_246 (O_246,N_49507,N_49916);
nand UO_247 (O_247,N_49992,N_49877);
nand UO_248 (O_248,N_49712,N_49666);
and UO_249 (O_249,N_49840,N_49644);
xor UO_250 (O_250,N_49763,N_49812);
nand UO_251 (O_251,N_49807,N_49679);
nor UO_252 (O_252,N_49690,N_49557);
and UO_253 (O_253,N_49614,N_49844);
nand UO_254 (O_254,N_49710,N_49598);
nor UO_255 (O_255,N_49985,N_49747);
nor UO_256 (O_256,N_49534,N_49542);
xor UO_257 (O_257,N_49518,N_49521);
and UO_258 (O_258,N_49723,N_49922);
or UO_259 (O_259,N_49890,N_49609);
and UO_260 (O_260,N_49832,N_49576);
nand UO_261 (O_261,N_49684,N_49560);
nor UO_262 (O_262,N_49926,N_49733);
or UO_263 (O_263,N_49806,N_49837);
and UO_264 (O_264,N_49860,N_49627);
and UO_265 (O_265,N_49639,N_49940);
nor UO_266 (O_266,N_49635,N_49665);
xnor UO_267 (O_267,N_49672,N_49774);
nand UO_268 (O_268,N_49671,N_49917);
nand UO_269 (O_269,N_49754,N_49767);
nand UO_270 (O_270,N_49723,N_49863);
and UO_271 (O_271,N_49781,N_49827);
nor UO_272 (O_272,N_49574,N_49854);
or UO_273 (O_273,N_49612,N_49775);
or UO_274 (O_274,N_49600,N_49550);
xnor UO_275 (O_275,N_49960,N_49885);
nand UO_276 (O_276,N_49764,N_49619);
nand UO_277 (O_277,N_49594,N_49571);
nand UO_278 (O_278,N_49546,N_49908);
nand UO_279 (O_279,N_49606,N_49638);
nor UO_280 (O_280,N_49757,N_49570);
xnor UO_281 (O_281,N_49965,N_49846);
and UO_282 (O_282,N_49528,N_49565);
nor UO_283 (O_283,N_49810,N_49985);
nand UO_284 (O_284,N_49682,N_49551);
xor UO_285 (O_285,N_49788,N_49928);
nand UO_286 (O_286,N_49696,N_49615);
nand UO_287 (O_287,N_49755,N_49624);
nand UO_288 (O_288,N_49989,N_49965);
nor UO_289 (O_289,N_49568,N_49517);
or UO_290 (O_290,N_49504,N_49758);
nand UO_291 (O_291,N_49967,N_49858);
xor UO_292 (O_292,N_49841,N_49506);
nand UO_293 (O_293,N_49547,N_49596);
and UO_294 (O_294,N_49750,N_49926);
and UO_295 (O_295,N_49525,N_49897);
nand UO_296 (O_296,N_49822,N_49876);
and UO_297 (O_297,N_49742,N_49880);
xor UO_298 (O_298,N_49773,N_49801);
or UO_299 (O_299,N_49811,N_49671);
nand UO_300 (O_300,N_49973,N_49841);
xor UO_301 (O_301,N_49825,N_49598);
or UO_302 (O_302,N_49996,N_49795);
or UO_303 (O_303,N_49951,N_49582);
xor UO_304 (O_304,N_49793,N_49600);
nor UO_305 (O_305,N_49957,N_49798);
and UO_306 (O_306,N_49648,N_49835);
nand UO_307 (O_307,N_49731,N_49504);
or UO_308 (O_308,N_49639,N_49892);
nor UO_309 (O_309,N_49950,N_49765);
nor UO_310 (O_310,N_49970,N_49999);
nor UO_311 (O_311,N_49502,N_49512);
nand UO_312 (O_312,N_49824,N_49793);
xnor UO_313 (O_313,N_49639,N_49686);
and UO_314 (O_314,N_49940,N_49925);
nand UO_315 (O_315,N_49844,N_49885);
and UO_316 (O_316,N_49675,N_49823);
and UO_317 (O_317,N_49701,N_49602);
nor UO_318 (O_318,N_49917,N_49851);
or UO_319 (O_319,N_49823,N_49749);
xor UO_320 (O_320,N_49550,N_49603);
or UO_321 (O_321,N_49915,N_49916);
xor UO_322 (O_322,N_49693,N_49797);
or UO_323 (O_323,N_49946,N_49653);
or UO_324 (O_324,N_49866,N_49726);
and UO_325 (O_325,N_49993,N_49524);
and UO_326 (O_326,N_49804,N_49533);
nand UO_327 (O_327,N_49977,N_49635);
nor UO_328 (O_328,N_49755,N_49989);
nand UO_329 (O_329,N_49712,N_49885);
or UO_330 (O_330,N_49570,N_49617);
nand UO_331 (O_331,N_49869,N_49668);
xor UO_332 (O_332,N_49679,N_49936);
or UO_333 (O_333,N_49616,N_49668);
nand UO_334 (O_334,N_49925,N_49666);
or UO_335 (O_335,N_49825,N_49701);
xor UO_336 (O_336,N_49809,N_49882);
and UO_337 (O_337,N_49731,N_49954);
nor UO_338 (O_338,N_49577,N_49749);
xor UO_339 (O_339,N_49589,N_49573);
and UO_340 (O_340,N_49714,N_49992);
and UO_341 (O_341,N_49933,N_49968);
xnor UO_342 (O_342,N_49714,N_49998);
nor UO_343 (O_343,N_49665,N_49562);
nor UO_344 (O_344,N_49934,N_49560);
xor UO_345 (O_345,N_49882,N_49790);
or UO_346 (O_346,N_49605,N_49829);
nor UO_347 (O_347,N_49691,N_49834);
or UO_348 (O_348,N_49844,N_49549);
xnor UO_349 (O_349,N_49511,N_49500);
or UO_350 (O_350,N_49714,N_49967);
nand UO_351 (O_351,N_49633,N_49565);
xor UO_352 (O_352,N_49879,N_49969);
and UO_353 (O_353,N_49838,N_49548);
and UO_354 (O_354,N_49833,N_49961);
nor UO_355 (O_355,N_49791,N_49771);
and UO_356 (O_356,N_49756,N_49878);
or UO_357 (O_357,N_49528,N_49890);
xnor UO_358 (O_358,N_49826,N_49525);
nor UO_359 (O_359,N_49689,N_49716);
or UO_360 (O_360,N_49770,N_49859);
nor UO_361 (O_361,N_49744,N_49890);
or UO_362 (O_362,N_49644,N_49969);
and UO_363 (O_363,N_49964,N_49949);
nand UO_364 (O_364,N_49964,N_49846);
and UO_365 (O_365,N_49730,N_49530);
nor UO_366 (O_366,N_49714,N_49552);
nor UO_367 (O_367,N_49774,N_49658);
or UO_368 (O_368,N_49798,N_49972);
nand UO_369 (O_369,N_49637,N_49652);
or UO_370 (O_370,N_49590,N_49827);
and UO_371 (O_371,N_49863,N_49932);
and UO_372 (O_372,N_49626,N_49816);
nand UO_373 (O_373,N_49586,N_49659);
xor UO_374 (O_374,N_49532,N_49562);
nand UO_375 (O_375,N_49935,N_49584);
or UO_376 (O_376,N_49749,N_49999);
and UO_377 (O_377,N_49670,N_49822);
nand UO_378 (O_378,N_49665,N_49877);
nor UO_379 (O_379,N_49700,N_49778);
nor UO_380 (O_380,N_49821,N_49671);
and UO_381 (O_381,N_49758,N_49950);
nor UO_382 (O_382,N_49502,N_49830);
or UO_383 (O_383,N_49920,N_49607);
nand UO_384 (O_384,N_49571,N_49604);
and UO_385 (O_385,N_49851,N_49550);
nor UO_386 (O_386,N_49793,N_49972);
nand UO_387 (O_387,N_49836,N_49892);
or UO_388 (O_388,N_49692,N_49743);
and UO_389 (O_389,N_49634,N_49761);
xnor UO_390 (O_390,N_49999,N_49516);
xor UO_391 (O_391,N_49607,N_49958);
and UO_392 (O_392,N_49988,N_49658);
nand UO_393 (O_393,N_49812,N_49504);
nand UO_394 (O_394,N_49897,N_49687);
nor UO_395 (O_395,N_49704,N_49619);
xnor UO_396 (O_396,N_49837,N_49808);
and UO_397 (O_397,N_49537,N_49855);
xor UO_398 (O_398,N_49554,N_49619);
xor UO_399 (O_399,N_49649,N_49657);
or UO_400 (O_400,N_49522,N_49738);
nand UO_401 (O_401,N_49729,N_49744);
and UO_402 (O_402,N_49501,N_49712);
nand UO_403 (O_403,N_49866,N_49903);
xnor UO_404 (O_404,N_49586,N_49754);
xor UO_405 (O_405,N_49694,N_49797);
or UO_406 (O_406,N_49542,N_49686);
xor UO_407 (O_407,N_49988,N_49690);
nand UO_408 (O_408,N_49737,N_49552);
xnor UO_409 (O_409,N_49780,N_49588);
xor UO_410 (O_410,N_49806,N_49753);
xnor UO_411 (O_411,N_49886,N_49957);
and UO_412 (O_412,N_49968,N_49608);
and UO_413 (O_413,N_49742,N_49777);
and UO_414 (O_414,N_49617,N_49590);
or UO_415 (O_415,N_49850,N_49545);
or UO_416 (O_416,N_49962,N_49509);
xnor UO_417 (O_417,N_49570,N_49949);
or UO_418 (O_418,N_49912,N_49541);
nor UO_419 (O_419,N_49999,N_49659);
nand UO_420 (O_420,N_49687,N_49944);
or UO_421 (O_421,N_49822,N_49584);
or UO_422 (O_422,N_49652,N_49969);
or UO_423 (O_423,N_49596,N_49562);
xnor UO_424 (O_424,N_49539,N_49923);
xor UO_425 (O_425,N_49827,N_49870);
xnor UO_426 (O_426,N_49729,N_49609);
nand UO_427 (O_427,N_49888,N_49533);
xnor UO_428 (O_428,N_49990,N_49889);
nand UO_429 (O_429,N_49504,N_49582);
or UO_430 (O_430,N_49611,N_49632);
nand UO_431 (O_431,N_49843,N_49531);
and UO_432 (O_432,N_49847,N_49921);
nand UO_433 (O_433,N_49775,N_49506);
nor UO_434 (O_434,N_49649,N_49652);
nor UO_435 (O_435,N_49998,N_49902);
nand UO_436 (O_436,N_49521,N_49756);
nand UO_437 (O_437,N_49721,N_49750);
or UO_438 (O_438,N_49521,N_49628);
and UO_439 (O_439,N_49500,N_49779);
and UO_440 (O_440,N_49828,N_49991);
nor UO_441 (O_441,N_49515,N_49976);
and UO_442 (O_442,N_49592,N_49594);
xor UO_443 (O_443,N_49528,N_49605);
nand UO_444 (O_444,N_49954,N_49659);
xor UO_445 (O_445,N_49700,N_49515);
xor UO_446 (O_446,N_49841,N_49582);
xor UO_447 (O_447,N_49537,N_49981);
and UO_448 (O_448,N_49623,N_49545);
or UO_449 (O_449,N_49648,N_49979);
or UO_450 (O_450,N_49860,N_49887);
nand UO_451 (O_451,N_49552,N_49902);
or UO_452 (O_452,N_49630,N_49552);
or UO_453 (O_453,N_49676,N_49910);
and UO_454 (O_454,N_49969,N_49898);
nand UO_455 (O_455,N_49746,N_49928);
xor UO_456 (O_456,N_49626,N_49625);
or UO_457 (O_457,N_49818,N_49902);
nor UO_458 (O_458,N_49686,N_49778);
nor UO_459 (O_459,N_49977,N_49712);
xnor UO_460 (O_460,N_49802,N_49970);
or UO_461 (O_461,N_49844,N_49866);
and UO_462 (O_462,N_49970,N_49888);
nor UO_463 (O_463,N_49693,N_49548);
nor UO_464 (O_464,N_49821,N_49581);
or UO_465 (O_465,N_49814,N_49557);
nor UO_466 (O_466,N_49559,N_49739);
xor UO_467 (O_467,N_49692,N_49508);
xnor UO_468 (O_468,N_49783,N_49964);
or UO_469 (O_469,N_49916,N_49506);
nand UO_470 (O_470,N_49612,N_49756);
and UO_471 (O_471,N_49572,N_49568);
and UO_472 (O_472,N_49964,N_49896);
nor UO_473 (O_473,N_49696,N_49693);
and UO_474 (O_474,N_49538,N_49884);
nand UO_475 (O_475,N_49908,N_49887);
xnor UO_476 (O_476,N_49905,N_49817);
nor UO_477 (O_477,N_49671,N_49751);
or UO_478 (O_478,N_49550,N_49989);
nand UO_479 (O_479,N_49919,N_49787);
nand UO_480 (O_480,N_49964,N_49583);
nor UO_481 (O_481,N_49986,N_49757);
xnor UO_482 (O_482,N_49899,N_49774);
nor UO_483 (O_483,N_49613,N_49633);
nand UO_484 (O_484,N_49520,N_49871);
nand UO_485 (O_485,N_49583,N_49872);
xnor UO_486 (O_486,N_49979,N_49793);
nand UO_487 (O_487,N_49538,N_49859);
and UO_488 (O_488,N_49834,N_49598);
xor UO_489 (O_489,N_49989,N_49994);
nand UO_490 (O_490,N_49502,N_49897);
or UO_491 (O_491,N_49662,N_49805);
or UO_492 (O_492,N_49708,N_49876);
or UO_493 (O_493,N_49658,N_49615);
and UO_494 (O_494,N_49861,N_49747);
xnor UO_495 (O_495,N_49509,N_49776);
or UO_496 (O_496,N_49928,N_49729);
nor UO_497 (O_497,N_49570,N_49826);
or UO_498 (O_498,N_49670,N_49956);
and UO_499 (O_499,N_49817,N_49751);
and UO_500 (O_500,N_49628,N_49789);
nor UO_501 (O_501,N_49612,N_49874);
or UO_502 (O_502,N_49872,N_49882);
nor UO_503 (O_503,N_49695,N_49691);
and UO_504 (O_504,N_49895,N_49672);
and UO_505 (O_505,N_49685,N_49803);
and UO_506 (O_506,N_49976,N_49969);
or UO_507 (O_507,N_49782,N_49528);
or UO_508 (O_508,N_49502,N_49583);
xnor UO_509 (O_509,N_49823,N_49667);
nand UO_510 (O_510,N_49658,N_49616);
and UO_511 (O_511,N_49783,N_49884);
or UO_512 (O_512,N_49507,N_49727);
and UO_513 (O_513,N_49595,N_49734);
nor UO_514 (O_514,N_49892,N_49840);
or UO_515 (O_515,N_49763,N_49739);
nand UO_516 (O_516,N_49527,N_49655);
or UO_517 (O_517,N_49776,N_49836);
nor UO_518 (O_518,N_49678,N_49790);
nand UO_519 (O_519,N_49985,N_49527);
nor UO_520 (O_520,N_49609,N_49819);
nor UO_521 (O_521,N_49763,N_49571);
xnor UO_522 (O_522,N_49828,N_49565);
or UO_523 (O_523,N_49835,N_49519);
xnor UO_524 (O_524,N_49862,N_49716);
and UO_525 (O_525,N_49815,N_49576);
nor UO_526 (O_526,N_49972,N_49984);
or UO_527 (O_527,N_49894,N_49656);
and UO_528 (O_528,N_49916,N_49780);
xnor UO_529 (O_529,N_49880,N_49749);
xnor UO_530 (O_530,N_49869,N_49814);
and UO_531 (O_531,N_49536,N_49819);
nor UO_532 (O_532,N_49702,N_49620);
nand UO_533 (O_533,N_49813,N_49940);
nor UO_534 (O_534,N_49755,N_49734);
nand UO_535 (O_535,N_49784,N_49996);
nor UO_536 (O_536,N_49794,N_49739);
or UO_537 (O_537,N_49909,N_49698);
nand UO_538 (O_538,N_49604,N_49688);
nand UO_539 (O_539,N_49748,N_49957);
nand UO_540 (O_540,N_49542,N_49535);
and UO_541 (O_541,N_49837,N_49619);
nand UO_542 (O_542,N_49682,N_49742);
xor UO_543 (O_543,N_49527,N_49909);
nor UO_544 (O_544,N_49869,N_49886);
xnor UO_545 (O_545,N_49533,N_49567);
or UO_546 (O_546,N_49724,N_49742);
nand UO_547 (O_547,N_49576,N_49556);
xor UO_548 (O_548,N_49939,N_49753);
nand UO_549 (O_549,N_49615,N_49909);
and UO_550 (O_550,N_49739,N_49771);
nor UO_551 (O_551,N_49802,N_49691);
xnor UO_552 (O_552,N_49924,N_49505);
nor UO_553 (O_553,N_49696,N_49945);
xor UO_554 (O_554,N_49646,N_49852);
or UO_555 (O_555,N_49606,N_49778);
and UO_556 (O_556,N_49813,N_49896);
and UO_557 (O_557,N_49532,N_49860);
xnor UO_558 (O_558,N_49711,N_49961);
nand UO_559 (O_559,N_49903,N_49839);
and UO_560 (O_560,N_49909,N_49915);
nand UO_561 (O_561,N_49752,N_49827);
and UO_562 (O_562,N_49705,N_49667);
nor UO_563 (O_563,N_49756,N_49803);
nor UO_564 (O_564,N_49847,N_49698);
xnor UO_565 (O_565,N_49913,N_49804);
and UO_566 (O_566,N_49789,N_49510);
nor UO_567 (O_567,N_49595,N_49733);
or UO_568 (O_568,N_49976,N_49991);
xnor UO_569 (O_569,N_49641,N_49811);
nand UO_570 (O_570,N_49603,N_49805);
nand UO_571 (O_571,N_49971,N_49736);
xor UO_572 (O_572,N_49943,N_49626);
and UO_573 (O_573,N_49890,N_49724);
and UO_574 (O_574,N_49842,N_49958);
nand UO_575 (O_575,N_49845,N_49767);
and UO_576 (O_576,N_49778,N_49785);
and UO_577 (O_577,N_49834,N_49547);
nor UO_578 (O_578,N_49832,N_49934);
and UO_579 (O_579,N_49765,N_49581);
nor UO_580 (O_580,N_49860,N_49677);
nor UO_581 (O_581,N_49704,N_49501);
xor UO_582 (O_582,N_49698,N_49850);
nor UO_583 (O_583,N_49584,N_49994);
xor UO_584 (O_584,N_49686,N_49616);
nor UO_585 (O_585,N_49717,N_49539);
and UO_586 (O_586,N_49586,N_49618);
nor UO_587 (O_587,N_49851,N_49670);
nand UO_588 (O_588,N_49860,N_49965);
xnor UO_589 (O_589,N_49762,N_49663);
xnor UO_590 (O_590,N_49817,N_49527);
nand UO_591 (O_591,N_49984,N_49944);
nand UO_592 (O_592,N_49513,N_49555);
nor UO_593 (O_593,N_49704,N_49964);
nor UO_594 (O_594,N_49866,N_49753);
nor UO_595 (O_595,N_49654,N_49799);
or UO_596 (O_596,N_49770,N_49834);
nand UO_597 (O_597,N_49997,N_49797);
and UO_598 (O_598,N_49527,N_49877);
and UO_599 (O_599,N_49713,N_49913);
or UO_600 (O_600,N_49667,N_49779);
xor UO_601 (O_601,N_49591,N_49579);
and UO_602 (O_602,N_49832,N_49810);
nor UO_603 (O_603,N_49943,N_49565);
or UO_604 (O_604,N_49594,N_49995);
and UO_605 (O_605,N_49922,N_49656);
or UO_606 (O_606,N_49733,N_49581);
nand UO_607 (O_607,N_49576,N_49941);
nor UO_608 (O_608,N_49754,N_49907);
nor UO_609 (O_609,N_49516,N_49842);
xor UO_610 (O_610,N_49864,N_49846);
nor UO_611 (O_611,N_49804,N_49906);
or UO_612 (O_612,N_49659,N_49928);
nor UO_613 (O_613,N_49761,N_49754);
or UO_614 (O_614,N_49634,N_49850);
or UO_615 (O_615,N_49668,N_49802);
nand UO_616 (O_616,N_49829,N_49817);
and UO_617 (O_617,N_49873,N_49541);
nor UO_618 (O_618,N_49538,N_49908);
nor UO_619 (O_619,N_49946,N_49570);
or UO_620 (O_620,N_49750,N_49795);
or UO_621 (O_621,N_49585,N_49515);
xor UO_622 (O_622,N_49878,N_49658);
nand UO_623 (O_623,N_49806,N_49874);
and UO_624 (O_624,N_49890,N_49850);
nor UO_625 (O_625,N_49931,N_49867);
nand UO_626 (O_626,N_49622,N_49742);
nor UO_627 (O_627,N_49582,N_49924);
xnor UO_628 (O_628,N_49977,N_49746);
or UO_629 (O_629,N_49876,N_49524);
nand UO_630 (O_630,N_49856,N_49922);
or UO_631 (O_631,N_49727,N_49854);
or UO_632 (O_632,N_49825,N_49969);
nor UO_633 (O_633,N_49901,N_49995);
nor UO_634 (O_634,N_49742,N_49979);
nand UO_635 (O_635,N_49786,N_49829);
nor UO_636 (O_636,N_49682,N_49501);
and UO_637 (O_637,N_49532,N_49887);
or UO_638 (O_638,N_49574,N_49779);
xor UO_639 (O_639,N_49865,N_49802);
and UO_640 (O_640,N_49714,N_49629);
and UO_641 (O_641,N_49963,N_49872);
nand UO_642 (O_642,N_49502,N_49915);
nand UO_643 (O_643,N_49751,N_49873);
and UO_644 (O_644,N_49863,N_49749);
xnor UO_645 (O_645,N_49601,N_49510);
xor UO_646 (O_646,N_49937,N_49885);
and UO_647 (O_647,N_49609,N_49516);
xor UO_648 (O_648,N_49788,N_49985);
xor UO_649 (O_649,N_49610,N_49813);
or UO_650 (O_650,N_49780,N_49995);
or UO_651 (O_651,N_49948,N_49869);
or UO_652 (O_652,N_49527,N_49953);
nor UO_653 (O_653,N_49812,N_49968);
or UO_654 (O_654,N_49545,N_49622);
xor UO_655 (O_655,N_49744,N_49978);
nor UO_656 (O_656,N_49540,N_49885);
nor UO_657 (O_657,N_49566,N_49594);
nand UO_658 (O_658,N_49755,N_49629);
nand UO_659 (O_659,N_49633,N_49980);
and UO_660 (O_660,N_49830,N_49905);
or UO_661 (O_661,N_49954,N_49703);
or UO_662 (O_662,N_49934,N_49919);
and UO_663 (O_663,N_49978,N_49571);
and UO_664 (O_664,N_49876,N_49792);
nor UO_665 (O_665,N_49936,N_49944);
and UO_666 (O_666,N_49961,N_49594);
nor UO_667 (O_667,N_49726,N_49712);
xnor UO_668 (O_668,N_49630,N_49625);
or UO_669 (O_669,N_49583,N_49678);
nor UO_670 (O_670,N_49878,N_49618);
or UO_671 (O_671,N_49577,N_49516);
xnor UO_672 (O_672,N_49731,N_49701);
and UO_673 (O_673,N_49585,N_49619);
or UO_674 (O_674,N_49666,N_49854);
xnor UO_675 (O_675,N_49576,N_49707);
or UO_676 (O_676,N_49655,N_49797);
nand UO_677 (O_677,N_49753,N_49649);
nor UO_678 (O_678,N_49930,N_49600);
nor UO_679 (O_679,N_49550,N_49531);
or UO_680 (O_680,N_49746,N_49504);
nand UO_681 (O_681,N_49846,N_49616);
nor UO_682 (O_682,N_49618,N_49770);
or UO_683 (O_683,N_49717,N_49712);
or UO_684 (O_684,N_49621,N_49855);
xnor UO_685 (O_685,N_49811,N_49564);
xor UO_686 (O_686,N_49917,N_49716);
nor UO_687 (O_687,N_49614,N_49510);
nor UO_688 (O_688,N_49791,N_49567);
xor UO_689 (O_689,N_49799,N_49744);
xnor UO_690 (O_690,N_49535,N_49887);
nand UO_691 (O_691,N_49609,N_49979);
nand UO_692 (O_692,N_49938,N_49681);
and UO_693 (O_693,N_49615,N_49501);
xnor UO_694 (O_694,N_49503,N_49899);
nor UO_695 (O_695,N_49964,N_49803);
and UO_696 (O_696,N_49511,N_49840);
nor UO_697 (O_697,N_49643,N_49805);
or UO_698 (O_698,N_49971,N_49557);
and UO_699 (O_699,N_49703,N_49869);
nand UO_700 (O_700,N_49906,N_49686);
and UO_701 (O_701,N_49795,N_49743);
and UO_702 (O_702,N_49748,N_49866);
nand UO_703 (O_703,N_49539,N_49814);
nor UO_704 (O_704,N_49648,N_49656);
nor UO_705 (O_705,N_49632,N_49784);
xor UO_706 (O_706,N_49907,N_49555);
and UO_707 (O_707,N_49988,N_49685);
nand UO_708 (O_708,N_49884,N_49800);
nor UO_709 (O_709,N_49806,N_49547);
xor UO_710 (O_710,N_49660,N_49899);
or UO_711 (O_711,N_49987,N_49504);
xor UO_712 (O_712,N_49883,N_49943);
and UO_713 (O_713,N_49635,N_49647);
and UO_714 (O_714,N_49521,N_49964);
or UO_715 (O_715,N_49514,N_49774);
xor UO_716 (O_716,N_49859,N_49874);
nor UO_717 (O_717,N_49626,N_49717);
or UO_718 (O_718,N_49896,N_49618);
and UO_719 (O_719,N_49705,N_49800);
or UO_720 (O_720,N_49893,N_49879);
or UO_721 (O_721,N_49692,N_49826);
or UO_722 (O_722,N_49700,N_49873);
nor UO_723 (O_723,N_49597,N_49834);
nor UO_724 (O_724,N_49922,N_49629);
and UO_725 (O_725,N_49945,N_49581);
or UO_726 (O_726,N_49882,N_49874);
nor UO_727 (O_727,N_49612,N_49723);
nor UO_728 (O_728,N_49962,N_49689);
xnor UO_729 (O_729,N_49527,N_49670);
or UO_730 (O_730,N_49798,N_49776);
and UO_731 (O_731,N_49506,N_49984);
xnor UO_732 (O_732,N_49681,N_49739);
or UO_733 (O_733,N_49548,N_49971);
or UO_734 (O_734,N_49764,N_49528);
and UO_735 (O_735,N_49516,N_49665);
nor UO_736 (O_736,N_49504,N_49567);
xnor UO_737 (O_737,N_49968,N_49645);
and UO_738 (O_738,N_49596,N_49663);
or UO_739 (O_739,N_49794,N_49596);
xnor UO_740 (O_740,N_49900,N_49582);
nand UO_741 (O_741,N_49872,N_49665);
nand UO_742 (O_742,N_49786,N_49884);
nand UO_743 (O_743,N_49702,N_49759);
nand UO_744 (O_744,N_49580,N_49602);
nand UO_745 (O_745,N_49793,N_49680);
or UO_746 (O_746,N_49534,N_49565);
nor UO_747 (O_747,N_49662,N_49633);
nor UO_748 (O_748,N_49984,N_49626);
and UO_749 (O_749,N_49985,N_49577);
or UO_750 (O_750,N_49564,N_49908);
or UO_751 (O_751,N_49861,N_49616);
and UO_752 (O_752,N_49705,N_49591);
nor UO_753 (O_753,N_49546,N_49955);
xnor UO_754 (O_754,N_49862,N_49949);
or UO_755 (O_755,N_49575,N_49807);
xor UO_756 (O_756,N_49635,N_49739);
and UO_757 (O_757,N_49593,N_49677);
or UO_758 (O_758,N_49867,N_49872);
or UO_759 (O_759,N_49766,N_49649);
nand UO_760 (O_760,N_49869,N_49645);
and UO_761 (O_761,N_49845,N_49756);
nand UO_762 (O_762,N_49683,N_49837);
and UO_763 (O_763,N_49916,N_49928);
and UO_764 (O_764,N_49568,N_49583);
nand UO_765 (O_765,N_49529,N_49605);
or UO_766 (O_766,N_49537,N_49881);
nand UO_767 (O_767,N_49584,N_49634);
or UO_768 (O_768,N_49945,N_49941);
nand UO_769 (O_769,N_49927,N_49914);
xnor UO_770 (O_770,N_49755,N_49679);
or UO_771 (O_771,N_49596,N_49803);
and UO_772 (O_772,N_49909,N_49531);
xor UO_773 (O_773,N_49562,N_49968);
xor UO_774 (O_774,N_49631,N_49509);
xnor UO_775 (O_775,N_49700,N_49928);
xnor UO_776 (O_776,N_49770,N_49797);
and UO_777 (O_777,N_49563,N_49644);
nor UO_778 (O_778,N_49647,N_49867);
xnor UO_779 (O_779,N_49757,N_49562);
nor UO_780 (O_780,N_49612,N_49840);
nand UO_781 (O_781,N_49584,N_49928);
or UO_782 (O_782,N_49530,N_49580);
nor UO_783 (O_783,N_49813,N_49887);
xor UO_784 (O_784,N_49683,N_49855);
xnor UO_785 (O_785,N_49587,N_49822);
and UO_786 (O_786,N_49762,N_49637);
nand UO_787 (O_787,N_49639,N_49574);
nand UO_788 (O_788,N_49844,N_49982);
and UO_789 (O_789,N_49991,N_49941);
nand UO_790 (O_790,N_49719,N_49590);
nand UO_791 (O_791,N_49974,N_49676);
nor UO_792 (O_792,N_49532,N_49697);
and UO_793 (O_793,N_49938,N_49620);
xor UO_794 (O_794,N_49942,N_49769);
xor UO_795 (O_795,N_49704,N_49930);
nor UO_796 (O_796,N_49653,N_49827);
nor UO_797 (O_797,N_49788,N_49813);
and UO_798 (O_798,N_49914,N_49824);
xnor UO_799 (O_799,N_49810,N_49936);
nand UO_800 (O_800,N_49827,N_49529);
xor UO_801 (O_801,N_49538,N_49594);
nor UO_802 (O_802,N_49796,N_49982);
nor UO_803 (O_803,N_49561,N_49593);
nand UO_804 (O_804,N_49892,N_49522);
or UO_805 (O_805,N_49520,N_49561);
nor UO_806 (O_806,N_49978,N_49811);
and UO_807 (O_807,N_49542,N_49912);
or UO_808 (O_808,N_49757,N_49936);
or UO_809 (O_809,N_49808,N_49720);
or UO_810 (O_810,N_49990,N_49714);
or UO_811 (O_811,N_49789,N_49596);
nor UO_812 (O_812,N_49720,N_49546);
nand UO_813 (O_813,N_49538,N_49756);
nor UO_814 (O_814,N_49642,N_49756);
nand UO_815 (O_815,N_49557,N_49578);
or UO_816 (O_816,N_49987,N_49664);
or UO_817 (O_817,N_49734,N_49544);
and UO_818 (O_818,N_49716,N_49811);
xnor UO_819 (O_819,N_49537,N_49701);
and UO_820 (O_820,N_49541,N_49927);
or UO_821 (O_821,N_49678,N_49965);
or UO_822 (O_822,N_49798,N_49791);
xor UO_823 (O_823,N_49709,N_49618);
and UO_824 (O_824,N_49894,N_49529);
nand UO_825 (O_825,N_49970,N_49959);
nor UO_826 (O_826,N_49895,N_49685);
xor UO_827 (O_827,N_49532,N_49650);
and UO_828 (O_828,N_49962,N_49752);
or UO_829 (O_829,N_49883,N_49840);
xnor UO_830 (O_830,N_49661,N_49617);
and UO_831 (O_831,N_49982,N_49645);
nor UO_832 (O_832,N_49934,N_49563);
nor UO_833 (O_833,N_49559,N_49893);
nand UO_834 (O_834,N_49954,N_49761);
nand UO_835 (O_835,N_49659,N_49765);
and UO_836 (O_836,N_49655,N_49823);
and UO_837 (O_837,N_49857,N_49823);
xor UO_838 (O_838,N_49558,N_49702);
nor UO_839 (O_839,N_49874,N_49541);
nand UO_840 (O_840,N_49802,N_49915);
nand UO_841 (O_841,N_49812,N_49632);
or UO_842 (O_842,N_49517,N_49760);
nor UO_843 (O_843,N_49879,N_49512);
and UO_844 (O_844,N_49535,N_49560);
and UO_845 (O_845,N_49682,N_49504);
nor UO_846 (O_846,N_49958,N_49686);
nand UO_847 (O_847,N_49733,N_49886);
nand UO_848 (O_848,N_49608,N_49576);
nor UO_849 (O_849,N_49596,N_49546);
nor UO_850 (O_850,N_49833,N_49511);
nand UO_851 (O_851,N_49835,N_49912);
nor UO_852 (O_852,N_49602,N_49630);
and UO_853 (O_853,N_49863,N_49909);
or UO_854 (O_854,N_49669,N_49931);
xnor UO_855 (O_855,N_49714,N_49931);
and UO_856 (O_856,N_49840,N_49786);
nor UO_857 (O_857,N_49915,N_49639);
xor UO_858 (O_858,N_49515,N_49961);
xnor UO_859 (O_859,N_49641,N_49666);
nand UO_860 (O_860,N_49747,N_49716);
nand UO_861 (O_861,N_49508,N_49698);
and UO_862 (O_862,N_49976,N_49844);
nor UO_863 (O_863,N_49635,N_49907);
and UO_864 (O_864,N_49648,N_49579);
and UO_865 (O_865,N_49866,N_49936);
xor UO_866 (O_866,N_49774,N_49545);
or UO_867 (O_867,N_49653,N_49937);
xnor UO_868 (O_868,N_49776,N_49844);
nand UO_869 (O_869,N_49505,N_49736);
nor UO_870 (O_870,N_49715,N_49881);
xor UO_871 (O_871,N_49905,N_49903);
and UO_872 (O_872,N_49850,N_49931);
nor UO_873 (O_873,N_49595,N_49983);
xor UO_874 (O_874,N_49626,N_49902);
or UO_875 (O_875,N_49836,N_49585);
or UO_876 (O_876,N_49947,N_49571);
and UO_877 (O_877,N_49878,N_49532);
nand UO_878 (O_878,N_49777,N_49637);
or UO_879 (O_879,N_49571,N_49525);
xor UO_880 (O_880,N_49627,N_49903);
nand UO_881 (O_881,N_49918,N_49505);
and UO_882 (O_882,N_49558,N_49640);
or UO_883 (O_883,N_49537,N_49776);
nor UO_884 (O_884,N_49814,N_49801);
or UO_885 (O_885,N_49670,N_49852);
nand UO_886 (O_886,N_49625,N_49859);
or UO_887 (O_887,N_49956,N_49792);
nor UO_888 (O_888,N_49775,N_49636);
or UO_889 (O_889,N_49910,N_49759);
nor UO_890 (O_890,N_49702,N_49582);
and UO_891 (O_891,N_49614,N_49684);
and UO_892 (O_892,N_49669,N_49594);
or UO_893 (O_893,N_49516,N_49547);
nand UO_894 (O_894,N_49655,N_49627);
nor UO_895 (O_895,N_49984,N_49666);
or UO_896 (O_896,N_49924,N_49616);
xor UO_897 (O_897,N_49533,N_49779);
nand UO_898 (O_898,N_49955,N_49602);
and UO_899 (O_899,N_49990,N_49988);
nand UO_900 (O_900,N_49720,N_49664);
nor UO_901 (O_901,N_49934,N_49791);
xnor UO_902 (O_902,N_49943,N_49953);
and UO_903 (O_903,N_49525,N_49870);
and UO_904 (O_904,N_49712,N_49826);
and UO_905 (O_905,N_49791,N_49767);
xor UO_906 (O_906,N_49630,N_49863);
nand UO_907 (O_907,N_49516,N_49919);
xor UO_908 (O_908,N_49538,N_49542);
nand UO_909 (O_909,N_49854,N_49890);
nor UO_910 (O_910,N_49718,N_49949);
nor UO_911 (O_911,N_49865,N_49503);
nor UO_912 (O_912,N_49839,N_49856);
nand UO_913 (O_913,N_49812,N_49795);
nor UO_914 (O_914,N_49585,N_49877);
nor UO_915 (O_915,N_49806,N_49795);
nor UO_916 (O_916,N_49535,N_49551);
nand UO_917 (O_917,N_49794,N_49915);
xnor UO_918 (O_918,N_49591,N_49661);
and UO_919 (O_919,N_49531,N_49634);
xnor UO_920 (O_920,N_49923,N_49951);
nor UO_921 (O_921,N_49601,N_49783);
nand UO_922 (O_922,N_49742,N_49881);
or UO_923 (O_923,N_49946,N_49613);
nor UO_924 (O_924,N_49584,N_49909);
xnor UO_925 (O_925,N_49791,N_49554);
and UO_926 (O_926,N_49620,N_49806);
or UO_927 (O_927,N_49739,N_49699);
and UO_928 (O_928,N_49608,N_49716);
and UO_929 (O_929,N_49502,N_49823);
and UO_930 (O_930,N_49558,N_49858);
and UO_931 (O_931,N_49874,N_49589);
and UO_932 (O_932,N_49701,N_49569);
nand UO_933 (O_933,N_49967,N_49551);
and UO_934 (O_934,N_49931,N_49612);
or UO_935 (O_935,N_49679,N_49702);
nor UO_936 (O_936,N_49699,N_49535);
nand UO_937 (O_937,N_49820,N_49906);
nand UO_938 (O_938,N_49882,N_49883);
nor UO_939 (O_939,N_49900,N_49668);
and UO_940 (O_940,N_49805,N_49616);
xnor UO_941 (O_941,N_49568,N_49815);
or UO_942 (O_942,N_49827,N_49561);
nor UO_943 (O_943,N_49522,N_49945);
and UO_944 (O_944,N_49981,N_49778);
xor UO_945 (O_945,N_49725,N_49956);
or UO_946 (O_946,N_49907,N_49957);
xnor UO_947 (O_947,N_49641,N_49997);
nand UO_948 (O_948,N_49550,N_49560);
or UO_949 (O_949,N_49721,N_49778);
or UO_950 (O_950,N_49929,N_49776);
nand UO_951 (O_951,N_49942,N_49937);
or UO_952 (O_952,N_49679,N_49613);
nor UO_953 (O_953,N_49698,N_49961);
and UO_954 (O_954,N_49599,N_49971);
nand UO_955 (O_955,N_49871,N_49841);
xor UO_956 (O_956,N_49807,N_49887);
nor UO_957 (O_957,N_49500,N_49861);
nand UO_958 (O_958,N_49838,N_49579);
xor UO_959 (O_959,N_49943,N_49799);
nand UO_960 (O_960,N_49757,N_49525);
or UO_961 (O_961,N_49822,N_49799);
or UO_962 (O_962,N_49745,N_49991);
and UO_963 (O_963,N_49837,N_49970);
nand UO_964 (O_964,N_49557,N_49734);
and UO_965 (O_965,N_49578,N_49963);
nand UO_966 (O_966,N_49762,N_49619);
xor UO_967 (O_967,N_49707,N_49744);
or UO_968 (O_968,N_49899,N_49859);
or UO_969 (O_969,N_49691,N_49830);
nand UO_970 (O_970,N_49685,N_49798);
nor UO_971 (O_971,N_49962,N_49992);
xor UO_972 (O_972,N_49608,N_49760);
or UO_973 (O_973,N_49975,N_49740);
nor UO_974 (O_974,N_49998,N_49904);
xor UO_975 (O_975,N_49747,N_49645);
nor UO_976 (O_976,N_49962,N_49779);
xnor UO_977 (O_977,N_49871,N_49573);
xor UO_978 (O_978,N_49665,N_49625);
xnor UO_979 (O_979,N_49899,N_49801);
nor UO_980 (O_980,N_49908,N_49775);
or UO_981 (O_981,N_49930,N_49682);
and UO_982 (O_982,N_49835,N_49770);
xor UO_983 (O_983,N_49635,N_49504);
nand UO_984 (O_984,N_49834,N_49985);
xor UO_985 (O_985,N_49601,N_49914);
or UO_986 (O_986,N_49928,N_49541);
nand UO_987 (O_987,N_49949,N_49577);
nor UO_988 (O_988,N_49604,N_49508);
and UO_989 (O_989,N_49850,N_49635);
or UO_990 (O_990,N_49773,N_49565);
and UO_991 (O_991,N_49756,N_49553);
nor UO_992 (O_992,N_49940,N_49894);
nand UO_993 (O_993,N_49523,N_49561);
nand UO_994 (O_994,N_49517,N_49850);
nand UO_995 (O_995,N_49514,N_49591);
xnor UO_996 (O_996,N_49544,N_49609);
or UO_997 (O_997,N_49603,N_49529);
nor UO_998 (O_998,N_49631,N_49758);
and UO_999 (O_999,N_49995,N_49799);
and UO_1000 (O_1000,N_49672,N_49652);
nor UO_1001 (O_1001,N_49524,N_49544);
nand UO_1002 (O_1002,N_49518,N_49600);
or UO_1003 (O_1003,N_49943,N_49720);
xnor UO_1004 (O_1004,N_49578,N_49707);
nand UO_1005 (O_1005,N_49514,N_49752);
and UO_1006 (O_1006,N_49900,N_49726);
or UO_1007 (O_1007,N_49628,N_49959);
and UO_1008 (O_1008,N_49589,N_49795);
and UO_1009 (O_1009,N_49645,N_49882);
xnor UO_1010 (O_1010,N_49766,N_49988);
xor UO_1011 (O_1011,N_49554,N_49989);
or UO_1012 (O_1012,N_49761,N_49555);
xnor UO_1013 (O_1013,N_49921,N_49980);
or UO_1014 (O_1014,N_49590,N_49959);
nand UO_1015 (O_1015,N_49585,N_49909);
xnor UO_1016 (O_1016,N_49835,N_49851);
or UO_1017 (O_1017,N_49711,N_49724);
nand UO_1018 (O_1018,N_49968,N_49844);
nand UO_1019 (O_1019,N_49753,N_49512);
and UO_1020 (O_1020,N_49574,N_49804);
and UO_1021 (O_1021,N_49895,N_49635);
nor UO_1022 (O_1022,N_49783,N_49625);
nand UO_1023 (O_1023,N_49782,N_49840);
and UO_1024 (O_1024,N_49564,N_49920);
xnor UO_1025 (O_1025,N_49965,N_49551);
nand UO_1026 (O_1026,N_49595,N_49586);
and UO_1027 (O_1027,N_49762,N_49657);
or UO_1028 (O_1028,N_49752,N_49724);
xnor UO_1029 (O_1029,N_49967,N_49979);
or UO_1030 (O_1030,N_49994,N_49781);
xor UO_1031 (O_1031,N_49673,N_49746);
xor UO_1032 (O_1032,N_49502,N_49883);
or UO_1033 (O_1033,N_49884,N_49731);
or UO_1034 (O_1034,N_49732,N_49837);
or UO_1035 (O_1035,N_49659,N_49919);
and UO_1036 (O_1036,N_49513,N_49504);
xnor UO_1037 (O_1037,N_49767,N_49841);
or UO_1038 (O_1038,N_49526,N_49514);
nor UO_1039 (O_1039,N_49614,N_49723);
and UO_1040 (O_1040,N_49978,N_49858);
and UO_1041 (O_1041,N_49836,N_49965);
nor UO_1042 (O_1042,N_49566,N_49748);
nor UO_1043 (O_1043,N_49898,N_49514);
and UO_1044 (O_1044,N_49698,N_49947);
nor UO_1045 (O_1045,N_49527,N_49514);
and UO_1046 (O_1046,N_49650,N_49597);
nor UO_1047 (O_1047,N_49949,N_49779);
or UO_1048 (O_1048,N_49989,N_49608);
nor UO_1049 (O_1049,N_49959,N_49773);
nor UO_1050 (O_1050,N_49893,N_49895);
or UO_1051 (O_1051,N_49659,N_49947);
nand UO_1052 (O_1052,N_49897,N_49507);
nand UO_1053 (O_1053,N_49864,N_49889);
or UO_1054 (O_1054,N_49683,N_49663);
and UO_1055 (O_1055,N_49663,N_49832);
xnor UO_1056 (O_1056,N_49967,N_49800);
and UO_1057 (O_1057,N_49558,N_49881);
and UO_1058 (O_1058,N_49525,N_49622);
nand UO_1059 (O_1059,N_49711,N_49526);
or UO_1060 (O_1060,N_49790,N_49633);
xor UO_1061 (O_1061,N_49714,N_49837);
and UO_1062 (O_1062,N_49583,N_49837);
and UO_1063 (O_1063,N_49804,N_49512);
or UO_1064 (O_1064,N_49642,N_49709);
xnor UO_1065 (O_1065,N_49910,N_49633);
and UO_1066 (O_1066,N_49623,N_49872);
and UO_1067 (O_1067,N_49626,N_49971);
and UO_1068 (O_1068,N_49969,N_49570);
and UO_1069 (O_1069,N_49578,N_49534);
nand UO_1070 (O_1070,N_49836,N_49659);
xnor UO_1071 (O_1071,N_49557,N_49721);
or UO_1072 (O_1072,N_49922,N_49837);
and UO_1073 (O_1073,N_49735,N_49940);
or UO_1074 (O_1074,N_49736,N_49899);
and UO_1075 (O_1075,N_49890,N_49885);
and UO_1076 (O_1076,N_49546,N_49906);
nor UO_1077 (O_1077,N_49513,N_49875);
nand UO_1078 (O_1078,N_49580,N_49622);
nor UO_1079 (O_1079,N_49654,N_49810);
or UO_1080 (O_1080,N_49903,N_49561);
nor UO_1081 (O_1081,N_49768,N_49992);
nand UO_1082 (O_1082,N_49748,N_49867);
nor UO_1083 (O_1083,N_49682,N_49794);
nand UO_1084 (O_1084,N_49861,N_49879);
nand UO_1085 (O_1085,N_49579,N_49517);
nand UO_1086 (O_1086,N_49820,N_49600);
and UO_1087 (O_1087,N_49989,N_49655);
xnor UO_1088 (O_1088,N_49983,N_49563);
or UO_1089 (O_1089,N_49949,N_49505);
or UO_1090 (O_1090,N_49930,N_49512);
xnor UO_1091 (O_1091,N_49583,N_49976);
and UO_1092 (O_1092,N_49744,N_49779);
xnor UO_1093 (O_1093,N_49974,N_49729);
nand UO_1094 (O_1094,N_49567,N_49647);
or UO_1095 (O_1095,N_49654,N_49867);
xnor UO_1096 (O_1096,N_49895,N_49537);
nor UO_1097 (O_1097,N_49546,N_49964);
and UO_1098 (O_1098,N_49867,N_49605);
nor UO_1099 (O_1099,N_49933,N_49805);
xor UO_1100 (O_1100,N_49767,N_49787);
nor UO_1101 (O_1101,N_49537,N_49676);
or UO_1102 (O_1102,N_49510,N_49890);
nor UO_1103 (O_1103,N_49561,N_49694);
nand UO_1104 (O_1104,N_49922,N_49630);
xnor UO_1105 (O_1105,N_49667,N_49908);
or UO_1106 (O_1106,N_49992,N_49668);
xor UO_1107 (O_1107,N_49518,N_49765);
nor UO_1108 (O_1108,N_49873,N_49660);
nor UO_1109 (O_1109,N_49945,N_49703);
xor UO_1110 (O_1110,N_49801,N_49528);
nor UO_1111 (O_1111,N_49761,N_49842);
nor UO_1112 (O_1112,N_49561,N_49908);
nor UO_1113 (O_1113,N_49660,N_49900);
xor UO_1114 (O_1114,N_49914,N_49813);
or UO_1115 (O_1115,N_49555,N_49522);
nor UO_1116 (O_1116,N_49645,N_49737);
or UO_1117 (O_1117,N_49671,N_49532);
and UO_1118 (O_1118,N_49790,N_49771);
or UO_1119 (O_1119,N_49819,N_49544);
xnor UO_1120 (O_1120,N_49803,N_49953);
nor UO_1121 (O_1121,N_49897,N_49753);
or UO_1122 (O_1122,N_49601,N_49528);
nand UO_1123 (O_1123,N_49608,N_49931);
xnor UO_1124 (O_1124,N_49519,N_49858);
nor UO_1125 (O_1125,N_49990,N_49930);
and UO_1126 (O_1126,N_49587,N_49897);
and UO_1127 (O_1127,N_49696,N_49583);
xnor UO_1128 (O_1128,N_49859,N_49796);
nor UO_1129 (O_1129,N_49735,N_49998);
nor UO_1130 (O_1130,N_49678,N_49868);
nand UO_1131 (O_1131,N_49661,N_49903);
and UO_1132 (O_1132,N_49610,N_49754);
nand UO_1133 (O_1133,N_49722,N_49923);
nor UO_1134 (O_1134,N_49736,N_49580);
nand UO_1135 (O_1135,N_49666,N_49715);
nand UO_1136 (O_1136,N_49900,N_49607);
nand UO_1137 (O_1137,N_49700,N_49643);
xor UO_1138 (O_1138,N_49884,N_49717);
nor UO_1139 (O_1139,N_49774,N_49942);
or UO_1140 (O_1140,N_49949,N_49629);
and UO_1141 (O_1141,N_49720,N_49617);
and UO_1142 (O_1142,N_49550,N_49976);
xor UO_1143 (O_1143,N_49647,N_49978);
and UO_1144 (O_1144,N_49645,N_49537);
nand UO_1145 (O_1145,N_49970,N_49890);
nor UO_1146 (O_1146,N_49907,N_49982);
or UO_1147 (O_1147,N_49952,N_49595);
and UO_1148 (O_1148,N_49629,N_49981);
or UO_1149 (O_1149,N_49990,N_49872);
xor UO_1150 (O_1150,N_49632,N_49979);
nand UO_1151 (O_1151,N_49674,N_49945);
or UO_1152 (O_1152,N_49606,N_49700);
nor UO_1153 (O_1153,N_49838,N_49692);
or UO_1154 (O_1154,N_49591,N_49726);
or UO_1155 (O_1155,N_49748,N_49500);
nand UO_1156 (O_1156,N_49951,N_49962);
nand UO_1157 (O_1157,N_49847,N_49980);
and UO_1158 (O_1158,N_49842,N_49541);
xor UO_1159 (O_1159,N_49954,N_49826);
or UO_1160 (O_1160,N_49996,N_49828);
nor UO_1161 (O_1161,N_49934,N_49883);
or UO_1162 (O_1162,N_49614,N_49594);
or UO_1163 (O_1163,N_49971,N_49891);
and UO_1164 (O_1164,N_49863,N_49990);
xnor UO_1165 (O_1165,N_49936,N_49786);
nand UO_1166 (O_1166,N_49512,N_49841);
or UO_1167 (O_1167,N_49881,N_49571);
nand UO_1168 (O_1168,N_49647,N_49577);
nor UO_1169 (O_1169,N_49504,N_49588);
nor UO_1170 (O_1170,N_49569,N_49612);
nor UO_1171 (O_1171,N_49962,N_49702);
xor UO_1172 (O_1172,N_49922,N_49541);
xnor UO_1173 (O_1173,N_49513,N_49680);
xnor UO_1174 (O_1174,N_49586,N_49623);
xor UO_1175 (O_1175,N_49983,N_49956);
xor UO_1176 (O_1176,N_49589,N_49989);
xnor UO_1177 (O_1177,N_49765,N_49996);
xnor UO_1178 (O_1178,N_49646,N_49804);
nor UO_1179 (O_1179,N_49688,N_49652);
nand UO_1180 (O_1180,N_49517,N_49897);
and UO_1181 (O_1181,N_49515,N_49630);
nand UO_1182 (O_1182,N_49969,N_49935);
and UO_1183 (O_1183,N_49749,N_49762);
and UO_1184 (O_1184,N_49654,N_49748);
xor UO_1185 (O_1185,N_49625,N_49850);
or UO_1186 (O_1186,N_49710,N_49722);
nor UO_1187 (O_1187,N_49615,N_49993);
xnor UO_1188 (O_1188,N_49707,N_49709);
and UO_1189 (O_1189,N_49985,N_49960);
xor UO_1190 (O_1190,N_49778,N_49727);
nand UO_1191 (O_1191,N_49513,N_49729);
and UO_1192 (O_1192,N_49845,N_49976);
or UO_1193 (O_1193,N_49998,N_49649);
or UO_1194 (O_1194,N_49562,N_49980);
nor UO_1195 (O_1195,N_49830,N_49827);
or UO_1196 (O_1196,N_49899,N_49776);
or UO_1197 (O_1197,N_49733,N_49762);
or UO_1198 (O_1198,N_49695,N_49766);
nor UO_1199 (O_1199,N_49935,N_49873);
nand UO_1200 (O_1200,N_49999,N_49615);
nand UO_1201 (O_1201,N_49847,N_49507);
or UO_1202 (O_1202,N_49749,N_49745);
nor UO_1203 (O_1203,N_49890,N_49851);
nand UO_1204 (O_1204,N_49686,N_49656);
or UO_1205 (O_1205,N_49981,N_49766);
xor UO_1206 (O_1206,N_49634,N_49664);
or UO_1207 (O_1207,N_49930,N_49620);
or UO_1208 (O_1208,N_49776,N_49788);
and UO_1209 (O_1209,N_49712,N_49701);
and UO_1210 (O_1210,N_49790,N_49750);
or UO_1211 (O_1211,N_49756,N_49761);
nand UO_1212 (O_1212,N_49997,N_49848);
xnor UO_1213 (O_1213,N_49659,N_49719);
and UO_1214 (O_1214,N_49722,N_49725);
or UO_1215 (O_1215,N_49802,N_49990);
nand UO_1216 (O_1216,N_49806,N_49847);
or UO_1217 (O_1217,N_49791,N_49698);
nand UO_1218 (O_1218,N_49561,N_49859);
or UO_1219 (O_1219,N_49672,N_49633);
xor UO_1220 (O_1220,N_49795,N_49684);
nand UO_1221 (O_1221,N_49760,N_49826);
xor UO_1222 (O_1222,N_49515,N_49933);
nor UO_1223 (O_1223,N_49650,N_49787);
xor UO_1224 (O_1224,N_49785,N_49788);
xor UO_1225 (O_1225,N_49737,N_49704);
or UO_1226 (O_1226,N_49781,N_49635);
nand UO_1227 (O_1227,N_49764,N_49979);
nand UO_1228 (O_1228,N_49571,N_49535);
and UO_1229 (O_1229,N_49966,N_49710);
and UO_1230 (O_1230,N_49908,N_49816);
xnor UO_1231 (O_1231,N_49820,N_49968);
xor UO_1232 (O_1232,N_49690,N_49864);
or UO_1233 (O_1233,N_49557,N_49614);
or UO_1234 (O_1234,N_49576,N_49739);
or UO_1235 (O_1235,N_49959,N_49935);
or UO_1236 (O_1236,N_49940,N_49956);
xnor UO_1237 (O_1237,N_49740,N_49689);
and UO_1238 (O_1238,N_49910,N_49831);
and UO_1239 (O_1239,N_49820,N_49547);
nand UO_1240 (O_1240,N_49528,N_49749);
and UO_1241 (O_1241,N_49732,N_49597);
or UO_1242 (O_1242,N_49682,N_49721);
nand UO_1243 (O_1243,N_49868,N_49774);
nand UO_1244 (O_1244,N_49670,N_49718);
xnor UO_1245 (O_1245,N_49657,N_49565);
nand UO_1246 (O_1246,N_49683,N_49593);
or UO_1247 (O_1247,N_49917,N_49644);
xnor UO_1248 (O_1248,N_49695,N_49515);
nor UO_1249 (O_1249,N_49954,N_49828);
or UO_1250 (O_1250,N_49931,N_49685);
nor UO_1251 (O_1251,N_49516,N_49542);
or UO_1252 (O_1252,N_49782,N_49771);
nand UO_1253 (O_1253,N_49542,N_49811);
xor UO_1254 (O_1254,N_49557,N_49566);
nand UO_1255 (O_1255,N_49689,N_49835);
or UO_1256 (O_1256,N_49697,N_49827);
nand UO_1257 (O_1257,N_49971,N_49674);
nand UO_1258 (O_1258,N_49744,N_49775);
nand UO_1259 (O_1259,N_49579,N_49504);
xor UO_1260 (O_1260,N_49767,N_49675);
xnor UO_1261 (O_1261,N_49580,N_49547);
nor UO_1262 (O_1262,N_49924,N_49774);
nand UO_1263 (O_1263,N_49569,N_49596);
and UO_1264 (O_1264,N_49570,N_49901);
xnor UO_1265 (O_1265,N_49577,N_49645);
xor UO_1266 (O_1266,N_49502,N_49854);
nand UO_1267 (O_1267,N_49566,N_49847);
or UO_1268 (O_1268,N_49822,N_49510);
nor UO_1269 (O_1269,N_49722,N_49836);
and UO_1270 (O_1270,N_49660,N_49787);
and UO_1271 (O_1271,N_49724,N_49591);
xnor UO_1272 (O_1272,N_49695,N_49910);
nand UO_1273 (O_1273,N_49708,N_49562);
nand UO_1274 (O_1274,N_49561,N_49739);
and UO_1275 (O_1275,N_49704,N_49648);
nor UO_1276 (O_1276,N_49785,N_49801);
xor UO_1277 (O_1277,N_49949,N_49827);
and UO_1278 (O_1278,N_49816,N_49722);
or UO_1279 (O_1279,N_49683,N_49878);
or UO_1280 (O_1280,N_49743,N_49519);
or UO_1281 (O_1281,N_49765,N_49792);
xnor UO_1282 (O_1282,N_49955,N_49524);
nand UO_1283 (O_1283,N_49828,N_49514);
and UO_1284 (O_1284,N_49652,N_49619);
nor UO_1285 (O_1285,N_49961,N_49598);
nor UO_1286 (O_1286,N_49793,N_49740);
and UO_1287 (O_1287,N_49949,N_49712);
and UO_1288 (O_1288,N_49738,N_49796);
xor UO_1289 (O_1289,N_49884,N_49559);
xor UO_1290 (O_1290,N_49610,N_49840);
nand UO_1291 (O_1291,N_49501,N_49562);
nand UO_1292 (O_1292,N_49868,N_49912);
nor UO_1293 (O_1293,N_49927,N_49791);
nand UO_1294 (O_1294,N_49975,N_49563);
nand UO_1295 (O_1295,N_49677,N_49820);
or UO_1296 (O_1296,N_49842,N_49902);
nor UO_1297 (O_1297,N_49767,N_49706);
nand UO_1298 (O_1298,N_49688,N_49984);
or UO_1299 (O_1299,N_49681,N_49855);
or UO_1300 (O_1300,N_49643,N_49682);
nor UO_1301 (O_1301,N_49597,N_49640);
nand UO_1302 (O_1302,N_49703,N_49766);
nand UO_1303 (O_1303,N_49639,N_49878);
xnor UO_1304 (O_1304,N_49978,N_49592);
nand UO_1305 (O_1305,N_49770,N_49636);
and UO_1306 (O_1306,N_49887,N_49990);
and UO_1307 (O_1307,N_49968,N_49963);
nor UO_1308 (O_1308,N_49780,N_49625);
nand UO_1309 (O_1309,N_49987,N_49751);
xor UO_1310 (O_1310,N_49877,N_49869);
nand UO_1311 (O_1311,N_49538,N_49778);
or UO_1312 (O_1312,N_49691,N_49503);
or UO_1313 (O_1313,N_49936,N_49701);
nor UO_1314 (O_1314,N_49722,N_49907);
and UO_1315 (O_1315,N_49613,N_49944);
xnor UO_1316 (O_1316,N_49746,N_49836);
xnor UO_1317 (O_1317,N_49709,N_49794);
nor UO_1318 (O_1318,N_49980,N_49995);
and UO_1319 (O_1319,N_49830,N_49657);
or UO_1320 (O_1320,N_49981,N_49945);
and UO_1321 (O_1321,N_49792,N_49775);
xnor UO_1322 (O_1322,N_49901,N_49874);
and UO_1323 (O_1323,N_49571,N_49536);
and UO_1324 (O_1324,N_49789,N_49757);
nand UO_1325 (O_1325,N_49808,N_49609);
nor UO_1326 (O_1326,N_49945,N_49574);
nand UO_1327 (O_1327,N_49949,N_49850);
xor UO_1328 (O_1328,N_49983,N_49836);
xor UO_1329 (O_1329,N_49812,N_49516);
or UO_1330 (O_1330,N_49562,N_49644);
xnor UO_1331 (O_1331,N_49714,N_49554);
xnor UO_1332 (O_1332,N_49793,N_49921);
xor UO_1333 (O_1333,N_49696,N_49750);
and UO_1334 (O_1334,N_49968,N_49590);
and UO_1335 (O_1335,N_49918,N_49540);
nor UO_1336 (O_1336,N_49884,N_49509);
nand UO_1337 (O_1337,N_49971,N_49632);
xor UO_1338 (O_1338,N_49819,N_49587);
and UO_1339 (O_1339,N_49687,N_49689);
nor UO_1340 (O_1340,N_49998,N_49677);
and UO_1341 (O_1341,N_49982,N_49914);
or UO_1342 (O_1342,N_49935,N_49877);
and UO_1343 (O_1343,N_49582,N_49944);
nor UO_1344 (O_1344,N_49617,N_49807);
and UO_1345 (O_1345,N_49565,N_49551);
xnor UO_1346 (O_1346,N_49614,N_49895);
and UO_1347 (O_1347,N_49810,N_49765);
nand UO_1348 (O_1348,N_49926,N_49741);
xnor UO_1349 (O_1349,N_49602,N_49686);
or UO_1350 (O_1350,N_49585,N_49525);
nand UO_1351 (O_1351,N_49686,N_49931);
nor UO_1352 (O_1352,N_49534,N_49665);
and UO_1353 (O_1353,N_49702,N_49824);
and UO_1354 (O_1354,N_49723,N_49704);
xor UO_1355 (O_1355,N_49896,N_49533);
nand UO_1356 (O_1356,N_49571,N_49876);
and UO_1357 (O_1357,N_49998,N_49597);
xnor UO_1358 (O_1358,N_49857,N_49770);
or UO_1359 (O_1359,N_49740,N_49538);
or UO_1360 (O_1360,N_49775,N_49674);
xor UO_1361 (O_1361,N_49816,N_49527);
nor UO_1362 (O_1362,N_49593,N_49565);
or UO_1363 (O_1363,N_49682,N_49951);
nor UO_1364 (O_1364,N_49928,N_49731);
nor UO_1365 (O_1365,N_49685,N_49584);
xor UO_1366 (O_1366,N_49960,N_49666);
xnor UO_1367 (O_1367,N_49894,N_49666);
xor UO_1368 (O_1368,N_49878,N_49535);
or UO_1369 (O_1369,N_49951,N_49976);
xor UO_1370 (O_1370,N_49995,N_49836);
or UO_1371 (O_1371,N_49834,N_49972);
nand UO_1372 (O_1372,N_49681,N_49902);
nand UO_1373 (O_1373,N_49893,N_49681);
nand UO_1374 (O_1374,N_49703,N_49768);
nand UO_1375 (O_1375,N_49803,N_49836);
xor UO_1376 (O_1376,N_49948,N_49611);
nand UO_1377 (O_1377,N_49668,N_49704);
or UO_1378 (O_1378,N_49827,N_49568);
nand UO_1379 (O_1379,N_49716,N_49529);
and UO_1380 (O_1380,N_49515,N_49502);
nand UO_1381 (O_1381,N_49937,N_49567);
or UO_1382 (O_1382,N_49980,N_49707);
nor UO_1383 (O_1383,N_49953,N_49549);
xnor UO_1384 (O_1384,N_49528,N_49607);
and UO_1385 (O_1385,N_49718,N_49838);
or UO_1386 (O_1386,N_49824,N_49815);
and UO_1387 (O_1387,N_49908,N_49508);
or UO_1388 (O_1388,N_49542,N_49500);
or UO_1389 (O_1389,N_49716,N_49704);
or UO_1390 (O_1390,N_49673,N_49669);
xor UO_1391 (O_1391,N_49515,N_49550);
or UO_1392 (O_1392,N_49867,N_49964);
nor UO_1393 (O_1393,N_49956,N_49767);
xor UO_1394 (O_1394,N_49528,N_49715);
nor UO_1395 (O_1395,N_49624,N_49903);
xor UO_1396 (O_1396,N_49712,N_49984);
nor UO_1397 (O_1397,N_49810,N_49709);
xor UO_1398 (O_1398,N_49712,N_49611);
and UO_1399 (O_1399,N_49864,N_49691);
nor UO_1400 (O_1400,N_49872,N_49813);
nor UO_1401 (O_1401,N_49894,N_49743);
xor UO_1402 (O_1402,N_49579,N_49635);
xor UO_1403 (O_1403,N_49833,N_49985);
nand UO_1404 (O_1404,N_49969,N_49773);
nor UO_1405 (O_1405,N_49706,N_49749);
or UO_1406 (O_1406,N_49874,N_49572);
nand UO_1407 (O_1407,N_49874,N_49830);
xor UO_1408 (O_1408,N_49706,N_49531);
or UO_1409 (O_1409,N_49686,N_49997);
and UO_1410 (O_1410,N_49839,N_49764);
and UO_1411 (O_1411,N_49571,N_49870);
and UO_1412 (O_1412,N_49545,N_49743);
nand UO_1413 (O_1413,N_49782,N_49629);
nand UO_1414 (O_1414,N_49628,N_49675);
or UO_1415 (O_1415,N_49765,N_49504);
or UO_1416 (O_1416,N_49761,N_49610);
nand UO_1417 (O_1417,N_49851,N_49610);
and UO_1418 (O_1418,N_49906,N_49544);
and UO_1419 (O_1419,N_49721,N_49523);
or UO_1420 (O_1420,N_49834,N_49524);
nor UO_1421 (O_1421,N_49941,N_49707);
and UO_1422 (O_1422,N_49954,N_49849);
nor UO_1423 (O_1423,N_49603,N_49736);
nor UO_1424 (O_1424,N_49701,N_49744);
nand UO_1425 (O_1425,N_49868,N_49762);
xnor UO_1426 (O_1426,N_49745,N_49622);
nor UO_1427 (O_1427,N_49870,N_49623);
or UO_1428 (O_1428,N_49669,N_49731);
nor UO_1429 (O_1429,N_49757,N_49580);
or UO_1430 (O_1430,N_49722,N_49928);
xor UO_1431 (O_1431,N_49640,N_49690);
or UO_1432 (O_1432,N_49544,N_49760);
or UO_1433 (O_1433,N_49900,N_49783);
and UO_1434 (O_1434,N_49934,N_49863);
and UO_1435 (O_1435,N_49917,N_49555);
xor UO_1436 (O_1436,N_49531,N_49841);
nand UO_1437 (O_1437,N_49805,N_49975);
nor UO_1438 (O_1438,N_49897,N_49577);
xor UO_1439 (O_1439,N_49882,N_49772);
or UO_1440 (O_1440,N_49998,N_49583);
nand UO_1441 (O_1441,N_49855,N_49964);
nand UO_1442 (O_1442,N_49998,N_49603);
or UO_1443 (O_1443,N_49660,N_49617);
nor UO_1444 (O_1444,N_49723,N_49526);
nor UO_1445 (O_1445,N_49628,N_49712);
and UO_1446 (O_1446,N_49773,N_49923);
nand UO_1447 (O_1447,N_49520,N_49553);
nand UO_1448 (O_1448,N_49690,N_49949);
xor UO_1449 (O_1449,N_49821,N_49689);
xor UO_1450 (O_1450,N_49680,N_49593);
and UO_1451 (O_1451,N_49727,N_49964);
or UO_1452 (O_1452,N_49785,N_49616);
or UO_1453 (O_1453,N_49789,N_49594);
nand UO_1454 (O_1454,N_49590,N_49824);
nand UO_1455 (O_1455,N_49580,N_49921);
and UO_1456 (O_1456,N_49781,N_49552);
nor UO_1457 (O_1457,N_49655,N_49819);
nand UO_1458 (O_1458,N_49589,N_49705);
nor UO_1459 (O_1459,N_49540,N_49654);
xnor UO_1460 (O_1460,N_49939,N_49793);
xor UO_1461 (O_1461,N_49506,N_49722);
nand UO_1462 (O_1462,N_49597,N_49535);
nand UO_1463 (O_1463,N_49553,N_49879);
and UO_1464 (O_1464,N_49653,N_49835);
or UO_1465 (O_1465,N_49937,N_49756);
xor UO_1466 (O_1466,N_49645,N_49909);
and UO_1467 (O_1467,N_49904,N_49508);
xnor UO_1468 (O_1468,N_49739,N_49608);
nand UO_1469 (O_1469,N_49802,N_49967);
nand UO_1470 (O_1470,N_49872,N_49678);
xor UO_1471 (O_1471,N_49537,N_49626);
nor UO_1472 (O_1472,N_49704,N_49580);
nor UO_1473 (O_1473,N_49945,N_49590);
nand UO_1474 (O_1474,N_49807,N_49995);
nor UO_1475 (O_1475,N_49834,N_49861);
xnor UO_1476 (O_1476,N_49522,N_49725);
nand UO_1477 (O_1477,N_49930,N_49980);
and UO_1478 (O_1478,N_49934,N_49940);
nand UO_1479 (O_1479,N_49969,N_49949);
and UO_1480 (O_1480,N_49964,N_49513);
xnor UO_1481 (O_1481,N_49612,N_49834);
xor UO_1482 (O_1482,N_49958,N_49797);
nand UO_1483 (O_1483,N_49633,N_49909);
or UO_1484 (O_1484,N_49505,N_49993);
nor UO_1485 (O_1485,N_49525,N_49918);
xor UO_1486 (O_1486,N_49629,N_49728);
nand UO_1487 (O_1487,N_49518,N_49591);
and UO_1488 (O_1488,N_49592,N_49817);
or UO_1489 (O_1489,N_49561,N_49754);
or UO_1490 (O_1490,N_49757,N_49823);
xnor UO_1491 (O_1491,N_49548,N_49759);
nor UO_1492 (O_1492,N_49612,N_49884);
nor UO_1493 (O_1493,N_49811,N_49795);
xnor UO_1494 (O_1494,N_49642,N_49740);
or UO_1495 (O_1495,N_49858,N_49636);
nor UO_1496 (O_1496,N_49509,N_49817);
or UO_1497 (O_1497,N_49704,N_49743);
nor UO_1498 (O_1498,N_49522,N_49878);
nand UO_1499 (O_1499,N_49588,N_49653);
or UO_1500 (O_1500,N_49711,N_49968);
nand UO_1501 (O_1501,N_49649,N_49733);
or UO_1502 (O_1502,N_49696,N_49646);
and UO_1503 (O_1503,N_49922,N_49964);
nand UO_1504 (O_1504,N_49776,N_49635);
or UO_1505 (O_1505,N_49935,N_49764);
xnor UO_1506 (O_1506,N_49852,N_49511);
or UO_1507 (O_1507,N_49996,N_49696);
nor UO_1508 (O_1508,N_49557,N_49577);
or UO_1509 (O_1509,N_49669,N_49582);
and UO_1510 (O_1510,N_49859,N_49818);
nor UO_1511 (O_1511,N_49778,N_49651);
nor UO_1512 (O_1512,N_49838,N_49625);
nor UO_1513 (O_1513,N_49565,N_49969);
nand UO_1514 (O_1514,N_49833,N_49684);
xor UO_1515 (O_1515,N_49668,N_49675);
or UO_1516 (O_1516,N_49694,N_49638);
nor UO_1517 (O_1517,N_49910,N_49996);
nand UO_1518 (O_1518,N_49509,N_49979);
and UO_1519 (O_1519,N_49690,N_49565);
nand UO_1520 (O_1520,N_49950,N_49503);
or UO_1521 (O_1521,N_49908,N_49979);
nand UO_1522 (O_1522,N_49621,N_49654);
xnor UO_1523 (O_1523,N_49825,N_49900);
nor UO_1524 (O_1524,N_49754,N_49775);
xnor UO_1525 (O_1525,N_49887,N_49609);
xnor UO_1526 (O_1526,N_49966,N_49852);
or UO_1527 (O_1527,N_49598,N_49896);
and UO_1528 (O_1528,N_49731,N_49981);
xnor UO_1529 (O_1529,N_49972,N_49783);
xor UO_1530 (O_1530,N_49936,N_49588);
xor UO_1531 (O_1531,N_49997,N_49780);
nor UO_1532 (O_1532,N_49943,N_49702);
nand UO_1533 (O_1533,N_49597,N_49906);
nor UO_1534 (O_1534,N_49617,N_49970);
and UO_1535 (O_1535,N_49945,N_49950);
or UO_1536 (O_1536,N_49581,N_49991);
xor UO_1537 (O_1537,N_49747,N_49772);
or UO_1538 (O_1538,N_49708,N_49960);
or UO_1539 (O_1539,N_49712,N_49627);
xnor UO_1540 (O_1540,N_49871,N_49943);
nor UO_1541 (O_1541,N_49983,N_49682);
xor UO_1542 (O_1542,N_49768,N_49889);
nor UO_1543 (O_1543,N_49986,N_49653);
and UO_1544 (O_1544,N_49738,N_49935);
nor UO_1545 (O_1545,N_49513,N_49582);
xnor UO_1546 (O_1546,N_49715,N_49581);
nor UO_1547 (O_1547,N_49577,N_49781);
nor UO_1548 (O_1548,N_49845,N_49783);
xor UO_1549 (O_1549,N_49713,N_49863);
nand UO_1550 (O_1550,N_49639,N_49501);
nor UO_1551 (O_1551,N_49988,N_49765);
nor UO_1552 (O_1552,N_49516,N_49599);
xor UO_1553 (O_1553,N_49793,N_49829);
nor UO_1554 (O_1554,N_49846,N_49679);
nand UO_1555 (O_1555,N_49779,N_49682);
nor UO_1556 (O_1556,N_49595,N_49737);
or UO_1557 (O_1557,N_49944,N_49852);
nor UO_1558 (O_1558,N_49747,N_49780);
and UO_1559 (O_1559,N_49774,N_49624);
nor UO_1560 (O_1560,N_49779,N_49903);
or UO_1561 (O_1561,N_49726,N_49888);
nand UO_1562 (O_1562,N_49915,N_49756);
xnor UO_1563 (O_1563,N_49568,N_49921);
or UO_1564 (O_1564,N_49640,N_49846);
xor UO_1565 (O_1565,N_49799,N_49552);
and UO_1566 (O_1566,N_49948,N_49738);
or UO_1567 (O_1567,N_49830,N_49677);
or UO_1568 (O_1568,N_49858,N_49712);
and UO_1569 (O_1569,N_49654,N_49615);
and UO_1570 (O_1570,N_49929,N_49748);
nor UO_1571 (O_1571,N_49700,N_49715);
and UO_1572 (O_1572,N_49506,N_49757);
nor UO_1573 (O_1573,N_49913,N_49999);
and UO_1574 (O_1574,N_49688,N_49581);
nor UO_1575 (O_1575,N_49894,N_49977);
or UO_1576 (O_1576,N_49773,N_49612);
or UO_1577 (O_1577,N_49753,N_49709);
or UO_1578 (O_1578,N_49577,N_49703);
xor UO_1579 (O_1579,N_49936,N_49893);
nand UO_1580 (O_1580,N_49968,N_49634);
nand UO_1581 (O_1581,N_49889,N_49695);
xor UO_1582 (O_1582,N_49984,N_49701);
nor UO_1583 (O_1583,N_49712,N_49851);
nand UO_1584 (O_1584,N_49597,N_49940);
and UO_1585 (O_1585,N_49626,N_49705);
nor UO_1586 (O_1586,N_49502,N_49617);
nand UO_1587 (O_1587,N_49743,N_49670);
nor UO_1588 (O_1588,N_49690,N_49919);
or UO_1589 (O_1589,N_49546,N_49779);
nand UO_1590 (O_1590,N_49544,N_49718);
and UO_1591 (O_1591,N_49708,N_49832);
and UO_1592 (O_1592,N_49521,N_49641);
xnor UO_1593 (O_1593,N_49872,N_49768);
nor UO_1594 (O_1594,N_49715,N_49931);
and UO_1595 (O_1595,N_49643,N_49621);
nand UO_1596 (O_1596,N_49836,N_49914);
and UO_1597 (O_1597,N_49729,N_49602);
xor UO_1598 (O_1598,N_49952,N_49859);
or UO_1599 (O_1599,N_49891,N_49669);
or UO_1600 (O_1600,N_49805,N_49922);
xnor UO_1601 (O_1601,N_49570,N_49547);
xnor UO_1602 (O_1602,N_49770,N_49869);
or UO_1603 (O_1603,N_49621,N_49750);
nor UO_1604 (O_1604,N_49604,N_49922);
nand UO_1605 (O_1605,N_49868,N_49669);
nand UO_1606 (O_1606,N_49538,N_49949);
nor UO_1607 (O_1607,N_49525,N_49947);
nor UO_1608 (O_1608,N_49552,N_49756);
nor UO_1609 (O_1609,N_49864,N_49926);
or UO_1610 (O_1610,N_49830,N_49721);
xor UO_1611 (O_1611,N_49705,N_49728);
nand UO_1612 (O_1612,N_49506,N_49517);
or UO_1613 (O_1613,N_49947,N_49961);
or UO_1614 (O_1614,N_49808,N_49977);
or UO_1615 (O_1615,N_49692,N_49969);
nor UO_1616 (O_1616,N_49944,N_49759);
nand UO_1617 (O_1617,N_49531,N_49859);
and UO_1618 (O_1618,N_49663,N_49983);
nor UO_1619 (O_1619,N_49792,N_49645);
xor UO_1620 (O_1620,N_49578,N_49651);
xor UO_1621 (O_1621,N_49733,N_49707);
and UO_1622 (O_1622,N_49892,N_49808);
nor UO_1623 (O_1623,N_49964,N_49957);
xnor UO_1624 (O_1624,N_49599,N_49514);
xnor UO_1625 (O_1625,N_49738,N_49730);
or UO_1626 (O_1626,N_49866,N_49688);
and UO_1627 (O_1627,N_49629,N_49910);
xor UO_1628 (O_1628,N_49775,N_49995);
or UO_1629 (O_1629,N_49949,N_49925);
nor UO_1630 (O_1630,N_49832,N_49770);
nand UO_1631 (O_1631,N_49864,N_49990);
and UO_1632 (O_1632,N_49760,N_49665);
nor UO_1633 (O_1633,N_49922,N_49618);
xnor UO_1634 (O_1634,N_49785,N_49544);
nand UO_1635 (O_1635,N_49820,N_49983);
nand UO_1636 (O_1636,N_49714,N_49526);
nor UO_1637 (O_1637,N_49702,N_49860);
nand UO_1638 (O_1638,N_49965,N_49746);
nor UO_1639 (O_1639,N_49567,N_49730);
or UO_1640 (O_1640,N_49864,N_49709);
nand UO_1641 (O_1641,N_49984,N_49861);
nor UO_1642 (O_1642,N_49849,N_49616);
xnor UO_1643 (O_1643,N_49540,N_49910);
xnor UO_1644 (O_1644,N_49812,N_49905);
xnor UO_1645 (O_1645,N_49954,N_49710);
nand UO_1646 (O_1646,N_49778,N_49853);
and UO_1647 (O_1647,N_49674,N_49934);
xor UO_1648 (O_1648,N_49709,N_49876);
and UO_1649 (O_1649,N_49558,N_49774);
xor UO_1650 (O_1650,N_49548,N_49764);
xnor UO_1651 (O_1651,N_49521,N_49787);
or UO_1652 (O_1652,N_49728,N_49716);
and UO_1653 (O_1653,N_49582,N_49798);
and UO_1654 (O_1654,N_49751,N_49942);
and UO_1655 (O_1655,N_49728,N_49611);
nor UO_1656 (O_1656,N_49863,N_49817);
or UO_1657 (O_1657,N_49980,N_49810);
nand UO_1658 (O_1658,N_49864,N_49813);
and UO_1659 (O_1659,N_49758,N_49805);
or UO_1660 (O_1660,N_49758,N_49864);
nor UO_1661 (O_1661,N_49748,N_49689);
or UO_1662 (O_1662,N_49674,N_49633);
nor UO_1663 (O_1663,N_49669,N_49575);
nand UO_1664 (O_1664,N_49570,N_49755);
and UO_1665 (O_1665,N_49516,N_49942);
nor UO_1666 (O_1666,N_49769,N_49999);
xnor UO_1667 (O_1667,N_49800,N_49750);
nand UO_1668 (O_1668,N_49621,N_49965);
or UO_1669 (O_1669,N_49603,N_49886);
and UO_1670 (O_1670,N_49982,N_49927);
or UO_1671 (O_1671,N_49948,N_49783);
xor UO_1672 (O_1672,N_49578,N_49982);
nor UO_1673 (O_1673,N_49738,N_49994);
nand UO_1674 (O_1674,N_49564,N_49963);
xnor UO_1675 (O_1675,N_49771,N_49703);
nand UO_1676 (O_1676,N_49573,N_49769);
or UO_1677 (O_1677,N_49645,N_49609);
nor UO_1678 (O_1678,N_49919,N_49709);
nand UO_1679 (O_1679,N_49529,N_49635);
or UO_1680 (O_1680,N_49530,N_49660);
and UO_1681 (O_1681,N_49959,N_49509);
and UO_1682 (O_1682,N_49805,N_49959);
nor UO_1683 (O_1683,N_49787,N_49539);
xor UO_1684 (O_1684,N_49891,N_49977);
nor UO_1685 (O_1685,N_49640,N_49612);
or UO_1686 (O_1686,N_49541,N_49563);
xor UO_1687 (O_1687,N_49991,N_49765);
or UO_1688 (O_1688,N_49734,N_49574);
and UO_1689 (O_1689,N_49680,N_49838);
xnor UO_1690 (O_1690,N_49764,N_49926);
and UO_1691 (O_1691,N_49710,N_49580);
xnor UO_1692 (O_1692,N_49872,N_49633);
xor UO_1693 (O_1693,N_49889,N_49508);
or UO_1694 (O_1694,N_49562,N_49550);
or UO_1695 (O_1695,N_49719,N_49669);
or UO_1696 (O_1696,N_49971,N_49827);
xnor UO_1697 (O_1697,N_49763,N_49748);
xnor UO_1698 (O_1698,N_49796,N_49934);
nor UO_1699 (O_1699,N_49677,N_49920);
nor UO_1700 (O_1700,N_49675,N_49798);
or UO_1701 (O_1701,N_49575,N_49654);
xor UO_1702 (O_1702,N_49537,N_49531);
xor UO_1703 (O_1703,N_49990,N_49707);
or UO_1704 (O_1704,N_49964,N_49527);
xnor UO_1705 (O_1705,N_49691,N_49866);
nand UO_1706 (O_1706,N_49751,N_49668);
and UO_1707 (O_1707,N_49987,N_49800);
xor UO_1708 (O_1708,N_49886,N_49739);
nor UO_1709 (O_1709,N_49691,N_49791);
nor UO_1710 (O_1710,N_49653,N_49647);
nand UO_1711 (O_1711,N_49594,N_49998);
xnor UO_1712 (O_1712,N_49943,N_49836);
nor UO_1713 (O_1713,N_49623,N_49566);
nor UO_1714 (O_1714,N_49710,N_49688);
and UO_1715 (O_1715,N_49648,N_49512);
nand UO_1716 (O_1716,N_49789,N_49765);
and UO_1717 (O_1717,N_49818,N_49561);
nor UO_1718 (O_1718,N_49550,N_49740);
nand UO_1719 (O_1719,N_49925,N_49564);
and UO_1720 (O_1720,N_49702,N_49601);
nor UO_1721 (O_1721,N_49578,N_49507);
nand UO_1722 (O_1722,N_49661,N_49778);
xnor UO_1723 (O_1723,N_49536,N_49764);
xnor UO_1724 (O_1724,N_49612,N_49762);
nand UO_1725 (O_1725,N_49768,N_49830);
nand UO_1726 (O_1726,N_49938,N_49511);
xnor UO_1727 (O_1727,N_49941,N_49502);
nand UO_1728 (O_1728,N_49806,N_49701);
xnor UO_1729 (O_1729,N_49881,N_49552);
or UO_1730 (O_1730,N_49911,N_49753);
xnor UO_1731 (O_1731,N_49791,N_49515);
xnor UO_1732 (O_1732,N_49567,N_49590);
nand UO_1733 (O_1733,N_49504,N_49740);
or UO_1734 (O_1734,N_49734,N_49545);
or UO_1735 (O_1735,N_49849,N_49551);
or UO_1736 (O_1736,N_49541,N_49966);
and UO_1737 (O_1737,N_49962,N_49909);
or UO_1738 (O_1738,N_49807,N_49583);
nor UO_1739 (O_1739,N_49597,N_49709);
nand UO_1740 (O_1740,N_49956,N_49591);
nor UO_1741 (O_1741,N_49615,N_49859);
nor UO_1742 (O_1742,N_49600,N_49606);
nand UO_1743 (O_1743,N_49794,N_49810);
xnor UO_1744 (O_1744,N_49907,N_49677);
nand UO_1745 (O_1745,N_49797,N_49630);
nand UO_1746 (O_1746,N_49993,N_49533);
nand UO_1747 (O_1747,N_49881,N_49531);
xnor UO_1748 (O_1748,N_49782,N_49892);
nor UO_1749 (O_1749,N_49805,N_49719);
xor UO_1750 (O_1750,N_49627,N_49831);
nor UO_1751 (O_1751,N_49847,N_49758);
xor UO_1752 (O_1752,N_49931,N_49937);
or UO_1753 (O_1753,N_49832,N_49550);
and UO_1754 (O_1754,N_49887,N_49888);
xor UO_1755 (O_1755,N_49809,N_49690);
xor UO_1756 (O_1756,N_49712,N_49973);
and UO_1757 (O_1757,N_49699,N_49615);
nor UO_1758 (O_1758,N_49576,N_49509);
nor UO_1759 (O_1759,N_49650,N_49823);
and UO_1760 (O_1760,N_49586,N_49957);
xnor UO_1761 (O_1761,N_49839,N_49962);
and UO_1762 (O_1762,N_49609,N_49830);
nand UO_1763 (O_1763,N_49911,N_49870);
nor UO_1764 (O_1764,N_49595,N_49639);
nor UO_1765 (O_1765,N_49676,N_49863);
nor UO_1766 (O_1766,N_49918,N_49849);
xor UO_1767 (O_1767,N_49787,N_49841);
xor UO_1768 (O_1768,N_49633,N_49620);
and UO_1769 (O_1769,N_49524,N_49537);
or UO_1770 (O_1770,N_49723,N_49501);
nor UO_1771 (O_1771,N_49651,N_49818);
or UO_1772 (O_1772,N_49952,N_49763);
xnor UO_1773 (O_1773,N_49508,N_49570);
xnor UO_1774 (O_1774,N_49917,N_49939);
nand UO_1775 (O_1775,N_49592,N_49885);
and UO_1776 (O_1776,N_49854,N_49923);
and UO_1777 (O_1777,N_49991,N_49532);
nand UO_1778 (O_1778,N_49851,N_49512);
and UO_1779 (O_1779,N_49652,N_49779);
and UO_1780 (O_1780,N_49500,N_49696);
xnor UO_1781 (O_1781,N_49695,N_49968);
or UO_1782 (O_1782,N_49925,N_49524);
nor UO_1783 (O_1783,N_49695,N_49712);
nor UO_1784 (O_1784,N_49631,N_49544);
nor UO_1785 (O_1785,N_49647,N_49587);
nand UO_1786 (O_1786,N_49506,N_49523);
and UO_1787 (O_1787,N_49953,N_49556);
and UO_1788 (O_1788,N_49930,N_49817);
xor UO_1789 (O_1789,N_49693,N_49709);
xor UO_1790 (O_1790,N_49894,N_49884);
or UO_1791 (O_1791,N_49664,N_49638);
and UO_1792 (O_1792,N_49513,N_49866);
nor UO_1793 (O_1793,N_49641,N_49663);
nand UO_1794 (O_1794,N_49822,N_49633);
or UO_1795 (O_1795,N_49502,N_49961);
nand UO_1796 (O_1796,N_49824,N_49915);
and UO_1797 (O_1797,N_49808,N_49729);
and UO_1798 (O_1798,N_49676,N_49845);
xor UO_1799 (O_1799,N_49688,N_49628);
xnor UO_1800 (O_1800,N_49716,N_49574);
or UO_1801 (O_1801,N_49927,N_49605);
xor UO_1802 (O_1802,N_49787,N_49600);
or UO_1803 (O_1803,N_49951,N_49908);
nand UO_1804 (O_1804,N_49711,N_49926);
nand UO_1805 (O_1805,N_49929,N_49916);
nor UO_1806 (O_1806,N_49668,N_49782);
nor UO_1807 (O_1807,N_49780,N_49972);
nand UO_1808 (O_1808,N_49615,N_49538);
or UO_1809 (O_1809,N_49608,N_49929);
xor UO_1810 (O_1810,N_49620,N_49713);
nor UO_1811 (O_1811,N_49546,N_49800);
xor UO_1812 (O_1812,N_49890,N_49660);
nand UO_1813 (O_1813,N_49892,N_49627);
nor UO_1814 (O_1814,N_49771,N_49875);
nor UO_1815 (O_1815,N_49695,N_49982);
or UO_1816 (O_1816,N_49509,N_49760);
nand UO_1817 (O_1817,N_49781,N_49527);
and UO_1818 (O_1818,N_49716,N_49589);
and UO_1819 (O_1819,N_49652,N_49979);
and UO_1820 (O_1820,N_49775,N_49948);
nand UO_1821 (O_1821,N_49580,N_49915);
and UO_1822 (O_1822,N_49726,N_49567);
and UO_1823 (O_1823,N_49784,N_49810);
and UO_1824 (O_1824,N_49779,N_49858);
and UO_1825 (O_1825,N_49630,N_49645);
or UO_1826 (O_1826,N_49938,N_49572);
xnor UO_1827 (O_1827,N_49956,N_49512);
nand UO_1828 (O_1828,N_49520,N_49918);
xnor UO_1829 (O_1829,N_49704,N_49998);
or UO_1830 (O_1830,N_49828,N_49835);
nor UO_1831 (O_1831,N_49977,N_49710);
and UO_1832 (O_1832,N_49775,N_49919);
nor UO_1833 (O_1833,N_49618,N_49527);
or UO_1834 (O_1834,N_49742,N_49788);
nor UO_1835 (O_1835,N_49557,N_49980);
nand UO_1836 (O_1836,N_49754,N_49838);
nor UO_1837 (O_1837,N_49511,N_49854);
xor UO_1838 (O_1838,N_49853,N_49945);
and UO_1839 (O_1839,N_49640,N_49768);
nor UO_1840 (O_1840,N_49985,N_49524);
nor UO_1841 (O_1841,N_49880,N_49888);
xnor UO_1842 (O_1842,N_49577,N_49854);
xnor UO_1843 (O_1843,N_49620,N_49838);
and UO_1844 (O_1844,N_49847,N_49871);
nand UO_1845 (O_1845,N_49846,N_49988);
nand UO_1846 (O_1846,N_49551,N_49971);
nand UO_1847 (O_1847,N_49721,N_49669);
xnor UO_1848 (O_1848,N_49659,N_49636);
and UO_1849 (O_1849,N_49555,N_49720);
and UO_1850 (O_1850,N_49666,N_49731);
and UO_1851 (O_1851,N_49836,N_49805);
or UO_1852 (O_1852,N_49651,N_49769);
or UO_1853 (O_1853,N_49737,N_49988);
nor UO_1854 (O_1854,N_49763,N_49889);
nand UO_1855 (O_1855,N_49500,N_49946);
or UO_1856 (O_1856,N_49595,N_49750);
or UO_1857 (O_1857,N_49815,N_49993);
nor UO_1858 (O_1858,N_49918,N_49574);
nand UO_1859 (O_1859,N_49548,N_49781);
xor UO_1860 (O_1860,N_49589,N_49846);
nor UO_1861 (O_1861,N_49585,N_49640);
nand UO_1862 (O_1862,N_49939,N_49816);
or UO_1863 (O_1863,N_49866,N_49899);
nor UO_1864 (O_1864,N_49542,N_49840);
nor UO_1865 (O_1865,N_49738,N_49798);
and UO_1866 (O_1866,N_49991,N_49889);
nor UO_1867 (O_1867,N_49524,N_49845);
xnor UO_1868 (O_1868,N_49679,N_49503);
or UO_1869 (O_1869,N_49623,N_49916);
nand UO_1870 (O_1870,N_49827,N_49714);
or UO_1871 (O_1871,N_49502,N_49642);
xor UO_1872 (O_1872,N_49542,N_49768);
xnor UO_1873 (O_1873,N_49764,N_49754);
nand UO_1874 (O_1874,N_49882,N_49665);
and UO_1875 (O_1875,N_49867,N_49894);
xor UO_1876 (O_1876,N_49899,N_49630);
xnor UO_1877 (O_1877,N_49850,N_49729);
xor UO_1878 (O_1878,N_49628,N_49754);
nor UO_1879 (O_1879,N_49713,N_49762);
or UO_1880 (O_1880,N_49837,N_49713);
nand UO_1881 (O_1881,N_49987,N_49733);
or UO_1882 (O_1882,N_49547,N_49951);
xnor UO_1883 (O_1883,N_49784,N_49711);
nand UO_1884 (O_1884,N_49924,N_49991);
and UO_1885 (O_1885,N_49512,N_49934);
or UO_1886 (O_1886,N_49594,N_49512);
xor UO_1887 (O_1887,N_49840,N_49876);
nand UO_1888 (O_1888,N_49641,N_49787);
nand UO_1889 (O_1889,N_49510,N_49889);
and UO_1890 (O_1890,N_49902,N_49865);
xor UO_1891 (O_1891,N_49760,N_49731);
nand UO_1892 (O_1892,N_49640,N_49632);
nand UO_1893 (O_1893,N_49961,N_49693);
nand UO_1894 (O_1894,N_49955,N_49667);
xor UO_1895 (O_1895,N_49738,N_49815);
nand UO_1896 (O_1896,N_49630,N_49779);
nor UO_1897 (O_1897,N_49885,N_49746);
and UO_1898 (O_1898,N_49639,N_49696);
nand UO_1899 (O_1899,N_49783,N_49621);
nor UO_1900 (O_1900,N_49961,N_49649);
nand UO_1901 (O_1901,N_49923,N_49879);
or UO_1902 (O_1902,N_49579,N_49667);
xnor UO_1903 (O_1903,N_49691,N_49653);
nor UO_1904 (O_1904,N_49722,N_49520);
nand UO_1905 (O_1905,N_49850,N_49706);
and UO_1906 (O_1906,N_49637,N_49857);
nor UO_1907 (O_1907,N_49940,N_49919);
nor UO_1908 (O_1908,N_49508,N_49574);
nand UO_1909 (O_1909,N_49725,N_49726);
and UO_1910 (O_1910,N_49915,N_49918);
nor UO_1911 (O_1911,N_49980,N_49845);
nand UO_1912 (O_1912,N_49543,N_49733);
nor UO_1913 (O_1913,N_49606,N_49597);
or UO_1914 (O_1914,N_49718,N_49686);
or UO_1915 (O_1915,N_49852,N_49751);
nor UO_1916 (O_1916,N_49736,N_49588);
xnor UO_1917 (O_1917,N_49880,N_49929);
or UO_1918 (O_1918,N_49546,N_49811);
xor UO_1919 (O_1919,N_49850,N_49921);
nand UO_1920 (O_1920,N_49872,N_49686);
and UO_1921 (O_1921,N_49822,N_49787);
or UO_1922 (O_1922,N_49866,N_49870);
xor UO_1923 (O_1923,N_49618,N_49686);
nand UO_1924 (O_1924,N_49547,N_49906);
and UO_1925 (O_1925,N_49629,N_49530);
and UO_1926 (O_1926,N_49600,N_49636);
nor UO_1927 (O_1927,N_49984,N_49593);
nand UO_1928 (O_1928,N_49855,N_49581);
xnor UO_1929 (O_1929,N_49814,N_49627);
or UO_1930 (O_1930,N_49764,N_49974);
nor UO_1931 (O_1931,N_49679,N_49723);
xor UO_1932 (O_1932,N_49914,N_49936);
nand UO_1933 (O_1933,N_49704,N_49961);
and UO_1934 (O_1934,N_49821,N_49789);
nor UO_1935 (O_1935,N_49887,N_49585);
xor UO_1936 (O_1936,N_49729,N_49818);
nand UO_1937 (O_1937,N_49557,N_49951);
xor UO_1938 (O_1938,N_49930,N_49555);
or UO_1939 (O_1939,N_49581,N_49644);
nor UO_1940 (O_1940,N_49994,N_49732);
nand UO_1941 (O_1941,N_49639,N_49998);
or UO_1942 (O_1942,N_49943,N_49979);
nor UO_1943 (O_1943,N_49840,N_49664);
nor UO_1944 (O_1944,N_49555,N_49964);
nor UO_1945 (O_1945,N_49869,N_49997);
nand UO_1946 (O_1946,N_49866,N_49534);
nand UO_1947 (O_1947,N_49803,N_49831);
xnor UO_1948 (O_1948,N_49988,N_49832);
nand UO_1949 (O_1949,N_49813,N_49629);
nand UO_1950 (O_1950,N_49981,N_49897);
or UO_1951 (O_1951,N_49606,N_49979);
or UO_1952 (O_1952,N_49530,N_49596);
nand UO_1953 (O_1953,N_49979,N_49526);
nand UO_1954 (O_1954,N_49815,N_49565);
nand UO_1955 (O_1955,N_49534,N_49718);
xor UO_1956 (O_1956,N_49850,N_49623);
xor UO_1957 (O_1957,N_49574,N_49933);
xnor UO_1958 (O_1958,N_49767,N_49505);
nor UO_1959 (O_1959,N_49678,N_49802);
nand UO_1960 (O_1960,N_49870,N_49655);
or UO_1961 (O_1961,N_49940,N_49830);
nor UO_1962 (O_1962,N_49989,N_49644);
nand UO_1963 (O_1963,N_49825,N_49665);
or UO_1964 (O_1964,N_49981,N_49608);
nand UO_1965 (O_1965,N_49782,N_49998);
and UO_1966 (O_1966,N_49800,N_49596);
or UO_1967 (O_1967,N_49772,N_49574);
nor UO_1968 (O_1968,N_49764,N_49725);
xor UO_1969 (O_1969,N_49859,N_49947);
and UO_1970 (O_1970,N_49790,N_49760);
xnor UO_1971 (O_1971,N_49963,N_49590);
and UO_1972 (O_1972,N_49883,N_49727);
xnor UO_1973 (O_1973,N_49795,N_49807);
nand UO_1974 (O_1974,N_49983,N_49628);
nand UO_1975 (O_1975,N_49995,N_49649);
nor UO_1976 (O_1976,N_49967,N_49993);
nor UO_1977 (O_1977,N_49877,N_49581);
and UO_1978 (O_1978,N_49632,N_49789);
and UO_1979 (O_1979,N_49560,N_49917);
and UO_1980 (O_1980,N_49650,N_49603);
xor UO_1981 (O_1981,N_49711,N_49566);
nand UO_1982 (O_1982,N_49588,N_49984);
xor UO_1983 (O_1983,N_49656,N_49530);
and UO_1984 (O_1984,N_49978,N_49726);
nand UO_1985 (O_1985,N_49545,N_49913);
or UO_1986 (O_1986,N_49649,N_49796);
nor UO_1987 (O_1987,N_49889,N_49934);
or UO_1988 (O_1988,N_49709,N_49848);
xnor UO_1989 (O_1989,N_49765,N_49971);
and UO_1990 (O_1990,N_49675,N_49600);
or UO_1991 (O_1991,N_49585,N_49955);
nand UO_1992 (O_1992,N_49506,N_49640);
xor UO_1993 (O_1993,N_49750,N_49589);
nand UO_1994 (O_1994,N_49813,N_49660);
nor UO_1995 (O_1995,N_49726,N_49768);
and UO_1996 (O_1996,N_49849,N_49766);
nand UO_1997 (O_1997,N_49902,N_49747);
nor UO_1998 (O_1998,N_49511,N_49649);
nand UO_1999 (O_1999,N_49625,N_49761);
nand UO_2000 (O_2000,N_49943,N_49638);
xor UO_2001 (O_2001,N_49720,N_49756);
nand UO_2002 (O_2002,N_49979,N_49990);
nor UO_2003 (O_2003,N_49892,N_49839);
or UO_2004 (O_2004,N_49854,N_49729);
or UO_2005 (O_2005,N_49927,N_49677);
nand UO_2006 (O_2006,N_49598,N_49584);
xnor UO_2007 (O_2007,N_49994,N_49948);
nor UO_2008 (O_2008,N_49979,N_49548);
or UO_2009 (O_2009,N_49638,N_49689);
and UO_2010 (O_2010,N_49669,N_49991);
or UO_2011 (O_2011,N_49693,N_49613);
or UO_2012 (O_2012,N_49529,N_49584);
xor UO_2013 (O_2013,N_49675,N_49654);
or UO_2014 (O_2014,N_49612,N_49937);
or UO_2015 (O_2015,N_49893,N_49734);
nor UO_2016 (O_2016,N_49728,N_49959);
and UO_2017 (O_2017,N_49721,N_49747);
xor UO_2018 (O_2018,N_49945,N_49882);
and UO_2019 (O_2019,N_49504,N_49533);
and UO_2020 (O_2020,N_49881,N_49926);
or UO_2021 (O_2021,N_49822,N_49871);
nor UO_2022 (O_2022,N_49650,N_49731);
nor UO_2023 (O_2023,N_49963,N_49893);
xor UO_2024 (O_2024,N_49732,N_49648);
xnor UO_2025 (O_2025,N_49526,N_49729);
xor UO_2026 (O_2026,N_49502,N_49927);
xnor UO_2027 (O_2027,N_49917,N_49935);
or UO_2028 (O_2028,N_49953,N_49547);
nand UO_2029 (O_2029,N_49747,N_49872);
and UO_2030 (O_2030,N_49852,N_49681);
nor UO_2031 (O_2031,N_49558,N_49603);
and UO_2032 (O_2032,N_49896,N_49854);
xor UO_2033 (O_2033,N_49992,N_49516);
xor UO_2034 (O_2034,N_49684,N_49847);
or UO_2035 (O_2035,N_49513,N_49855);
nor UO_2036 (O_2036,N_49619,N_49669);
nand UO_2037 (O_2037,N_49850,N_49570);
xnor UO_2038 (O_2038,N_49957,N_49554);
or UO_2039 (O_2039,N_49514,N_49662);
nor UO_2040 (O_2040,N_49623,N_49908);
and UO_2041 (O_2041,N_49658,N_49989);
or UO_2042 (O_2042,N_49866,N_49948);
and UO_2043 (O_2043,N_49530,N_49848);
nand UO_2044 (O_2044,N_49864,N_49530);
and UO_2045 (O_2045,N_49578,N_49545);
or UO_2046 (O_2046,N_49918,N_49861);
or UO_2047 (O_2047,N_49614,N_49796);
xnor UO_2048 (O_2048,N_49809,N_49773);
nor UO_2049 (O_2049,N_49826,N_49831);
xnor UO_2050 (O_2050,N_49629,N_49771);
and UO_2051 (O_2051,N_49958,N_49826);
nor UO_2052 (O_2052,N_49799,N_49519);
nor UO_2053 (O_2053,N_49621,N_49743);
and UO_2054 (O_2054,N_49950,N_49521);
nand UO_2055 (O_2055,N_49788,N_49605);
and UO_2056 (O_2056,N_49742,N_49556);
or UO_2057 (O_2057,N_49704,N_49801);
or UO_2058 (O_2058,N_49726,N_49782);
nor UO_2059 (O_2059,N_49788,N_49957);
nand UO_2060 (O_2060,N_49919,N_49629);
and UO_2061 (O_2061,N_49723,N_49984);
xor UO_2062 (O_2062,N_49673,N_49864);
nor UO_2063 (O_2063,N_49902,N_49786);
and UO_2064 (O_2064,N_49659,N_49757);
or UO_2065 (O_2065,N_49779,N_49554);
xor UO_2066 (O_2066,N_49779,N_49615);
nand UO_2067 (O_2067,N_49820,N_49861);
nor UO_2068 (O_2068,N_49815,N_49928);
nand UO_2069 (O_2069,N_49507,N_49986);
and UO_2070 (O_2070,N_49709,N_49659);
nor UO_2071 (O_2071,N_49876,N_49745);
nand UO_2072 (O_2072,N_49618,N_49529);
or UO_2073 (O_2073,N_49522,N_49715);
nor UO_2074 (O_2074,N_49603,N_49863);
xor UO_2075 (O_2075,N_49790,N_49935);
nand UO_2076 (O_2076,N_49599,N_49880);
nand UO_2077 (O_2077,N_49542,N_49552);
nand UO_2078 (O_2078,N_49544,N_49968);
and UO_2079 (O_2079,N_49659,N_49516);
nor UO_2080 (O_2080,N_49847,N_49737);
or UO_2081 (O_2081,N_49626,N_49751);
or UO_2082 (O_2082,N_49768,N_49808);
xor UO_2083 (O_2083,N_49533,N_49840);
or UO_2084 (O_2084,N_49803,N_49637);
xor UO_2085 (O_2085,N_49943,N_49887);
nand UO_2086 (O_2086,N_49821,N_49986);
and UO_2087 (O_2087,N_49662,N_49972);
nor UO_2088 (O_2088,N_49661,N_49589);
nor UO_2089 (O_2089,N_49933,N_49818);
or UO_2090 (O_2090,N_49597,N_49804);
nand UO_2091 (O_2091,N_49820,N_49928);
and UO_2092 (O_2092,N_49927,N_49845);
nand UO_2093 (O_2093,N_49945,N_49680);
xor UO_2094 (O_2094,N_49671,N_49983);
and UO_2095 (O_2095,N_49852,N_49665);
or UO_2096 (O_2096,N_49647,N_49924);
nor UO_2097 (O_2097,N_49561,N_49706);
nand UO_2098 (O_2098,N_49785,N_49701);
xor UO_2099 (O_2099,N_49758,N_49961);
or UO_2100 (O_2100,N_49577,N_49828);
nand UO_2101 (O_2101,N_49582,N_49891);
nand UO_2102 (O_2102,N_49642,N_49568);
and UO_2103 (O_2103,N_49966,N_49943);
and UO_2104 (O_2104,N_49972,N_49733);
nor UO_2105 (O_2105,N_49937,N_49573);
nor UO_2106 (O_2106,N_49506,N_49717);
and UO_2107 (O_2107,N_49949,N_49913);
or UO_2108 (O_2108,N_49740,N_49866);
xor UO_2109 (O_2109,N_49856,N_49985);
and UO_2110 (O_2110,N_49855,N_49897);
or UO_2111 (O_2111,N_49986,N_49609);
and UO_2112 (O_2112,N_49711,N_49983);
nor UO_2113 (O_2113,N_49635,N_49761);
and UO_2114 (O_2114,N_49943,N_49717);
and UO_2115 (O_2115,N_49975,N_49859);
nor UO_2116 (O_2116,N_49634,N_49828);
nor UO_2117 (O_2117,N_49822,N_49707);
nand UO_2118 (O_2118,N_49978,N_49948);
and UO_2119 (O_2119,N_49944,N_49961);
xor UO_2120 (O_2120,N_49605,N_49941);
or UO_2121 (O_2121,N_49695,N_49655);
or UO_2122 (O_2122,N_49691,N_49803);
xnor UO_2123 (O_2123,N_49962,N_49676);
or UO_2124 (O_2124,N_49573,N_49824);
nor UO_2125 (O_2125,N_49963,N_49735);
nor UO_2126 (O_2126,N_49675,N_49690);
nand UO_2127 (O_2127,N_49757,N_49542);
and UO_2128 (O_2128,N_49679,N_49995);
and UO_2129 (O_2129,N_49746,N_49657);
nand UO_2130 (O_2130,N_49736,N_49657);
nor UO_2131 (O_2131,N_49729,N_49542);
xnor UO_2132 (O_2132,N_49674,N_49816);
or UO_2133 (O_2133,N_49925,N_49594);
xor UO_2134 (O_2134,N_49747,N_49785);
xnor UO_2135 (O_2135,N_49634,N_49715);
nand UO_2136 (O_2136,N_49606,N_49853);
or UO_2137 (O_2137,N_49824,N_49973);
nor UO_2138 (O_2138,N_49684,N_49672);
or UO_2139 (O_2139,N_49521,N_49634);
or UO_2140 (O_2140,N_49529,N_49961);
or UO_2141 (O_2141,N_49983,N_49731);
nand UO_2142 (O_2142,N_49685,N_49732);
or UO_2143 (O_2143,N_49936,N_49925);
nand UO_2144 (O_2144,N_49860,N_49632);
nor UO_2145 (O_2145,N_49890,N_49739);
nor UO_2146 (O_2146,N_49941,N_49514);
or UO_2147 (O_2147,N_49912,N_49926);
nand UO_2148 (O_2148,N_49716,N_49519);
nor UO_2149 (O_2149,N_49755,N_49938);
or UO_2150 (O_2150,N_49929,N_49582);
and UO_2151 (O_2151,N_49561,N_49862);
xor UO_2152 (O_2152,N_49634,N_49872);
nor UO_2153 (O_2153,N_49901,N_49584);
nand UO_2154 (O_2154,N_49538,N_49786);
and UO_2155 (O_2155,N_49828,N_49697);
nand UO_2156 (O_2156,N_49689,N_49551);
nand UO_2157 (O_2157,N_49910,N_49588);
nor UO_2158 (O_2158,N_49539,N_49758);
xnor UO_2159 (O_2159,N_49699,N_49686);
and UO_2160 (O_2160,N_49520,N_49718);
and UO_2161 (O_2161,N_49870,N_49855);
xor UO_2162 (O_2162,N_49730,N_49545);
nor UO_2163 (O_2163,N_49751,N_49984);
or UO_2164 (O_2164,N_49526,N_49972);
xnor UO_2165 (O_2165,N_49544,N_49716);
xnor UO_2166 (O_2166,N_49880,N_49500);
and UO_2167 (O_2167,N_49563,N_49687);
nor UO_2168 (O_2168,N_49755,N_49743);
nor UO_2169 (O_2169,N_49864,N_49932);
or UO_2170 (O_2170,N_49551,N_49807);
and UO_2171 (O_2171,N_49939,N_49575);
nor UO_2172 (O_2172,N_49900,N_49705);
nand UO_2173 (O_2173,N_49869,N_49807);
nand UO_2174 (O_2174,N_49718,N_49727);
xnor UO_2175 (O_2175,N_49554,N_49860);
nor UO_2176 (O_2176,N_49722,N_49599);
nand UO_2177 (O_2177,N_49962,N_49939);
and UO_2178 (O_2178,N_49776,N_49587);
xor UO_2179 (O_2179,N_49621,N_49777);
nor UO_2180 (O_2180,N_49952,N_49521);
nand UO_2181 (O_2181,N_49532,N_49520);
or UO_2182 (O_2182,N_49569,N_49837);
nand UO_2183 (O_2183,N_49649,N_49992);
or UO_2184 (O_2184,N_49924,N_49567);
or UO_2185 (O_2185,N_49523,N_49871);
nand UO_2186 (O_2186,N_49865,N_49815);
nand UO_2187 (O_2187,N_49851,N_49741);
xnor UO_2188 (O_2188,N_49748,N_49975);
or UO_2189 (O_2189,N_49627,N_49816);
xnor UO_2190 (O_2190,N_49832,N_49755);
xor UO_2191 (O_2191,N_49788,N_49961);
nor UO_2192 (O_2192,N_49833,N_49583);
or UO_2193 (O_2193,N_49922,N_49783);
or UO_2194 (O_2194,N_49587,N_49561);
xor UO_2195 (O_2195,N_49564,N_49893);
nand UO_2196 (O_2196,N_49530,N_49842);
nor UO_2197 (O_2197,N_49848,N_49830);
or UO_2198 (O_2198,N_49809,N_49738);
nor UO_2199 (O_2199,N_49859,N_49846);
xor UO_2200 (O_2200,N_49997,N_49800);
nand UO_2201 (O_2201,N_49915,N_49652);
or UO_2202 (O_2202,N_49698,N_49598);
nand UO_2203 (O_2203,N_49933,N_49599);
nor UO_2204 (O_2204,N_49668,N_49912);
or UO_2205 (O_2205,N_49866,N_49614);
nand UO_2206 (O_2206,N_49687,N_49972);
or UO_2207 (O_2207,N_49972,N_49851);
nor UO_2208 (O_2208,N_49600,N_49628);
xnor UO_2209 (O_2209,N_49895,N_49863);
and UO_2210 (O_2210,N_49764,N_49769);
and UO_2211 (O_2211,N_49737,N_49927);
xnor UO_2212 (O_2212,N_49696,N_49593);
nor UO_2213 (O_2213,N_49943,N_49505);
xor UO_2214 (O_2214,N_49575,N_49871);
or UO_2215 (O_2215,N_49709,N_49534);
nor UO_2216 (O_2216,N_49831,N_49666);
nor UO_2217 (O_2217,N_49845,N_49745);
or UO_2218 (O_2218,N_49589,N_49523);
or UO_2219 (O_2219,N_49953,N_49580);
xnor UO_2220 (O_2220,N_49976,N_49775);
nand UO_2221 (O_2221,N_49648,N_49723);
nor UO_2222 (O_2222,N_49791,N_49921);
and UO_2223 (O_2223,N_49803,N_49798);
nand UO_2224 (O_2224,N_49510,N_49936);
or UO_2225 (O_2225,N_49914,N_49708);
and UO_2226 (O_2226,N_49514,N_49543);
nor UO_2227 (O_2227,N_49896,N_49737);
or UO_2228 (O_2228,N_49620,N_49866);
nor UO_2229 (O_2229,N_49851,N_49540);
nor UO_2230 (O_2230,N_49535,N_49934);
nand UO_2231 (O_2231,N_49792,N_49666);
xor UO_2232 (O_2232,N_49713,N_49524);
and UO_2233 (O_2233,N_49823,N_49778);
nand UO_2234 (O_2234,N_49845,N_49797);
and UO_2235 (O_2235,N_49750,N_49501);
and UO_2236 (O_2236,N_49580,N_49777);
nand UO_2237 (O_2237,N_49961,N_49524);
and UO_2238 (O_2238,N_49690,N_49758);
and UO_2239 (O_2239,N_49602,N_49803);
or UO_2240 (O_2240,N_49778,N_49585);
or UO_2241 (O_2241,N_49860,N_49528);
or UO_2242 (O_2242,N_49592,N_49577);
and UO_2243 (O_2243,N_49778,N_49898);
or UO_2244 (O_2244,N_49729,N_49633);
nand UO_2245 (O_2245,N_49502,N_49708);
nand UO_2246 (O_2246,N_49586,N_49554);
nor UO_2247 (O_2247,N_49882,N_49977);
and UO_2248 (O_2248,N_49586,N_49693);
and UO_2249 (O_2249,N_49835,N_49787);
or UO_2250 (O_2250,N_49788,N_49510);
nor UO_2251 (O_2251,N_49786,N_49731);
xor UO_2252 (O_2252,N_49509,N_49644);
nor UO_2253 (O_2253,N_49814,N_49621);
nand UO_2254 (O_2254,N_49692,N_49903);
or UO_2255 (O_2255,N_49753,N_49914);
nand UO_2256 (O_2256,N_49518,N_49638);
xnor UO_2257 (O_2257,N_49645,N_49967);
and UO_2258 (O_2258,N_49989,N_49565);
and UO_2259 (O_2259,N_49771,N_49588);
xnor UO_2260 (O_2260,N_49666,N_49790);
and UO_2261 (O_2261,N_49552,N_49782);
nand UO_2262 (O_2262,N_49899,N_49548);
nand UO_2263 (O_2263,N_49985,N_49939);
nor UO_2264 (O_2264,N_49871,N_49800);
and UO_2265 (O_2265,N_49998,N_49817);
or UO_2266 (O_2266,N_49538,N_49776);
or UO_2267 (O_2267,N_49825,N_49681);
xor UO_2268 (O_2268,N_49834,N_49777);
and UO_2269 (O_2269,N_49750,N_49671);
nand UO_2270 (O_2270,N_49571,N_49549);
or UO_2271 (O_2271,N_49719,N_49950);
nor UO_2272 (O_2272,N_49572,N_49574);
or UO_2273 (O_2273,N_49502,N_49958);
nor UO_2274 (O_2274,N_49953,N_49718);
nand UO_2275 (O_2275,N_49519,N_49666);
nor UO_2276 (O_2276,N_49989,N_49522);
nor UO_2277 (O_2277,N_49768,N_49968);
nand UO_2278 (O_2278,N_49746,N_49713);
xnor UO_2279 (O_2279,N_49917,N_49768);
nor UO_2280 (O_2280,N_49714,N_49572);
and UO_2281 (O_2281,N_49932,N_49769);
nand UO_2282 (O_2282,N_49824,N_49585);
xor UO_2283 (O_2283,N_49818,N_49816);
xnor UO_2284 (O_2284,N_49736,N_49832);
xor UO_2285 (O_2285,N_49714,N_49807);
xor UO_2286 (O_2286,N_49606,N_49898);
nand UO_2287 (O_2287,N_49764,N_49815);
nand UO_2288 (O_2288,N_49742,N_49595);
nand UO_2289 (O_2289,N_49875,N_49861);
and UO_2290 (O_2290,N_49568,N_49590);
and UO_2291 (O_2291,N_49974,N_49553);
nor UO_2292 (O_2292,N_49971,N_49741);
xor UO_2293 (O_2293,N_49850,N_49705);
nand UO_2294 (O_2294,N_49969,N_49960);
nand UO_2295 (O_2295,N_49755,N_49635);
nor UO_2296 (O_2296,N_49611,N_49920);
nand UO_2297 (O_2297,N_49572,N_49660);
nor UO_2298 (O_2298,N_49719,N_49774);
and UO_2299 (O_2299,N_49648,N_49650);
nand UO_2300 (O_2300,N_49962,N_49888);
nand UO_2301 (O_2301,N_49603,N_49713);
nor UO_2302 (O_2302,N_49935,N_49671);
or UO_2303 (O_2303,N_49543,N_49924);
xnor UO_2304 (O_2304,N_49830,N_49542);
and UO_2305 (O_2305,N_49523,N_49528);
xor UO_2306 (O_2306,N_49970,N_49942);
nand UO_2307 (O_2307,N_49629,N_49723);
xnor UO_2308 (O_2308,N_49521,N_49621);
nand UO_2309 (O_2309,N_49545,N_49722);
or UO_2310 (O_2310,N_49661,N_49773);
xor UO_2311 (O_2311,N_49607,N_49851);
and UO_2312 (O_2312,N_49616,N_49650);
nor UO_2313 (O_2313,N_49749,N_49519);
nor UO_2314 (O_2314,N_49685,N_49990);
or UO_2315 (O_2315,N_49655,N_49606);
nand UO_2316 (O_2316,N_49776,N_49558);
nand UO_2317 (O_2317,N_49970,N_49994);
and UO_2318 (O_2318,N_49763,N_49536);
nor UO_2319 (O_2319,N_49836,N_49673);
xnor UO_2320 (O_2320,N_49937,N_49858);
and UO_2321 (O_2321,N_49876,N_49652);
nand UO_2322 (O_2322,N_49756,N_49633);
nor UO_2323 (O_2323,N_49991,N_49672);
nand UO_2324 (O_2324,N_49672,N_49760);
nor UO_2325 (O_2325,N_49818,N_49549);
nor UO_2326 (O_2326,N_49664,N_49938);
or UO_2327 (O_2327,N_49740,N_49515);
nor UO_2328 (O_2328,N_49727,N_49872);
or UO_2329 (O_2329,N_49888,N_49909);
nand UO_2330 (O_2330,N_49871,N_49538);
xnor UO_2331 (O_2331,N_49723,N_49517);
nor UO_2332 (O_2332,N_49944,N_49957);
nand UO_2333 (O_2333,N_49926,N_49955);
nor UO_2334 (O_2334,N_49538,N_49507);
or UO_2335 (O_2335,N_49747,N_49681);
or UO_2336 (O_2336,N_49998,N_49822);
nand UO_2337 (O_2337,N_49998,N_49544);
nor UO_2338 (O_2338,N_49890,N_49500);
and UO_2339 (O_2339,N_49877,N_49531);
or UO_2340 (O_2340,N_49979,N_49744);
nor UO_2341 (O_2341,N_49642,N_49749);
or UO_2342 (O_2342,N_49682,N_49689);
or UO_2343 (O_2343,N_49767,N_49567);
and UO_2344 (O_2344,N_49975,N_49951);
nor UO_2345 (O_2345,N_49871,N_49926);
or UO_2346 (O_2346,N_49823,N_49522);
nand UO_2347 (O_2347,N_49889,N_49676);
and UO_2348 (O_2348,N_49630,N_49607);
xnor UO_2349 (O_2349,N_49856,N_49630);
or UO_2350 (O_2350,N_49580,N_49504);
or UO_2351 (O_2351,N_49876,N_49549);
nand UO_2352 (O_2352,N_49521,N_49653);
or UO_2353 (O_2353,N_49837,N_49759);
and UO_2354 (O_2354,N_49577,N_49881);
nand UO_2355 (O_2355,N_49920,N_49680);
nand UO_2356 (O_2356,N_49715,N_49941);
xor UO_2357 (O_2357,N_49535,N_49698);
and UO_2358 (O_2358,N_49892,N_49651);
and UO_2359 (O_2359,N_49695,N_49984);
and UO_2360 (O_2360,N_49794,N_49652);
nand UO_2361 (O_2361,N_49843,N_49986);
xor UO_2362 (O_2362,N_49717,N_49671);
or UO_2363 (O_2363,N_49544,N_49963);
nor UO_2364 (O_2364,N_49917,N_49725);
nand UO_2365 (O_2365,N_49774,N_49679);
xnor UO_2366 (O_2366,N_49933,N_49891);
or UO_2367 (O_2367,N_49857,N_49785);
or UO_2368 (O_2368,N_49870,N_49898);
nor UO_2369 (O_2369,N_49809,N_49653);
nor UO_2370 (O_2370,N_49609,N_49923);
nor UO_2371 (O_2371,N_49909,N_49846);
xor UO_2372 (O_2372,N_49975,N_49591);
xor UO_2373 (O_2373,N_49603,N_49546);
and UO_2374 (O_2374,N_49514,N_49548);
nand UO_2375 (O_2375,N_49676,N_49781);
xnor UO_2376 (O_2376,N_49961,N_49965);
and UO_2377 (O_2377,N_49692,N_49843);
nand UO_2378 (O_2378,N_49996,N_49854);
nand UO_2379 (O_2379,N_49669,N_49802);
xnor UO_2380 (O_2380,N_49619,N_49577);
nand UO_2381 (O_2381,N_49563,N_49939);
xnor UO_2382 (O_2382,N_49737,N_49584);
or UO_2383 (O_2383,N_49978,N_49638);
nand UO_2384 (O_2384,N_49614,N_49656);
nor UO_2385 (O_2385,N_49658,N_49519);
xnor UO_2386 (O_2386,N_49539,N_49904);
xnor UO_2387 (O_2387,N_49896,N_49855);
xnor UO_2388 (O_2388,N_49518,N_49923);
or UO_2389 (O_2389,N_49995,N_49616);
xor UO_2390 (O_2390,N_49606,N_49614);
or UO_2391 (O_2391,N_49831,N_49862);
nor UO_2392 (O_2392,N_49854,N_49525);
or UO_2393 (O_2393,N_49822,N_49791);
nand UO_2394 (O_2394,N_49540,N_49835);
and UO_2395 (O_2395,N_49694,N_49919);
nand UO_2396 (O_2396,N_49902,N_49665);
or UO_2397 (O_2397,N_49651,N_49985);
nor UO_2398 (O_2398,N_49678,N_49918);
nor UO_2399 (O_2399,N_49509,N_49597);
nor UO_2400 (O_2400,N_49503,N_49607);
nand UO_2401 (O_2401,N_49736,N_49768);
nor UO_2402 (O_2402,N_49607,N_49910);
or UO_2403 (O_2403,N_49715,N_49928);
xnor UO_2404 (O_2404,N_49500,N_49571);
xor UO_2405 (O_2405,N_49621,N_49914);
and UO_2406 (O_2406,N_49885,N_49679);
and UO_2407 (O_2407,N_49920,N_49998);
xor UO_2408 (O_2408,N_49998,N_49936);
nand UO_2409 (O_2409,N_49517,N_49854);
and UO_2410 (O_2410,N_49945,N_49786);
or UO_2411 (O_2411,N_49523,N_49569);
nand UO_2412 (O_2412,N_49816,N_49717);
xnor UO_2413 (O_2413,N_49790,N_49897);
nand UO_2414 (O_2414,N_49885,N_49998);
nor UO_2415 (O_2415,N_49534,N_49549);
or UO_2416 (O_2416,N_49862,N_49868);
nand UO_2417 (O_2417,N_49698,N_49792);
nand UO_2418 (O_2418,N_49999,N_49733);
nand UO_2419 (O_2419,N_49659,N_49640);
xnor UO_2420 (O_2420,N_49651,N_49890);
nand UO_2421 (O_2421,N_49616,N_49591);
xor UO_2422 (O_2422,N_49849,N_49613);
or UO_2423 (O_2423,N_49642,N_49679);
and UO_2424 (O_2424,N_49999,N_49822);
nor UO_2425 (O_2425,N_49913,N_49856);
and UO_2426 (O_2426,N_49987,N_49775);
nor UO_2427 (O_2427,N_49702,N_49937);
and UO_2428 (O_2428,N_49793,N_49992);
or UO_2429 (O_2429,N_49680,N_49621);
nand UO_2430 (O_2430,N_49852,N_49925);
nand UO_2431 (O_2431,N_49697,N_49955);
or UO_2432 (O_2432,N_49576,N_49938);
xor UO_2433 (O_2433,N_49765,N_49651);
nand UO_2434 (O_2434,N_49976,N_49901);
or UO_2435 (O_2435,N_49751,N_49693);
xnor UO_2436 (O_2436,N_49792,N_49589);
or UO_2437 (O_2437,N_49644,N_49838);
nor UO_2438 (O_2438,N_49590,N_49912);
nor UO_2439 (O_2439,N_49819,N_49512);
and UO_2440 (O_2440,N_49568,N_49756);
nor UO_2441 (O_2441,N_49650,N_49800);
nor UO_2442 (O_2442,N_49721,N_49650);
and UO_2443 (O_2443,N_49717,N_49675);
nor UO_2444 (O_2444,N_49766,N_49808);
xor UO_2445 (O_2445,N_49609,N_49920);
nor UO_2446 (O_2446,N_49624,N_49968);
xnor UO_2447 (O_2447,N_49573,N_49940);
xnor UO_2448 (O_2448,N_49982,N_49838);
xnor UO_2449 (O_2449,N_49516,N_49611);
nand UO_2450 (O_2450,N_49513,N_49845);
or UO_2451 (O_2451,N_49765,N_49841);
xor UO_2452 (O_2452,N_49716,N_49956);
nand UO_2453 (O_2453,N_49523,N_49909);
xor UO_2454 (O_2454,N_49879,N_49676);
xor UO_2455 (O_2455,N_49953,N_49974);
nand UO_2456 (O_2456,N_49585,N_49899);
or UO_2457 (O_2457,N_49758,N_49818);
nand UO_2458 (O_2458,N_49881,N_49896);
xor UO_2459 (O_2459,N_49644,N_49709);
or UO_2460 (O_2460,N_49698,N_49808);
or UO_2461 (O_2461,N_49510,N_49754);
nor UO_2462 (O_2462,N_49976,N_49786);
nand UO_2463 (O_2463,N_49870,N_49651);
or UO_2464 (O_2464,N_49566,N_49849);
or UO_2465 (O_2465,N_49666,N_49902);
or UO_2466 (O_2466,N_49652,N_49747);
nand UO_2467 (O_2467,N_49671,N_49557);
nor UO_2468 (O_2468,N_49853,N_49933);
xor UO_2469 (O_2469,N_49594,N_49588);
nor UO_2470 (O_2470,N_49838,N_49868);
xnor UO_2471 (O_2471,N_49578,N_49734);
nand UO_2472 (O_2472,N_49776,N_49665);
nor UO_2473 (O_2473,N_49654,N_49897);
xor UO_2474 (O_2474,N_49877,N_49620);
or UO_2475 (O_2475,N_49608,N_49609);
or UO_2476 (O_2476,N_49889,N_49702);
and UO_2477 (O_2477,N_49881,N_49541);
or UO_2478 (O_2478,N_49664,N_49543);
nor UO_2479 (O_2479,N_49744,N_49527);
or UO_2480 (O_2480,N_49625,N_49533);
xor UO_2481 (O_2481,N_49765,N_49766);
nor UO_2482 (O_2482,N_49706,N_49854);
nor UO_2483 (O_2483,N_49972,N_49617);
or UO_2484 (O_2484,N_49775,N_49594);
xnor UO_2485 (O_2485,N_49581,N_49533);
nor UO_2486 (O_2486,N_49716,N_49847);
xnor UO_2487 (O_2487,N_49930,N_49595);
nand UO_2488 (O_2488,N_49753,N_49671);
and UO_2489 (O_2489,N_49517,N_49984);
xnor UO_2490 (O_2490,N_49685,N_49846);
nor UO_2491 (O_2491,N_49758,N_49520);
xnor UO_2492 (O_2492,N_49532,N_49847);
and UO_2493 (O_2493,N_49715,N_49614);
or UO_2494 (O_2494,N_49683,N_49786);
nand UO_2495 (O_2495,N_49894,N_49941);
and UO_2496 (O_2496,N_49605,N_49700);
nor UO_2497 (O_2497,N_49562,N_49985);
nor UO_2498 (O_2498,N_49829,N_49642);
nor UO_2499 (O_2499,N_49773,N_49616);
and UO_2500 (O_2500,N_49846,N_49579);
nor UO_2501 (O_2501,N_49538,N_49540);
nor UO_2502 (O_2502,N_49922,N_49527);
and UO_2503 (O_2503,N_49792,N_49602);
nand UO_2504 (O_2504,N_49824,N_49596);
xnor UO_2505 (O_2505,N_49645,N_49800);
xor UO_2506 (O_2506,N_49614,N_49858);
nor UO_2507 (O_2507,N_49988,N_49720);
and UO_2508 (O_2508,N_49790,N_49693);
and UO_2509 (O_2509,N_49620,N_49773);
nand UO_2510 (O_2510,N_49554,N_49634);
nor UO_2511 (O_2511,N_49942,N_49753);
and UO_2512 (O_2512,N_49596,N_49739);
xnor UO_2513 (O_2513,N_49539,N_49943);
or UO_2514 (O_2514,N_49911,N_49666);
nand UO_2515 (O_2515,N_49931,N_49530);
nand UO_2516 (O_2516,N_49626,N_49792);
nor UO_2517 (O_2517,N_49645,N_49912);
nand UO_2518 (O_2518,N_49959,N_49514);
and UO_2519 (O_2519,N_49838,N_49511);
nor UO_2520 (O_2520,N_49986,N_49514);
or UO_2521 (O_2521,N_49731,N_49623);
xnor UO_2522 (O_2522,N_49599,N_49579);
xor UO_2523 (O_2523,N_49708,N_49890);
nor UO_2524 (O_2524,N_49532,N_49578);
or UO_2525 (O_2525,N_49842,N_49771);
nand UO_2526 (O_2526,N_49671,N_49619);
nand UO_2527 (O_2527,N_49576,N_49789);
nor UO_2528 (O_2528,N_49609,N_49599);
nor UO_2529 (O_2529,N_49622,N_49692);
nand UO_2530 (O_2530,N_49502,N_49801);
or UO_2531 (O_2531,N_49693,N_49828);
xor UO_2532 (O_2532,N_49726,N_49769);
and UO_2533 (O_2533,N_49587,N_49824);
and UO_2534 (O_2534,N_49778,N_49819);
nand UO_2535 (O_2535,N_49975,N_49702);
or UO_2536 (O_2536,N_49736,N_49992);
nor UO_2537 (O_2537,N_49961,N_49702);
xor UO_2538 (O_2538,N_49662,N_49913);
and UO_2539 (O_2539,N_49576,N_49638);
nor UO_2540 (O_2540,N_49600,N_49999);
xnor UO_2541 (O_2541,N_49877,N_49834);
nand UO_2542 (O_2542,N_49608,N_49829);
and UO_2543 (O_2543,N_49817,N_49546);
and UO_2544 (O_2544,N_49808,N_49854);
xor UO_2545 (O_2545,N_49570,N_49590);
nor UO_2546 (O_2546,N_49611,N_49972);
or UO_2547 (O_2547,N_49643,N_49585);
and UO_2548 (O_2548,N_49648,N_49709);
and UO_2549 (O_2549,N_49537,N_49570);
xor UO_2550 (O_2550,N_49937,N_49905);
or UO_2551 (O_2551,N_49874,N_49940);
and UO_2552 (O_2552,N_49817,N_49660);
and UO_2553 (O_2553,N_49601,N_49993);
nor UO_2554 (O_2554,N_49610,N_49565);
nor UO_2555 (O_2555,N_49902,N_49522);
xor UO_2556 (O_2556,N_49710,N_49544);
or UO_2557 (O_2557,N_49565,N_49733);
nor UO_2558 (O_2558,N_49561,N_49755);
and UO_2559 (O_2559,N_49916,N_49955);
and UO_2560 (O_2560,N_49988,N_49522);
nor UO_2561 (O_2561,N_49886,N_49882);
and UO_2562 (O_2562,N_49988,N_49665);
nand UO_2563 (O_2563,N_49573,N_49748);
xnor UO_2564 (O_2564,N_49784,N_49915);
xnor UO_2565 (O_2565,N_49636,N_49773);
nor UO_2566 (O_2566,N_49684,N_49591);
or UO_2567 (O_2567,N_49760,N_49735);
nand UO_2568 (O_2568,N_49687,N_49596);
or UO_2569 (O_2569,N_49872,N_49645);
nand UO_2570 (O_2570,N_49620,N_49858);
nand UO_2571 (O_2571,N_49761,N_49500);
xnor UO_2572 (O_2572,N_49518,N_49645);
xor UO_2573 (O_2573,N_49872,N_49550);
xnor UO_2574 (O_2574,N_49630,N_49828);
nand UO_2575 (O_2575,N_49753,N_49867);
nand UO_2576 (O_2576,N_49815,N_49528);
nor UO_2577 (O_2577,N_49898,N_49592);
nand UO_2578 (O_2578,N_49793,N_49618);
or UO_2579 (O_2579,N_49989,N_49987);
nor UO_2580 (O_2580,N_49573,N_49696);
and UO_2581 (O_2581,N_49746,N_49897);
or UO_2582 (O_2582,N_49821,N_49816);
nor UO_2583 (O_2583,N_49617,N_49813);
xnor UO_2584 (O_2584,N_49697,N_49690);
nor UO_2585 (O_2585,N_49691,N_49657);
xnor UO_2586 (O_2586,N_49650,N_49606);
nand UO_2587 (O_2587,N_49550,N_49703);
nand UO_2588 (O_2588,N_49519,N_49622);
or UO_2589 (O_2589,N_49570,N_49555);
and UO_2590 (O_2590,N_49916,N_49548);
and UO_2591 (O_2591,N_49934,N_49835);
xor UO_2592 (O_2592,N_49733,N_49977);
nand UO_2593 (O_2593,N_49664,N_49567);
xnor UO_2594 (O_2594,N_49729,N_49525);
nand UO_2595 (O_2595,N_49582,N_49958);
xor UO_2596 (O_2596,N_49861,N_49823);
nor UO_2597 (O_2597,N_49723,N_49580);
nor UO_2598 (O_2598,N_49590,N_49981);
or UO_2599 (O_2599,N_49600,N_49505);
or UO_2600 (O_2600,N_49734,N_49800);
and UO_2601 (O_2601,N_49819,N_49972);
or UO_2602 (O_2602,N_49755,N_49932);
and UO_2603 (O_2603,N_49653,N_49561);
and UO_2604 (O_2604,N_49755,N_49908);
and UO_2605 (O_2605,N_49598,N_49758);
xor UO_2606 (O_2606,N_49806,N_49708);
nand UO_2607 (O_2607,N_49808,N_49704);
and UO_2608 (O_2608,N_49938,N_49863);
or UO_2609 (O_2609,N_49818,N_49773);
and UO_2610 (O_2610,N_49879,N_49669);
xnor UO_2611 (O_2611,N_49573,N_49859);
xor UO_2612 (O_2612,N_49726,N_49713);
or UO_2613 (O_2613,N_49552,N_49871);
and UO_2614 (O_2614,N_49757,N_49937);
and UO_2615 (O_2615,N_49717,N_49773);
xor UO_2616 (O_2616,N_49598,N_49869);
xor UO_2617 (O_2617,N_49970,N_49693);
or UO_2618 (O_2618,N_49676,N_49644);
or UO_2619 (O_2619,N_49760,N_49758);
and UO_2620 (O_2620,N_49600,N_49552);
nor UO_2621 (O_2621,N_49812,N_49760);
nand UO_2622 (O_2622,N_49926,N_49787);
nor UO_2623 (O_2623,N_49636,N_49712);
xnor UO_2624 (O_2624,N_49780,N_49742);
or UO_2625 (O_2625,N_49642,N_49943);
nand UO_2626 (O_2626,N_49613,N_49851);
and UO_2627 (O_2627,N_49667,N_49514);
nor UO_2628 (O_2628,N_49533,N_49942);
xor UO_2629 (O_2629,N_49844,N_49865);
and UO_2630 (O_2630,N_49637,N_49935);
xor UO_2631 (O_2631,N_49859,N_49973);
nor UO_2632 (O_2632,N_49503,N_49875);
nand UO_2633 (O_2633,N_49513,N_49742);
or UO_2634 (O_2634,N_49948,N_49532);
xnor UO_2635 (O_2635,N_49956,N_49989);
or UO_2636 (O_2636,N_49651,N_49991);
or UO_2637 (O_2637,N_49613,N_49845);
and UO_2638 (O_2638,N_49668,N_49640);
nor UO_2639 (O_2639,N_49957,N_49623);
nor UO_2640 (O_2640,N_49552,N_49795);
or UO_2641 (O_2641,N_49671,N_49758);
nand UO_2642 (O_2642,N_49693,N_49619);
and UO_2643 (O_2643,N_49847,N_49836);
xor UO_2644 (O_2644,N_49671,N_49896);
xnor UO_2645 (O_2645,N_49802,N_49567);
or UO_2646 (O_2646,N_49605,N_49751);
and UO_2647 (O_2647,N_49689,N_49501);
and UO_2648 (O_2648,N_49821,N_49603);
and UO_2649 (O_2649,N_49922,N_49594);
nand UO_2650 (O_2650,N_49925,N_49566);
xor UO_2651 (O_2651,N_49988,N_49796);
nand UO_2652 (O_2652,N_49796,N_49790);
or UO_2653 (O_2653,N_49881,N_49692);
nor UO_2654 (O_2654,N_49516,N_49768);
nand UO_2655 (O_2655,N_49930,N_49652);
and UO_2656 (O_2656,N_49964,N_49713);
or UO_2657 (O_2657,N_49523,N_49639);
or UO_2658 (O_2658,N_49774,N_49861);
xor UO_2659 (O_2659,N_49994,N_49886);
xnor UO_2660 (O_2660,N_49582,N_49657);
nor UO_2661 (O_2661,N_49534,N_49902);
xnor UO_2662 (O_2662,N_49855,N_49772);
nor UO_2663 (O_2663,N_49511,N_49956);
xnor UO_2664 (O_2664,N_49508,N_49887);
nor UO_2665 (O_2665,N_49760,N_49915);
nor UO_2666 (O_2666,N_49741,N_49605);
and UO_2667 (O_2667,N_49749,N_49981);
nand UO_2668 (O_2668,N_49999,N_49893);
and UO_2669 (O_2669,N_49843,N_49775);
xor UO_2670 (O_2670,N_49895,N_49729);
nor UO_2671 (O_2671,N_49835,N_49721);
nor UO_2672 (O_2672,N_49850,N_49816);
and UO_2673 (O_2673,N_49709,N_49773);
or UO_2674 (O_2674,N_49882,N_49593);
nand UO_2675 (O_2675,N_49626,N_49572);
xor UO_2676 (O_2676,N_49879,N_49773);
and UO_2677 (O_2677,N_49920,N_49676);
and UO_2678 (O_2678,N_49518,N_49918);
nand UO_2679 (O_2679,N_49506,N_49991);
xnor UO_2680 (O_2680,N_49780,N_49552);
nand UO_2681 (O_2681,N_49654,N_49659);
nor UO_2682 (O_2682,N_49874,N_49567);
nand UO_2683 (O_2683,N_49964,N_49716);
or UO_2684 (O_2684,N_49881,N_49628);
or UO_2685 (O_2685,N_49633,N_49918);
or UO_2686 (O_2686,N_49882,N_49694);
or UO_2687 (O_2687,N_49838,N_49909);
nand UO_2688 (O_2688,N_49673,N_49742);
or UO_2689 (O_2689,N_49750,N_49617);
xor UO_2690 (O_2690,N_49789,N_49903);
xnor UO_2691 (O_2691,N_49836,N_49952);
or UO_2692 (O_2692,N_49518,N_49659);
nor UO_2693 (O_2693,N_49858,N_49654);
xnor UO_2694 (O_2694,N_49533,N_49913);
xnor UO_2695 (O_2695,N_49529,N_49919);
nor UO_2696 (O_2696,N_49520,N_49942);
and UO_2697 (O_2697,N_49899,N_49638);
and UO_2698 (O_2698,N_49801,N_49886);
or UO_2699 (O_2699,N_49554,N_49766);
or UO_2700 (O_2700,N_49566,N_49834);
and UO_2701 (O_2701,N_49622,N_49564);
and UO_2702 (O_2702,N_49548,N_49731);
nor UO_2703 (O_2703,N_49979,N_49531);
or UO_2704 (O_2704,N_49910,N_49852);
nor UO_2705 (O_2705,N_49993,N_49785);
and UO_2706 (O_2706,N_49685,N_49526);
or UO_2707 (O_2707,N_49668,N_49868);
xnor UO_2708 (O_2708,N_49666,N_49771);
nand UO_2709 (O_2709,N_49553,N_49748);
nor UO_2710 (O_2710,N_49545,N_49827);
nand UO_2711 (O_2711,N_49958,N_49991);
and UO_2712 (O_2712,N_49952,N_49810);
nand UO_2713 (O_2713,N_49552,N_49804);
or UO_2714 (O_2714,N_49522,N_49559);
nor UO_2715 (O_2715,N_49987,N_49872);
and UO_2716 (O_2716,N_49903,N_49811);
nor UO_2717 (O_2717,N_49811,N_49786);
xnor UO_2718 (O_2718,N_49821,N_49511);
nor UO_2719 (O_2719,N_49589,N_49743);
xnor UO_2720 (O_2720,N_49919,N_49710);
and UO_2721 (O_2721,N_49535,N_49731);
xor UO_2722 (O_2722,N_49766,N_49546);
and UO_2723 (O_2723,N_49814,N_49725);
nand UO_2724 (O_2724,N_49591,N_49897);
xnor UO_2725 (O_2725,N_49999,N_49664);
or UO_2726 (O_2726,N_49502,N_49963);
and UO_2727 (O_2727,N_49842,N_49641);
xnor UO_2728 (O_2728,N_49635,N_49999);
xor UO_2729 (O_2729,N_49947,N_49670);
or UO_2730 (O_2730,N_49718,N_49577);
and UO_2731 (O_2731,N_49611,N_49801);
and UO_2732 (O_2732,N_49721,N_49876);
and UO_2733 (O_2733,N_49974,N_49589);
nor UO_2734 (O_2734,N_49695,N_49503);
nor UO_2735 (O_2735,N_49895,N_49657);
nand UO_2736 (O_2736,N_49617,N_49644);
or UO_2737 (O_2737,N_49784,N_49901);
nand UO_2738 (O_2738,N_49741,N_49695);
and UO_2739 (O_2739,N_49582,N_49750);
xnor UO_2740 (O_2740,N_49840,N_49707);
nor UO_2741 (O_2741,N_49911,N_49893);
or UO_2742 (O_2742,N_49519,N_49946);
and UO_2743 (O_2743,N_49591,N_49758);
or UO_2744 (O_2744,N_49883,N_49968);
nor UO_2745 (O_2745,N_49517,N_49740);
nand UO_2746 (O_2746,N_49700,N_49847);
xor UO_2747 (O_2747,N_49801,N_49574);
nor UO_2748 (O_2748,N_49963,N_49679);
and UO_2749 (O_2749,N_49642,N_49998);
xor UO_2750 (O_2750,N_49977,N_49691);
nand UO_2751 (O_2751,N_49970,N_49616);
nand UO_2752 (O_2752,N_49997,N_49957);
xnor UO_2753 (O_2753,N_49932,N_49577);
nand UO_2754 (O_2754,N_49652,N_49677);
nand UO_2755 (O_2755,N_49940,N_49538);
nand UO_2756 (O_2756,N_49692,N_49982);
or UO_2757 (O_2757,N_49591,N_49985);
xnor UO_2758 (O_2758,N_49895,N_49600);
or UO_2759 (O_2759,N_49542,N_49595);
nor UO_2760 (O_2760,N_49925,N_49899);
nand UO_2761 (O_2761,N_49809,N_49584);
nand UO_2762 (O_2762,N_49576,N_49679);
or UO_2763 (O_2763,N_49510,N_49604);
and UO_2764 (O_2764,N_49738,N_49816);
nand UO_2765 (O_2765,N_49533,N_49737);
or UO_2766 (O_2766,N_49628,N_49975);
or UO_2767 (O_2767,N_49735,N_49739);
xnor UO_2768 (O_2768,N_49633,N_49680);
or UO_2769 (O_2769,N_49603,N_49909);
nor UO_2770 (O_2770,N_49858,N_49582);
xor UO_2771 (O_2771,N_49597,N_49731);
and UO_2772 (O_2772,N_49824,N_49884);
nand UO_2773 (O_2773,N_49874,N_49614);
or UO_2774 (O_2774,N_49653,N_49818);
nor UO_2775 (O_2775,N_49621,N_49837);
nor UO_2776 (O_2776,N_49865,N_49738);
and UO_2777 (O_2777,N_49656,N_49854);
xnor UO_2778 (O_2778,N_49762,N_49886);
xor UO_2779 (O_2779,N_49544,N_49596);
or UO_2780 (O_2780,N_49581,N_49970);
or UO_2781 (O_2781,N_49548,N_49735);
and UO_2782 (O_2782,N_49522,N_49732);
and UO_2783 (O_2783,N_49661,N_49622);
nand UO_2784 (O_2784,N_49555,N_49576);
nor UO_2785 (O_2785,N_49651,N_49658);
nand UO_2786 (O_2786,N_49908,N_49824);
and UO_2787 (O_2787,N_49715,N_49567);
nor UO_2788 (O_2788,N_49572,N_49897);
xnor UO_2789 (O_2789,N_49536,N_49981);
or UO_2790 (O_2790,N_49670,N_49807);
and UO_2791 (O_2791,N_49961,N_49673);
nand UO_2792 (O_2792,N_49740,N_49947);
nor UO_2793 (O_2793,N_49875,N_49795);
and UO_2794 (O_2794,N_49782,N_49868);
nand UO_2795 (O_2795,N_49938,N_49702);
or UO_2796 (O_2796,N_49965,N_49978);
nor UO_2797 (O_2797,N_49659,N_49918);
nand UO_2798 (O_2798,N_49529,N_49917);
or UO_2799 (O_2799,N_49956,N_49759);
xor UO_2800 (O_2800,N_49822,N_49969);
nand UO_2801 (O_2801,N_49588,N_49858);
nand UO_2802 (O_2802,N_49839,N_49656);
xnor UO_2803 (O_2803,N_49678,N_49748);
xor UO_2804 (O_2804,N_49986,N_49574);
nand UO_2805 (O_2805,N_49573,N_49694);
xor UO_2806 (O_2806,N_49630,N_49736);
xnor UO_2807 (O_2807,N_49859,N_49783);
xnor UO_2808 (O_2808,N_49774,N_49525);
nor UO_2809 (O_2809,N_49965,N_49857);
or UO_2810 (O_2810,N_49503,N_49633);
xnor UO_2811 (O_2811,N_49535,N_49846);
xor UO_2812 (O_2812,N_49554,N_49852);
xor UO_2813 (O_2813,N_49789,N_49995);
xor UO_2814 (O_2814,N_49747,N_49887);
or UO_2815 (O_2815,N_49690,N_49505);
nor UO_2816 (O_2816,N_49647,N_49966);
xor UO_2817 (O_2817,N_49582,N_49936);
or UO_2818 (O_2818,N_49621,N_49931);
or UO_2819 (O_2819,N_49634,N_49743);
and UO_2820 (O_2820,N_49680,N_49960);
nor UO_2821 (O_2821,N_49862,N_49614);
nor UO_2822 (O_2822,N_49555,N_49620);
nand UO_2823 (O_2823,N_49680,N_49957);
nand UO_2824 (O_2824,N_49614,N_49809);
or UO_2825 (O_2825,N_49527,N_49554);
xor UO_2826 (O_2826,N_49531,N_49530);
or UO_2827 (O_2827,N_49946,N_49791);
or UO_2828 (O_2828,N_49650,N_49903);
xnor UO_2829 (O_2829,N_49971,N_49857);
nor UO_2830 (O_2830,N_49581,N_49808);
nand UO_2831 (O_2831,N_49556,N_49504);
nor UO_2832 (O_2832,N_49553,N_49548);
nor UO_2833 (O_2833,N_49690,N_49774);
nor UO_2834 (O_2834,N_49672,N_49720);
and UO_2835 (O_2835,N_49743,N_49875);
and UO_2836 (O_2836,N_49803,N_49696);
nand UO_2837 (O_2837,N_49924,N_49850);
xnor UO_2838 (O_2838,N_49911,N_49603);
xnor UO_2839 (O_2839,N_49798,N_49680);
nor UO_2840 (O_2840,N_49864,N_49941);
xor UO_2841 (O_2841,N_49636,N_49976);
or UO_2842 (O_2842,N_49620,N_49777);
xor UO_2843 (O_2843,N_49756,N_49844);
xor UO_2844 (O_2844,N_49830,N_49924);
nand UO_2845 (O_2845,N_49873,N_49687);
and UO_2846 (O_2846,N_49858,N_49878);
xnor UO_2847 (O_2847,N_49649,N_49817);
xor UO_2848 (O_2848,N_49543,N_49523);
or UO_2849 (O_2849,N_49973,N_49950);
and UO_2850 (O_2850,N_49707,N_49885);
nor UO_2851 (O_2851,N_49901,N_49892);
nand UO_2852 (O_2852,N_49649,N_49623);
or UO_2853 (O_2853,N_49738,N_49543);
nor UO_2854 (O_2854,N_49732,N_49913);
or UO_2855 (O_2855,N_49742,N_49512);
and UO_2856 (O_2856,N_49839,N_49702);
or UO_2857 (O_2857,N_49819,N_49641);
xor UO_2858 (O_2858,N_49997,N_49568);
nor UO_2859 (O_2859,N_49667,N_49590);
and UO_2860 (O_2860,N_49993,N_49940);
nand UO_2861 (O_2861,N_49585,N_49660);
and UO_2862 (O_2862,N_49975,N_49541);
and UO_2863 (O_2863,N_49990,N_49967);
and UO_2864 (O_2864,N_49512,N_49666);
or UO_2865 (O_2865,N_49859,N_49650);
or UO_2866 (O_2866,N_49515,N_49931);
or UO_2867 (O_2867,N_49510,N_49548);
nand UO_2868 (O_2868,N_49696,N_49717);
nor UO_2869 (O_2869,N_49834,N_49707);
or UO_2870 (O_2870,N_49653,N_49918);
and UO_2871 (O_2871,N_49506,N_49524);
and UO_2872 (O_2872,N_49672,N_49727);
xnor UO_2873 (O_2873,N_49944,N_49794);
and UO_2874 (O_2874,N_49569,N_49787);
nand UO_2875 (O_2875,N_49873,N_49784);
nor UO_2876 (O_2876,N_49622,N_49571);
nand UO_2877 (O_2877,N_49935,N_49852);
nand UO_2878 (O_2878,N_49904,N_49824);
xnor UO_2879 (O_2879,N_49824,N_49922);
nand UO_2880 (O_2880,N_49602,N_49642);
xnor UO_2881 (O_2881,N_49563,N_49668);
xor UO_2882 (O_2882,N_49828,N_49775);
and UO_2883 (O_2883,N_49613,N_49972);
xnor UO_2884 (O_2884,N_49575,N_49706);
xor UO_2885 (O_2885,N_49628,N_49617);
nor UO_2886 (O_2886,N_49703,N_49587);
xor UO_2887 (O_2887,N_49759,N_49715);
or UO_2888 (O_2888,N_49681,N_49537);
or UO_2889 (O_2889,N_49626,N_49574);
nor UO_2890 (O_2890,N_49687,N_49893);
xnor UO_2891 (O_2891,N_49913,N_49798);
and UO_2892 (O_2892,N_49793,N_49789);
or UO_2893 (O_2893,N_49991,N_49637);
or UO_2894 (O_2894,N_49630,N_49866);
and UO_2895 (O_2895,N_49564,N_49624);
and UO_2896 (O_2896,N_49620,N_49784);
xor UO_2897 (O_2897,N_49999,N_49978);
nand UO_2898 (O_2898,N_49646,N_49584);
or UO_2899 (O_2899,N_49639,N_49875);
and UO_2900 (O_2900,N_49944,N_49555);
nand UO_2901 (O_2901,N_49649,N_49540);
or UO_2902 (O_2902,N_49751,N_49706);
nand UO_2903 (O_2903,N_49570,N_49709);
nor UO_2904 (O_2904,N_49765,N_49911);
and UO_2905 (O_2905,N_49923,N_49573);
or UO_2906 (O_2906,N_49883,N_49916);
or UO_2907 (O_2907,N_49705,N_49889);
and UO_2908 (O_2908,N_49518,N_49676);
nand UO_2909 (O_2909,N_49523,N_49799);
nand UO_2910 (O_2910,N_49642,N_49952);
nand UO_2911 (O_2911,N_49801,N_49566);
nand UO_2912 (O_2912,N_49643,N_49966);
nor UO_2913 (O_2913,N_49809,N_49701);
nand UO_2914 (O_2914,N_49555,N_49931);
nand UO_2915 (O_2915,N_49726,N_49761);
or UO_2916 (O_2916,N_49779,N_49976);
or UO_2917 (O_2917,N_49774,N_49645);
nor UO_2918 (O_2918,N_49721,N_49848);
xnor UO_2919 (O_2919,N_49925,N_49688);
or UO_2920 (O_2920,N_49849,N_49999);
xnor UO_2921 (O_2921,N_49761,N_49686);
and UO_2922 (O_2922,N_49759,N_49716);
nand UO_2923 (O_2923,N_49530,N_49684);
or UO_2924 (O_2924,N_49927,N_49690);
nor UO_2925 (O_2925,N_49932,N_49833);
and UO_2926 (O_2926,N_49777,N_49573);
and UO_2927 (O_2927,N_49932,N_49578);
nand UO_2928 (O_2928,N_49793,N_49981);
nor UO_2929 (O_2929,N_49938,N_49721);
or UO_2930 (O_2930,N_49531,N_49690);
nor UO_2931 (O_2931,N_49551,N_49981);
nand UO_2932 (O_2932,N_49592,N_49832);
xnor UO_2933 (O_2933,N_49725,N_49668);
xor UO_2934 (O_2934,N_49730,N_49895);
xnor UO_2935 (O_2935,N_49681,N_49887);
nand UO_2936 (O_2936,N_49643,N_49664);
and UO_2937 (O_2937,N_49842,N_49605);
xor UO_2938 (O_2938,N_49744,N_49641);
or UO_2939 (O_2939,N_49865,N_49876);
or UO_2940 (O_2940,N_49685,N_49694);
or UO_2941 (O_2941,N_49698,N_49675);
nor UO_2942 (O_2942,N_49785,N_49882);
and UO_2943 (O_2943,N_49567,N_49982);
or UO_2944 (O_2944,N_49906,N_49726);
xnor UO_2945 (O_2945,N_49980,N_49601);
and UO_2946 (O_2946,N_49796,N_49633);
or UO_2947 (O_2947,N_49730,N_49776);
nor UO_2948 (O_2948,N_49566,N_49678);
nand UO_2949 (O_2949,N_49762,N_49795);
xor UO_2950 (O_2950,N_49844,N_49663);
and UO_2951 (O_2951,N_49738,N_49826);
or UO_2952 (O_2952,N_49924,N_49737);
or UO_2953 (O_2953,N_49929,N_49619);
and UO_2954 (O_2954,N_49977,N_49517);
xnor UO_2955 (O_2955,N_49951,N_49504);
nor UO_2956 (O_2956,N_49554,N_49758);
nor UO_2957 (O_2957,N_49753,N_49899);
and UO_2958 (O_2958,N_49905,N_49938);
and UO_2959 (O_2959,N_49544,N_49598);
nand UO_2960 (O_2960,N_49821,N_49646);
xnor UO_2961 (O_2961,N_49935,N_49655);
and UO_2962 (O_2962,N_49890,N_49916);
nand UO_2963 (O_2963,N_49706,N_49598);
xor UO_2964 (O_2964,N_49637,N_49957);
and UO_2965 (O_2965,N_49518,N_49967);
nor UO_2966 (O_2966,N_49838,N_49720);
and UO_2967 (O_2967,N_49807,N_49565);
and UO_2968 (O_2968,N_49844,N_49845);
nor UO_2969 (O_2969,N_49679,N_49960);
nand UO_2970 (O_2970,N_49574,N_49611);
nand UO_2971 (O_2971,N_49668,N_49609);
or UO_2972 (O_2972,N_49550,N_49585);
nand UO_2973 (O_2973,N_49909,N_49743);
or UO_2974 (O_2974,N_49525,N_49812);
and UO_2975 (O_2975,N_49516,N_49545);
xnor UO_2976 (O_2976,N_49758,N_49792);
nand UO_2977 (O_2977,N_49844,N_49704);
xor UO_2978 (O_2978,N_49785,N_49844);
and UO_2979 (O_2979,N_49561,N_49606);
or UO_2980 (O_2980,N_49504,N_49653);
xnor UO_2981 (O_2981,N_49703,N_49841);
xnor UO_2982 (O_2982,N_49575,N_49634);
nand UO_2983 (O_2983,N_49731,N_49557);
nor UO_2984 (O_2984,N_49990,N_49687);
nand UO_2985 (O_2985,N_49633,N_49882);
nand UO_2986 (O_2986,N_49586,N_49991);
xor UO_2987 (O_2987,N_49600,N_49673);
or UO_2988 (O_2988,N_49876,N_49868);
and UO_2989 (O_2989,N_49983,N_49738);
xnor UO_2990 (O_2990,N_49915,N_49614);
xor UO_2991 (O_2991,N_49682,N_49925);
nor UO_2992 (O_2992,N_49983,N_49880);
and UO_2993 (O_2993,N_49661,N_49642);
xnor UO_2994 (O_2994,N_49715,N_49938);
and UO_2995 (O_2995,N_49947,N_49509);
xnor UO_2996 (O_2996,N_49736,N_49742);
and UO_2997 (O_2997,N_49877,N_49544);
xnor UO_2998 (O_2998,N_49956,N_49761);
or UO_2999 (O_2999,N_49980,N_49765);
nor UO_3000 (O_3000,N_49636,N_49519);
and UO_3001 (O_3001,N_49825,N_49730);
and UO_3002 (O_3002,N_49994,N_49545);
xor UO_3003 (O_3003,N_49782,N_49908);
nor UO_3004 (O_3004,N_49505,N_49616);
nand UO_3005 (O_3005,N_49623,N_49723);
xnor UO_3006 (O_3006,N_49606,N_49542);
nand UO_3007 (O_3007,N_49716,N_49777);
or UO_3008 (O_3008,N_49715,N_49718);
nor UO_3009 (O_3009,N_49674,N_49773);
xnor UO_3010 (O_3010,N_49822,N_49945);
or UO_3011 (O_3011,N_49958,N_49696);
nor UO_3012 (O_3012,N_49895,N_49865);
and UO_3013 (O_3013,N_49604,N_49533);
or UO_3014 (O_3014,N_49984,N_49735);
nor UO_3015 (O_3015,N_49574,N_49810);
nor UO_3016 (O_3016,N_49555,N_49653);
nand UO_3017 (O_3017,N_49549,N_49916);
xor UO_3018 (O_3018,N_49686,N_49967);
xor UO_3019 (O_3019,N_49574,N_49647);
nor UO_3020 (O_3020,N_49515,N_49602);
xnor UO_3021 (O_3021,N_49899,N_49860);
nand UO_3022 (O_3022,N_49750,N_49622);
nor UO_3023 (O_3023,N_49707,N_49726);
xnor UO_3024 (O_3024,N_49918,N_49914);
and UO_3025 (O_3025,N_49781,N_49790);
or UO_3026 (O_3026,N_49730,N_49910);
or UO_3027 (O_3027,N_49836,N_49642);
xor UO_3028 (O_3028,N_49536,N_49508);
and UO_3029 (O_3029,N_49875,N_49891);
xnor UO_3030 (O_3030,N_49747,N_49594);
nor UO_3031 (O_3031,N_49767,N_49768);
nand UO_3032 (O_3032,N_49715,N_49827);
nand UO_3033 (O_3033,N_49595,N_49699);
nand UO_3034 (O_3034,N_49648,N_49757);
or UO_3035 (O_3035,N_49785,N_49935);
or UO_3036 (O_3036,N_49882,N_49839);
nand UO_3037 (O_3037,N_49943,N_49792);
nor UO_3038 (O_3038,N_49593,N_49968);
xor UO_3039 (O_3039,N_49957,N_49813);
and UO_3040 (O_3040,N_49771,N_49761);
nand UO_3041 (O_3041,N_49690,N_49728);
or UO_3042 (O_3042,N_49748,N_49930);
xor UO_3043 (O_3043,N_49651,N_49697);
and UO_3044 (O_3044,N_49534,N_49994);
nor UO_3045 (O_3045,N_49838,N_49857);
nor UO_3046 (O_3046,N_49600,N_49748);
xnor UO_3047 (O_3047,N_49729,N_49847);
nor UO_3048 (O_3048,N_49923,N_49904);
or UO_3049 (O_3049,N_49783,N_49912);
and UO_3050 (O_3050,N_49547,N_49732);
or UO_3051 (O_3051,N_49548,N_49508);
and UO_3052 (O_3052,N_49848,N_49525);
xor UO_3053 (O_3053,N_49771,N_49759);
or UO_3054 (O_3054,N_49644,N_49940);
and UO_3055 (O_3055,N_49970,N_49969);
and UO_3056 (O_3056,N_49646,N_49726);
or UO_3057 (O_3057,N_49845,N_49538);
and UO_3058 (O_3058,N_49903,N_49717);
xor UO_3059 (O_3059,N_49619,N_49816);
nor UO_3060 (O_3060,N_49719,N_49961);
nand UO_3061 (O_3061,N_49546,N_49611);
nor UO_3062 (O_3062,N_49638,N_49831);
nor UO_3063 (O_3063,N_49708,N_49978);
or UO_3064 (O_3064,N_49653,N_49554);
nor UO_3065 (O_3065,N_49957,N_49987);
nand UO_3066 (O_3066,N_49832,N_49737);
xor UO_3067 (O_3067,N_49724,N_49944);
or UO_3068 (O_3068,N_49727,N_49838);
and UO_3069 (O_3069,N_49983,N_49845);
and UO_3070 (O_3070,N_49694,N_49759);
nand UO_3071 (O_3071,N_49994,N_49748);
and UO_3072 (O_3072,N_49746,N_49969);
xnor UO_3073 (O_3073,N_49832,N_49731);
nor UO_3074 (O_3074,N_49839,N_49569);
xnor UO_3075 (O_3075,N_49774,N_49884);
xor UO_3076 (O_3076,N_49688,N_49552);
xor UO_3077 (O_3077,N_49762,N_49656);
and UO_3078 (O_3078,N_49911,N_49649);
or UO_3079 (O_3079,N_49810,N_49979);
xnor UO_3080 (O_3080,N_49769,N_49592);
nor UO_3081 (O_3081,N_49570,N_49705);
and UO_3082 (O_3082,N_49886,N_49963);
and UO_3083 (O_3083,N_49874,N_49838);
nand UO_3084 (O_3084,N_49654,N_49989);
or UO_3085 (O_3085,N_49563,N_49596);
nor UO_3086 (O_3086,N_49681,N_49849);
xnor UO_3087 (O_3087,N_49648,N_49513);
or UO_3088 (O_3088,N_49778,N_49909);
nand UO_3089 (O_3089,N_49725,N_49736);
or UO_3090 (O_3090,N_49691,N_49769);
nor UO_3091 (O_3091,N_49815,N_49783);
nand UO_3092 (O_3092,N_49620,N_49534);
and UO_3093 (O_3093,N_49645,N_49561);
nand UO_3094 (O_3094,N_49745,N_49706);
xor UO_3095 (O_3095,N_49545,N_49904);
nor UO_3096 (O_3096,N_49674,N_49569);
nor UO_3097 (O_3097,N_49529,N_49639);
or UO_3098 (O_3098,N_49896,N_49653);
or UO_3099 (O_3099,N_49693,N_49509);
nand UO_3100 (O_3100,N_49825,N_49835);
nor UO_3101 (O_3101,N_49946,N_49752);
nand UO_3102 (O_3102,N_49591,N_49944);
nor UO_3103 (O_3103,N_49980,N_49715);
nor UO_3104 (O_3104,N_49784,N_49725);
xor UO_3105 (O_3105,N_49946,N_49575);
nor UO_3106 (O_3106,N_49853,N_49615);
nor UO_3107 (O_3107,N_49571,N_49591);
nand UO_3108 (O_3108,N_49829,N_49674);
nor UO_3109 (O_3109,N_49529,N_49519);
nor UO_3110 (O_3110,N_49757,N_49874);
xor UO_3111 (O_3111,N_49992,N_49661);
or UO_3112 (O_3112,N_49732,N_49734);
and UO_3113 (O_3113,N_49606,N_49532);
nand UO_3114 (O_3114,N_49765,N_49663);
nor UO_3115 (O_3115,N_49628,N_49696);
nor UO_3116 (O_3116,N_49676,N_49739);
and UO_3117 (O_3117,N_49777,N_49536);
or UO_3118 (O_3118,N_49598,N_49553);
nand UO_3119 (O_3119,N_49560,N_49830);
xnor UO_3120 (O_3120,N_49963,N_49748);
nor UO_3121 (O_3121,N_49698,N_49721);
xor UO_3122 (O_3122,N_49532,N_49977);
xor UO_3123 (O_3123,N_49983,N_49651);
nor UO_3124 (O_3124,N_49595,N_49973);
nor UO_3125 (O_3125,N_49892,N_49579);
xnor UO_3126 (O_3126,N_49844,N_49725);
and UO_3127 (O_3127,N_49716,N_49507);
nor UO_3128 (O_3128,N_49849,N_49705);
nand UO_3129 (O_3129,N_49840,N_49715);
nor UO_3130 (O_3130,N_49806,N_49867);
xnor UO_3131 (O_3131,N_49746,N_49559);
and UO_3132 (O_3132,N_49639,N_49836);
xnor UO_3133 (O_3133,N_49916,N_49713);
nor UO_3134 (O_3134,N_49608,N_49779);
or UO_3135 (O_3135,N_49850,N_49504);
nor UO_3136 (O_3136,N_49520,N_49779);
or UO_3137 (O_3137,N_49775,N_49762);
and UO_3138 (O_3138,N_49695,N_49624);
or UO_3139 (O_3139,N_49615,N_49926);
xor UO_3140 (O_3140,N_49566,N_49910);
and UO_3141 (O_3141,N_49920,N_49870);
xor UO_3142 (O_3142,N_49547,N_49569);
or UO_3143 (O_3143,N_49947,N_49671);
nand UO_3144 (O_3144,N_49828,N_49642);
nand UO_3145 (O_3145,N_49920,N_49997);
or UO_3146 (O_3146,N_49718,N_49561);
or UO_3147 (O_3147,N_49625,N_49708);
nor UO_3148 (O_3148,N_49985,N_49564);
xor UO_3149 (O_3149,N_49798,N_49766);
and UO_3150 (O_3150,N_49652,N_49626);
nand UO_3151 (O_3151,N_49636,N_49997);
nand UO_3152 (O_3152,N_49922,N_49988);
or UO_3153 (O_3153,N_49701,N_49833);
or UO_3154 (O_3154,N_49807,N_49977);
nand UO_3155 (O_3155,N_49835,N_49638);
nor UO_3156 (O_3156,N_49764,N_49982);
nand UO_3157 (O_3157,N_49669,N_49941);
nand UO_3158 (O_3158,N_49818,N_49820);
nand UO_3159 (O_3159,N_49536,N_49972);
nor UO_3160 (O_3160,N_49916,N_49523);
or UO_3161 (O_3161,N_49590,N_49725);
xnor UO_3162 (O_3162,N_49950,N_49594);
nand UO_3163 (O_3163,N_49991,N_49862);
nor UO_3164 (O_3164,N_49941,N_49819);
nand UO_3165 (O_3165,N_49599,N_49791);
or UO_3166 (O_3166,N_49870,N_49903);
or UO_3167 (O_3167,N_49856,N_49887);
nor UO_3168 (O_3168,N_49774,N_49984);
or UO_3169 (O_3169,N_49587,N_49608);
nand UO_3170 (O_3170,N_49995,N_49638);
xnor UO_3171 (O_3171,N_49909,N_49958);
nand UO_3172 (O_3172,N_49992,N_49966);
nor UO_3173 (O_3173,N_49829,N_49904);
nor UO_3174 (O_3174,N_49907,N_49963);
or UO_3175 (O_3175,N_49891,N_49621);
nand UO_3176 (O_3176,N_49984,N_49817);
xnor UO_3177 (O_3177,N_49940,N_49918);
nor UO_3178 (O_3178,N_49624,N_49533);
nor UO_3179 (O_3179,N_49810,N_49859);
nand UO_3180 (O_3180,N_49770,N_49841);
nor UO_3181 (O_3181,N_49715,N_49783);
or UO_3182 (O_3182,N_49602,N_49513);
nand UO_3183 (O_3183,N_49970,N_49611);
and UO_3184 (O_3184,N_49874,N_49721);
and UO_3185 (O_3185,N_49720,N_49512);
nand UO_3186 (O_3186,N_49767,N_49918);
nor UO_3187 (O_3187,N_49956,N_49984);
or UO_3188 (O_3188,N_49824,N_49696);
nor UO_3189 (O_3189,N_49841,N_49858);
xor UO_3190 (O_3190,N_49987,N_49502);
nor UO_3191 (O_3191,N_49966,N_49907);
nor UO_3192 (O_3192,N_49907,N_49651);
or UO_3193 (O_3193,N_49576,N_49895);
nor UO_3194 (O_3194,N_49977,N_49723);
or UO_3195 (O_3195,N_49718,N_49621);
nor UO_3196 (O_3196,N_49826,N_49829);
xor UO_3197 (O_3197,N_49788,N_49553);
nand UO_3198 (O_3198,N_49786,N_49831);
nand UO_3199 (O_3199,N_49837,N_49617);
or UO_3200 (O_3200,N_49741,N_49573);
nor UO_3201 (O_3201,N_49580,N_49596);
xnor UO_3202 (O_3202,N_49501,N_49782);
xnor UO_3203 (O_3203,N_49776,N_49939);
and UO_3204 (O_3204,N_49904,N_49882);
nor UO_3205 (O_3205,N_49721,N_49796);
xor UO_3206 (O_3206,N_49917,N_49834);
or UO_3207 (O_3207,N_49871,N_49599);
and UO_3208 (O_3208,N_49870,N_49816);
xnor UO_3209 (O_3209,N_49980,N_49506);
and UO_3210 (O_3210,N_49571,N_49765);
nand UO_3211 (O_3211,N_49827,N_49746);
nor UO_3212 (O_3212,N_49820,N_49797);
or UO_3213 (O_3213,N_49578,N_49971);
nand UO_3214 (O_3214,N_49576,N_49552);
nand UO_3215 (O_3215,N_49885,N_49869);
nor UO_3216 (O_3216,N_49910,N_49558);
nand UO_3217 (O_3217,N_49538,N_49809);
or UO_3218 (O_3218,N_49641,N_49843);
xnor UO_3219 (O_3219,N_49931,N_49826);
nand UO_3220 (O_3220,N_49567,N_49892);
nor UO_3221 (O_3221,N_49920,N_49536);
or UO_3222 (O_3222,N_49532,N_49555);
xnor UO_3223 (O_3223,N_49575,N_49812);
xor UO_3224 (O_3224,N_49829,N_49726);
xnor UO_3225 (O_3225,N_49598,N_49592);
or UO_3226 (O_3226,N_49920,N_49942);
nor UO_3227 (O_3227,N_49822,N_49968);
nor UO_3228 (O_3228,N_49682,N_49840);
nor UO_3229 (O_3229,N_49961,N_49563);
xnor UO_3230 (O_3230,N_49936,N_49927);
xnor UO_3231 (O_3231,N_49777,N_49922);
or UO_3232 (O_3232,N_49606,N_49971);
nand UO_3233 (O_3233,N_49573,N_49513);
or UO_3234 (O_3234,N_49556,N_49963);
xor UO_3235 (O_3235,N_49916,N_49960);
and UO_3236 (O_3236,N_49961,N_49663);
or UO_3237 (O_3237,N_49502,N_49728);
or UO_3238 (O_3238,N_49912,N_49913);
and UO_3239 (O_3239,N_49620,N_49501);
xnor UO_3240 (O_3240,N_49500,N_49932);
xor UO_3241 (O_3241,N_49660,N_49923);
and UO_3242 (O_3242,N_49618,N_49923);
nor UO_3243 (O_3243,N_49708,N_49847);
xnor UO_3244 (O_3244,N_49755,N_49864);
nand UO_3245 (O_3245,N_49588,N_49870);
and UO_3246 (O_3246,N_49984,N_49546);
nor UO_3247 (O_3247,N_49733,N_49964);
xnor UO_3248 (O_3248,N_49525,N_49616);
nand UO_3249 (O_3249,N_49598,N_49797);
nand UO_3250 (O_3250,N_49716,N_49521);
and UO_3251 (O_3251,N_49504,N_49865);
nand UO_3252 (O_3252,N_49693,N_49872);
nand UO_3253 (O_3253,N_49756,N_49926);
xnor UO_3254 (O_3254,N_49546,N_49583);
or UO_3255 (O_3255,N_49715,N_49505);
xnor UO_3256 (O_3256,N_49716,N_49996);
and UO_3257 (O_3257,N_49584,N_49880);
or UO_3258 (O_3258,N_49590,N_49872);
nor UO_3259 (O_3259,N_49918,N_49978);
and UO_3260 (O_3260,N_49890,N_49948);
xor UO_3261 (O_3261,N_49878,N_49539);
nand UO_3262 (O_3262,N_49666,N_49858);
nand UO_3263 (O_3263,N_49789,N_49620);
and UO_3264 (O_3264,N_49592,N_49705);
nand UO_3265 (O_3265,N_49620,N_49628);
nor UO_3266 (O_3266,N_49630,N_49999);
nor UO_3267 (O_3267,N_49998,N_49949);
nor UO_3268 (O_3268,N_49901,N_49609);
and UO_3269 (O_3269,N_49728,N_49760);
and UO_3270 (O_3270,N_49583,N_49968);
nand UO_3271 (O_3271,N_49603,N_49669);
and UO_3272 (O_3272,N_49814,N_49779);
nand UO_3273 (O_3273,N_49523,N_49980);
nand UO_3274 (O_3274,N_49745,N_49616);
xnor UO_3275 (O_3275,N_49759,N_49608);
nor UO_3276 (O_3276,N_49978,N_49912);
nand UO_3277 (O_3277,N_49743,N_49973);
or UO_3278 (O_3278,N_49926,N_49768);
or UO_3279 (O_3279,N_49566,N_49598);
and UO_3280 (O_3280,N_49697,N_49814);
and UO_3281 (O_3281,N_49506,N_49657);
and UO_3282 (O_3282,N_49567,N_49875);
xnor UO_3283 (O_3283,N_49757,N_49677);
nand UO_3284 (O_3284,N_49941,N_49799);
xnor UO_3285 (O_3285,N_49583,N_49630);
nor UO_3286 (O_3286,N_49869,N_49728);
xnor UO_3287 (O_3287,N_49982,N_49643);
nand UO_3288 (O_3288,N_49913,N_49825);
or UO_3289 (O_3289,N_49831,N_49750);
xor UO_3290 (O_3290,N_49858,N_49864);
or UO_3291 (O_3291,N_49659,N_49599);
or UO_3292 (O_3292,N_49875,N_49781);
and UO_3293 (O_3293,N_49556,N_49832);
or UO_3294 (O_3294,N_49653,N_49670);
nor UO_3295 (O_3295,N_49973,N_49739);
xor UO_3296 (O_3296,N_49750,N_49722);
xor UO_3297 (O_3297,N_49522,N_49797);
xor UO_3298 (O_3298,N_49583,N_49588);
or UO_3299 (O_3299,N_49817,N_49693);
xor UO_3300 (O_3300,N_49733,N_49912);
nor UO_3301 (O_3301,N_49913,N_49675);
nor UO_3302 (O_3302,N_49934,N_49860);
nor UO_3303 (O_3303,N_49985,N_49898);
and UO_3304 (O_3304,N_49555,N_49741);
xnor UO_3305 (O_3305,N_49517,N_49701);
and UO_3306 (O_3306,N_49526,N_49792);
or UO_3307 (O_3307,N_49895,N_49561);
or UO_3308 (O_3308,N_49701,N_49768);
xor UO_3309 (O_3309,N_49786,N_49573);
nand UO_3310 (O_3310,N_49517,N_49784);
xor UO_3311 (O_3311,N_49609,N_49825);
or UO_3312 (O_3312,N_49526,N_49506);
nand UO_3313 (O_3313,N_49859,N_49580);
and UO_3314 (O_3314,N_49978,N_49941);
nor UO_3315 (O_3315,N_49940,N_49789);
or UO_3316 (O_3316,N_49520,N_49792);
nor UO_3317 (O_3317,N_49763,N_49940);
and UO_3318 (O_3318,N_49835,N_49855);
xnor UO_3319 (O_3319,N_49856,N_49596);
xor UO_3320 (O_3320,N_49940,N_49678);
nand UO_3321 (O_3321,N_49656,N_49788);
or UO_3322 (O_3322,N_49923,N_49752);
nor UO_3323 (O_3323,N_49562,N_49512);
and UO_3324 (O_3324,N_49823,N_49854);
nor UO_3325 (O_3325,N_49867,N_49561);
or UO_3326 (O_3326,N_49693,N_49979);
and UO_3327 (O_3327,N_49724,N_49989);
and UO_3328 (O_3328,N_49731,N_49999);
xnor UO_3329 (O_3329,N_49675,N_49985);
or UO_3330 (O_3330,N_49922,N_49941);
nor UO_3331 (O_3331,N_49569,N_49848);
and UO_3332 (O_3332,N_49915,N_49721);
nand UO_3333 (O_3333,N_49893,N_49558);
or UO_3334 (O_3334,N_49759,N_49594);
nand UO_3335 (O_3335,N_49812,N_49910);
xor UO_3336 (O_3336,N_49574,N_49579);
nor UO_3337 (O_3337,N_49571,N_49942);
and UO_3338 (O_3338,N_49715,N_49901);
and UO_3339 (O_3339,N_49929,N_49931);
nor UO_3340 (O_3340,N_49577,N_49846);
and UO_3341 (O_3341,N_49602,N_49617);
xor UO_3342 (O_3342,N_49886,N_49740);
nand UO_3343 (O_3343,N_49684,N_49513);
or UO_3344 (O_3344,N_49699,N_49751);
or UO_3345 (O_3345,N_49547,N_49986);
nor UO_3346 (O_3346,N_49856,N_49905);
xor UO_3347 (O_3347,N_49801,N_49809);
xor UO_3348 (O_3348,N_49977,N_49628);
nand UO_3349 (O_3349,N_49901,N_49946);
or UO_3350 (O_3350,N_49785,N_49835);
xor UO_3351 (O_3351,N_49912,N_49946);
and UO_3352 (O_3352,N_49694,N_49906);
nor UO_3353 (O_3353,N_49507,N_49896);
nand UO_3354 (O_3354,N_49784,N_49954);
or UO_3355 (O_3355,N_49965,N_49810);
or UO_3356 (O_3356,N_49774,N_49532);
nor UO_3357 (O_3357,N_49988,N_49918);
or UO_3358 (O_3358,N_49886,N_49547);
nor UO_3359 (O_3359,N_49686,N_49951);
and UO_3360 (O_3360,N_49815,N_49548);
nand UO_3361 (O_3361,N_49562,N_49726);
nand UO_3362 (O_3362,N_49568,N_49844);
or UO_3363 (O_3363,N_49876,N_49657);
xnor UO_3364 (O_3364,N_49888,N_49685);
or UO_3365 (O_3365,N_49716,N_49578);
and UO_3366 (O_3366,N_49668,N_49804);
xor UO_3367 (O_3367,N_49998,N_49635);
nor UO_3368 (O_3368,N_49768,N_49769);
xor UO_3369 (O_3369,N_49605,N_49609);
xnor UO_3370 (O_3370,N_49954,N_49817);
nor UO_3371 (O_3371,N_49640,N_49770);
xor UO_3372 (O_3372,N_49563,N_49950);
and UO_3373 (O_3373,N_49667,N_49786);
and UO_3374 (O_3374,N_49567,N_49876);
or UO_3375 (O_3375,N_49927,N_49885);
or UO_3376 (O_3376,N_49786,N_49898);
nand UO_3377 (O_3377,N_49970,N_49881);
or UO_3378 (O_3378,N_49664,N_49952);
xor UO_3379 (O_3379,N_49914,N_49782);
xnor UO_3380 (O_3380,N_49547,N_49545);
nand UO_3381 (O_3381,N_49691,N_49901);
or UO_3382 (O_3382,N_49965,N_49969);
nand UO_3383 (O_3383,N_49575,N_49655);
and UO_3384 (O_3384,N_49628,N_49911);
nand UO_3385 (O_3385,N_49536,N_49604);
or UO_3386 (O_3386,N_49952,N_49936);
nor UO_3387 (O_3387,N_49753,N_49588);
nand UO_3388 (O_3388,N_49828,N_49802);
or UO_3389 (O_3389,N_49835,N_49809);
and UO_3390 (O_3390,N_49620,N_49573);
xnor UO_3391 (O_3391,N_49515,N_49683);
or UO_3392 (O_3392,N_49923,N_49840);
and UO_3393 (O_3393,N_49594,N_49687);
nand UO_3394 (O_3394,N_49547,N_49521);
and UO_3395 (O_3395,N_49554,N_49635);
or UO_3396 (O_3396,N_49728,N_49618);
xnor UO_3397 (O_3397,N_49658,N_49640);
and UO_3398 (O_3398,N_49587,N_49948);
xnor UO_3399 (O_3399,N_49879,N_49763);
or UO_3400 (O_3400,N_49613,N_49833);
nor UO_3401 (O_3401,N_49867,N_49899);
nor UO_3402 (O_3402,N_49697,N_49844);
nand UO_3403 (O_3403,N_49963,N_49611);
xnor UO_3404 (O_3404,N_49930,N_49853);
nor UO_3405 (O_3405,N_49634,N_49579);
nand UO_3406 (O_3406,N_49753,N_49507);
nand UO_3407 (O_3407,N_49789,N_49937);
nand UO_3408 (O_3408,N_49847,N_49531);
or UO_3409 (O_3409,N_49986,N_49777);
nor UO_3410 (O_3410,N_49613,N_49500);
nor UO_3411 (O_3411,N_49745,N_49947);
xnor UO_3412 (O_3412,N_49836,N_49694);
nand UO_3413 (O_3413,N_49770,N_49886);
and UO_3414 (O_3414,N_49826,N_49771);
xnor UO_3415 (O_3415,N_49859,N_49769);
nand UO_3416 (O_3416,N_49834,N_49823);
nor UO_3417 (O_3417,N_49890,N_49828);
and UO_3418 (O_3418,N_49994,N_49787);
xor UO_3419 (O_3419,N_49653,N_49936);
xnor UO_3420 (O_3420,N_49819,N_49744);
nor UO_3421 (O_3421,N_49505,N_49758);
or UO_3422 (O_3422,N_49514,N_49922);
xor UO_3423 (O_3423,N_49593,N_49666);
xor UO_3424 (O_3424,N_49827,N_49689);
nand UO_3425 (O_3425,N_49960,N_49596);
nand UO_3426 (O_3426,N_49599,N_49519);
and UO_3427 (O_3427,N_49664,N_49588);
nor UO_3428 (O_3428,N_49923,N_49895);
nor UO_3429 (O_3429,N_49752,N_49733);
nand UO_3430 (O_3430,N_49615,N_49953);
nor UO_3431 (O_3431,N_49763,N_49637);
or UO_3432 (O_3432,N_49723,N_49815);
nand UO_3433 (O_3433,N_49926,N_49893);
nand UO_3434 (O_3434,N_49514,N_49938);
and UO_3435 (O_3435,N_49724,N_49607);
nor UO_3436 (O_3436,N_49858,N_49660);
and UO_3437 (O_3437,N_49572,N_49573);
and UO_3438 (O_3438,N_49959,N_49579);
and UO_3439 (O_3439,N_49911,N_49808);
and UO_3440 (O_3440,N_49770,N_49998);
nor UO_3441 (O_3441,N_49890,N_49781);
nand UO_3442 (O_3442,N_49519,N_49576);
and UO_3443 (O_3443,N_49858,N_49646);
xnor UO_3444 (O_3444,N_49955,N_49996);
or UO_3445 (O_3445,N_49916,N_49694);
nor UO_3446 (O_3446,N_49543,N_49990);
nand UO_3447 (O_3447,N_49710,N_49898);
xor UO_3448 (O_3448,N_49931,N_49750);
and UO_3449 (O_3449,N_49750,N_49839);
nand UO_3450 (O_3450,N_49797,N_49637);
and UO_3451 (O_3451,N_49690,N_49871);
or UO_3452 (O_3452,N_49819,N_49893);
nand UO_3453 (O_3453,N_49773,N_49631);
and UO_3454 (O_3454,N_49520,N_49937);
or UO_3455 (O_3455,N_49606,N_49826);
nor UO_3456 (O_3456,N_49828,N_49955);
nor UO_3457 (O_3457,N_49553,N_49872);
nor UO_3458 (O_3458,N_49890,N_49737);
xor UO_3459 (O_3459,N_49567,N_49984);
nand UO_3460 (O_3460,N_49654,N_49649);
nor UO_3461 (O_3461,N_49514,N_49580);
xnor UO_3462 (O_3462,N_49946,N_49738);
xor UO_3463 (O_3463,N_49572,N_49520);
nand UO_3464 (O_3464,N_49664,N_49973);
or UO_3465 (O_3465,N_49855,N_49938);
nand UO_3466 (O_3466,N_49864,N_49788);
nor UO_3467 (O_3467,N_49913,N_49961);
nand UO_3468 (O_3468,N_49709,N_49958);
xnor UO_3469 (O_3469,N_49859,N_49928);
nor UO_3470 (O_3470,N_49904,N_49510);
or UO_3471 (O_3471,N_49934,N_49664);
xor UO_3472 (O_3472,N_49643,N_49854);
or UO_3473 (O_3473,N_49878,N_49812);
xor UO_3474 (O_3474,N_49827,N_49594);
and UO_3475 (O_3475,N_49525,N_49511);
nor UO_3476 (O_3476,N_49642,N_49707);
or UO_3477 (O_3477,N_49552,N_49578);
nand UO_3478 (O_3478,N_49784,N_49503);
nor UO_3479 (O_3479,N_49630,N_49636);
and UO_3480 (O_3480,N_49648,N_49635);
xnor UO_3481 (O_3481,N_49684,N_49547);
nor UO_3482 (O_3482,N_49623,N_49779);
xor UO_3483 (O_3483,N_49942,N_49992);
xnor UO_3484 (O_3484,N_49704,N_49907);
or UO_3485 (O_3485,N_49647,N_49738);
xor UO_3486 (O_3486,N_49775,N_49779);
or UO_3487 (O_3487,N_49757,N_49594);
nor UO_3488 (O_3488,N_49871,N_49851);
nand UO_3489 (O_3489,N_49687,N_49753);
and UO_3490 (O_3490,N_49740,N_49805);
nand UO_3491 (O_3491,N_49751,N_49810);
xor UO_3492 (O_3492,N_49580,N_49702);
and UO_3493 (O_3493,N_49866,N_49743);
and UO_3494 (O_3494,N_49694,N_49731);
or UO_3495 (O_3495,N_49636,N_49542);
or UO_3496 (O_3496,N_49747,N_49528);
nor UO_3497 (O_3497,N_49986,N_49740);
nor UO_3498 (O_3498,N_49923,N_49797);
or UO_3499 (O_3499,N_49859,N_49648);
and UO_3500 (O_3500,N_49749,N_49554);
nand UO_3501 (O_3501,N_49791,N_49574);
nor UO_3502 (O_3502,N_49726,N_49817);
xor UO_3503 (O_3503,N_49940,N_49890);
or UO_3504 (O_3504,N_49822,N_49943);
nand UO_3505 (O_3505,N_49616,N_49956);
xnor UO_3506 (O_3506,N_49688,N_49980);
xor UO_3507 (O_3507,N_49572,N_49818);
nor UO_3508 (O_3508,N_49809,N_49739);
nand UO_3509 (O_3509,N_49649,N_49616);
or UO_3510 (O_3510,N_49601,N_49527);
or UO_3511 (O_3511,N_49924,N_49518);
nor UO_3512 (O_3512,N_49727,N_49997);
or UO_3513 (O_3513,N_49867,N_49840);
xor UO_3514 (O_3514,N_49557,N_49809);
or UO_3515 (O_3515,N_49983,N_49514);
xnor UO_3516 (O_3516,N_49694,N_49584);
xnor UO_3517 (O_3517,N_49739,N_49504);
and UO_3518 (O_3518,N_49592,N_49977);
and UO_3519 (O_3519,N_49837,N_49924);
xor UO_3520 (O_3520,N_49768,N_49534);
and UO_3521 (O_3521,N_49572,N_49765);
or UO_3522 (O_3522,N_49851,N_49630);
nor UO_3523 (O_3523,N_49616,N_49571);
and UO_3524 (O_3524,N_49648,N_49651);
or UO_3525 (O_3525,N_49978,N_49892);
nand UO_3526 (O_3526,N_49823,N_49970);
nand UO_3527 (O_3527,N_49983,N_49878);
or UO_3528 (O_3528,N_49526,N_49527);
nor UO_3529 (O_3529,N_49634,N_49533);
nand UO_3530 (O_3530,N_49710,N_49934);
xor UO_3531 (O_3531,N_49763,N_49709);
or UO_3532 (O_3532,N_49638,N_49525);
nor UO_3533 (O_3533,N_49885,N_49818);
xor UO_3534 (O_3534,N_49897,N_49820);
nor UO_3535 (O_3535,N_49678,N_49632);
nand UO_3536 (O_3536,N_49703,N_49845);
nor UO_3537 (O_3537,N_49774,N_49906);
and UO_3538 (O_3538,N_49910,N_49621);
nand UO_3539 (O_3539,N_49631,N_49765);
xor UO_3540 (O_3540,N_49986,N_49605);
nor UO_3541 (O_3541,N_49587,N_49978);
nand UO_3542 (O_3542,N_49954,N_49983);
nand UO_3543 (O_3543,N_49916,N_49765);
xor UO_3544 (O_3544,N_49880,N_49815);
nand UO_3545 (O_3545,N_49927,N_49979);
xnor UO_3546 (O_3546,N_49676,N_49746);
xor UO_3547 (O_3547,N_49884,N_49826);
and UO_3548 (O_3548,N_49712,N_49524);
and UO_3549 (O_3549,N_49939,N_49623);
and UO_3550 (O_3550,N_49622,N_49973);
or UO_3551 (O_3551,N_49721,N_49761);
xnor UO_3552 (O_3552,N_49559,N_49635);
and UO_3553 (O_3553,N_49966,N_49726);
xnor UO_3554 (O_3554,N_49822,N_49509);
nand UO_3555 (O_3555,N_49665,N_49670);
nor UO_3556 (O_3556,N_49636,N_49514);
nor UO_3557 (O_3557,N_49574,N_49979);
or UO_3558 (O_3558,N_49690,N_49905);
nor UO_3559 (O_3559,N_49912,N_49823);
or UO_3560 (O_3560,N_49770,N_49847);
xor UO_3561 (O_3561,N_49745,N_49700);
and UO_3562 (O_3562,N_49634,N_49767);
and UO_3563 (O_3563,N_49917,N_49518);
and UO_3564 (O_3564,N_49557,N_49800);
xnor UO_3565 (O_3565,N_49873,N_49678);
and UO_3566 (O_3566,N_49813,N_49929);
nand UO_3567 (O_3567,N_49953,N_49600);
or UO_3568 (O_3568,N_49682,N_49757);
and UO_3569 (O_3569,N_49737,N_49757);
and UO_3570 (O_3570,N_49976,N_49559);
or UO_3571 (O_3571,N_49551,N_49856);
and UO_3572 (O_3572,N_49625,N_49512);
and UO_3573 (O_3573,N_49783,N_49898);
and UO_3574 (O_3574,N_49561,N_49640);
and UO_3575 (O_3575,N_49954,N_49720);
xnor UO_3576 (O_3576,N_49595,N_49628);
nand UO_3577 (O_3577,N_49962,N_49727);
and UO_3578 (O_3578,N_49883,N_49650);
xnor UO_3579 (O_3579,N_49903,N_49897);
xor UO_3580 (O_3580,N_49755,N_49729);
or UO_3581 (O_3581,N_49996,N_49627);
nand UO_3582 (O_3582,N_49608,N_49874);
nand UO_3583 (O_3583,N_49860,N_49578);
and UO_3584 (O_3584,N_49792,N_49550);
nor UO_3585 (O_3585,N_49720,N_49857);
and UO_3586 (O_3586,N_49617,N_49526);
and UO_3587 (O_3587,N_49539,N_49685);
and UO_3588 (O_3588,N_49831,N_49756);
and UO_3589 (O_3589,N_49538,N_49754);
and UO_3590 (O_3590,N_49942,N_49530);
or UO_3591 (O_3591,N_49922,N_49878);
nor UO_3592 (O_3592,N_49805,N_49693);
and UO_3593 (O_3593,N_49510,N_49625);
or UO_3594 (O_3594,N_49649,N_49783);
or UO_3595 (O_3595,N_49643,N_49703);
or UO_3596 (O_3596,N_49713,N_49599);
or UO_3597 (O_3597,N_49925,N_49813);
or UO_3598 (O_3598,N_49591,N_49882);
xnor UO_3599 (O_3599,N_49962,N_49807);
nor UO_3600 (O_3600,N_49649,N_49890);
or UO_3601 (O_3601,N_49836,N_49577);
nor UO_3602 (O_3602,N_49955,N_49838);
and UO_3603 (O_3603,N_49935,N_49685);
or UO_3604 (O_3604,N_49615,N_49617);
nor UO_3605 (O_3605,N_49867,N_49578);
nand UO_3606 (O_3606,N_49757,N_49692);
and UO_3607 (O_3607,N_49686,N_49950);
xor UO_3608 (O_3608,N_49936,N_49647);
xnor UO_3609 (O_3609,N_49929,N_49573);
nor UO_3610 (O_3610,N_49929,N_49787);
or UO_3611 (O_3611,N_49834,N_49670);
nor UO_3612 (O_3612,N_49892,N_49677);
and UO_3613 (O_3613,N_49932,N_49729);
nor UO_3614 (O_3614,N_49952,N_49641);
nor UO_3615 (O_3615,N_49503,N_49898);
nor UO_3616 (O_3616,N_49722,N_49531);
and UO_3617 (O_3617,N_49891,N_49792);
or UO_3618 (O_3618,N_49918,N_49877);
or UO_3619 (O_3619,N_49586,N_49787);
xnor UO_3620 (O_3620,N_49545,N_49702);
xor UO_3621 (O_3621,N_49972,N_49586);
nand UO_3622 (O_3622,N_49720,N_49991);
nand UO_3623 (O_3623,N_49578,N_49682);
nand UO_3624 (O_3624,N_49895,N_49621);
nor UO_3625 (O_3625,N_49625,N_49515);
nand UO_3626 (O_3626,N_49819,N_49988);
nand UO_3627 (O_3627,N_49920,N_49701);
xnor UO_3628 (O_3628,N_49945,N_49541);
nand UO_3629 (O_3629,N_49722,N_49645);
nand UO_3630 (O_3630,N_49790,N_49741);
and UO_3631 (O_3631,N_49754,N_49782);
nand UO_3632 (O_3632,N_49959,N_49769);
nand UO_3633 (O_3633,N_49756,N_49580);
nor UO_3634 (O_3634,N_49716,N_49872);
nor UO_3635 (O_3635,N_49849,N_49892);
or UO_3636 (O_3636,N_49790,N_49869);
nor UO_3637 (O_3637,N_49564,N_49542);
and UO_3638 (O_3638,N_49710,N_49858);
and UO_3639 (O_3639,N_49597,N_49531);
xor UO_3640 (O_3640,N_49599,N_49680);
and UO_3641 (O_3641,N_49693,N_49680);
or UO_3642 (O_3642,N_49576,N_49790);
xnor UO_3643 (O_3643,N_49962,N_49898);
or UO_3644 (O_3644,N_49598,N_49935);
or UO_3645 (O_3645,N_49840,N_49808);
and UO_3646 (O_3646,N_49847,N_49935);
and UO_3647 (O_3647,N_49915,N_49813);
nand UO_3648 (O_3648,N_49737,N_49638);
or UO_3649 (O_3649,N_49665,N_49716);
nor UO_3650 (O_3650,N_49734,N_49999);
or UO_3651 (O_3651,N_49637,N_49794);
or UO_3652 (O_3652,N_49514,N_49897);
and UO_3653 (O_3653,N_49639,N_49867);
xnor UO_3654 (O_3654,N_49975,N_49560);
and UO_3655 (O_3655,N_49749,N_49881);
and UO_3656 (O_3656,N_49656,N_49941);
or UO_3657 (O_3657,N_49561,N_49932);
and UO_3658 (O_3658,N_49533,N_49945);
xor UO_3659 (O_3659,N_49625,N_49799);
and UO_3660 (O_3660,N_49900,N_49809);
nand UO_3661 (O_3661,N_49691,N_49821);
nand UO_3662 (O_3662,N_49833,N_49944);
or UO_3663 (O_3663,N_49896,N_49552);
or UO_3664 (O_3664,N_49871,N_49591);
and UO_3665 (O_3665,N_49712,N_49509);
xnor UO_3666 (O_3666,N_49916,N_49710);
nor UO_3667 (O_3667,N_49795,N_49551);
or UO_3668 (O_3668,N_49889,N_49838);
nand UO_3669 (O_3669,N_49579,N_49687);
nand UO_3670 (O_3670,N_49542,N_49652);
nor UO_3671 (O_3671,N_49560,N_49778);
xor UO_3672 (O_3672,N_49680,N_49855);
and UO_3673 (O_3673,N_49957,N_49847);
or UO_3674 (O_3674,N_49985,N_49618);
and UO_3675 (O_3675,N_49935,N_49828);
nor UO_3676 (O_3676,N_49513,N_49765);
nor UO_3677 (O_3677,N_49928,N_49679);
nor UO_3678 (O_3678,N_49963,N_49826);
nand UO_3679 (O_3679,N_49842,N_49804);
and UO_3680 (O_3680,N_49940,N_49799);
xnor UO_3681 (O_3681,N_49939,N_49790);
or UO_3682 (O_3682,N_49754,N_49642);
nand UO_3683 (O_3683,N_49791,N_49757);
nand UO_3684 (O_3684,N_49531,N_49552);
xor UO_3685 (O_3685,N_49997,N_49578);
nor UO_3686 (O_3686,N_49624,N_49876);
nand UO_3687 (O_3687,N_49579,N_49899);
xor UO_3688 (O_3688,N_49857,N_49580);
or UO_3689 (O_3689,N_49540,N_49900);
and UO_3690 (O_3690,N_49537,N_49949);
nand UO_3691 (O_3691,N_49598,N_49638);
xor UO_3692 (O_3692,N_49743,N_49939);
nand UO_3693 (O_3693,N_49724,N_49561);
or UO_3694 (O_3694,N_49664,N_49645);
xor UO_3695 (O_3695,N_49873,N_49592);
nand UO_3696 (O_3696,N_49534,N_49863);
xor UO_3697 (O_3697,N_49888,N_49833);
and UO_3698 (O_3698,N_49800,N_49756);
and UO_3699 (O_3699,N_49663,N_49741);
nand UO_3700 (O_3700,N_49933,N_49929);
xor UO_3701 (O_3701,N_49814,N_49956);
or UO_3702 (O_3702,N_49817,N_49573);
xnor UO_3703 (O_3703,N_49693,N_49774);
nand UO_3704 (O_3704,N_49584,N_49560);
or UO_3705 (O_3705,N_49947,N_49906);
and UO_3706 (O_3706,N_49906,N_49802);
nand UO_3707 (O_3707,N_49921,N_49532);
nor UO_3708 (O_3708,N_49958,N_49981);
xor UO_3709 (O_3709,N_49992,N_49765);
or UO_3710 (O_3710,N_49604,N_49719);
and UO_3711 (O_3711,N_49875,N_49729);
nand UO_3712 (O_3712,N_49688,N_49886);
nand UO_3713 (O_3713,N_49977,N_49908);
nor UO_3714 (O_3714,N_49983,N_49871);
nand UO_3715 (O_3715,N_49699,N_49667);
nand UO_3716 (O_3716,N_49963,N_49593);
nor UO_3717 (O_3717,N_49877,N_49833);
and UO_3718 (O_3718,N_49845,N_49839);
and UO_3719 (O_3719,N_49914,N_49584);
nand UO_3720 (O_3720,N_49902,N_49956);
nor UO_3721 (O_3721,N_49599,N_49622);
nand UO_3722 (O_3722,N_49803,N_49788);
and UO_3723 (O_3723,N_49737,N_49664);
xnor UO_3724 (O_3724,N_49940,N_49865);
nand UO_3725 (O_3725,N_49525,N_49722);
and UO_3726 (O_3726,N_49914,N_49910);
xnor UO_3727 (O_3727,N_49636,N_49973);
xnor UO_3728 (O_3728,N_49606,N_49957);
and UO_3729 (O_3729,N_49507,N_49571);
nor UO_3730 (O_3730,N_49539,N_49628);
or UO_3731 (O_3731,N_49700,N_49843);
nand UO_3732 (O_3732,N_49928,N_49706);
nor UO_3733 (O_3733,N_49542,N_49506);
nand UO_3734 (O_3734,N_49857,N_49799);
nand UO_3735 (O_3735,N_49715,N_49674);
and UO_3736 (O_3736,N_49561,N_49958);
nand UO_3737 (O_3737,N_49856,N_49803);
nor UO_3738 (O_3738,N_49801,N_49509);
nand UO_3739 (O_3739,N_49684,N_49676);
xnor UO_3740 (O_3740,N_49738,N_49547);
or UO_3741 (O_3741,N_49728,N_49596);
xnor UO_3742 (O_3742,N_49721,N_49819);
nor UO_3743 (O_3743,N_49802,N_49952);
or UO_3744 (O_3744,N_49986,N_49990);
xnor UO_3745 (O_3745,N_49662,N_49657);
xnor UO_3746 (O_3746,N_49577,N_49583);
and UO_3747 (O_3747,N_49641,N_49591);
nand UO_3748 (O_3748,N_49608,N_49586);
nor UO_3749 (O_3749,N_49680,N_49617);
nand UO_3750 (O_3750,N_49622,N_49838);
nor UO_3751 (O_3751,N_49586,N_49859);
or UO_3752 (O_3752,N_49640,N_49977);
xor UO_3753 (O_3753,N_49728,N_49976);
xnor UO_3754 (O_3754,N_49698,N_49760);
or UO_3755 (O_3755,N_49627,N_49598);
nand UO_3756 (O_3756,N_49503,N_49729);
xnor UO_3757 (O_3757,N_49674,N_49739);
and UO_3758 (O_3758,N_49657,N_49931);
xnor UO_3759 (O_3759,N_49676,N_49599);
nor UO_3760 (O_3760,N_49676,N_49504);
or UO_3761 (O_3761,N_49524,N_49514);
or UO_3762 (O_3762,N_49688,N_49957);
nand UO_3763 (O_3763,N_49811,N_49952);
nand UO_3764 (O_3764,N_49715,N_49693);
nor UO_3765 (O_3765,N_49942,N_49729);
and UO_3766 (O_3766,N_49922,N_49950);
and UO_3767 (O_3767,N_49762,N_49820);
or UO_3768 (O_3768,N_49526,N_49974);
and UO_3769 (O_3769,N_49682,N_49826);
nor UO_3770 (O_3770,N_49716,N_49688);
xor UO_3771 (O_3771,N_49549,N_49979);
and UO_3772 (O_3772,N_49875,N_49836);
xnor UO_3773 (O_3773,N_49686,N_49824);
nor UO_3774 (O_3774,N_49743,N_49687);
or UO_3775 (O_3775,N_49977,N_49985);
or UO_3776 (O_3776,N_49676,N_49927);
nor UO_3777 (O_3777,N_49546,N_49731);
and UO_3778 (O_3778,N_49955,N_49686);
nand UO_3779 (O_3779,N_49891,N_49994);
nand UO_3780 (O_3780,N_49674,N_49546);
and UO_3781 (O_3781,N_49617,N_49809);
nand UO_3782 (O_3782,N_49544,N_49775);
and UO_3783 (O_3783,N_49753,N_49761);
and UO_3784 (O_3784,N_49524,N_49963);
or UO_3785 (O_3785,N_49620,N_49673);
or UO_3786 (O_3786,N_49940,N_49585);
nand UO_3787 (O_3787,N_49829,N_49922);
and UO_3788 (O_3788,N_49736,N_49592);
xor UO_3789 (O_3789,N_49552,N_49668);
xnor UO_3790 (O_3790,N_49909,N_49927);
nand UO_3791 (O_3791,N_49884,N_49935);
xor UO_3792 (O_3792,N_49724,N_49811);
nor UO_3793 (O_3793,N_49898,N_49674);
nor UO_3794 (O_3794,N_49776,N_49782);
nor UO_3795 (O_3795,N_49652,N_49611);
and UO_3796 (O_3796,N_49675,N_49543);
or UO_3797 (O_3797,N_49877,N_49813);
and UO_3798 (O_3798,N_49609,N_49742);
xor UO_3799 (O_3799,N_49923,N_49832);
and UO_3800 (O_3800,N_49929,N_49952);
or UO_3801 (O_3801,N_49560,N_49703);
or UO_3802 (O_3802,N_49663,N_49510);
xnor UO_3803 (O_3803,N_49645,N_49751);
and UO_3804 (O_3804,N_49865,N_49959);
xnor UO_3805 (O_3805,N_49632,N_49973);
and UO_3806 (O_3806,N_49597,N_49561);
and UO_3807 (O_3807,N_49909,N_49640);
or UO_3808 (O_3808,N_49900,N_49830);
or UO_3809 (O_3809,N_49975,N_49535);
nor UO_3810 (O_3810,N_49907,N_49918);
or UO_3811 (O_3811,N_49652,N_49855);
nand UO_3812 (O_3812,N_49647,N_49779);
or UO_3813 (O_3813,N_49725,N_49620);
nand UO_3814 (O_3814,N_49954,N_49992);
xor UO_3815 (O_3815,N_49584,N_49902);
nand UO_3816 (O_3816,N_49749,N_49944);
and UO_3817 (O_3817,N_49764,N_49517);
nor UO_3818 (O_3818,N_49604,N_49784);
and UO_3819 (O_3819,N_49867,N_49879);
xnor UO_3820 (O_3820,N_49838,N_49509);
or UO_3821 (O_3821,N_49659,N_49984);
xor UO_3822 (O_3822,N_49545,N_49760);
xnor UO_3823 (O_3823,N_49954,N_49873);
xor UO_3824 (O_3824,N_49571,N_49659);
or UO_3825 (O_3825,N_49830,N_49597);
nor UO_3826 (O_3826,N_49654,N_49600);
nand UO_3827 (O_3827,N_49619,N_49526);
and UO_3828 (O_3828,N_49658,N_49667);
nor UO_3829 (O_3829,N_49566,N_49567);
or UO_3830 (O_3830,N_49762,N_49597);
and UO_3831 (O_3831,N_49593,N_49682);
and UO_3832 (O_3832,N_49742,N_49921);
or UO_3833 (O_3833,N_49916,N_49993);
nor UO_3834 (O_3834,N_49982,N_49933);
xor UO_3835 (O_3835,N_49625,N_49870);
nor UO_3836 (O_3836,N_49596,N_49561);
nor UO_3837 (O_3837,N_49552,N_49832);
and UO_3838 (O_3838,N_49844,N_49577);
nor UO_3839 (O_3839,N_49864,N_49694);
xor UO_3840 (O_3840,N_49740,N_49546);
xnor UO_3841 (O_3841,N_49732,N_49777);
or UO_3842 (O_3842,N_49571,N_49891);
and UO_3843 (O_3843,N_49895,N_49676);
xnor UO_3844 (O_3844,N_49510,N_49628);
nand UO_3845 (O_3845,N_49858,N_49742);
or UO_3846 (O_3846,N_49651,N_49776);
nand UO_3847 (O_3847,N_49931,N_49920);
or UO_3848 (O_3848,N_49793,N_49631);
nand UO_3849 (O_3849,N_49654,N_49826);
nor UO_3850 (O_3850,N_49554,N_49863);
xor UO_3851 (O_3851,N_49895,N_49656);
nand UO_3852 (O_3852,N_49576,N_49852);
nor UO_3853 (O_3853,N_49909,N_49575);
xnor UO_3854 (O_3854,N_49728,N_49601);
and UO_3855 (O_3855,N_49538,N_49600);
or UO_3856 (O_3856,N_49939,N_49914);
nor UO_3857 (O_3857,N_49733,N_49654);
or UO_3858 (O_3858,N_49785,N_49508);
nand UO_3859 (O_3859,N_49931,N_49626);
or UO_3860 (O_3860,N_49808,N_49884);
and UO_3861 (O_3861,N_49757,N_49544);
and UO_3862 (O_3862,N_49953,N_49755);
nor UO_3863 (O_3863,N_49700,N_49707);
and UO_3864 (O_3864,N_49850,N_49906);
xnor UO_3865 (O_3865,N_49841,N_49624);
nand UO_3866 (O_3866,N_49576,N_49714);
and UO_3867 (O_3867,N_49916,N_49759);
nor UO_3868 (O_3868,N_49682,N_49971);
or UO_3869 (O_3869,N_49711,N_49812);
nor UO_3870 (O_3870,N_49507,N_49787);
xnor UO_3871 (O_3871,N_49602,N_49550);
and UO_3872 (O_3872,N_49821,N_49807);
or UO_3873 (O_3873,N_49675,N_49925);
and UO_3874 (O_3874,N_49536,N_49533);
nor UO_3875 (O_3875,N_49942,N_49891);
and UO_3876 (O_3876,N_49939,N_49515);
and UO_3877 (O_3877,N_49558,N_49971);
nor UO_3878 (O_3878,N_49529,N_49884);
or UO_3879 (O_3879,N_49879,N_49715);
and UO_3880 (O_3880,N_49755,N_49690);
and UO_3881 (O_3881,N_49753,N_49795);
and UO_3882 (O_3882,N_49751,N_49778);
and UO_3883 (O_3883,N_49784,N_49982);
nand UO_3884 (O_3884,N_49677,N_49747);
nand UO_3885 (O_3885,N_49963,N_49779);
nand UO_3886 (O_3886,N_49601,N_49949);
xor UO_3887 (O_3887,N_49974,N_49985);
xor UO_3888 (O_3888,N_49964,N_49833);
nor UO_3889 (O_3889,N_49632,N_49845);
xor UO_3890 (O_3890,N_49831,N_49633);
xnor UO_3891 (O_3891,N_49814,N_49853);
or UO_3892 (O_3892,N_49796,N_49822);
and UO_3893 (O_3893,N_49997,N_49913);
or UO_3894 (O_3894,N_49761,N_49556);
xor UO_3895 (O_3895,N_49932,N_49990);
xor UO_3896 (O_3896,N_49537,N_49604);
nand UO_3897 (O_3897,N_49797,N_49829);
nand UO_3898 (O_3898,N_49870,N_49644);
nor UO_3899 (O_3899,N_49653,N_49695);
nor UO_3900 (O_3900,N_49749,N_49768);
or UO_3901 (O_3901,N_49599,N_49583);
and UO_3902 (O_3902,N_49644,N_49638);
nor UO_3903 (O_3903,N_49624,N_49675);
nand UO_3904 (O_3904,N_49587,N_49772);
and UO_3905 (O_3905,N_49767,N_49838);
xor UO_3906 (O_3906,N_49648,N_49692);
nor UO_3907 (O_3907,N_49979,N_49754);
or UO_3908 (O_3908,N_49850,N_49880);
nand UO_3909 (O_3909,N_49893,N_49568);
and UO_3910 (O_3910,N_49509,N_49967);
nand UO_3911 (O_3911,N_49998,N_49795);
xnor UO_3912 (O_3912,N_49748,N_49522);
or UO_3913 (O_3913,N_49879,N_49531);
or UO_3914 (O_3914,N_49952,N_49577);
nand UO_3915 (O_3915,N_49867,N_49575);
nor UO_3916 (O_3916,N_49603,N_49999);
nand UO_3917 (O_3917,N_49883,N_49663);
xor UO_3918 (O_3918,N_49569,N_49894);
and UO_3919 (O_3919,N_49738,N_49621);
and UO_3920 (O_3920,N_49745,N_49986);
and UO_3921 (O_3921,N_49970,N_49811);
or UO_3922 (O_3922,N_49689,N_49616);
nor UO_3923 (O_3923,N_49561,N_49664);
nor UO_3924 (O_3924,N_49569,N_49731);
xor UO_3925 (O_3925,N_49828,N_49721);
nand UO_3926 (O_3926,N_49665,N_49914);
and UO_3927 (O_3927,N_49567,N_49735);
nor UO_3928 (O_3928,N_49820,N_49663);
xnor UO_3929 (O_3929,N_49601,N_49963);
nor UO_3930 (O_3930,N_49520,N_49676);
and UO_3931 (O_3931,N_49746,N_49666);
xor UO_3932 (O_3932,N_49790,N_49647);
nor UO_3933 (O_3933,N_49582,N_49717);
and UO_3934 (O_3934,N_49869,N_49989);
and UO_3935 (O_3935,N_49800,N_49608);
nand UO_3936 (O_3936,N_49508,N_49596);
and UO_3937 (O_3937,N_49928,N_49877);
and UO_3938 (O_3938,N_49784,N_49839);
nand UO_3939 (O_3939,N_49800,N_49725);
and UO_3940 (O_3940,N_49629,N_49963);
nor UO_3941 (O_3941,N_49988,N_49907);
xnor UO_3942 (O_3942,N_49597,N_49889);
and UO_3943 (O_3943,N_49639,N_49554);
or UO_3944 (O_3944,N_49855,N_49674);
and UO_3945 (O_3945,N_49882,N_49890);
or UO_3946 (O_3946,N_49621,N_49726);
xor UO_3947 (O_3947,N_49755,N_49904);
xnor UO_3948 (O_3948,N_49601,N_49637);
or UO_3949 (O_3949,N_49551,N_49505);
nor UO_3950 (O_3950,N_49928,N_49656);
nor UO_3951 (O_3951,N_49852,N_49585);
nand UO_3952 (O_3952,N_49623,N_49664);
or UO_3953 (O_3953,N_49992,N_49546);
or UO_3954 (O_3954,N_49871,N_49988);
or UO_3955 (O_3955,N_49805,N_49593);
or UO_3956 (O_3956,N_49866,N_49958);
nand UO_3957 (O_3957,N_49783,N_49581);
nand UO_3958 (O_3958,N_49526,N_49574);
or UO_3959 (O_3959,N_49562,N_49908);
xor UO_3960 (O_3960,N_49973,N_49619);
xor UO_3961 (O_3961,N_49989,N_49903);
nand UO_3962 (O_3962,N_49931,N_49567);
nand UO_3963 (O_3963,N_49815,N_49657);
nor UO_3964 (O_3964,N_49967,N_49508);
or UO_3965 (O_3965,N_49661,N_49842);
nor UO_3966 (O_3966,N_49893,N_49840);
or UO_3967 (O_3967,N_49506,N_49515);
nand UO_3968 (O_3968,N_49682,N_49803);
nor UO_3969 (O_3969,N_49969,N_49992);
nor UO_3970 (O_3970,N_49502,N_49884);
nor UO_3971 (O_3971,N_49954,N_49755);
or UO_3972 (O_3972,N_49613,N_49842);
xnor UO_3973 (O_3973,N_49931,N_49888);
or UO_3974 (O_3974,N_49571,N_49980);
xor UO_3975 (O_3975,N_49724,N_49901);
or UO_3976 (O_3976,N_49546,N_49570);
or UO_3977 (O_3977,N_49898,N_49603);
or UO_3978 (O_3978,N_49698,N_49881);
nand UO_3979 (O_3979,N_49740,N_49799);
nand UO_3980 (O_3980,N_49650,N_49760);
xnor UO_3981 (O_3981,N_49753,N_49740);
nand UO_3982 (O_3982,N_49738,N_49787);
xnor UO_3983 (O_3983,N_49638,N_49868);
nor UO_3984 (O_3984,N_49790,N_49583);
xnor UO_3985 (O_3985,N_49778,N_49855);
and UO_3986 (O_3986,N_49925,N_49610);
nand UO_3987 (O_3987,N_49515,N_49845);
and UO_3988 (O_3988,N_49705,N_49693);
nor UO_3989 (O_3989,N_49511,N_49967);
or UO_3990 (O_3990,N_49781,N_49581);
or UO_3991 (O_3991,N_49652,N_49556);
or UO_3992 (O_3992,N_49967,N_49694);
nor UO_3993 (O_3993,N_49530,N_49610);
and UO_3994 (O_3994,N_49623,N_49729);
xnor UO_3995 (O_3995,N_49620,N_49757);
nor UO_3996 (O_3996,N_49951,N_49806);
nand UO_3997 (O_3997,N_49676,N_49639);
and UO_3998 (O_3998,N_49844,N_49705);
or UO_3999 (O_3999,N_49871,N_49842);
or UO_4000 (O_4000,N_49747,N_49846);
xnor UO_4001 (O_4001,N_49911,N_49993);
xnor UO_4002 (O_4002,N_49536,N_49619);
nand UO_4003 (O_4003,N_49942,N_49615);
and UO_4004 (O_4004,N_49701,N_49639);
and UO_4005 (O_4005,N_49833,N_49654);
or UO_4006 (O_4006,N_49721,N_49993);
nor UO_4007 (O_4007,N_49859,N_49604);
xnor UO_4008 (O_4008,N_49607,N_49521);
and UO_4009 (O_4009,N_49919,N_49751);
and UO_4010 (O_4010,N_49582,N_49633);
nor UO_4011 (O_4011,N_49602,N_49637);
xor UO_4012 (O_4012,N_49633,N_49742);
or UO_4013 (O_4013,N_49588,N_49632);
nand UO_4014 (O_4014,N_49565,N_49543);
and UO_4015 (O_4015,N_49779,N_49873);
xor UO_4016 (O_4016,N_49521,N_49657);
and UO_4017 (O_4017,N_49708,N_49686);
nand UO_4018 (O_4018,N_49658,N_49629);
or UO_4019 (O_4019,N_49516,N_49975);
or UO_4020 (O_4020,N_49606,N_49900);
and UO_4021 (O_4021,N_49888,N_49644);
and UO_4022 (O_4022,N_49581,N_49663);
xor UO_4023 (O_4023,N_49935,N_49722);
nand UO_4024 (O_4024,N_49759,N_49776);
and UO_4025 (O_4025,N_49723,N_49769);
nor UO_4026 (O_4026,N_49765,N_49650);
and UO_4027 (O_4027,N_49651,N_49967);
or UO_4028 (O_4028,N_49582,N_49902);
nand UO_4029 (O_4029,N_49743,N_49965);
nand UO_4030 (O_4030,N_49913,N_49765);
nor UO_4031 (O_4031,N_49941,N_49905);
and UO_4032 (O_4032,N_49702,N_49946);
xnor UO_4033 (O_4033,N_49642,N_49627);
or UO_4034 (O_4034,N_49805,N_49886);
and UO_4035 (O_4035,N_49895,N_49604);
xnor UO_4036 (O_4036,N_49561,N_49931);
nand UO_4037 (O_4037,N_49994,N_49899);
nor UO_4038 (O_4038,N_49934,N_49637);
or UO_4039 (O_4039,N_49539,N_49514);
and UO_4040 (O_4040,N_49819,N_49899);
xnor UO_4041 (O_4041,N_49526,N_49502);
nand UO_4042 (O_4042,N_49774,N_49524);
nand UO_4043 (O_4043,N_49507,N_49794);
and UO_4044 (O_4044,N_49782,N_49811);
xor UO_4045 (O_4045,N_49956,N_49859);
nand UO_4046 (O_4046,N_49557,N_49526);
and UO_4047 (O_4047,N_49951,N_49728);
xnor UO_4048 (O_4048,N_49522,N_49994);
xor UO_4049 (O_4049,N_49633,N_49704);
nor UO_4050 (O_4050,N_49993,N_49530);
xor UO_4051 (O_4051,N_49881,N_49568);
or UO_4052 (O_4052,N_49531,N_49578);
or UO_4053 (O_4053,N_49666,N_49538);
xor UO_4054 (O_4054,N_49665,N_49730);
nand UO_4055 (O_4055,N_49505,N_49737);
and UO_4056 (O_4056,N_49661,N_49613);
or UO_4057 (O_4057,N_49547,N_49862);
nand UO_4058 (O_4058,N_49945,N_49629);
nor UO_4059 (O_4059,N_49856,N_49813);
nand UO_4060 (O_4060,N_49663,N_49747);
nand UO_4061 (O_4061,N_49532,N_49538);
or UO_4062 (O_4062,N_49648,N_49688);
nor UO_4063 (O_4063,N_49902,N_49564);
nor UO_4064 (O_4064,N_49618,N_49798);
xnor UO_4065 (O_4065,N_49879,N_49684);
nand UO_4066 (O_4066,N_49956,N_49921);
nor UO_4067 (O_4067,N_49568,N_49650);
xnor UO_4068 (O_4068,N_49566,N_49919);
nand UO_4069 (O_4069,N_49623,N_49695);
nor UO_4070 (O_4070,N_49944,N_49882);
nor UO_4071 (O_4071,N_49592,N_49779);
nor UO_4072 (O_4072,N_49797,N_49745);
xnor UO_4073 (O_4073,N_49523,N_49534);
or UO_4074 (O_4074,N_49696,N_49766);
and UO_4075 (O_4075,N_49911,N_49658);
xor UO_4076 (O_4076,N_49502,N_49947);
xnor UO_4077 (O_4077,N_49625,N_49754);
and UO_4078 (O_4078,N_49830,N_49799);
or UO_4079 (O_4079,N_49887,N_49922);
nor UO_4080 (O_4080,N_49584,N_49978);
and UO_4081 (O_4081,N_49577,N_49797);
and UO_4082 (O_4082,N_49749,N_49843);
nand UO_4083 (O_4083,N_49569,N_49754);
nor UO_4084 (O_4084,N_49913,N_49610);
xnor UO_4085 (O_4085,N_49957,N_49561);
xor UO_4086 (O_4086,N_49775,N_49823);
nand UO_4087 (O_4087,N_49945,N_49843);
and UO_4088 (O_4088,N_49998,N_49705);
xnor UO_4089 (O_4089,N_49944,N_49519);
nor UO_4090 (O_4090,N_49972,N_49594);
or UO_4091 (O_4091,N_49654,N_49598);
xnor UO_4092 (O_4092,N_49718,N_49922);
and UO_4093 (O_4093,N_49614,N_49786);
nor UO_4094 (O_4094,N_49750,N_49734);
or UO_4095 (O_4095,N_49660,N_49522);
xor UO_4096 (O_4096,N_49899,N_49798);
xor UO_4097 (O_4097,N_49692,N_49594);
or UO_4098 (O_4098,N_49960,N_49504);
xnor UO_4099 (O_4099,N_49535,N_49602);
or UO_4100 (O_4100,N_49549,N_49536);
and UO_4101 (O_4101,N_49705,N_49647);
or UO_4102 (O_4102,N_49520,N_49652);
nor UO_4103 (O_4103,N_49539,N_49809);
nand UO_4104 (O_4104,N_49585,N_49569);
or UO_4105 (O_4105,N_49802,N_49791);
nor UO_4106 (O_4106,N_49550,N_49718);
nor UO_4107 (O_4107,N_49710,N_49655);
or UO_4108 (O_4108,N_49656,N_49580);
and UO_4109 (O_4109,N_49528,N_49642);
nor UO_4110 (O_4110,N_49518,N_49636);
nand UO_4111 (O_4111,N_49552,N_49731);
or UO_4112 (O_4112,N_49580,N_49739);
nor UO_4113 (O_4113,N_49582,N_49511);
xor UO_4114 (O_4114,N_49939,N_49769);
nand UO_4115 (O_4115,N_49856,N_49579);
nand UO_4116 (O_4116,N_49588,N_49596);
nor UO_4117 (O_4117,N_49645,N_49838);
or UO_4118 (O_4118,N_49875,N_49678);
xnor UO_4119 (O_4119,N_49764,N_49903);
or UO_4120 (O_4120,N_49938,N_49942);
xor UO_4121 (O_4121,N_49565,N_49793);
and UO_4122 (O_4122,N_49673,N_49801);
nor UO_4123 (O_4123,N_49755,N_49516);
or UO_4124 (O_4124,N_49941,N_49839);
nand UO_4125 (O_4125,N_49787,N_49679);
xnor UO_4126 (O_4126,N_49528,N_49538);
or UO_4127 (O_4127,N_49790,N_49710);
xor UO_4128 (O_4128,N_49788,N_49618);
xor UO_4129 (O_4129,N_49627,N_49848);
nand UO_4130 (O_4130,N_49686,N_49893);
and UO_4131 (O_4131,N_49967,N_49736);
nor UO_4132 (O_4132,N_49822,N_49538);
or UO_4133 (O_4133,N_49514,N_49966);
nand UO_4134 (O_4134,N_49565,N_49579);
or UO_4135 (O_4135,N_49783,N_49893);
xnor UO_4136 (O_4136,N_49824,N_49763);
nor UO_4137 (O_4137,N_49969,N_49675);
nor UO_4138 (O_4138,N_49798,N_49797);
or UO_4139 (O_4139,N_49727,N_49933);
and UO_4140 (O_4140,N_49993,N_49695);
nor UO_4141 (O_4141,N_49535,N_49842);
or UO_4142 (O_4142,N_49507,N_49589);
xnor UO_4143 (O_4143,N_49881,N_49655);
xor UO_4144 (O_4144,N_49572,N_49787);
and UO_4145 (O_4145,N_49561,N_49515);
or UO_4146 (O_4146,N_49709,N_49670);
nor UO_4147 (O_4147,N_49810,N_49684);
or UO_4148 (O_4148,N_49722,N_49698);
nand UO_4149 (O_4149,N_49840,N_49515);
nand UO_4150 (O_4150,N_49935,N_49500);
nor UO_4151 (O_4151,N_49519,N_49550);
or UO_4152 (O_4152,N_49721,N_49849);
and UO_4153 (O_4153,N_49939,N_49927);
nand UO_4154 (O_4154,N_49982,N_49662);
and UO_4155 (O_4155,N_49791,N_49708);
nor UO_4156 (O_4156,N_49944,N_49781);
nor UO_4157 (O_4157,N_49900,N_49724);
or UO_4158 (O_4158,N_49717,N_49914);
nand UO_4159 (O_4159,N_49831,N_49598);
xnor UO_4160 (O_4160,N_49558,N_49547);
xnor UO_4161 (O_4161,N_49543,N_49778);
xor UO_4162 (O_4162,N_49881,N_49993);
nand UO_4163 (O_4163,N_49538,N_49753);
and UO_4164 (O_4164,N_49660,N_49644);
and UO_4165 (O_4165,N_49759,N_49628);
and UO_4166 (O_4166,N_49878,N_49527);
and UO_4167 (O_4167,N_49711,N_49785);
xor UO_4168 (O_4168,N_49571,N_49731);
xnor UO_4169 (O_4169,N_49617,N_49673);
nor UO_4170 (O_4170,N_49538,N_49819);
and UO_4171 (O_4171,N_49984,N_49891);
and UO_4172 (O_4172,N_49733,N_49602);
or UO_4173 (O_4173,N_49784,N_49947);
nor UO_4174 (O_4174,N_49553,N_49856);
and UO_4175 (O_4175,N_49820,N_49959);
xnor UO_4176 (O_4176,N_49814,N_49848);
and UO_4177 (O_4177,N_49659,N_49628);
nor UO_4178 (O_4178,N_49551,N_49686);
xnor UO_4179 (O_4179,N_49827,N_49572);
and UO_4180 (O_4180,N_49558,N_49533);
and UO_4181 (O_4181,N_49544,N_49522);
nand UO_4182 (O_4182,N_49885,N_49537);
nor UO_4183 (O_4183,N_49594,N_49621);
and UO_4184 (O_4184,N_49685,N_49799);
nor UO_4185 (O_4185,N_49858,N_49836);
xnor UO_4186 (O_4186,N_49909,N_49837);
or UO_4187 (O_4187,N_49575,N_49630);
xnor UO_4188 (O_4188,N_49891,N_49857);
xnor UO_4189 (O_4189,N_49672,N_49710);
or UO_4190 (O_4190,N_49506,N_49921);
nor UO_4191 (O_4191,N_49522,N_49686);
nand UO_4192 (O_4192,N_49961,N_49891);
or UO_4193 (O_4193,N_49811,N_49625);
and UO_4194 (O_4194,N_49881,N_49823);
nor UO_4195 (O_4195,N_49819,N_49523);
nand UO_4196 (O_4196,N_49546,N_49879);
nand UO_4197 (O_4197,N_49621,N_49617);
and UO_4198 (O_4198,N_49812,N_49989);
or UO_4199 (O_4199,N_49575,N_49625);
and UO_4200 (O_4200,N_49675,N_49958);
xnor UO_4201 (O_4201,N_49912,N_49670);
nor UO_4202 (O_4202,N_49890,N_49824);
xor UO_4203 (O_4203,N_49963,N_49532);
nor UO_4204 (O_4204,N_49895,N_49864);
and UO_4205 (O_4205,N_49890,N_49853);
nor UO_4206 (O_4206,N_49882,N_49967);
and UO_4207 (O_4207,N_49930,N_49855);
nor UO_4208 (O_4208,N_49890,N_49787);
nor UO_4209 (O_4209,N_49670,N_49961);
nand UO_4210 (O_4210,N_49959,N_49536);
and UO_4211 (O_4211,N_49592,N_49763);
xnor UO_4212 (O_4212,N_49614,N_49629);
and UO_4213 (O_4213,N_49503,N_49756);
and UO_4214 (O_4214,N_49652,N_49680);
nor UO_4215 (O_4215,N_49930,N_49689);
or UO_4216 (O_4216,N_49769,N_49952);
nor UO_4217 (O_4217,N_49702,N_49966);
or UO_4218 (O_4218,N_49843,N_49685);
xor UO_4219 (O_4219,N_49854,N_49720);
or UO_4220 (O_4220,N_49767,N_49847);
and UO_4221 (O_4221,N_49972,N_49567);
xor UO_4222 (O_4222,N_49617,N_49567);
nand UO_4223 (O_4223,N_49988,N_49986);
nor UO_4224 (O_4224,N_49859,N_49936);
nor UO_4225 (O_4225,N_49747,N_49830);
and UO_4226 (O_4226,N_49873,N_49920);
nor UO_4227 (O_4227,N_49537,N_49900);
xnor UO_4228 (O_4228,N_49782,N_49656);
or UO_4229 (O_4229,N_49947,N_49500);
nor UO_4230 (O_4230,N_49728,N_49779);
and UO_4231 (O_4231,N_49533,N_49745);
or UO_4232 (O_4232,N_49744,N_49943);
and UO_4233 (O_4233,N_49831,N_49799);
and UO_4234 (O_4234,N_49577,N_49770);
nand UO_4235 (O_4235,N_49576,N_49650);
nor UO_4236 (O_4236,N_49795,N_49593);
nand UO_4237 (O_4237,N_49933,N_49532);
nor UO_4238 (O_4238,N_49920,N_49901);
nor UO_4239 (O_4239,N_49920,N_49666);
xnor UO_4240 (O_4240,N_49824,N_49978);
nand UO_4241 (O_4241,N_49776,N_49930);
nor UO_4242 (O_4242,N_49521,N_49629);
nand UO_4243 (O_4243,N_49685,N_49701);
nor UO_4244 (O_4244,N_49839,N_49662);
and UO_4245 (O_4245,N_49653,N_49503);
or UO_4246 (O_4246,N_49754,N_49994);
xnor UO_4247 (O_4247,N_49582,N_49537);
xor UO_4248 (O_4248,N_49866,N_49682);
nand UO_4249 (O_4249,N_49759,N_49650);
nor UO_4250 (O_4250,N_49594,N_49786);
or UO_4251 (O_4251,N_49977,N_49929);
or UO_4252 (O_4252,N_49844,N_49909);
nand UO_4253 (O_4253,N_49557,N_49618);
nor UO_4254 (O_4254,N_49845,N_49526);
nand UO_4255 (O_4255,N_49776,N_49657);
and UO_4256 (O_4256,N_49739,N_49808);
nand UO_4257 (O_4257,N_49931,N_49700);
nand UO_4258 (O_4258,N_49708,N_49700);
and UO_4259 (O_4259,N_49516,N_49798);
and UO_4260 (O_4260,N_49517,N_49611);
xnor UO_4261 (O_4261,N_49822,N_49927);
xor UO_4262 (O_4262,N_49557,N_49568);
xor UO_4263 (O_4263,N_49945,N_49753);
nor UO_4264 (O_4264,N_49571,N_49778);
and UO_4265 (O_4265,N_49812,N_49694);
xnor UO_4266 (O_4266,N_49905,N_49649);
or UO_4267 (O_4267,N_49859,N_49916);
nor UO_4268 (O_4268,N_49821,N_49690);
and UO_4269 (O_4269,N_49740,N_49818);
nand UO_4270 (O_4270,N_49831,N_49528);
or UO_4271 (O_4271,N_49656,N_49722);
nand UO_4272 (O_4272,N_49516,N_49897);
xnor UO_4273 (O_4273,N_49779,N_49969);
and UO_4274 (O_4274,N_49949,N_49508);
xor UO_4275 (O_4275,N_49670,N_49848);
nor UO_4276 (O_4276,N_49962,N_49517);
nor UO_4277 (O_4277,N_49946,N_49732);
nor UO_4278 (O_4278,N_49925,N_49830);
and UO_4279 (O_4279,N_49869,N_49619);
xor UO_4280 (O_4280,N_49849,N_49690);
and UO_4281 (O_4281,N_49721,N_49908);
and UO_4282 (O_4282,N_49615,N_49690);
nand UO_4283 (O_4283,N_49652,N_49538);
xor UO_4284 (O_4284,N_49610,N_49763);
and UO_4285 (O_4285,N_49869,N_49747);
nand UO_4286 (O_4286,N_49506,N_49962);
nand UO_4287 (O_4287,N_49924,N_49976);
xor UO_4288 (O_4288,N_49850,N_49576);
nand UO_4289 (O_4289,N_49802,N_49511);
xnor UO_4290 (O_4290,N_49647,N_49602);
xor UO_4291 (O_4291,N_49675,N_49984);
or UO_4292 (O_4292,N_49682,N_49882);
xor UO_4293 (O_4293,N_49568,N_49991);
and UO_4294 (O_4294,N_49942,N_49934);
or UO_4295 (O_4295,N_49911,N_49522);
nor UO_4296 (O_4296,N_49541,N_49513);
and UO_4297 (O_4297,N_49979,N_49601);
nor UO_4298 (O_4298,N_49759,N_49583);
nand UO_4299 (O_4299,N_49801,N_49877);
nor UO_4300 (O_4300,N_49596,N_49871);
nand UO_4301 (O_4301,N_49636,N_49791);
xnor UO_4302 (O_4302,N_49556,N_49935);
or UO_4303 (O_4303,N_49861,N_49522);
nor UO_4304 (O_4304,N_49702,N_49579);
xnor UO_4305 (O_4305,N_49850,N_49864);
nand UO_4306 (O_4306,N_49821,N_49758);
nor UO_4307 (O_4307,N_49883,N_49787);
and UO_4308 (O_4308,N_49714,N_49868);
or UO_4309 (O_4309,N_49973,N_49875);
xor UO_4310 (O_4310,N_49686,N_49665);
xor UO_4311 (O_4311,N_49585,N_49910);
nand UO_4312 (O_4312,N_49717,N_49562);
or UO_4313 (O_4313,N_49926,N_49652);
nand UO_4314 (O_4314,N_49506,N_49578);
and UO_4315 (O_4315,N_49552,N_49532);
nor UO_4316 (O_4316,N_49635,N_49920);
nor UO_4317 (O_4317,N_49877,N_49818);
nor UO_4318 (O_4318,N_49712,N_49515);
nor UO_4319 (O_4319,N_49818,N_49794);
nor UO_4320 (O_4320,N_49615,N_49936);
nand UO_4321 (O_4321,N_49683,N_49850);
and UO_4322 (O_4322,N_49786,N_49928);
xnor UO_4323 (O_4323,N_49849,N_49916);
xnor UO_4324 (O_4324,N_49600,N_49678);
nand UO_4325 (O_4325,N_49591,N_49652);
or UO_4326 (O_4326,N_49781,N_49813);
xnor UO_4327 (O_4327,N_49667,N_49868);
or UO_4328 (O_4328,N_49883,N_49757);
and UO_4329 (O_4329,N_49892,N_49602);
nand UO_4330 (O_4330,N_49757,N_49826);
xnor UO_4331 (O_4331,N_49927,N_49554);
nor UO_4332 (O_4332,N_49668,N_49845);
or UO_4333 (O_4333,N_49586,N_49888);
or UO_4334 (O_4334,N_49795,N_49892);
nor UO_4335 (O_4335,N_49513,N_49830);
xor UO_4336 (O_4336,N_49753,N_49800);
and UO_4337 (O_4337,N_49879,N_49636);
nor UO_4338 (O_4338,N_49662,N_49631);
nand UO_4339 (O_4339,N_49661,N_49831);
or UO_4340 (O_4340,N_49875,N_49822);
or UO_4341 (O_4341,N_49971,N_49580);
nand UO_4342 (O_4342,N_49717,N_49899);
xnor UO_4343 (O_4343,N_49732,N_49996);
or UO_4344 (O_4344,N_49931,N_49919);
or UO_4345 (O_4345,N_49609,N_49970);
or UO_4346 (O_4346,N_49545,N_49539);
or UO_4347 (O_4347,N_49788,N_49760);
and UO_4348 (O_4348,N_49871,N_49700);
or UO_4349 (O_4349,N_49511,N_49705);
and UO_4350 (O_4350,N_49775,N_49740);
xor UO_4351 (O_4351,N_49934,N_49702);
nand UO_4352 (O_4352,N_49525,N_49617);
nor UO_4353 (O_4353,N_49925,N_49656);
or UO_4354 (O_4354,N_49558,N_49571);
and UO_4355 (O_4355,N_49802,N_49974);
or UO_4356 (O_4356,N_49651,N_49540);
nand UO_4357 (O_4357,N_49859,N_49732);
nor UO_4358 (O_4358,N_49528,N_49998);
or UO_4359 (O_4359,N_49572,N_49527);
or UO_4360 (O_4360,N_49773,N_49815);
xnor UO_4361 (O_4361,N_49630,N_49714);
nor UO_4362 (O_4362,N_49699,N_49641);
nand UO_4363 (O_4363,N_49889,N_49750);
and UO_4364 (O_4364,N_49961,N_49895);
nor UO_4365 (O_4365,N_49897,N_49858);
or UO_4366 (O_4366,N_49629,N_49817);
or UO_4367 (O_4367,N_49781,N_49582);
and UO_4368 (O_4368,N_49940,N_49992);
nand UO_4369 (O_4369,N_49925,N_49542);
nand UO_4370 (O_4370,N_49708,N_49837);
nand UO_4371 (O_4371,N_49603,N_49846);
nand UO_4372 (O_4372,N_49600,N_49941);
xnor UO_4373 (O_4373,N_49640,N_49758);
xnor UO_4374 (O_4374,N_49987,N_49806);
xor UO_4375 (O_4375,N_49745,N_49861);
or UO_4376 (O_4376,N_49698,N_49845);
and UO_4377 (O_4377,N_49800,N_49628);
nor UO_4378 (O_4378,N_49869,N_49836);
nor UO_4379 (O_4379,N_49768,N_49881);
nor UO_4380 (O_4380,N_49834,N_49722);
xnor UO_4381 (O_4381,N_49638,N_49695);
nor UO_4382 (O_4382,N_49687,N_49745);
nand UO_4383 (O_4383,N_49925,N_49771);
nand UO_4384 (O_4384,N_49541,N_49956);
nor UO_4385 (O_4385,N_49656,N_49914);
xor UO_4386 (O_4386,N_49796,N_49789);
nand UO_4387 (O_4387,N_49850,N_49828);
or UO_4388 (O_4388,N_49972,N_49635);
or UO_4389 (O_4389,N_49999,N_49678);
xor UO_4390 (O_4390,N_49588,N_49859);
nand UO_4391 (O_4391,N_49558,N_49907);
and UO_4392 (O_4392,N_49707,N_49758);
nand UO_4393 (O_4393,N_49731,N_49867);
and UO_4394 (O_4394,N_49909,N_49945);
and UO_4395 (O_4395,N_49873,N_49680);
nand UO_4396 (O_4396,N_49819,N_49584);
nand UO_4397 (O_4397,N_49627,N_49746);
or UO_4398 (O_4398,N_49876,N_49838);
nand UO_4399 (O_4399,N_49975,N_49831);
nand UO_4400 (O_4400,N_49588,N_49556);
nor UO_4401 (O_4401,N_49869,N_49523);
xor UO_4402 (O_4402,N_49819,N_49571);
nor UO_4403 (O_4403,N_49684,N_49884);
nor UO_4404 (O_4404,N_49897,N_49633);
nand UO_4405 (O_4405,N_49924,N_49733);
nand UO_4406 (O_4406,N_49992,N_49601);
xnor UO_4407 (O_4407,N_49511,N_49831);
xnor UO_4408 (O_4408,N_49792,N_49838);
nand UO_4409 (O_4409,N_49702,N_49641);
and UO_4410 (O_4410,N_49862,N_49966);
xnor UO_4411 (O_4411,N_49500,N_49843);
nand UO_4412 (O_4412,N_49700,N_49948);
xor UO_4413 (O_4413,N_49617,N_49583);
and UO_4414 (O_4414,N_49628,N_49994);
nand UO_4415 (O_4415,N_49988,N_49775);
nor UO_4416 (O_4416,N_49947,N_49515);
nand UO_4417 (O_4417,N_49687,N_49612);
xor UO_4418 (O_4418,N_49696,N_49980);
or UO_4419 (O_4419,N_49500,N_49958);
nor UO_4420 (O_4420,N_49815,N_49902);
and UO_4421 (O_4421,N_49817,N_49912);
xor UO_4422 (O_4422,N_49538,N_49877);
or UO_4423 (O_4423,N_49621,N_49935);
or UO_4424 (O_4424,N_49762,N_49968);
nand UO_4425 (O_4425,N_49816,N_49543);
nand UO_4426 (O_4426,N_49934,N_49815);
nor UO_4427 (O_4427,N_49520,N_49588);
or UO_4428 (O_4428,N_49762,N_49682);
and UO_4429 (O_4429,N_49916,N_49598);
xnor UO_4430 (O_4430,N_49749,N_49615);
nor UO_4431 (O_4431,N_49904,N_49594);
and UO_4432 (O_4432,N_49501,N_49881);
or UO_4433 (O_4433,N_49576,N_49935);
nor UO_4434 (O_4434,N_49506,N_49852);
nand UO_4435 (O_4435,N_49773,N_49678);
xor UO_4436 (O_4436,N_49870,N_49864);
and UO_4437 (O_4437,N_49827,N_49613);
nor UO_4438 (O_4438,N_49745,N_49939);
nand UO_4439 (O_4439,N_49559,N_49923);
or UO_4440 (O_4440,N_49857,N_49753);
nand UO_4441 (O_4441,N_49790,N_49605);
xor UO_4442 (O_4442,N_49670,N_49794);
xor UO_4443 (O_4443,N_49586,N_49764);
or UO_4444 (O_4444,N_49739,N_49833);
and UO_4445 (O_4445,N_49718,N_49968);
nand UO_4446 (O_4446,N_49512,N_49584);
nand UO_4447 (O_4447,N_49827,N_49769);
and UO_4448 (O_4448,N_49576,N_49537);
nand UO_4449 (O_4449,N_49953,N_49944);
xnor UO_4450 (O_4450,N_49825,N_49972);
nor UO_4451 (O_4451,N_49708,N_49852);
and UO_4452 (O_4452,N_49796,N_49643);
and UO_4453 (O_4453,N_49777,N_49816);
xnor UO_4454 (O_4454,N_49861,N_49873);
xnor UO_4455 (O_4455,N_49643,N_49564);
or UO_4456 (O_4456,N_49894,N_49854);
nand UO_4457 (O_4457,N_49979,N_49828);
or UO_4458 (O_4458,N_49778,N_49926);
or UO_4459 (O_4459,N_49503,N_49768);
nand UO_4460 (O_4460,N_49740,N_49583);
and UO_4461 (O_4461,N_49804,N_49722);
or UO_4462 (O_4462,N_49941,N_49873);
or UO_4463 (O_4463,N_49851,N_49788);
nor UO_4464 (O_4464,N_49617,N_49871);
or UO_4465 (O_4465,N_49590,N_49966);
nor UO_4466 (O_4466,N_49670,N_49544);
or UO_4467 (O_4467,N_49525,N_49701);
or UO_4468 (O_4468,N_49555,N_49695);
or UO_4469 (O_4469,N_49637,N_49767);
and UO_4470 (O_4470,N_49633,N_49854);
and UO_4471 (O_4471,N_49651,N_49547);
or UO_4472 (O_4472,N_49761,N_49665);
nand UO_4473 (O_4473,N_49817,N_49664);
or UO_4474 (O_4474,N_49650,N_49501);
nor UO_4475 (O_4475,N_49997,N_49979);
nand UO_4476 (O_4476,N_49958,N_49913);
nand UO_4477 (O_4477,N_49658,N_49547);
and UO_4478 (O_4478,N_49596,N_49690);
nand UO_4479 (O_4479,N_49692,N_49725);
or UO_4480 (O_4480,N_49635,N_49960);
xor UO_4481 (O_4481,N_49936,N_49854);
nand UO_4482 (O_4482,N_49923,N_49736);
or UO_4483 (O_4483,N_49854,N_49604);
or UO_4484 (O_4484,N_49747,N_49678);
xor UO_4485 (O_4485,N_49849,N_49711);
and UO_4486 (O_4486,N_49865,N_49900);
xnor UO_4487 (O_4487,N_49536,N_49558);
nand UO_4488 (O_4488,N_49859,N_49797);
nand UO_4489 (O_4489,N_49882,N_49864);
nand UO_4490 (O_4490,N_49960,N_49932);
and UO_4491 (O_4491,N_49643,N_49588);
nor UO_4492 (O_4492,N_49825,N_49684);
nor UO_4493 (O_4493,N_49983,N_49971);
and UO_4494 (O_4494,N_49549,N_49889);
nor UO_4495 (O_4495,N_49899,N_49543);
nor UO_4496 (O_4496,N_49807,N_49968);
nor UO_4497 (O_4497,N_49941,N_49979);
nor UO_4498 (O_4498,N_49549,N_49644);
or UO_4499 (O_4499,N_49662,N_49951);
nand UO_4500 (O_4500,N_49958,N_49809);
xnor UO_4501 (O_4501,N_49666,N_49862);
or UO_4502 (O_4502,N_49938,N_49726);
nor UO_4503 (O_4503,N_49760,N_49841);
nor UO_4504 (O_4504,N_49766,N_49532);
xor UO_4505 (O_4505,N_49666,N_49868);
nor UO_4506 (O_4506,N_49769,N_49786);
nand UO_4507 (O_4507,N_49750,N_49554);
and UO_4508 (O_4508,N_49986,N_49834);
and UO_4509 (O_4509,N_49832,N_49610);
and UO_4510 (O_4510,N_49555,N_49505);
or UO_4511 (O_4511,N_49639,N_49580);
nor UO_4512 (O_4512,N_49591,N_49825);
or UO_4513 (O_4513,N_49754,N_49619);
and UO_4514 (O_4514,N_49663,N_49885);
and UO_4515 (O_4515,N_49779,N_49524);
nor UO_4516 (O_4516,N_49930,N_49639);
or UO_4517 (O_4517,N_49928,N_49540);
and UO_4518 (O_4518,N_49954,N_49691);
or UO_4519 (O_4519,N_49844,N_49609);
nand UO_4520 (O_4520,N_49760,N_49919);
nand UO_4521 (O_4521,N_49573,N_49978);
xnor UO_4522 (O_4522,N_49594,N_49825);
or UO_4523 (O_4523,N_49884,N_49686);
xnor UO_4524 (O_4524,N_49892,N_49575);
nor UO_4525 (O_4525,N_49935,N_49900);
nor UO_4526 (O_4526,N_49932,N_49614);
nor UO_4527 (O_4527,N_49617,N_49965);
xor UO_4528 (O_4528,N_49766,N_49871);
and UO_4529 (O_4529,N_49587,N_49677);
nor UO_4530 (O_4530,N_49947,N_49755);
nor UO_4531 (O_4531,N_49851,N_49918);
xor UO_4532 (O_4532,N_49911,N_49887);
xor UO_4533 (O_4533,N_49838,N_49564);
nand UO_4534 (O_4534,N_49634,N_49547);
xnor UO_4535 (O_4535,N_49608,N_49941);
xnor UO_4536 (O_4536,N_49539,N_49962);
nand UO_4537 (O_4537,N_49573,N_49738);
nand UO_4538 (O_4538,N_49748,N_49727);
xnor UO_4539 (O_4539,N_49962,N_49958);
and UO_4540 (O_4540,N_49723,N_49807);
nor UO_4541 (O_4541,N_49739,N_49690);
or UO_4542 (O_4542,N_49518,N_49990);
nand UO_4543 (O_4543,N_49627,N_49717);
xor UO_4544 (O_4544,N_49661,N_49517);
or UO_4545 (O_4545,N_49874,N_49699);
xnor UO_4546 (O_4546,N_49901,N_49520);
or UO_4547 (O_4547,N_49632,N_49785);
or UO_4548 (O_4548,N_49530,N_49978);
and UO_4549 (O_4549,N_49534,N_49689);
or UO_4550 (O_4550,N_49560,N_49842);
and UO_4551 (O_4551,N_49805,N_49906);
nor UO_4552 (O_4552,N_49548,N_49995);
xor UO_4553 (O_4553,N_49941,N_49659);
nor UO_4554 (O_4554,N_49897,N_49510);
xor UO_4555 (O_4555,N_49887,N_49678);
nand UO_4556 (O_4556,N_49544,N_49803);
xnor UO_4557 (O_4557,N_49516,N_49985);
xnor UO_4558 (O_4558,N_49739,N_49680);
and UO_4559 (O_4559,N_49922,N_49552);
nor UO_4560 (O_4560,N_49893,N_49760);
nor UO_4561 (O_4561,N_49972,N_49669);
and UO_4562 (O_4562,N_49510,N_49599);
and UO_4563 (O_4563,N_49945,N_49544);
or UO_4564 (O_4564,N_49683,N_49669);
nor UO_4565 (O_4565,N_49713,N_49877);
nand UO_4566 (O_4566,N_49741,N_49771);
and UO_4567 (O_4567,N_49792,N_49502);
xor UO_4568 (O_4568,N_49737,N_49613);
and UO_4569 (O_4569,N_49657,N_49849);
and UO_4570 (O_4570,N_49596,N_49565);
nor UO_4571 (O_4571,N_49888,N_49688);
or UO_4572 (O_4572,N_49716,N_49979);
xor UO_4573 (O_4573,N_49693,N_49794);
nor UO_4574 (O_4574,N_49842,N_49538);
and UO_4575 (O_4575,N_49528,N_49991);
nor UO_4576 (O_4576,N_49729,N_49975);
nor UO_4577 (O_4577,N_49891,N_49505);
xnor UO_4578 (O_4578,N_49511,N_49850);
nand UO_4579 (O_4579,N_49600,N_49728);
xor UO_4580 (O_4580,N_49638,N_49915);
xor UO_4581 (O_4581,N_49729,N_49793);
nand UO_4582 (O_4582,N_49603,N_49600);
and UO_4583 (O_4583,N_49562,N_49913);
nand UO_4584 (O_4584,N_49510,N_49606);
xor UO_4585 (O_4585,N_49918,N_49605);
nand UO_4586 (O_4586,N_49573,N_49614);
and UO_4587 (O_4587,N_49857,N_49521);
and UO_4588 (O_4588,N_49929,N_49615);
nor UO_4589 (O_4589,N_49626,N_49794);
nand UO_4590 (O_4590,N_49905,N_49823);
xnor UO_4591 (O_4591,N_49740,N_49955);
and UO_4592 (O_4592,N_49511,N_49693);
xnor UO_4593 (O_4593,N_49810,N_49796);
nor UO_4594 (O_4594,N_49637,N_49802);
and UO_4595 (O_4595,N_49754,N_49504);
nor UO_4596 (O_4596,N_49892,N_49712);
nand UO_4597 (O_4597,N_49894,N_49918);
or UO_4598 (O_4598,N_49909,N_49959);
nor UO_4599 (O_4599,N_49987,N_49869);
nand UO_4600 (O_4600,N_49692,N_49792);
and UO_4601 (O_4601,N_49569,N_49660);
nor UO_4602 (O_4602,N_49655,N_49752);
nand UO_4603 (O_4603,N_49518,N_49716);
nor UO_4604 (O_4604,N_49597,N_49704);
or UO_4605 (O_4605,N_49693,N_49746);
nor UO_4606 (O_4606,N_49512,N_49569);
and UO_4607 (O_4607,N_49506,N_49790);
nor UO_4608 (O_4608,N_49505,N_49990);
nand UO_4609 (O_4609,N_49892,N_49878);
and UO_4610 (O_4610,N_49700,N_49610);
and UO_4611 (O_4611,N_49819,N_49907);
xor UO_4612 (O_4612,N_49694,N_49549);
or UO_4613 (O_4613,N_49711,N_49943);
or UO_4614 (O_4614,N_49513,N_49901);
nand UO_4615 (O_4615,N_49615,N_49736);
xor UO_4616 (O_4616,N_49922,N_49649);
nand UO_4617 (O_4617,N_49931,N_49739);
nand UO_4618 (O_4618,N_49547,N_49602);
nor UO_4619 (O_4619,N_49762,N_49596);
xnor UO_4620 (O_4620,N_49912,N_49601);
or UO_4621 (O_4621,N_49500,N_49578);
nand UO_4622 (O_4622,N_49917,N_49887);
nand UO_4623 (O_4623,N_49687,N_49892);
or UO_4624 (O_4624,N_49789,N_49751);
nand UO_4625 (O_4625,N_49555,N_49545);
nand UO_4626 (O_4626,N_49760,N_49590);
or UO_4627 (O_4627,N_49628,N_49605);
or UO_4628 (O_4628,N_49513,N_49897);
or UO_4629 (O_4629,N_49636,N_49841);
and UO_4630 (O_4630,N_49986,N_49847);
nor UO_4631 (O_4631,N_49573,N_49903);
nand UO_4632 (O_4632,N_49519,N_49653);
nand UO_4633 (O_4633,N_49645,N_49580);
or UO_4634 (O_4634,N_49569,N_49704);
and UO_4635 (O_4635,N_49968,N_49676);
and UO_4636 (O_4636,N_49818,N_49948);
xor UO_4637 (O_4637,N_49568,N_49634);
and UO_4638 (O_4638,N_49920,N_49685);
and UO_4639 (O_4639,N_49865,N_49662);
and UO_4640 (O_4640,N_49947,N_49896);
or UO_4641 (O_4641,N_49576,N_49833);
nand UO_4642 (O_4642,N_49637,N_49548);
and UO_4643 (O_4643,N_49728,N_49550);
and UO_4644 (O_4644,N_49678,N_49950);
or UO_4645 (O_4645,N_49969,N_49788);
nor UO_4646 (O_4646,N_49824,N_49555);
xnor UO_4647 (O_4647,N_49606,N_49547);
and UO_4648 (O_4648,N_49561,N_49652);
and UO_4649 (O_4649,N_49534,N_49916);
xor UO_4650 (O_4650,N_49600,N_49544);
nor UO_4651 (O_4651,N_49578,N_49902);
or UO_4652 (O_4652,N_49899,N_49748);
and UO_4653 (O_4653,N_49946,N_49910);
nand UO_4654 (O_4654,N_49856,N_49780);
and UO_4655 (O_4655,N_49719,N_49536);
nor UO_4656 (O_4656,N_49678,N_49537);
nor UO_4657 (O_4657,N_49577,N_49838);
nand UO_4658 (O_4658,N_49554,N_49981);
nor UO_4659 (O_4659,N_49649,N_49627);
xor UO_4660 (O_4660,N_49950,N_49961);
or UO_4661 (O_4661,N_49939,N_49789);
nand UO_4662 (O_4662,N_49973,N_49555);
or UO_4663 (O_4663,N_49945,N_49554);
nand UO_4664 (O_4664,N_49785,N_49849);
nor UO_4665 (O_4665,N_49726,N_49793);
xnor UO_4666 (O_4666,N_49641,N_49765);
nand UO_4667 (O_4667,N_49983,N_49981);
or UO_4668 (O_4668,N_49839,N_49658);
nor UO_4669 (O_4669,N_49536,N_49919);
and UO_4670 (O_4670,N_49542,N_49578);
nor UO_4671 (O_4671,N_49757,N_49897);
and UO_4672 (O_4672,N_49805,N_49925);
nor UO_4673 (O_4673,N_49715,N_49824);
xor UO_4674 (O_4674,N_49959,N_49671);
and UO_4675 (O_4675,N_49858,N_49551);
nor UO_4676 (O_4676,N_49586,N_49795);
and UO_4677 (O_4677,N_49832,N_49815);
and UO_4678 (O_4678,N_49504,N_49984);
xor UO_4679 (O_4679,N_49981,N_49944);
nand UO_4680 (O_4680,N_49692,N_49986);
nand UO_4681 (O_4681,N_49941,N_49990);
nor UO_4682 (O_4682,N_49515,N_49973);
xnor UO_4683 (O_4683,N_49501,N_49910);
or UO_4684 (O_4684,N_49927,N_49746);
nor UO_4685 (O_4685,N_49926,N_49584);
xnor UO_4686 (O_4686,N_49632,N_49531);
xor UO_4687 (O_4687,N_49970,N_49674);
or UO_4688 (O_4688,N_49754,N_49916);
xnor UO_4689 (O_4689,N_49884,N_49641);
nor UO_4690 (O_4690,N_49985,N_49652);
or UO_4691 (O_4691,N_49536,N_49913);
xnor UO_4692 (O_4692,N_49934,N_49700);
nor UO_4693 (O_4693,N_49696,N_49999);
nand UO_4694 (O_4694,N_49988,N_49638);
nor UO_4695 (O_4695,N_49548,N_49772);
nand UO_4696 (O_4696,N_49860,N_49759);
nor UO_4697 (O_4697,N_49613,N_49888);
xor UO_4698 (O_4698,N_49701,N_49554);
xor UO_4699 (O_4699,N_49551,N_49744);
or UO_4700 (O_4700,N_49953,N_49699);
or UO_4701 (O_4701,N_49678,N_49770);
nand UO_4702 (O_4702,N_49514,N_49850);
or UO_4703 (O_4703,N_49877,N_49607);
and UO_4704 (O_4704,N_49514,N_49900);
and UO_4705 (O_4705,N_49558,N_49507);
or UO_4706 (O_4706,N_49553,N_49740);
and UO_4707 (O_4707,N_49987,N_49838);
nand UO_4708 (O_4708,N_49580,N_49780);
and UO_4709 (O_4709,N_49611,N_49579);
xnor UO_4710 (O_4710,N_49778,N_49514);
nor UO_4711 (O_4711,N_49821,N_49566);
and UO_4712 (O_4712,N_49603,N_49928);
xor UO_4713 (O_4713,N_49580,N_49582);
and UO_4714 (O_4714,N_49779,N_49539);
and UO_4715 (O_4715,N_49924,N_49682);
and UO_4716 (O_4716,N_49566,N_49700);
and UO_4717 (O_4717,N_49657,N_49664);
or UO_4718 (O_4718,N_49716,N_49744);
nand UO_4719 (O_4719,N_49688,N_49725);
nor UO_4720 (O_4720,N_49673,N_49826);
or UO_4721 (O_4721,N_49835,N_49979);
xor UO_4722 (O_4722,N_49704,N_49900);
nand UO_4723 (O_4723,N_49665,N_49743);
and UO_4724 (O_4724,N_49949,N_49988);
nand UO_4725 (O_4725,N_49825,N_49567);
or UO_4726 (O_4726,N_49886,N_49511);
or UO_4727 (O_4727,N_49505,N_49984);
nand UO_4728 (O_4728,N_49721,N_49797);
xor UO_4729 (O_4729,N_49537,N_49593);
xor UO_4730 (O_4730,N_49754,N_49845);
xnor UO_4731 (O_4731,N_49521,N_49616);
and UO_4732 (O_4732,N_49748,N_49895);
or UO_4733 (O_4733,N_49894,N_49739);
nand UO_4734 (O_4734,N_49870,N_49642);
and UO_4735 (O_4735,N_49543,N_49640);
nand UO_4736 (O_4736,N_49529,N_49703);
or UO_4737 (O_4737,N_49884,N_49879);
xnor UO_4738 (O_4738,N_49613,N_49706);
nor UO_4739 (O_4739,N_49849,N_49968);
or UO_4740 (O_4740,N_49515,N_49614);
or UO_4741 (O_4741,N_49914,N_49713);
nor UO_4742 (O_4742,N_49554,N_49668);
nand UO_4743 (O_4743,N_49915,N_49796);
and UO_4744 (O_4744,N_49635,N_49615);
xnor UO_4745 (O_4745,N_49835,N_49639);
nor UO_4746 (O_4746,N_49690,N_49664);
or UO_4747 (O_4747,N_49812,N_49510);
xnor UO_4748 (O_4748,N_49878,N_49584);
nand UO_4749 (O_4749,N_49991,N_49679);
nand UO_4750 (O_4750,N_49678,N_49750);
and UO_4751 (O_4751,N_49560,N_49866);
nand UO_4752 (O_4752,N_49763,N_49833);
or UO_4753 (O_4753,N_49553,N_49753);
and UO_4754 (O_4754,N_49839,N_49900);
xor UO_4755 (O_4755,N_49957,N_49820);
and UO_4756 (O_4756,N_49651,N_49681);
nand UO_4757 (O_4757,N_49895,N_49808);
or UO_4758 (O_4758,N_49952,N_49875);
or UO_4759 (O_4759,N_49621,N_49959);
nand UO_4760 (O_4760,N_49680,N_49591);
nor UO_4761 (O_4761,N_49854,N_49959);
xnor UO_4762 (O_4762,N_49612,N_49813);
nor UO_4763 (O_4763,N_49798,N_49925);
and UO_4764 (O_4764,N_49812,N_49540);
or UO_4765 (O_4765,N_49976,N_49918);
and UO_4766 (O_4766,N_49514,N_49880);
or UO_4767 (O_4767,N_49891,N_49919);
nand UO_4768 (O_4768,N_49991,N_49792);
and UO_4769 (O_4769,N_49958,N_49548);
and UO_4770 (O_4770,N_49578,N_49584);
xor UO_4771 (O_4771,N_49821,N_49764);
and UO_4772 (O_4772,N_49793,N_49685);
xor UO_4773 (O_4773,N_49841,N_49695);
and UO_4774 (O_4774,N_49662,N_49661);
nor UO_4775 (O_4775,N_49508,N_49966);
xnor UO_4776 (O_4776,N_49866,N_49507);
nor UO_4777 (O_4777,N_49897,N_49992);
and UO_4778 (O_4778,N_49986,N_49577);
and UO_4779 (O_4779,N_49536,N_49924);
or UO_4780 (O_4780,N_49996,N_49718);
xnor UO_4781 (O_4781,N_49512,N_49692);
nand UO_4782 (O_4782,N_49641,N_49519);
or UO_4783 (O_4783,N_49883,N_49935);
nor UO_4784 (O_4784,N_49690,N_49533);
or UO_4785 (O_4785,N_49803,N_49783);
and UO_4786 (O_4786,N_49956,N_49520);
or UO_4787 (O_4787,N_49872,N_49741);
xnor UO_4788 (O_4788,N_49581,N_49766);
and UO_4789 (O_4789,N_49561,N_49670);
and UO_4790 (O_4790,N_49786,N_49807);
and UO_4791 (O_4791,N_49563,N_49640);
and UO_4792 (O_4792,N_49745,N_49974);
nand UO_4793 (O_4793,N_49710,N_49678);
nand UO_4794 (O_4794,N_49945,N_49701);
nor UO_4795 (O_4795,N_49595,N_49513);
nor UO_4796 (O_4796,N_49572,N_49887);
nand UO_4797 (O_4797,N_49755,N_49902);
nor UO_4798 (O_4798,N_49768,N_49594);
xnor UO_4799 (O_4799,N_49961,N_49847);
xnor UO_4800 (O_4800,N_49517,N_49942);
nand UO_4801 (O_4801,N_49672,N_49545);
and UO_4802 (O_4802,N_49930,N_49800);
or UO_4803 (O_4803,N_49676,N_49750);
xnor UO_4804 (O_4804,N_49659,N_49889);
and UO_4805 (O_4805,N_49557,N_49819);
nor UO_4806 (O_4806,N_49955,N_49844);
nor UO_4807 (O_4807,N_49732,N_49519);
xor UO_4808 (O_4808,N_49810,N_49877);
nor UO_4809 (O_4809,N_49535,N_49805);
nand UO_4810 (O_4810,N_49531,N_49963);
nor UO_4811 (O_4811,N_49735,N_49941);
or UO_4812 (O_4812,N_49587,N_49809);
or UO_4813 (O_4813,N_49592,N_49844);
or UO_4814 (O_4814,N_49656,N_49695);
nand UO_4815 (O_4815,N_49765,N_49512);
nand UO_4816 (O_4816,N_49621,N_49929);
or UO_4817 (O_4817,N_49834,N_49974);
nand UO_4818 (O_4818,N_49782,N_49948);
xnor UO_4819 (O_4819,N_49562,N_49606);
nand UO_4820 (O_4820,N_49581,N_49847);
and UO_4821 (O_4821,N_49535,N_49823);
nand UO_4822 (O_4822,N_49710,N_49902);
and UO_4823 (O_4823,N_49882,N_49816);
nor UO_4824 (O_4824,N_49798,N_49835);
and UO_4825 (O_4825,N_49629,N_49589);
xnor UO_4826 (O_4826,N_49876,N_49839);
and UO_4827 (O_4827,N_49654,N_49961);
nand UO_4828 (O_4828,N_49896,N_49628);
nor UO_4829 (O_4829,N_49880,N_49812);
and UO_4830 (O_4830,N_49548,N_49749);
nand UO_4831 (O_4831,N_49665,N_49660);
nand UO_4832 (O_4832,N_49989,N_49761);
xnor UO_4833 (O_4833,N_49906,N_49893);
nor UO_4834 (O_4834,N_49745,N_49747);
or UO_4835 (O_4835,N_49989,N_49711);
xor UO_4836 (O_4836,N_49525,N_49599);
or UO_4837 (O_4837,N_49941,N_49877);
nor UO_4838 (O_4838,N_49587,N_49511);
nand UO_4839 (O_4839,N_49527,N_49783);
nand UO_4840 (O_4840,N_49965,N_49849);
nand UO_4841 (O_4841,N_49912,N_49806);
nor UO_4842 (O_4842,N_49623,N_49661);
nand UO_4843 (O_4843,N_49910,N_49669);
or UO_4844 (O_4844,N_49835,N_49758);
or UO_4845 (O_4845,N_49850,N_49765);
xnor UO_4846 (O_4846,N_49885,N_49557);
nand UO_4847 (O_4847,N_49536,N_49589);
or UO_4848 (O_4848,N_49690,N_49691);
nor UO_4849 (O_4849,N_49555,N_49853);
nand UO_4850 (O_4850,N_49640,N_49991);
nand UO_4851 (O_4851,N_49685,N_49500);
nor UO_4852 (O_4852,N_49979,N_49671);
nand UO_4853 (O_4853,N_49510,N_49722);
xor UO_4854 (O_4854,N_49894,N_49544);
nor UO_4855 (O_4855,N_49668,N_49528);
nor UO_4856 (O_4856,N_49841,N_49643);
or UO_4857 (O_4857,N_49864,N_49752);
xor UO_4858 (O_4858,N_49855,N_49821);
nor UO_4859 (O_4859,N_49742,N_49515);
xnor UO_4860 (O_4860,N_49994,N_49905);
nor UO_4861 (O_4861,N_49621,N_49924);
nor UO_4862 (O_4862,N_49614,N_49990);
and UO_4863 (O_4863,N_49850,N_49830);
nand UO_4864 (O_4864,N_49736,N_49800);
and UO_4865 (O_4865,N_49628,N_49649);
xnor UO_4866 (O_4866,N_49989,N_49844);
and UO_4867 (O_4867,N_49841,N_49704);
xnor UO_4868 (O_4868,N_49893,N_49580);
nor UO_4869 (O_4869,N_49986,N_49545);
or UO_4870 (O_4870,N_49836,N_49866);
xor UO_4871 (O_4871,N_49641,N_49985);
nand UO_4872 (O_4872,N_49798,N_49769);
or UO_4873 (O_4873,N_49656,N_49804);
or UO_4874 (O_4874,N_49855,N_49612);
or UO_4875 (O_4875,N_49514,N_49725);
xor UO_4876 (O_4876,N_49570,N_49573);
and UO_4877 (O_4877,N_49624,N_49706);
nand UO_4878 (O_4878,N_49785,N_49627);
nor UO_4879 (O_4879,N_49615,N_49846);
nor UO_4880 (O_4880,N_49609,N_49949);
xnor UO_4881 (O_4881,N_49625,N_49896);
and UO_4882 (O_4882,N_49911,N_49797);
and UO_4883 (O_4883,N_49738,N_49871);
nand UO_4884 (O_4884,N_49973,N_49782);
and UO_4885 (O_4885,N_49578,N_49899);
or UO_4886 (O_4886,N_49823,N_49933);
and UO_4887 (O_4887,N_49645,N_49734);
nor UO_4888 (O_4888,N_49861,N_49935);
nor UO_4889 (O_4889,N_49855,N_49988);
xor UO_4890 (O_4890,N_49503,N_49832);
nor UO_4891 (O_4891,N_49595,N_49898);
nand UO_4892 (O_4892,N_49779,N_49727);
xor UO_4893 (O_4893,N_49896,N_49891);
or UO_4894 (O_4894,N_49778,N_49753);
xor UO_4895 (O_4895,N_49528,N_49563);
nand UO_4896 (O_4896,N_49815,N_49613);
or UO_4897 (O_4897,N_49642,N_49753);
nor UO_4898 (O_4898,N_49633,N_49609);
xor UO_4899 (O_4899,N_49775,N_49569);
nand UO_4900 (O_4900,N_49548,N_49539);
and UO_4901 (O_4901,N_49974,N_49988);
nand UO_4902 (O_4902,N_49707,N_49999);
or UO_4903 (O_4903,N_49642,N_49706);
nand UO_4904 (O_4904,N_49510,N_49734);
nand UO_4905 (O_4905,N_49753,N_49766);
and UO_4906 (O_4906,N_49868,N_49608);
nand UO_4907 (O_4907,N_49996,N_49853);
or UO_4908 (O_4908,N_49513,N_49860);
and UO_4909 (O_4909,N_49542,N_49677);
xor UO_4910 (O_4910,N_49811,N_49529);
and UO_4911 (O_4911,N_49693,N_49545);
nor UO_4912 (O_4912,N_49784,N_49548);
and UO_4913 (O_4913,N_49943,N_49800);
nand UO_4914 (O_4914,N_49636,N_49978);
or UO_4915 (O_4915,N_49777,N_49502);
nor UO_4916 (O_4916,N_49629,N_49730);
xnor UO_4917 (O_4917,N_49532,N_49852);
or UO_4918 (O_4918,N_49966,N_49505);
nor UO_4919 (O_4919,N_49652,N_49993);
xnor UO_4920 (O_4920,N_49864,N_49629);
nor UO_4921 (O_4921,N_49998,N_49593);
and UO_4922 (O_4922,N_49693,N_49792);
xnor UO_4923 (O_4923,N_49746,N_49564);
nand UO_4924 (O_4924,N_49559,N_49892);
nand UO_4925 (O_4925,N_49625,N_49822);
or UO_4926 (O_4926,N_49974,N_49778);
nand UO_4927 (O_4927,N_49638,N_49647);
xnor UO_4928 (O_4928,N_49917,N_49774);
nor UO_4929 (O_4929,N_49589,N_49849);
and UO_4930 (O_4930,N_49521,N_49949);
nand UO_4931 (O_4931,N_49568,N_49941);
nor UO_4932 (O_4932,N_49742,N_49815);
xor UO_4933 (O_4933,N_49681,N_49599);
nand UO_4934 (O_4934,N_49956,N_49536);
or UO_4935 (O_4935,N_49771,N_49601);
and UO_4936 (O_4936,N_49721,N_49739);
and UO_4937 (O_4937,N_49665,N_49971);
nor UO_4938 (O_4938,N_49829,N_49995);
xnor UO_4939 (O_4939,N_49878,N_49614);
nand UO_4940 (O_4940,N_49606,N_49949);
nand UO_4941 (O_4941,N_49760,N_49855);
nand UO_4942 (O_4942,N_49718,N_49783);
or UO_4943 (O_4943,N_49910,N_49699);
nand UO_4944 (O_4944,N_49924,N_49501);
xor UO_4945 (O_4945,N_49786,N_49601);
nor UO_4946 (O_4946,N_49824,N_49786);
nor UO_4947 (O_4947,N_49759,N_49984);
xor UO_4948 (O_4948,N_49986,N_49727);
xor UO_4949 (O_4949,N_49665,N_49616);
and UO_4950 (O_4950,N_49678,N_49541);
and UO_4951 (O_4951,N_49850,N_49856);
or UO_4952 (O_4952,N_49810,N_49766);
nor UO_4953 (O_4953,N_49916,N_49583);
xor UO_4954 (O_4954,N_49666,N_49564);
or UO_4955 (O_4955,N_49560,N_49896);
and UO_4956 (O_4956,N_49920,N_49608);
xor UO_4957 (O_4957,N_49697,N_49672);
and UO_4958 (O_4958,N_49623,N_49871);
or UO_4959 (O_4959,N_49794,N_49872);
nand UO_4960 (O_4960,N_49537,N_49972);
nand UO_4961 (O_4961,N_49778,N_49701);
nand UO_4962 (O_4962,N_49674,N_49730);
nor UO_4963 (O_4963,N_49646,N_49930);
xor UO_4964 (O_4964,N_49832,N_49574);
xor UO_4965 (O_4965,N_49728,N_49797);
nand UO_4966 (O_4966,N_49792,N_49572);
or UO_4967 (O_4967,N_49784,N_49720);
and UO_4968 (O_4968,N_49541,N_49867);
xor UO_4969 (O_4969,N_49822,N_49971);
nor UO_4970 (O_4970,N_49651,N_49691);
xor UO_4971 (O_4971,N_49774,N_49823);
nand UO_4972 (O_4972,N_49791,N_49686);
nand UO_4973 (O_4973,N_49899,N_49745);
nor UO_4974 (O_4974,N_49680,N_49578);
or UO_4975 (O_4975,N_49522,N_49978);
or UO_4976 (O_4976,N_49889,N_49761);
nor UO_4977 (O_4977,N_49959,N_49806);
or UO_4978 (O_4978,N_49837,N_49627);
or UO_4979 (O_4979,N_49510,N_49726);
nand UO_4980 (O_4980,N_49817,N_49608);
nor UO_4981 (O_4981,N_49536,N_49591);
nor UO_4982 (O_4982,N_49794,N_49852);
nor UO_4983 (O_4983,N_49672,N_49772);
and UO_4984 (O_4984,N_49513,N_49885);
and UO_4985 (O_4985,N_49684,N_49543);
or UO_4986 (O_4986,N_49784,N_49967);
xor UO_4987 (O_4987,N_49562,N_49735);
nor UO_4988 (O_4988,N_49661,N_49557);
and UO_4989 (O_4989,N_49854,N_49913);
or UO_4990 (O_4990,N_49747,N_49588);
xor UO_4991 (O_4991,N_49877,N_49999);
xor UO_4992 (O_4992,N_49860,N_49997);
or UO_4993 (O_4993,N_49589,N_49617);
and UO_4994 (O_4994,N_49589,N_49787);
nor UO_4995 (O_4995,N_49630,N_49584);
xor UO_4996 (O_4996,N_49926,N_49586);
xnor UO_4997 (O_4997,N_49977,N_49587);
and UO_4998 (O_4998,N_49900,N_49723);
nor UO_4999 (O_4999,N_49609,N_49973);
endmodule